module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 ,
    pi131 , pi132 , pi133 , pi134 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 ,
    pi130 , pi131 , pi132 , pi133 , pi134 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ;
  wire n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018,
    n1019, n1020, n1021, n1022, n1023, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108,
    n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411,
    n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441,
    n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471,
    n1472, n1473, n1474, n1475, n1476, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1624,
    n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642,
    n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654,
    n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672,
    n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721,
    n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751,
    n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782,
    n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812,
    n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1843,
    n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861,
    n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873,
    n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2062,
    n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086,
    n2087, n2088, n2089, n2090, n2091, n2092,
    n2093, n2094, n2095, n2096, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122,
    n2123, n2124, n2125, n2126, n2127, n2128,
    n2129, n2130, n2131, n2132, n2133, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141,
    n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153,
    n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183,
    n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2225, n2226, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233,
    n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2276, n2277, n2278,
    n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303,
    n2304, n2305, n2306, n2307, n2308, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341,
    n2342, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386,
    n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2395, n2396, n2397, n2398, n2399,
    n2400, n2401, n2402, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424,
    n2425, n2426, n2427, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2480, n2481, n2482,
    n2483, n2484, n2485, n2486, n2487, n2488,
    n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2497, n2498, n2499, n2500, n2501,
    n2502, n2503, n2504, n2505, n2506, n2507,
    n2508, n2509, n2510, n2511, n2512, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2582, n2583, n2584,
    n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596,
    n2597, n2599, n2600, n2601, n2602, n2603,
    n2604, n2605, n2606, n2607, n2608, n2609,
    n2610, n2611, n2612, n2613, n2614, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641,
    n2642, n2643, n2644, n2645, n2646, n2647,
    n2648, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2684, n2685, n2686,
    n2687, n2688, n2689, n2690, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2701, n2702, n2703, n2704, n2705,
    n2706, n2707, n2708, n2709, n2710, n2711,
    n2712, n2713, n2714, n2715, n2716, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2735, n2736, n2737,
    n2738, n2739, n2740, n2741, n2742, n2743,
    n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794,
    n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2803, n2804, n2805, n2806, n2807,
    n2808, n2809, n2810, n2811, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851,
    n2852, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896,
    n2897, n2898, n2899, n2900, n2901, n2902,
    n2903, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915,
    n2916, n2917, n2918, n2919, n2920, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2939, n2940, n2941,
    n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953,
    n2954, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2997, n2998,
    n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3007, n3008, n3009, n3010, n3011,
    n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3024,
    n3025, n3027, n3028, n3030, n3031, n3033,
    n3034, n3036, n3037, n3039, n3040, n3042,
    n3043, n3045, n3046, n3048, n3049, n3051,
    n3052, n3054, n3055, n3057, n3058, n3060,
    n3061, n3063, n3064, n3066, n3067, n3069,
    n3070, n3072, n3073, n3075, n3076, n3078,
    n3079, n3081, n3082, n3084, n3085, n3087,
    n3088, n3090, n3091, n3093, n3094, n3096,
    n3097, n3099, n3100, n3102, n3103, n3105,
    n3106, n3108, n3109, n3111, n3112, n3114,
    n3115, n3117, n3118, n3120, n3121, n3123,
    n3124, n3126, n3127, n3129, n3130, n3132,
    n3133, n3135, n3136, n3138, n3139, n3141,
    n3142, n3144, n3145, n3147, n3148, n3150,
    n3151, n3153, n3154, n3156, n3157, n3159,
    n3160, n3162, n3163, n3165, n3166, n3168,
    n3169, n3171, n3172, n3174, n3175, n3177,
    n3178, n3180, n3181, n3183, n3184, n3186,
    n3187, n3189, n3190, n3192, n3193, n3195,
    n3196, n3198, n3199, n3201, n3202, n3204,
    n3205, n3207, n3208, n3210, n3211, n3213,
    n3214;
  assign n264 = ~pi132  & pi133 ;
  assign n265 = pi130  & ~pi131 ;
  assign n266 = pi89  & pi128 ;
  assign n267 = pi90  & ~pi128 ;
  assign n268 = ~n266 & ~n267;
  assign n269 = pi129  & ~n268;
  assign n270 = pi92  & ~pi128 ;
  assign n271 = pi91  & pi128 ;
  assign n272 = ~n270 & ~n271;
  assign n273 = ~pi129  & ~n272;
  assign n274 = ~n269 & ~n273;
  assign n275 = n265 & ~n274;
  assign n276 = ~pi130  & pi131 ;
  assign n277 = pi85  & pi128 ;
  assign n278 = pi86  & ~pi128 ;
  assign n279 = ~n277 & ~n278;
  assign n280 = pi129  & ~n279;
  assign n281 = pi88  & ~pi128 ;
  assign n282 = pi87  & pi128 ;
  assign n283 = ~n281 & ~n282;
  assign n284 = ~pi129  & ~n283;
  assign n285 = ~n280 & ~n284;
  assign n286 = n276 & ~n285;
  assign n287 = ~pi130  & ~pi131 ;
  assign n288 = pi93  & pi128 ;
  assign n289 = pi94  & ~pi128 ;
  assign n290 = ~n288 & ~n289;
  assign n291 = pi129  & ~n290;
  assign n292 = pi96  & ~pi128 ;
  assign n293 = pi95  & pi128 ;
  assign n294 = ~n292 & ~n293;
  assign n295 = ~pi129  & ~n294;
  assign n296 = ~n291 & ~n295;
  assign n297 = n287 & ~n296;
  assign n298 = pi130  & pi131 ;
  assign n299 = pi81  & pi128 ;
  assign n300 = pi82  & ~pi128 ;
  assign n301 = ~n299 & ~n300;
  assign n302 = pi129  & ~n301;
  assign n303 = pi84  & ~pi128 ;
  assign n304 = pi83  & pi128 ;
  assign n305 = ~n303 & ~n304;
  assign n306 = ~pi129  & ~n305;
  assign n307 = ~n302 & ~n306;
  assign n308 = n298 & ~n307;
  assign n309 = ~n297 & ~n308;
  assign n310 = ~n286 & n309;
  assign n311 = ~n275 & n310;
  assign n312 = n264 & ~n311;
  assign n313 = pi132  & ~pi133 ;
  assign n314 = pi105  & pi128 ;
  assign n315 = pi106  & ~pi128 ;
  assign n316 = ~n314 & ~n315;
  assign n317 = pi129  & ~n316;
  assign n318 = pi108  & ~pi128 ;
  assign n319 = pi107  & pi128 ;
  assign n320 = ~n318 & ~n319;
  assign n321 = ~pi129  & ~n320;
  assign n322 = ~n317 & ~n321;
  assign n323 = n265 & ~n322;
  assign n324 = pi101  & pi128 ;
  assign n325 = pi102  & ~pi128 ;
  assign n326 = ~n324 & ~n325;
  assign n327 = pi129  & ~n326;
  assign n328 = pi104  & ~pi128 ;
  assign n329 = pi103  & pi128 ;
  assign n330 = ~n328 & ~n329;
  assign n331 = ~pi129  & ~n330;
  assign n332 = ~n327 & ~n331;
  assign n333 = n276 & ~n332;
  assign n334 = pi109  & pi128 ;
  assign n335 = pi110  & ~pi128 ;
  assign n336 = ~n334 & ~n335;
  assign n337 = pi129  & ~n336;
  assign n338 = pi112  & ~pi128 ;
  assign n339 = pi111  & pi128 ;
  assign n340 = ~n338 & ~n339;
  assign n341 = ~pi129  & ~n340;
  assign n342 = ~n337 & ~n341;
  assign n343 = n287 & ~n342;
  assign n344 = pi97  & pi128 ;
  assign n345 = pi98  & ~pi128 ;
  assign n346 = ~n344 & ~n345;
  assign n347 = pi129  & ~n346;
  assign n348 = pi100  & ~pi128 ;
  assign n349 = pi99  & pi128 ;
  assign n350 = ~n348 & ~n349;
  assign n351 = ~pi129  & ~n350;
  assign n352 = ~n347 & ~n351;
  assign n353 = n298 & ~n352;
  assign n354 = ~n343 & ~n353;
  assign n355 = ~n333 & n354;
  assign n356 = ~n323 & n355;
  assign n357 = n313 & ~n356;
  assign n358 = pi132  & pi133 ;
  assign n359 = pi73  & pi128 ;
  assign n360 = pi74  & ~pi128 ;
  assign n361 = ~n359 & ~n360;
  assign n362 = pi129  & ~n361;
  assign n363 = pi76  & ~pi128 ;
  assign n364 = pi75  & pi128 ;
  assign n365 = ~n363 & ~n364;
  assign n366 = ~pi129  & ~n365;
  assign n367 = ~n362 & ~n366;
  assign n368 = n265 & ~n367;
  assign n369 = pi69  & pi128 ;
  assign n370 = pi70  & ~pi128 ;
  assign n371 = ~n369 & ~n370;
  assign n372 = pi129  & ~n371;
  assign n373 = pi72  & ~pi128 ;
  assign n374 = pi71  & pi128 ;
  assign n375 = ~n373 & ~n374;
  assign n376 = ~pi129  & ~n375;
  assign n377 = ~n372 & ~n376;
  assign n378 = n276 & ~n377;
  assign n379 = pi77  & pi128 ;
  assign n380 = pi78  & ~pi128 ;
  assign n381 = ~n379 & ~n380;
  assign n382 = pi129  & ~n381;
  assign n383 = pi80  & ~pi128 ;
  assign n384 = pi79  & pi128 ;
  assign n385 = ~n383 & ~n384;
  assign n386 = ~pi129  & ~n385;
  assign n387 = ~n382 & ~n386;
  assign n388 = n287 & ~n387;
  assign n389 = pi65  & pi128 ;
  assign n390 = pi66  & ~pi128 ;
  assign n391 = ~n389 & ~n390;
  assign n392 = pi129  & ~n391;
  assign n393 = pi68  & ~pi128 ;
  assign n394 = pi67  & pi128 ;
  assign n395 = ~n393 & ~n394;
  assign n396 = ~pi129  & ~n395;
  assign n397 = ~n392 & ~n396;
  assign n398 = n298 & ~n397;
  assign n399 = ~n388 & ~n398;
  assign n400 = ~n378 & n399;
  assign n401 = ~n368 & n400;
  assign n402 = n358 & ~n401;
  assign n403 = ~pi132  & ~pi133 ;
  assign n404 = pi121  & pi128 ;
  assign n405 = pi122  & ~pi128 ;
  assign n406 = ~n404 & ~n405;
  assign n407 = pi129  & ~n406;
  assign n408 = pi124  & ~pi128 ;
  assign n409 = pi123  & pi128 ;
  assign n410 = ~n408 & ~n409;
  assign n411 = ~pi129  & ~n410;
  assign n412 = ~n407 & ~n411;
  assign n413 = n265 & ~n412;
  assign n414 = pi117  & pi128 ;
  assign n415 = pi118  & ~pi128 ;
  assign n416 = ~n414 & ~n415;
  assign n417 = pi129  & ~n416;
  assign n418 = pi120  & ~pi128 ;
  assign n419 = pi119  & pi128 ;
  assign n420 = ~n418 & ~n419;
  assign n421 = ~pi129  & ~n420;
  assign n422 = ~n417 & ~n421;
  assign n423 = n276 & ~n422;
  assign n424 = pi125  & pi128 ;
  assign n425 = pi126  & ~pi128 ;
  assign n426 = ~n424 & ~n425;
  assign n427 = pi129  & ~n426;
  assign n428 = pi0  & ~pi128 ;
  assign n429 = pi127  & pi128 ;
  assign n430 = ~n428 & ~n429;
  assign n431 = ~pi129  & ~n430;
  assign n432 = ~n427 & ~n431;
  assign n433 = n287 & ~n432;
  assign n434 = pi113  & pi128 ;
  assign n435 = pi114  & ~pi128 ;
  assign n436 = ~n434 & ~n435;
  assign n437 = pi129  & ~n436;
  assign n438 = pi116  & ~pi128 ;
  assign n439 = pi115  & pi128 ;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~pi129  & ~n440;
  assign n442 = ~n437 & ~n441;
  assign n443 = n298 & ~n442;
  assign n444 = ~n433 & ~n443;
  assign n445 = ~n423 & n444;
  assign n446 = ~n413 & n445;
  assign n447 = n403 & ~n446;
  assign n448 = ~n402 & ~n447;
  assign n449 = ~n357 & n448;
  assign n450 = ~n312 & n449;
  assign n451 = ~pi134  & ~n450;
  assign n452 = pi25  & pi128 ;
  assign n453 = pi26  & ~pi128 ;
  assign n454 = ~n452 & ~n453;
  assign n455 = pi129  & ~n454;
  assign n456 = pi28  & ~pi128 ;
  assign n457 = pi27  & pi128 ;
  assign n458 = ~n456 & ~n457;
  assign n459 = ~pi129  & ~n458;
  assign n460 = ~n455 & ~n459;
  assign n461 = n265 & ~n460;
  assign n462 = pi21  & pi128 ;
  assign n463 = pi22  & ~pi128 ;
  assign n464 = ~n462 & ~n463;
  assign n465 = pi129  & ~n464;
  assign n466 = pi24  & ~pi128 ;
  assign n467 = pi23  & pi128 ;
  assign n468 = ~n466 & ~n467;
  assign n469 = ~pi129  & ~n468;
  assign n470 = ~n465 & ~n469;
  assign n471 = n276 & ~n470;
  assign n472 = pi29  & pi128 ;
  assign n473 = pi30  & ~pi128 ;
  assign n474 = ~n472 & ~n473;
  assign n475 = pi129  & ~n474;
  assign n476 = pi32  & ~pi128 ;
  assign n477 = pi31  & pi128 ;
  assign n478 = ~n476 & ~n477;
  assign n479 = ~pi129  & ~n478;
  assign n480 = ~n475 & ~n479;
  assign n481 = n287 & ~n480;
  assign n482 = pi17  & pi128 ;
  assign n483 = pi18  & ~pi128 ;
  assign n484 = ~n482 & ~n483;
  assign n485 = pi129  & ~n484;
  assign n486 = pi20  & ~pi128 ;
  assign n487 = pi19  & pi128 ;
  assign n488 = ~n486 & ~n487;
  assign n489 = ~pi129  & ~n488;
  assign n490 = ~n485 & ~n489;
  assign n491 = n298 & ~n490;
  assign n492 = ~n481 & ~n491;
  assign n493 = ~n471 & n492;
  assign n494 = ~n461 & n493;
  assign n495 = n264 & ~n494;
  assign n496 = pi41  & pi128 ;
  assign n497 = pi42  & ~pi128 ;
  assign n498 = ~n496 & ~n497;
  assign n499 = pi129  & ~n498;
  assign n500 = pi44  & ~pi128 ;
  assign n501 = pi43  & pi128 ;
  assign n502 = ~n500 & ~n501;
  assign n503 = ~pi129  & ~n502;
  assign n504 = ~n499 & ~n503;
  assign n505 = n265 & ~n504;
  assign n506 = pi40  & ~pi128 ;
  assign n507 = pi39  & pi128 ;
  assign n508 = ~n506 & ~n507;
  assign n509 = ~pi129  & ~n508;
  assign n510 = pi37  & pi128 ;
  assign n511 = pi38  & ~pi128 ;
  assign n512 = ~n510 & ~n511;
  assign n513 = pi129  & ~n512;
  assign n514 = ~n509 & ~n513;
  assign n515 = n276 & ~n514;
  assign n516 = pi45  & pi128 ;
  assign n517 = pi46  & ~pi128 ;
  assign n518 = ~n516 & ~n517;
  assign n519 = pi129  & ~n518;
  assign n520 = pi48  & ~pi128 ;
  assign n521 = pi47  & pi128 ;
  assign n522 = ~n520 & ~n521;
  assign n523 = ~pi129  & ~n522;
  assign n524 = ~n519 & ~n523;
  assign n525 = n287 & ~n524;
  assign n526 = pi33  & pi128 ;
  assign n527 = pi34  & ~pi128 ;
  assign n528 = ~n526 & ~n527;
  assign n529 = pi129  & ~n528;
  assign n530 = pi36  & ~pi128 ;
  assign n531 = pi35  & pi128 ;
  assign n532 = ~n530 & ~n531;
  assign n533 = ~pi129  & ~n532;
  assign n534 = ~n529 & ~n533;
  assign n535 = n298 & ~n534;
  assign n536 = ~n525 & ~n535;
  assign n537 = ~n515 & n536;
  assign n538 = ~n505 & n537;
  assign n539 = n313 & ~n538;
  assign n540 = pi9  & pi128 ;
  assign n541 = pi10  & ~pi128 ;
  assign n542 = ~n540 & ~n541;
  assign n543 = pi129  & ~n542;
  assign n544 = pi12  & ~pi128 ;
  assign n545 = pi11  & pi128 ;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~pi129  & ~n546;
  assign n548 = ~n543 & ~n547;
  assign n549 = n265 & ~n548;
  assign n550 = pi5  & pi128 ;
  assign n551 = pi6  & ~pi128 ;
  assign n552 = ~n550 & ~n551;
  assign n553 = pi129  & ~n552;
  assign n554 = pi8  & ~pi128 ;
  assign n555 = pi7  & pi128 ;
  assign n556 = ~n554 & ~n555;
  assign n557 = ~pi129  & ~n556;
  assign n558 = ~n553 & ~n557;
  assign n559 = n276 & ~n558;
  assign n560 = pi13  & pi128 ;
  assign n561 = pi14  & ~pi128 ;
  assign n562 = ~n560 & ~n561;
  assign n563 = pi129  & ~n562;
  assign n564 = pi16  & ~pi128 ;
  assign n565 = pi15  & pi128 ;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~pi129  & ~n566;
  assign n568 = ~n563 & ~n567;
  assign n569 = n287 & ~n568;
  assign n570 = pi1  & pi128 ;
  assign n571 = pi2  & ~pi128 ;
  assign n572 = ~n570 & ~n571;
  assign n573 = pi129  & ~n572;
  assign n574 = pi4  & ~pi128 ;
  assign n575 = pi3  & pi128 ;
  assign n576 = ~n574 & ~n575;
  assign n577 = ~pi129  & ~n576;
  assign n578 = ~n573 & ~n577;
  assign n579 = n298 & ~n578;
  assign n580 = ~n569 & ~n579;
  assign n581 = ~n559 & n580;
  assign n582 = ~n549 & n581;
  assign n583 = n358 & ~n582;
  assign n584 = pi57  & pi128 ;
  assign n585 = pi58  & ~pi128 ;
  assign n586 = ~n584 & ~n585;
  assign n587 = pi129  & ~n586;
  assign n588 = pi60  & ~pi128 ;
  assign n589 = pi59  & pi128 ;
  assign n590 = ~n588 & ~n589;
  assign n591 = ~pi129  & ~n590;
  assign n592 = ~n587 & ~n591;
  assign n593 = n265 & ~n592;
  assign n594 = pi53  & pi128 ;
  assign n595 = pi54  & ~pi128 ;
  assign n596 = ~n594 & ~n595;
  assign n597 = pi129  & ~n596;
  assign n598 = pi56  & ~pi128 ;
  assign n599 = pi55  & pi128 ;
  assign n600 = ~n598 & ~n599;
  assign n601 = ~pi129  & ~n600;
  assign n602 = ~n597 & ~n601;
  assign n603 = n276 & ~n602;
  assign n604 = pi61  & pi128 ;
  assign n605 = pi62  & ~pi128 ;
  assign n606 = ~n604 & ~n605;
  assign n607 = pi129  & ~n606;
  assign n608 = pi64  & ~pi128 ;
  assign n609 = pi63  & pi128 ;
  assign n610 = ~n608 & ~n609;
  assign n611 = ~pi129  & ~n610;
  assign n612 = ~n607 & ~n611;
  assign n613 = n287 & ~n612;
  assign n614 = pi49  & pi128 ;
  assign n615 = pi50  & ~pi128 ;
  assign n616 = ~n614 & ~n615;
  assign n617 = pi129  & ~n616;
  assign n618 = pi52  & ~pi128 ;
  assign n619 = pi51  & pi128 ;
  assign n620 = ~n618 & ~n619;
  assign n621 = ~pi129  & ~n620;
  assign n622 = ~n617 & ~n621;
  assign n623 = n298 & ~n622;
  assign n624 = ~n613 & ~n623;
  assign n625 = ~n603 & n624;
  assign n626 = ~n593 & n625;
  assign n627 = n403 & ~n626;
  assign n628 = ~n583 & ~n627;
  assign n629 = ~n539 & n628;
  assign n630 = ~n495 & n629;
  assign n631 = pi134  & ~n630;
  assign po0  = n451 | n631;
  assign n633 = pi93  & ~pi128 ;
  assign n634 = pi92  & pi128 ;
  assign n635 = ~n633 & ~n634;
  assign n636 = ~pi129  & ~n635;
  assign n637 = pi90  & pi128 ;
  assign n638 = pi91  & ~pi128 ;
  assign n639 = ~n637 & ~n638;
  assign n640 = pi129  & ~n639;
  assign n641 = ~n636 & ~n640;
  assign n642 = n265 & ~n641;
  assign n643 = pi89  & ~pi128 ;
  assign n644 = pi88  & pi128 ;
  assign n645 = ~n643 & ~n644;
  assign n646 = ~pi129  & ~n645;
  assign n647 = pi86  & pi128 ;
  assign n648 = pi87  & ~pi128 ;
  assign n649 = ~n647 & ~n648;
  assign n650 = pi129  & ~n649;
  assign n651 = ~n646 & ~n650;
  assign n652 = n276 & ~n651;
  assign n653 = pi97  & ~pi128 ;
  assign n654 = pi96  & pi128 ;
  assign n655 = ~n653 & ~n654;
  assign n656 = ~pi129  & ~n655;
  assign n657 = pi94  & pi128 ;
  assign n658 = pi95  & ~pi128 ;
  assign n659 = ~n657 & ~n658;
  assign n660 = pi129  & ~n659;
  assign n661 = ~n656 & ~n660;
  assign n662 = n287 & ~n661;
  assign n663 = pi85  & ~pi128 ;
  assign n664 = pi84  & pi128 ;
  assign n665 = ~n663 & ~n664;
  assign n666 = ~pi129  & ~n665;
  assign n667 = pi82  & pi128 ;
  assign n668 = pi83  & ~pi128 ;
  assign n669 = ~n667 & ~n668;
  assign n670 = pi129  & ~n669;
  assign n671 = ~n666 & ~n670;
  assign n672 = n298 & ~n671;
  assign n673 = ~n662 & ~n672;
  assign n674 = ~n652 & n673;
  assign n675 = ~n642 & n674;
  assign n676 = n264 & ~n675;
  assign n677 = pi109  & ~pi128 ;
  assign n678 = pi108  & pi128 ;
  assign n679 = ~n677 & ~n678;
  assign n680 = ~pi129  & ~n679;
  assign n681 = pi106  & pi128 ;
  assign n682 = pi107  & ~pi128 ;
  assign n683 = ~n681 & ~n682;
  assign n684 = pi129  & ~n683;
  assign n685 = ~n680 & ~n684;
  assign n686 = n265 & ~n685;
  assign n687 = pi105  & ~pi128 ;
  assign n688 = pi104  & pi128 ;
  assign n689 = ~n687 & ~n688;
  assign n690 = ~pi129  & ~n689;
  assign n691 = pi102  & pi128 ;
  assign n692 = pi103  & ~pi128 ;
  assign n693 = ~n691 & ~n692;
  assign n694 = pi129  & ~n693;
  assign n695 = ~n690 & ~n694;
  assign n696 = n276 & ~n695;
  assign n697 = pi113  & ~pi128 ;
  assign n698 = pi112  & pi128 ;
  assign n699 = ~n697 & ~n698;
  assign n700 = ~pi129  & ~n699;
  assign n701 = pi110  & pi128 ;
  assign n702 = pi111  & ~pi128 ;
  assign n703 = ~n701 & ~n702;
  assign n704 = pi129  & ~n703;
  assign n705 = ~n700 & ~n704;
  assign n706 = n287 & ~n705;
  assign n707 = pi101  & ~pi128 ;
  assign n708 = pi100  & pi128 ;
  assign n709 = ~n707 & ~n708;
  assign n710 = ~pi129  & ~n709;
  assign n711 = pi98  & pi128 ;
  assign n712 = pi99  & ~pi128 ;
  assign n713 = ~n711 & ~n712;
  assign n714 = pi129  & ~n713;
  assign n715 = ~n710 & ~n714;
  assign n716 = n298 & ~n715;
  assign n717 = ~n706 & ~n716;
  assign n718 = ~n696 & n717;
  assign n719 = ~n686 & n718;
  assign n720 = n313 & ~n719;
  assign n721 = pi77  & ~pi128 ;
  assign n722 = pi76  & pi128 ;
  assign n723 = ~n721 & ~n722;
  assign n724 = ~pi129  & ~n723;
  assign n725 = pi74  & pi128 ;
  assign n726 = pi75  & ~pi128 ;
  assign n727 = ~n725 & ~n726;
  assign n728 = pi129  & ~n727;
  assign n729 = ~n724 & ~n728;
  assign n730 = n265 & ~n729;
  assign n731 = pi73  & ~pi128 ;
  assign n732 = pi72  & pi128 ;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~pi129  & ~n733;
  assign n735 = pi70  & pi128 ;
  assign n736 = pi71  & ~pi128 ;
  assign n737 = ~n735 & ~n736;
  assign n738 = pi129  & ~n737;
  assign n739 = ~n734 & ~n738;
  assign n740 = n276 & ~n739;
  assign n741 = pi81  & ~pi128 ;
  assign n742 = pi80  & pi128 ;
  assign n743 = ~n741 & ~n742;
  assign n744 = ~pi129  & ~n743;
  assign n745 = pi78  & pi128 ;
  assign n746 = pi79  & ~pi128 ;
  assign n747 = ~n745 & ~n746;
  assign n748 = pi129  & ~n747;
  assign n749 = ~n744 & ~n748;
  assign n750 = n287 & ~n749;
  assign n751 = pi69  & ~pi128 ;
  assign n752 = pi68  & pi128 ;
  assign n753 = ~n751 & ~n752;
  assign n754 = ~pi129  & ~n753;
  assign n755 = pi66  & pi128 ;
  assign n756 = pi67  & ~pi128 ;
  assign n757 = ~n755 & ~n756;
  assign n758 = pi129  & ~n757;
  assign n759 = ~n754 & ~n758;
  assign n760 = n298 & ~n759;
  assign n761 = ~n750 & ~n760;
  assign n762 = ~n740 & n761;
  assign n763 = ~n730 & n762;
  assign n764 = n358 & ~n763;
  assign n765 = pi125  & ~pi128 ;
  assign n766 = pi124  & pi128 ;
  assign n767 = ~n765 & ~n766;
  assign n768 = ~pi129  & ~n767;
  assign n769 = pi122  & pi128 ;
  assign n770 = pi123  & ~pi128 ;
  assign n771 = ~n769 & ~n770;
  assign n772 = pi129  & ~n771;
  assign n773 = ~n768 & ~n772;
  assign n774 = n265 & ~n773;
  assign n775 = pi121  & ~pi128 ;
  assign n776 = pi120  & pi128 ;
  assign n777 = ~n775 & ~n776;
  assign n778 = ~pi129  & ~n777;
  assign n779 = pi118  & pi128 ;
  assign n780 = pi119  & ~pi128 ;
  assign n781 = ~n779 & ~n780;
  assign n782 = pi129  & ~n781;
  assign n783 = ~n778 & ~n782;
  assign n784 = n276 & ~n783;
  assign n785 = pi1  & ~pi128 ;
  assign n786 = pi0  & pi128 ;
  assign n787 = ~n785 & ~n786;
  assign n788 = ~pi129  & ~n787;
  assign n789 = pi126  & pi128 ;
  assign n790 = pi127  & ~pi128 ;
  assign n791 = ~n789 & ~n790;
  assign n792 = pi129  & ~n791;
  assign n793 = ~n788 & ~n792;
  assign n794 = n287 & ~n793;
  assign n795 = pi117  & ~pi128 ;
  assign n796 = pi116  & pi128 ;
  assign n797 = ~n795 & ~n796;
  assign n798 = ~pi129  & ~n797;
  assign n799 = pi114  & pi128 ;
  assign n800 = pi115  & ~pi128 ;
  assign n801 = ~n799 & ~n800;
  assign n802 = pi129  & ~n801;
  assign n803 = ~n798 & ~n802;
  assign n804 = n298 & ~n803;
  assign n805 = ~n794 & ~n804;
  assign n806 = ~n784 & n805;
  assign n807 = ~n774 & n806;
  assign n808 = n403 & ~n807;
  assign n809 = ~n764 & ~n808;
  assign n810 = ~n720 & n809;
  assign n811 = ~n676 & n810;
  assign n812 = ~pi134  & ~n811;
  assign n813 = pi13  & ~pi128 ;
  assign n814 = pi12  & pi128 ;
  assign n815 = ~n813 & ~n814;
  assign n816 = ~pi129  & ~n815;
  assign n817 = pi10  & pi128 ;
  assign n818 = pi11  & ~pi128 ;
  assign n819 = ~n817 & ~n818;
  assign n820 = pi129  & ~n819;
  assign n821 = ~n816 & ~n820;
  assign n822 = n265 & ~n821;
  assign n823 = pi9  & ~pi128 ;
  assign n824 = pi8  & pi128 ;
  assign n825 = ~n823 & ~n824;
  assign n826 = ~pi129  & ~n825;
  assign n827 = pi6  & pi128 ;
  assign n828 = pi7  & ~pi128 ;
  assign n829 = ~n827 & ~n828;
  assign n830 = pi129  & ~n829;
  assign n831 = ~n826 & ~n830;
  assign n832 = n276 & ~n831;
  assign n833 = pi17  & ~pi128 ;
  assign n834 = pi16  & pi128 ;
  assign n835 = ~n833 & ~n834;
  assign n836 = ~pi129  & ~n835;
  assign n837 = pi14  & pi128 ;
  assign n838 = pi15  & ~pi128 ;
  assign n839 = ~n837 & ~n838;
  assign n840 = pi129  & ~n839;
  assign n841 = ~n836 & ~n840;
  assign n842 = n287 & ~n841;
  assign n843 = pi5  & ~pi128 ;
  assign n844 = pi4  & pi128 ;
  assign n845 = ~n843 & ~n844;
  assign n846 = ~pi129  & ~n845;
  assign n847 = pi2  & pi128 ;
  assign n848 = pi3  & ~pi128 ;
  assign n849 = ~n847 & ~n848;
  assign n850 = pi129  & ~n849;
  assign n851 = ~n846 & ~n850;
  assign n852 = n298 & ~n851;
  assign n853 = ~n842 & ~n852;
  assign n854 = ~n832 & n853;
  assign n855 = ~n822 & n854;
  assign n856 = n358 & ~n855;
  assign n857 = pi29  & ~pi128 ;
  assign n858 = pi28  & pi128 ;
  assign n859 = ~n857 & ~n858;
  assign n860 = ~pi129  & ~n859;
  assign n861 = pi26  & pi128 ;
  assign n862 = pi27  & ~pi128 ;
  assign n863 = ~n861 & ~n862;
  assign n864 = pi129  & ~n863;
  assign n865 = ~n860 & ~n864;
  assign n866 = n265 & ~n865;
  assign n867 = pi25  & ~pi128 ;
  assign n868 = pi24  & pi128 ;
  assign n869 = ~n867 & ~n868;
  assign n870 = ~pi129  & ~n869;
  assign n871 = pi22  & pi128 ;
  assign n872 = pi23  & ~pi128 ;
  assign n873 = ~n871 & ~n872;
  assign n874 = pi129  & ~n873;
  assign n875 = ~n870 & ~n874;
  assign n876 = n276 & ~n875;
  assign n877 = pi33  & ~pi128 ;
  assign n878 = pi32  & pi128 ;
  assign n879 = ~n877 & ~n878;
  assign n880 = ~pi129  & ~n879;
  assign n881 = pi30  & pi128 ;
  assign n882 = pi31  & ~pi128 ;
  assign n883 = ~n881 & ~n882;
  assign n884 = pi129  & ~n883;
  assign n885 = ~n880 & ~n884;
  assign n886 = n287 & ~n885;
  assign n887 = pi21  & ~pi128 ;
  assign n888 = pi20  & pi128 ;
  assign n889 = ~n887 & ~n888;
  assign n890 = ~pi129  & ~n889;
  assign n891 = pi18  & pi128 ;
  assign n892 = pi19  & ~pi128 ;
  assign n893 = ~n891 & ~n892;
  assign n894 = pi129  & ~n893;
  assign n895 = ~n890 & ~n894;
  assign n896 = n298 & ~n895;
  assign n897 = ~n886 & ~n896;
  assign n898 = ~n876 & n897;
  assign n899 = ~n866 & n898;
  assign n900 = n264 & ~n899;
  assign n901 = pi61  & ~pi128 ;
  assign n902 = pi60  & pi128 ;
  assign n903 = ~n901 & ~n902;
  assign n904 = ~pi129  & ~n903;
  assign n905 = pi58  & pi128 ;
  assign n906 = pi59  & ~pi128 ;
  assign n907 = ~n905 & ~n906;
  assign n908 = pi129  & ~n907;
  assign n909 = ~n904 & ~n908;
  assign n910 = n265 & ~n909;
  assign n911 = pi57  & ~pi128 ;
  assign n912 = pi56  & pi128 ;
  assign n913 = ~n911 & ~n912;
  assign n914 = ~pi129  & ~n913;
  assign n915 = pi54  & pi128 ;
  assign n916 = pi55  & ~pi128 ;
  assign n917 = ~n915 & ~n916;
  assign n918 = pi129  & ~n917;
  assign n919 = ~n914 & ~n918;
  assign n920 = n276 & ~n919;
  assign n921 = pi65  & ~pi128 ;
  assign n922 = pi64  & pi128 ;
  assign n923 = ~n921 & ~n922;
  assign n924 = ~pi129  & ~n923;
  assign n925 = pi62  & pi128 ;
  assign n926 = pi63  & ~pi128 ;
  assign n927 = ~n925 & ~n926;
  assign n928 = pi129  & ~n927;
  assign n929 = ~n924 & ~n928;
  assign n930 = n287 & ~n929;
  assign n931 = pi53  & ~pi128 ;
  assign n932 = pi52  & pi128 ;
  assign n933 = ~n931 & ~n932;
  assign n934 = ~pi129  & ~n933;
  assign n935 = pi50  & pi128 ;
  assign n936 = pi51  & ~pi128 ;
  assign n937 = ~n935 & ~n936;
  assign n938 = pi129  & ~n937;
  assign n939 = ~n934 & ~n938;
  assign n940 = n298 & ~n939;
  assign n941 = ~n930 & ~n940;
  assign n942 = ~n920 & n941;
  assign n943 = ~n910 & n942;
  assign n944 = n403 & ~n943;
  assign n945 = pi42  & pi128 ;
  assign n946 = pi43  & ~pi128 ;
  assign n947 = ~n945 & ~n946;
  assign n948 = pi129  & ~n947;
  assign n949 = pi45  & ~pi128 ;
  assign n950 = pi44  & pi128 ;
  assign n951 = ~n949 & ~n950;
  assign n952 = ~pi129  & ~n951;
  assign n953 = ~n948 & ~n952;
  assign n954 = n265 & ~n953;
  assign n955 = pi41  & ~pi128 ;
  assign n956 = pi40  & pi128 ;
  assign n957 = ~n955 & ~n956;
  assign n958 = ~pi129  & ~n957;
  assign n959 = pi39  & ~pi128 ;
  assign n960 = pi38  & pi128 ;
  assign n961 = ~n959 & ~n960;
  assign n962 = pi129  & ~n961;
  assign n963 = ~n958 & ~n962;
  assign n964 = n276 & ~n963;
  assign n965 = pi49  & ~pi128 ;
  assign n966 = pi48  & pi128 ;
  assign n967 = ~n965 & ~n966;
  assign n968 = ~pi129  & ~n967;
  assign n969 = pi46  & pi128 ;
  assign n970 = pi47  & ~pi128 ;
  assign n971 = ~n969 & ~n970;
  assign n972 = pi129  & ~n971;
  assign n973 = ~n968 & ~n972;
  assign n974 = n287 & ~n973;
  assign n975 = pi37  & ~pi128 ;
  assign n976 = pi36  & pi128 ;
  assign n977 = ~n975 & ~n976;
  assign n978 = ~pi129  & ~n977;
  assign n979 = pi34  & pi128 ;
  assign n980 = pi35  & ~pi128 ;
  assign n981 = ~n979 & ~n980;
  assign n982 = pi129  & ~n981;
  assign n983 = ~n978 & ~n982;
  assign n984 = n298 & ~n983;
  assign n985 = ~n974 & ~n984;
  assign n986 = ~n964 & n985;
  assign n987 = ~n954 & n986;
  assign n988 = n313 & ~n987;
  assign n989 = ~n944 & ~n988;
  assign n990 = ~n900 & n989;
  assign n991 = ~n856 & n990;
  assign n992 = pi134  & ~n991;
  assign po1  = n812 | n992;
  assign n994 = ~pi129  & ~n290;
  assign n995 = pi129  & ~n272;
  assign n996 = ~n994 & ~n995;
  assign n997 = n265 & ~n996;
  assign n998 = ~pi129  & ~n268;
  assign n999 = pi129  & ~n283;
  assign n1000 = ~n998 & ~n999;
  assign n1001 = n276 & ~n1000;
  assign n1002 = ~pi129  & ~n346;
  assign n1003 = pi129  & ~n294;
  assign n1004 = ~n1002 & ~n1003;
  assign n1005 = n287 & ~n1004;
  assign n1006 = ~pi129  & ~n279;
  assign n1007 = pi129  & ~n305;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = n298 & ~n1008;
  assign n1010 = ~n1005 & ~n1009;
  assign n1011 = ~n1001 & n1010;
  assign n1012 = ~n997 & n1011;
  assign n1013 = n264 & ~n1012;
  assign n1014 = ~pi129  & ~n336;
  assign n1015 = pi129  & ~n320;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = n265 & ~n1016;
  assign n1018 = ~pi129  & ~n316;
  assign n1019 = pi129  & ~n330;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = n276 & ~n1020;
  assign n1022 = ~pi129  & ~n436;
  assign n1023 = pi129  & ~n340;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = n287 & ~n1024;
  assign n1026 = ~pi129  & ~n326;
  assign n1027 = pi129  & ~n350;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = n298 & ~n1028;
  assign n1030 = ~n1025 & ~n1029;
  assign n1031 = ~n1021 & n1030;
  assign n1032 = ~n1017 & n1031;
  assign n1033 = n313 & ~n1032;
  assign n1034 = ~pi129  & ~n381;
  assign n1035 = pi129  & ~n365;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = n265 & ~n1036;
  assign n1038 = ~pi129  & ~n361;
  assign n1039 = pi129  & ~n375;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = n276 & ~n1040;
  assign n1042 = ~pi129  & ~n301;
  assign n1043 = pi129  & ~n385;
  assign n1044 = ~n1042 & ~n1043;
  assign n1045 = n287 & ~n1044;
  assign n1046 = ~pi129  & ~n371;
  assign n1047 = pi129  & ~n395;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = n298 & ~n1048;
  assign n1050 = ~n1045 & ~n1049;
  assign n1051 = ~n1041 & n1050;
  assign n1052 = ~n1037 & n1051;
  assign n1053 = n358 & ~n1052;
  assign n1054 = ~pi129  & ~n426;
  assign n1055 = pi129  & ~n410;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = n265 & ~n1056;
  assign n1058 = ~pi129  & ~n406;
  assign n1059 = pi129  & ~n420;
  assign n1060 = ~n1058 & ~n1059;
  assign n1061 = n276 & ~n1060;
  assign n1062 = ~pi129  & ~n572;
  assign n1063 = pi129  & ~n430;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = n287 & ~n1064;
  assign n1066 = ~pi129  & ~n416;
  assign n1067 = pi129  & ~n440;
  assign n1068 = ~n1066 & ~n1067;
  assign n1069 = n298 & ~n1068;
  assign n1070 = ~n1065 & ~n1069;
  assign n1071 = ~n1061 & n1070;
  assign n1072 = ~n1057 & n1071;
  assign n1073 = n403 & ~n1072;
  assign n1074 = ~n1053 & ~n1073;
  assign n1075 = ~n1033 & n1074;
  assign n1076 = ~n1013 & n1075;
  assign n1077 = ~pi134  & ~n1076;
  assign n1078 = ~pi129  & ~n562;
  assign n1079 = pi129  & ~n546;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = n265 & ~n1080;
  assign n1082 = ~pi129  & ~n542;
  assign n1083 = pi129  & ~n556;
  assign n1084 = ~n1082 & ~n1083;
  assign n1085 = n276 & ~n1084;
  assign n1086 = ~pi129  & ~n484;
  assign n1087 = pi129  & ~n566;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = n287 & ~n1088;
  assign n1090 = ~pi129  & ~n552;
  assign n1091 = pi129  & ~n576;
  assign n1092 = ~n1090 & ~n1091;
  assign n1093 = n298 & ~n1092;
  assign n1094 = ~n1089 & ~n1093;
  assign n1095 = ~n1085 & n1094;
  assign n1096 = ~n1081 & n1095;
  assign n1097 = n358 & ~n1096;
  assign n1098 = ~pi129  & ~n474;
  assign n1099 = pi129  & ~n458;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = n265 & ~n1100;
  assign n1102 = ~pi129  & ~n454;
  assign n1103 = pi129  & ~n468;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = n276 & ~n1104;
  assign n1106 = ~pi129  & ~n528;
  assign n1107 = pi129  & ~n478;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = n287 & ~n1108;
  assign n1110 = ~pi129  & ~n464;
  assign n1111 = pi129  & ~n488;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = n298 & ~n1112;
  assign n1114 = ~n1109 & ~n1113;
  assign n1115 = ~n1105 & n1114;
  assign n1116 = ~n1101 & n1115;
  assign n1117 = n264 & ~n1116;
  assign n1118 = ~pi129  & ~n606;
  assign n1119 = pi129  & ~n590;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = n265 & ~n1120;
  assign n1122 = ~pi129  & ~n586;
  assign n1123 = pi129  & ~n600;
  assign n1124 = ~n1122 & ~n1123;
  assign n1125 = n276 & ~n1124;
  assign n1126 = ~pi129  & ~n391;
  assign n1127 = pi129  & ~n610;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = n287 & ~n1128;
  assign n1130 = ~pi129  & ~n596;
  assign n1131 = pi129  & ~n620;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = n298 & ~n1132;
  assign n1134 = ~n1129 & ~n1133;
  assign n1135 = ~n1125 & n1134;
  assign n1136 = ~n1121 & n1135;
  assign n1137 = n403 & ~n1136;
  assign n1138 = pi129  & ~n502;
  assign n1139 = ~pi129  & ~n518;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = n265 & ~n1140;
  assign n1142 = ~pi129  & ~n498;
  assign n1143 = pi129  & ~n508;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = n276 & ~n1144;
  assign n1146 = ~pi129  & ~n616;
  assign n1147 = pi129  & ~n522;
  assign n1148 = ~n1146 & ~n1147;
  assign n1149 = n287 & ~n1148;
  assign n1150 = ~pi129  & ~n512;
  assign n1151 = pi129  & ~n532;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = n298 & ~n1152;
  assign n1154 = ~n1149 & ~n1153;
  assign n1155 = ~n1145 & n1154;
  assign n1156 = ~n1141 & n1155;
  assign n1157 = n313 & ~n1156;
  assign n1158 = ~n1137 & ~n1157;
  assign n1159 = ~n1117 & n1158;
  assign n1160 = ~n1097 & n1159;
  assign n1161 = pi134  & ~n1160;
  assign po2  = n1077 | n1161;
  assign n1163 = ~pi129  & ~n659;
  assign n1164 = pi129  & ~n635;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = n265 & ~n1165;
  assign n1167 = ~pi129  & ~n639;
  assign n1168 = pi129  & ~n645;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = n276 & ~n1169;
  assign n1171 = ~pi129  & ~n713;
  assign n1172 = pi129  & ~n655;
  assign n1173 = ~n1171 & ~n1172;
  assign n1174 = n287 & ~n1173;
  assign n1175 = ~pi129  & ~n649;
  assign n1176 = pi129  & ~n665;
  assign n1177 = ~n1175 & ~n1176;
  assign n1178 = n298 & ~n1177;
  assign n1179 = ~n1174 & ~n1178;
  assign n1180 = ~n1170 & n1179;
  assign n1181 = ~n1166 & n1180;
  assign n1182 = n264 & ~n1181;
  assign n1183 = ~pi129  & ~n747;
  assign n1184 = pi129  & ~n723;
  assign n1185 = ~n1183 & ~n1184;
  assign n1186 = n265 & ~n1185;
  assign n1187 = ~pi129  & ~n727;
  assign n1188 = pi129  & ~n733;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = n276 & ~n1189;
  assign n1191 = ~pi129  & ~n669;
  assign n1192 = pi129  & ~n743;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = n287 & ~n1193;
  assign n1195 = ~pi129  & ~n737;
  assign n1196 = pi129  & ~n753;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = n298 & ~n1197;
  assign n1199 = ~n1194 & ~n1198;
  assign n1200 = ~n1190 & n1199;
  assign n1201 = ~n1186 & n1200;
  assign n1202 = n358 & ~n1201;
  assign n1203 = ~pi129  & ~n703;
  assign n1204 = pi129  & ~n679;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = n265 & ~n1205;
  assign n1207 = ~pi129  & ~n683;
  assign n1208 = pi129  & ~n689;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = n276 & ~n1209;
  assign n1211 = ~pi129  & ~n801;
  assign n1212 = pi129  & ~n699;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = n287 & ~n1213;
  assign n1215 = ~pi129  & ~n693;
  assign n1216 = pi129  & ~n709;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = n298 & ~n1217;
  assign n1219 = ~n1214 & ~n1218;
  assign n1220 = ~n1210 & n1219;
  assign n1221 = ~n1206 & n1220;
  assign n1222 = n313 & ~n1221;
  assign n1223 = ~pi129  & ~n791;
  assign n1224 = pi129  & ~n767;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = n265 & ~n1225;
  assign n1227 = ~pi129  & ~n771;
  assign n1228 = pi129  & ~n777;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = n276 & ~n1229;
  assign n1231 = ~pi129  & ~n849;
  assign n1232 = pi129  & ~n787;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = n287 & ~n1233;
  assign n1235 = ~pi129  & ~n781;
  assign n1236 = pi129  & ~n797;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = n298 & ~n1237;
  assign n1239 = ~n1234 & ~n1238;
  assign n1240 = ~n1230 & n1239;
  assign n1241 = ~n1226 & n1240;
  assign n1242 = n403 & ~n1241;
  assign n1243 = ~n1222 & ~n1242;
  assign n1244 = ~n1202 & n1243;
  assign n1245 = ~n1182 & n1244;
  assign n1246 = ~pi134  & ~n1245;
  assign n1247 = pi129  & ~n951;
  assign n1248 = ~pi129  & ~n971;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = n265 & ~n1249;
  assign n1251 = ~pi129  & ~n947;
  assign n1252 = pi129  & ~n957;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = n276 & ~n1253;
  assign n1255 = ~pi129  & ~n937;
  assign n1256 = pi129  & ~n967;
  assign n1257 = ~n1255 & ~n1256;
  assign n1258 = n287 & ~n1257;
  assign n1259 = ~pi129  & ~n961;
  assign n1260 = pi129  & ~n977;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = n298 & ~n1261;
  assign n1263 = ~n1258 & ~n1262;
  assign n1264 = ~n1254 & n1263;
  assign n1265 = ~n1250 & n1264;
  assign n1266 = n313 & ~n1265;
  assign n1267 = ~pi129  & ~n883;
  assign n1268 = pi129  & ~n859;
  assign n1269 = ~n1267 & ~n1268;
  assign n1270 = n265 & ~n1269;
  assign n1271 = ~pi129  & ~n863;
  assign n1272 = pi129  & ~n869;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = n276 & ~n1273;
  assign n1275 = ~pi129  & ~n981;
  assign n1276 = pi129  & ~n879;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = n287 & ~n1277;
  assign n1279 = ~pi129  & ~n873;
  assign n1280 = pi129  & ~n889;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = n298 & ~n1281;
  assign n1283 = ~n1278 & ~n1282;
  assign n1284 = ~n1274 & n1283;
  assign n1285 = ~n1270 & n1284;
  assign n1286 = n264 & ~n1285;
  assign n1287 = ~pi129  & ~n927;
  assign n1288 = pi129  & ~n903;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = n265 & ~n1289;
  assign n1291 = ~pi129  & ~n907;
  assign n1292 = pi129  & ~n913;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = n276 & ~n1293;
  assign n1295 = ~pi129  & ~n757;
  assign n1296 = pi129  & ~n923;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = n287 & ~n1297;
  assign n1299 = ~pi129  & ~n917;
  assign n1300 = pi129  & ~n933;
  assign n1301 = ~n1299 & ~n1300;
  assign n1302 = n298 & ~n1301;
  assign n1303 = ~n1298 & ~n1302;
  assign n1304 = ~n1294 & n1303;
  assign n1305 = ~n1290 & n1304;
  assign n1306 = n403 & ~n1305;
  assign n1307 = ~pi129  & ~n839;
  assign n1308 = pi129  & ~n815;
  assign n1309 = ~n1307 & ~n1308;
  assign n1310 = n265 & ~n1309;
  assign n1311 = ~pi129  & ~n819;
  assign n1312 = pi129  & ~n825;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = n276 & ~n1313;
  assign n1315 = ~pi129  & ~n893;
  assign n1316 = pi129  & ~n835;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = n287 & ~n1317;
  assign n1319 = ~pi129  & ~n829;
  assign n1320 = pi129  & ~n845;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = n298 & ~n1321;
  assign n1323 = ~n1318 & ~n1322;
  assign n1324 = ~n1314 & n1323;
  assign n1325 = ~n1310 & n1324;
  assign n1326 = n358 & ~n1325;
  assign n1327 = ~n1306 & ~n1326;
  assign n1328 = ~n1286 & n1327;
  assign n1329 = ~n1266 & n1328;
  assign n1330 = pi134  & ~n1329;
  assign po3  = n1246 | n1330;
  assign n1332 = n265 & ~n296;
  assign n1333 = ~n274 & n276;
  assign n1334 = n287 & ~n352;
  assign n1335 = ~n285 & n298;
  assign n1336 = ~n1334 & ~n1335;
  assign n1337 = ~n1333 & n1336;
  assign n1338 = ~n1332 & n1337;
  assign n1339 = n264 & ~n1338;
  assign n1340 = n265 & ~n342;
  assign n1341 = n276 & ~n322;
  assign n1342 = n287 & ~n442;
  assign n1343 = n298 & ~n332;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = ~n1341 & n1344;
  assign n1346 = ~n1340 & n1345;
  assign n1347 = n313 & ~n1346;
  assign n1348 = n265 & ~n387;
  assign n1349 = n276 & ~n367;
  assign n1350 = n287 & ~n307;
  assign n1351 = n298 & ~n377;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = ~n1349 & n1352;
  assign n1354 = ~n1348 & n1353;
  assign n1355 = n358 & ~n1354;
  assign n1356 = n265 & ~n432;
  assign n1357 = n276 & ~n412;
  assign n1358 = n287 & ~n578;
  assign n1359 = n298 & ~n422;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = ~n1357 & n1360;
  assign n1362 = ~n1356 & n1361;
  assign n1363 = n403 & ~n1362;
  assign n1364 = ~n1355 & ~n1363;
  assign n1365 = ~n1347 & n1364;
  assign n1366 = ~n1339 & n1365;
  assign n1367 = ~pi134  & ~n1366;
  assign n1368 = n265 & ~n612;
  assign n1369 = n276 & ~n592;
  assign n1370 = n287 & ~n397;
  assign n1371 = n298 & ~n602;
  assign n1372 = ~n1370 & ~n1371;
  assign n1373 = ~n1369 & n1372;
  assign n1374 = ~n1368 & n1373;
  assign n1375 = n403 & ~n1374;
  assign n1376 = n265 & ~n568;
  assign n1377 = n276 & ~n548;
  assign n1378 = n287 & ~n490;
  assign n1379 = n298 & ~n558;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = ~n1377 & n1380;
  assign n1382 = ~n1376 & n1381;
  assign n1383 = n358 & ~n1382;
  assign n1384 = n265 & ~n524;
  assign n1385 = n276 & ~n504;
  assign n1386 = n287 & ~n622;
  assign n1387 = n298 & ~n514;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = ~n1385 & n1388;
  assign n1390 = ~n1384 & n1389;
  assign n1391 = n313 & ~n1390;
  assign n1392 = n265 & ~n480;
  assign n1393 = n276 & ~n460;
  assign n1394 = n287 & ~n534;
  assign n1395 = n298 & ~n470;
  assign n1396 = ~n1394 & ~n1395;
  assign n1397 = ~n1393 & n1396;
  assign n1398 = ~n1392 & n1397;
  assign n1399 = n264 & ~n1398;
  assign n1400 = ~n1391 & ~n1399;
  assign n1401 = ~n1383 & n1400;
  assign n1402 = ~n1375 & n1401;
  assign n1403 = pi134  & ~n1402;
  assign po4  = n1367 | n1403;
  assign n1405 = n265 & ~n661;
  assign n1406 = n276 & ~n641;
  assign n1407 = n287 & ~n715;
  assign n1408 = n298 & ~n651;
  assign n1409 = ~n1407 & ~n1408;
  assign n1410 = ~n1406 & n1409;
  assign n1411 = ~n1405 & n1410;
  assign n1412 = n264 & ~n1411;
  assign n1413 = n265 & ~n705;
  assign n1414 = n276 & ~n685;
  assign n1415 = n287 & ~n803;
  assign n1416 = n298 & ~n695;
  assign n1417 = ~n1415 & ~n1416;
  assign n1418 = ~n1414 & n1417;
  assign n1419 = ~n1413 & n1418;
  assign n1420 = n313 & ~n1419;
  assign n1421 = n265 & ~n749;
  assign n1422 = n276 & ~n729;
  assign n1423 = n287 & ~n671;
  assign n1424 = n298 & ~n739;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = ~n1422 & n1425;
  assign n1427 = ~n1421 & n1426;
  assign n1428 = n358 & ~n1427;
  assign n1429 = n265 & ~n793;
  assign n1430 = n276 & ~n773;
  assign n1431 = n287 & ~n851;
  assign n1432 = n298 & ~n783;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = ~n1430 & n1433;
  assign n1435 = ~n1429 & n1434;
  assign n1436 = n403 & ~n1435;
  assign n1437 = ~n1428 & ~n1436;
  assign n1438 = ~n1420 & n1437;
  assign n1439 = ~n1412 & n1438;
  assign n1440 = ~pi134  & ~n1439;
  assign n1441 = n265 & ~n929;
  assign n1442 = n276 & ~n909;
  assign n1443 = n287 & ~n759;
  assign n1444 = n298 & ~n919;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = ~n1442 & n1445;
  assign n1447 = ~n1441 & n1446;
  assign n1448 = n403 & ~n1447;
  assign n1449 = n265 & ~n841;
  assign n1450 = n276 & ~n821;
  assign n1451 = n287 & ~n895;
  assign n1452 = n298 & ~n831;
  assign n1453 = ~n1451 & ~n1452;
  assign n1454 = ~n1450 & n1453;
  assign n1455 = ~n1449 & n1454;
  assign n1456 = n358 & ~n1455;
  assign n1457 = n265 & ~n973;
  assign n1458 = n276 & ~n953;
  assign n1459 = n287 & ~n939;
  assign n1460 = n298 & ~n963;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = ~n1458 & n1461;
  assign n1463 = ~n1457 & n1462;
  assign n1464 = n313 & ~n1463;
  assign n1465 = n265 & ~n885;
  assign n1466 = n276 & ~n865;
  assign n1467 = n287 & ~n983;
  assign n1468 = n298 & ~n875;
  assign n1469 = ~n1467 & ~n1468;
  assign n1470 = ~n1466 & n1469;
  assign n1471 = ~n1465 & n1470;
  assign n1472 = n264 & ~n1471;
  assign n1473 = ~n1464 & ~n1472;
  assign n1474 = ~n1456 & n1473;
  assign n1475 = ~n1448 & n1474;
  assign n1476 = pi134  & ~n1475;
  assign po5  = n1440 | n1476;
  assign n1478 = n265 & ~n1004;
  assign n1479 = n276 & ~n996;
  assign n1480 = n287 & ~n1028;
  assign n1481 = n298 & ~n1000;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = ~n1479 & n1482;
  assign n1484 = ~n1478 & n1483;
  assign n1485 = n264 & ~n1484;
  assign n1486 = n265 & ~n1024;
  assign n1487 = n276 & ~n1016;
  assign n1488 = n287 & ~n1068;
  assign n1489 = n298 & ~n1020;
  assign n1490 = ~n1488 & ~n1489;
  assign n1491 = ~n1487 & n1490;
  assign n1492 = ~n1486 & n1491;
  assign n1493 = n313 & ~n1492;
  assign n1494 = n265 & ~n1044;
  assign n1495 = n276 & ~n1036;
  assign n1496 = n287 & ~n1008;
  assign n1497 = n298 & ~n1040;
  assign n1498 = ~n1496 & ~n1497;
  assign n1499 = ~n1495 & n1498;
  assign n1500 = ~n1494 & n1499;
  assign n1501 = n358 & ~n1500;
  assign n1502 = n265 & ~n1064;
  assign n1503 = n276 & ~n1056;
  assign n1504 = n287 & ~n1092;
  assign n1505 = n298 & ~n1060;
  assign n1506 = ~n1504 & ~n1505;
  assign n1507 = ~n1503 & n1506;
  assign n1508 = ~n1502 & n1507;
  assign n1509 = n403 & ~n1508;
  assign n1510 = ~n1501 & ~n1509;
  assign n1511 = ~n1493 & n1510;
  assign n1512 = ~n1485 & n1511;
  assign n1513 = ~pi134  & ~n1512;
  assign n1514 = n265 & ~n1128;
  assign n1515 = n276 & ~n1120;
  assign n1516 = n287 & ~n1048;
  assign n1517 = n298 & ~n1124;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = ~n1515 & n1518;
  assign n1520 = ~n1514 & n1519;
  assign n1521 = n403 & ~n1520;
  assign n1522 = n265 & ~n1088;
  assign n1523 = n276 & ~n1080;
  assign n1524 = n287 & ~n1112;
  assign n1525 = n298 & ~n1084;
  assign n1526 = ~n1524 & ~n1525;
  assign n1527 = ~n1523 & n1526;
  assign n1528 = ~n1522 & n1527;
  assign n1529 = n358 & ~n1528;
  assign n1530 = n265 & ~n1148;
  assign n1531 = n276 & ~n1140;
  assign n1532 = n287 & ~n1132;
  assign n1533 = n298 & ~n1144;
  assign n1534 = ~n1532 & ~n1533;
  assign n1535 = ~n1531 & n1534;
  assign n1536 = ~n1530 & n1535;
  assign n1537 = n313 & ~n1536;
  assign n1538 = n265 & ~n1108;
  assign n1539 = n276 & ~n1100;
  assign n1540 = n287 & ~n1152;
  assign n1541 = n298 & ~n1104;
  assign n1542 = ~n1540 & ~n1541;
  assign n1543 = ~n1539 & n1542;
  assign n1544 = ~n1538 & n1543;
  assign n1545 = n264 & ~n1544;
  assign n1546 = ~n1537 & ~n1545;
  assign n1547 = ~n1529 & n1546;
  assign n1548 = ~n1521 & n1547;
  assign n1549 = pi134  & ~n1548;
  assign po6  = n1513 | n1549;
  assign n1551 = n265 & ~n1173;
  assign n1552 = n276 & ~n1165;
  assign n1553 = n287 & ~n1217;
  assign n1554 = n298 & ~n1169;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = ~n1552 & n1555;
  assign n1557 = ~n1551 & n1556;
  assign n1558 = n264 & ~n1557;
  assign n1559 = n265 & ~n1213;
  assign n1560 = n276 & ~n1205;
  assign n1561 = n287 & ~n1237;
  assign n1562 = n298 & ~n1209;
  assign n1563 = ~n1561 & ~n1562;
  assign n1564 = ~n1560 & n1563;
  assign n1565 = ~n1559 & n1564;
  assign n1566 = n313 & ~n1565;
  assign n1567 = n265 & ~n1193;
  assign n1568 = n276 & ~n1185;
  assign n1569 = n287 & ~n1177;
  assign n1570 = n298 & ~n1189;
  assign n1571 = ~n1569 & ~n1570;
  assign n1572 = ~n1568 & n1571;
  assign n1573 = ~n1567 & n1572;
  assign n1574 = n358 & ~n1573;
  assign n1575 = n265 & ~n1233;
  assign n1576 = n276 & ~n1225;
  assign n1577 = n287 & ~n1321;
  assign n1578 = n298 & ~n1229;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = ~n1576 & n1579;
  assign n1581 = ~n1575 & n1580;
  assign n1582 = n403 & ~n1581;
  assign n1583 = ~n1574 & ~n1582;
  assign n1584 = ~n1566 & n1583;
  assign n1585 = ~n1558 & n1584;
  assign n1586 = ~pi134  & ~n1585;
  assign n1587 = n265 & ~n1297;
  assign n1588 = n276 & ~n1289;
  assign n1589 = n287 & ~n1197;
  assign n1590 = n298 & ~n1293;
  assign n1591 = ~n1589 & ~n1590;
  assign n1592 = ~n1588 & n1591;
  assign n1593 = ~n1587 & n1592;
  assign n1594 = n403 & ~n1593;
  assign n1595 = n265 & ~n1317;
  assign n1596 = n276 & ~n1309;
  assign n1597 = n287 & ~n1281;
  assign n1598 = n298 & ~n1313;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = ~n1596 & n1599;
  assign n1601 = ~n1595 & n1600;
  assign n1602 = n358 & ~n1601;
  assign n1603 = n276 & ~n1249;
  assign n1604 = n287 & ~n1301;
  assign n1605 = n265 & ~n1257;
  assign n1606 = n298 & ~n1253;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = ~n1604 & n1607;
  assign n1609 = ~n1603 & n1608;
  assign n1610 = n313 & ~n1609;
  assign n1611 = n265 & ~n1277;
  assign n1612 = n276 & ~n1269;
  assign n1613 = n287 & ~n1261;
  assign n1614 = n298 & ~n1273;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n1612 & n1615;
  assign n1617 = ~n1611 & n1616;
  assign n1618 = n264 & ~n1617;
  assign n1619 = ~n1610 & ~n1618;
  assign n1620 = ~n1602 & n1619;
  assign n1621 = ~n1594 & n1620;
  assign n1622 = pi134  & ~n1621;
  assign po7  = n1586 | n1622;
  assign n1624 = n265 & ~n352;
  assign n1625 = n276 & ~n296;
  assign n1626 = n287 & ~n332;
  assign n1627 = ~n274 & n298;
  assign n1628 = ~n1626 & ~n1627;
  assign n1629 = ~n1625 & n1628;
  assign n1630 = ~n1624 & n1629;
  assign n1631 = n264 & ~n1630;
  assign n1632 = n265 & ~n442;
  assign n1633 = n276 & ~n342;
  assign n1634 = n287 & ~n422;
  assign n1635 = n298 & ~n322;
  assign n1636 = ~n1634 & ~n1635;
  assign n1637 = ~n1633 & n1636;
  assign n1638 = ~n1632 & n1637;
  assign n1639 = n313 & ~n1638;
  assign n1640 = n265 & ~n307;
  assign n1641 = n276 & ~n387;
  assign n1642 = ~n285 & n287;
  assign n1643 = n298 & ~n367;
  assign n1644 = ~n1642 & ~n1643;
  assign n1645 = ~n1641 & n1644;
  assign n1646 = ~n1640 & n1645;
  assign n1647 = n358 & ~n1646;
  assign n1648 = n265 & ~n578;
  assign n1649 = n276 & ~n432;
  assign n1650 = n287 & ~n558;
  assign n1651 = n298 & ~n412;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = ~n1649 & n1652;
  assign n1654 = ~n1648 & n1653;
  assign n1655 = n403 & ~n1654;
  assign n1656 = ~n1647 & ~n1655;
  assign n1657 = ~n1639 & n1656;
  assign n1658 = ~n1631 & n1657;
  assign n1659 = ~pi134  & ~n1658;
  assign n1660 = n265 & ~n397;
  assign n1661 = n276 & ~n612;
  assign n1662 = n287 & ~n377;
  assign n1663 = n298 & ~n592;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = ~n1661 & n1664;
  assign n1666 = ~n1660 & n1665;
  assign n1667 = n403 & ~n1666;
  assign n1668 = n265 & ~n490;
  assign n1669 = n276 & ~n568;
  assign n1670 = n287 & ~n470;
  assign n1671 = n298 & ~n548;
  assign n1672 = ~n1670 & ~n1671;
  assign n1673 = ~n1669 & n1672;
  assign n1674 = ~n1668 & n1673;
  assign n1675 = n358 & ~n1674;
  assign n1676 = n265 & ~n622;
  assign n1677 = n276 & ~n524;
  assign n1678 = n287 & ~n602;
  assign n1679 = n298 & ~n504;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = ~n1677 & n1680;
  assign n1682 = ~n1676 & n1681;
  assign n1683 = n313 & ~n1682;
  assign n1684 = n265 & ~n534;
  assign n1685 = n276 & ~n480;
  assign n1686 = n287 & ~n514;
  assign n1687 = n298 & ~n460;
  assign n1688 = ~n1686 & ~n1687;
  assign n1689 = ~n1685 & n1688;
  assign n1690 = ~n1684 & n1689;
  assign n1691 = n264 & ~n1690;
  assign n1692 = ~n1683 & ~n1691;
  assign n1693 = ~n1675 & n1692;
  assign n1694 = ~n1667 & n1693;
  assign n1695 = pi134  & ~n1694;
  assign po8  = n1659 | n1695;
  assign n1697 = n265 & ~n715;
  assign n1698 = n276 & ~n661;
  assign n1699 = n287 & ~n695;
  assign n1700 = n298 & ~n641;
  assign n1701 = ~n1699 & ~n1700;
  assign n1702 = ~n1698 & n1701;
  assign n1703 = ~n1697 & n1702;
  assign n1704 = n264 & ~n1703;
  assign n1705 = n265 & ~n803;
  assign n1706 = n276 & ~n705;
  assign n1707 = n287 & ~n783;
  assign n1708 = n298 & ~n685;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = ~n1706 & n1709;
  assign n1711 = ~n1705 & n1710;
  assign n1712 = n313 & ~n1711;
  assign n1713 = n265 & ~n671;
  assign n1714 = n276 & ~n749;
  assign n1715 = n287 & ~n651;
  assign n1716 = n298 & ~n729;
  assign n1717 = ~n1715 & ~n1716;
  assign n1718 = ~n1714 & n1717;
  assign n1719 = ~n1713 & n1718;
  assign n1720 = n358 & ~n1719;
  assign n1721 = n265 & ~n851;
  assign n1722 = n276 & ~n793;
  assign n1723 = n287 & ~n831;
  assign n1724 = n298 & ~n773;
  assign n1725 = ~n1723 & ~n1724;
  assign n1726 = ~n1722 & n1725;
  assign n1727 = ~n1721 & n1726;
  assign n1728 = n403 & ~n1727;
  assign n1729 = ~n1720 & ~n1728;
  assign n1730 = ~n1712 & n1729;
  assign n1731 = ~n1704 & n1730;
  assign n1732 = ~pi134  & ~n1731;
  assign n1733 = n265 & ~n759;
  assign n1734 = n276 & ~n929;
  assign n1735 = n287 & ~n739;
  assign n1736 = n298 & ~n909;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = ~n1734 & n1737;
  assign n1739 = ~n1733 & n1738;
  assign n1740 = n403 & ~n1739;
  assign n1741 = n265 & ~n895;
  assign n1742 = n276 & ~n841;
  assign n1743 = n287 & ~n875;
  assign n1744 = n298 & ~n821;
  assign n1745 = ~n1743 & ~n1744;
  assign n1746 = ~n1742 & n1745;
  assign n1747 = ~n1741 & n1746;
  assign n1748 = n358 & ~n1747;
  assign n1749 = n265 & ~n939;
  assign n1750 = n276 & ~n973;
  assign n1751 = n287 & ~n919;
  assign n1752 = n298 & ~n953;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = ~n1750 & n1753;
  assign n1755 = ~n1749 & n1754;
  assign n1756 = n313 & ~n1755;
  assign n1757 = n265 & ~n983;
  assign n1758 = n276 & ~n885;
  assign n1759 = n287 & ~n963;
  assign n1760 = n298 & ~n865;
  assign n1761 = ~n1759 & ~n1760;
  assign n1762 = ~n1758 & n1761;
  assign n1763 = ~n1757 & n1762;
  assign n1764 = n264 & ~n1763;
  assign n1765 = ~n1756 & ~n1764;
  assign n1766 = ~n1748 & n1765;
  assign n1767 = ~n1740 & n1766;
  assign n1768 = pi134  & ~n1767;
  assign po9  = n1732 | n1768;
  assign n1770 = n265 & ~n1028;
  assign n1771 = n276 & ~n1004;
  assign n1772 = n287 & ~n1020;
  assign n1773 = n298 & ~n996;
  assign n1774 = ~n1772 & ~n1773;
  assign n1775 = ~n1771 & n1774;
  assign n1776 = ~n1770 & n1775;
  assign n1777 = n264 & ~n1776;
  assign n1778 = n265 & ~n1068;
  assign n1779 = n276 & ~n1024;
  assign n1780 = n287 & ~n1060;
  assign n1781 = n298 & ~n1016;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = ~n1779 & n1782;
  assign n1784 = ~n1778 & n1783;
  assign n1785 = n313 & ~n1784;
  assign n1786 = n265 & ~n1008;
  assign n1787 = n276 & ~n1044;
  assign n1788 = n287 & ~n1000;
  assign n1789 = n298 & ~n1036;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = ~n1787 & n1790;
  assign n1792 = ~n1786 & n1791;
  assign n1793 = n358 & ~n1792;
  assign n1794 = n265 & ~n1092;
  assign n1795 = n276 & ~n1064;
  assign n1796 = n287 & ~n1084;
  assign n1797 = n298 & ~n1056;
  assign n1798 = ~n1796 & ~n1797;
  assign n1799 = ~n1795 & n1798;
  assign n1800 = ~n1794 & n1799;
  assign n1801 = n403 & ~n1800;
  assign n1802 = ~n1793 & ~n1801;
  assign n1803 = ~n1785 & n1802;
  assign n1804 = ~n1777 & n1803;
  assign n1805 = ~pi134  & ~n1804;
  assign n1806 = n265 & ~n1048;
  assign n1807 = n276 & ~n1128;
  assign n1808 = n287 & ~n1040;
  assign n1809 = n298 & ~n1120;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = ~n1807 & n1810;
  assign n1812 = ~n1806 & n1811;
  assign n1813 = n403 & ~n1812;
  assign n1814 = n265 & ~n1112;
  assign n1815 = n276 & ~n1088;
  assign n1816 = n287 & ~n1104;
  assign n1817 = n298 & ~n1080;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = ~n1815 & n1818;
  assign n1820 = ~n1814 & n1819;
  assign n1821 = n358 & ~n1820;
  assign n1822 = n265 & ~n1132;
  assign n1823 = n276 & ~n1148;
  assign n1824 = n287 & ~n1124;
  assign n1825 = n298 & ~n1140;
  assign n1826 = ~n1824 & ~n1825;
  assign n1827 = ~n1823 & n1826;
  assign n1828 = ~n1822 & n1827;
  assign n1829 = n313 & ~n1828;
  assign n1830 = n265 & ~n1152;
  assign n1831 = n276 & ~n1108;
  assign n1832 = n287 & ~n1144;
  assign n1833 = n298 & ~n1100;
  assign n1834 = ~n1832 & ~n1833;
  assign n1835 = ~n1831 & n1834;
  assign n1836 = ~n1830 & n1835;
  assign n1837 = n264 & ~n1836;
  assign n1838 = ~n1829 & ~n1837;
  assign n1839 = ~n1821 & n1838;
  assign n1840 = ~n1813 & n1839;
  assign n1841 = pi134  & ~n1840;
  assign po10  = n1805 | n1841;
  assign n1843 = n265 & ~n1217;
  assign n1844 = n276 & ~n1173;
  assign n1845 = n287 & ~n1209;
  assign n1846 = n298 & ~n1165;
  assign n1847 = ~n1845 & ~n1846;
  assign n1848 = ~n1844 & n1847;
  assign n1849 = ~n1843 & n1848;
  assign n1850 = n264 & ~n1849;
  assign n1851 = n265 & ~n1237;
  assign n1852 = n276 & ~n1213;
  assign n1853 = n287 & ~n1229;
  assign n1854 = n298 & ~n1205;
  assign n1855 = ~n1853 & ~n1854;
  assign n1856 = ~n1852 & n1855;
  assign n1857 = ~n1851 & n1856;
  assign n1858 = n313 & ~n1857;
  assign n1859 = n265 & ~n1177;
  assign n1860 = n276 & ~n1193;
  assign n1861 = n287 & ~n1169;
  assign n1862 = n298 & ~n1185;
  assign n1863 = ~n1861 & ~n1862;
  assign n1864 = ~n1860 & n1863;
  assign n1865 = ~n1859 & n1864;
  assign n1866 = n358 & ~n1865;
  assign n1867 = n265 & ~n1321;
  assign n1868 = n276 & ~n1233;
  assign n1869 = n287 & ~n1313;
  assign n1870 = n298 & ~n1225;
  assign n1871 = ~n1869 & ~n1870;
  assign n1872 = ~n1868 & n1871;
  assign n1873 = ~n1867 & n1872;
  assign n1874 = n403 & ~n1873;
  assign n1875 = ~n1866 & ~n1874;
  assign n1876 = ~n1858 & n1875;
  assign n1877 = ~n1850 & n1876;
  assign n1878 = ~pi134  & ~n1877;
  assign n1879 = n265 & ~n1197;
  assign n1880 = n276 & ~n1297;
  assign n1881 = n287 & ~n1189;
  assign n1882 = n298 & ~n1289;
  assign n1883 = ~n1881 & ~n1882;
  assign n1884 = ~n1880 & n1883;
  assign n1885 = ~n1879 & n1884;
  assign n1886 = n403 & ~n1885;
  assign n1887 = n265 & ~n1281;
  assign n1888 = n276 & ~n1317;
  assign n1889 = n287 & ~n1273;
  assign n1890 = n298 & ~n1309;
  assign n1891 = ~n1889 & ~n1890;
  assign n1892 = ~n1888 & n1891;
  assign n1893 = ~n1887 & n1892;
  assign n1894 = n358 & ~n1893;
  assign n1895 = n276 & ~n1257;
  assign n1896 = n265 & ~n1301;
  assign n1897 = n287 & ~n1293;
  assign n1898 = n298 & ~n1249;
  assign n1899 = ~n1897 & ~n1898;
  assign n1900 = ~n1896 & n1899;
  assign n1901 = ~n1895 & n1900;
  assign n1902 = n313 & ~n1901;
  assign n1903 = n265 & ~n1261;
  assign n1904 = n276 & ~n1277;
  assign n1905 = n287 & ~n1253;
  assign n1906 = n298 & ~n1269;
  assign n1907 = ~n1905 & ~n1906;
  assign n1908 = ~n1904 & n1907;
  assign n1909 = ~n1903 & n1908;
  assign n1910 = n264 & ~n1909;
  assign n1911 = ~n1902 & ~n1910;
  assign n1912 = ~n1894 & n1911;
  assign n1913 = ~n1886 & n1912;
  assign n1914 = pi134  & ~n1913;
  assign po11  = n1878 | n1914;
  assign n1916 = n265 & ~n332;
  assign n1917 = n276 & ~n352;
  assign n1918 = n287 & ~n322;
  assign n1919 = ~n296 & n298;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = ~n1917 & n1920;
  assign n1922 = ~n1916 & n1921;
  assign n1923 = n264 & ~n1922;
  assign n1924 = n265 & ~n422;
  assign n1925 = n276 & ~n442;
  assign n1926 = n287 & ~n412;
  assign n1927 = n298 & ~n342;
  assign n1928 = ~n1926 & ~n1927;
  assign n1929 = ~n1925 & n1928;
  assign n1930 = ~n1924 & n1929;
  assign n1931 = n313 & ~n1930;
  assign n1932 = n265 & ~n285;
  assign n1933 = n276 & ~n307;
  assign n1934 = ~n274 & n287;
  assign n1935 = n298 & ~n387;
  assign n1936 = ~n1934 & ~n1935;
  assign n1937 = ~n1933 & n1936;
  assign n1938 = ~n1932 & n1937;
  assign n1939 = n358 & ~n1938;
  assign n1940 = n265 & ~n558;
  assign n1941 = n276 & ~n578;
  assign n1942 = n287 & ~n548;
  assign n1943 = n298 & ~n432;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = ~n1941 & n1944;
  assign n1946 = ~n1940 & n1945;
  assign n1947 = n403 & ~n1946;
  assign n1948 = ~n1939 & ~n1947;
  assign n1949 = ~n1931 & n1948;
  assign n1950 = ~n1923 & n1949;
  assign n1951 = ~pi134  & ~n1950;
  assign n1952 = n265 & ~n377;
  assign n1953 = n276 & ~n397;
  assign n1954 = n287 & ~n367;
  assign n1955 = n298 & ~n612;
  assign n1956 = ~n1954 & ~n1955;
  assign n1957 = ~n1953 & n1956;
  assign n1958 = ~n1952 & n1957;
  assign n1959 = n403 & ~n1958;
  assign n1960 = n265 & ~n470;
  assign n1961 = n276 & ~n490;
  assign n1962 = n287 & ~n460;
  assign n1963 = n298 & ~n568;
  assign n1964 = ~n1962 & ~n1963;
  assign n1965 = ~n1961 & n1964;
  assign n1966 = ~n1960 & n1965;
  assign n1967 = n358 & ~n1966;
  assign n1968 = n265 & ~n602;
  assign n1969 = n276 & ~n622;
  assign n1970 = n287 & ~n592;
  assign n1971 = n298 & ~n524;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = ~n1969 & n1972;
  assign n1974 = ~n1968 & n1973;
  assign n1975 = n313 & ~n1974;
  assign n1976 = n265 & ~n514;
  assign n1977 = n276 & ~n534;
  assign n1978 = n287 & ~n504;
  assign n1979 = n298 & ~n480;
  assign n1980 = ~n1978 & ~n1979;
  assign n1981 = ~n1977 & n1980;
  assign n1982 = ~n1976 & n1981;
  assign n1983 = n264 & ~n1982;
  assign n1984 = ~n1975 & ~n1983;
  assign n1985 = ~n1967 & n1984;
  assign n1986 = ~n1959 & n1985;
  assign n1987 = pi134  & ~n1986;
  assign po12  = n1951 | n1987;
  assign n1989 = n265 & ~n695;
  assign n1990 = n276 & ~n715;
  assign n1991 = n287 & ~n685;
  assign n1992 = n298 & ~n661;
  assign n1993 = ~n1991 & ~n1992;
  assign n1994 = ~n1990 & n1993;
  assign n1995 = ~n1989 & n1994;
  assign n1996 = n264 & ~n1995;
  assign n1997 = n265 & ~n783;
  assign n1998 = n276 & ~n803;
  assign n1999 = n287 & ~n773;
  assign n2000 = n298 & ~n705;
  assign n2001 = ~n1999 & ~n2000;
  assign n2002 = ~n1998 & n2001;
  assign n2003 = ~n1997 & n2002;
  assign n2004 = n313 & ~n2003;
  assign n2005 = n265 & ~n651;
  assign n2006 = n276 & ~n671;
  assign n2007 = n287 & ~n641;
  assign n2008 = n298 & ~n749;
  assign n2009 = ~n2007 & ~n2008;
  assign n2010 = ~n2006 & n2009;
  assign n2011 = ~n2005 & n2010;
  assign n2012 = n358 & ~n2011;
  assign n2013 = n265 & ~n831;
  assign n2014 = n276 & ~n851;
  assign n2015 = n287 & ~n821;
  assign n2016 = n298 & ~n793;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = ~n2014 & n2017;
  assign n2019 = ~n2013 & n2018;
  assign n2020 = n403 & ~n2019;
  assign n2021 = ~n2012 & ~n2020;
  assign n2022 = ~n2004 & n2021;
  assign n2023 = ~n1996 & n2022;
  assign n2024 = ~pi134  & ~n2023;
  assign n2025 = n265 & ~n739;
  assign n2026 = n276 & ~n759;
  assign n2027 = n287 & ~n729;
  assign n2028 = n298 & ~n929;
  assign n2029 = ~n2027 & ~n2028;
  assign n2030 = ~n2026 & n2029;
  assign n2031 = ~n2025 & n2030;
  assign n2032 = n403 & ~n2031;
  assign n2033 = n265 & ~n875;
  assign n2034 = n276 & ~n895;
  assign n2035 = n287 & ~n865;
  assign n2036 = n298 & ~n841;
  assign n2037 = ~n2035 & ~n2036;
  assign n2038 = ~n2034 & n2037;
  assign n2039 = ~n2033 & n2038;
  assign n2040 = n358 & ~n2039;
  assign n2041 = n265 & ~n919;
  assign n2042 = n276 & ~n939;
  assign n2043 = n287 & ~n909;
  assign n2044 = n298 & ~n973;
  assign n2045 = ~n2043 & ~n2044;
  assign n2046 = ~n2042 & n2045;
  assign n2047 = ~n2041 & n2046;
  assign n2048 = n313 & ~n2047;
  assign n2049 = n265 & ~n963;
  assign n2050 = n276 & ~n983;
  assign n2051 = n287 & ~n953;
  assign n2052 = n298 & ~n885;
  assign n2053 = ~n2051 & ~n2052;
  assign n2054 = ~n2050 & n2053;
  assign n2055 = ~n2049 & n2054;
  assign n2056 = n264 & ~n2055;
  assign n2057 = ~n2048 & ~n2056;
  assign n2058 = ~n2040 & n2057;
  assign n2059 = ~n2032 & n2058;
  assign n2060 = pi134  & ~n2059;
  assign po13  = n2024 | n2060;
  assign n2062 = n265 & ~n1020;
  assign n2063 = n276 & ~n1028;
  assign n2064 = n287 & ~n1016;
  assign n2065 = n298 & ~n1004;
  assign n2066 = ~n2064 & ~n2065;
  assign n2067 = ~n2063 & n2066;
  assign n2068 = ~n2062 & n2067;
  assign n2069 = n264 & ~n2068;
  assign n2070 = n265 & ~n1060;
  assign n2071 = n276 & ~n1068;
  assign n2072 = n287 & ~n1056;
  assign n2073 = n298 & ~n1024;
  assign n2074 = ~n2072 & ~n2073;
  assign n2075 = ~n2071 & n2074;
  assign n2076 = ~n2070 & n2075;
  assign n2077 = n313 & ~n2076;
  assign n2078 = n265 & ~n1000;
  assign n2079 = n276 & ~n1008;
  assign n2080 = n287 & ~n996;
  assign n2081 = n298 & ~n1044;
  assign n2082 = ~n2080 & ~n2081;
  assign n2083 = ~n2079 & n2082;
  assign n2084 = ~n2078 & n2083;
  assign n2085 = n358 & ~n2084;
  assign n2086 = n265 & ~n1084;
  assign n2087 = n276 & ~n1092;
  assign n2088 = n287 & ~n1080;
  assign n2089 = n298 & ~n1064;
  assign n2090 = ~n2088 & ~n2089;
  assign n2091 = ~n2087 & n2090;
  assign n2092 = ~n2086 & n2091;
  assign n2093 = n403 & ~n2092;
  assign n2094 = ~n2085 & ~n2093;
  assign n2095 = ~n2077 & n2094;
  assign n2096 = ~n2069 & n2095;
  assign n2097 = ~pi134  & ~n2096;
  assign n2098 = n265 & ~n1040;
  assign n2099 = n276 & ~n1048;
  assign n2100 = n287 & ~n1036;
  assign n2101 = n298 & ~n1128;
  assign n2102 = ~n2100 & ~n2101;
  assign n2103 = ~n2099 & n2102;
  assign n2104 = ~n2098 & n2103;
  assign n2105 = n403 & ~n2104;
  assign n2106 = n265 & ~n1104;
  assign n2107 = n276 & ~n1112;
  assign n2108 = n287 & ~n1100;
  assign n2109 = n298 & ~n1088;
  assign n2110 = ~n2108 & ~n2109;
  assign n2111 = ~n2107 & n2110;
  assign n2112 = ~n2106 & n2111;
  assign n2113 = n358 & ~n2112;
  assign n2114 = n265 & ~n1124;
  assign n2115 = n276 & ~n1132;
  assign n2116 = n287 & ~n1120;
  assign n2117 = n298 & ~n1148;
  assign n2118 = ~n2116 & ~n2117;
  assign n2119 = ~n2115 & n2118;
  assign n2120 = ~n2114 & n2119;
  assign n2121 = n313 & ~n2120;
  assign n2122 = n265 & ~n1144;
  assign n2123 = n276 & ~n1152;
  assign n2124 = n287 & ~n1140;
  assign n2125 = n298 & ~n1108;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = ~n2123 & n2126;
  assign n2128 = ~n2122 & n2127;
  assign n2129 = n264 & ~n2128;
  assign n2130 = ~n2121 & ~n2129;
  assign n2131 = ~n2113 & n2130;
  assign n2132 = ~n2105 & n2131;
  assign n2133 = pi134  & ~n2132;
  assign po14  = n2097 | n2133;
  assign n2135 = n265 & ~n1209;
  assign n2136 = n276 & ~n1217;
  assign n2137 = n287 & ~n1205;
  assign n2138 = n298 & ~n1173;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140 = ~n2136 & n2139;
  assign n2141 = ~n2135 & n2140;
  assign n2142 = n264 & ~n2141;
  assign n2143 = n265 & ~n1229;
  assign n2144 = n276 & ~n1237;
  assign n2145 = n287 & ~n1225;
  assign n2146 = n298 & ~n1213;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = ~n2144 & n2147;
  assign n2149 = ~n2143 & n2148;
  assign n2150 = n313 & ~n2149;
  assign n2151 = n265 & ~n1169;
  assign n2152 = n276 & ~n1177;
  assign n2153 = n287 & ~n1165;
  assign n2154 = n298 & ~n1193;
  assign n2155 = ~n2153 & ~n2154;
  assign n2156 = ~n2152 & n2155;
  assign n2157 = ~n2151 & n2156;
  assign n2158 = n358 & ~n2157;
  assign n2159 = n265 & ~n1313;
  assign n2160 = n276 & ~n1321;
  assign n2161 = n287 & ~n1309;
  assign n2162 = n298 & ~n1233;
  assign n2163 = ~n2161 & ~n2162;
  assign n2164 = ~n2160 & n2163;
  assign n2165 = ~n2159 & n2164;
  assign n2166 = n403 & ~n2165;
  assign n2167 = ~n2158 & ~n2166;
  assign n2168 = ~n2150 & n2167;
  assign n2169 = ~n2142 & n2168;
  assign n2170 = ~pi134  & ~n2169;
  assign n2171 = n265 & ~n1189;
  assign n2172 = n276 & ~n1197;
  assign n2173 = n287 & ~n1185;
  assign n2174 = n298 & ~n1297;
  assign n2175 = ~n2173 & ~n2174;
  assign n2176 = ~n2172 & n2175;
  assign n2177 = ~n2171 & n2176;
  assign n2178 = n403 & ~n2177;
  assign n2179 = n265 & ~n1273;
  assign n2180 = n276 & ~n1281;
  assign n2181 = n287 & ~n1269;
  assign n2182 = n298 & ~n1317;
  assign n2183 = ~n2181 & ~n2182;
  assign n2184 = ~n2180 & n2183;
  assign n2185 = ~n2179 & n2184;
  assign n2186 = n358 & ~n2185;
  assign n2187 = n265 & ~n1293;
  assign n2188 = n276 & ~n1301;
  assign n2189 = n287 & ~n1289;
  assign n2190 = n298 & ~n1257;
  assign n2191 = ~n2189 & ~n2190;
  assign n2192 = ~n2188 & n2191;
  assign n2193 = ~n2187 & n2192;
  assign n2194 = n313 & ~n2193;
  assign n2195 = n265 & ~n1253;
  assign n2196 = n276 & ~n1261;
  assign n2197 = n287 & ~n1249;
  assign n2198 = n298 & ~n1277;
  assign n2199 = ~n2197 & ~n2198;
  assign n2200 = ~n2196 & n2199;
  assign n2201 = ~n2195 & n2200;
  assign n2202 = n264 & ~n2201;
  assign n2203 = ~n2194 & ~n2202;
  assign n2204 = ~n2186 & n2203;
  assign n2205 = ~n2178 & n2204;
  assign n2206 = pi134  & ~n2205;
  assign po15  = n2170 | n2206;
  assign n2208 = n264 & ~n356;
  assign n2209 = n313 & ~n446;
  assign n2210 = ~n311 & n358;
  assign n2211 = n403 & ~n582;
  assign n2212 = ~n2210 & ~n2211;
  assign n2213 = ~n2209 & n2212;
  assign n2214 = ~n2208 & n2213;
  assign n2215 = ~pi134  & ~n2214;
  assign n2216 = n358 & ~n494;
  assign n2217 = n264 & ~n538;
  assign n2218 = ~n401 & n403;
  assign n2219 = n313 & ~n626;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = ~n2217 & n2220;
  assign n2222 = ~n2216 & n2221;
  assign n2223 = pi134  & ~n2222;
  assign po16  = n2215 | n2223;
  assign n2225 = n264 & ~n719;
  assign n2226 = n313 & ~n807;
  assign n2227 = n358 & ~n675;
  assign n2228 = n403 & ~n855;
  assign n2229 = ~n2227 & ~n2228;
  assign n2230 = ~n2226 & n2229;
  assign n2231 = ~n2225 & n2230;
  assign n2232 = ~pi134  & ~n2231;
  assign n2233 = n403 & ~n763;
  assign n2234 = n358 & ~n899;
  assign n2235 = n313 & ~n943;
  assign n2236 = n264 & ~n987;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = ~n2234 & n2237;
  assign n2239 = ~n2233 & n2238;
  assign n2240 = pi134  & ~n2239;
  assign po17  = n2232 | n2240;
  assign n2242 = n264 & ~n1032;
  assign n2243 = n313 & ~n1072;
  assign n2244 = n358 & ~n1012;
  assign n2245 = n403 & ~n1096;
  assign n2246 = ~n2244 & ~n2245;
  assign n2247 = ~n2243 & n2246;
  assign n2248 = ~n2242 & n2247;
  assign n2249 = ~pi134  & ~n2248;
  assign n2250 = n403 & ~n1052;
  assign n2251 = n358 & ~n1116;
  assign n2252 = n313 & ~n1136;
  assign n2253 = n264 & ~n1156;
  assign n2254 = ~n2252 & ~n2253;
  assign n2255 = ~n2251 & n2254;
  assign n2256 = ~n2250 & n2255;
  assign n2257 = pi134  & ~n2256;
  assign po18  = n2249 | n2257;
  assign n2259 = n358 & ~n1181;
  assign n2260 = n403 & ~n1325;
  assign n2261 = n264 & ~n1221;
  assign n2262 = n313 & ~n1241;
  assign n2263 = ~n2261 & ~n2262;
  assign n2264 = ~n2260 & n2263;
  assign n2265 = ~n2259 & n2264;
  assign n2266 = ~pi134  & ~n2265;
  assign n2267 = n403 & ~n1201;
  assign n2268 = n264 & ~n1265;
  assign n2269 = n313 & ~n1305;
  assign n2270 = n358 & ~n1285;
  assign n2271 = ~n2269 & ~n2270;
  assign n2272 = ~n2268 & n2271;
  assign n2273 = ~n2267 & n2272;
  assign n2274 = pi134  & ~n2273;
  assign po19  = n2266 | n2274;
  assign n2276 = n264 & ~n1346;
  assign n2277 = n313 & ~n1362;
  assign n2278 = n358 & ~n1338;
  assign n2279 = n403 & ~n1382;
  assign n2280 = ~n2278 & ~n2279;
  assign n2281 = ~n2277 & n2280;
  assign n2282 = ~n2276 & n2281;
  assign n2283 = ~pi134  & ~n2282;
  assign n2284 = n264 & ~n1390;
  assign n2285 = n313 & ~n1374;
  assign n2286 = n403 & ~n1354;
  assign n2287 = n358 & ~n1398;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = ~n2285 & n2288;
  assign n2290 = ~n2284 & n2289;
  assign n2291 = pi134  & ~n2290;
  assign po20  = n2283 | n2291;
  assign n2293 = n264 & ~n1419;
  assign n2294 = n313 & ~n1435;
  assign n2295 = n358 & ~n1411;
  assign n2296 = n403 & ~n1455;
  assign n2297 = ~n2295 & ~n2296;
  assign n2298 = ~n2294 & n2297;
  assign n2299 = ~n2293 & n2298;
  assign n2300 = ~pi134  & ~n2299;
  assign n2301 = n264 & ~n1463;
  assign n2302 = n313 & ~n1447;
  assign n2303 = n403 & ~n1427;
  assign n2304 = n358 & ~n1471;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = ~n2302 & n2305;
  assign n2307 = ~n2301 & n2306;
  assign n2308 = pi134  & ~n2307;
  assign po21  = n2300 | n2308;
  assign n2310 = n264 & ~n1492;
  assign n2311 = n313 & ~n1508;
  assign n2312 = n358 & ~n1484;
  assign n2313 = n403 & ~n1528;
  assign n2314 = ~n2312 & ~n2313;
  assign n2315 = ~n2311 & n2314;
  assign n2316 = ~n2310 & n2315;
  assign n2317 = ~pi134  & ~n2316;
  assign n2318 = n264 & ~n1536;
  assign n2319 = n313 & ~n1520;
  assign n2320 = n403 & ~n1500;
  assign n2321 = n358 & ~n1544;
  assign n2322 = ~n2320 & ~n2321;
  assign n2323 = ~n2319 & n2322;
  assign n2324 = ~n2318 & n2323;
  assign n2325 = pi134  & ~n2324;
  assign po22  = n2317 | n2325;
  assign n2327 = n403 & ~n1601;
  assign n2328 = n264 & ~n1565;
  assign n2329 = n358 & ~n1557;
  assign n2330 = n313 & ~n1581;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = ~n2328 & n2331;
  assign n2333 = ~n2327 & n2332;
  assign n2334 = ~pi134  & ~n2333;
  assign n2335 = n313 & ~n1593;
  assign n2336 = n403 & ~n1573;
  assign n2337 = n264 & ~n1609;
  assign n2338 = n358 & ~n1617;
  assign n2339 = ~n2337 & ~n2338;
  assign n2340 = ~n2336 & n2339;
  assign n2341 = ~n2335 & n2340;
  assign n2342 = pi134  & ~n2341;
  assign po23  = n2334 | n2342;
  assign n2344 = n403 & ~n1674;
  assign n2345 = n264 & ~n1638;
  assign n2346 = n358 & ~n1630;
  assign n2347 = n313 & ~n1654;
  assign n2348 = ~n2346 & ~n2347;
  assign n2349 = ~n2345 & n2348;
  assign n2350 = ~n2344 & n2349;
  assign n2351 = ~pi134  & ~n2350;
  assign n2352 = n313 & ~n1666;
  assign n2353 = n403 & ~n1646;
  assign n2354 = n264 & ~n1682;
  assign n2355 = n358 & ~n1690;
  assign n2356 = ~n2354 & ~n2355;
  assign n2357 = ~n2353 & n2356;
  assign n2358 = ~n2352 & n2357;
  assign n2359 = pi134  & ~n2358;
  assign po24  = n2351 | n2359;
  assign n2361 = n403 & ~n1747;
  assign n2362 = n264 & ~n1711;
  assign n2363 = n358 & ~n1703;
  assign n2364 = n313 & ~n1727;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = ~n2362 & n2365;
  assign n2367 = ~n2361 & n2366;
  assign n2368 = ~pi134  & ~n2367;
  assign n2369 = n313 & ~n1739;
  assign n2370 = n403 & ~n1719;
  assign n2371 = n264 & ~n1755;
  assign n2372 = n358 & ~n1763;
  assign n2373 = ~n2371 & ~n2372;
  assign n2374 = ~n2370 & n2373;
  assign n2375 = ~n2369 & n2374;
  assign n2376 = pi134  & ~n2375;
  assign po25  = n2368 | n2376;
  assign n2378 = n264 & ~n1784;
  assign n2379 = n313 & ~n1800;
  assign n2380 = n358 & ~n1776;
  assign n2381 = n403 & ~n1820;
  assign n2382 = ~n2380 & ~n2381;
  assign n2383 = ~n2379 & n2382;
  assign n2384 = ~n2378 & n2383;
  assign n2385 = ~pi134  & ~n2384;
  assign n2386 = n313 & ~n1812;
  assign n2387 = n403 & ~n1792;
  assign n2388 = n264 & ~n1828;
  assign n2389 = n358 & ~n1836;
  assign n2390 = ~n2388 & ~n2389;
  assign n2391 = ~n2387 & n2390;
  assign n2392 = ~n2386 & n2391;
  assign n2393 = pi134  & ~n2392;
  assign po26  = n2385 | n2393;
  assign n2395 = n264 & ~n1857;
  assign n2396 = n313 & ~n1873;
  assign n2397 = n358 & ~n1849;
  assign n2398 = n403 & ~n1893;
  assign n2399 = ~n2397 & ~n2398;
  assign n2400 = ~n2396 & n2399;
  assign n2401 = ~n2395 & n2400;
  assign n2402 = ~pi134  & ~n2401;
  assign n2403 = n313 & ~n1885;
  assign n2404 = n403 & ~n1865;
  assign n2405 = n264 & ~n1901;
  assign n2406 = n358 & ~n1909;
  assign n2407 = ~n2405 & ~n2406;
  assign n2408 = ~n2404 & n2407;
  assign n2409 = ~n2403 & n2408;
  assign n2410 = pi134  & ~n2409;
  assign po27  = n2402 | n2410;
  assign n2412 = n264 & ~n1930;
  assign n2413 = n313 & ~n1946;
  assign n2414 = n358 & ~n1922;
  assign n2415 = n403 & ~n1966;
  assign n2416 = ~n2414 & ~n2415;
  assign n2417 = ~n2413 & n2416;
  assign n2418 = ~n2412 & n2417;
  assign n2419 = ~pi134  & ~n2418;
  assign n2420 = n313 & ~n1958;
  assign n2421 = n403 & ~n1938;
  assign n2422 = n264 & ~n1974;
  assign n2423 = n358 & ~n1982;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = ~n2421 & n2424;
  assign n2426 = ~n2420 & n2425;
  assign n2427 = pi134  & ~n2426;
  assign po28  = n2419 | n2427;
  assign n2429 = n264 & ~n2003;
  assign n2430 = n313 & ~n2019;
  assign n2431 = n358 & ~n1995;
  assign n2432 = n403 & ~n2039;
  assign n2433 = ~n2431 & ~n2432;
  assign n2434 = ~n2430 & n2433;
  assign n2435 = ~n2429 & n2434;
  assign n2436 = ~pi134  & ~n2435;
  assign n2437 = n313 & ~n2031;
  assign n2438 = n403 & ~n2011;
  assign n2439 = n264 & ~n2047;
  assign n2440 = n358 & ~n2055;
  assign n2441 = ~n2439 & ~n2440;
  assign n2442 = ~n2438 & n2441;
  assign n2443 = ~n2437 & n2442;
  assign n2444 = pi134  & ~n2443;
  assign po29  = n2436 | n2444;
  assign n2446 = n264 & ~n2076;
  assign n2447 = n313 & ~n2092;
  assign n2448 = n358 & ~n2068;
  assign n2449 = n403 & ~n2112;
  assign n2450 = ~n2448 & ~n2449;
  assign n2451 = ~n2447 & n2450;
  assign n2452 = ~n2446 & n2451;
  assign n2453 = ~pi134  & ~n2452;
  assign n2454 = n313 & ~n2104;
  assign n2455 = n403 & ~n2084;
  assign n2456 = n264 & ~n2120;
  assign n2457 = n358 & ~n2128;
  assign n2458 = ~n2456 & ~n2457;
  assign n2459 = ~n2455 & n2458;
  assign n2460 = ~n2454 & n2459;
  assign n2461 = pi134  & ~n2460;
  assign po30  = n2453 | n2461;
  assign n2463 = n264 & ~n2149;
  assign n2464 = n313 & ~n2165;
  assign n2465 = n358 & ~n2141;
  assign n2466 = n403 & ~n2185;
  assign n2467 = ~n2465 & ~n2466;
  assign n2468 = ~n2464 & n2467;
  assign n2469 = ~n2463 & n2468;
  assign n2470 = ~pi134  & ~n2469;
  assign n2471 = n313 & ~n2177;
  assign n2472 = n403 & ~n2157;
  assign n2473 = n264 & ~n2193;
  assign n2474 = n358 & ~n2201;
  assign n2475 = ~n2473 & ~n2474;
  assign n2476 = ~n2472 & n2475;
  assign n2477 = ~n2471 & n2476;
  assign n2478 = pi134  & ~n2477;
  assign po31  = n2470 | n2478;
  assign n2480 = n264 & ~n446;
  assign n2481 = n313 & ~n582;
  assign n2482 = ~n356 & n358;
  assign n2483 = n403 & ~n494;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = ~n2481 & n2484;
  assign n2486 = ~n2480 & n2485;
  assign n2487 = ~pi134  & ~n2486;
  assign n2488 = ~n311 & n403;
  assign n2489 = n358 & ~n538;
  assign n2490 = n313 & ~n401;
  assign n2491 = n264 & ~n626;
  assign n2492 = ~n2490 & ~n2491;
  assign n2493 = ~n2489 & n2492;
  assign n2494 = ~n2488 & n2493;
  assign n2495 = pi134  & ~n2494;
  assign po32  = n2487 | n2495;
  assign n2497 = n264 & ~n807;
  assign n2498 = n313 & ~n855;
  assign n2499 = n358 & ~n719;
  assign n2500 = n403 & ~n899;
  assign n2501 = ~n2499 & ~n2500;
  assign n2502 = ~n2498 & n2501;
  assign n2503 = ~n2497 & n2502;
  assign n2504 = ~pi134  & ~n2503;
  assign n2505 = n313 & ~n763;
  assign n2506 = n403 & ~n675;
  assign n2507 = n264 & ~n943;
  assign n2508 = n358 & ~n987;
  assign n2509 = ~n2507 & ~n2508;
  assign n2510 = ~n2506 & n2509;
  assign n2511 = ~n2505 & n2510;
  assign n2512 = pi134  & ~n2511;
  assign po33  = n2504 | n2512;
  assign n2514 = n264 & ~n1072;
  assign n2515 = n313 & ~n1096;
  assign n2516 = n358 & ~n1032;
  assign n2517 = n403 & ~n1116;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = ~n2515 & n2518;
  assign n2520 = ~n2514 & n2519;
  assign n2521 = ~pi134  & ~n2520;
  assign n2522 = n313 & ~n1052;
  assign n2523 = n403 & ~n1012;
  assign n2524 = n264 & ~n1136;
  assign n2525 = n358 & ~n1156;
  assign n2526 = ~n2524 & ~n2525;
  assign n2527 = ~n2523 & n2526;
  assign n2528 = ~n2522 & n2527;
  assign n2529 = pi134  & ~n2528;
  assign po34  = n2521 | n2529;
  assign n2531 = n403 & ~n1285;
  assign n2532 = n313 & ~n1325;
  assign n2533 = n358 & ~n1221;
  assign n2534 = n264 & ~n1241;
  assign n2535 = ~n2533 & ~n2534;
  assign n2536 = ~n2532 & n2535;
  assign n2537 = ~n2531 & n2536;
  assign n2538 = ~pi134  & ~n2537;
  assign n2539 = n403 & ~n1181;
  assign n2540 = n313 & ~n1201;
  assign n2541 = n264 & ~n1305;
  assign n2542 = n358 & ~n1265;
  assign n2543 = ~n2541 & ~n2542;
  assign n2544 = ~n2540 & n2543;
  assign n2545 = ~n2539 & n2544;
  assign n2546 = pi134  & ~n2545;
  assign po35  = n2538 | n2546;
  assign n2548 = n264 & ~n1362;
  assign n2549 = n313 & ~n1382;
  assign n2550 = n358 & ~n1346;
  assign n2551 = n403 & ~n1398;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = ~n2549 & n2552;
  assign n2554 = ~n2548 & n2553;
  assign n2555 = ~pi134  & ~n2554;
  assign n2556 = n403 & ~n1338;
  assign n2557 = n358 & ~n1390;
  assign n2558 = n313 & ~n1354;
  assign n2559 = n264 & ~n1374;
  assign n2560 = ~n2558 & ~n2559;
  assign n2561 = ~n2557 & n2560;
  assign n2562 = ~n2556 & n2561;
  assign n2563 = pi134  & ~n2562;
  assign po36  = n2555 | n2563;
  assign n2565 = n264 & ~n1435;
  assign n2566 = n313 & ~n1455;
  assign n2567 = n358 & ~n1419;
  assign n2568 = n403 & ~n1471;
  assign n2569 = ~n2567 & ~n2568;
  assign n2570 = ~n2566 & n2569;
  assign n2571 = ~n2565 & n2570;
  assign n2572 = ~pi134  & ~n2571;
  assign n2573 = n403 & ~n1411;
  assign n2574 = n358 & ~n1463;
  assign n2575 = n313 & ~n1427;
  assign n2576 = n264 & ~n1447;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = ~n2574 & n2577;
  assign n2579 = ~n2573 & n2578;
  assign n2580 = pi134  & ~n2579;
  assign po37  = n2572 | n2580;
  assign n2582 = n264 & ~n1508;
  assign n2583 = n313 & ~n1528;
  assign n2584 = n358 & ~n1492;
  assign n2585 = n403 & ~n1544;
  assign n2586 = ~n2584 & ~n2585;
  assign n2587 = ~n2583 & n2586;
  assign n2588 = ~n2582 & n2587;
  assign n2589 = ~pi134  & ~n2588;
  assign n2590 = n403 & ~n1484;
  assign n2591 = n358 & ~n1536;
  assign n2592 = n313 & ~n1500;
  assign n2593 = n264 & ~n1520;
  assign n2594 = ~n2592 & ~n2593;
  assign n2595 = ~n2591 & n2594;
  assign n2596 = ~n2590 & n2595;
  assign n2597 = pi134  & ~n2596;
  assign po38  = n2589 | n2597;
  assign n2599 = n403 & ~n1617;
  assign n2600 = n358 & ~n1565;
  assign n2601 = n313 & ~n1601;
  assign n2602 = n264 & ~n1581;
  assign n2603 = ~n2601 & ~n2602;
  assign n2604 = ~n2600 & n2603;
  assign n2605 = ~n2599 & n2604;
  assign n2606 = ~pi134  & ~n2605;
  assign n2607 = n264 & ~n1593;
  assign n2608 = n313 & ~n1573;
  assign n2609 = n358 & ~n1609;
  assign n2610 = n403 & ~n1557;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = ~n2608 & n2611;
  assign n2613 = ~n2607 & n2612;
  assign n2614 = pi134  & ~n2613;
  assign po39  = n2606 | n2614;
  assign n2616 = n403 & ~n1690;
  assign n2617 = n358 & ~n1638;
  assign n2618 = n313 & ~n1674;
  assign n2619 = n264 & ~n1654;
  assign n2620 = ~n2618 & ~n2619;
  assign n2621 = ~n2617 & n2620;
  assign n2622 = ~n2616 & n2621;
  assign n2623 = ~pi134  & ~n2622;
  assign n2624 = n264 & ~n1666;
  assign n2625 = n313 & ~n1646;
  assign n2626 = n358 & ~n1682;
  assign n2627 = n403 & ~n1630;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = ~n2625 & n2628;
  assign n2630 = ~n2624 & n2629;
  assign n2631 = pi134  & ~n2630;
  assign po40  = n2623 | n2631;
  assign n2633 = n403 & ~n1763;
  assign n2634 = n358 & ~n1711;
  assign n2635 = n313 & ~n1747;
  assign n2636 = n264 & ~n1727;
  assign n2637 = ~n2635 & ~n2636;
  assign n2638 = ~n2634 & n2637;
  assign n2639 = ~n2633 & n2638;
  assign n2640 = ~pi134  & ~n2639;
  assign n2641 = n264 & ~n1739;
  assign n2642 = n313 & ~n1719;
  assign n2643 = n358 & ~n1755;
  assign n2644 = n403 & ~n1703;
  assign n2645 = ~n2643 & ~n2644;
  assign n2646 = ~n2642 & n2645;
  assign n2647 = ~n2641 & n2646;
  assign n2648 = pi134  & ~n2647;
  assign po41  = n2640 | n2648;
  assign n2650 = n264 & ~n1800;
  assign n2651 = n313 & ~n1820;
  assign n2652 = n358 & ~n1784;
  assign n2653 = n403 & ~n1836;
  assign n2654 = ~n2652 & ~n2653;
  assign n2655 = ~n2651 & n2654;
  assign n2656 = ~n2650 & n2655;
  assign n2657 = ~pi134  & ~n2656;
  assign n2658 = n264 & ~n1812;
  assign n2659 = n313 & ~n1792;
  assign n2660 = n358 & ~n1828;
  assign n2661 = n403 & ~n1776;
  assign n2662 = ~n2660 & ~n2661;
  assign n2663 = ~n2659 & n2662;
  assign n2664 = ~n2658 & n2663;
  assign n2665 = pi134  & ~n2664;
  assign po42  = n2657 | n2665;
  assign n2667 = n264 & ~n1873;
  assign n2668 = n313 & ~n1893;
  assign n2669 = n358 & ~n1857;
  assign n2670 = n403 & ~n1909;
  assign n2671 = ~n2669 & ~n2670;
  assign n2672 = ~n2668 & n2671;
  assign n2673 = ~n2667 & n2672;
  assign n2674 = ~pi134  & ~n2673;
  assign n2675 = n264 & ~n1885;
  assign n2676 = n313 & ~n1865;
  assign n2677 = n358 & ~n1901;
  assign n2678 = n403 & ~n1849;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = ~n2676 & n2679;
  assign n2681 = ~n2675 & n2680;
  assign n2682 = pi134  & ~n2681;
  assign po43  = n2674 | n2682;
  assign n2684 = n264 & ~n1946;
  assign n2685 = n313 & ~n1966;
  assign n2686 = n358 & ~n1930;
  assign n2687 = n403 & ~n1982;
  assign n2688 = ~n2686 & ~n2687;
  assign n2689 = ~n2685 & n2688;
  assign n2690 = ~n2684 & n2689;
  assign n2691 = ~pi134  & ~n2690;
  assign n2692 = n264 & ~n1958;
  assign n2693 = n313 & ~n1938;
  assign n2694 = n358 & ~n1974;
  assign n2695 = n403 & ~n1922;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = ~n2693 & n2696;
  assign n2698 = ~n2692 & n2697;
  assign n2699 = pi134  & ~n2698;
  assign po44  = n2691 | n2699;
  assign n2701 = n264 & ~n2019;
  assign n2702 = n313 & ~n2039;
  assign n2703 = n358 & ~n2003;
  assign n2704 = n403 & ~n2055;
  assign n2705 = ~n2703 & ~n2704;
  assign n2706 = ~n2702 & n2705;
  assign n2707 = ~n2701 & n2706;
  assign n2708 = ~pi134  & ~n2707;
  assign n2709 = n264 & ~n2031;
  assign n2710 = n313 & ~n2011;
  assign n2711 = n358 & ~n2047;
  assign n2712 = n403 & ~n1995;
  assign n2713 = ~n2711 & ~n2712;
  assign n2714 = ~n2710 & n2713;
  assign n2715 = ~n2709 & n2714;
  assign n2716 = pi134  & ~n2715;
  assign po45  = n2708 | n2716;
  assign n2718 = n264 & ~n2092;
  assign n2719 = n313 & ~n2112;
  assign n2720 = n358 & ~n2076;
  assign n2721 = n403 & ~n2128;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = ~n2719 & n2722;
  assign n2724 = ~n2718 & n2723;
  assign n2725 = ~pi134  & ~n2724;
  assign n2726 = n264 & ~n2104;
  assign n2727 = n313 & ~n2084;
  assign n2728 = n358 & ~n2120;
  assign n2729 = n403 & ~n2068;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = ~n2727 & n2730;
  assign n2732 = ~n2726 & n2731;
  assign n2733 = pi134  & ~n2732;
  assign po46  = n2725 | n2733;
  assign n2735 = n264 & ~n2165;
  assign n2736 = n313 & ~n2185;
  assign n2737 = n358 & ~n2149;
  assign n2738 = n403 & ~n2201;
  assign n2739 = ~n2737 & ~n2738;
  assign n2740 = ~n2736 & n2739;
  assign n2741 = ~n2735 & n2740;
  assign n2742 = ~pi134  & ~n2741;
  assign n2743 = n264 & ~n2177;
  assign n2744 = n313 & ~n2157;
  assign n2745 = n358 & ~n2193;
  assign n2746 = n403 & ~n2141;
  assign n2747 = ~n2745 & ~n2746;
  assign n2748 = ~n2744 & n2747;
  assign n2749 = ~n2743 & n2748;
  assign n2750 = pi134  & ~n2749;
  assign po47  = n2742 | n2750;
  assign n2752 = n264 & ~n582;
  assign n2753 = n313 & ~n494;
  assign n2754 = n358 & ~n446;
  assign n2755 = n403 & ~n538;
  assign n2756 = ~n2754 & ~n2755;
  assign n2757 = ~n2753 & n2756;
  assign n2758 = ~n2752 & n2757;
  assign n2759 = ~pi134  & ~n2758;
  assign n2760 = ~n311 & n313;
  assign n2761 = ~n356 & n403;
  assign n2762 = n264 & ~n401;
  assign n2763 = n358 & ~n626;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = ~n2761 & n2764;
  assign n2766 = ~n2760 & n2765;
  assign n2767 = pi134  & ~n2766;
  assign po48  = n2759 | n2767;
  assign n2769 = n264 & ~n855;
  assign n2770 = n313 & ~n899;
  assign n2771 = n358 & ~n807;
  assign n2772 = n403 & ~n987;
  assign n2773 = ~n2771 & ~n2772;
  assign n2774 = ~n2770 & n2773;
  assign n2775 = ~n2769 & n2774;
  assign n2776 = ~pi134  & ~n2775;
  assign n2777 = n264 & ~n763;
  assign n2778 = n313 & ~n675;
  assign n2779 = n358 & ~n943;
  assign n2780 = n403 & ~n719;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = ~n2778 & n2781;
  assign n2783 = ~n2777 & n2782;
  assign n2784 = pi134  & ~n2783;
  assign po49  = n2776 | n2784;
  assign n2786 = n264 & ~n1096;
  assign n2787 = n313 & ~n1116;
  assign n2788 = n358 & ~n1072;
  assign n2789 = n403 & ~n1156;
  assign n2790 = ~n2788 & ~n2789;
  assign n2791 = ~n2787 & n2790;
  assign n2792 = ~n2786 & n2791;
  assign n2793 = ~pi134  & ~n2792;
  assign n2794 = n264 & ~n1052;
  assign n2795 = n313 & ~n1012;
  assign n2796 = n358 & ~n1136;
  assign n2797 = n403 & ~n1032;
  assign n2798 = ~n2796 & ~n2797;
  assign n2799 = ~n2795 & n2798;
  assign n2800 = ~n2794 & n2799;
  assign n2801 = pi134  & ~n2800;
  assign po50  = n2793 | n2801;
  assign n2803 = n313 & ~n1285;
  assign n2804 = n264 & ~n1325;
  assign n2805 = n403 & ~n1265;
  assign n2806 = n358 & ~n1241;
  assign n2807 = ~n2805 & ~n2806;
  assign n2808 = ~n2804 & n2807;
  assign n2809 = ~n2803 & n2808;
  assign n2810 = ~pi134  & ~n2809;
  assign n2811 = n403 & ~n1221;
  assign n2812 = n313 & ~n1181;
  assign n2813 = n358 & ~n1305;
  assign n2814 = n264 & ~n1201;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = ~n2812 & n2815;
  assign n2817 = ~n2811 & n2816;
  assign n2818 = pi134  & ~n2817;
  assign po51  = n2810 | n2818;
  assign n2820 = n358 & ~n1362;
  assign n2821 = n264 & ~n1382;
  assign n2822 = n403 & ~n1390;
  assign n2823 = n313 & ~n1398;
  assign n2824 = ~n2822 & ~n2823;
  assign n2825 = ~n2821 & n2824;
  assign n2826 = ~n2820 & n2825;
  assign n2827 = ~pi134  & ~n2826;
  assign n2828 = n313 & ~n1338;
  assign n2829 = n358 & ~n1374;
  assign n2830 = n264 & ~n1354;
  assign n2831 = n403 & ~n1346;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = ~n2829 & n2832;
  assign n2834 = ~n2828 & n2833;
  assign n2835 = pi134  & ~n2834;
  assign po52  = n2827 | n2835;
  assign n2837 = n358 & ~n1435;
  assign n2838 = n264 & ~n1455;
  assign n2839 = n403 & ~n1463;
  assign n2840 = n313 & ~n1471;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = ~n2838 & n2841;
  assign n2843 = ~n2837 & n2842;
  assign n2844 = ~pi134  & ~n2843;
  assign n2845 = n313 & ~n1411;
  assign n2846 = n358 & ~n1447;
  assign n2847 = n264 & ~n1427;
  assign n2848 = n403 & ~n1419;
  assign n2849 = ~n2847 & ~n2848;
  assign n2850 = ~n2846 & n2849;
  assign n2851 = ~n2845 & n2850;
  assign n2852 = pi134  & ~n2851;
  assign po53  = n2844 | n2852;
  assign n2854 = n358 & ~n1508;
  assign n2855 = n264 & ~n1528;
  assign n2856 = n403 & ~n1536;
  assign n2857 = n313 & ~n1544;
  assign n2858 = ~n2856 & ~n2857;
  assign n2859 = ~n2855 & n2858;
  assign n2860 = ~n2854 & n2859;
  assign n2861 = ~pi134  & ~n2860;
  assign n2862 = n313 & ~n1484;
  assign n2863 = n358 & ~n1520;
  assign n2864 = n264 & ~n1500;
  assign n2865 = n403 & ~n1492;
  assign n2866 = ~n2864 & ~n2865;
  assign n2867 = ~n2863 & n2866;
  assign n2868 = ~n2862 & n2867;
  assign n2869 = pi134  & ~n2868;
  assign po54  = n2861 | n2869;
  assign n2871 = n264 & ~n1601;
  assign n2872 = n313 & ~n1617;
  assign n2873 = n403 & ~n1609;
  assign n2874 = n358 & ~n1581;
  assign n2875 = ~n2873 & ~n2874;
  assign n2876 = ~n2872 & n2875;
  assign n2877 = ~n2871 & n2876;
  assign n2878 = ~pi134  & ~n2877;
  assign n2879 = n264 & ~n1573;
  assign n2880 = n313 & ~n1557;
  assign n2881 = n358 & ~n1593;
  assign n2882 = n403 & ~n1565;
  assign n2883 = ~n2881 & ~n2882;
  assign n2884 = ~n2880 & n2883;
  assign n2885 = ~n2879 & n2884;
  assign n2886 = pi134  & ~n2885;
  assign po55  = n2878 | n2886;
  assign n2888 = n264 & ~n1674;
  assign n2889 = n313 & ~n1690;
  assign n2890 = n403 & ~n1682;
  assign n2891 = n358 & ~n1654;
  assign n2892 = ~n2890 & ~n2891;
  assign n2893 = ~n2889 & n2892;
  assign n2894 = ~n2888 & n2893;
  assign n2895 = ~pi134  & ~n2894;
  assign n2896 = n264 & ~n1646;
  assign n2897 = n313 & ~n1630;
  assign n2898 = n358 & ~n1666;
  assign n2899 = n403 & ~n1638;
  assign n2900 = ~n2898 & ~n2899;
  assign n2901 = ~n2897 & n2900;
  assign n2902 = ~n2896 & n2901;
  assign n2903 = pi134  & ~n2902;
  assign po56  = n2895 | n2903;
  assign n2905 = n264 & ~n1747;
  assign n2906 = n313 & ~n1763;
  assign n2907 = n403 & ~n1755;
  assign n2908 = n358 & ~n1727;
  assign n2909 = ~n2907 & ~n2908;
  assign n2910 = ~n2906 & n2909;
  assign n2911 = ~n2905 & n2910;
  assign n2912 = ~pi134  & ~n2911;
  assign n2913 = n264 & ~n1719;
  assign n2914 = n313 & ~n1703;
  assign n2915 = n358 & ~n1739;
  assign n2916 = n403 & ~n1711;
  assign n2917 = ~n2915 & ~n2916;
  assign n2918 = ~n2914 & n2917;
  assign n2919 = ~n2913 & n2918;
  assign n2920 = pi134  & ~n2919;
  assign po57  = n2912 | n2920;
  assign n2922 = n358 & ~n1800;
  assign n2923 = n264 & ~n1820;
  assign n2924 = n403 & ~n1828;
  assign n2925 = n313 & ~n1836;
  assign n2926 = ~n2924 & ~n2925;
  assign n2927 = ~n2923 & n2926;
  assign n2928 = ~n2922 & n2927;
  assign n2929 = ~pi134  & ~n2928;
  assign n2930 = n264 & ~n1792;
  assign n2931 = n313 & ~n1776;
  assign n2932 = n358 & ~n1812;
  assign n2933 = n403 & ~n1784;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = ~n2931 & n2934;
  assign n2936 = ~n2930 & n2935;
  assign n2937 = pi134  & ~n2936;
  assign po58  = n2929 | n2937;
  assign n2939 = n358 & ~n1873;
  assign n2940 = n264 & ~n1893;
  assign n2941 = n403 & ~n1901;
  assign n2942 = n313 & ~n1909;
  assign n2943 = ~n2941 & ~n2942;
  assign n2944 = ~n2940 & n2943;
  assign n2945 = ~n2939 & n2944;
  assign n2946 = ~pi134  & ~n2945;
  assign n2947 = n264 & ~n1865;
  assign n2948 = n313 & ~n1849;
  assign n2949 = n358 & ~n1885;
  assign n2950 = n403 & ~n1857;
  assign n2951 = ~n2949 & ~n2950;
  assign n2952 = ~n2948 & n2951;
  assign n2953 = ~n2947 & n2952;
  assign n2954 = pi134  & ~n2953;
  assign po59  = n2946 | n2954;
  assign n2956 = n358 & ~n1946;
  assign n2957 = n264 & ~n1966;
  assign n2958 = n403 & ~n1974;
  assign n2959 = n313 & ~n1982;
  assign n2960 = ~n2958 & ~n2959;
  assign n2961 = ~n2957 & n2960;
  assign n2962 = ~n2956 & n2961;
  assign n2963 = ~pi134  & ~n2962;
  assign n2964 = n264 & ~n1938;
  assign n2965 = n313 & ~n1922;
  assign n2966 = n358 & ~n1958;
  assign n2967 = n403 & ~n1930;
  assign n2968 = ~n2966 & ~n2967;
  assign n2969 = ~n2965 & n2968;
  assign n2970 = ~n2964 & n2969;
  assign n2971 = pi134  & ~n2970;
  assign po60  = n2963 | n2971;
  assign n2973 = n358 & ~n2019;
  assign n2974 = n264 & ~n2039;
  assign n2975 = n403 & ~n2047;
  assign n2976 = n313 & ~n2055;
  assign n2977 = ~n2975 & ~n2976;
  assign n2978 = ~n2974 & n2977;
  assign n2979 = ~n2973 & n2978;
  assign n2980 = ~pi134  & ~n2979;
  assign n2981 = n264 & ~n2011;
  assign n2982 = n313 & ~n1995;
  assign n2983 = n358 & ~n2031;
  assign n2984 = n403 & ~n2003;
  assign n2985 = ~n2983 & ~n2984;
  assign n2986 = ~n2982 & n2985;
  assign n2987 = ~n2981 & n2986;
  assign n2988 = pi134  & ~n2987;
  assign po61  = n2980 | n2988;
  assign n2990 = n358 & ~n2092;
  assign n2991 = n264 & ~n2112;
  assign n2992 = n403 & ~n2120;
  assign n2993 = n313 & ~n2128;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = ~n2991 & n2994;
  assign n2996 = ~n2990 & n2995;
  assign n2997 = ~pi134  & ~n2996;
  assign n2998 = n264 & ~n2084;
  assign n2999 = n313 & ~n2068;
  assign n3000 = n358 & ~n2104;
  assign n3001 = n403 & ~n2076;
  assign n3002 = ~n3000 & ~n3001;
  assign n3003 = ~n2999 & n3002;
  assign n3004 = ~n2998 & n3003;
  assign n3005 = pi134  & ~n3004;
  assign po62  = n2997 | n3005;
  assign n3007 = n358 & ~n2165;
  assign n3008 = n264 & ~n2185;
  assign n3009 = n403 & ~n2193;
  assign n3010 = n313 & ~n2201;
  assign n3011 = ~n3009 & ~n3010;
  assign n3012 = ~n3008 & n3011;
  assign n3013 = ~n3007 & n3012;
  assign n3014 = ~pi134  & ~n3013;
  assign n3015 = n264 & ~n2157;
  assign n3016 = n313 & ~n2141;
  assign n3017 = n358 & ~n2177;
  assign n3018 = n403 & ~n2149;
  assign n3019 = ~n3017 & ~n3018;
  assign n3020 = ~n3016 & n3019;
  assign n3021 = ~n3015 & n3020;
  assign n3022 = pi134  & ~n3021;
  assign po63  = n3014 | n3022;
  assign n3024 = ~pi134  & ~n630;
  assign n3025 = pi134  & ~n450;
  assign po64  = n3024 | n3025;
  assign n3027 = ~pi134  & ~n991;
  assign n3028 = pi134  & ~n811;
  assign po65  = n3027 | n3028;
  assign n3030 = ~pi134  & ~n1160;
  assign n3031 = pi134  & ~n1076;
  assign po66  = n3030 | n3031;
  assign n3033 = ~pi134  & ~n1329;
  assign n3034 = pi134  & ~n1245;
  assign po67  = n3033 | n3034;
  assign n3036 = ~pi134  & ~n1402;
  assign n3037 = pi134  & ~n1366;
  assign po68  = n3036 | n3037;
  assign n3039 = ~pi134  & ~n1475;
  assign n3040 = pi134  & ~n1439;
  assign po69  = n3039 | n3040;
  assign n3042 = ~pi134  & ~n1548;
  assign n3043 = pi134  & ~n1512;
  assign po70  = n3042 | n3043;
  assign n3045 = ~pi134  & ~n1621;
  assign n3046 = pi134  & ~n1585;
  assign po71  = n3045 | n3046;
  assign n3048 = ~pi134  & ~n1694;
  assign n3049 = pi134  & ~n1658;
  assign po72  = n3048 | n3049;
  assign n3051 = ~pi134  & ~n1767;
  assign n3052 = pi134  & ~n1731;
  assign po73  = n3051 | n3052;
  assign n3054 = ~pi134  & ~n1840;
  assign n3055 = pi134  & ~n1804;
  assign po74  = n3054 | n3055;
  assign n3057 = ~pi134  & ~n1913;
  assign n3058 = pi134  & ~n1877;
  assign po75  = n3057 | n3058;
  assign n3060 = ~pi134  & ~n1986;
  assign n3061 = pi134  & ~n1950;
  assign po76  = n3060 | n3061;
  assign n3063 = ~pi134  & ~n2059;
  assign n3064 = pi134  & ~n2023;
  assign po77  = n3063 | n3064;
  assign n3066 = ~pi134  & ~n2132;
  assign n3067 = pi134  & ~n2096;
  assign po78  = n3066 | n3067;
  assign n3069 = ~pi134  & ~n2205;
  assign n3070 = pi134  & ~n2169;
  assign po79  = n3069 | n3070;
  assign n3072 = ~pi134  & ~n2222;
  assign n3073 = pi134  & ~n2214;
  assign po80  = n3072 | n3073;
  assign n3075 = ~pi134  & ~n2239;
  assign n3076 = pi134  & ~n2231;
  assign po81  = n3075 | n3076;
  assign n3078 = ~pi134  & ~n2256;
  assign n3079 = pi134  & ~n2248;
  assign po82  = n3078 | n3079;
  assign n3081 = ~pi134  & ~n2273;
  assign n3082 = pi134  & ~n2265;
  assign po83  = n3081 | n3082;
  assign n3084 = ~pi134  & ~n2290;
  assign n3085 = pi134  & ~n2282;
  assign po84  = n3084 | n3085;
  assign n3087 = ~pi134  & ~n2307;
  assign n3088 = pi134  & ~n2299;
  assign po85  = n3087 | n3088;
  assign n3090 = ~pi134  & ~n2324;
  assign n3091 = pi134  & ~n2316;
  assign po86  = n3090 | n3091;
  assign n3093 = ~pi134  & ~n2341;
  assign n3094 = pi134  & ~n2333;
  assign po87  = n3093 | n3094;
  assign n3096 = ~pi134  & ~n2358;
  assign n3097 = pi134  & ~n2350;
  assign po88  = n3096 | n3097;
  assign n3099 = ~pi134  & ~n2375;
  assign n3100 = pi134  & ~n2367;
  assign po89  = n3099 | n3100;
  assign n3102 = ~pi134  & ~n2392;
  assign n3103 = pi134  & ~n2384;
  assign po90  = n3102 | n3103;
  assign n3105 = ~pi134  & ~n2409;
  assign n3106 = pi134  & ~n2401;
  assign po91  = n3105 | n3106;
  assign n3108 = ~pi134  & ~n2426;
  assign n3109 = pi134  & ~n2418;
  assign po92  = n3108 | n3109;
  assign n3111 = ~pi134  & ~n2443;
  assign n3112 = pi134  & ~n2435;
  assign po93  = n3111 | n3112;
  assign n3114 = ~pi134  & ~n2460;
  assign n3115 = pi134  & ~n2452;
  assign po94  = n3114 | n3115;
  assign n3117 = ~pi134  & ~n2477;
  assign n3118 = pi134  & ~n2469;
  assign po95  = n3117 | n3118;
  assign n3120 = ~pi134  & ~n2494;
  assign n3121 = pi134  & ~n2486;
  assign po96  = n3120 | n3121;
  assign n3123 = ~pi134  & ~n2511;
  assign n3124 = pi134  & ~n2503;
  assign po97  = n3123 | n3124;
  assign n3126 = ~pi134  & ~n2528;
  assign n3127 = pi134  & ~n2520;
  assign po98  = n3126 | n3127;
  assign n3129 = ~pi134  & ~n2545;
  assign n3130 = pi134  & ~n2537;
  assign po99  = n3129 | n3130;
  assign n3132 = ~pi134  & ~n2562;
  assign n3133 = pi134  & ~n2554;
  assign po100  = n3132 | n3133;
  assign n3135 = ~pi134  & ~n2579;
  assign n3136 = pi134  & ~n2571;
  assign po101  = n3135 | n3136;
  assign n3138 = ~pi134  & ~n2596;
  assign n3139 = pi134  & ~n2588;
  assign po102  = n3138 | n3139;
  assign n3141 = ~pi134  & ~n2613;
  assign n3142 = pi134  & ~n2605;
  assign po103  = n3141 | n3142;
  assign n3144 = ~pi134  & ~n2630;
  assign n3145 = pi134  & ~n2622;
  assign po104  = n3144 | n3145;
  assign n3147 = ~pi134  & ~n2647;
  assign n3148 = pi134  & ~n2639;
  assign po105  = n3147 | n3148;
  assign n3150 = ~pi134  & ~n2664;
  assign n3151 = pi134  & ~n2656;
  assign po106  = n3150 | n3151;
  assign n3153 = ~pi134  & ~n2681;
  assign n3154 = pi134  & ~n2673;
  assign po107  = n3153 | n3154;
  assign n3156 = ~pi134  & ~n2698;
  assign n3157 = pi134  & ~n2690;
  assign po108  = n3156 | n3157;
  assign n3159 = ~pi134  & ~n2715;
  assign n3160 = pi134  & ~n2707;
  assign po109  = n3159 | n3160;
  assign n3162 = ~pi134  & ~n2732;
  assign n3163 = pi134  & ~n2724;
  assign po110  = n3162 | n3163;
  assign n3165 = ~pi134  & ~n2749;
  assign n3166 = pi134  & ~n2741;
  assign po111  = n3165 | n3166;
  assign n3168 = ~pi134  & ~n2766;
  assign n3169 = pi134  & ~n2758;
  assign po112  = n3168 | n3169;
  assign n3171 = ~pi134  & ~n2783;
  assign n3172 = pi134  & ~n2775;
  assign po113  = n3171 | n3172;
  assign n3174 = ~pi134  & ~n2800;
  assign n3175 = pi134  & ~n2792;
  assign po114  = n3174 | n3175;
  assign n3177 = ~pi134  & ~n2817;
  assign n3178 = pi134  & ~n2809;
  assign po115  = n3177 | n3178;
  assign n3180 = ~pi134  & ~n2834;
  assign n3181 = pi134  & ~n2826;
  assign po116  = n3180 | n3181;
  assign n3183 = ~pi134  & ~n2851;
  assign n3184 = pi134  & ~n2843;
  assign po117  = n3183 | n3184;
  assign n3186 = ~pi134  & ~n2868;
  assign n3187 = pi134  & ~n2860;
  assign po118  = n3186 | n3187;
  assign n3189 = ~pi134  & ~n2885;
  assign n3190 = pi134  & ~n2877;
  assign po119  = n3189 | n3190;
  assign n3192 = ~pi134  & ~n2902;
  assign n3193 = pi134  & ~n2894;
  assign po120  = n3192 | n3193;
  assign n3195 = ~pi134  & ~n2919;
  assign n3196 = pi134  & ~n2911;
  assign po121  = n3195 | n3196;
  assign n3198 = ~pi134  & ~n2936;
  assign n3199 = pi134  & ~n2928;
  assign po122  = n3198 | n3199;
  assign n3201 = ~pi134  & ~n2953;
  assign n3202 = pi134  & ~n2945;
  assign po123  = n3201 | n3202;
  assign n3204 = ~pi134  & ~n2970;
  assign n3205 = pi134  & ~n2962;
  assign po124  = n3204 | n3205;
  assign n3207 = ~pi134  & ~n2987;
  assign n3208 = pi134  & ~n2979;
  assign po125  = n3207 | n3208;
  assign n3210 = ~pi134  & ~n3004;
  assign n3211 = pi134  & ~n2996;
  assign po126  = n3210 | n3211;
  assign n3213 = ~pi134  & ~n3021;
  assign n3214 = pi134  & ~n3013;
  assign po127  = n3213 | n3214;
endmodule
