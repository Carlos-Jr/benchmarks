module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411,
    n412, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n448, n449, n450,
    n451, n452, n453, n454, n455, n456, n457,
    n458, n459, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n476, n477, n478, n479, n480,
    n481, n482, n483, n485, n486, n487, n488,
    n489, n490, n491, n492, n494, n495, n496,
    n497, n498, n499, n500, n501, n503, n504,
    n505, n506, n507, n508, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n520,
    n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n532, n533, n534, n535,
    n536, n537, n538, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n562, n563, n564, n565,
    n566, n567, n569, n570, n571, n572, n573,
    n574, n575, n577, n578, n579, n580, n581,
    n582, n583, n585, n586, n587, n588, n589,
    n590, n591, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n619, n620,
    n621, n622, n623, n624, n625, n627, n628,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n694,
    n695, n696, n697, n698, n699, n700, n701,
    n702, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n786, n787, n788, n789,
    n790, n791, n793, n794, n795, n796, n797,
    n798, n800, n801, n802, n803, n804, n805,
    n807, n808, n809, n810, n811, n812, n814,
    n815, n816, n817, n818, n819, n821, n822,
    n823, n824, n825, n826, n828, n829, n830,
    n831, n832, n833, n835, n836, n837, n838,
    n839, n840, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n859, n860, n861,
    n862, n863, n864, n865, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883,
    n885, n886, n887, n888, n889, n890, n891,
    n892, n893, n894, n895, n896, n897, n898,
    n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958,
    n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n981, n982,
    n983, n984, n985, n986, n987, n988, n989,
    n990, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1019, n1020, n1021, n1023, n1024,
    n1025, n1027, n1028, n1029, n1030, n1031,
    n1033, n1036, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1103, n1104, n1105,
    n1107, n1108, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1120,
    n1121, n1122, n1123, n1125, n1126, n1127,
    n1128, n1130, n1131, n1132, n1133, n1135,
    n1136, n1137, n1138, n1139, n1141, n1142,
    n1143, n1145, n1146, n1147, n1148, n1150,
    n1151, n1152, n1153, n1155, n1156, n1157,
    n1158, n1160, n1161, n1162, n1163, n1165,
    n1166, n1167, n1169, n1170, n1171, n1173,
    n1174, n1175, n1177, n1178, n1179, n1181,
    n1182, n1183, n1185, n1186, n1187, n1189,
    n1190, n1191, n1192, n1193, n1195, n1196,
    n1197, n1199, n1200, n1201, n1203, n1204,
    n1205, n1207, n1208, n1209, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1230, n1231,
    n1232, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1242, n1243, n1244, n1246,
    n1247, n1248, n1250, n1251, n1252, n1253,
    n1254, n1256, n1257, n1258, n1260, n1261,
    n1262, n1264, n1265, n1266, n1268, n1269,
    n1270, n1272, n1273, n1274, n1276, n1277,
    n1278, n1279, n1280, n1281, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1291,
    n1292, n1293, n1295, n1296, n1297, n1299,
    n1300, n1301, n1303, n1304, n1305, n1307,
    n1308, n1309, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390,
    n1392, n1393, n1394, n1395, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1433, n1434, n1435, n1436,
    n1438, n1439, n1440, n1441, n1443, n1444,
    n1445, n1446, n1448, n1449, n1450, n1451,
    n1453, n1454, n1455, n1456, n1457, n1459,
    n1460, n1461, n1462, n1464, n1465, n1466,
    n1467, n1468, n1471, n1472, n1473, n1474,
    n1475, n1478, n1479, n1480, n1482, n1487,
    n1488, n1490;
  assign n291 = ~pi5 & ~pi22;
  assign n292 = ~pi9 & ~pi11;
  assign n293 = n291 & n292;
  assign n294 = ~pi4 & ~pi19;
  assign n295 = ~pi18 & n294;
  assign n296 = ~pi16 & n295;
  assign n297 = n293 & n296;
  assign n298 = ~pi17 & ~pi21;
  assign n299 = ~pi8 & n298;
  assign n300 = ~pi14 & n299;
  assign n301 = ~pi6 & ~pi12;
  assign n302 = ~pi7 & n301;
  assign n303 = ~pi13 & n302;
  assign n304 = n300 & n303;
  assign n305 = n297 & n304;
  assign n306 = pi54 & ~n305;
  assign n307 = ~pi0 & ~n306;
  assign n308 = n291 & ~n292;
  assign n309 = ~pi56 & n308;
  assign n310 = ~pi56 & ~n291;
  assign n311 = ~pi8 & ~pi21;
  assign n312 = ~pi7 & pi13;
  assign n313 = n311 & n312;
  assign n314 = ~pi7 & n311;
  assign n315 = pi7 & ~n311;
  assign n316 = ~n314 & ~n315;
  assign n317 = pi8 & pi21;
  assign n318 = ~pi13 & ~n317;
  assign n319 = n316 & n318;
  assign n320 = ~n313 & ~n319;
  assign n321 = ~pi14 & ~n320;
  assign n322 = ~pi13 & pi14;
  assign n323 = n314 & n322;
  assign n324 = ~n321 & ~n323;
  assign n325 = ~pi10 & ~n324;
  assign n326 = ~pi13 & ~pi14;
  assign n327 = pi10 & n326;
  assign n328 = n314 & n327;
  assign n329 = ~n325 & ~n328;
  assign n330 = n291 & ~n329;
  assign n331 = n296 & n330;
  assign n332 = ~pi17 & n331;
  assign n333 = n301 & n332;
  assign n334 = ~n310 & ~n333;
  assign n335 = n292 & ~n334;
  assign n336 = ~n309 & ~n335;
  assign n337 = pi54 & ~n336;
  assign n338 = ~n307 & ~n337;
  assign n339 = ~pi129 & ~n338;
  assign po15 = pi3 | ~n339;
  assign n341 = ~pi11 & ~pi12;
  assign n342 = n311 & n341;
  assign n343 = n296 & n342;
  assign n344 = ~pi7 & ~pi13;
  assign n345 = ~pi5 & ~pi6;
  assign n346 = n344 & n345;
  assign n347 = ~pi10 & ~pi22;
  assign n348 = n326 & n347;
  assign n349 = n346 & n348;
  assign n350 = n343 & n349;
  assign n351 = ~pi17 & pi54;
  assign n352 = ~n350 & n351;
  assign n353 = ~pi1 & ~n352;
  assign n354 = ~pi14 & pi54;
  assign n355 = ~pi8 & ~pi11;
  assign n356 = n298 & n355;
  assign n357 = ~pi5 & n301;
  assign n358 = pi5 & ~n301;
  assign n359 = ~n357 & ~n358;
  assign n360 = pi6 & pi12;
  assign n361 = ~pi7 & ~n360;
  assign n362 = n359 & n361;
  assign n363 = pi7 & n357;
  assign n364 = ~n362 & ~n363;
  assign n365 = ~pi13 & ~n364;
  assign n366 = n312 & n357;
  assign n367 = ~n365 & ~n366;
  assign n368 = ~pi9 & ~n367;
  assign n369 = n344 & n357;
  assign n370 = pi9 & n369;
  assign n371 = ~n368 & ~n370;
  assign n372 = n296 & ~n371;
  assign n373 = n356 & n372;
  assign n374 = n354 & n373;
  assign n375 = n347 & n374;
  assign n376 = ~n353 & ~n375;
  assign n377 = ~pi129 & ~n376;
  assign po16 = pi3 | ~n377;
  assign n379 = pi122 & pi127;
  assign n380 = ~pi43 & ~pi47;
  assign n381 = ~pi48 & n380;
  assign n382 = ~pi46 & ~pi50;
  assign n383 = ~pi41 & n382;
  assign n384 = n381 & n383;
  assign n385 = ~pi2 & ~pi45;
  assign n386 = ~pi24 & ~pi49;
  assign n387 = ~pi15 & n386;
  assign n388 = ~pi20 & n387;
  assign n389 = n385 & n388;
  assign n390 = n384 & n389;
  assign n391 = pi82 & ~n390;
  assign n392 = ~pi42 & ~pi44;
  assign n393 = ~pi38 & ~pi40;
  assign n394 = n392 & n393;
  assign n395 = pi82 & ~n394;
  assign n396 = ~n391 & ~n395;
  assign n397 = ~n379 & n396;
  assign n398 = ~pi65 & n397;
  assign n399 = ~pi47 & ~pi48;
  assign n400 = ~pi45 & n399;
  assign n401 = ~pi41 & ~pi46;
  assign n402 = ~pi43 & n401;
  assign n403 = n400 & n402;
  assign n404 = ~pi50 & n394;
  assign n405 = n386 & n404;
  assign n406 = n403 & n405;
  assign n407 = n388 & n406;
  assign n408 = pi82 & ~n407;
  assign n409 = ~pi82 & n379;
  assign n410 = ~n408 & ~n409;
  assign n411 = pi2 & ~n410;
  assign n412 = ~n398 & ~n411;
  assign po17 = ~pi129 & ~n412;
  assign n414 = ~pi9 & ~pi14;
  assign n415 = n347 & n414;
  assign n416 = n346 & n415;
  assign n417 = ~pi17 & n343;
  assign n418 = n416 & n417;
  assign n419 = ~pi61 & ~pi118;
  assign n420 = ~n418 & n419;
  assign n421 = pi0 & ~pi123;
  assign n422 = ~pi113 & n421;
  assign n423 = ~n420 & ~n422;
  assign po18 = ~pi129 & ~n423;
  assign n425 = ~pi9 & ~pi22;
  assign n426 = n327 & n425;
  assign n427 = n369 & n426;
  assign n428 = ~pi16 & pi54;
  assign n429 = n295 & n428;
  assign n430 = n356 & n429;
  assign n431 = n427 & n430;
  assign n432 = pi4 & ~pi54;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~pi129 & ~n433;
  assign po19 = ~pi3 & n434;
  assign n436 = pi5 & ~pi54;
  assign n437 = ~pi25 & ~pi29;
  assign n438 = pi28 & n437;
  assign n439 = n302 & n438;
  assign n440 = ~pi13 & n415;
  assign n441 = n439 & n440;
  assign n442 = ~pi5 & ~pi59;
  assign n443 = n430 & n442;
  assign n444 = n441 & n443;
  assign n445 = ~n436 & ~n444;
  assign n446 = ~pi129 & ~n445;
  assign po20 = ~pi3 & n446;
  assign n448 = pi6 & ~pi54;
  assign n449 = ~pi5 & ~pi7;
  assign n450 = pi25 & ~pi29;
  assign n451 = ~pi28 & n450;
  assign n452 = ~pi12 & n451;
  assign n453 = n449 & n452;
  assign n454 = n440 & n453;
  assign n455 = ~pi6 & ~pi59;
  assign n456 = n430 & n455;
  assign n457 = n454 & n456;
  assign n458 = ~n448 & ~n457;
  assign n459 = ~pi129 & ~n458;
  assign po21 = ~pi3 & n459;
  assign n461 = pi7 & ~pi54;
  assign n462 = ~pi7 & n294;
  assign n463 = n428 & n462;
  assign n464 = pi8 & ~pi18;
  assign n465 = n298 & n464;
  assign n466 = n463 & n465;
  assign n467 = ~pi6 & n341;
  assign n468 = ~pi9 & ~pi10;
  assign n469 = n326 & n468;
  assign n470 = n467 & n469;
  assign n471 = n291 & n470;
  assign n472 = n466 & n471;
  assign n473 = ~n461 & ~n472;
  assign n474 = ~pi129 & ~n473;
  assign po22 = ~pi3 & n474;
  assign n476 = pi8 & ~pi54;
  assign n477 = n369 & n415;
  assign n478 = n296 & n351;
  assign n479 = pi21 & n355;
  assign n480 = n478 & n479;
  assign n481 = n477 & n480;
  assign n482 = ~n476 & ~n481;
  assign n483 = ~pi129 & ~n482;
  assign po23 = ~pi3 & n483;
  assign n485 = pi9 & ~pi54;
  assign n486 = pi11 & ~pi12;
  assign n487 = n349 & n486;
  assign n488 = ~pi9 & n299;
  assign n489 = n429 & n488;
  assign n490 = n487 & n489;
  assign n491 = ~n485 & ~n490;
  assign n492 = ~pi129 & ~n491;
  assign po24 = ~pi3 & n492;
  assign n494 = pi10 & ~pi54;
  assign n495 = ~pi10 & n299;
  assign n496 = n429 & n495;
  assign n497 = pi14 & n293;
  assign n498 = n303 & n497;
  assign n499 = n496 & n498;
  assign n500 = ~n494 & ~n499;
  assign n501 = ~pi129 & ~n500;
  assign po25 = ~pi3 & n501;
  assign n503 = pi11 & ~pi54;
  assign n504 = pi22 & n469;
  assign n505 = n369 & n504;
  assign n506 = n430 & n505;
  assign n507 = ~n503 & ~n506;
  assign n508 = ~pi129 & ~n507;
  assign po26 = ~pi3 & n508;
  assign n510 = pi12 & ~pi54;
  assign n511 = ~pi12 & n294;
  assign n512 = n428 & n511;
  assign n513 = pi18 & n299;
  assign n514 = n512 & n513;
  assign n515 = ~pi11 & n416;
  assign n516 = n514 & n515;
  assign n517 = ~n510 & ~n516;
  assign n518 = ~pi129 & ~n517;
  assign po27 = ~pi3 & n518;
  assign n520 = pi13 & ~pi54;
  assign n521 = ~pi13 & ~pi59;
  assign n522 = n430 & n521;
  assign n523 = ~pi25 & ~pi28;
  assign n524 = ~pi7 & n523;
  assign n525 = n357 & n524;
  assign n526 = pi29 & n415;
  assign n527 = n525 & n526;
  assign n528 = n522 & n527;
  assign n529 = ~n520 & ~n528;
  assign n530 = ~pi129 & ~n529;
  assign po28 = ~pi3 & n530;
  assign n532 = pi14 & ~pi54;
  assign n533 = n300 & n429;
  assign n534 = ~pi10 & n293;
  assign n535 = n366 & n534;
  assign n536 = n533 & n535;
  assign n537 = ~n532 & ~n536;
  assign n538 = ~pi129 & ~n537;
  assign po29 = ~pi3 & n538;
  assign n540 = ~pi40 & n392;
  assign n541 = ~pi38 & ~pi50;
  assign n542 = ~pi46 & n541;
  assign n543 = n540 & n542;
  assign n544 = n403 & n543;
  assign n545 = n387 & n544;
  assign n546 = pi82 & ~n545;
  assign n547 = ~n379 & ~n546;
  assign n548 = ~pi70 & n547;
  assign n549 = pi15 & ~n406;
  assign n550 = n383 & n394;
  assign n551 = ~pi43 & n550;
  assign n552 = ~pi2 & ~pi20;
  assign n553 = n387 & ~n552;
  assign n554 = n551 & n553;
  assign n555 = n400 & n554;
  assign n556 = ~n549 & ~n555;
  assign n557 = pi82 & ~n556;
  assign n558 = pi15 & n409;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~n548 & n559;
  assign po30 = ~pi129 & ~n560;
  assign n562 = pi16 & ~pi54;
  assign n563 = pi6 & n365;
  assign n564 = n415 & n563;
  assign n565 = n430 & n564;
  assign n566 = ~n562 & ~n565;
  assign n567 = ~pi129 & ~n566;
  assign po31 = ~pi3 & n567;
  assign n569 = pi17 & ~pi54;
  assign n570 = n440 & n525;
  assign n571 = ~pi29 & pi59;
  assign n572 = n430 & n571;
  assign n573 = n570 & n572;
  assign n574 = ~n569 & ~n573;
  assign n575 = ~pi129 & ~n574;
  assign po32 = ~pi3 & n575;
  assign n577 = pi18 & ~pi54;
  assign n578 = pi16 & pi54;
  assign n579 = n295 & n578;
  assign n580 = n356 & n579;
  assign n581 = n477 & n580;
  assign n582 = ~n577 & ~n581;
  assign n583 = ~pi129 & ~n582;
  assign po33 = ~pi3 & n583;
  assign n585 = pi19 & ~pi54;
  assign n586 = ~pi11 & n311;
  assign n587 = pi17 & n586;
  assign n588 = n429 & n587;
  assign n589 = n477 & n588;
  assign n590 = ~n585 & ~n589;
  assign n591 = ~pi129 & ~n590;
  assign po34 = ~pi3 & n591;
  assign n593 = ~n379 & ~n408;
  assign n594 = ~pi71 & n593;
  assign n595 = ~pi24 & n403;
  assign n596 = ~pi15 & ~pi49;
  assign n597 = n404 & n596;
  assign n598 = n595 & n597;
  assign n599 = pi20 & ~n598;
  assign n600 = pi2 & n407;
  assign n601 = ~n599 & ~n600;
  assign n602 = pi82 & ~n601;
  assign n603 = pi20 & n409;
  assign n604 = ~n602 & ~n603;
  assign n605 = ~n594 & n604;
  assign po35 = ~pi129 & ~n605;
  assign n607 = pi21 & ~pi54;
  assign n608 = ~pi17 & ~pi18;
  assign n609 = n355 & n608;
  assign n610 = ~pi4 & ~pi16;
  assign n611 = ~pi21 & pi54;
  assign n612 = pi19 & n611;
  assign n613 = n610 & n612;
  assign n614 = n609 & n613;
  assign n615 = n477 & n614;
  assign n616 = ~n607 & ~n615;
  assign n617 = ~pi129 & ~n616;
  assign po36 = ~pi3 & n617;
  assign n619 = pi22 & ~pi54;
  assign n620 = ~pi22 & n299;
  assign n621 = n429 & n620;
  assign n622 = n362 & n470;
  assign n623 = n621 & n622;
  assign n624 = ~n619 & ~n623;
  assign n625 = ~pi129 & ~n624;
  assign po37 = ~pi3 & n625;
  assign n627 = ~pi23 & pi55;
  assign n628 = ~pi129 & ~n627;
  assign po38 = pi61 & n628;
  assign n630 = pi82 & ~n544;
  assign n631 = n552 & n596;
  assign n632 = pi82 & ~n631;
  assign n633 = n379 & ~n632;
  assign n634 = ~n630 & ~n633;
  assign n635 = ~pi24 & ~n634;
  assign n636 = n385 & n399;
  assign n637 = n631 & n636;
  assign n638 = n551 & n637;
  assign n639 = pi82 & ~n638;
  assign n640 = ~n379 & ~n639;
  assign n641 = pi63 & n640;
  assign n642 = pi24 & pi82;
  assign n643 = n404 & n642;
  assign n644 = n403 & n643;
  assign n645 = ~pi129 & ~n644;
  assign n646 = ~n641 & n645;
  assign po39 = ~n635 & n646;
  assign n648 = pi85 & pi116;
  assign n649 = pi85 & ~pi116;
  assign n650 = ~pi110 & ~n649;
  assign n651 = ~pi96 & n650;
  assign n652 = ~n648 & ~n651;
  assign n653 = pi100 & ~n652;
  assign n654 = pi25 & ~pi116;
  assign n655 = pi85 & n654;
  assign n656 = ~n653 & ~n655;
  assign n657 = ~pi26 & ~n656;
  assign n658 = ~pi95 & ~pi100;
  assign n659 = ~pi97 & n658;
  assign n660 = ~pi110 & ~n659;
  assign n661 = pi25 & ~n660;
  assign n662 = pi26 & pi116;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~pi39 & ~pi52;
  assign n665 = ~pi51 & n664;
  assign n666 = ~n663 & ~n665;
  assign n667 = pi26 & n654;
  assign n668 = ~n666 & ~n667;
  assign n669 = ~pi85 & ~n668;
  assign n670 = ~n657 & ~n669;
  assign n671 = ~pi27 & ~n670;
  assign n672 = pi116 & n665;
  assign n673 = ~n654 & ~n672;
  assign n674 = pi27 & ~n673;
  assign n675 = n661 & n665;
  assign n676 = ~n674 & ~n675;
  assign n677 = ~pi26 & ~pi85;
  assign n678 = ~n676 & n677;
  assign n679 = ~n671 & ~n678;
  assign n680 = ~pi53 & ~n679;
  assign n681 = pi53 & ~pi85;
  assign n682 = ~pi27 & n681;
  assign n683 = n654 & ~n667;
  assign n684 = n682 & n683;
  assign n685 = ~n680 & ~n684;
  assign n686 = ~pi58 & ~n685;
  assign n687 = ~pi27 & ~pi85;
  assign n688 = ~pi53 & pi58;
  assign n689 = n687 & n688;
  assign n690 = n683 & n689;
  assign n691 = ~n686 & ~n690;
  assign n692 = ~pi129 & ~n691;
  assign po40 = ~pi3 & n692;
  assign n694 = ~n652 & ~n662;
  assign n695 = pi100 & n694;
  assign n696 = ~pi85 & ~n672;
  assign n697 = pi26 & n696;
  assign n698 = ~n695 & ~n697;
  assign n699 = ~pi129 & ~n698;
  assign n700 = ~pi3 & n699;
  assign n701 = ~pi53 & ~pi58;
  assign n702 = ~pi27 & n701;
  assign po41 = n700 & n702;
  assign n704 = pi95 & ~pi96;
  assign n705 = pi27 & pi116;
  assign n706 = n650 & ~n705;
  assign n707 = n704 & n706;
  assign n708 = ~pi27 & n648;
  assign n709 = ~n707 & ~n708;
  assign n710 = ~pi100 & ~n709;
  assign n711 = pi27 & n696;
  assign n712 = ~n710 & ~n711;
  assign n713 = ~pi129 & ~n712;
  assign n714 = ~pi3 & n713;
  assign n715 = ~pi26 & n701;
  assign po42 = n714 & n715;
  assign n717 = ~pi26 & ~n665;
  assign n718 = ~pi27 & n665;
  assign n719 = ~n717 & ~n718;
  assign n720 = ~n660 & ~n719;
  assign n721 = pi26 & ~pi27;
  assign n722 = ~pi26 & pi27;
  assign n723 = ~n721 & ~n722;
  assign n724 = ~pi116 & ~n723;
  assign n725 = ~n720 & ~n724;
  assign n726 = pi28 & ~n725;
  assign n727 = ~pi26 & ~pi100;
  assign n728 = ~pi110 & n727;
  assign n729 = n704 & n728;
  assign n730 = n662 & n665;
  assign n731 = ~n729 & ~n730;
  assign n732 = ~pi27 & ~n731;
  assign n733 = n705 & n717;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~n726 & n734;
  assign n736 = ~pi85 & ~n735;
  assign n737 = pi28 & ~pi116;
  assign n738 = ~pi100 & pi116;
  assign n739 = ~n737 & ~n738;
  assign n740 = pi85 & ~n739;
  assign n741 = ~pi26 & ~pi27;
  assign n742 = n740 & n741;
  assign n743 = ~n736 & ~n742;
  assign n744 = ~pi53 & ~n743;
  assign n745 = ~pi27 & pi28;
  assign n746 = ~pi116 & n745;
  assign n747 = ~pi26 & n681;
  assign n748 = n746 & n747;
  assign n749 = ~n744 & ~n748;
  assign n750 = ~pi58 & ~n749;
  assign n751 = n677 & n688;
  assign n752 = n746 & n751;
  assign n753 = ~n750 & ~n752;
  assign n754 = ~pi129 & ~n753;
  assign po43 = ~pi3 & n754;
  assign n756 = pi58 & pi116;
  assign n757 = ~pi58 & ~pi110;
  assign n758 = ~pi96 & n757;
  assign n759 = n658 & n758;
  assign n760 = ~n756 & ~n759;
  assign n761 = ~pi53 & ~n760;
  assign n762 = pi97 & n761;
  assign n763 = pi53 & ~pi58;
  assign n764 = ~n688 & ~n763;
  assign n765 = ~pi116 & ~n764;
  assign n766 = ~n660 & n701;
  assign n767 = ~n765 & ~n766;
  assign n768 = pi29 & ~n767;
  assign n769 = ~n762 & ~n768;
  assign n770 = ~pi27 & ~n769;
  assign n771 = pi29 & ~pi116;
  assign n772 = pi27 & n771;
  assign n773 = n701 & n772;
  assign n774 = ~n770 & ~n773;
  assign n775 = ~pi85 & ~n774;
  assign n776 = pi85 & n702;
  assign n777 = n771 & n776;
  assign n778 = ~n775 & ~n777;
  assign n779 = ~pi26 & ~n778;
  assign n780 = ~pi85 & n701;
  assign n781 = n721 & n780;
  assign n782 = n771 & n781;
  assign n783 = ~n779 & ~n782;
  assign n784 = ~pi129 & ~n783;
  assign po44 = ~pi3 & n784;
  assign n786 = pi30 & ~pi109;
  assign n787 = pi60 & pi109;
  assign n788 = ~n786 & ~n787;
  assign n789 = ~pi106 & ~n788;
  assign n790 = pi88 & pi106;
  assign n791 = ~n789 & ~n790;
  assign po45 = ~pi129 & ~n791;
  assign n793 = pi89 & pi106;
  assign n794 = pi30 & pi109;
  assign n795 = pi31 & ~pi109;
  assign n796 = ~n794 & ~n795;
  assign n797 = ~pi106 & ~n796;
  assign n798 = ~n793 & ~n797;
  assign po46 = ~pi129 & ~n798;
  assign n800 = pi99 & pi106;
  assign n801 = pi31 & pi109;
  assign n802 = pi32 & ~pi109;
  assign n803 = ~n801 & ~n802;
  assign n804 = ~pi106 & ~n803;
  assign n805 = ~n800 & ~n804;
  assign po47 = ~pi129 & ~n805;
  assign n807 = pi90 & pi106;
  assign n808 = pi32 & pi109;
  assign n809 = pi33 & ~pi109;
  assign n810 = ~n808 & ~n809;
  assign n811 = ~pi106 & ~n810;
  assign n812 = ~n807 & ~n811;
  assign po48 = ~pi129 & ~n812;
  assign n814 = pi91 & pi106;
  assign n815 = pi33 & pi109;
  assign n816 = pi34 & ~pi109;
  assign n817 = ~n815 & ~n816;
  assign n818 = ~pi106 & ~n817;
  assign n819 = ~n814 & ~n818;
  assign po49 = ~pi129 & ~n819;
  assign n821 = pi92 & pi106;
  assign n822 = pi34 & pi109;
  assign n823 = pi35 & ~pi109;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~pi106 & ~n824;
  assign n826 = ~n821 & ~n825;
  assign po50 = ~pi129 & ~n826;
  assign n828 = pi98 & pi106;
  assign n829 = pi35 & pi109;
  assign n830 = pi36 & ~pi109;
  assign n831 = ~n829 & ~n830;
  assign n832 = ~pi106 & ~n831;
  assign n833 = ~n828 & ~n832;
  assign po51 = ~pi129 & ~n833;
  assign n835 = pi93 & pi106;
  assign n836 = pi36 & pi109;
  assign n837 = pi37 & ~pi109;
  assign n838 = ~n836 & ~n837;
  assign n839 = ~pi106 & ~n838;
  assign n840 = ~n835 & ~n839;
  assign po52 = ~pi129 & ~n840;
  assign n842 = pi82 & ~n540;
  assign n843 = n379 & ~n391;
  assign n844 = ~n842 & ~n843;
  assign n845 = ~pi38 & ~n844;
  assign n846 = ~pi45 & ~pi48;
  assign n847 = ~pi24 & n631;
  assign n848 = n846 & n847;
  assign n849 = n380 & n383;
  assign n850 = n540 & n849;
  assign n851 = n848 & n850;
  assign n852 = pi82 & ~n851;
  assign n853 = ~n379 & ~n852;
  assign n854 = pi74 & n853;
  assign n855 = n395 & n540;
  assign n856 = ~pi129 & ~n855;
  assign n857 = ~n854 & n856;
  assign po53 = ~n845 & n857;
  assign n859 = ~pi51 & pi109;
  assign n860 = n664 & n859;
  assign n861 = ~pi106 & ~n860;
  assign n862 = ~pi51 & ~pi52;
  assign n863 = pi109 & n862;
  assign n864 = pi39 & ~n863;
  assign n865 = n861 & ~n864;
  assign po54 = ~pi129 & ~n865;
  assign n867 = pi82 & ~n392;
  assign n868 = n381 & n389;
  assign n869 = n402 & n541;
  assign n870 = n868 & n869;
  assign n871 = pi82 & ~n870;
  assign n872 = n379 & ~n871;
  assign n873 = ~n867 & ~n872;
  assign n874 = ~pi40 & ~n873;
  assign n875 = n392 & n542;
  assign n876 = ~pi41 & n868;
  assign n877 = n875 & n876;
  assign n878 = pi82 & ~n877;
  assign n879 = ~n379 & ~n878;
  assign n880 = pi73 & n879;
  assign n881 = n842 & ~n867;
  assign n882 = ~pi129 & ~n881;
  assign n883 = ~n880 & n882;
  assign po55 = ~n874 & n883;
  assign n885 = pi82 & ~n543;
  assign n886 = pi82 & ~n868;
  assign n887 = n379 & ~n886;
  assign n888 = ~n885 & ~n887;
  assign n889 = ~pi41 & ~n888;
  assign n890 = n380 & n543;
  assign n891 = n848 & n890;
  assign n892 = pi82 & ~n891;
  assign n893 = ~n379 & ~n892;
  assign n894 = pi76 & n893;
  assign n895 = pi82 & ~n550;
  assign n896 = n543 & n895;
  assign n897 = ~pi129 & ~n896;
  assign n898 = ~n894 & n897;
  assign po56 = ~n889 & n898;
  assign n900 = pi44 & pi82;
  assign n901 = n382 & n393;
  assign n902 = n876 & n901;
  assign n903 = pi82 & ~n902;
  assign n904 = n379 & ~n903;
  assign n905 = ~n900 & ~n904;
  assign n906 = ~pi42 & ~n905;
  assign n907 = ~pi44 & n393;
  assign n908 = n849 & n907;
  assign n909 = n848 & n908;
  assign n910 = pi82 & ~n909;
  assign n911 = ~n379 & ~n910;
  assign n912 = pi72 & n911;
  assign n913 = ~pi44 & pi82;
  assign n914 = pi42 & n913;
  assign n915 = ~pi129 & ~n914;
  assign n916 = ~n912 & n915;
  assign po57 = ~n906 & n916;
  assign n918 = n388 & n636;
  assign n919 = pi82 & ~n918;
  assign n920 = n379 & ~n919;
  assign n921 = ~n895 & ~n920;
  assign n922 = ~pi43 & ~n921;
  assign n923 = ~n919 & n921;
  assign n924 = pi77 & n923;
  assign n925 = pi82 & ~n551;
  assign n926 = n550 & n925;
  assign n927 = ~pi129 & ~n926;
  assign n928 = ~n924 & n927;
  assign po58 = ~n922 & n928;
  assign n930 = ~pi40 & ~pi42;
  assign n931 = ~pi38 & n930;
  assign n932 = n849 & n931;
  assign n933 = n848 & n932;
  assign n934 = pi82 & ~n933;
  assign n935 = pi67 & ~n379;
  assign n936 = ~pi44 & n379;
  assign n937 = ~n935 & ~n936;
  assign n938 = ~n934 & ~n937;
  assign n939 = ~pi129 & ~n900;
  assign po59 = ~n938 & n939;
  assign n941 = pi82 & ~n847;
  assign n942 = n379 & ~n941;
  assign n943 = pi48 & n931;
  assign n944 = n913 & n943;
  assign n945 = pi47 & n930;
  assign n946 = n913 & n945;
  assign n947 = ~n925 & ~n946;
  assign n948 = ~n944 & n947;
  assign n949 = ~n942 & n948;
  assign n950 = ~pi45 & ~n949;
  assign n951 = n399 & n847;
  assign n952 = n551 & n951;
  assign n953 = pi82 & ~n952;
  assign n954 = ~n379 & ~n953;
  assign n955 = pi68 & n954;
  assign n956 = n630 & n948;
  assign n957 = ~pi129 & ~n956;
  assign n958 = ~n955 & n957;
  assign po60 = ~n950 & n958;
  assign n960 = pi82 & ~n404;
  assign n961 = pi82 & ~n876;
  assign n962 = n379 & ~n961;
  assign n963 = ~n960 & ~n962;
  assign n964 = ~pi46 & ~n963;
  assign n965 = ~n961 & n963;
  assign n966 = pi75 & n965;
  assign n967 = n404 & n885;
  assign n968 = ~pi129 & ~n967;
  assign n969 = ~n966 & n968;
  assign po61 = ~n964 & n969;
  assign n971 = pi82 & ~n848;
  assign n972 = n379 & ~n971;
  assign n973 = ~n925 & ~n972;
  assign n974 = ~pi47 & ~n973;
  assign n975 = ~n971 & n973;
  assign n976 = pi64 & n975;
  assign n977 = n869 & n946;
  assign n978 = ~pi129 & ~n977;
  assign n979 = ~n976 & n978;
  assign po62 = ~n974 & n979;
  assign n981 = ~pi47 & n389;
  assign n982 = n551 & n981;
  assign n983 = pi82 & ~n982;
  assign n984 = ~n379 & ~n983;
  assign n985 = pi62 & n984;
  assign n986 = n849 & n944;
  assign n987 = ~pi129 & ~n986;
  assign n988 = ~n985 & n987;
  assign n989 = ~n887 & n947;
  assign n990 = ~pi48 & ~n989;
  assign po63 = n988 & ~n990;
  assign n992 = pi82 & ~n406;
  assign n993 = ~n379 & ~n992;
  assign n994 = ~pi69 & n993;
  assign n995 = n404 & n595;
  assign n996 = pi49 & ~n995;
  assign n997 = ~pi50 & ~n631;
  assign n998 = n406 & n997;
  assign n999 = ~n996 & ~n998;
  assign n1000 = pi82 & ~n999;
  assign n1001 = pi49 & n409;
  assign n1002 = ~n1000 & ~n1001;
  assign n1003 = ~n994 & n1002;
  assign po64 = ~pi129 & ~n1003;
  assign n1005 = n402 & n918;
  assign n1006 = pi82 & ~n1005;
  assign n1007 = n379 & ~n1006;
  assign n1008 = ~n395 & ~n1007;
  assign n1009 = ~pi50 & ~n1008;
  assign n1010 = n394 & n631;
  assign n1011 = n595 & n1010;
  assign n1012 = pi82 & ~n1011;
  assign n1013 = ~n379 & ~n1012;
  assign n1014 = pi66 & n1013;
  assign n1015 = n394 & n960;
  assign n1016 = ~pi129 & ~n1015;
  assign n1017 = ~n1014 & n1016;
  assign po65 = ~n1009 & n1017;
  assign n1019 = pi51 & ~pi109;
  assign n1020 = ~n859 & ~n1019;
  assign n1021 = ~pi106 & n1020;
  assign po66 = ~pi129 & ~n1021;
  assign n1023 = pi52 & ~n859;
  assign n1024 = ~pi106 & ~n863;
  assign n1025 = ~n1023 & n1024;
  assign po67 = ~pi129 & ~n1025;
  assign n1027 = ~pi116 & n763;
  assign n1028 = ~n762 & ~n1027;
  assign n1029 = ~pi129 & ~n1028;
  assign n1030 = ~pi3 & n1029;
  assign n1031 = n687 & n1030;
  assign po68 = ~pi26 & n1031;
  assign n1033 = n923 & ~n925;
  assign po69 = pi129 | n1033;
  assign po129 = pi123 | pi129;
  assign n1036 = pi114 & ~pi122;
  assign po70 = ~po129 & n1036;
  assign n1038 = ~pi26 & pi58;
  assign n1039 = n662 & ~n756;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = pi94 & ~n1040;
  assign n1042 = pi58 & ~pi116;
  assign n1043 = pi37 & ~pi116;
  assign n1044 = ~n1038 & ~n1043;
  assign n1045 = ~n1042 & ~n1044;
  assign n1046 = ~n1041 & ~n1045;
  assign n1047 = ~pi53 & ~n1046;
  assign n1048 = ~pi26 & pi37;
  assign n1049 = ~pi58 & n1048;
  assign n1050 = ~n1047 & ~n1049;
  assign n1051 = ~pi85 & ~n1050;
  assign n1052 = n701 & n1048;
  assign n1053 = ~n1051 & ~n1052;
  assign n1054 = ~pi27 & ~n1053;
  assign n1055 = n780 & n1048;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = ~pi129 & ~n1056;
  assign po71 = ~pi3 & n1057;
  assign n1059 = ~pi26 & ~pi53;
  assign n1060 = pi26 & pi53;
  assign n1061 = ~pi85 & ~n1060;
  assign n1062 = ~n1059 & ~n1061;
  assign n1063 = ~pi58 & ~n1062;
  assign n1064 = ~pi85 & n1059;
  assign n1065 = ~pi116 & n1064;
  assign n1066 = ~n1063 & ~n1065;
  assign n1067 = pi57 & ~n1066;
  assign n1068 = pi60 & n756;
  assign n1069 = n1064 & n1068;
  assign n1070 = ~n1067 & ~n1069;
  assign n1071 = ~pi27 & ~n1070;
  assign n1072 = pi57 & ~pi58;
  assign n1073 = n1064 & n1072;
  assign n1074 = ~n1071 & ~n1073;
  assign n1075 = ~pi129 & ~n1074;
  assign po72 = ~pi3 & n1075;
  assign n1077 = n741 & n1042;
  assign n1078 = ~pi58 & ~n723;
  assign n1079 = n672 & n1078;
  assign n1080 = ~n1077 & ~n1079;
  assign n1081 = ~pi129 & ~n1080;
  assign n1082 = ~pi3 & n1081;
  assign n1083 = ~pi53 & n1082;
  assign po73 = ~pi85 & n1083;
  assign n1085 = pi59 & ~n767;
  assign n1086 = n660 & n701;
  assign n1087 = pi96 & n1086;
  assign n1088 = ~n1085 & ~n1087;
  assign n1089 = ~pi85 & ~n1088;
  assign n1090 = pi59 & ~pi116;
  assign n1091 = pi85 & n701;
  assign n1092 = n1090 & n1091;
  assign n1093 = ~n1089 & ~n1092;
  assign n1094 = ~pi27 & ~n1093;
  assign n1095 = pi27 & n780;
  assign n1096 = n1090 & n1095;
  assign n1097 = ~n1094 & ~n1096;
  assign n1098 = ~pi26 & ~n1097;
  assign n1099 = n781 & n1090;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = ~pi129 & ~n1100;
  assign po74 = ~pi3 & n1101;
  assign n1103 = ~pi117 & ~pi122;
  assign n1104 = pi60 & ~n1103;
  assign n1105 = pi123 & n1103;
  assign po75 = n1104 | n1105;
  assign n1107 = ~pi114 & pi123;
  assign n1108 = ~pi122 & n1107;
  assign po76 = ~pi129 & n1108;
  assign n1110 = pi136 & ~pi137;
  assign n1111 = pi132 & pi133;
  assign n1112 = pi131 & n1111;
  assign n1113 = ~pi138 & n1112;
  assign n1114 = n1110 & n1113;
  assign n1115 = pi62 & ~n1114;
  assign n1116 = ~pi140 & n1110;
  assign n1117 = n1113 & n1116;
  assign n1118 = ~n1115 & ~n1117;
  assign po77 = pi129 | n1118;
  assign n1120 = pi63 & ~n1114;
  assign n1121 = ~pi142 & n1110;
  assign n1122 = n1113 & n1121;
  assign n1123 = ~n1120 & ~n1122;
  assign po78 = pi129 | n1123;
  assign n1125 = pi64 & ~n1114;
  assign n1126 = ~pi139 & n1110;
  assign n1127 = n1113 & n1126;
  assign n1128 = ~n1125 & ~n1127;
  assign po79 = pi129 | n1128;
  assign n1130 = pi65 & ~n1114;
  assign n1131 = ~pi146 & n1110;
  assign n1132 = n1113 & n1131;
  assign n1133 = ~n1130 & ~n1132;
  assign po80 = pi129 | n1133;
  assign n1135 = ~pi136 & ~pi137;
  assign n1136 = n1113 & n1135;
  assign n1137 = pi66 & ~n1136;
  assign n1138 = ~pi143 & n1136;
  assign n1139 = ~n1137 & ~n1138;
  assign po81 = pi129 | n1139;
  assign n1141 = pi67 & ~n1136;
  assign n1142 = ~pi139 & n1136;
  assign n1143 = ~n1141 & ~n1142;
  assign po82 = pi129 | n1143;
  assign n1145 = pi68 & ~n1114;
  assign n1146 = ~pi141 & n1110;
  assign n1147 = n1113 & n1146;
  assign n1148 = ~n1145 & ~n1147;
  assign po83 = pi129 | n1148;
  assign n1150 = pi69 & ~n1114;
  assign n1151 = ~pi143 & n1110;
  assign n1152 = n1113 & n1151;
  assign n1153 = ~n1150 & ~n1152;
  assign po84 = pi129 | n1153;
  assign n1155 = pi70 & ~n1114;
  assign n1156 = ~pi144 & n1110;
  assign n1157 = n1113 & n1156;
  assign n1158 = ~n1155 & ~n1157;
  assign po85 = pi129 | n1158;
  assign n1160 = pi71 & ~n1114;
  assign n1161 = ~pi145 & n1110;
  assign n1162 = n1113 & n1161;
  assign n1163 = ~n1160 & ~n1162;
  assign po86 = pi129 | n1163;
  assign n1165 = pi72 & ~n1136;
  assign n1166 = ~pi140 & n1136;
  assign n1167 = ~n1165 & ~n1166;
  assign po87 = pi129 | n1167;
  assign n1169 = pi73 & ~n1136;
  assign n1170 = ~pi141 & n1136;
  assign n1171 = ~n1169 & ~n1170;
  assign po88 = pi129 | n1171;
  assign n1173 = pi74 & ~n1136;
  assign n1174 = ~pi142 & n1136;
  assign n1175 = ~n1173 & ~n1174;
  assign po89 = pi129 | n1175;
  assign n1177 = pi75 & ~n1136;
  assign n1178 = ~pi144 & n1136;
  assign n1179 = ~n1177 & ~n1178;
  assign po90 = pi129 | n1179;
  assign n1181 = pi76 & ~n1136;
  assign n1182 = ~pi145 & n1136;
  assign n1183 = ~n1181 & ~n1182;
  assign po91 = pi129 | n1183;
  assign n1185 = pi77 & ~n1136;
  assign n1186 = ~pi146 & n1136;
  assign n1187 = ~n1185 & ~n1186;
  assign po92 = pi129 | n1187;
  assign n1189 = ~pi136 & pi137;
  assign n1190 = n1113 & n1189;
  assign n1191 = pi78 & ~n1190;
  assign n1192 = pi142 & n1190;
  assign n1193 = ~n1191 & ~n1192;
  assign po93 = ~pi129 & ~n1193;
  assign n1195 = pi79 & ~n1190;
  assign n1196 = pi143 & n1190;
  assign n1197 = ~n1195 & ~n1196;
  assign po94 = ~pi129 & ~n1197;
  assign n1199 = pi80 & ~n1190;
  assign n1200 = pi144 & n1190;
  assign n1201 = ~n1199 & ~n1200;
  assign po95 = ~pi129 & ~n1201;
  assign n1203 = pi81 & ~n1190;
  assign n1204 = pi145 & n1190;
  assign n1205 = ~n1203 & ~n1204;
  assign po96 = ~pi129 & ~n1205;
  assign n1207 = pi82 & ~n1190;
  assign n1208 = pi146 & n1190;
  assign n1209 = ~n1207 & ~n1208;
  assign po97 = ~pi129 & ~n1209;
  assign n1211 = pi89 & pi138;
  assign n1212 = ~pi62 & ~pi138;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = pi136 & ~n1213;
  assign n1215 = pi119 & pi138;
  assign n1216 = ~pi72 & ~pi138;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = ~pi136 & ~n1217;
  assign n1219 = ~n1214 & ~n1218;
  assign n1220 = ~pi137 & ~n1219;
  assign n1221 = ~pi115 & pi138;
  assign n1222 = pi87 & ~pi138;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = ~pi136 & ~n1223;
  assign n1225 = pi136 & ~pi138;
  assign n1226 = pi31 & n1225;
  assign n1227 = ~n1224 & ~n1226;
  assign n1228 = pi137 & ~n1227;
  assign po98 = n1220 | n1228;
  assign n1230 = pi84 & ~n1190;
  assign n1231 = pi141 & n1190;
  assign n1232 = ~n1230 & ~n1231;
  assign po99 = ~pi129 & ~n1232;
  assign n1234 = ~pi85 & ~n659;
  assign n1235 = ~pi110 & n1234;
  assign n1236 = pi96 & n1235;
  assign n1237 = ~n649 & ~n1236;
  assign n1238 = ~pi129 & ~n1237;
  assign n1239 = ~pi3 & n1238;
  assign n1240 = n702 & n1239;
  assign po100 = ~pi26 & n1240;
  assign n1242 = pi86 & ~n1190;
  assign n1243 = pi139 & n1190;
  assign n1244 = ~n1242 & ~n1243;
  assign po101 = ~pi129 & ~n1244;
  assign n1246 = pi87 & ~n1190;
  assign n1247 = pi140 & n1190;
  assign n1248 = ~n1246 & ~n1247;
  assign po102 = ~pi129 & ~n1248;
  assign n1250 = pi136 & pi137;
  assign n1251 = n1113 & n1250;
  assign n1252 = pi88 & ~n1251;
  assign n1253 = pi139 & n1251;
  assign n1254 = ~n1252 & ~n1253;
  assign po103 = ~pi129 & ~n1254;
  assign n1256 = pi89 & ~n1251;
  assign n1257 = pi140 & n1251;
  assign n1258 = ~n1256 & ~n1257;
  assign po104 = ~pi129 & ~n1258;
  assign n1260 = pi90 & ~n1251;
  assign n1261 = pi142 & n1251;
  assign n1262 = ~n1260 & ~n1261;
  assign po105 = ~pi129 & ~n1262;
  assign n1264 = pi91 & ~n1251;
  assign n1265 = pi143 & n1251;
  assign n1266 = ~n1264 & ~n1265;
  assign po106 = ~pi129 & ~n1266;
  assign n1268 = pi92 & ~n1251;
  assign n1269 = pi144 & n1251;
  assign n1270 = ~n1268 & ~n1269;
  assign po107 = ~pi129 & ~n1270;
  assign n1272 = pi93 & ~n1251;
  assign n1273 = pi146 & n1251;
  assign n1274 = ~n1272 & ~n1273;
  assign po108 = ~pi129 & ~n1274;
  assign n1276 = pi82 & pi138;
  assign n1277 = n1135 & n1276;
  assign n1278 = n1112 & n1277;
  assign n1279 = pi94 & ~n1278;
  assign n1280 = pi142 & n1278;
  assign n1281 = ~n1279 & ~n1280;
  assign po109 = ~pi129 & ~n1281;
  assign n1283 = ~pi3 & ~n1112;
  assign n1284 = ~pi110 & n1283;
  assign n1285 = n1112 & ~n1277;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = pi95 & ~n1286;
  assign n1288 = pi143 & n1278;
  assign n1289 = ~n1287 & ~n1288;
  assign po110 = ~pi129 & ~n1289;
  assign n1291 = pi96 & ~n1286;
  assign n1292 = pi146 & n1278;
  assign n1293 = ~n1291 & ~n1292;
  assign po111 = ~pi129 & ~n1293;
  assign n1295 = pi97 & ~n1286;
  assign n1296 = pi145 & n1278;
  assign n1297 = ~n1295 & ~n1296;
  assign po112 = ~pi129 & ~n1297;
  assign n1299 = pi98 & ~n1251;
  assign n1300 = pi145 & n1251;
  assign n1301 = ~n1299 & ~n1300;
  assign po113 = ~pi129 & ~n1301;
  assign n1303 = pi99 & ~n1251;
  assign n1304 = pi141 & n1251;
  assign n1305 = ~n1303 & ~n1304;
  assign po114 = ~pi129 & ~n1305;
  assign n1307 = pi100 & ~n1286;
  assign n1308 = pi144 & n1278;
  assign n1309 = ~n1307 & ~n1308;
  assign po115 = ~pi129 & ~n1309;
  assign n1311 = pi124 & pi138;
  assign n1312 = ~pi77 & ~pi138;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = ~pi136 & ~n1313;
  assign n1315 = ~pi65 & ~pi138;
  assign n1316 = pi93 & pi138;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = pi136 & ~n1317;
  assign n1319 = ~n1314 & ~n1318;
  assign n1320 = ~pi137 & ~n1319;
  assign n1321 = pi37 & n1225;
  assign n1322 = pi96 & pi138;
  assign n1323 = pi82 & ~pi138;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = ~pi136 & ~n1324;
  assign n1326 = ~n1321 & ~n1325;
  assign n1327 = pi137 & ~n1326;
  assign po116 = n1320 | n1327;
  assign n1329 = pi91 & n1110;
  assign n1330 = pi95 & n1189;
  assign n1331 = ~n1329 & ~n1330;
  assign n1332 = pi138 & ~n1331;
  assign n1333 = pi79 & ~pi136;
  assign n1334 = pi34 & pi136;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = pi137 & ~n1335;
  assign n1337 = ~pi69 & pi136;
  assign n1338 = ~pi66 & ~pi136;
  assign n1339 = ~n1337 & ~n1338;
  assign n1340 = ~pi137 & ~n1339;
  assign n1341 = ~n1336 & ~n1340;
  assign n1342 = ~pi138 & ~n1341;
  assign po117 = n1332 | n1342;
  assign n1344 = pi90 & n1110;
  assign n1345 = pi94 & n1189;
  assign n1346 = ~n1344 & ~n1345;
  assign n1347 = pi138 & ~n1346;
  assign n1348 = pi78 & ~pi136;
  assign n1349 = pi33 & pi136;
  assign n1350 = ~n1348 & ~n1349;
  assign n1351 = pi137 & ~n1350;
  assign n1352 = ~pi63 & pi136;
  assign n1353 = ~pi74 & ~pi136;
  assign n1354 = ~n1352 & ~n1353;
  assign n1355 = ~pi137 & ~n1354;
  assign n1356 = ~n1351 & ~n1355;
  assign n1357 = ~pi138 & ~n1356;
  assign po118 = n1347 | n1357;
  assign n1359 = pi99 & n1110;
  assign n1360 = ~pi112 & n1189;
  assign n1361 = ~n1359 & ~n1360;
  assign n1362 = pi138 & ~n1361;
  assign n1363 = ~pi68 & pi136;
  assign n1364 = ~pi73 & ~pi136;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = ~pi137 & ~n1365;
  assign n1367 = pi84 & ~pi136;
  assign n1368 = pi32 & pi136;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = pi137 & ~n1369;
  assign n1371 = ~n1366 & ~n1370;
  assign n1372 = ~pi138 & ~n1371;
  assign po119 = n1362 | n1372;
  assign n1374 = pi92 & pi138;
  assign n1375 = ~pi70 & ~pi138;
  assign n1376 = ~n1374 & ~n1375;
  assign n1377 = pi136 & ~n1376;
  assign n1378 = pi125 & pi138;
  assign n1379 = ~pi75 & ~pi138;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = ~pi136 & ~n1380;
  assign n1382 = ~n1377 & ~n1381;
  assign n1383 = ~pi137 & ~n1382;
  assign n1384 = pi80 & ~pi138;
  assign n1385 = pi100 & pi138;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = ~pi136 & ~n1386;
  assign n1388 = pi35 & n1225;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = pi137 & ~n1389;
  assign po120 = n1383 | n1390;
  assign n1392 = n715 & n1235;
  assign n1393 = ~pi27 & n1392;
  assign n1394 = ~n648 & ~n1393;
  assign n1395 = ~pi129 & ~n1394;
  assign po121 = ~pi3 & n1395;
  assign n1397 = pi98 & pi138;
  assign n1398 = ~pi71 & ~pi138;
  assign n1399 = ~n1397 & ~n1398;
  assign n1400 = pi136 & ~n1399;
  assign n1401 = ~pi76 & ~pi138;
  assign n1402 = pi23 & pi138;
  assign n1403 = ~n1401 & ~n1402;
  assign n1404 = ~pi136 & ~n1403;
  assign n1405 = ~n1400 & ~n1404;
  assign n1406 = ~pi137 & ~n1405;
  assign n1407 = pi36 & n1225;
  assign n1408 = pi81 & ~pi138;
  assign n1409 = pi97 & pi138;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~pi136 & ~n1410;
  assign n1412 = ~n1407 & ~n1411;
  assign n1413 = pi137 & ~n1412;
  assign po122 = n1406 | n1413;
  assign n1415 = pi88 & pi138;
  assign n1416 = ~pi64 & ~pi138;
  assign n1417 = ~n1415 & ~n1416;
  assign n1418 = pi136 & ~n1417;
  assign n1419 = pi120 & pi138;
  assign n1420 = ~pi67 & ~pi138;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = ~pi136 & ~n1421;
  assign n1423 = ~n1418 & ~n1422;
  assign n1424 = ~pi137 & ~n1423;
  assign n1425 = pi86 & ~pi138;
  assign n1426 = pi111 & pi138;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = ~pi136 & ~n1427;
  assign n1429 = pi30 & n1225;
  assign n1430 = ~n1428 & ~n1429;
  assign n1431 = pi137 & ~n1430;
  assign po123 = n1424 | n1431;
  assign n1433 = ~n665 & n722;
  assign n1434 = ~n721 & ~n1433;
  assign n1435 = ~pi129 & ~n1434;
  assign n1436 = ~pi3 & n1435;
  assign po124 = pi116 & n1436;
  assign n1438 = ~pi97 & n688;
  assign n1439 = ~n763 & ~n1438;
  assign n1440 = ~pi129 & ~n1439;
  assign n1441 = ~pi3 & n1440;
  assign po125 = pi116 & n1441;
  assign n1443 = pi111 & ~n1277;
  assign n1444 = pi139 & n1277;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = n1112 & ~n1445;
  assign po126 = ~pi129 & n1446;
  assign n1448 = ~pi112 & ~n1277;
  assign n1449 = pi141 & n1277;
  assign n1450 = ~n1448 & ~n1449;
  assign n1451 = n1112 & ~n1450;
  assign po127 = ~pi129 & n1451;
  assign n1453 = ~pi54 & ~pi113;
  assign n1454 = ~pi11 & ~pi22;
  assign n1455 = pi54 & ~n1454;
  assign n1456 = ~n1453 & ~n1455;
  assign n1457 = ~pi129 & ~n1456;
  assign po128 = ~pi3 & n1457;
  assign n1459 = ~pi115 & ~n1277;
  assign n1460 = pi140 & n1277;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = n1112 & ~n1461;
  assign po130 = ~pi129 & n1462;
  assign n1464 = ~pi4 & ~pi12;
  assign n1465 = ~pi7 & ~pi9;
  assign n1466 = n1464 & n1465;
  assign n1467 = ~pi129 & ~n1466;
  assign n1468 = ~pi3 & n1467;
  assign po131 = pi54 & n1468;
  assign po132 = ~pi122 | pi129;
  assign n1471 = ~pi54 & pi118;
  assign n1472 = pi29 & n523;
  assign n1473 = pi54 & ~pi59;
  assign n1474 = n1472 & n1473;
  assign n1475 = ~n1471 & ~n1474;
  assign po133 = ~pi129 & ~n1475;
  assign po134 = ~pi129 & ~n658;
  assign n1478 = ~pi110 & ~pi120;
  assign n1479 = ~pi3 & n1478;
  assign n1480 = ~pi129 & ~n1479;
  assign po135 = ~pi111 & n1480;
  assign n1482 = pi81 & pi120;
  assign po136 = ~pi129 & n1482;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi57 & ~pi129;
  assign n1487 = ~pi96 & pi125;
  assign n1488 = ~pi3 & ~n1487;
  assign po140 = ~pi129 & ~n1488;
  assign n1490 = ~pi126 & pi132;
  assign po141 = pi133 & n1490;
  assign po12 = 1'b1;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
endmodule
