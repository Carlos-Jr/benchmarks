module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 ,
    po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 ,
    po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 ,
    po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 ,
    po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 ,
    po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 ,
    po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 ,
    po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 ,
    po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 ,
    po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ;
  output po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 ,
    po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 ,
    po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 ,
    po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 ,
    po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 ,
    po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 ,
    po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 ,
    po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 ,
    po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 ,
    po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ;
  wire n194, n196, n197, n198, n200, n201, n202,
    n203, n204, n205, n206, n207, n209, n210,
    n211, n212, n213, n214, n215, n216, n217,
    n218, n219, n220, n221, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n291,
    n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n362, n363,
    n364, n365, n366, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391,
    n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n455, n456,
    n457, n458, n459, n460, n461, n462, n463,
    n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n505, n506,
    n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555,
    n556, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811,
    n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825,
    n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847,
    n848, n849, n850, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n861,
    n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889,
    n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n904,
    n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925,
    n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068,
    n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159,
    n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372,
    n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402,
    n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432,
    n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444,
    n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511,
    n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541,
    n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572,
    n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602,
    n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614,
    n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632,
    n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681,
    n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711,
    n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741,
    n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1771,
    n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056,
    n2057, n2058, n2059, n2060, n2061, n2062,
    n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086,
    n2087, n2088, n2089, n2090, n2091, n2092,
    n2093, n2094, n2095, n2096, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122,
    n2123, n2124, n2125, n2126, n2127, n2128,
    n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2150, n2151, n2152,
    n2153, n2154, n2155, n2156, n2157, n2158,
    n2159, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183,
    n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213,
    n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231,
    n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273,
    n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291,
    n2292, n2293, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376,
    n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388,
    n2389, n2390, n2391, n2392, n2393, n2394,
    n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406,
    n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424,
    n2425, n2426, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461,
    n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521,
    n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551,
    n2552, n2553, n2554, n2555, n2556, n2557,
    n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569,
    n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872,
    n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884,
    n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896,
    n2897, n2898, n2899, n2900, n2901, n2902,
    n2903, n2904, n2905, n2906, n2907, n2908,
    n2909, n2910, n2911, n2912, n2913, n2914,
    n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926,
    n2927, n2928, n2929, n2930, n2931, n2932,
    n2933, n2934, n2935, n2936, n2937, n2938,
    n2939, n2940, n2941, n2942, n2943, n2944,
    n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956,
    n2957, n2958, n2959, n2960, n2961, n2962,
    n2963, n2964, n2965, n2966, n2967, n2968,
    n2969, n2970, n2971, n2972, n2973, n2974,
    n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986,
    n2987, n2988, n2989, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2997, n2998,
    n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016,
    n3017, n3018, n3019, n3021, n3022, n3023,
    n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035,
    n3036, n3037, n3038, n3039, n3040, n3041,
    n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053,
    n3054, n3055, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3065,
    n3066, n3067, n3068, n3069, n3070, n3071,
    n3072, n3073, n3074, n3075, n3076, n3077,
    n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3095,
    n3096, n3097, n3098, n3099, n3100, n3101,
    n3102, n3103, n3104, n3105, n3106, n3107,
    n3108, n3109, n3110, n3111, n3112, n3113,
    n3114, n3115, n3116, n3117, n3118, n3119,
    n3120, n3121, n3122, n3123, n3124, n3125,
    n3126, n3127, n3128, n3129, n3130, n3131,
    n3132, n3133, n3134, n3135, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143,
    n3144, n3145, n3146, n3147, n3148, n3149,
    n3150, n3151, n3152, n3153, n3154, n3155,
    n3156, n3157, n3158, n3159, n3160, n3161,
    n3162, n3163, n3164, n3165, n3166, n3167,
    n3168, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179,
    n3180, n3181, n3182, n3183, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282,
    n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300,
    n3301, n3302, n3303, n3304, n3305, n3306,
    n3307, n3308, n3309, n3310, n3311, n3312,
    n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324,
    n3325, n3326, n3327, n3328, n3329, n3330,
    n3331, n3332, n3333, n3334, n3335, n3336,
    n3337, n3338, n3339, n3340, n3341, n3342,
    n3343, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3684, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3862,
    n3863, n3864, n3865, n3866, n3867, n3868,
    n3869, n3870, n3871, n3872, n3873, n3874,
    n3875, n3876, n3877, n3878, n3879, n3880,
    n3881, n3882, n3883, n3884, n3885, n3886,
    n3887, n3888, n3889, n3890, n3891, n3892,
    n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3902, n3903, n3904,
    n3905, n3906, n3907, n3908, n3909, n3910,
    n3911, n3912, n3913, n3914, n3915, n3916,
    n3917, n3918, n3919, n3920, n3921, n3922,
    n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934,
    n3935, n3936, n3937, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006,
    n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036,
    n4037, n4038, n4039, n4041, n4042, n4043,
    n4044, n4045, n4046, n4047, n4048, n4049,
    n4050, n4051, n4052, n4053, n4054, n4055,
    n4056, n4057, n4058, n4059, n4060, n4061,
    n4062, n4063, n4064, n4065, n4066, n4067,
    n4068, n4069, n4070, n4071, n4072, n4073,
    n4074, n4075, n4076, n4077, n4078, n4079,
    n4080, n4081, n4082, n4083, n4084, n4085,
    n4086, n4087, n4088, n4089, n4090, n4091,
    n4092, n4093, n4094, n4095, n4096, n4097,
    n4098, n4099, n4100, n4101, n4102, n4103,
    n4104, n4105, n4106, n4107, n4108, n4109,
    n4110, n4111, n4112, n4113, n4114, n4115,
    n4116, n4117, n4118, n4119, n4120, n4121,
    n4122, n4123, n4124, n4125, n4126, n4127,
    n4128, n4129, n4130, n4131, n4132, n4133,
    n4134, n4135, n4136, n4137, n4138, n4139,
    n4140, n4141, n4142, n4143, n4144, n4145,
    n4146, n4147, n4148, n4149, n4150, n4151,
    n4152, n4153, n4154, n4155, n4156, n4157,
    n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181,
    n4182, n4183, n4184, n4185, n4186, n4187,
    n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217,
    n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4228, n4229, n4230,
    n4231, n4232, n4233, n4234, n4235, n4236,
    n4237, n4238, n4239, n4240, n4241, n4242,
    n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254,
    n4255, n4256, n4257, n4258, n4259, n4260,
    n4261, n4262, n4263, n4264, n4265, n4266,
    n4267, n4268, n4269, n4270, n4271, n4272,
    n4273, n4274, n4275, n4276, n4277, n4278,
    n4279, n4280, n4281, n4282, n4283, n4284,
    n4285, n4286, n4287, n4288, n4289, n4290,
    n4291, n4292, n4293, n4294, n4295, n4296,
    n4297, n4298, n4299, n4300, n4301, n4302,
    n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314,
    n4315, n4316, n4317, n4318, n4319, n4320,
    n4321, n4322, n4323, n4324, n4325, n4326,
    n4327, n4328, n4329, n4330, n4331, n4332,
    n4333, n4334, n4335, n4336, n4337, n4338,
    n4339, n4340, n4341, n4342, n4343, n4344,
    n4345, n4346, n4347, n4348, n4349, n4350,
    n4351, n4352, n4353, n4354, n4355, n4356,
    n4357, n4358, n4359, n4360, n4361, n4362,
    n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392,
    n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4416, n4417,
    n4418, n4419, n4420, n4421, n4422, n4423,
    n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4432, n4433, n4434, n4435,
    n4436, n4437, n4438, n4439, n4440, n4441,
    n4442, n4443, n4444, n4445, n4446, n4447,
    n4448, n4449, n4450, n4451, n4452, n4453,
    n4454, n4455, n4456, n4457, n4458, n4459,
    n4460, n4461, n4462, n4463, n4464, n4465,
    n4466, n4467, n4468, n4469, n4470, n4471,
    n4472, n4473, n4474, n4475, n4476, n4477,
    n4478, n4479, n4480, n4481, n4482, n4483,
    n4484, n4485, n4486, n4487, n4488, n4489,
    n4490, n4491, n4492, n4493, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501,
    n4502, n4503, n4504, n4505, n4506, n4507,
    n4508, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525,
    n4526, n4527, n4528, n4529, n4530, n4531,
    n4532, n4533, n4534, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622,
    n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682,
    n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700,
    n4701, n4702, n4703, n4704, n4705, n4706,
    n4707, n4708, n4709, n4710, n4711, n4712,
    n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724,
    n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742,
    n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802,
    n4803, n4804, n4805, n4806, n4807, n4809,
    n4810, n4811, n4812, n4813, n4814, n4815,
    n4816, n4817, n4818, n4819, n4820, n4821,
    n4822, n4823, n4824, n4825, n4826, n4827,
    n4828, n4829, n4830, n4831, n4832, n4833,
    n4834, n4835, n4836, n4837, n4838, n4839,
    n4840, n4841, n4842, n4843, n4844, n4845,
    n4846, n4847, n4848, n4849, n4850, n4851,
    n4852, n4853, n4854, n4855, n4856, n4857,
    n4858, n4859, n4860, n4861, n4862, n4863,
    n4864, n4865, n4866, n4867, n4868, n4869,
    n4870, n4871, n4872, n4873, n4874, n4875,
    n4876, n4877, n4878, n4879, n4880, n4881,
    n4882, n4883, n4884, n4885, n4886, n4887,
    n4888, n4889, n4890, n4891, n4892, n4893,
    n4894, n4895, n4896, n4897, n4898, n4899,
    n4900, n4901, n4902, n4903, n4904, n4905,
    n4906, n4907, n4908, n4909, n4910, n4911,
    n4912, n4913, n4914, n4915, n4916, n4917,
    n4918, n4919, n4920, n4921, n4922, n4923,
    n4924, n4925, n4926, n4927, n4928, n4929,
    n4930, n4931, n4932, n4933, n4934, n4935,
    n4936, n4937, n4938, n4939, n4940, n4941,
    n4942, n4943, n4944, n4945, n4946, n4947,
    n4948, n4949, n4950, n4951, n4952, n4953,
    n4954, n4955, n4956, n4957, n4958, n4959,
    n4960, n4961, n4962, n4963, n4964, n4965,
    n4966, n4967, n4968, n4969, n4970, n4971,
    n4972, n4973, n4974, n4975, n4976, n4977,
    n4978, n4979, n4980, n4981, n4982, n4983,
    n4984, n4985, n4986, n4987, n4988, n4989,
    n4990, n4991, n4992, n4993, n4994, n4995,
    n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5003, n5004, n5005, n5006, n5007,
    n5008, n5009, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019,
    n5020, n5021, n5022, n5024, n5025, n5026,
    n5027, n5028, n5029, n5030, n5031, n5032,
    n5033, n5034, n5035, n5036, n5037, n5038,
    n5039, n5040, n5041, n5042, n5043, n5044,
    n5045, n5046, n5047, n5048, n5049, n5050,
    n5051, n5052, n5053, n5054, n5055, n5056,
    n5057, n5058, n5059, n5060, n5061, n5062,
    n5063, n5064, n5065, n5066, n5067, n5068,
    n5069, n5070, n5071, n5072, n5073, n5074,
    n5075, n5076, n5077, n5078, n5079, n5080,
    n5081, n5082, n5083, n5084, n5085, n5086,
    n5087, n5088, n5089, n5090, n5091, n5092,
    n5093, n5094, n5095, n5096, n5097, n5098,
    n5099, n5100, n5101, n5102, n5103, n5104,
    n5105, n5106, n5107, n5108, n5109, n5110,
    n5111, n5112, n5113, n5114, n5115, n5116,
    n5117, n5118, n5119, n5120, n5121, n5122,
    n5123, n5124, n5125, n5126, n5127, n5128,
    n5129, n5130, n5131, n5132, n5133, n5134,
    n5135, n5136, n5137, n5138, n5139, n5140,
    n5141, n5142, n5143, n5144, n5145, n5146,
    n5147, n5148, n5149, n5150, n5151, n5152,
    n5153, n5154, n5155, n5156, n5157, n5158,
    n5159, n5160, n5161, n5162, n5163, n5164,
    n5165, n5166, n5167, n5168, n5169, n5170,
    n5171, n5172, n5173, n5174, n5175, n5176,
    n5177, n5178, n5179, n5180, n5181, n5182,
    n5183, n5184, n5185, n5186, n5187, n5188,
    n5189, n5190, n5191, n5192, n5193, n5194,
    n5195, n5196, n5197, n5198, n5199, n5200,
    n5201, n5202, n5203, n5204, n5205, n5206,
    n5207, n5208, n5209, n5210, n5211, n5212,
    n5213, n5214, n5215, n5216, n5217, n5218,
    n5219, n5220, n5221, n5222, n5223, n5224,
    n5225, n5226, n5227, n5229, n5230, n5231,
    n5232, n5233, n5234, n5235, n5236, n5237,
    n5238, n5239, n5240, n5241, n5242, n5243,
    n5244, n5245, n5246, n5247, n5248, n5249,
    n5250, n5251, n5252, n5253, n5254, n5255,
    n5256, n5257, n5258, n5259, n5260, n5261,
    n5262, n5263, n5264, n5265, n5266, n5267,
    n5268, n5269, n5270, n5271, n5272, n5273,
    n5274, n5275, n5276, n5277, n5278, n5279,
    n5280, n5281, n5282, n5283, n5284, n5285,
    n5286, n5287, n5288, n5289, n5290, n5291,
    n5292, n5293, n5294, n5295, n5296, n5297,
    n5298, n5299, n5300, n5301, n5302, n5303,
    n5304, n5305, n5306, n5307, n5308, n5309,
    n5310, n5311, n5312, n5313, n5314, n5315,
    n5316, n5317, n5318, n5319, n5320, n5321,
    n5322, n5323, n5324, n5325, n5326, n5327,
    n5328, n5329, n5330, n5331, n5332, n5333,
    n5334, n5335, n5336, n5337, n5338, n5339,
    n5340, n5341, n5342, n5343, n5344, n5345,
    n5346, n5347, n5348, n5349, n5350, n5351,
    n5352, n5353, n5354, n5355, n5356, n5357,
    n5358, n5359, n5360, n5361, n5362, n5363,
    n5364, n5365, n5366, n5367, n5368, n5369,
    n5370, n5371, n5372, n5373, n5374, n5375,
    n5376, n5377, n5378, n5379, n5380, n5381,
    n5382, n5383, n5384, n5385, n5386, n5387,
    n5388, n5389, n5390, n5391, n5392, n5393,
    n5394, n5395, n5396, n5397, n5398, n5399,
    n5400, n5401, n5402, n5403, n5404, n5405,
    n5406, n5407, n5408, n5409, n5410, n5411,
    n5412, n5413, n5414, n5415, n5416, n5417,
    n5418, n5419, n5420, n5421, n5422, n5423,
    n5424, n5425, n5426, n5427, n5428, n5429,
    n5430, n5431, n5432, n5433, n5434, n5435,
    n5436, n5437, n5438, n5439, n5440, n5441,
    n5443, n5444, n5445, n5446, n5447, n5448,
    n5449, n5450, n5451, n5452, n5453, n5454,
    n5455, n5456, n5457, n5458, n5459, n5460,
    n5461, n5462, n5463, n5464, n5465, n5466,
    n5467, n5468, n5469, n5470, n5471, n5472,
    n5473, n5474, n5475, n5476, n5477, n5478,
    n5479, n5480, n5481, n5482, n5483, n5484,
    n5485, n5486, n5487, n5488, n5489, n5490,
    n5491, n5492, n5493, n5494, n5495, n5496,
    n5497, n5498, n5499, n5500, n5501, n5502,
    n5503, n5504, n5505, n5506, n5507, n5508,
    n5509, n5510, n5511, n5512, n5513, n5514,
    n5515, n5516, n5517, n5518, n5519, n5520,
    n5521, n5522, n5523, n5524, n5525, n5526,
    n5527, n5528, n5529, n5530, n5531, n5532,
    n5533, n5534, n5535, n5536, n5537, n5538,
    n5539, n5540, n5541, n5542, n5543, n5544,
    n5545, n5546, n5547, n5548, n5549, n5550,
    n5551, n5552, n5553, n5554, n5555, n5556,
    n5557, n5558, n5559, n5560, n5561, n5562,
    n5563, n5564, n5565, n5566, n5567, n5568,
    n5569, n5570, n5571, n5572, n5573, n5574,
    n5575, n5576, n5577, n5578, n5579, n5580,
    n5581, n5582, n5583, n5584, n5585, n5586,
    n5587, n5588, n5589, n5590, n5591, n5592,
    n5593, n5594, n5595, n5596, n5597, n5598,
    n5599, n5600, n5601, n5602, n5603, n5604,
    n5605, n5606, n5607, n5608, n5609, n5610,
    n5611, n5612, n5613, n5614, n5615, n5616,
    n5617, n5618, n5619, n5620, n5621, n5622,
    n5623, n5624, n5625, n5626, n5627, n5628,
    n5629, n5630, n5631, n5632, n5633, n5634,
    n5635, n5636, n5637, n5638, n5639, n5640,
    n5641, n5642, n5643, n5644, n5645, n5646,
    n5647, n5648, n5649, n5650, n5651, n5652,
    n5653, n5654, n5655, n5656, n5657, n5658,
    n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5667, n5668, n5669, n5670, n5671,
    n5672, n5673, n5674, n5675, n5676, n5677,
    n5678, n5679, n5680, n5681, n5682, n5683,
    n5684, n5685, n5686, n5687, n5688, n5689,
    n5690, n5691, n5692, n5693, n5694, n5695,
    n5696, n5697, n5698, n5699, n5700, n5701,
    n5702, n5703, n5704, n5705, n5706, n5707,
    n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5715, n5716, n5717, n5718, n5719,
    n5720, n5721, n5722, n5723, n5724, n5725,
    n5726, n5727, n5728, n5729, n5730, n5731,
    n5732, n5733, n5734, n5735, n5736, n5737,
    n5738, n5739, n5740, n5741, n5742, n5743,
    n5744, n5745, n5746, n5747, n5748, n5749,
    n5750, n5751, n5752, n5753, n5754, n5755,
    n5756, n5757, n5758, n5759, n5760, n5761,
    n5762, n5763, n5764, n5765, n5766, n5767,
    n5768, n5769, n5770, n5771, n5772, n5773,
    n5774, n5775, n5776, n5777, n5778, n5779,
    n5780, n5781, n5782, n5783, n5784, n5785,
    n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5794, n5795, n5796, n5797,
    n5798, n5799, n5800, n5801, n5802, n5803,
    n5804, n5805, n5806, n5807, n5808, n5809,
    n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5817, n5818, n5819, n5820, n5821,
    n5822, n5823, n5824, n5825, n5826, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833,
    n5834, n5835, n5836, n5837, n5838, n5839,
    n5840, n5841, n5842, n5843, n5844, n5845,
    n5846, n5847, n5848, n5849, n5850, n5851,
    n5852, n5853, n5854, n5855, n5856, n5857,
    n5858, n5859, n5860, n5861, n5862, n5863,
    n5864, n5865, n5866, n5867, n5868, n5869,
    n5870, n5871, n5872, n5873, n5874, n5875,
    n5876, n5877, n5878, n5879, n5880, n5881,
    n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894,
    n5895, n5896, n5897, n5898, n5899, n5900,
    n5901, n5902, n5903, n5904, n5905, n5906,
    n5907, n5908, n5909, n5910, n5911, n5912,
    n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924,
    n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954,
    n5955, n5956, n5957, n5958, n5959, n5960,
    n5961, n5962, n5963, n5964, n5965, n5966,
    n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984,
    n5985, n5986, n5987, n5988, n5989, n5990,
    n5991, n5992, n5993, n5994, n5995, n5996,
    n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008,
    n6009, n6010, n6011, n6012, n6013, n6014,
    n6015, n6016, n6017, n6018, n6019, n6020,
    n6021, n6022, n6023, n6024, n6025, n6026,
    n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038,
    n6039, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050,
    n6051, n6052, n6053, n6054, n6055, n6056,
    n6057, n6058, n6059, n6060, n6061, n6062,
    n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074,
    n6075, n6076, n6077, n6078, n6079, n6080,
    n6081, n6082, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6090, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6107, n6108, n6109, n6110, n6111,
    n6112, n6113, n6114, n6115, n6116, n6117,
    n6118, n6119, n6120, n6121, n6122, n6123,
    n6124, n6125, n6126, n6127, n6128, n6129,
    n6130, n6131, n6132, n6133, n6134, n6135,
    n6136, n6137, n6138, n6139, n6140, n6141,
    n6142, n6143, n6144, n6145, n6146, n6147,
    n6148, n6149, n6150, n6151, n6152, n6153,
    n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6165,
    n6166, n6167, n6168, n6169, n6170, n6171,
    n6172, n6173, n6174, n6175, n6176, n6177,
    n6178, n6179, n6180, n6181, n6182, n6183,
    n6184, n6185, n6186, n6187, n6188, n6189,
    n6190, n6191, n6192, n6193, n6194, n6195,
    n6196, n6197, n6198, n6199, n6200, n6201,
    n6202, n6203, n6204, n6205, n6206, n6207,
    n6208, n6209, n6210, n6211, n6212, n6213,
    n6214, n6215, n6216, n6217, n6218, n6219,
    n6220, n6221, n6222, n6223, n6224, n6225,
    n6226, n6227, n6228, n6229, n6230, n6231,
    n6232, n6233, n6234, n6235, n6236, n6237,
    n6238, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255,
    n6256, n6257, n6258, n6259, n6260, n6261,
    n6262, n6263, n6264, n6265, n6266, n6267,
    n6268, n6269, n6270, n6271, n6272, n6273,
    n6274, n6275, n6276, n6277, n6278, n6279,
    n6280, n6281, n6282, n6283, n6284, n6285,
    n6286, n6287, n6288, n6289, n6290, n6291,
    n6292, n6293, n6294, n6295, n6296, n6297,
    n6298, n6299, n6300, n6301, n6302, n6303,
    n6304, n6305, n6306, n6307, n6308, n6309,
    n6310, n6311, n6312, n6313, n6314, n6315,
    n6316, n6317, n6318, n6319, n6320, n6321,
    n6322, n6323, n6324, n6325, n6326, n6327,
    n6328, n6329, n6330, n6331, n6332, n6333,
    n6334, n6335, n6336, n6337, n6339, n6340,
    n6341, n6342, n6343, n6344, n6345, n6346,
    n6347, n6348, n6349, n6350, n6351, n6352,
    n6353, n6354, n6355, n6356, n6357, n6358,
    n6359, n6360, n6361, n6362, n6363, n6364,
    n6365, n6366, n6367, n6368, n6369, n6370,
    n6371, n6372, n6373, n6374, n6375, n6376,
    n6377, n6378, n6379, n6380, n6381, n6382,
    n6383, n6384, n6385, n6386, n6387, n6388,
    n6389, n6390, n6391, n6392, n6393, n6394,
    n6395, n6396, n6397, n6398, n6399, n6400,
    n6401, n6402, n6403, n6404, n6405, n6406,
    n6407, n6408, n6409, n6410, n6411, n6412,
    n6413, n6414, n6415, n6416, n6417, n6418,
    n6419, n6420, n6421, n6422, n6423, n6424,
    n6425, n6426, n6427, n6428, n6429, n6430,
    n6431, n6432, n6433, n6434, n6435, n6436,
    n6437, n6438, n6439, n6440, n6441, n6442,
    n6443, n6444, n6445, n6446, n6447, n6448,
    n6449, n6450, n6451, n6452, n6453, n6454,
    n6455, n6456, n6457, n6458, n6459, n6460,
    n6461, n6462, n6463, n6464, n6465, n6466,
    n6467, n6468, n6469, n6470, n6471, n6472,
    n6473, n6474, n6475, n6476, n6477, n6478,
    n6479, n6480, n6481, n6482, n6483, n6484,
    n6485, n6486, n6487, n6488, n6489, n6490,
    n6491, n6492, n6493, n6494, n6495, n6496,
    n6497, n6498, n6499, n6500, n6501, n6502,
    n6503, n6504, n6505, n6506, n6507, n6508,
    n6509, n6510, n6511, n6512, n6513, n6514,
    n6515, n6516, n6517, n6518, n6519, n6520,
    n6521, n6522, n6523, n6524, n6525, n6526,
    n6527, n6528, n6529, n6530, n6531, n6532,
    n6533, n6534, n6535, n6536, n6537, n6538,
    n6539, n6540, n6541, n6542, n6543, n6544,
    n6545, n6546, n6547, n6548, n6549, n6550,
    n6551, n6552, n6553, n6554, n6555, n6556,
    n6557, n6558, n6559, n6560, n6561, n6562,
    n6563, n6564, n6565, n6566, n6567, n6568,
    n6569, n6570, n6571, n6572, n6573, n6575,
    n6576, n6577, n6578, n6579, n6580, n6581,
    n6582, n6583, n6584, n6585, n6586, n6587,
    n6588, n6589, n6590, n6591, n6592, n6593,
    n6594, n6595, n6596, n6597, n6598, n6599,
    n6600, n6601, n6602, n6603, n6604, n6605,
    n6606, n6607, n6608, n6609, n6610, n6611,
    n6612, n6613, n6614, n6615, n6616, n6617,
    n6618, n6619, n6620, n6621, n6622, n6623,
    n6624, n6625, n6626, n6627, n6628, n6629,
    n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641,
    n6642, n6643, n6644, n6645, n6646, n6647,
    n6648, n6649, n6650, n6651, n6652, n6653,
    n6654, n6655, n6656, n6657, n6658, n6659,
    n6660, n6661, n6662, n6663, n6664, n6665,
    n6666, n6667, n6668, n6669, n6670, n6671,
    n6672, n6673, n6674, n6675, n6676, n6677,
    n6678, n6679, n6680, n6681, n6682, n6683,
    n6684, n6685, n6686, n6687, n6688, n6689,
    n6690, n6691, n6692, n6693, n6694, n6695,
    n6696, n6697, n6698, n6699, n6700, n6701,
    n6702, n6703, n6704, n6705, n6706, n6707,
    n6708, n6709, n6710, n6711, n6712, n6713,
    n6714, n6715, n6716, n6717, n6718, n6719,
    n6720, n6721, n6722, n6723, n6724, n6725,
    n6726, n6727, n6728, n6729, n6730, n6731,
    n6732, n6733, n6734, n6735, n6736, n6737,
    n6738, n6739, n6740, n6741, n6742, n6743,
    n6744, n6745, n6746, n6747, n6748, n6749,
    n6750, n6751, n6752, n6753, n6754, n6755,
    n6756, n6757, n6758, n6759, n6760, n6761,
    n6762, n6763, n6764, n6765, n6766, n6767,
    n6768, n6769, n6770, n6771, n6772, n6773,
    n6774, n6775, n6776, n6777, n6778, n6779,
    n6780, n6781, n6782, n6783, n6784, n6785,
    n6786, n6787, n6788, n6789, n6790, n6791,
    n6792, n6793, n6794, n6795, n6796, n6797,
    n6798, n6799, n6800, n6801, n6802, n6803,
    n6804, n6805, n6806, n6807, n6808, n6809,
    n6810, n6811, n6812, n6813, n6814, n6815,
    n6816, n6817, n6818, n6819, n6820, n6821,
    n6823, n6824, n6825, n6826, n6827, n6828,
    n6829, n6830, n6831, n6832, n6833, n6834,
    n6835, n6836, n6837, n6838, n6839, n6840,
    n6841, n6842, n6843, n6844, n6845, n6846,
    n6847, n6848, n6849, n6850, n6851, n6852,
    n6853, n6854, n6855, n6856, n6857, n6858,
    n6859, n6860, n6861, n6862, n6863, n6864,
    n6865, n6866, n6867, n6868, n6869, n6870,
    n6871, n6872, n6873, n6874, n6875, n6876,
    n6877, n6878, n6879, n6880, n6881, n6882,
    n6883, n6884, n6885, n6886, n6887, n6888,
    n6889, n6890, n6891, n6892, n6893, n6894,
    n6895, n6896, n6897, n6898, n6899, n6900,
    n6901, n6902, n6903, n6904, n6905, n6906,
    n6907, n6908, n6909, n6910, n6911, n6912,
    n6913, n6914, n6915, n6916, n6917, n6918,
    n6919, n6920, n6921, n6922, n6923, n6924,
    n6925, n6926, n6927, n6928, n6929, n6930,
    n6931, n6932, n6933, n6934, n6935, n6936,
    n6937, n6938, n6939, n6940, n6941, n6942,
    n6943, n6944, n6945, n6946, n6947, n6948,
    n6949, n6950, n6951, n6952, n6953, n6954,
    n6955, n6956, n6957, n6958, n6959, n6960,
    n6961, n6962, n6963, n6964, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972,
    n6973, n6974, n6975, n6976, n6977, n6978,
    n6979, n6980, n6981, n6982, n6983, n6984,
    n6985, n6986, n6987, n6988, n6989, n6990,
    n6991, n6992, n6993, n6994, n6995, n6996,
    n6997, n6998, n6999, n7000, n7001, n7002,
    n7003, n7004, n7005, n7006, n7007, n7008,
    n7009, n7010, n7011, n7012, n7013, n7014,
    n7015, n7016, n7017, n7018, n7019, n7020,
    n7021, n7022, n7023, n7024, n7025, n7026,
    n7027, n7028, n7029, n7030, n7031, n7032,
    n7033, n7034, n7035, n7036, n7037, n7038,
    n7039, n7040, n7041, n7042, n7043, n7044,
    n7045, n7046, n7047, n7048, n7049, n7050,
    n7051, n7052, n7053, n7054, n7055, n7056,
    n7057, n7058, n7059, n7060, n7061, n7062,
    n7063, n7064, n7066, n7067, n7068, n7069,
    n7070, n7071, n7072, n7073, n7074, n7075,
    n7076, n7077, n7078, n7079, n7080, n7081,
    n7082, n7083, n7084, n7085, n7086, n7087,
    n7088, n7089, n7090, n7091, n7092, n7093,
    n7094, n7095, n7096, n7097, n7098, n7099,
    n7100, n7101, n7102, n7103, n7104, n7105,
    n7106, n7107, n7108, n7109, n7110, n7111,
    n7112, n7113, n7114, n7115, n7116, n7117,
    n7118, n7119, n7120, n7121, n7122, n7123,
    n7124, n7125, n7126, n7127, n7128, n7129,
    n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7137, n7138, n7139, n7140, n7141,
    n7142, n7143, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153,
    n7154, n7155, n7156, n7157, n7158, n7159,
    n7160, n7161, n7162, n7163, n7164, n7165,
    n7166, n7167, n7168, n7169, n7170, n7171,
    n7172, n7173, n7174, n7175, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7194, n7195,
    n7196, n7197, n7198, n7199, n7200, n7201,
    n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7227, n7228, n7229, n7230, n7231,
    n7232, n7233, n7234, n7235, n7236, n7237,
    n7238, n7239, n7240, n7241, n7242, n7243,
    n7244, n7245, n7246, n7247, n7248, n7249,
    n7250, n7251, n7252, n7253, n7254, n7255,
    n7256, n7257, n7258, n7259, n7260, n7261,
    n7262, n7263, n7264, n7265, n7266, n7267,
    n7268, n7269, n7270, n7271, n7272, n7273,
    n7274, n7275, n7276, n7277, n7278, n7279,
    n7280, n7281, n7282, n7283, n7284, n7285,
    n7286, n7287, n7288, n7289, n7290, n7291,
    n7292, n7293, n7294, n7295, n7296, n7297,
    n7298, n7299, n7300, n7301, n7302, n7303,
    n7304, n7305, n7306, n7307, n7308, n7309,
    n7310, n7311, n7312, n7313, n7314, n7315,
    n7316, n7317, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352,
    n7353, n7354, n7355, n7356, n7357, n7358,
    n7359, n7360, n7361, n7362, n7363, n7364,
    n7365, n7366, n7367, n7368, n7369, n7370,
    n7371, n7372, n7373, n7374, n7375, n7376,
    n7377, n7378, n7379, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400,
    n7401, n7402, n7403, n7404, n7405, n7406,
    n7407, n7408, n7409, n7410, n7411, n7412,
    n7413, n7414, n7415, n7416, n7417, n7418,
    n7419, n7420, n7421, n7422, n7423, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430,
    n7431, n7432, n7433, n7434, n7435, n7436,
    n7437, n7438, n7439, n7440, n7441, n7442,
    n7443, n7444, n7445, n7446, n7447, n7448,
    n7449, n7450, n7451, n7452, n7453, n7454,
    n7455, n7456, n7457, n7458, n7459, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466,
    n7467, n7468, n7469, n7470, n7471, n7472,
    n7473, n7474, n7475, n7476, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484,
    n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496,
    n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514,
    n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526,
    n7527, n7528, n7529, n7530, n7531, n7532,
    n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556,
    n7557, n7558, n7559, n7560, n7561, n7562,
    n7563, n7564, n7565, n7566, n7567, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581,
    n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611,
    n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653,
    n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683,
    n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713,
    n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7721, n7722, n7723, n7724, n7725,
    n7726, n7727, n7728, n7729, n7730, n7731,
    n7732, n7733, n7734, n7735, n7736, n7737,
    n7738, n7739, n7740, n7741, n7742, n7743,
    n7744, n7745, n7746, n7747, n7748, n7749,
    n7750, n7751, n7752, n7753, n7754, n7755,
    n7756, n7757, n7758, n7759, n7760, n7761,
    n7762, n7763, n7764, n7765, n7766, n7767,
    n7768, n7769, n7770, n7771, n7772, n7773,
    n7774, n7775, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785,
    n7786, n7787, n7788, n7789, n7790, n7791,
    n7792, n7793, n7794, n7795, n7796, n7797,
    n7798, n7799, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821,
    n7822, n7823, n7824, n7825, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834,
    n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852,
    n7853, n7854, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912,
    n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966,
    n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056,
    n8057, n8058, n8059, n8060, n8061, n8062,
    n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8085, n8086, n8087,
    n8088, n8089, n8090, n8091, n8092, n8093,
    n8094, n8095, n8096, n8097, n8098, n8099,
    n8100, n8101, n8102, n8103, n8104, n8105,
    n8106, n8107, n8108, n8109, n8110, n8111,
    n8112, n8113, n8114, n8115, n8116, n8117,
    n8118, n8119, n8120, n8121, n8122, n8123,
    n8124, n8125, n8126, n8127, n8128, n8129,
    n8130, n8131, n8132, n8133, n8134, n8135,
    n8136, n8137, n8138, n8139, n8140, n8141,
    n8142, n8143, n8144, n8145, n8146, n8147,
    n8148, n8149, n8150, n8151, n8152, n8153,
    n8154, n8155, n8156, n8157, n8158, n8159,
    n8160, n8161, n8162, n8163, n8164, n8165,
    n8166, n8167, n8168, n8169, n8170, n8171,
    n8172, n8173, n8174, n8175, n8176, n8177,
    n8178, n8179, n8180, n8181, n8182, n8183,
    n8184, n8185, n8186, n8187, n8188, n8189,
    n8190, n8191, n8192, n8193, n8194, n8195,
    n8196, n8197, n8198, n8199, n8200, n8201,
    n8202, n8203, n8204, n8205, n8206, n8207,
    n8208, n8209, n8210, n8211, n8212, n8213,
    n8214, n8215, n8216, n8217, n8218, n8219,
    n8220, n8221, n8222, n8223, n8224, n8225,
    n8226, n8227, n8228, n8229, n8230, n8231,
    n8232, n8233, n8234, n8235, n8236, n8237,
    n8238, n8239, n8240, n8241, n8242, n8243,
    n8244, n8245, n8246, n8247, n8248, n8249,
    n8250, n8251, n8252, n8253, n8254, n8255,
    n8256, n8257, n8258, n8259, n8260, n8261,
    n8262, n8263, n8264, n8265, n8266, n8267,
    n8268, n8269, n8270, n8271, n8272, n8273,
    n8274, n8275, n8276, n8277, n8278, n8279,
    n8280, n8281, n8282, n8283, n8284, n8285,
    n8286, n8287, n8288, n8289, n8290, n8291,
    n8292, n8293, n8294, n8295, n8296, n8297,
    n8298, n8299, n8300, n8301, n8302, n8303,
    n8304, n8305, n8306, n8307, n8308, n8309,
    n8310, n8311, n8312, n8313, n8314, n8315,
    n8316, n8317, n8318, n8319, n8320, n8321,
    n8322, n8323, n8324, n8325, n8326, n8327,
    n8328, n8329, n8330, n8331, n8332, n8333,
    n8334, n8335, n8336, n8337, n8338, n8339,
    n8340, n8341, n8342, n8343, n8344, n8345,
    n8346, n8347, n8348, n8349, n8350, n8351,
    n8352, n8353, n8354, n8355, n8356, n8357,
    n8359, n8360, n8361, n8362, n8363, n8364,
    n8365, n8366, n8367, n8368, n8369, n8370,
    n8371, n8372, n8373, n8374, n8375, n8376,
    n8377, n8378, n8379, n8380, n8381, n8382,
    n8383, n8384, n8385, n8386, n8387, n8388,
    n8389, n8390, n8391, n8392, n8393, n8394,
    n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8403, n8404, n8405, n8406,
    n8407, n8408, n8409, n8410, n8411, n8412,
    n8413, n8414, n8415, n8416, n8417, n8418,
    n8419, n8420, n8421, n8422, n8423, n8424,
    n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8434, n8435, n8436,
    n8437, n8438, n8439, n8440, n8441, n8442,
    n8443, n8444, n8445, n8446, n8447, n8448,
    n8449, n8450, n8451, n8452, n8453, n8454,
    n8455, n8456, n8457, n8458, n8459, n8460,
    n8461, n8462, n8463, n8464, n8465, n8466,
    n8467, n8468, n8469, n8470, n8471, n8472,
    n8473, n8474, n8475, n8476, n8477, n8478,
    n8479, n8480, n8481, n8482, n8483, n8484,
    n8485, n8486, n8487, n8488, n8489, n8490,
    n8491, n8492, n8493, n8494, n8495, n8496,
    n8497, n8498, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508,
    n8509, n8510, n8511, n8512, n8513, n8514,
    n8515, n8516, n8517, n8518, n8519, n8520,
    n8521, n8522, n8523, n8524, n8525, n8526,
    n8527, n8528, n8529, n8530, n8531, n8532,
    n8533, n8534, n8535, n8536, n8537, n8538,
    n8539, n8540, n8541, n8542, n8543, n8544,
    n8545, n8546, n8547, n8548, n8549, n8550,
    n8551, n8552, n8553, n8554, n8555, n8556,
    n8557, n8558, n8559, n8560, n8561, n8562,
    n8563, n8564, n8565, n8566, n8567, n8568,
    n8569, n8570, n8571, n8572, n8573, n8574,
    n8575, n8576, n8577, n8578, n8579, n8580,
    n8581, n8582, n8583, n8584, n8585, n8586,
    n8587, n8588, n8589, n8590, n8591, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598,
    n8599, n8600, n8601, n8602, n8603, n8604,
    n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8613, n8614, n8615, n8616,
    n8617, n8618, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8632, n8633, n8634, n8635,
    n8636, n8637, n8638, n8639, n8640, n8641,
    n8642, n8643, n8644, n8645, n8646, n8647,
    n8648, n8649, n8650, n8651, n8652, n8653,
    n8654, n8655, n8656, n8657, n8658, n8659,
    n8660, n8661, n8662, n8663, n8664, n8665,
    n8666, n8667, n8668, n8669, n8670, n8671,
    n8672, n8673, n8674, n8675, n8676, n8677,
    n8678, n8679, n8680, n8681, n8682, n8683,
    n8684, n8685, n8686, n8687, n8688, n8689,
    n8690, n8691, n8692, n8693, n8694, n8695,
    n8696, n8697, n8698, n8699, n8700, n8701,
    n8702, n8703, n8704, n8705, n8706, n8707,
    n8708, n8709, n8710, n8711, n8712, n8713,
    n8714, n8715, n8716, n8717, n8718, n8719,
    n8720, n8721, n8722, n8723, n8724, n8725,
    n8726, n8727, n8728, n8729, n8730, n8731,
    n8732, n8733, n8734, n8735, n8736, n8737,
    n8738, n8739, n8740, n8741, n8742, n8743,
    n8744, n8745, n8746, n8747, n8748, n8749,
    n8750, n8751, n8752, n8753, n8754, n8755,
    n8756, n8757, n8758, n8759, n8760, n8761,
    n8762, n8763, n8764, n8765, n8766, n8767,
    n8768, n8769, n8770, n8771, n8772, n8773,
    n8774, n8775, n8776, n8777, n8778, n8779,
    n8780, n8781, n8782, n8783, n8784, n8785,
    n8786, n8787, n8788, n8789, n8790, n8791,
    n8792, n8793, n8794, n8795, n8796, n8797,
    n8798, n8799, n8800, n8801, n8802, n8803,
    n8804, n8805, n8806, n8807, n8808, n8809,
    n8810, n8811, n8812, n8813, n8814, n8815,
    n8816, n8817, n8818, n8819, n8820, n8821,
    n8822, n8823, n8824, n8825, n8826, n8827,
    n8828, n8829, n8830, n8831, n8832, n8833,
    n8834, n8835, n8836, n8837, n8838, n8839,
    n8840, n8841, n8842, n8843, n8844, n8845,
    n8846, n8847, n8848, n8849, n8850, n8851,
    n8852, n8853, n8854, n8855, n8856, n8857,
    n8858, n8859, n8860, n8861, n8862, n8863,
    n8864, n8865, n8866, n8867, n8868, n8869,
    n8870, n8871, n8872, n8873, n8874, n8875,
    n8876, n8877, n8878, n8879, n8880, n8881,
    n8882, n8883, n8884, n8885, n8886, n8887,
    n8888, n8889, n8890, n8891, n8892, n8893,
    n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905,
    n8906, n8907, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8917, n8918,
    n8919, n8920, n8921, n8922, n8923, n8924,
    n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936,
    n8937, n8938, n8939, n8940, n8941, n8942,
    n8943, n8944, n8945, n8946, n8947, n8948,
    n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966,
    n8967, n8968, n8969, n8970, n8971, n8972,
    n8973, n8974, n8975, n8976, n8977, n8978,
    n8979, n8980, n8981, n8982, n8983, n8984,
    n8985, n8986, n8987, n8988, n8989, n8990,
    n8991, n8992, n8993, n8994, n8995, n8996,
    n8997, n8998, n8999, n9000, n9001, n9002,
    n9003, n9004, n9005, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9017, n9018, n9019, n9020,
    n9021, n9022, n9023, n9024, n9025, n9026,
    n9027, n9028, n9029, n9030, n9031, n9032,
    n9033, n9034, n9035, n9036, n9037, n9038,
    n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050,
    n9051, n9052, n9053, n9054, n9055, n9056,
    n9057, n9058, n9059, n9060, n9061, n9062,
    n9063, n9064, n9065, n9066, n9067, n9068,
    n9069, n9070, n9071, n9072, n9073, n9074,
    n9075, n9076, n9077, n9078, n9079, n9080,
    n9081, n9082, n9083, n9084, n9085, n9086,
    n9087, n9088, n9089, n9090, n9091, n9092,
    n9093, n9094, n9095, n9096, n9097, n9098,
    n9099, n9100, n9101, n9102, n9103, n9104,
    n9105, n9106, n9107, n9108, n9109, n9110,
    n9111, n9112, n9113, n9114, n9115, n9116,
    n9117, n9118, n9119, n9120, n9121, n9122,
    n9123, n9124, n9125, n9126, n9127, n9128,
    n9129, n9130, n9131, n9132, n9133, n9134,
    n9135, n9136, n9137, n9138, n9139, n9140,
    n9141, n9142, n9143, n9144, n9145, n9146,
    n9147, n9148, n9149, n9150, n9151, n9152,
    n9153, n9154, n9155, n9156, n9157, n9158,
    n9159, n9160, n9161, n9162, n9163, n9164,
    n9165, n9166, n9167, n9168, n9169, n9170,
    n9171, n9172, n9173, n9174, n9175, n9176,
    n9177, n9178, n9179, n9180, n9181, n9182,
    n9183, n9184, n9186, n9187, n9188, n9189,
    n9190, n9191, n9192, n9193, n9194, n9195,
    n9196, n9197, n9198, n9199, n9200, n9201,
    n9202, n9203, n9204, n9205, n9206, n9207,
    n9208, n9209, n9210, n9211, n9212, n9213,
    n9214, n9215, n9216, n9217, n9218, n9219,
    n9220, n9221, n9222, n9223, n9224, n9225,
    n9226, n9227, n9228, n9229, n9230, n9231,
    n9232, n9233, n9234, n9235, n9236, n9237,
    n9238, n9239, n9240, n9241, n9242, n9243,
    n9244, n9245, n9246, n9247, n9248, n9249,
    n9250, n9251, n9252, n9253, n9254, n9255,
    n9256, n9257, n9258, n9259, n9260, n9261,
    n9262, n9263, n9264, n9265, n9266, n9267,
    n9268, n9269, n9270, n9271, n9272, n9273,
    n9274, n9275, n9276, n9277, n9278, n9279,
    n9280, n9281, n9282, n9283, n9284, n9285,
    n9286, n9287, n9288, n9289, n9290, n9291,
    n9292, n9293, n9294, n9295, n9296, n9297,
    n9298, n9299, n9300, n9301, n9302, n9303,
    n9304, n9305, n9306, n9307, n9308, n9309,
    n9310, n9311, n9312, n9313, n9314, n9315,
    n9316, n9317, n9318, n9319, n9320, n9321,
    n9322, n9323, n9324, n9325, n9326, n9327,
    n9328, n9329, n9330, n9331, n9332, n9333,
    n9334, n9335, n9336, n9337, n9338, n9339,
    n9340, n9341, n9342, n9343, n9344, n9345,
    n9346, n9347, n9348, n9349, n9350, n9351,
    n9352, n9353, n9354, n9355, n9356, n9357,
    n9358, n9359, n9360, n9361, n9362, n9363,
    n9364, n9365, n9366, n9367, n9368, n9369,
    n9370, n9371, n9372, n9373, n9374, n9375,
    n9376, n9377, n9378, n9379, n9380, n9381,
    n9382, n9383, n9384, n9385, n9386, n9387,
    n9388, n9389, n9390, n9391, n9392, n9393,
    n9394, n9395, n9396, n9397, n9398, n9399,
    n9400, n9401, n9402, n9403, n9404, n9405,
    n9406, n9407, n9408, n9409, n9410, n9411,
    n9412, n9413, n9414, n9415, n9416, n9417,
    n9418, n9419, n9420, n9421, n9422, n9423,
    n9424, n9425, n9426, n9427, n9428, n9429,
    n9430, n9431, n9432, n9433, n9434, n9435,
    n9436, n9437, n9438, n9439, n9440, n9441,
    n9442, n9443, n9444, n9445, n9446, n9447,
    n9448, n9449, n9450, n9451, n9452, n9453,
    n9454, n9455, n9456, n9457, n9458, n9460,
    n9461, n9462, n9463, n9464, n9465, n9466,
    n9467, n9468, n9469, n9470, n9471, n9472,
    n9473, n9474, n9475, n9476, n9477, n9478,
    n9479, n9480, n9481, n9482, n9483, n9484,
    n9485, n9486, n9487, n9488, n9489, n9490,
    n9491, n9492, n9493, n9494, n9495, n9496,
    n9497, n9498, n9499, n9500, n9501, n9502,
    n9503, n9504, n9505, n9506, n9507, n9508,
    n9509, n9510, n9511, n9512, n9513, n9514,
    n9515, n9516, n9517, n9518, n9519, n9520,
    n9521, n9522, n9523, n9524, n9525, n9526,
    n9527, n9528, n9529, n9530, n9531, n9532,
    n9533, n9534, n9535, n9536, n9537, n9538,
    n9539, n9540, n9541, n9542, n9543, n9544,
    n9545, n9546, n9547, n9548, n9549, n9550,
    n9551, n9552, n9553, n9554, n9555, n9556,
    n9557, n9558, n9559, n9560, n9561, n9562,
    n9563, n9564, n9565, n9566, n9567, n9568,
    n9569, n9570, n9571, n9572, n9573, n9574,
    n9575, n9576, n9577, n9578, n9579, n9580,
    n9581, n9582, n9583, n9584, n9585, n9586,
    n9587, n9588, n9589, n9590, n9591, n9592,
    n9593, n9594, n9595, n9596, n9597, n9598,
    n9599, n9600, n9601, n9602, n9603, n9604,
    n9605, n9606, n9607, n9608, n9609, n9610,
    n9611, n9612, n9613, n9614, n9615, n9616,
    n9617, n9618, n9619, n9620, n9621, n9622,
    n9623, n9624, n9625, n9626, n9627, n9628,
    n9629, n9630, n9631, n9632, n9633, n9634,
    n9635, n9636, n9637, n9638, n9639, n9640,
    n9641, n9642, n9643, n9644, n9645, n9646,
    n9647, n9648, n9649, n9650, n9651, n9652,
    n9653, n9654, n9655, n9656, n9657, n9658,
    n9659, n9660, n9661, n9662, n9663, n9664,
    n9665, n9666, n9667, n9668, n9669, n9670,
    n9671, n9672, n9673, n9674, n9675, n9676,
    n9677, n9678, n9679, n9680, n9681, n9682,
    n9683, n9684, n9685, n9686, n9687, n9688,
    n9689, n9690, n9691, n9692, n9693, n9694,
    n9695, n9696, n9697, n9698, n9699, n9700,
    n9701, n9702, n9703, n9704, n9705, n9706,
    n9707, n9708, n9709, n9710, n9711, n9712,
    n9713, n9714, n9715, n9716, n9717, n9718,
    n9719, n9720, n9721, n9722, n9723, n9724,
    n9725, n9726, n9727, n9729, n9730, n9731,
    n9732, n9733, n9734, n9735, n9736, n9737,
    n9738, n9739, n9740, n9741, n9742, n9743,
    n9744, n9745, n9746, n9747, n9748, n9749,
    n9750, n9751, n9752, n9753, n9754, n9755,
    n9756, n9757, n9758, n9759, n9760, n9761,
    n9762, n9763, n9764, n9765, n9766, n9767,
    n9768, n9769, n9770, n9771, n9772, n9773,
    n9774, n9775, n9776, n9777, n9778, n9779,
    n9780, n9781, n9782, n9783, n9784, n9785,
    n9786, n9787, n9788, n9789, n9790, n9791,
    n9792, n9793, n9794, n9795, n9796, n9797,
    n9798, n9799, n9800, n9801, n9802, n9803,
    n9804, n9805, n9806, n9807, n9808, n9809,
    n9810, n9811, n9812, n9813, n9814, n9815,
    n9816, n9817, n9818, n9819, n9820, n9821,
    n9822, n9823, n9824, n9825, n9826, n9827,
    n9828, n9829, n9830, n9831, n9832, n9833,
    n9834, n9835, n9836, n9837, n9838, n9839,
    n9840, n9841, n9842, n9843, n9844, n9845,
    n9846, n9847, n9848, n9849, n9850, n9851,
    n9852, n9853, n9854, n9855, n9856, n9857,
    n9858, n9859, n9860, n9861, n9862, n9863,
    n9864, n9865, n9866, n9867, n9868, n9869,
    n9870, n9871, n9872, n9873, n9874, n9875,
    n9876, n9877, n9878, n9879, n9880, n9881,
    n9882, n9883, n9884, n9885, n9886, n9887,
    n9888, n9889, n9890, n9891, n9892, n9893,
    n9894, n9895, n9896, n9897, n9898, n9899,
    n9900, n9901, n9902, n9903, n9904, n9905,
    n9906, n9907, n9908, n9909, n9910, n9911,
    n9912, n9913, n9914, n9915, n9916, n9917,
    n9918, n9919, n9920, n9921, n9922, n9923,
    n9924, n9925, n9926, n9927, n9928, n9929,
    n9930, n9931, n9932, n9933, n9934, n9935,
    n9936, n9937, n9938, n9939, n9940, n9941,
    n9942, n9943, n9944, n9945, n9946, n9947,
    n9948, n9949, n9950, n9951, n9952, n9953,
    n9954, n9955, n9956, n9957, n9958, n9959,
    n9960, n9961, n9962, n9963, n9964, n9965,
    n9966, n9967, n9968, n9969, n9970, n9971,
    n9972, n9973, n9974, n9975, n9976, n9977,
    n9978, n9979, n9980, n9981, n9982, n9983,
    n9984, n9985, n9986, n9987, n9988, n9990,
    n9991, n9992, n9993, n9994, n9995, n9996,
    n9997, n9998, n9999, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026,
    n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044,
    n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062,
    n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074,
    n10075, n10076, n10077, n10078, n10079, n10080,
    n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092,
    n10093, n10094, n10095, n10096, n10097, n10098,
    n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116,
    n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134,
    n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146,
    n10147, n10148, n10149, n10150, n10151, n10152,
    n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170,
    n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188,
    n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200,
    n10201, n10202, n10203, n10204, n10205, n10206,
    n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218,
    n10219, n10220, n10221, n10222, n10223, n10224,
    n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236,
    n10237, n10238, n10239, n10241, n10242, n10243,
    n10244, n10245, n10246, n10247, n10248, n10249,
    n10250, n10251, n10252, n10253, n10254, n10255,
    n10256, n10257, n10258, n10259, n10260, n10261,
    n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10269, n10270, n10271, n10272, n10273,
    n10274, n10275, n10276, n10277, n10278, n10279,
    n10280, n10281, n10282, n10283, n10284, n10285,
    n10286, n10287, n10288, n10289, n10290, n10291,
    n10292, n10293, n10294, n10295, n10296, n10297,
    n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309,
    n10310, n10311, n10312, n10313, n10314, n10315,
    n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327,
    n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345,
    n10346, n10347, n10348, n10349, n10350, n10351,
    n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363,
    n10364, n10365, n10366, n10367, n10368, n10369,
    n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381,
    n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10395, n10396, n10397, n10398, n10399,
    n10400, n10401, n10402, n10403, n10404, n10405,
    n10406, n10407, n10408, n10409, n10410, n10411,
    n10412, n10413, n10414, n10415, n10416, n10417,
    n10418, n10419, n10420, n10421, n10422, n10423,
    n10424, n10425, n10426, n10427, n10428, n10429,
    n10430, n10431, n10432, n10433, n10434, n10435,
    n10436, n10437, n10438, n10439, n10440, n10441,
    n10442, n10443, n10444, n10445, n10446, n10447,
    n10448, n10449, n10450, n10451, n10452, n10453,
    n10454, n10455, n10456, n10457, n10458, n10459,
    n10460, n10461, n10462, n10463, n10464, n10465,
    n10466, n10467, n10468, n10469, n10470, n10471,
    n10472, n10473, n10474, n10475, n10476, n10477,
    n10478, n10479, n10480, n10481, n10482, n10483,
    n10484, n10485, n10486, n10487, n10488, n10489,
    n10490, n10491, n10492, n10493, n10495, n10496,
    n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508,
    n10509, n10510, n10511, n10512, n10513, n10514,
    n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10530, n10531, n10532,
    n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544,
    n10545, n10546, n10547, n10548, n10549, n10550,
    n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562,
    n10563, n10564, n10565, n10566, n10567, n10568,
    n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580,
    n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592,
    n10593, n10594, n10595, n10596, n10597, n10598,
    n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610,
    n10611, n10612, n10613, n10614, n10615, n10616,
    n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634,
    n10635, n10636, n10637, n10638, n10639, n10640,
    n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10651, n10652,
    n10653, n10654, n10655, n10656, n10657, n10658,
    n10659, n10660, n10661, n10662, n10663, n10664,
    n10665, n10666, n10667, n10668, n10669, n10670,
    n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10680, n10681, n10682,
    n10683, n10684, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10698, n10699, n10700,
    n10701, n10702, n10703, n10704, n10705, n10706,
    n10707, n10708, n10709, n10710, n10711, n10712,
    n10713, n10714, n10715, n10716, n10717, n10718,
    n10719, n10720, n10721, n10722, n10723, n10724,
    n10725, n10726, n10727, n10728, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736,
    n10737, n10738, n10739, n10740, n10741, n10742,
    n10743, n10745, n10746, n10747, n10748, n10749,
    n10750, n10751, n10752, n10753, n10754, n10755,
    n10756, n10757, n10758, n10759, n10760, n10761,
    n10762, n10763, n10764, n10765, n10766, n10767,
    n10768, n10769, n10770, n10771, n10772, n10773,
    n10774, n10775, n10776, n10777, n10778, n10779,
    n10780, n10781, n10782, n10783, n10784, n10785,
    n10786, n10787, n10788, n10789, n10790, n10791,
    n10792, n10793, n10794, n10795, n10796, n10797,
    n10798, n10799, n10800, n10801, n10802, n10803,
    n10804, n10805, n10806, n10807, n10808, n10809,
    n10810, n10811, n10812, n10813, n10814, n10815,
    n10816, n10817, n10818, n10819, n10820, n10821,
    n10822, n10823, n10824, n10825, n10826, n10827,
    n10828, n10829, n10830, n10831, n10832, n10833,
    n10834, n10835, n10836, n10837, n10838, n10839,
    n10840, n10841, n10842, n10843, n10844, n10845,
    n10846, n10847, n10848, n10849, n10850, n10851,
    n10852, n10853, n10854, n10855, n10856, n10857,
    n10858, n10859, n10860, n10861, n10862, n10863,
    n10864, n10865, n10866, n10867, n10868, n10869,
    n10870, n10871, n10872, n10873, n10874, n10875,
    n10876, n10877, n10878, n10879, n10880, n10881,
    n10882, n10883, n10884, n10885, n10886, n10887,
    n10888, n10889, n10890, n10891, n10892, n10893,
    n10894, n10895, n10896, n10897, n10898, n10899,
    n10900, n10901, n10902, n10903, n10904, n10905,
    n10906, n10907, n10908, n10909, n10910, n10911,
    n10912, n10913, n10914, n10915, n10916, n10917,
    n10918, n10919, n10920, n10921, n10922, n10923,
    n10924, n10925, n10926, n10927, n10928, n10929,
    n10930, n10931, n10932, n10933, n10934, n10935,
    n10936, n10937, n10938, n10939, n10940, n10941,
    n10942, n10943, n10944, n10945, n10946, n10947,
    n10948, n10949, n10950, n10951, n10952, n10953,
    n10954, n10955, n10956, n10957, n10958, n10959,
    n10960, n10961, n10962, n10963, n10964, n10965,
    n10966, n10967, n10968, n10969, n10970, n10971,
    n10972, n10973, n10974, n10975, n10976, n10977,
    n10978, n10979, n10980, n10981, n10982, n10984,
    n10985, n10986, n10987, n10988, n10989, n10990,
    n10991, n10992, n10993, n10994, n10995, n10996,
    n10997, n10998, n10999, n11000, n11001, n11002,
    n11003, n11004, n11005, n11006, n11007, n11008,
    n11009, n11010, n11011, n11012, n11013, n11014,
    n11015, n11016, n11017, n11018, n11019, n11020,
    n11021, n11022, n11023, n11024, n11025, n11026,
    n11027, n11028, n11029, n11030, n11031, n11032,
    n11033, n11034, n11035, n11036, n11037, n11038,
    n11039, n11040, n11041, n11042, n11043, n11044,
    n11045, n11046, n11047, n11048, n11049, n11050,
    n11051, n11052, n11053, n11054, n11055, n11056,
    n11057, n11058, n11059, n11060, n11061, n11062,
    n11063, n11064, n11065, n11066, n11067, n11068,
    n11069, n11070, n11071, n11072, n11073, n11074,
    n11075, n11076, n11077, n11078, n11079, n11080,
    n11081, n11082, n11083, n11084, n11085, n11086,
    n11087, n11088, n11089, n11090, n11091, n11092,
    n11093, n11094, n11095, n11096, n11097, n11098,
    n11099, n11100, n11101, n11102, n11103, n11104,
    n11105, n11106, n11107, n11108, n11109, n11110,
    n11111, n11112, n11113, n11114, n11115, n11116,
    n11117, n11118, n11119, n11120, n11121, n11122,
    n11123, n11124, n11125, n11126, n11127, n11128,
    n11129, n11130, n11131, n11132, n11133, n11134,
    n11135, n11136, n11137, n11138, n11139, n11140,
    n11141, n11142, n11143, n11144, n11145, n11146,
    n11147, n11148, n11149, n11150, n11151, n11152,
    n11153, n11154, n11155, n11156, n11157, n11158,
    n11159, n11160, n11161, n11162, n11163, n11164,
    n11165, n11166, n11167, n11168, n11169, n11170,
    n11171, n11172, n11173, n11174, n11175, n11176,
    n11177, n11178, n11179, n11180, n11181, n11182,
    n11183, n11184, n11185, n11186, n11187, n11188,
    n11189, n11190, n11191, n11192, n11193, n11194,
    n11195, n11196, n11197, n11198, n11199, n11200,
    n11201, n11202, n11203, n11204, n11205, n11206,
    n11207, n11208, n11209, n11210, n11211, n11212,
    n11213, n11214, n11215, n11216, n11217, n11218,
    n11219, n11221, n11222, n11223, n11224, n11225,
    n11226, n11227, n11228, n11229, n11230, n11231,
    n11232, n11233, n11234, n11235, n11236, n11237,
    n11238, n11239, n11240, n11241, n11242, n11243,
    n11244, n11245, n11246, n11247, n11248, n11249,
    n11250, n11251, n11252, n11253, n11254, n11255,
    n11256, n11257, n11258, n11259, n11260, n11261,
    n11262, n11263, n11264, n11265, n11266, n11267,
    n11268, n11269, n11270, n11271, n11272, n11273,
    n11274, n11275, n11276, n11277, n11278, n11279,
    n11280, n11281, n11282, n11283, n11284, n11285,
    n11286, n11287, n11288, n11289, n11290, n11291,
    n11292, n11293, n11294, n11295, n11296, n11297,
    n11298, n11299, n11300, n11301, n11302, n11303,
    n11304, n11305, n11306, n11307, n11308, n11309,
    n11310, n11311, n11312, n11313, n11314, n11315,
    n11316, n11317, n11318, n11319, n11320, n11321,
    n11322, n11323, n11324, n11325, n11326, n11327,
    n11328, n11329, n11330, n11331, n11332, n11333,
    n11334, n11335, n11336, n11337, n11338, n11339,
    n11340, n11341, n11342, n11343, n11344, n11345,
    n11346, n11347, n11348, n11349, n11350, n11351,
    n11352, n11353, n11354, n11355, n11356, n11357,
    n11358, n11359, n11360, n11361, n11362, n11363,
    n11364, n11365, n11366, n11367, n11368, n11369,
    n11370, n11371, n11372, n11373, n11374, n11375,
    n11376, n11377, n11378, n11379, n11380, n11381,
    n11382, n11383, n11384, n11385, n11386, n11387,
    n11388, n11389, n11390, n11391, n11392, n11393,
    n11394, n11395, n11396, n11397, n11398, n11399,
    n11400, n11401, n11402, n11403, n11404, n11405,
    n11406, n11407, n11408, n11409, n11410, n11411,
    n11412, n11413, n11414, n11415, n11416, n11417,
    n11418, n11419, n11420, n11421, n11422, n11423,
    n11424, n11425, n11426, n11427, n11428, n11429,
    n11430, n11431, n11432, n11433, n11434, n11435,
    n11436, n11437, n11438, n11439, n11440, n11441,
    n11442, n11443, n11444, n11445, n11446, n11447,
    n11448, n11449, n11450, n11451, n11452, n11453,
    n11455, n11456, n11457, n11458, n11459, n11460,
    n11461, n11462, n11463, n11464, n11465, n11466,
    n11467, n11468, n11469, n11470, n11471, n11472,
    n11473, n11474, n11475, n11476, n11477, n11478,
    n11479, n11480, n11481, n11482, n11483, n11484,
    n11485, n11486, n11487, n11488, n11489, n11490,
    n11491, n11492, n11493, n11494, n11495, n11496,
    n11497, n11498, n11499, n11500, n11501, n11502,
    n11503, n11504, n11505, n11506, n11507, n11508,
    n11509, n11510, n11511, n11512, n11513, n11514,
    n11515, n11516, n11517, n11518, n11519, n11520,
    n11521, n11522, n11523, n11524, n11525, n11526,
    n11527, n11528, n11529, n11530, n11531, n11532,
    n11533, n11534, n11535, n11536, n11537, n11538,
    n11539, n11540, n11541, n11542, n11543, n11544,
    n11545, n11546, n11547, n11548, n11549, n11550,
    n11551, n11552, n11553, n11554, n11555, n11556,
    n11557, n11558, n11559, n11560, n11561, n11562,
    n11563, n11564, n11565, n11566, n11567, n11568,
    n11569, n11570, n11571, n11572, n11573, n11574,
    n11575, n11576, n11577, n11578, n11579, n11580,
    n11581, n11582, n11583, n11584, n11585, n11586,
    n11587, n11588, n11589, n11590, n11591, n11592,
    n11593, n11594, n11595, n11596, n11597, n11598,
    n11599, n11600, n11601, n11602, n11603, n11604,
    n11605, n11606, n11607, n11608, n11609, n11610,
    n11611, n11612, n11613, n11614, n11615, n11616,
    n11617, n11618, n11619, n11620, n11621, n11622,
    n11623, n11624, n11625, n11626, n11627, n11628,
    n11629, n11630, n11631, n11632, n11633, n11634,
    n11635, n11636, n11637, n11638, n11639, n11640,
    n11641, n11642, n11643, n11644, n11645, n11646,
    n11647, n11648, n11649, n11650, n11651, n11652,
    n11653, n11654, n11655, n11656, n11657, n11658,
    n11659, n11660, n11661, n11662, n11663, n11664,
    n11665, n11666, n11667, n11668, n11669, n11670,
    n11671, n11672, n11673, n11674, n11675, n11676,
    n11677, n11678, n11679, n11680, n11682, n11683,
    n11684, n11685, n11686, n11687, n11688, n11689,
    n11690, n11691, n11692, n11693, n11694, n11695,
    n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11704, n11705, n11706, n11707,
    n11708, n11709, n11710, n11711, n11712, n11713,
    n11714, n11715, n11716, n11717, n11718, n11719,
    n11720, n11721, n11722, n11723, n11724, n11725,
    n11726, n11727, n11728, n11729, n11730, n11731,
    n11732, n11733, n11734, n11735, n11736, n11737,
    n11738, n11739, n11740, n11741, n11742, n11743,
    n11744, n11745, n11746, n11747, n11748, n11749,
    n11750, n11751, n11752, n11753, n11754, n11755,
    n11756, n11757, n11758, n11759, n11760, n11761,
    n11762, n11763, n11764, n11765, n11766, n11767,
    n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779,
    n11780, n11781, n11782, n11783, n11784, n11785,
    n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797,
    n11798, n11799, n11800, n11801, n11802, n11803,
    n11804, n11805, n11806, n11807, n11808, n11809,
    n11810, n11811, n11812, n11813, n11814, n11815,
    n11816, n11817, n11818, n11819, n11820, n11821,
    n11822, n11823, n11824, n11825, n11826, n11827,
    n11828, n11829, n11830, n11831, n11832, n11833,
    n11834, n11835, n11836, n11837, n11838, n11839,
    n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11849, n11850, n11851,
    n11852, n11853, n11854, n11855, n11856, n11857,
    n11858, n11859, n11860, n11861, n11862, n11863,
    n11864, n11865, n11866, n11867, n11868, n11869,
    n11870, n11871, n11872, n11873, n11874, n11875,
    n11876, n11877, n11878, n11879, n11880, n11881,
    n11882, n11883, n11884, n11885, n11886, n11887,
    n11888, n11889, n11890, n11891, n11892, n11893,
    n11894, n11895, n11896, n11897, n11898, n11899,
    n11900, n11901, n11902, n11903, n11904, n11905,
    n11906, n11907, n11908, n11909, n11910, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044,
    n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12128, n12129,
    n12130, n12131, n12132, n12133, n12134, n12135,
    n12136, n12137, n12138, n12139, n12140, n12141,
    n12142, n12143, n12144, n12145, n12146, n12147,
    n12148, n12149, n12150, n12151, n12152, n12153,
    n12154, n12155, n12156, n12157, n12158, n12159,
    n12160, n12161, n12162, n12163, n12164, n12165,
    n12166, n12167, n12168, n12169, n12170, n12171,
    n12172, n12173, n12174, n12175, n12176, n12177,
    n12178, n12179, n12180, n12181, n12182, n12183,
    n12184, n12185, n12186, n12187, n12188, n12189,
    n12190, n12191, n12192, n12193, n12194, n12195,
    n12196, n12197, n12198, n12199, n12200, n12201,
    n12202, n12203, n12204, n12205, n12206, n12207,
    n12208, n12209, n12210, n12211, n12212, n12213,
    n12214, n12215, n12216, n12217, n12218, n12219,
    n12220, n12221, n12222, n12223, n12224, n12225,
    n12226, n12227, n12228, n12229, n12230, n12231,
    n12232, n12233, n12234, n12235, n12236, n12237,
    n12238, n12239, n12240, n12241, n12242, n12243,
    n12244, n12245, n12246, n12247, n12248, n12249,
    n12250, n12251, n12252, n12253, n12254, n12255,
    n12256, n12257, n12258, n12259, n12260, n12261,
    n12262, n12263, n12264, n12265, n12266, n12267,
    n12268, n12269, n12270, n12271, n12272, n12273,
    n12274, n12275, n12276, n12277, n12278, n12279,
    n12280, n12281, n12282, n12283, n12284, n12285,
    n12286, n12287, n12288, n12289, n12290, n12291,
    n12292, n12293, n12294, n12295, n12296, n12297,
    n12298, n12299, n12300, n12301, n12302, n12303,
    n12304, n12305, n12306, n12307, n12308, n12309,
    n12310, n12311, n12312, n12313, n12314, n12315,
    n12316, n12317, n12318, n12319, n12320, n12321,
    n12322, n12323, n12324, n12325, n12326, n12327,
    n12328, n12329, n12330, n12331, n12332, n12333,
    n12334, n12335, n12336, n12337, n12338, n12339,
    n12340, n12341, n12342, n12344, n12345, n12346,
    n12347, n12348, n12349, n12350, n12351, n12352,
    n12353, n12354, n12355, n12356, n12357, n12358,
    n12359, n12360, n12361, n12362, n12363, n12364,
    n12365, n12366, n12367, n12368, n12369, n12370,
    n12371, n12372, n12373, n12374, n12375, n12376,
    n12377, n12378, n12379, n12380, n12381, n12382,
    n12383, n12384, n12385, n12386, n12387, n12388,
    n12389, n12390, n12391, n12392, n12393, n12394,
    n12395, n12396, n12397, n12398, n12399, n12400,
    n12401, n12402, n12403, n12404, n12405, n12406,
    n12407, n12408, n12409, n12410, n12411, n12412,
    n12413, n12414, n12415, n12416, n12417, n12418,
    n12419, n12420, n12421, n12422, n12423, n12424,
    n12425, n12426, n12427, n12428, n12429, n12430,
    n12431, n12432, n12433, n12434, n12435, n12436,
    n12437, n12438, n12439, n12440, n12441, n12442,
    n12443, n12444, n12445, n12446, n12447, n12448,
    n12449, n12450, n12451, n12452, n12453, n12454,
    n12455, n12456, n12457, n12458, n12459, n12460,
    n12461, n12462, n12463, n12464, n12465, n12466,
    n12467, n12468, n12469, n12470, n12471, n12472,
    n12473, n12474, n12475, n12476, n12477, n12478,
    n12479, n12480, n12481, n12482, n12483, n12484,
    n12485, n12486, n12487, n12488, n12489, n12490,
    n12491, n12492, n12493, n12494, n12495, n12496,
    n12497, n12498, n12499, n12500, n12501, n12502,
    n12503, n12504, n12505, n12506, n12507, n12508,
    n12509, n12510, n12511, n12512, n12513, n12514,
    n12515, n12516, n12517, n12518, n12519, n12520,
    n12521, n12522, n12523, n12524, n12525, n12526,
    n12527, n12528, n12529, n12530, n12531, n12532,
    n12533, n12534, n12535, n12536, n12537, n12538,
    n12539, n12540, n12541, n12542, n12543, n12544,
    n12545, n12546, n12547, n12548, n12549, n12550,
    n12552, n12553, n12554, n12555, n12556, n12557,
    n12558, n12559, n12560, n12561, n12562, n12563,
    n12564, n12565, n12566, n12567, n12568, n12569,
    n12570, n12571, n12572, n12573, n12574, n12575,
    n12576, n12577, n12578, n12579, n12580, n12581,
    n12582, n12583, n12584, n12585, n12586, n12587,
    n12588, n12589, n12590, n12591, n12592, n12593,
    n12594, n12595, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12604, n12605,
    n12606, n12607, n12608, n12609, n12610, n12611,
    n12612, n12613, n12614, n12615, n12616, n12617,
    n12618, n12619, n12620, n12621, n12622, n12623,
    n12624, n12625, n12626, n12627, n12628, n12629,
    n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641,
    n12642, n12643, n12644, n12645, n12646, n12647,
    n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659,
    n12660, n12661, n12662, n12663, n12664, n12665,
    n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677,
    n12678, n12679, n12680, n12681, n12682, n12683,
    n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12691, n12692, n12693, n12694, n12695,
    n12696, n12697, n12698, n12699, n12700, n12701,
    n12702, n12703, n12704, n12705, n12706, n12707,
    n12708, n12709, n12710, n12711, n12712, n12713,
    n12714, n12715, n12716, n12717, n12718, n12719,
    n12720, n12721, n12722, n12723, n12724, n12725,
    n12726, n12727, n12728, n12729, n12730, n12731,
    n12732, n12733, n12734, n12735, n12736, n12737,
    n12738, n12739, n12740, n12741, n12742, n12743,
    n12744, n12745, n12746, n12747, n12748, n12749,
    n12750, n12751, n12752, n12753, n12754, n12755,
    n12756, n12757, n12759, n12760, n12761, n12762,
    n12763, n12764, n12765, n12766, n12767, n12768,
    n12769, n12770, n12771, n12772, n12773, n12774,
    n12775, n12776, n12777, n12778, n12779, n12780,
    n12781, n12782, n12783, n12784, n12785, n12786,
    n12787, n12788, n12789, n12790, n12791, n12792,
    n12793, n12794, n12795, n12796, n12797, n12798,
    n12799, n12800, n12801, n12802, n12803, n12804,
    n12805, n12806, n12807, n12808, n12809, n12810,
    n12811, n12812, n12813, n12814, n12815, n12816,
    n12817, n12818, n12819, n12820, n12821, n12822,
    n12823, n12824, n12825, n12826, n12827, n12828,
    n12829, n12830, n12831, n12832, n12833, n12834,
    n12835, n12836, n12837, n12838, n12839, n12840,
    n12841, n12842, n12843, n12844, n12845, n12846,
    n12847, n12848, n12849, n12850, n12851, n12852,
    n12853, n12854, n12855, n12856, n12857, n12858,
    n12859, n12860, n12861, n12862, n12863, n12864,
    n12865, n12866, n12867, n12868, n12869, n12870,
    n12871, n12872, n12873, n12874, n12875, n12876,
    n12877, n12878, n12879, n12880, n12881, n12882,
    n12883, n12884, n12885, n12886, n12887, n12888,
    n12889, n12890, n12891, n12892, n12893, n12894,
    n12895, n12896, n12897, n12898, n12899, n12900,
    n12901, n12902, n12903, n12904, n12905, n12906,
    n12907, n12908, n12909, n12910, n12911, n12912,
    n12913, n12914, n12915, n12916, n12917, n12918,
    n12919, n12920, n12921, n12922, n12923, n12924,
    n12925, n12926, n12927, n12928, n12929, n12930,
    n12931, n12932, n12933, n12934, n12935, n12936,
    n12937, n12938, n12939, n12940, n12941, n12942,
    n12943, n12944, n12945, n12946, n12947, n12948,
    n12949, n12950, n12951, n12952, n12953, n12954,
    n12956, n12957, n12958, n12959, n12960, n12961,
    n12962, n12963, n12964, n12965, n12966, n12967,
    n12968, n12969, n12970, n12971, n12972, n12973,
    n12974, n12975, n12976, n12977, n12978, n12979,
    n12980, n12981, n12982, n12983, n12984, n12985,
    n12986, n12987, n12988, n12989, n12990, n12991,
    n12992, n12993, n12994, n12995, n12996, n12997,
    n12998, n12999, n13000, n13001, n13002, n13003,
    n13004, n13005, n13006, n13007, n13008, n13009,
    n13010, n13011, n13012, n13013, n13014, n13015,
    n13016, n13017, n13018, n13019, n13020, n13021,
    n13022, n13023, n13024, n13025, n13026, n13027,
    n13028, n13029, n13030, n13031, n13032, n13033,
    n13034, n13035, n13036, n13037, n13038, n13039,
    n13040, n13041, n13042, n13043, n13044, n13045,
    n13046, n13047, n13048, n13049, n13050, n13051,
    n13052, n13053, n13054, n13055, n13056, n13057,
    n13058, n13059, n13060, n13061, n13062, n13063,
    n13064, n13065, n13066, n13067, n13068, n13069,
    n13070, n13071, n13072, n13073, n13074, n13075,
    n13076, n13077, n13078, n13079, n13080, n13081,
    n13082, n13083, n13084, n13085, n13086, n13087,
    n13088, n13089, n13090, n13091, n13092, n13093,
    n13094, n13095, n13096, n13097, n13098, n13099,
    n13100, n13101, n13102, n13103, n13104, n13105,
    n13106, n13107, n13108, n13109, n13110, n13111,
    n13112, n13113, n13114, n13115, n13116, n13117,
    n13118, n13119, n13120, n13121, n13122, n13123,
    n13124, n13125, n13126, n13127, n13128, n13129,
    n13130, n13131, n13132, n13133, n13134, n13135,
    n13136, n13137, n13138, n13139, n13140, n13141,
    n13142, n13143, n13144, n13145, n13146, n13147,
    n13148, n13149, n13150, n13151, n13152, n13153,
    n13154, n13155, n13156, n13157, n13158, n13159,
    n13160, n13162, n13163, n13164, n13165, n13166,
    n13167, n13168, n13169, n13170, n13171, n13172,
    n13173, n13174, n13175, n13176, n13177, n13178,
    n13179, n13180, n13181, n13182, n13183, n13184,
    n13185, n13186, n13187, n13188, n13189, n13190,
    n13191, n13192, n13193, n13194, n13195, n13196,
    n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214,
    n13215, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232,
    n13233, n13234, n13235, n13236, n13237, n13238,
    n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250,
    n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13300, n13301, n13302, n13303, n13304,
    n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n13319, n13320, n13321, n13322,
    n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334,
    n13335, n13336, n13337, n13338, n13339, n13340,
    n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352,
    n13353, n13355, n13356, n13357, n13358, n13359,
    n13360, n13361, n13362, n13363, n13364, n13365,
    n13366, n13367, n13368, n13369, n13370, n13371,
    n13372, n13373, n13374, n13375, n13376, n13377,
    n13378, n13379, n13380, n13381, n13382, n13383,
    n13384, n13385, n13386, n13387, n13388, n13389,
    n13390, n13391, n13392, n13393, n13394, n13395,
    n13396, n13397, n13398, n13399, n13400, n13401,
    n13402, n13403, n13404, n13405, n13406, n13407,
    n13408, n13409, n13410, n13411, n13412, n13413,
    n13414, n13415, n13416, n13417, n13418, n13419,
    n13420, n13421, n13422, n13423, n13424, n13425,
    n13426, n13427, n13428, n13429, n13430, n13431,
    n13432, n13433, n13434, n13435, n13436, n13437,
    n13438, n13439, n13440, n13441, n13442, n13443,
    n13444, n13445, n13446, n13447, n13448, n13449,
    n13450, n13451, n13452, n13453, n13454, n13455,
    n13456, n13457, n13458, n13459, n13460, n13461,
    n13462, n13463, n13464, n13465, n13466, n13467,
    n13468, n13469, n13470, n13471, n13472, n13473,
    n13474, n13475, n13476, n13477, n13478, n13479,
    n13480, n13481, n13482, n13483, n13484, n13485,
    n13486, n13487, n13488, n13489, n13490, n13491,
    n13492, n13493, n13494, n13495, n13496, n13497,
    n13498, n13499, n13500, n13501, n13502, n13503,
    n13504, n13505, n13506, n13507, n13508, n13509,
    n13510, n13511, n13512, n13513, n13514, n13515,
    n13516, n13517, n13518, n13519, n13520, n13521,
    n13522, n13523, n13524, n13525, n13526, n13527,
    n13528, n13529, n13530, n13531, n13532, n13533,
    n13534, n13535, n13536, n13537, n13538, n13539,
    n13540, n13541, n13542, n13543, n13544, n13545,
    n13546, n13548, n13549, n13550, n13551, n13552,
    n13553, n13554, n13555, n13556, n13557, n13558,
    n13559, n13560, n13561, n13562, n13563, n13564,
    n13565, n13566, n13567, n13568, n13569, n13570,
    n13571, n13572, n13573, n13574, n13575, n13576,
    n13577, n13578, n13579, n13580, n13581, n13582,
    n13583, n13584, n13585, n13586, n13587, n13588,
    n13589, n13590, n13591, n13592, n13593, n13594,
    n13595, n13596, n13597, n13598, n13599, n13600,
    n13601, n13602, n13603, n13604, n13605, n13606,
    n13607, n13608, n13609, n13610, n13611, n13612,
    n13613, n13614, n13615, n13616, n13617, n13618,
    n13619, n13620, n13621, n13622, n13623, n13624,
    n13625, n13626, n13627, n13628, n13629, n13630,
    n13631, n13632, n13633, n13634, n13635, n13636,
    n13637, n13638, n13639, n13640, n13641, n13642,
    n13643, n13644, n13645, n13646, n13647, n13648,
    n13649, n13650, n13651, n13652, n13653, n13654,
    n13655, n13656, n13657, n13658, n13659, n13660,
    n13661, n13662, n13663, n13664, n13665, n13666,
    n13667, n13668, n13669, n13670, n13671, n13672,
    n13673, n13674, n13675, n13676, n13677, n13678,
    n13679, n13680, n13681, n13682, n13683, n13684,
    n13685, n13686, n13687, n13688, n13689, n13690,
    n13691, n13692, n13693, n13694, n13695, n13696,
    n13697, n13698, n13699, n13700, n13701, n13702,
    n13703, n13704, n13705, n13706, n13707, n13708,
    n13709, n13710, n13711, n13712, n13713, n13714,
    n13715, n13716, n13717, n13718, n13719, n13720,
    n13721, n13722, n13723, n13724, n13725, n13726,
    n13727, n13728, n13729, n13730, n13731, n13732,
    n13734, n13735, n13736, n13737, n13738, n13739,
    n13740, n13741, n13742, n13743, n13744, n13745,
    n13746, n13747, n13748, n13749, n13750, n13751,
    n13752, n13753, n13754, n13755, n13756, n13757,
    n13758, n13759, n13760, n13761, n13762, n13763,
    n13764, n13765, n13766, n13767, n13768, n13769,
    n13770, n13771, n13772, n13773, n13774, n13775,
    n13776, n13777, n13778, n13779, n13780, n13781,
    n13782, n13783, n13784, n13785, n13786, n13787,
    n13788, n13789, n13790, n13791, n13792, n13793,
    n13794, n13795, n13796, n13797, n13798, n13799,
    n13800, n13801, n13802, n13803, n13804, n13805,
    n13806, n13807, n13808, n13809, n13810, n13811,
    n13812, n13813, n13814, n13815, n13816, n13817,
    n13818, n13819, n13820, n13821, n13822, n13823,
    n13824, n13825, n13826, n13827, n13828, n13829,
    n13830, n13831, n13832, n13833, n13834, n13835,
    n13836, n13837, n13838, n13839, n13840, n13841,
    n13842, n13843, n13844, n13845, n13846, n13847,
    n13848, n13849, n13850, n13851, n13852, n13853,
    n13854, n13855, n13856, n13857, n13858, n13859,
    n13860, n13861, n13862, n13863, n13864, n13865,
    n13866, n13867, n13868, n13869, n13870, n13871,
    n13872, n13873, n13874, n13875, n13876, n13877,
    n13878, n13879, n13880, n13881, n13882, n13883,
    n13884, n13885, n13886, n13887, n13888, n13889,
    n13890, n13891, n13892, n13893, n13894, n13895,
    n13896, n13897, n13898, n13899, n13900, n13901,
    n13902, n13903, n13904, n13905, n13906, n13907,
    n13908, n13909, n13910, n13911, n13912, n13913,
    n13914, n13915, n13916, n13917, n13919, n13920,
    n13921, n13922, n13923, n13924, n13925, n13926,
    n13927, n13928, n13929, n13930, n13931, n13932,
    n13933, n13934, n13935, n13936, n13937, n13938,
    n13939, n13940, n13941, n13942, n13943, n13944,
    n13945, n13946, n13947, n13948, n13949, n13950,
    n13951, n13952, n13953, n13954, n13955, n13956,
    n13957, n13958, n13959, n13960, n13961, n13962,
    n13963, n13964, n13965, n13966, n13967, n13968,
    n13969, n13970, n13971, n13972, n13973, n13974,
    n13975, n13976, n13977, n13978, n13979, n13980,
    n13981, n13982, n13983, n13984, n13985, n13986,
    n13987, n13988, n13989, n13990, n13991, n13992,
    n13993, n13994, n13995, n13996, n13997, n13998,
    n13999, n14000, n14001, n14002, n14003, n14004,
    n14005, n14006, n14007, n14008, n14009, n14010,
    n14011, n14012, n14013, n14014, n14015, n14016,
    n14017, n14018, n14019, n14020, n14021, n14022,
    n14023, n14024, n14025, n14026, n14027, n14028,
    n14029, n14030, n14031, n14032, n14033, n14034,
    n14035, n14036, n14037, n14038, n14039, n14040,
    n14041, n14042, n14043, n14044, n14045, n14046,
    n14047, n14048, n14049, n14050, n14051, n14052,
    n14053, n14054, n14055, n14056, n14057, n14058,
    n14059, n14060, n14061, n14062, n14063, n14064,
    n14065, n14066, n14067, n14068, n14069, n14070,
    n14071, n14072, n14073, n14074, n14075, n14076,
    n14077, n14078, n14079, n14080, n14081, n14082,
    n14083, n14084, n14085, n14086, n14087, n14088,
    n14089, n14090, n14091, n14093, n14094, n14095,
    n14096, n14097, n14098, n14099, n14100, n14101,
    n14102, n14103, n14104, n14105, n14106, n14107,
    n14108, n14109, n14110, n14111, n14112, n14113,
    n14114, n14115, n14116, n14117, n14118, n14119,
    n14120, n14121, n14122, n14123, n14124, n14125,
    n14126, n14127, n14128, n14129, n14130, n14131,
    n14132, n14133, n14134, n14135, n14136, n14137,
    n14138, n14139, n14140, n14141, n14142, n14143,
    n14144, n14145, n14146, n14147, n14148, n14149,
    n14150, n14151, n14152, n14153, n14154, n14155,
    n14156, n14157, n14158, n14159, n14160, n14161,
    n14162, n14163, n14164, n14165, n14166, n14167,
    n14168, n14169, n14170, n14171, n14172, n14173,
    n14174, n14175, n14176, n14177, n14178, n14179,
    n14180, n14181, n14182, n14183, n14184, n14185,
    n14186, n14187, n14188, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197,
    n14198, n14199, n14200, n14201, n14202, n14203,
    n14204, n14205, n14206, n14207, n14208, n14209,
    n14210, n14211, n14212, n14213, n14214, n14215,
    n14216, n14217, n14218, n14219, n14220, n14221,
    n14222, n14223, n14224, n14225, n14226, n14227,
    n14228, n14229, n14230, n14231, n14232, n14233,
    n14234, n14235, n14236, n14237, n14238, n14239,
    n14240, n14241, n14242, n14243, n14244, n14245,
    n14246, n14247, n14248, n14249, n14250, n14251,
    n14252, n14253, n14254, n14255, n14256, n14257,
    n14258, n14259, n14260, n14261, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14329, n14330,
    n14331, n14332, n14333, n14334, n14335, n14336,
    n14337, n14338, n14339, n14340, n14341, n14342,
    n14343, n14344, n14345, n14346, n14347, n14348,
    n14349, n14350, n14351, n14352, n14353, n14354,
    n14355, n14356, n14357, n14358, n14359, n14360,
    n14361, n14362, n14363, n14364, n14365, n14366,
    n14367, n14368, n14369, n14370, n14371, n14372,
    n14373, n14374, n14375, n14376, n14377, n14378,
    n14379, n14380, n14381, n14382, n14383, n14384,
    n14385, n14386, n14387, n14388, n14389, n14390,
    n14391, n14392, n14393, n14394, n14395, n14396,
    n14397, n14398, n14399, n14400, n14401, n14402,
    n14403, n14404, n14405, n14406, n14407, n14408,
    n14409, n14410, n14411, n14412, n14413, n14414,
    n14415, n14416, n14417, n14418, n14419, n14420,
    n14421, n14422, n14423, n14424, n14425, n14426,
    n14427, n14428, n14430, n14431, n14432, n14433,
    n14434, n14435, n14436, n14437, n14438, n14439,
    n14440, n14441, n14442, n14443, n14444, n14445,
    n14446, n14447, n14448, n14449, n14450, n14451,
    n14452, n14453, n14454, n14455, n14456, n14457,
    n14458, n14459, n14460, n14461, n14462, n14463,
    n14464, n14465, n14466, n14467, n14468, n14469,
    n14470, n14471, n14472, n14473, n14474, n14475,
    n14476, n14477, n14478, n14479, n14480, n14481,
    n14482, n14483, n14484, n14485, n14486, n14487,
    n14488, n14489, n14490, n14491, n14492, n14493,
    n14494, n14495, n14496, n14497, n14498, n14499,
    n14500, n14501, n14502, n14503, n14504, n14505,
    n14506, n14507, n14508, n14509, n14510, n14511,
    n14512, n14513, n14514, n14515, n14516, n14517,
    n14518, n14519, n14520, n14521, n14522, n14523,
    n14524, n14525, n14526, n14527, n14528, n14529,
    n14530, n14531, n14532, n14533, n14534, n14535,
    n14536, n14537, n14538, n14539, n14540, n14541,
    n14542, n14543, n14544, n14545, n14546, n14547,
    n14548, n14549, n14550, n14551, n14552, n14553,
    n14554, n14555, n14556, n14557, n14558, n14559,
    n14560, n14561, n14562, n14563, n14564, n14565,
    n14566, n14567, n14568, n14569, n14570, n14571,
    n14572, n14573, n14574, n14575, n14576, n14577,
    n14578, n14579, n14580, n14581, n14582, n14583,
    n14584, n14585, n14586, n14587, n14588, n14589,
    n14590, n14591, n14592, n14593, n14594, n14595,
    n14596, n14598, n14599, n14600, n14601, n14602,
    n14603, n14604, n14605, n14606, n14607, n14608,
    n14609, n14610, n14611, n14612, n14613, n14614,
    n14615, n14616, n14617, n14618, n14619, n14620,
    n14621, n14622, n14623, n14624, n14625, n14626,
    n14627, n14628, n14629, n14630, n14631, n14632,
    n14633, n14634, n14635, n14636, n14637, n14638,
    n14639, n14640, n14641, n14642, n14643, n14644,
    n14645, n14646, n14647, n14648, n14649, n14650,
    n14651, n14652, n14653, n14654, n14655, n14656,
    n14657, n14658, n14659, n14660, n14661, n14662,
    n14663, n14664, n14665, n14666, n14667, n14668,
    n14669, n14670, n14671, n14672, n14673, n14674,
    n14675, n14676, n14677, n14678, n14679, n14680,
    n14681, n14682, n14683, n14684, n14685, n14686,
    n14687, n14688, n14689, n14690, n14691, n14692,
    n14693, n14694, n14695, n14696, n14697, n14698,
    n14699, n14700, n14701, n14702, n14703, n14704,
    n14705, n14706, n14707, n14708, n14709, n14710,
    n14711, n14712, n14713, n14714, n14715, n14716,
    n14717, n14718, n14719, n14720, n14721, n14722,
    n14723, n14724, n14725, n14726, n14727, n14728,
    n14729, n14730, n14731, n14732, n14733, n14734,
    n14735, n14736, n14737, n14738, n14739, n14740,
    n14741, n14742, n14743, n14744, n14745, n14746,
    n14747, n14748, n14749, n14750, n14751, n14752,
    n14753, n14755, n14756, n14757, n14758, n14759,
    n14760, n14761, n14762, n14763, n14764, n14765,
    n14766, n14767, n14768, n14769, n14770, n14771,
    n14772, n14773, n14774, n14775, n14776, n14777,
    n14778, n14779, n14780, n14781, n14782, n14783,
    n14784, n14785, n14786, n14787, n14788, n14789,
    n14790, n14791, n14792, n14793, n14794, n14795,
    n14796, n14797, n14798, n14799, n14800, n14801,
    n14802, n14803, n14804, n14805, n14806, n14807,
    n14808, n14809, n14810, n14811, n14812, n14813,
    n14814, n14815, n14816, n14817, n14818, n14819,
    n14820, n14821, n14822, n14823, n14824, n14825,
    n14826, n14827, n14828, n14829, n14830, n14831,
    n14832, n14833, n14834, n14835, n14836, n14837,
    n14838, n14839, n14840, n14841, n14842, n14843,
    n14844, n14845, n14846, n14847, n14848, n14849,
    n14850, n14851, n14852, n14853, n14854, n14855,
    n14856, n14857, n14858, n14859, n14860, n14861,
    n14862, n14863, n14864, n14865, n14866, n14867,
    n14868, n14869, n14870, n14871, n14872, n14873,
    n14874, n14875, n14876, n14877, n14878, n14879,
    n14880, n14881, n14882, n14883, n14884, n14885,
    n14886, n14887, n14888, n14889, n14890, n14891,
    n14892, n14893, n14894, n14895, n14896, n14897,
    n14898, n14899, n14900, n14901, n14902, n14903,
    n14904, n14905, n14906, n14907, n14908, n14909,
    n14910, n14911, n14913, n14914, n14915, n14916,
    n14917, n14918, n14919, n14920, n14921, n14922,
    n14923, n14924, n14925, n14926, n14927, n14928,
    n14929, n14930, n14931, n14932, n14933, n14934,
    n14935, n14936, n14937, n14938, n14939, n14940,
    n14941, n14942, n14943, n14944, n14945, n14946,
    n14947, n14948, n14949, n14950, n14951, n14952,
    n14953, n14954, n14955, n14956, n14957, n14958,
    n14959, n14960, n14961, n14962, n14963, n14964,
    n14965, n14966, n14967, n14968, n14969, n14970,
    n14971, n14972, n14973, n14974, n14975, n14976,
    n14977, n14978, n14979, n14980, n14981, n14982,
    n14983, n14984, n14985, n14986, n14987, n14988,
    n14989, n14990, n14991, n14992, n14993, n14994,
    n14995, n14996, n14997, n14998, n14999, n15000,
    n15001, n15002, n15003, n15004, n15005, n15006,
    n15007, n15008, n15009, n15010, n15011, n15012,
    n15013, n15014, n15015, n15016, n15017, n15018,
    n15019, n15020, n15021, n15022, n15023, n15024,
    n15025, n15026, n15027, n15028, n15029, n15030,
    n15031, n15032, n15033, n15034, n15035, n15036,
    n15037, n15038, n15039, n15040, n15041, n15042,
    n15043, n15044, n15045, n15046, n15047, n15048,
    n15049, n15050, n15051, n15052, n15053, n15054,
    n15055, n15056, n15057, n15058, n15059, n15061,
    n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073,
    n15074, n15075, n15076, n15077, n15078, n15079,
    n15080, n15081, n15082, n15083, n15084, n15085,
    n15086, n15087, n15088, n15089, n15090, n15091,
    n15092, n15093, n15094, n15095, n15096, n15097,
    n15098, n15099, n15100, n15101, n15102, n15103,
    n15104, n15105, n15106, n15107, n15108, n15109,
    n15110, n15111, n15112, n15113, n15114, n15115,
    n15116, n15117, n15118, n15119, n15120, n15121,
    n15122, n15123, n15124, n15125, n15126, n15127,
    n15128, n15129, n15130, n15131, n15132, n15133,
    n15134, n15135, n15136, n15137, n15138, n15139,
    n15140, n15141, n15142, n15143, n15144, n15145,
    n15146, n15147, n15148, n15149, n15150, n15151,
    n15152, n15153, n15154, n15155, n15156, n15157,
    n15158, n15159, n15160, n15161, n15162, n15163,
    n15164, n15165, n15166, n15167, n15168, n15169,
    n15170, n15171, n15172, n15173, n15174, n15175,
    n15176, n15177, n15178, n15179, n15180, n15181,
    n15182, n15183, n15184, n15185, n15186, n15187,
    n15188, n15189, n15190, n15191, n15192, n15193,
    n15194, n15195, n15196, n15197, n15198, n15199,
    n15200, n15201, n15202, n15203, n15204, n15205,
    n15206, n15208, n15209, n15210, n15211, n15212,
    n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230,
    n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248,
    n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260,
    n15261, n15262, n15263, n15264, n15265, n15266,
    n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278,
    n15279, n15280, n15281, n15282, n15283, n15284,
    n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296,
    n15297, n15298, n15299, n15300, n15301, n15302,
    n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314,
    n15315, n15316, n15317, n15318, n15319, n15320,
    n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332,
    n15333, n15334, n15335, n15336, n15337, n15338,
    n15339, n15340, n15341, n15342, n15344, n15345,
    n15346, n15347, n15348, n15349, n15350, n15351,
    n15352, n15353, n15354, n15355, n15356, n15357,
    n15358, n15359, n15360, n15361, n15362, n15363,
    n15364, n15365, n15366, n15367, n15368, n15369,
    n15370, n15371, n15372, n15373, n15374, n15375,
    n15376, n15377, n15378, n15379, n15380, n15381,
    n15382, n15383, n15384, n15385, n15386, n15387,
    n15388, n15389, n15390, n15391, n15392, n15393,
    n15394, n15395, n15396, n15397, n15398, n15399,
    n15400, n15401, n15402, n15403, n15404, n15405,
    n15406, n15407, n15408, n15409, n15410, n15411,
    n15412, n15413, n15414, n15415, n15416, n15417,
    n15418, n15419, n15420, n15421, n15422, n15423,
    n15424, n15425, n15426, n15427, n15428, n15429,
    n15430, n15431, n15432, n15433, n15434, n15435,
    n15436, n15437, n15438, n15439, n15440, n15441,
    n15442, n15443, n15444, n15445, n15446, n15447,
    n15448, n15449, n15450, n15451, n15452, n15453,
    n15454, n15455, n15456, n15457, n15458, n15459,
    n15460, n15461, n15462, n15463, n15464, n15465,
    n15466, n15467, n15468, n15469, n15470, n15471,
    n15472, n15473, n15474, n15475, n15476, n15477,
    n15478, n15479, n15480, n15481, n15482, n15484,
    n15485, n15486, n15487, n15488, n15489, n15490,
    n15491, n15492, n15493, n15494, n15495, n15496,
    n15497, n15498, n15499, n15500, n15501, n15502,
    n15503, n15504, n15505, n15506, n15507, n15508,
    n15509, n15510, n15511, n15512, n15513, n15514,
    n15515, n15516, n15517, n15518, n15519, n15520,
    n15521, n15522, n15523, n15524, n15525, n15526,
    n15527, n15528, n15529, n15530, n15531, n15532,
    n15533, n15534, n15535, n15536, n15537, n15538,
    n15539, n15540, n15541, n15542, n15543, n15544,
    n15545, n15546, n15547, n15548, n15549, n15550,
    n15551, n15552, n15553, n15554, n15555, n15556,
    n15557, n15558, n15559, n15560, n15561, n15562,
    n15563, n15564, n15565, n15566, n15567, n15568,
    n15569, n15570, n15571, n15572, n15573, n15574,
    n15575, n15576, n15577, n15578, n15579, n15580,
    n15581, n15582, n15583, n15584, n15585, n15586,
    n15587, n15588, n15589, n15590, n15591, n15592,
    n15593, n15594, n15595, n15596, n15597, n15598,
    n15599, n15600, n15601, n15602, n15603, n15604,
    n15605, n15606, n15607, n15608, n15609, n15610,
    n15611, n15612, n15613, n15614, n15616, n15617,
    n15618, n15619, n15620, n15621, n15622, n15623,
    n15624, n15625, n15626, n15627, n15628, n15629,
    n15630, n15631, n15632, n15633, n15634, n15635,
    n15636, n15637, n15638, n15639, n15640, n15641,
    n15642, n15643, n15644, n15645, n15646, n15647,
    n15648, n15649, n15650, n15651, n15652, n15653,
    n15654, n15655, n15656, n15657, n15658, n15659,
    n15660, n15661, n15662, n15663, n15664, n15665,
    n15666, n15667, n15668, n15669, n15670, n15671,
    n15672, n15673, n15674, n15675, n15676, n15677,
    n15678, n15679, n15680, n15681, n15682, n15683,
    n15684, n15685, n15686, n15687, n15688, n15689,
    n15690, n15691, n15692, n15693, n15694, n15695,
    n15696, n15697, n15698, n15699, n15700, n15701,
    n15702, n15703, n15704, n15705, n15706, n15707,
    n15708, n15709, n15710, n15711, n15712, n15713,
    n15714, n15715, n15716, n15717, n15718, n15719,
    n15720, n15721, n15722, n15723, n15724, n15725,
    n15726, n15727, n15728, n15729, n15730, n15731,
    n15732, n15733, n15734, n15735, n15736, n15737,
    n15738, n15739, n15740, n15741, n15743, n15744,
    n15745, n15746, n15747, n15748, n15749, n15750,
    n15751, n15752, n15753, n15754, n15755, n15756,
    n15757, n15758, n15759, n15760, n15761, n15762,
    n15763, n15764, n15765, n15766, n15767, n15768,
    n15769, n15770, n15771, n15772, n15773, n15774,
    n15775, n15776, n15777, n15778, n15779, n15780,
    n15781, n15782, n15783, n15784, n15785, n15786,
    n15787, n15788, n15789, n15790, n15791, n15792,
    n15793, n15794, n15795, n15796, n15797, n15798,
    n15799, n15800, n15801, n15802, n15803, n15804,
    n15805, n15806, n15807, n15808, n15809, n15810,
    n15811, n15812, n15813, n15814, n15815, n15816,
    n15817, n15818, n15819, n15820, n15821, n15822,
    n15823, n15824, n15825, n15826, n15827, n15828,
    n15829, n15830, n15831, n15832, n15833, n15834,
    n15835, n15836, n15837, n15838, n15839, n15840,
    n15841, n15842, n15843, n15844, n15845, n15846,
    n15847, n15848, n15849, n15850, n15851, n15852,
    n15853, n15854, n15855, n15856, n15857, n15858,
    n15859, n15860, n15862, n15863, n15864, n15865,
    n15866, n15867, n15868, n15869, n15870, n15871,
    n15872, n15873, n15874, n15875, n15876, n15877,
    n15878, n15879, n15880, n15881, n15882, n15883,
    n15884, n15885, n15886, n15887, n15888, n15889,
    n15890, n15891, n15892, n15893, n15894, n15895,
    n15896, n15897, n15898, n15899, n15900, n15901,
    n15902, n15903, n15904, n15905, n15906, n15907,
    n15908, n15909, n15910, n15911, n15912, n15913,
    n15914, n15915, n15916, n15917, n15918, n15919,
    n15920, n15921, n15922, n15923, n15924, n15925,
    n15926, n15927, n15928, n15929, n15930, n15931,
    n15932, n15933, n15934, n15935, n15936, n15937,
    n15938, n15939, n15940, n15941, n15942, n15943,
    n15944, n15945, n15946, n15947, n15948, n15949,
    n15950, n15951, n15952, n15953, n15954, n15955,
    n15956, n15957, n15958, n15959, n15960, n15961,
    n15962, n15963, n15964, n15965, n15966, n15967,
    n15968, n15969, n15970, n15971, n15972, n15973,
    n15974, n15975, n15976, n15977, n15978, n15979,
    n15980, n15981, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998,
    n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016,
    n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034,
    n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088,
    n16089, n16090, n16092, n16093, n16094, n16095,
    n16096, n16097, n16098, n16099, n16100, n16101,
    n16102, n16103, n16104, n16105, n16106, n16107,
    n16108, n16109, n16110, n16111, n16112, n16113,
    n16114, n16115, n16116, n16117, n16118, n16119,
    n16120, n16121, n16122, n16123, n16124, n16125,
    n16126, n16127, n16128, n16129, n16130, n16131,
    n16132, n16133, n16134, n16135, n16136, n16137,
    n16138, n16139, n16140, n16141, n16142, n16143,
    n16144, n16145, n16146, n16147, n16148, n16149,
    n16150, n16151, n16152, n16153, n16154, n16155,
    n16156, n16157, n16158, n16159, n16160, n16161,
    n16162, n16163, n16164, n16165, n16166, n16167,
    n16168, n16169, n16170, n16171, n16172, n16173,
    n16174, n16175, n16176, n16177, n16178, n16179,
    n16180, n16181, n16182, n16183, n16184, n16185,
    n16186, n16187, n16188, n16189, n16190, n16191,
    n16192, n16193, n16194, n16195, n16196, n16197,
    n16198, n16199, n16200, n16201, n16202, n16203,
    n16204, n16205, n16207, n16208, n16209, n16210,
    n16211, n16212, n16213, n16214, n16215, n16216,
    n16217, n16218, n16219, n16220, n16221, n16222,
    n16223, n16224, n16225, n16226, n16227, n16228,
    n16229, n16230, n16231, n16232, n16233, n16234,
    n16235, n16236, n16237, n16238, n16239, n16240,
    n16241, n16242, n16243, n16244, n16245, n16246,
    n16247, n16248, n16249, n16250, n16251, n16252,
    n16253, n16254, n16255, n16256, n16257, n16258,
    n16259, n16260, n16261, n16262, n16263, n16264,
    n16265, n16266, n16267, n16268, n16269, n16270,
    n16271, n16272, n16273, n16274, n16275, n16276,
    n16277, n16278, n16279, n16280, n16281, n16282,
    n16283, n16284, n16285, n16286, n16287, n16288,
    n16289, n16290, n16291, n16292, n16293, n16294,
    n16295, n16296, n16297, n16298, n16299, n16300,
    n16301, n16302, n16303, n16304, n16305, n16306,
    n16307, n16308, n16309, n16310, n16311, n16312,
    n16313, n16314, n16316, n16317, n16318, n16319,
    n16320, n16321, n16322, n16323, n16324, n16325,
    n16326, n16327, n16328, n16329, n16330, n16331,
    n16332, n16333, n16334, n16335, n16336, n16337,
    n16338, n16339, n16340, n16341, n16342, n16343,
    n16344, n16345, n16346, n16347, n16348, n16349,
    n16350, n16351, n16352, n16353, n16354, n16355,
    n16356, n16357, n16358, n16359, n16360, n16361,
    n16362, n16363, n16364, n16365, n16366, n16367,
    n16368, n16369, n16370, n16371, n16372, n16373,
    n16374, n16375, n16376, n16377, n16378, n16379,
    n16380, n16381, n16382, n16383, n16384, n16385,
    n16386, n16387, n16388, n16389, n16390, n16391,
    n16392, n16393, n16394, n16395, n16396, n16397,
    n16398, n16399, n16400, n16401, n16402, n16403,
    n16404, n16405, n16406, n16407, n16408, n16409,
    n16410, n16411, n16412, n16413, n16414, n16415,
    n16416, n16418, n16419, n16420, n16421, n16422,
    n16423, n16424, n16425, n16426, n16427, n16428,
    n16429, n16430, n16431, n16432, n16433, n16434,
    n16435, n16436, n16437, n16438, n16439, n16440,
    n16441, n16442, n16443, n16444, n16445, n16446,
    n16447, n16448, n16449, n16450, n16451, n16452,
    n16453, n16454, n16455, n16456, n16457, n16458,
    n16459, n16460, n16461, n16462, n16463, n16464,
    n16465, n16466, n16467, n16468, n16469, n16470,
    n16471, n16472, n16473, n16474, n16475, n16476,
    n16477, n16478, n16479, n16480, n16481, n16482,
    n16483, n16484, n16485, n16486, n16487, n16488,
    n16489, n16490, n16491, n16492, n16493, n16494,
    n16495, n16496, n16497, n16498, n16499, n16500,
    n16501, n16502, n16503, n16504, n16505, n16506,
    n16507, n16508, n16509, n16511, n16512, n16513,
    n16514, n16515, n16516, n16517, n16518, n16519,
    n16520, n16521, n16522, n16523, n16524, n16525,
    n16526, n16527, n16528, n16529, n16530, n16531,
    n16532, n16533, n16534, n16535, n16536, n16537,
    n16538, n16539, n16540, n16541, n16542, n16543,
    n16544, n16545, n16546, n16547, n16548, n16549,
    n16550, n16551, n16552, n16553, n16554, n16555,
    n16556, n16557, n16558, n16559, n16560, n16561,
    n16562, n16563, n16564, n16565, n16566, n16567,
    n16568, n16569, n16570, n16571, n16572, n16573,
    n16574, n16575, n16576, n16577, n16578, n16579,
    n16580, n16581, n16582, n16583, n16584, n16585,
    n16586, n16587, n16588, n16589, n16590, n16591,
    n16592, n16593, n16594, n16595, n16596, n16597,
    n16598, n16599, n16600, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622,
    n16623, n16624, n16625, n16626, n16627, n16628,
    n16629, n16630, n16631, n16632, n16633, n16634,
    n16635, n16636, n16637, n16638, n16639, n16640,
    n16641, n16642, n16643, n16644, n16645, n16646,
    n16647, n16648, n16649, n16650, n16651, n16652,
    n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664,
    n16665, n16666, n16667, n16668, n16669, n16670,
    n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682,
    n16683, n16684, n16685, n16686, n16688, n16689,
    n16690, n16691, n16692, n16693, n16694, n16695,
    n16696, n16697, n16698, n16699, n16700, n16701,
    n16702, n16703, n16704, n16705, n16706, n16707,
    n16708, n16709, n16710, n16711, n16712, n16713,
    n16714, n16715, n16716, n16717, n16718, n16719,
    n16720, n16721, n16722, n16723, n16724, n16725,
    n16726, n16727, n16728, n16729, n16730, n16731,
    n16732, n16733, n16734, n16735, n16736, n16737,
    n16738, n16739, n16740, n16741, n16742, n16743,
    n16744, n16745, n16746, n16747, n16748, n16749,
    n16750, n16751, n16752, n16753, n16754, n16755,
    n16756, n16757, n16758, n16759, n16760, n16761,
    n16762, n16763, n16764, n16765, n16766, n16767,
    n16768, n16769, n16770, n16772, n16773, n16774,
    n16775, n16776, n16777, n16778, n16779, n16780,
    n16781, n16782, n16783, n16784, n16785, n16786,
    n16787, n16788, n16789, n16790, n16791, n16792,
    n16793, n16794, n16795, n16796, n16797, n16798,
    n16799, n16800, n16801, n16802, n16803, n16804,
    n16805, n16806, n16807, n16808, n16809, n16810,
    n16811, n16812, n16813, n16814, n16815, n16816,
    n16817, n16818, n16819, n16820, n16821, n16822,
    n16823, n16824, n16825, n16826, n16827, n16828,
    n16829, n16830, n16831, n16832, n16833, n16834,
    n16835, n16836, n16837, n16838, n16839, n16840,
    n16841, n16842, n16843, n16844, n16845, n16846,
    n16847, n16848, n16849, n16851, n16852, n16853,
    n16854, n16855, n16856, n16857, n16858, n16859,
    n16860, n16861, n16862, n16863, n16864, n16865,
    n16866, n16867, n16868, n16869, n16870, n16871,
    n16872, n16873, n16874, n16875, n16876, n16877,
    n16878, n16879, n16880, n16881, n16882, n16883,
    n16884, n16885, n16886, n16887, n16888, n16889,
    n16890, n16891, n16892, n16893, n16894, n16895,
    n16896, n16897, n16898, n16899, n16900, n16901,
    n16902, n16903, n16904, n16905, n16906, n16907,
    n16908, n16909, n16910, n16911, n16912, n16913,
    n16914, n16915, n16916, n16917, n16918, n16919,
    n16920, n16921, n16922, n16923, n16924, n16926,
    n16927, n16928, n16929, n16930, n16931, n16932,
    n16933, n16934, n16935, n16936, n16937, n16938,
    n16939, n16940, n16941, n16942, n16943, n16944,
    n16945, n16946, n16947, n16948, n16949, n16950,
    n16951, n16952, n16953, n16954, n16955, n16956,
    n16957, n16958, n16959, n16960, n16961, n16962,
    n16963, n16964, n16965, n16966, n16967, n16968,
    n16969, n16970, n16971, n16972, n16973, n16974,
    n16975, n16976, n16977, n16978, n16979, n16980,
    n16981, n16982, n16983, n16984, n16985, n16986,
    n16987, n16988, n16989, n16990, n16991, n16992,
    n16993, n16994, n16996, n16997, n16998, n16999,
    n17000, n17001, n17002, n17003, n17004, n17005,
    n17006, n17007, n17008, n17009, n17010, n17011,
    n17012, n17013, n17014, n17015, n17016, n17017,
    n17018, n17019, n17020, n17021, n17022, n17023,
    n17024, n17025, n17026, n17027, n17028, n17029,
    n17030, n17031, n17032, n17033, n17034, n17035,
    n17036, n17037, n17038, n17039, n17040, n17041,
    n17042, n17043, n17044, n17045, n17046, n17047,
    n17048, n17049, n17050, n17051, n17052, n17053,
    n17054, n17055, n17056, n17057, n17058, n17059,
    n17060, n17061, n17063, n17064, n17065, n17066,
    n17067, n17068, n17069, n17070, n17071, n17072,
    n17073, n17074, n17075, n17076, n17077, n17078,
    n17079, n17080, n17081, n17082, n17083, n17084,
    n17085, n17086, n17087, n17088, n17089, n17090,
    n17091, n17092, n17093, n17094, n17095, n17096,
    n17097, n17098, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108,
    n17109, n17110, n17111, n17112, n17113, n17114,
    n17115, n17116, n17117, n17118, n17119, n17121,
    n17122, n17123, n17124, n17125, n17126, n17127,
    n17128, n17129, n17130, n17131, n17132, n17133,
    n17134, n17135, n17136, n17137, n17138, n17139,
    n17140, n17141, n17142, n17143, n17144, n17145,
    n17146, n17147, n17148, n17149, n17150, n17151,
    n17152, n17153, n17154, n17155, n17156, n17157,
    n17158, n17159, n17160, n17161, n17162, n17163,
    n17164, n17165, n17166, n17167, n17168, n17169,
    n17170, n17171, n17172, n17173, n17174, n17175,
    n17176, n17177, n17178, n17180, n17181, n17182,
    n17183, n17184, n17185, n17186, n17187, n17188,
    n17189, n17190, n17191, n17192, n17193, n17194,
    n17195, n17196, n17197, n17198, n17199, n17200,
    n17201, n17202, n17203, n17204, n17205, n17206,
    n17207, n17208, n17209, n17210, n17211, n17212,
    n17213, n17214, n17215, n17216, n17217, n17218,
    n17219, n17220, n17221, n17222, n17223, n17224,
    n17225, n17226, n17227, n17228, n17229, n17230,
    n17231, n17232, n17234, n17235, n17236, n17237,
    n17238, n17239, n17240, n17241, n17242, n17243,
    n17244, n17245, n17246, n17247, n17248, n17249,
    n17250, n17251, n17252, n17253, n17254, n17255,
    n17256, n17257, n17258, n17259, n17260, n17261,
    n17262, n17263, n17264, n17265, n17266, n17267,
    n17268, n17269, n17270, n17271, n17272, n17273,
    n17274, n17275, n17276, n17277, n17278, n17279,
    n17280, n17282, n17283, n17284, n17285, n17286,
    n17287, n17288, n17289, n17290, n17291, n17292,
    n17293, n17294, n17295, n17296, n17297, n17298,
    n17299, n17300, n17301, n17302, n17303, n17304,
    n17305, n17306, n17307, n17308, n17309, n17310,
    n17311, n17312, n17313, n17314, n17315, n17316,
    n17317, n17318, n17319, n17320, n17321, n17322,
    n17323, n17324, n17325, n17327, n17328, n17329,
    n17330, n17331, n17332, n17333, n17334, n17335,
    n17336, n17337, n17338, n17339, n17340, n17341,
    n17342, n17343, n17344, n17345, n17346, n17347,
    n17348, n17349, n17350, n17351, n17352, n17353,
    n17354, n17355, n17356, n17357, n17358, n17359,
    n17360, n17361, n17362, n17363, n17364, n17365,
    n17366, n17367, n17368, n17369, n17371, n17372,
    n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384,
    n17385, n17386, n17387, n17388, n17389, n17390,
    n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402,
    n17403, n17404, n17406, n17407, n17408, n17409,
    n17410, n17411, n17412, n17413, n17414, n17415,
    n17416, n17417, n17418, n17419, n17420, n17421,
    n17422, n17423, n17424, n17425, n17426, n17427,
    n17428, n17429, n17430, n17431, n17432, n17433,
    n17434, n17435, n17436, n17437, n17438, n17440,
    n17441, n17442, n17443, n17444, n17445, n17446,
    n17447, n17448, n17449, n17450, n17451, n17452,
    n17453, n17454, n17455, n17456, n17457, n17458,
    n17459, n17460, n17461, n17462, n17463, n17464,
    n17466, n17467, n17468, n17469, n17470, n17471,
    n17472, n17473, n17474, n17475, n17476, n17477,
    n17478, n17479, n17480, n17481, n17482, n17484,
    n17485, n17486, n17487, n17488, n17489, n17490,
    n17491, n17492, n17493, n17494, n17495, n17496,
    n17497, n17498, n17499, n17500, n17501, n17503,
    n17504, n17505, n17506, n17507, n17508, n17509,
    n17510, n17511, n17512, n17513, n17515, n17516,
    n17517, n17518, n17519, n17520, n17521, n17523,
    n17524, n17525, n17526;
  assign n194 = pi0  & pi1 ;
  assign po2  = pi1  & ~n194;
  assign n196 = pi0  & pi2 ;
  assign n197 = n194 & n196;
  assign n198 = ~n194 & ~n196;
  assign po3  = ~n197 & ~n198;
  assign n200 = pi1  & pi2 ;
  assign n201 = pi2  & ~n200;
  assign n202 = pi0  & pi3 ;
  assign n203 = ~n201 & ~n202;
  assign n204 = n201 & n202;
  assign n205 = ~n203 & ~n204;
  assign n206 = n197 & ~n205;
  assign n207 = ~n197 & n205;
  assign po4  = n206 | n207;
  assign n209 = pi3  & pi4 ;
  assign n210 = n194 & n209;
  assign n211 = pi1  & pi3 ;
  assign n212 = pi0  & pi4 ;
  assign n213 = ~n211 & ~n212;
  assign n214 = ~n210 & ~n213;
  assign n215 = ~n200 & ~n214;
  assign n216 = n200 & n214;
  assign n217 = ~n215 & ~n216;
  assign n218 = pi2  & pi3 ;
  assign n219 = pi0  & n218;
  assign n220 = ~n217 & ~n219;
  assign n221 = n217 & n219;
  assign po5  = ~n220 & ~n221;
  assign n223 = pi1  & pi4 ;
  assign n224 = pi0  & pi5 ;
  assign n225 = ~n223 & ~n224;
  assign n226 = pi4  & pi5 ;
  assign n227 = n194 & n226;
  assign n228 = n210 & ~n227;
  assign n229 = ~n227 & ~n228;
  assign n230 = ~n225 & n229;
  assign n231 = n210 & ~n228;
  assign n232 = ~n230 & ~n231;
  assign n233 = pi3  & ~n218;
  assign n234 = n232 & ~n233;
  assign n235 = ~n232 & n233;
  assign n236 = ~n234 & ~n235;
  assign n237 = ~n216 & ~n221;
  assign n238 = ~n236 & n237;
  assign n239 = ~n234 & ~n237;
  assign po6  = ~n238 & ~n239;
  assign n241 = ~n235 & ~n239;
  assign n242 = pi6  & n219;
  assign n243 = pi0  & pi6 ;
  assign n244 = ~n242 & n243;
  assign n245 = n218 & ~n242;
  assign n246 = ~n244 & ~n245;
  assign n247 = n200 & n226;
  assign n248 = pi1  & pi5 ;
  assign n249 = pi2  & pi4 ;
  assign n250 = ~n248 & ~n249;
  assign n251 = ~n247 & ~n250;
  assign n252 = n246 & ~n251;
  assign n253 = ~n246 & n251;
  assign n254 = ~n252 & ~n253;
  assign n255 = n229 & ~n254;
  assign n256 = ~n229 & n254;
  assign n257 = ~n255 & ~n256;
  assign n258 = n241 & ~n257;
  assign n259 = ~n241 & ~n255;
  assign n260 = ~n256 & n259;
  assign po7  = ~n258 & ~n260;
  assign n262 = pi2  & pi5 ;
  assign n263 = ~n209 & ~n262;
  assign n264 = n218 & n226;
  assign n265 = pi0  & pi7 ;
  assign n266 = ~n263 & n265;
  assign n267 = ~n264 & n266;
  assign n268 = ~n264 & ~n267;
  assign n269 = ~n263 & n268;
  assign n270 = n265 & ~n267;
  assign n271 = ~n269 & ~n270;
  assign n272 = ~n242 & ~n253;
  assign n273 = pi1  & pi6 ;
  assign n274 = n247 & ~n273;
  assign n275 = n247 & ~n274;
  assign n276 = ~pi4  & ~n273;
  assign n277 = pi4  & n273;
  assign n278 = ~n276 & ~n277;
  assign n279 = ~n274 & n278;
  assign n280 = ~n275 & ~n279;
  assign n281 = ~n272 & ~n280;
  assign n282 = n272 & n280;
  assign n283 = ~n281 & ~n282;
  assign n284 = n271 & ~n283;
  assign n285 = ~n271 & n283;
  assign n286 = ~n284 & ~n285;
  assign n287 = ~n256 & ~n259;
  assign n288 = ~n286 & n287;
  assign n289 = n286 & ~n287;
  assign po8  = ~n288 & ~n289;
  assign n291 = ~n274 & ~n281;
  assign n292 = pi1  & pi7 ;
  assign n293 = pi3  & pi5 ;
  assign n294 = n292 & n293;
  assign n295 = n292 & ~n294;
  assign n296 = n293 & ~n294;
  assign n297 = ~n295 & ~n296;
  assign n298 = ~n268 & ~n297;
  assign n299 = ~n268 & ~n298;
  assign n300 = ~n297 & ~n298;
  assign n301 = ~n299 & ~n300;
  assign n302 = pi0  & pi8 ;
  assign n303 = pi2  & pi6 ;
  assign n304 = ~n302 & ~n303;
  assign n305 = pi6  & pi8 ;
  assign n306 = n196 & n305;
  assign n307 = n277 & ~n304;
  assign n308 = ~n306 & n307;
  assign n309 = ~n306 & ~n308;
  assign n310 = ~n304 & n309;
  assign n311 = n277 & ~n308;
  assign n312 = ~n310 & ~n311;
  assign n313 = ~n301 & ~n312;
  assign n314 = n301 & n312;
  assign n315 = ~n313 & ~n314;
  assign n316 = n291 & ~n315;
  assign n317 = ~n291 & n315;
  assign n318 = ~n316 & ~n317;
  assign n319 = ~n285 & ~n289;
  assign n320 = ~n318 & n319;
  assign n321 = n318 & ~n319;
  assign po9  = ~n320 & ~n321;
  assign n323 = ~n298 & ~n313;
  assign n324 = pi3  & pi6 ;
  assign n325 = ~n226 & ~n324;
  assign n326 = pi5  & pi6 ;
  assign n327 = n209 & n326;
  assign n328 = pi2  & pi7 ;
  assign n329 = ~n325 & n328;
  assign n330 = ~n327 & n329;
  assign n331 = ~n327 & ~n330;
  assign n332 = ~n325 & n331;
  assign n333 = n328 & ~n330;
  assign n334 = ~n332 & ~n333;
  assign n335 = ~n309 & ~n334;
  assign n336 = ~n309 & ~n335;
  assign n337 = ~n334 & ~n335;
  assign n338 = ~n336 & ~n337;
  assign n339 = pi0  & pi9 ;
  assign n340 = n294 & ~n339;
  assign n341 = ~n294 & n339;
  assign n342 = ~n340 & ~n341;
  assign n343 = pi5  & pi8 ;
  assign n344 = pi1  & n343;
  assign n345 = pi5  & ~n344;
  assign n346 = pi1  & pi8 ;
  assign n347 = ~n344 & n346;
  assign n348 = ~n345 & ~n347;
  assign n349 = ~n342 & ~n348;
  assign n350 = n342 & n348;
  assign n351 = ~n349 & ~n350;
  assign n352 = ~n338 & n351;
  assign n353 = n338 & ~n351;
  assign n354 = ~n352 & ~n353;
  assign n355 = ~n323 & n354;
  assign n356 = n323 & ~n354;
  assign n357 = ~n355 & ~n356;
  assign n358 = ~n317 & ~n321;
  assign n359 = ~n357 & n358;
  assign n360 = n357 & ~n358;
  assign po10  = ~n359 & ~n360;
  assign n362 = ~n335 & ~n352;
  assign n363 = pi2  & pi8 ;
  assign n364 = pi0  & pi10 ;
  assign n365 = pi3  & pi7 ;
  assign n366 = n364 & n365;
  assign n367 = ~n364 & ~n365;
  assign n368 = n363 & ~n366;
  assign n369 = ~n367 & n368;
  assign n370 = n363 & ~n369;
  assign n371 = ~n366 & ~n369;
  assign n372 = ~n367 & n371;
  assign n373 = ~n370 & ~n372;
  assign n374 = n294 & n339;
  assign n375 = ~n349 & ~n374;
  assign n376 = ~n373 & n375;
  assign n377 = n373 & ~n375;
  assign n378 = ~n376 & ~n377;
  assign n379 = pi9  & n277;
  assign n380 = pi1  & pi9 ;
  assign n381 = pi4  & pi6 ;
  assign n382 = ~n380 & ~n381;
  assign n383 = ~n379 & ~n382;
  assign n384 = n344 & n383;
  assign n385 = n344 & ~n384;
  assign n386 = n383 & ~n384;
  assign n387 = ~n385 & ~n386;
  assign n388 = ~n331 & ~n387;
  assign n389 = n331 & ~n385;
  assign n390 = ~n386 & n389;
  assign n391 = ~n388 & ~n390;
  assign n392 = ~n378 & n391;
  assign n393 = n378 & ~n391;
  assign n394 = ~n392 & ~n393;
  assign n395 = n362 & ~n394;
  assign n396 = ~n362 & n394;
  assign n397 = ~n395 & ~n396;
  assign n398 = ~n355 & ~n360;
  assign n399 = ~n397 & n398;
  assign n400 = ~n395 & ~n398;
  assign n401 = ~n396 & n400;
  assign po11  = ~n399 & ~n401;
  assign n403 = ~n373 & ~n375;
  assign n404 = ~n392 & ~n403;
  assign n405 = pi10  & n273;
  assign n406 = pi6  & ~n405;
  assign n407 = pi1  & pi10 ;
  assign n408 = ~n405 & n407;
  assign n409 = ~n406 & ~n408;
  assign n410 = ~n371 & ~n409;
  assign n411 = ~n371 & ~n410;
  assign n412 = ~n409 & ~n410;
  assign n413 = ~n411 & ~n412;
  assign n414 = pi8  & pi9 ;
  assign n415 = n218 & n414;
  assign n416 = pi2  & pi9 ;
  assign n417 = pi3  & pi8 ;
  assign n418 = ~n416 & ~n417;
  assign n419 = ~n415 & ~n418;
  assign n420 = n379 & n419;
  assign n421 = n379 & ~n420;
  assign n422 = ~n415 & ~n420;
  assign n423 = ~n418 & n422;
  assign n424 = ~n421 & ~n423;
  assign n425 = ~n413 & ~n424;
  assign n426 = ~n413 & ~n425;
  assign n427 = ~n424 & ~n425;
  assign n428 = ~n426 & ~n427;
  assign n429 = ~n384 & ~n388;
  assign n430 = pi4  & pi7 ;
  assign n431 = ~n326 & ~n430;
  assign n432 = pi6  & pi7 ;
  assign n433 = n226 & n432;
  assign n434 = pi0  & pi11 ;
  assign n435 = ~n431 & n434;
  assign n436 = ~n433 & n435;
  assign n437 = ~n433 & ~n436;
  assign n438 = ~n431 & n437;
  assign n439 = n434 & ~n436;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~n429 & ~n440;
  assign n442 = ~n429 & ~n441;
  assign n443 = ~n440 & ~n441;
  assign n444 = ~n442 & ~n443;
  assign n445 = ~n428 & ~n444;
  assign n446 = n428 & n444;
  assign n447 = ~n445 & ~n446;
  assign n448 = n404 & ~n447;
  assign n449 = ~n404 & n447;
  assign n450 = ~n448 & ~n449;
  assign n451 = ~n396 & ~n400;
  assign n452 = ~n450 & n451;
  assign n453 = n450 & ~n451;
  assign po12  = ~n452 & ~n453;
  assign n455 = ~n441 & ~n445;
  assign n456 = n422 & n437;
  assign n457 = ~n422 & ~n437;
  assign n458 = ~n456 & ~n457;
  assign n459 = pi3  & pi9 ;
  assign n460 = pi10  & pi12 ;
  assign n461 = n196 & n460;
  assign n462 = pi0  & pi12 ;
  assign n463 = pi2  & pi10 ;
  assign n464 = ~n462 & ~n463;
  assign n465 = n459 & ~n461;
  assign n466 = ~n464 & n465;
  assign n467 = n459 & ~n466;
  assign n468 = ~n461 & ~n466;
  assign n469 = ~n464 & n468;
  assign n470 = ~n467 & ~n469;
  assign n471 = n458 & ~n470;
  assign n472 = n458 & ~n471;
  assign n473 = ~n470 & ~n471;
  assign n474 = ~n472 & ~n473;
  assign n475 = ~n410 & ~n425;
  assign n476 = pi4  & pi8 ;
  assign n477 = ~n405 & ~n476;
  assign n478 = n405 & n476;
  assign n479 = pi5  & pi11 ;
  assign n480 = n292 & n479;
  assign n481 = pi5  & pi7 ;
  assign n482 = pi1  & pi11 ;
  assign n483 = ~n481 & ~n482;
  assign n484 = ~n480 & ~n483;
  assign n485 = ~n477 & ~n478;
  assign n486 = n484 & n485;
  assign n487 = ~n478 & ~n486;
  assign n488 = ~n477 & n487;
  assign n489 = n484 & ~n486;
  assign n490 = ~n488 & ~n489;
  assign n491 = ~n475 & ~n490;
  assign n492 = n475 & n490;
  assign n493 = ~n491 & ~n492;
  assign n494 = ~n474 & n493;
  assign n495 = n474 & ~n493;
  assign n496 = ~n494 & ~n495;
  assign n497 = n455 & ~n496;
  assign n498 = ~n455 & n496;
  assign n499 = ~n497 & ~n498;
  assign n500 = ~n449 & ~n453;
  assign n501 = ~n499 & n500;
  assign n502 = ~n497 & ~n500;
  assign n503 = ~n498 & n502;
  assign po13  = ~n501 & ~n503;
  assign n505 = pi3  & pi10 ;
  assign n506 = pi9  & pi13 ;
  assign n507 = n212 & n506;
  assign n508 = pi0  & pi13 ;
  assign n509 = pi4  & pi9 ;
  assign n510 = ~n508 & ~n509;
  assign n511 = n505 & ~n507;
  assign n512 = ~n510 & n511;
  assign n513 = n505 & ~n512;
  assign n514 = ~n507 & ~n512;
  assign n515 = ~n510 & n514;
  assign n516 = ~n513 & ~n515;
  assign n517 = n487 & ~n516;
  assign n518 = ~n487 & n516;
  assign n519 = ~n517 & ~n518;
  assign n520 = pi2  & pi11 ;
  assign n521 = pi7  & pi8 ;
  assign n522 = n326 & n521;
  assign n523 = ~n343 & ~n432;
  assign n524 = n520 & ~n522;
  assign n525 = ~n523 & n524;
  assign n526 = n520 & ~n525;
  assign n527 = ~n522 & ~n525;
  assign n528 = ~n523 & n527;
  assign n529 = ~n526 & ~n528;
  assign n530 = ~n519 & ~n529;
  assign n531 = n519 & n529;
  assign n532 = ~n530 & ~n531;
  assign n533 = ~n457 & ~n471;
  assign n534 = ~pi12  & n480;
  assign n535 = pi12  & n292;
  assign n536 = pi1  & pi12 ;
  assign n537 = ~pi7  & ~n536;
  assign n538 = ~n535 & ~n537;
  assign n539 = ~n480 & ~n538;
  assign n540 = ~n534 & ~n539;
  assign n541 = ~n468 & n540;
  assign n542 = n468 & ~n540;
  assign n543 = ~n541 & ~n542;
  assign n544 = n533 & ~n543;
  assign n545 = ~n533 & n543;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~n491 & ~n494;
  assign n548 = ~n546 & n547;
  assign n549 = n546 & ~n547;
  assign n550 = ~n548 & ~n549;
  assign n551 = ~n532 & ~n550;
  assign n552 = n532 & n550;
  assign n553 = ~n551 & ~n552;
  assign n554 = ~n498 & ~n502;
  assign n555 = ~n553 & n554;
  assign n556 = n553 & ~n554;
  assign po14  = ~n555 & ~n556;
  assign n558 = ~n545 & ~n549;
  assign n559 = pi1  & pi13 ;
  assign n560 = ~n305 & ~n559;
  assign n561 = n305 & n559;
  assign n562 = ~n560 & ~n561;
  assign n563 = ~n527 & n562;
  assign n564 = ~n527 & ~n563;
  assign n565 = n562 & ~n563;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~n514 & ~n566;
  assign n568 = ~n514 & ~n567;
  assign n569 = ~n566 & ~n567;
  assign n570 = ~n568 & ~n569;
  assign n571 = ~n487 & ~n516;
  assign n572 = ~n530 & ~n571;
  assign n573 = n570 & n572;
  assign n574 = ~n570 & ~n572;
  assign n575 = ~n573 & ~n574;
  assign n576 = pi2  & pi12 ;
  assign n577 = pi3  & pi11 ;
  assign n578 = ~n576 & ~n577;
  assign n579 = pi11  & pi12 ;
  assign n580 = n218 & n579;
  assign n581 = pi0  & pi14 ;
  assign n582 = ~n578 & n581;
  assign n583 = ~n580 & n582;
  assign n584 = ~n580 & ~n583;
  assign n585 = ~n578 & n584;
  assign n586 = n581 & ~n583;
  assign n587 = ~n585 & ~n586;
  assign n588 = pi4  & pi10 ;
  assign n589 = pi5  & pi9 ;
  assign n590 = ~n588 & ~n589;
  assign n591 = pi9  & pi10 ;
  assign n592 = n226 & n591;
  assign n593 = n535 & ~n590;
  assign n594 = ~n592 & n593;
  assign n595 = n535 & ~n594;
  assign n596 = ~n592 & ~n594;
  assign n597 = ~n590 & n596;
  assign n598 = ~n595 & ~n597;
  assign n599 = ~n587 & ~n598;
  assign n600 = ~n587 & ~n599;
  assign n601 = ~n598 & ~n599;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~n534 & ~n541;
  assign n604 = n602 & n603;
  assign n605 = ~n602 & ~n603;
  assign n606 = ~n604 & ~n605;
  assign n607 = n575 & ~n606;
  assign n608 = ~n575 & n606;
  assign n609 = ~n607 & ~n608;
  assign n610 = ~n558 & ~n609;
  assign n611 = n558 & n609;
  assign n612 = ~n610 & ~n611;
  assign n613 = ~n552 & ~n556;
  assign n614 = ~n612 & n613;
  assign n615 = ~n611 & ~n613;
  assign n616 = ~n610 & n615;
  assign po15  = ~n614 & ~n616;
  assign n618 = ~n610 & ~n615;
  assign n619 = pi4  & pi11 ;
  assign n620 = ~n561 & ~n619;
  assign n621 = n561 & n619;
  assign n622 = pi1  & pi14 ;
  assign n623 = pi8  & ~n622;
  assign n624 = ~pi8  & n622;
  assign n625 = ~n623 & ~n624;
  assign n626 = ~n620 & ~n621;
  assign n627 = ~n625 & n626;
  assign n628 = ~n621 & ~n627;
  assign n629 = ~n620 & n628;
  assign n630 = ~n625 & ~n627;
  assign n631 = ~n629 & ~n630;
  assign n632 = pi2  & pi13 ;
  assign n633 = pi6  & pi9 ;
  assign n634 = n521 & n633;
  assign n635 = ~n521 & ~n633;
  assign n636 = n632 & ~n634;
  assign n637 = ~n635 & n636;
  assign n638 = n632 & ~n637;
  assign n639 = ~n634 & ~n637;
  assign n640 = ~n635 & n639;
  assign n641 = ~n638 & ~n640;
  assign n642 = ~n631 & ~n641;
  assign n643 = ~n631 & ~n642;
  assign n644 = ~n641 & ~n642;
  assign n645 = ~n643 & ~n644;
  assign n646 = ~n563 & ~n567;
  assign n647 = n645 & n646;
  assign n648 = ~n645 & ~n646;
  assign n649 = ~n647 & ~n648;
  assign n650 = n584 & n596;
  assign n651 = ~n584 & ~n596;
  assign n652 = ~n650 & ~n651;
  assign n653 = pi5  & pi10 ;
  assign n654 = pi0  & pi15 ;
  assign n655 = pi3  & pi12 ;
  assign n656 = n654 & n655;
  assign n657 = ~n654 & ~n655;
  assign n658 = n653 & ~n656;
  assign n659 = ~n657 & n658;
  assign n660 = n653 & ~n659;
  assign n661 = ~n656 & ~n659;
  assign n662 = ~n657 & n661;
  assign n663 = ~n660 & ~n662;
  assign n664 = n652 & ~n663;
  assign n665 = n652 & ~n664;
  assign n666 = ~n663 & ~n664;
  assign n667 = ~n665 & ~n666;
  assign n668 = ~n599 & ~n605;
  assign n669 = n667 & n668;
  assign n670 = ~n667 & ~n668;
  assign n671 = ~n669 & ~n670;
  assign n672 = n649 & ~n671;
  assign n673 = ~n649 & n671;
  assign n674 = ~n672 & ~n673;
  assign n675 = ~n573 & ~n607;
  assign n676 = ~n674 & n675;
  assign n677 = n674 & ~n675;
  assign n678 = ~n676 & ~n677;
  assign n679 = ~n618 & ~n678;
  assign n680 = n618 & n678;
  assign po16  = n679 | n680;
  assign n682 = n628 & n661;
  assign n683 = ~n628 & ~n661;
  assign n684 = ~n682 & ~n683;
  assign n685 = pi6  & pi16 ;
  assign n686 = n364 & n685;
  assign n687 = pi0  & pi16 ;
  assign n688 = pi6  & pi10 ;
  assign n689 = ~n687 & ~n688;
  assign n690 = n479 & ~n686;
  assign n691 = ~n689 & n690;
  assign n692 = n479 & ~n691;
  assign n693 = ~n686 & ~n691;
  assign n694 = ~n689 & n693;
  assign n695 = ~n692 & ~n694;
  assign n696 = n684 & ~n695;
  assign n697 = n684 & ~n696;
  assign n698 = ~n695 & ~n696;
  assign n699 = ~n697 & ~n698;
  assign n700 = ~n642 & ~n648;
  assign n701 = n699 & n700;
  assign n702 = ~n699 & ~n700;
  assign n703 = ~n701 & ~n702;
  assign n704 = ~n651 & ~n664;
  assign n705 = pi4  & pi12 ;
  assign n706 = pi13  & pi14 ;
  assign n707 = n218 & n706;
  assign n708 = pi3  & pi13 ;
  assign n709 = pi2  & pi14 ;
  assign n710 = ~n708 & ~n709;
  assign n711 = n705 & ~n707;
  assign n712 = ~n710 & n711;
  assign n713 = n705 & ~n712;
  assign n714 = ~n707 & ~n712;
  assign n715 = ~n710 & n714;
  assign n716 = ~n713 & ~n715;
  assign n717 = ~n704 & ~n716;
  assign n718 = ~n704 & ~n717;
  assign n719 = ~n716 & ~n717;
  assign n720 = ~n718 & ~n719;
  assign n721 = pi8  & n622;
  assign n722 = pi7  & pi9 ;
  assign n723 = pi1  & pi15 ;
  assign n724 = n722 & n723;
  assign n725 = ~n722 & ~n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = n721 & n726;
  assign n728 = n721 & ~n727;
  assign n729 = ~n721 & n726;
  assign n730 = ~n728 & ~n729;
  assign n731 = ~n639 & ~n730;
  assign n732 = ~n639 & ~n731;
  assign n733 = ~n730 & ~n731;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~n720 & ~n734;
  assign n736 = ~n720 & ~n735;
  assign n737 = ~n734 & ~n735;
  assign n738 = ~n736 & ~n737;
  assign n739 = ~n703 & n738;
  assign n740 = n703 & ~n738;
  assign n741 = ~n739 & ~n740;
  assign n742 = ~n669 & ~n673;
  assign n743 = n741 & n742;
  assign n744 = ~n741 & ~n742;
  assign n745 = ~n743 & ~n744;
  assign n746 = ~n618 & ~n677;
  assign n747 = ~n676 & ~n746;
  assign n748 = ~n745 & n747;
  assign n749 = n745 & ~n747;
  assign po17  = ~n748 & ~n749;
  assign n751 = ~n702 & ~n740;
  assign n752 = pi5  & pi12 ;
  assign n753 = pi0  & pi17 ;
  assign n754 = ~n752 & ~n753;
  assign n755 = n752 & n753;
  assign n756 = n724 & ~n754;
  assign n757 = ~n755 & n756;
  assign n758 = ~n755 & ~n757;
  assign n759 = ~n754 & n758;
  assign n760 = n724 & ~n757;
  assign n761 = ~n759 & ~n760;
  assign n762 = pi3  & pi14 ;
  assign n763 = n521 & n591;
  assign n764 = pi7  & pi10 ;
  assign n765 = ~n414 & ~n764;
  assign n766 = n762 & ~n763;
  assign n767 = ~n765 & n766;
  assign n768 = n762 & ~n767;
  assign n769 = ~n763 & ~n767;
  assign n770 = ~n765 & n769;
  assign n771 = ~n768 & ~n770;
  assign n772 = ~n761 & ~n771;
  assign n773 = ~n761 & ~n772;
  assign n774 = ~n771 & ~n772;
  assign n775 = ~n773 & ~n774;
  assign n776 = pi6  & pi11 ;
  assign n777 = pi13  & pi15 ;
  assign n778 = n249 & n777;
  assign n779 = pi2  & pi15 ;
  assign n780 = pi4  & pi13 ;
  assign n781 = ~n779 & ~n780;
  assign n782 = n776 & ~n778;
  assign n783 = ~n781 & n782;
  assign n784 = n776 & ~n783;
  assign n785 = ~n778 & ~n783;
  assign n786 = ~n781 & n785;
  assign n787 = ~n784 & ~n786;
  assign n788 = ~n775 & ~n787;
  assign n789 = ~n775 & ~n788;
  assign n790 = ~n787 & ~n788;
  assign n791 = ~n789 & ~n790;
  assign n792 = ~n717 & ~n735;
  assign n793 = n791 & n792;
  assign n794 = ~n791 & ~n792;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~n727 & ~n731;
  assign n797 = ~n683 & ~n696;
  assign n798 = n796 & n797;
  assign n799 = ~n796 & ~n797;
  assign n800 = ~n798 & ~n799;
  assign n801 = pi1  & pi16 ;
  assign n802 = ~pi9  & ~n801;
  assign n803 = pi9  & pi16 ;
  assign n804 = pi1  & n803;
  assign n805 = ~n802 & ~n804;
  assign n806 = ~n714 & n805;
  assign n807 = ~n714 & ~n806;
  assign n808 = n805 & ~n806;
  assign n809 = ~n807 & ~n808;
  assign n810 = ~n693 & ~n809;
  assign n811 = ~n693 & ~n810;
  assign n812 = ~n809 & ~n810;
  assign n813 = ~n811 & ~n812;
  assign n814 = ~n800 & n813;
  assign n815 = n800 & ~n813;
  assign n816 = ~n814 & ~n815;
  assign n817 = n795 & n816;
  assign n818 = ~n795 & ~n816;
  assign n819 = ~n817 & ~n818;
  assign n820 = ~n751 & n819;
  assign n821 = n751 & ~n819;
  assign n822 = ~n820 & ~n821;
  assign n823 = ~n743 & ~n749;
  assign n824 = ~n822 & n823;
  assign n825 = n822 & ~n823;
  assign po18  = ~n824 & ~n825;
  assign n827 = ~n794 & ~n817;
  assign n828 = pi0  & pi18 ;
  assign n829 = pi5  & pi13 ;
  assign n830 = ~n828 & ~n829;
  assign n831 = n828 & n829;
  assign n832 = pi7  & pi11 ;
  assign n833 = ~n830 & n832;
  assign n834 = ~n831 & n833;
  assign n835 = ~n831 & ~n834;
  assign n836 = ~n830 & n835;
  assign n837 = n832 & ~n834;
  assign n838 = ~n836 & ~n837;
  assign n839 = pi4  & pi14 ;
  assign n840 = pi15  & pi16 ;
  assign n841 = n218 & n840;
  assign n842 = pi3  & pi15 ;
  assign n843 = pi2  & pi16 ;
  assign n844 = ~n842 & ~n843;
  assign n845 = n839 & ~n841;
  assign n846 = ~n844 & n845;
  assign n847 = n839 & ~n846;
  assign n848 = ~n841 & ~n846;
  assign n849 = ~n844 & n848;
  assign n850 = ~n847 & ~n849;
  assign n851 = ~n838 & ~n850;
  assign n852 = ~n838 & ~n851;
  assign n853 = ~n850 & ~n851;
  assign n854 = ~n852 & ~n853;
  assign n855 = pi8  & pi10 ;
  assign n856 = pi1  & pi17 ;
  assign n857 = n855 & n856;
  assign n858 = n855 & ~n857;
  assign n859 = ~n855 & n856;
  assign n860 = ~n858 & ~n859;
  assign n861 = pi6  & pi12 ;
  assign n862 = ~n804 & ~n861;
  assign n863 = n804 & n861;
  assign n864 = ~n862 & ~n863;
  assign n865 = ~n860 & n864;
  assign n866 = ~n860 & ~n865;
  assign n867 = ~n863 & ~n865;
  assign n868 = ~n862 & n867;
  assign n869 = ~n866 & ~n868;
  assign n870 = ~n854 & ~n869;
  assign n871 = ~n854 & ~n870;
  assign n872 = ~n869 & ~n870;
  assign n873 = ~n871 & ~n872;
  assign n874 = ~n799 & ~n815;
  assign n875 = ~n873 & ~n874;
  assign n876 = ~n873 & ~n875;
  assign n877 = ~n874 & ~n875;
  assign n878 = ~n876 & ~n877;
  assign n879 = n769 & n785;
  assign n880 = ~n769 & ~n785;
  assign n881 = ~n879 & ~n880;
  assign n882 = n758 & ~n881;
  assign n883 = ~n758 & n881;
  assign n884 = ~n882 & ~n883;
  assign n885 = ~n806 & ~n810;
  assign n886 = ~n772 & ~n788;
  assign n887 = n885 & n886;
  assign n888 = ~n885 & ~n886;
  assign n889 = ~n887 & ~n888;
  assign n890 = n884 & n889;
  assign n891 = ~n884 & ~n889;
  assign n892 = ~n890 & ~n891;
  assign n893 = ~n878 & n892;
  assign n894 = n878 & ~n892;
  assign n895 = ~n893 & ~n894;
  assign n896 = ~n827 & n895;
  assign n897 = n827 & ~n895;
  assign n898 = ~n896 & ~n897;
  assign n899 = ~n820 & ~n825;
  assign n900 = ~n898 & n899;
  assign n901 = ~n897 & ~n899;
  assign n902 = ~n896 & n901;
  assign po19  = ~n900 & ~n902;
  assign n904 = n835 & n867;
  assign n905 = ~n835 & ~n867;
  assign n906 = ~n904 & ~n905;
  assign n907 = pi3  & pi16 ;
  assign n908 = pi8  & pi11 ;
  assign n909 = n591 & n908;
  assign n910 = ~n591 & ~n908;
  assign n911 = n907 & ~n909;
  assign n912 = ~n910 & n911;
  assign n913 = n907 & ~n912;
  assign n914 = ~n909 & ~n912;
  assign n915 = ~n910 & n914;
  assign n916 = ~n913 & ~n915;
  assign n917 = n906 & ~n916;
  assign n918 = n906 & ~n917;
  assign n919 = ~n916 & ~n917;
  assign n920 = ~n918 & ~n919;
  assign n921 = ~n851 & ~n870;
  assign n922 = pi1  & pi18 ;
  assign n923 = n857 & ~n922;
  assign n924 = n857 & ~n923;
  assign n925 = ~pi10  & ~n922;
  assign n926 = pi10  & n922;
  assign n927 = ~n925 & ~n926;
  assign n928 = ~n923 & n927;
  assign n929 = ~n924 & ~n928;
  assign n930 = ~n848 & ~n929;
  assign n931 = n848 & n929;
  assign n932 = ~n930 & ~n931;
  assign n933 = ~n921 & n932;
  assign n934 = n921 & ~n932;
  assign n935 = ~n933 & ~n934;
  assign n936 = ~n920 & n935;
  assign n937 = n920 & ~n935;
  assign n938 = ~n936 & ~n937;
  assign n939 = pi2  & pi17 ;
  assign n940 = pi4  & pi15 ;
  assign n941 = ~n939 & ~n940;
  assign n942 = pi15  & pi17 ;
  assign n943 = n249 & n942;
  assign n944 = pi0  & pi19 ;
  assign n945 = ~n941 & n944;
  assign n946 = ~n943 & n945;
  assign n947 = ~n943 & ~n946;
  assign n948 = ~n941 & n947;
  assign n949 = n944 & ~n946;
  assign n950 = ~n948 & ~n949;
  assign n951 = pi5  & pi14 ;
  assign n952 = pi12  & pi13 ;
  assign n953 = n432 & n952;
  assign n954 = pi6  & pi13 ;
  assign n955 = pi7  & pi12 ;
  assign n956 = ~n954 & ~n955;
  assign n957 = n951 & ~n953;
  assign n958 = ~n956 & n957;
  assign n959 = n951 & ~n958;
  assign n960 = ~n953 & ~n958;
  assign n961 = ~n956 & n960;
  assign n962 = ~n959 & ~n961;
  assign n963 = ~n950 & ~n962;
  assign n964 = ~n950 & ~n963;
  assign n965 = ~n962 & ~n963;
  assign n966 = ~n964 & ~n965;
  assign n967 = ~n880 & ~n883;
  assign n968 = n966 & n967;
  assign n969 = ~n966 & ~n967;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~n888 & ~n890;
  assign n972 = n970 & ~n971;
  assign n973 = ~n970 & n971;
  assign n974 = ~n972 & ~n973;
  assign n975 = n938 & n974;
  assign n976 = ~n938 & ~n974;
  assign n977 = ~n975 & ~n976;
  assign n978 = ~n875 & ~n893;
  assign n979 = ~n977 & n978;
  assign n980 = n977 & ~n978;
  assign n981 = ~n979 & ~n980;
  assign n982 = ~n896 & ~n901;
  assign n983 = ~n981 & n982;
  assign n984 = n981 & ~n982;
  assign po20  = ~n983 & ~n984;
  assign n986 = ~n972 & ~n975;
  assign n987 = ~n923 & ~n930;
  assign n988 = pi2  & pi18 ;
  assign n989 = pi16  & pi17 ;
  assign n990 = n209 & n989;
  assign n991 = pi3  & pi17 ;
  assign n992 = pi4  & pi16 ;
  assign n993 = ~n991 & ~n992;
  assign n994 = n988 & ~n990;
  assign n995 = ~n993 & n994;
  assign n996 = n988 & ~n995;
  assign n997 = ~n990 & ~n995;
  assign n998 = ~n993 & n997;
  assign n999 = ~n996 & ~n998;
  assign n1000 = ~n987 & ~n999;
  assign n1001 = ~n987 & ~n1000;
  assign n1002 = ~n999 & ~n1000;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = ~n905 & ~n917;
  assign n1005 = n1003 & n1004;
  assign n1006 = ~n1003 & ~n1004;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = ~n933 & ~n936;
  assign n1009 = ~n1007 & n1008;
  assign n1010 = n1007 & ~n1008;
  assign n1011 = ~n1009 & ~n1010;
  assign n1012 = pi9  & pi11 ;
  assign n1013 = pi1  & pi19 ;
  assign n1014 = ~n1012 & ~n1013;
  assign n1015 = n1012 & n1013;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = ~n914 & n1016;
  assign n1018 = ~n914 & ~n1017;
  assign n1019 = n1016 & ~n1017;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = ~n947 & ~n1020;
  assign n1022 = ~n947 & ~n1021;
  assign n1023 = ~n1020 & ~n1021;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = ~n963 & ~n969;
  assign n1026 = n1024 & n1025;
  assign n1027 = ~n1024 & ~n1025;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = pi0  & pi20 ;
  assign n1030 = pi7  & pi13 ;
  assign n1031 = ~n1029 & ~n1030;
  assign n1032 = n1029 & n1030;
  assign n1033 = ~n1031 & ~n1032;
  assign n1034 = n926 & n1033;
  assign n1035 = ~n926 & ~n1033;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = ~n960 & n1036;
  assign n1038 = n960 & ~n1036;
  assign n1039 = ~n1037 & ~n1038;
  assign n1040 = pi8  & pi12 ;
  assign n1041 = pi14  & pi15 ;
  assign n1042 = n326 & n1041;
  assign n1043 = pi5  & pi15 ;
  assign n1044 = pi6  & pi14 ;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = n1040 & ~n1042;
  assign n1047 = ~n1045 & n1046;
  assign n1048 = n1040 & ~n1047;
  assign n1049 = ~n1042 & ~n1047;
  assign n1050 = ~n1045 & n1049;
  assign n1051 = ~n1048 & ~n1050;
  assign n1052 = n1039 & ~n1051;
  assign n1053 = n1039 & ~n1052;
  assign n1054 = ~n1051 & ~n1052;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = n1028 & ~n1055;
  assign n1057 = ~n1028 & n1055;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = n1011 & n1058;
  assign n1060 = n1011 & ~n1059;
  assign n1061 = n1058 & ~n1059;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~n986 & ~n1062;
  assign n1064 = n986 & n1062;
  assign n1065 = ~n1063 & ~n1064;
  assign n1066 = ~n980 & ~n984;
  assign n1067 = n1065 & ~n1066;
  assign n1068 = ~n1065 & n1066;
  assign po21  = ~n1067 & ~n1068;
  assign n1070 = ~n1010 & ~n1059;
  assign n1071 = n997 & n1049;
  assign n1072 = ~n997 & ~n1049;
  assign n1073 = ~n1071 & ~n1072;
  assign n1074 = ~n1032 & ~n1034;
  assign n1075 = ~n1073 & n1074;
  assign n1076 = n1073 & ~n1074;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~n1000 & ~n1006;
  assign n1079 = ~n1077 & n1078;
  assign n1080 = n1077 & ~n1078;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = pi2  & pi19 ;
  assign n1083 = pi3  & pi18 ;
  assign n1084 = ~n1082 & ~n1083;
  assign n1085 = pi18  & pi19 ;
  assign n1086 = n218 & n1085;
  assign n1087 = pi5  & pi16 ;
  assign n1088 = ~n1084 & n1087;
  assign n1089 = ~n1086 & n1088;
  assign n1090 = ~n1086 & ~n1089;
  assign n1091 = ~n1084 & n1090;
  assign n1092 = n1087 & ~n1089;
  assign n1093 = ~n1091 & ~n1092;
  assign n1094 = pi6  & pi15 ;
  assign n1095 = n521 & n706;
  assign n1096 = pi7  & pi14 ;
  assign n1097 = pi8  & pi13 ;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = n1094 & ~n1095;
  assign n1100 = ~n1098 & n1099;
  assign n1101 = n1094 & ~n1100;
  assign n1102 = ~n1095 & ~n1100;
  assign n1103 = ~n1098 & n1102;
  assign n1104 = ~n1101 & ~n1103;
  assign n1105 = ~n1093 & ~n1104;
  assign n1106 = ~n1093 & ~n1105;
  assign n1107 = ~n1104 & ~n1105;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = pi4  & pi17 ;
  assign n1110 = n579 & n591;
  assign n1111 = pi10  & pi11 ;
  assign n1112 = pi9  & pi12 ;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = n1109 & ~n1110;
  assign n1115 = ~n1113 & n1114;
  assign n1116 = n1109 & ~n1115;
  assign n1117 = ~n1110 & ~n1115;
  assign n1118 = ~n1113 & n1117;
  assign n1119 = ~n1116 & ~n1118;
  assign n1120 = ~n1108 & ~n1119;
  assign n1121 = ~n1108 & ~n1120;
  assign n1122 = ~n1119 & ~n1120;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = ~n1081 & n1123;
  assign n1125 = n1081 & ~n1123;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = ~n1017 & ~n1021;
  assign n1128 = pi0  & pi21 ;
  assign n1129 = n1015 & ~n1128;
  assign n1130 = ~n1015 & n1128;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = pi1  & pi20 ;
  assign n1133 = pi11  & n1132;
  assign n1134 = pi11  & ~n1133;
  assign n1135 = n1132 & ~n1133;
  assign n1136 = ~n1134 & ~n1135;
  assign n1137 = ~n1131 & ~n1136;
  assign n1138 = n1131 & n1136;
  assign n1139 = ~n1137 & ~n1138;
  assign n1140 = n1127 & ~n1139;
  assign n1141 = ~n1127 & n1139;
  assign n1142 = ~n1140 & ~n1141;
  assign n1143 = ~n1037 & ~n1052;
  assign n1144 = ~n1142 & n1143;
  assign n1145 = n1142 & ~n1143;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = ~n1027 & ~n1056;
  assign n1148 = n1146 & ~n1147;
  assign n1149 = ~n1146 & n1147;
  assign n1150 = ~n1148 & ~n1149;
  assign n1151 = n1126 & n1150;
  assign n1152 = ~n1126 & ~n1150;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~n1070 & n1153;
  assign n1155 = n1070 & ~n1153;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = ~n1063 & ~n1067;
  assign n1158 = ~n1156 & n1157;
  assign n1159 = n1156 & ~n1157;
  assign po22  = ~n1158 & ~n1159;
  assign n1161 = ~n1148 & ~n1151;
  assign n1162 = n1090 & n1102;
  assign n1163 = ~n1090 & ~n1102;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = n1015 & n1128;
  assign n1166 = ~n1137 & ~n1165;
  assign n1167 = ~n1164 & n1166;
  assign n1168 = n1164 & ~n1166;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = ~n1141 & ~n1145;
  assign n1171 = ~n1169 & n1170;
  assign n1172 = n1169 & ~n1170;
  assign n1173 = ~n1171 & ~n1172;
  assign n1174 = pi7  & pi15 ;
  assign n1175 = pi8  & pi14 ;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = n521 & n1041;
  assign n1178 = pi0  & pi22 ;
  assign n1179 = ~n1176 & n1178;
  assign n1180 = ~n1177 & n1179;
  assign n1181 = ~n1177 & ~n1180;
  assign n1182 = ~n1176 & n1181;
  assign n1183 = n1178 & ~n1180;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = pi2  & pi20 ;
  assign n1186 = n685 & n1185;
  assign n1187 = ~n685 & ~n1185;
  assign n1188 = n506 & ~n1186;
  assign n1189 = ~n1187 & n1188;
  assign n1190 = n506 & ~n1189;
  assign n1191 = ~n1186 & ~n1189;
  assign n1192 = ~n1187 & n1191;
  assign n1193 = ~n1190 & ~n1192;
  assign n1194 = ~n1184 & ~n1193;
  assign n1195 = ~n1184 & ~n1194;
  assign n1196 = ~n1193 & ~n1194;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = pi3  & pi19 ;
  assign n1199 = pi17  & pi18 ;
  assign n1200 = n226 & n1199;
  assign n1201 = pi5  & pi17 ;
  assign n1202 = pi4  & pi18 ;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = n1198 & ~n1200;
  assign n1205 = ~n1203 & n1204;
  assign n1206 = n1198 & ~n1205;
  assign n1207 = ~n1200 & ~n1205;
  assign n1208 = ~n1203 & n1207;
  assign n1209 = ~n1206 & ~n1208;
  assign n1210 = ~n1197 & ~n1209;
  assign n1211 = ~n1197 & ~n1210;
  assign n1212 = ~n1209 & ~n1210;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = ~n1173 & n1213;
  assign n1215 = n1173 & ~n1213;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = ~n1080 & ~n1125;
  assign n1218 = ~n1105 & ~n1120;
  assign n1219 = ~n1072 & ~n1076;
  assign n1220 = pi1  & pi21 ;
  assign n1221 = n460 & n1220;
  assign n1222 = ~n460 & ~n1220;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = n1133 & n1223;
  assign n1225 = ~n1133 & ~n1223;
  assign n1226 = ~n1224 & ~n1225;
  assign n1227 = ~n1117 & n1226;
  assign n1228 = n1117 & ~n1226;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~n1219 & n1229;
  assign n1231 = ~n1219 & ~n1230;
  assign n1232 = n1229 & ~n1230;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = ~n1218 & ~n1233;
  assign n1235 = n1218 & n1233;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = ~n1217 & n1236;
  assign n1238 = ~n1217 & ~n1237;
  assign n1239 = n1236 & ~n1237;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = n1216 & ~n1240;
  assign n1242 = ~n1216 & n1240;
  assign n1243 = ~n1241 & ~n1242;
  assign n1244 = ~n1161 & n1243;
  assign n1245 = n1161 & ~n1243;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = ~n1154 & ~n1159;
  assign n1248 = ~n1246 & n1247;
  assign n1249 = ~n1245 & ~n1247;
  assign n1250 = ~n1244 & n1249;
  assign po23  = ~n1248 & ~n1250;
  assign n1252 = ~n1237 & ~n1241;
  assign n1253 = ~n1230 & ~n1234;
  assign n1254 = pi3  & pi20 ;
  assign n1255 = pi5  & pi18 ;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = pi18  & pi20 ;
  assign n1258 = n293 & n1257;
  assign n1259 = pi6  & pi17 ;
  assign n1260 = ~n1256 & n1259;
  assign n1261 = ~n1258 & n1260;
  assign n1262 = ~n1258 & ~n1261;
  assign n1263 = ~n1256 & n1262;
  assign n1264 = n1259 & ~n1261;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = pi4  & pi19 ;
  assign n1267 = n952 & n1111;
  assign n1268 = pi10  & pi13 ;
  assign n1269 = ~n579 & ~n1268;
  assign n1270 = n1266 & ~n1267;
  assign n1271 = ~n1269 & n1270;
  assign n1272 = n1266 & ~n1271;
  assign n1273 = ~n1267 & ~n1271;
  assign n1274 = ~n1269 & n1273;
  assign n1275 = ~n1272 & ~n1274;
  assign n1276 = ~n1265 & ~n1275;
  assign n1277 = ~n1265 & ~n1276;
  assign n1278 = ~n1275 & ~n1276;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = ~n1224 & ~n1227;
  assign n1281 = n1279 & n1280;
  assign n1282 = ~n1279 & ~n1280;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = pi0  & pi23 ;
  assign n1285 = pi2  & pi21 ;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = pi21  & pi23 ;
  assign n1288 = n196 & n1287;
  assign n1289 = n1221 & ~n1286;
  assign n1290 = ~n1288 & n1289;
  assign n1291 = ~n1288 & ~n1290;
  assign n1292 = ~n1286 & n1291;
  assign n1293 = n1221 & ~n1290;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = n1181 & ~n1294;
  assign n1296 = ~n1181 & n1294;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = pi7  & pi16 ;
  assign n1299 = n414 & n1041;
  assign n1300 = pi8  & pi15 ;
  assign n1301 = pi9  & pi14 ;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = n1298 & ~n1299;
  assign n1304 = ~n1302 & n1303;
  assign n1305 = n1298 & ~n1304;
  assign n1306 = ~n1299 & ~n1304;
  assign n1307 = ~n1302 & n1306;
  assign n1308 = ~n1305 & ~n1307;
  assign n1309 = ~n1297 & ~n1308;
  assign n1310 = n1297 & n1308;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = ~n1283 & ~n1311;
  assign n1313 = n1283 & n1311;
  assign n1314 = ~n1312 & ~n1313;
  assign n1315 = ~n1253 & n1314;
  assign n1316 = n1253 & ~n1314;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = ~n1172 & ~n1215;
  assign n1319 = ~n1163 & ~n1168;
  assign n1320 = ~n1194 & ~n1210;
  assign n1321 = n1319 & n1320;
  assign n1322 = ~n1319 & ~n1320;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = pi1  & pi22 ;
  assign n1325 = pi12  & n1324;
  assign n1326 = ~pi12  & ~n1324;
  assign n1327 = ~n1325 & ~n1326;
  assign n1328 = n1207 & ~n1327;
  assign n1329 = ~n1207 & n1327;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = ~n1191 & n1330;
  assign n1332 = n1191 & ~n1330;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = n1323 & n1333;
  assign n1335 = ~n1323 & ~n1333;
  assign n1336 = ~n1334 & ~n1335;
  assign n1337 = ~n1318 & n1336;
  assign n1338 = n1318 & ~n1336;
  assign n1339 = ~n1337 & ~n1338;
  assign n1340 = n1317 & n1339;
  assign n1341 = ~n1317 & ~n1339;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = n1252 & ~n1342;
  assign n1344 = ~n1252 & n1342;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = ~n1244 & ~n1249;
  assign n1347 = ~n1345 & n1346;
  assign n1348 = n1345 & ~n1346;
  assign po24  = ~n1347 & ~n1348;
  assign n1350 = ~n1337 & ~n1340;
  assign n1351 = ~n1313 & ~n1315;
  assign n1352 = n1262 & n1273;
  assign n1353 = ~n1262 & ~n1273;
  assign n1354 = ~n1352 & ~n1353;
  assign n1355 = n1306 & ~n1354;
  assign n1356 = ~n1306 & n1354;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = ~n1276 & ~n1282;
  assign n1359 = ~n1181 & ~n1294;
  assign n1360 = ~n1309 & ~n1359;
  assign n1361 = n1358 & n1360;
  assign n1362 = ~n1358 & ~n1360;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = n1357 & n1363;
  assign n1365 = ~n1357 & ~n1363;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~n1351 & n1366;
  assign n1368 = ~n1351 & ~n1367;
  assign n1369 = n1366 & ~n1367;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = pi0  & pi24 ;
  assign n1372 = n1325 & n1371;
  assign n1373 = n1325 & ~n1372;
  assign n1374 = ~n1325 & n1371;
  assign n1375 = ~n1373 & ~n1374;
  assign n1376 = pi1  & pi23 ;
  assign n1377 = pi11  & pi13 ;
  assign n1378 = n1376 & n1377;
  assign n1379 = n1376 & ~n1378;
  assign n1380 = n1377 & ~n1378;
  assign n1381 = ~n1379 & ~n1380;
  assign n1382 = ~n1375 & ~n1381;
  assign n1383 = ~n1375 & ~n1382;
  assign n1384 = ~n1381 & ~n1382;
  assign n1385 = ~n1383 & ~n1384;
  assign n1386 = pi7  & pi17 ;
  assign n1387 = pi18  & pi22 ;
  assign n1388 = n303 & n1387;
  assign n1389 = pi2  & pi22 ;
  assign n1390 = pi6  & pi18 ;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = n1386 & ~n1388;
  assign n1393 = ~n1391 & n1392;
  assign n1394 = n1386 & ~n1393;
  assign n1395 = ~n1388 & ~n1393;
  assign n1396 = ~n1391 & n1395;
  assign n1397 = ~n1394 & ~n1396;
  assign n1398 = ~n1385 & ~n1397;
  assign n1399 = ~n1385 & ~n1398;
  assign n1400 = ~n1397 & ~n1398;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = ~n1329 & ~n1331;
  assign n1403 = n1401 & n1402;
  assign n1404 = ~n1401 & ~n1402;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = pi3  & pi21 ;
  assign n1407 = pi19  & pi20 ;
  assign n1408 = n226 & n1407;
  assign n1409 = pi4  & pi20 ;
  assign n1410 = pi5  & pi19 ;
  assign n1411 = ~n1409 & ~n1410;
  assign n1412 = n1406 & ~n1408;
  assign n1413 = ~n1411 & n1412;
  assign n1414 = n1406 & ~n1413;
  assign n1415 = ~n1408 & ~n1413;
  assign n1416 = ~n1411 & n1415;
  assign n1417 = ~n1414 & ~n1416;
  assign n1418 = n1291 & ~n1417;
  assign n1419 = ~n1291 & n1417;
  assign n1420 = ~n1418 & ~n1419;
  assign n1421 = pi8  & pi16 ;
  assign n1422 = n591 & n1041;
  assign n1423 = pi9  & pi15 ;
  assign n1424 = pi10  & pi14 ;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = n1421 & ~n1422;
  assign n1427 = ~n1425 & n1426;
  assign n1428 = n1421 & ~n1427;
  assign n1429 = ~n1422 & ~n1427;
  assign n1430 = ~n1425 & n1429;
  assign n1431 = ~n1428 & ~n1430;
  assign n1432 = ~n1420 & ~n1431;
  assign n1433 = n1420 & n1431;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = ~n1405 & ~n1434;
  assign n1436 = n1405 & n1434;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = ~n1322 & ~n1334;
  assign n1439 = n1437 & ~n1438;
  assign n1440 = ~n1437 & n1438;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = ~n1370 & n1441;
  assign n1443 = n1370 & ~n1441;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = ~n1350 & n1444;
  assign n1446 = n1350 & ~n1444;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~n1344 & ~n1348;
  assign n1449 = ~n1447 & n1448;
  assign n1450 = ~n1446 & ~n1448;
  assign n1451 = ~n1445 & n1450;
  assign po25  = ~n1449 & ~n1451;
  assign n1453 = ~n1367 & ~n1442;
  assign n1454 = pi0  & pi25 ;
  assign n1455 = pi2  & pi23 ;
  assign n1456 = ~n1454 & ~n1455;
  assign n1457 = pi23  & pi25 ;
  assign n1458 = n196 & n1457;
  assign n1459 = pi10  & pi15 ;
  assign n1460 = ~n1456 & n1459;
  assign n1461 = ~n1458 & n1460;
  assign n1462 = ~n1458 & ~n1461;
  assign n1463 = ~n1456 & n1462;
  assign n1464 = n1459 & ~n1461;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = pi7  & pi18 ;
  assign n1467 = n414 & n989;
  assign n1468 = pi8  & pi17 ;
  assign n1469 = ~n803 & ~n1468;
  assign n1470 = n1466 & ~n1467;
  assign n1471 = ~n1469 & n1470;
  assign n1472 = n1466 & ~n1471;
  assign n1473 = ~n1467 & ~n1471;
  assign n1474 = ~n1469 & n1473;
  assign n1475 = ~n1472 & ~n1474;
  assign n1476 = ~n1465 & ~n1475;
  assign n1477 = ~n1465 & ~n1476;
  assign n1478 = ~n1475 & ~n1476;
  assign n1479 = ~n1477 & ~n1478;
  assign n1480 = pi6  & pi19 ;
  assign n1481 = pi21  & pi22 ;
  assign n1482 = n209 & n1481;
  assign n1483 = pi3  & pi22 ;
  assign n1484 = pi4  & pi21 ;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = n1480 & ~n1482;
  assign n1487 = ~n1485 & n1486;
  assign n1488 = n1480 & ~n1487;
  assign n1489 = ~n1482 & ~n1487;
  assign n1490 = ~n1485 & n1489;
  assign n1491 = ~n1488 & ~n1490;
  assign n1492 = ~n1479 & ~n1491;
  assign n1493 = ~n1479 & ~n1492;
  assign n1494 = ~n1491 & ~n1492;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = ~n1362 & ~n1364;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = ~n1495 & ~n1497;
  assign n1499 = ~n1496 & ~n1497;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = pi1  & pi24 ;
  assign n1502 = pi13  & n1501;
  assign n1503 = ~pi13  & ~n1501;
  assign n1504 = ~n1502 & ~n1503;
  assign n1505 = n1378 & n1504;
  assign n1506 = ~n1378 & ~n1504;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = ~n1415 & n1507;
  assign n1509 = n1415 & ~n1507;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = ~n1353 & ~n1356;
  assign n1512 = pi5  & pi20 ;
  assign n1513 = pi11  & pi14 ;
  assign n1514 = n952 & n1513;
  assign n1515 = ~n952 & ~n1513;
  assign n1516 = n1512 & ~n1514;
  assign n1517 = ~n1515 & n1516;
  assign n1518 = n1512 & ~n1517;
  assign n1519 = ~n1514 & ~n1517;
  assign n1520 = ~n1515 & n1519;
  assign n1521 = ~n1518 & ~n1520;
  assign n1522 = ~n1511 & ~n1521;
  assign n1523 = ~n1511 & ~n1522;
  assign n1524 = ~n1521 & ~n1522;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = n1510 & ~n1525;
  assign n1527 = n1510 & ~n1526;
  assign n1528 = ~n1525 & ~n1526;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = ~n1500 & ~n1529;
  assign n1531 = ~n1500 & ~n1530;
  assign n1532 = ~n1529 & ~n1530;
  assign n1533 = ~n1531 & ~n1532;
  assign n1534 = n1395 & n1429;
  assign n1535 = ~n1395 & ~n1429;
  assign n1536 = ~n1534 & ~n1535;
  assign n1537 = ~n1372 & ~n1382;
  assign n1538 = ~n1536 & n1537;
  assign n1539 = n1536 & ~n1537;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = ~n1291 & ~n1417;
  assign n1542 = ~n1432 & ~n1541;
  assign n1543 = ~n1540 & n1542;
  assign n1544 = n1540 & ~n1542;
  assign n1545 = ~n1543 & ~n1544;
  assign n1546 = ~n1398 & ~n1404;
  assign n1547 = ~n1545 & n1546;
  assign n1548 = n1545 & ~n1546;
  assign n1549 = ~n1547 & ~n1548;
  assign n1550 = ~n1436 & ~n1439;
  assign n1551 = n1549 & ~n1550;
  assign n1552 = n1549 & ~n1551;
  assign n1553 = ~n1550 & ~n1551;
  assign n1554 = ~n1552 & ~n1553;
  assign n1555 = ~n1533 & ~n1554;
  assign n1556 = n1533 & n1554;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = n1453 & ~n1557;
  assign n1559 = ~n1453 & n1557;
  assign n1560 = ~n1558 & ~n1559;
  assign n1561 = ~n1445 & ~n1450;
  assign n1562 = ~n1560 & n1561;
  assign n1563 = n1560 & ~n1561;
  assign po26  = ~n1562 & ~n1563;
  assign n1565 = ~n1551 & ~n1555;
  assign n1566 = pi3  & pi23 ;
  assign n1567 = pi7  & pi19 ;
  assign n1568 = ~n1566 & ~n1567;
  assign n1569 = n1566 & n1567;
  assign n1570 = pi2  & pi24 ;
  assign n1571 = ~n1568 & n1570;
  assign n1572 = ~n1569 & n1571;
  assign n1573 = ~n1569 & ~n1572;
  assign n1574 = ~n1568 & n1573;
  assign n1575 = n1570 & ~n1572;
  assign n1576 = ~n1574 & ~n1575;
  assign n1577 = pi9  & pi17 ;
  assign n1578 = n840 & n1111;
  assign n1579 = pi11  & pi15 ;
  assign n1580 = pi10  & pi16 ;
  assign n1581 = ~n1579 & ~n1580;
  assign n1582 = n1577 & ~n1578;
  assign n1583 = ~n1581 & n1582;
  assign n1584 = n1577 & ~n1583;
  assign n1585 = ~n1578 & ~n1583;
  assign n1586 = ~n1581 & n1585;
  assign n1587 = ~n1584 & ~n1586;
  assign n1588 = ~n1576 & ~n1587;
  assign n1589 = ~n1576 & ~n1588;
  assign n1590 = ~n1587 & ~n1588;
  assign n1591 = ~n1589 & ~n1590;
  assign n1592 = pi4  & pi22 ;
  assign n1593 = pi20  & pi21 ;
  assign n1594 = n326 & n1593;
  assign n1595 = pi5  & pi21 ;
  assign n1596 = pi6  & pi20 ;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = n1592 & ~n1594;
  assign n1599 = ~n1597 & n1598;
  assign n1600 = n1592 & ~n1599;
  assign n1601 = ~n1594 & ~n1599;
  assign n1602 = ~n1597 & n1601;
  assign n1603 = ~n1600 & ~n1602;
  assign n1604 = ~n1591 & ~n1603;
  assign n1605 = ~n1591 & ~n1604;
  assign n1606 = ~n1603 & ~n1604;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = ~n1544 & ~n1548;
  assign n1609 = n1607 & n1608;
  assign n1610 = ~n1607 & ~n1608;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = ~n1535 & ~n1539;
  assign n1613 = ~n1505 & ~n1508;
  assign n1614 = n1612 & n1613;
  assign n1615 = ~n1612 & ~n1613;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = n1462 & n1473;
  assign n1618 = ~n1462 & ~n1473;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = pi0  & pi26 ;
  assign n1621 = pi8  & pi18 ;
  assign n1622 = n1620 & n1621;
  assign n1623 = ~n1620 & ~n1621;
  assign n1624 = n1502 & ~n1622;
  assign n1625 = ~n1623 & n1624;
  assign n1626 = n1502 & ~n1625;
  assign n1627 = ~n1622 & ~n1625;
  assign n1628 = ~n1623 & n1627;
  assign n1629 = ~n1626 & ~n1628;
  assign n1630 = n1619 & ~n1629;
  assign n1631 = n1619 & ~n1630;
  assign n1632 = ~n1629 & ~n1630;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = n1616 & ~n1633;
  assign n1635 = ~n1616 & n1633;
  assign n1636 = ~n1634 & ~n1635;
  assign n1637 = n1611 & n1636;
  assign n1638 = n1611 & ~n1637;
  assign n1639 = n1636 & ~n1637;
  assign n1640 = ~n1638 & ~n1639;
  assign n1641 = ~n1497 & ~n1530;
  assign n1642 = ~n1522 & ~n1526;
  assign n1643 = ~n1476 & ~n1492;
  assign n1644 = pi12  & pi14 ;
  assign n1645 = pi1  & pi25 ;
  assign n1646 = ~n1644 & ~n1645;
  assign n1647 = n1644 & n1645;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = ~n1519 & n1648;
  assign n1650 = ~n1519 & ~n1649;
  assign n1651 = n1648 & ~n1649;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = ~n1489 & ~n1652;
  assign n1654 = n1489 & n1652;
  assign n1655 = ~n1653 & ~n1654;
  assign n1656 = ~n1643 & n1655;
  assign n1657 = n1643 & ~n1655;
  assign n1658 = ~n1656 & ~n1657;
  assign n1659 = ~n1642 & n1658;
  assign n1660 = n1642 & ~n1658;
  assign n1661 = ~n1659 & ~n1660;
  assign n1662 = ~n1641 & n1661;
  assign n1663 = n1641 & ~n1661;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = ~n1640 & ~n1664;
  assign n1666 = n1640 & n1664;
  assign n1667 = ~n1665 & ~n1666;
  assign n1668 = ~n1565 & ~n1667;
  assign n1669 = n1565 & n1667;
  assign n1670 = ~n1668 & ~n1669;
  assign n1671 = ~n1559 & ~n1563;
  assign n1672 = ~n1670 & n1671;
  assign n1673 = n1670 & ~n1671;
  assign po27  = ~n1672 & ~n1673;
  assign n1675 = ~n1610 & ~n1637;
  assign n1676 = pi4  & pi23 ;
  assign n1677 = pi6  & pi21 ;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = n1676 & n1677;
  assign n1680 = pi3  & pi24 ;
  assign n1681 = ~n1678 & n1680;
  assign n1682 = ~n1679 & n1681;
  assign n1683 = ~n1679 & ~n1682;
  assign n1684 = ~n1678 & n1683;
  assign n1685 = n1680 & ~n1682;
  assign n1686 = ~n1684 & ~n1685;
  assign n1687 = pi5  & pi22 ;
  assign n1688 = n952 & n1041;
  assign n1689 = pi12  & pi15 ;
  assign n1690 = ~n706 & ~n1689;
  assign n1691 = n1687 & ~n1688;
  assign n1692 = ~n1690 & n1691;
  assign n1693 = n1687 & ~n1692;
  assign n1694 = ~n1688 & ~n1692;
  assign n1695 = ~n1690 & n1694;
  assign n1696 = ~n1693 & ~n1695;
  assign n1697 = ~n1686 & ~n1696;
  assign n1698 = ~n1686 & ~n1697;
  assign n1699 = ~n1696 & ~n1697;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = pi0  & pi27 ;
  assign n1702 = n1647 & ~n1701;
  assign n1703 = ~n1647 & n1701;
  assign n1704 = ~n1702 & ~n1703;
  assign n1705 = pi26  & n622;
  assign n1706 = pi14  & ~n1705;
  assign n1707 = pi1  & pi26 ;
  assign n1708 = ~n1705 & n1707;
  assign n1709 = ~n1706 & ~n1708;
  assign n1710 = ~n1704 & ~n1709;
  assign n1711 = n1704 & n1709;
  assign n1712 = ~n1710 & ~n1711;
  assign n1713 = n1700 & n1712;
  assign n1714 = ~n1700 & ~n1712;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = n1585 & n1601;
  assign n1717 = ~n1585 & ~n1601;
  assign n1718 = ~n1716 & ~n1717;
  assign n1719 = n1573 & ~n1718;
  assign n1720 = ~n1573 & n1718;
  assign n1721 = ~n1719 & ~n1720;
  assign n1722 = ~n1615 & ~n1634;
  assign n1723 = n1721 & ~n1722;
  assign n1724 = ~n1721 & n1722;
  assign n1725 = ~n1723 & ~n1724;
  assign n1726 = ~n1715 & n1725;
  assign n1727 = n1715 & ~n1725;
  assign n1728 = ~n1726 & ~n1727;
  assign n1729 = ~n1675 & n1728;
  assign n1730 = n1675 & ~n1728;
  assign n1731 = ~n1729 & ~n1730;
  assign n1732 = pi11  & pi16 ;
  assign n1733 = pi20  & pi25 ;
  assign n1734 = n328 & n1733;
  assign n1735 = pi2  & pi25 ;
  assign n1736 = pi7  & pi20 ;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = ~n1734 & ~n1737;
  assign n1739 = ~n1732 & ~n1738;
  assign n1740 = n1732 & n1738;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = ~n1627 & n1741;
  assign n1743 = n1627 & ~n1741;
  assign n1744 = ~n1742 & ~n1743;
  assign n1745 = pi8  & pi19 ;
  assign n1746 = n591 & n1199;
  assign n1747 = pi10  & pi17 ;
  assign n1748 = pi9  & pi18 ;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = n1745 & ~n1746;
  assign n1751 = ~n1749 & n1750;
  assign n1752 = n1745 & ~n1751;
  assign n1753 = ~n1746 & ~n1751;
  assign n1754 = ~n1749 & n1753;
  assign n1755 = ~n1752 & ~n1754;
  assign n1756 = n1744 & ~n1755;
  assign n1757 = n1744 & ~n1756;
  assign n1758 = ~n1755 & ~n1756;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = ~n1656 & ~n1659;
  assign n1761 = n1759 & n1760;
  assign n1762 = ~n1759 & ~n1760;
  assign n1763 = ~n1761 & ~n1762;
  assign n1764 = ~n1649 & ~n1653;
  assign n1765 = ~n1618 & ~n1630;
  assign n1766 = n1764 & n1765;
  assign n1767 = ~n1764 & ~n1765;
  assign n1768 = ~n1766 & ~n1767;
  assign n1769 = ~n1588 & ~n1604;
  assign n1770 = ~n1768 & n1769;
  assign n1771 = n1768 & ~n1769;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = n1763 & n1772;
  assign n1774 = ~n1763 & ~n1772;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = n1731 & n1775;
  assign n1777 = ~n1731 & ~n1775;
  assign n1778 = ~n1776 & ~n1777;
  assign n1779 = ~n1663 & ~n1666;
  assign n1780 = n1778 & n1779;
  assign n1781 = ~n1778 & ~n1779;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = ~n1668 & ~n1673;
  assign n1784 = ~n1782 & n1783;
  assign n1785 = n1782 & ~n1783;
  assign po28  = ~n1784 & ~n1785;
  assign n1787 = ~n1723 & ~n1726;
  assign n1788 = pi8  & pi20 ;
  assign n1789 = pi24  & pi25 ;
  assign n1790 = n209 & n1789;
  assign n1791 = pi3  & pi25 ;
  assign n1792 = pi4  & pi24 ;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = n1788 & ~n1790;
  assign n1795 = ~n1793 & n1794;
  assign n1796 = n1788 & ~n1795;
  assign n1797 = ~n1790 & ~n1795;
  assign n1798 = ~n1793 & n1797;
  assign n1799 = ~n1796 & ~n1798;
  assign n1800 = n1647 & n1701;
  assign n1801 = ~n1710 & ~n1800;
  assign n1802 = ~n1799 & n1801;
  assign n1803 = n1799 & ~n1801;
  assign n1804 = ~n1802 & ~n1803;
  assign n1805 = pi7  & pi21 ;
  assign n1806 = pi22  & pi23 ;
  assign n1807 = n326 & n1806;
  assign n1808 = pi5  & pi23 ;
  assign n1809 = pi6  & pi22 ;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = n1805 & ~n1807;
  assign n1812 = ~n1810 & n1811;
  assign n1813 = n1805 & ~n1812;
  assign n1814 = ~n1807 & ~n1812;
  assign n1815 = ~n1810 & n1814;
  assign n1816 = ~n1813 & ~n1815;
  assign n1817 = ~n1804 & ~n1816;
  assign n1818 = n1804 & n1816;
  assign n1819 = ~n1817 & ~n1818;
  assign n1820 = n1787 & ~n1819;
  assign n1821 = ~n1787 & n1819;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = ~n1700 & n1712;
  assign n1824 = ~n1697 & ~n1823;
  assign n1825 = ~n1742 & ~n1756;
  assign n1826 = pi1  & pi27 ;
  assign n1827 = n777 & n1826;
  assign n1828 = ~n777 & ~n1826;
  assign n1829 = ~n1827 & ~n1828;
  assign n1830 = n1705 & n1829;
  assign n1831 = n1705 & ~n1830;
  assign n1832 = ~n1705 & n1829;
  assign n1833 = ~n1831 & ~n1832;
  assign n1834 = ~n1694 & ~n1833;
  assign n1835 = n1694 & n1833;
  assign n1836 = ~n1834 & ~n1835;
  assign n1837 = ~n1825 & n1836;
  assign n1838 = n1825 & ~n1836;
  assign n1839 = ~n1837 & ~n1838;
  assign n1840 = ~n1824 & n1839;
  assign n1841 = n1824 & ~n1839;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = n1822 & n1842;
  assign n1844 = ~n1822 & ~n1842;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = ~n1729 & ~n1776;
  assign n1847 = ~n1762 & ~n1773;
  assign n1848 = n1683 & n1753;
  assign n1849 = ~n1683 & ~n1753;
  assign n1850 = ~n1848 & ~n1849;
  assign n1851 = ~n1734 & ~n1740;
  assign n1852 = ~n1850 & n1851;
  assign n1853 = n1850 & ~n1851;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = ~n1767 & ~n1771;
  assign n1856 = ~n1854 & n1855;
  assign n1857 = n1854 & ~n1855;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = pi0  & pi28 ;
  assign n1860 = pi12  & pi16 ;
  assign n1861 = ~n1859 & ~n1860;
  assign n1862 = n1859 & n1860;
  assign n1863 = pi11  & pi17 ;
  assign n1864 = ~n1861 & n1863;
  assign n1865 = ~n1862 & n1864;
  assign n1866 = ~n1862 & ~n1865;
  assign n1867 = ~n1861 & n1866;
  assign n1868 = n1863 & ~n1865;
  assign n1869 = ~n1867 & ~n1868;
  assign n1870 = pi2  & pi26 ;
  assign n1871 = n591 & n1085;
  assign n1872 = pi9  & pi19 ;
  assign n1873 = pi10  & pi18 ;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = n1870 & ~n1871;
  assign n1876 = ~n1874 & n1875;
  assign n1877 = n1870 & ~n1876;
  assign n1878 = ~n1871 & ~n1876;
  assign n1879 = ~n1874 & n1878;
  assign n1880 = ~n1877 & ~n1879;
  assign n1881 = ~n1869 & ~n1880;
  assign n1882 = ~n1869 & ~n1881;
  assign n1883 = ~n1880 & ~n1881;
  assign n1884 = ~n1882 & ~n1883;
  assign n1885 = ~n1717 & ~n1720;
  assign n1886 = n1884 & n1885;
  assign n1887 = ~n1884 & ~n1885;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = n1858 & n1888;
  assign n1890 = ~n1858 & ~n1888;
  assign n1891 = ~n1889 & ~n1890;
  assign n1892 = ~n1847 & n1891;
  assign n1893 = n1847 & ~n1891;
  assign n1894 = ~n1892 & ~n1893;
  assign n1895 = ~n1846 & n1894;
  assign n1896 = n1846 & ~n1894;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = ~n1845 & ~n1897;
  assign n1899 = n1845 & n1897;
  assign n1900 = ~n1898 & ~n1899;
  assign n1901 = ~n1780 & ~n1785;
  assign n1902 = ~n1900 & n1901;
  assign n1903 = n1900 & ~n1901;
  assign po29  = ~n1902 & ~n1903;
  assign n1905 = ~n1892 & ~n1895;
  assign n1906 = ~n1857 & ~n1889;
  assign n1907 = ~n1837 & ~n1840;
  assign n1908 = n1906 & n1907;
  assign n1909 = ~n1906 & ~n1907;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = ~n1881 & ~n1887;
  assign n1912 = ~n1799 & ~n1801;
  assign n1913 = ~n1817 & ~n1912;
  assign n1914 = n1911 & n1913;
  assign n1915 = ~n1911 & ~n1913;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = n1866 & n1878;
  assign n1918 = ~n1866 & ~n1878;
  assign n1919 = ~n1917 & ~n1918;
  assign n1920 = pi0  & pi29 ;
  assign n1921 = pi2  & pi27 ;
  assign n1922 = ~n1920 & ~n1921;
  assign n1923 = pi27  & pi29 ;
  assign n1924 = n196 & n1923;
  assign n1925 = n1827 & ~n1922;
  assign n1926 = ~n1924 & n1925;
  assign n1927 = n1827 & ~n1926;
  assign n1928 = ~n1924 & ~n1926;
  assign n1929 = ~n1922 & n1928;
  assign n1930 = ~n1927 & ~n1929;
  assign n1931 = n1919 & ~n1930;
  assign n1932 = n1919 & ~n1931;
  assign n1933 = ~n1930 & ~n1931;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = n1916 & ~n1934;
  assign n1936 = ~n1916 & n1934;
  assign n1937 = ~n1935 & ~n1936;
  assign n1938 = n1910 & n1937;
  assign n1939 = n1910 & ~n1938;
  assign n1940 = n1937 & ~n1938;
  assign n1941 = ~n1939 & ~n1940;
  assign n1942 = ~n1821 & ~n1843;
  assign n1943 = ~n1830 & ~n1834;
  assign n1944 = pi6  & pi23 ;
  assign n1945 = pi13  & pi16 ;
  assign n1946 = n1041 & n1945;
  assign n1947 = ~n1041 & ~n1945;
  assign n1948 = n1944 & ~n1946;
  assign n1949 = ~n1947 & n1948;
  assign n1950 = n1944 & ~n1949;
  assign n1951 = ~n1946 & ~n1949;
  assign n1952 = ~n1947 & n1951;
  assign n1953 = ~n1950 & ~n1952;
  assign n1954 = ~n1943 & ~n1953;
  assign n1955 = ~n1943 & ~n1954;
  assign n1956 = ~n1953 & ~n1954;
  assign n1957 = ~n1955 & ~n1956;
  assign n1958 = ~n1849 & ~n1853;
  assign n1959 = n1957 & n1958;
  assign n1960 = ~n1957 & ~n1958;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = pi3  & pi26 ;
  assign n1963 = pi8  & pi21 ;
  assign n1964 = ~n1962 & ~n1963;
  assign n1965 = pi21  & pi26 ;
  assign n1966 = n417 & n1965;
  assign n1967 = pi12  & pi17 ;
  assign n1968 = ~n1964 & n1967;
  assign n1969 = ~n1966 & n1968;
  assign n1970 = ~n1966 & ~n1969;
  assign n1971 = ~n1964 & n1970;
  assign n1972 = n1967 & ~n1969;
  assign n1973 = ~n1971 & ~n1972;
  assign n1974 = pi9  & pi20 ;
  assign n1975 = n1085 & n1111;
  assign n1976 = pi10  & pi19 ;
  assign n1977 = pi11  & pi18 ;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = n1974 & ~n1975;
  assign n1980 = ~n1978 & n1979;
  assign n1981 = n1974 & ~n1980;
  assign n1982 = ~n1975 & ~n1980;
  assign n1983 = ~n1978 & n1982;
  assign n1984 = ~n1981 & ~n1983;
  assign n1985 = ~n1973 & ~n1984;
  assign n1986 = ~n1973 & ~n1985;
  assign n1987 = ~n1984 & ~n1985;
  assign n1988 = ~n1986 & ~n1987;
  assign n1989 = pi4  & pi25 ;
  assign n1990 = pi22  & pi24 ;
  assign n1991 = n481 & n1990;
  assign n1992 = pi7  & pi22 ;
  assign n1993 = pi5  & pi24 ;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = n1989 & ~n1991;
  assign n1996 = ~n1994 & n1995;
  assign n1997 = n1989 & ~n1996;
  assign n1998 = ~n1991 & ~n1996;
  assign n1999 = ~n1994 & n1998;
  assign n2000 = ~n1997 & ~n1999;
  assign n2001 = ~n1988 & ~n2000;
  assign n2002 = ~n1988 & ~n2001;
  assign n2003 = ~n2000 & ~n2001;
  assign n2004 = ~n2002 & ~n2003;
  assign n2005 = pi28  & n723;
  assign n2006 = pi1  & pi28 ;
  assign n2007 = ~pi15  & ~n2006;
  assign n2008 = ~n2005 & ~n2007;
  assign n2009 = n1814 & ~n2008;
  assign n2010 = ~n1814 & n2008;
  assign n2011 = ~n2009 & ~n2010;
  assign n2012 = ~n1797 & n2011;
  assign n2013 = n1797 & ~n2011;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = ~n2004 & n2014;
  assign n2016 = n2004 & ~n2014;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = n1961 & n2017;
  assign n2019 = ~n1961 & ~n2017;
  assign n2020 = ~n2018 & ~n2019;
  assign n2021 = ~n1942 & n2020;
  assign n2022 = ~n1942 & ~n2021;
  assign n2023 = n2020 & ~n2021;
  assign n2024 = ~n2022 & ~n2023;
  assign n2025 = ~n1941 & ~n2024;
  assign n2026 = n1941 & n2024;
  assign n2027 = ~n2025 & ~n2026;
  assign n2028 = ~n1905 & n2027;
  assign n2029 = n1905 & ~n2027;
  assign n2030 = ~n2028 & ~n2029;
  assign n2031 = ~n1899 & ~n1903;
  assign n2032 = ~n2030 & n2031;
  assign n2033 = n2030 & ~n2031;
  assign po30  = ~n2032 & ~n2033;
  assign n2035 = ~n2021 & ~n2025;
  assign n2036 = pi0  & pi30 ;
  assign n2037 = n2005 & n2036;
  assign n2038 = n2005 & ~n2037;
  assign n2039 = ~n2005 & n2036;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = pi1  & pi29 ;
  assign n2042 = pi14  & pi16 ;
  assign n2043 = n2041 & n2042;
  assign n2044 = n2041 & ~n2043;
  assign n2045 = n2042 & ~n2043;
  assign n2046 = ~n2044 & ~n2045;
  assign n2047 = ~n2040 & ~n2046;
  assign n2048 = ~n2040 & ~n2047;
  assign n2049 = ~n2046 & ~n2047;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = ~n2010 & ~n2012;
  assign n2052 = n2050 & n2051;
  assign n2053 = ~n2050 & ~n2051;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = ~n1918 & ~n1931;
  assign n2056 = ~n2054 & n2055;
  assign n2057 = n2054 & ~n2055;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = ~n2015 & ~n2018;
  assign n2060 = ~n2058 & n2059;
  assign n2061 = n2058 & ~n2059;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = n1951 & n1998;
  assign n2064 = ~n1951 & ~n1998;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = pi13  & pi17 ;
  assign n2067 = pi2  & pi28 ;
  assign n2068 = pi9  & pi21 ;
  assign n2069 = n2067 & n2068;
  assign n2070 = ~n2067 & ~n2068;
  assign n2071 = n2066 & ~n2069;
  assign n2072 = ~n2070 & n2071;
  assign n2073 = n2066 & ~n2072;
  assign n2074 = ~n2069 & ~n2072;
  assign n2075 = ~n2070 & n2074;
  assign n2076 = ~n2073 & ~n2075;
  assign n2077 = n2065 & ~n2076;
  assign n2078 = n2065 & ~n2077;
  assign n2079 = ~n2076 & ~n2077;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = ~n1985 & ~n2001;
  assign n2082 = n2080 & n2081;
  assign n2083 = ~n2080 & ~n2081;
  assign n2084 = ~n2082 & ~n2083;
  assign n2085 = n1970 & n1982;
  assign n2086 = ~n1970 & ~n1982;
  assign n2087 = ~n2085 & ~n2086;
  assign n2088 = n1928 & ~n2087;
  assign n2089 = ~n1928 & n2087;
  assign n2090 = ~n2088 & ~n2089;
  assign n2091 = n2084 & n2090;
  assign n2092 = ~n2084 & ~n2090;
  assign n2093 = ~n2091 & ~n2092;
  assign n2094 = n2062 & n2093;
  assign n2095 = ~n2062 & ~n2093;
  assign n2096 = ~n2094 & ~n2095;
  assign n2097 = ~n1909 & ~n1938;
  assign n2098 = pi4  & pi26 ;
  assign n2099 = pi8  & pi22 ;
  assign n2100 = ~n2098 & ~n2099;
  assign n2101 = n2098 & n2099;
  assign n2102 = pi3  & pi27 ;
  assign n2103 = ~n2100 & n2102;
  assign n2104 = ~n2101 & n2103;
  assign n2105 = ~n2101 & ~n2104;
  assign n2106 = ~n2100 & n2105;
  assign n2107 = n2102 & ~n2104;
  assign n2108 = ~n2106 & ~n2107;
  assign n2109 = pi5  & pi25 ;
  assign n2110 = pi23  & pi24 ;
  assign n2111 = n432 & n2110;
  assign n2112 = pi6  & pi24 ;
  assign n2113 = pi7  & pi23 ;
  assign n2114 = ~n2112 & ~n2113;
  assign n2115 = n2109 & ~n2111;
  assign n2116 = ~n2114 & n2115;
  assign n2117 = n2109 & ~n2116;
  assign n2118 = ~n2111 & ~n2116;
  assign n2119 = ~n2114 & n2118;
  assign n2120 = ~n2117 & ~n2119;
  assign n2121 = ~n2108 & ~n2120;
  assign n2122 = ~n2108 & ~n2121;
  assign n2123 = ~n2120 & ~n2121;
  assign n2124 = ~n2122 & ~n2123;
  assign n2125 = pi10  & pi20 ;
  assign n2126 = n579 & n1085;
  assign n2127 = pi11  & pi19 ;
  assign n2128 = pi12  & pi18 ;
  assign n2129 = ~n2127 & ~n2128;
  assign n2130 = n2125 & ~n2126;
  assign n2131 = ~n2129 & n2130;
  assign n2132 = n2125 & ~n2131;
  assign n2133 = ~n2126 & ~n2131;
  assign n2134 = ~n2129 & n2133;
  assign n2135 = ~n2132 & ~n2134;
  assign n2136 = ~n2124 & ~n2135;
  assign n2137 = ~n2124 & ~n2136;
  assign n2138 = ~n2135 & ~n2136;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140 = ~n1954 & ~n1960;
  assign n2141 = n2139 & n2140;
  assign n2142 = ~n2139 & ~n2140;
  assign n2143 = ~n2141 & ~n2142;
  assign n2144 = ~n1915 & ~n1935;
  assign n2145 = n2143 & ~n2144;
  assign n2146 = ~n2143 & n2144;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = ~n2097 & n2147;
  assign n2149 = n2097 & ~n2147;
  assign n2150 = ~n2148 & ~n2149;
  assign n2151 = n2096 & n2150;
  assign n2152 = ~n2096 & ~n2150;
  assign n2153 = ~n2151 & ~n2152;
  assign n2154 = ~n2035 & n2153;
  assign n2155 = n2035 & ~n2153;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = ~n2028 & ~n2033;
  assign n2158 = ~n2156 & n2157;
  assign n2159 = n2156 & ~n2157;
  assign po31  = ~n2158 & ~n2159;
  assign n2161 = ~n2148 & ~n2151;
  assign n2162 = ~n2061 & ~n2094;
  assign n2163 = ~n2083 & ~n2091;
  assign n2164 = pi5  & pi26 ;
  assign n2165 = pi7  & pi24 ;
  assign n2166 = ~n2164 & ~n2165;
  assign n2167 = pi24  & pi26 ;
  assign n2168 = n481 & n2167;
  assign n2169 = pi8  & pi23 ;
  assign n2170 = ~n2166 & n2169;
  assign n2171 = ~n2168 & n2170;
  assign n2172 = ~n2168 & ~n2171;
  assign n2173 = ~n2166 & n2172;
  assign n2174 = n2169 & ~n2171;
  assign n2175 = ~n2173 & ~n2174;
  assign n2176 = pi6  & pi25 ;
  assign n2177 = n989 & n1041;
  assign n2178 = pi14  & pi17 ;
  assign n2179 = ~n840 & ~n2178;
  assign n2180 = n2176 & ~n2177;
  assign n2181 = ~n2179 & n2180;
  assign n2182 = n2176 & ~n2181;
  assign n2183 = ~n2177 & ~n2181;
  assign n2184 = ~n2179 & n2183;
  assign n2185 = ~n2182 & ~n2184;
  assign n2186 = ~n2175 & ~n2185;
  assign n2187 = ~n2175 & ~n2186;
  assign n2188 = ~n2185 & ~n2186;
  assign n2189 = ~n2187 & ~n2188;
  assign n2190 = pi2  & pi29 ;
  assign n2191 = pi27  & pi28 ;
  assign n2192 = n209 & n2191;
  assign n2193 = pi3  & pi28 ;
  assign n2194 = pi4  & pi27 ;
  assign n2195 = ~n2193 & ~n2194;
  assign n2196 = n2190 & ~n2192;
  assign n2197 = ~n2195 & n2196;
  assign n2198 = n2190 & ~n2197;
  assign n2199 = ~n2192 & ~n2197;
  assign n2200 = ~n2195 & n2199;
  assign n2201 = ~n2198 & ~n2200;
  assign n2202 = ~n2189 & ~n2201;
  assign n2203 = ~n2189 & ~n2202;
  assign n2204 = ~n2201 & ~n2202;
  assign n2205 = ~n2203 & ~n2204;
  assign n2206 = pi0  & pi31 ;
  assign n2207 = pi9  & pi22 ;
  assign n2208 = ~n2206 & ~n2207;
  assign n2209 = pi22  & pi31 ;
  assign n2210 = n339 & n2209;
  assign n2211 = pi10  & pi21 ;
  assign n2212 = ~n2208 & n2211;
  assign n2213 = ~n2210 & n2212;
  assign n2214 = ~n2210 & ~n2213;
  assign n2215 = ~n2208 & n2214;
  assign n2216 = n2211 & ~n2213;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = ~n2037 & ~n2047;
  assign n2219 = pi11  & pi20 ;
  assign n2220 = n952 & n1085;
  assign n2221 = pi12  & pi19 ;
  assign n2222 = pi13  & pi18 ;
  assign n2223 = ~n2221 & ~n2222;
  assign n2224 = n2219 & ~n2220;
  assign n2225 = ~n2223 & n2224;
  assign n2226 = n2219 & ~n2225;
  assign n2227 = ~n2220 & ~n2225;
  assign n2228 = ~n2223 & n2227;
  assign n2229 = ~n2226 & ~n2228;
  assign n2230 = ~n2218 & ~n2229;
  assign n2231 = ~n2218 & ~n2230;
  assign n2232 = ~n2229 & ~n2230;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = ~n2217 & ~n2233;
  assign n2235 = n2217 & n2233;
  assign n2236 = ~n2234 & ~n2235;
  assign n2237 = ~n2205 & n2236;
  assign n2238 = n2205 & ~n2236;
  assign n2239 = ~n2237 & ~n2238;
  assign n2240 = ~n2163 & n2239;
  assign n2241 = n2163 & ~n2239;
  assign n2242 = ~n2240 & ~n2241;
  assign n2243 = ~n2162 & n2242;
  assign n2244 = n2162 & ~n2242;
  assign n2245 = ~n2243 & ~n2244;
  assign n2246 = ~n2142 & ~n2145;
  assign n2247 = ~n2064 & ~n2077;
  assign n2248 = ~n2086 & ~n2089;
  assign n2249 = n2247 & n2248;
  assign n2250 = ~n2247 & ~n2248;
  assign n2251 = ~n2249 & ~n2250;
  assign n2252 = pi1  & pi30 ;
  assign n2253 = pi16  & n2252;
  assign n2254 = ~pi16  & ~n2252;
  assign n2255 = ~n2253 & ~n2254;
  assign n2256 = n2043 & n2255;
  assign n2257 = ~n2043 & ~n2255;
  assign n2258 = ~n2256 & ~n2257;
  assign n2259 = ~n2118 & n2258;
  assign n2260 = n2118 & ~n2258;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = n2251 & n2261;
  assign n2263 = ~n2251 & ~n2261;
  assign n2264 = ~n2262 & ~n2263;
  assign n2265 = n2246 & ~n2264;
  assign n2266 = ~n2246 & n2264;
  assign n2267 = ~n2265 & ~n2266;
  assign n2268 = n2074 & n2105;
  assign n2269 = ~n2074 & ~n2105;
  assign n2270 = ~n2268 & ~n2269;
  assign n2271 = n2133 & ~n2270;
  assign n2272 = ~n2133 & n2270;
  assign n2273 = ~n2271 & ~n2272;
  assign n2274 = ~n2121 & ~n2136;
  assign n2275 = ~n2273 & n2274;
  assign n2276 = n2273 & ~n2274;
  assign n2277 = ~n2275 & ~n2276;
  assign n2278 = ~n2053 & ~n2057;
  assign n2279 = ~n2277 & n2278;
  assign n2280 = n2277 & ~n2278;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = n2267 & n2281;
  assign n2283 = ~n2267 & ~n2281;
  assign n2284 = ~n2282 & ~n2283;
  assign n2285 = n2245 & n2284;
  assign n2286 = ~n2245 & ~n2284;
  assign n2287 = ~n2285 & ~n2286;
  assign n2288 = ~n2161 & n2287;
  assign n2289 = n2161 & ~n2287;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = ~n2154 & ~n2159;
  assign n2292 = ~n2290 & n2291;
  assign n2293 = n2290 & ~n2291;
  assign po32  = ~n2292 & ~n2293;
  assign n2295 = ~n2243 & ~n2285;
  assign n2296 = ~n2266 & ~n2282;
  assign n2297 = ~n2276 & ~n2280;
  assign n2298 = pi5  & pi27 ;
  assign n2299 = pi4  & pi28 ;
  assign n2300 = ~n2298 & ~n2299;
  assign n2301 = n226 & n2191;
  assign n2302 = pi9  & pi23 ;
  assign n2303 = ~n2300 & n2302;
  assign n2304 = ~n2301 & n2303;
  assign n2305 = ~n2301 & ~n2304;
  assign n2306 = ~n2300 & n2305;
  assign n2307 = n2302 & ~n2304;
  assign n2308 = ~n2306 & ~n2307;
  assign n2309 = pi8  & pi24 ;
  assign n2310 = pi25  & pi26 ;
  assign n2311 = n432 & n2310;
  assign n2312 = pi6  & pi26 ;
  assign n2313 = pi7  & pi25 ;
  assign n2314 = ~n2312 & ~n2313;
  assign n2315 = n2309 & ~n2311;
  assign n2316 = ~n2314 & n2315;
  assign n2317 = n2309 & ~n2316;
  assign n2318 = ~n2311 & ~n2316;
  assign n2319 = ~n2314 & n2318;
  assign n2320 = ~n2317 & ~n2319;
  assign n2321 = ~n2308 & ~n2320;
  assign n2322 = ~n2308 & ~n2321;
  assign n2323 = ~n2320 & ~n2321;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = ~n2256 & ~n2259;
  assign n2326 = n2324 & n2325;
  assign n2327 = ~n2324 & ~n2325;
  assign n2328 = ~n2326 & ~n2327;
  assign n2329 = pi0  & pi32 ;
  assign n2330 = pi2  & pi30 ;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = pi30  & pi32 ;
  assign n2333 = n196 & n2332;
  assign n2334 = n2253 & ~n2331;
  assign n2335 = ~n2333 & n2334;
  assign n2336 = ~n2333 & ~n2335;
  assign n2337 = ~n2331 & n2336;
  assign n2338 = n2253 & ~n2335;
  assign n2339 = ~n2337 & ~n2338;
  assign n2340 = pi11  & pi21 ;
  assign n2341 = n952 & n1407;
  assign n2342 = pi12  & pi20 ;
  assign n2343 = pi13  & pi19 ;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = n2340 & ~n2341;
  assign n2346 = ~n2344 & n2345;
  assign n2347 = n2340 & ~n2346;
  assign n2348 = ~n2341 & ~n2346;
  assign n2349 = ~n2344 & n2348;
  assign n2350 = ~n2347 & ~n2349;
  assign n2351 = ~n2339 & ~n2350;
  assign n2352 = ~n2339 & ~n2351;
  assign n2353 = ~n2350 & ~n2351;
  assign n2354 = ~n2352 & ~n2353;
  assign n2355 = pi14  & pi18 ;
  assign n2356 = pi3  & pi29 ;
  assign n2357 = pi10  & pi22 ;
  assign n2358 = n2356 & n2357;
  assign n2359 = ~n2356 & ~n2357;
  assign n2360 = n2355 & ~n2358;
  assign n2361 = ~n2359 & n2360;
  assign n2362 = n2355 & ~n2361;
  assign n2363 = ~n2358 & ~n2361;
  assign n2364 = ~n2359 & n2363;
  assign n2365 = ~n2362 & ~n2364;
  assign n2366 = ~n2354 & ~n2365;
  assign n2367 = ~n2354 & ~n2366;
  assign n2368 = ~n2365 & ~n2366;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = ~n2328 & n2369;
  assign n2371 = n2328 & ~n2369;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = ~n2297 & n2372;
  assign n2374 = n2297 & ~n2372;
  assign n2375 = ~n2373 & ~n2374;
  assign n2376 = ~n2296 & n2375;
  assign n2377 = n2296 & ~n2375;
  assign n2378 = ~n2376 & ~n2377;
  assign n2379 = ~n2250 & ~n2262;
  assign n2380 = n2214 & n2227;
  assign n2381 = ~n2214 & ~n2227;
  assign n2382 = ~n2380 & ~n2381;
  assign n2383 = n2199 & ~n2382;
  assign n2384 = ~n2199 & n2382;
  assign n2385 = ~n2383 & ~n2384;
  assign n2386 = pi1  & pi31 ;
  assign n2387 = ~n942 & ~n2386;
  assign n2388 = n942 & n2386;
  assign n2389 = ~n2387 & ~n2388;
  assign n2390 = n2183 & ~n2389;
  assign n2391 = ~n2183 & n2389;
  assign n2392 = ~n2390 & ~n2391;
  assign n2393 = ~n2172 & n2392;
  assign n2394 = n2172 & ~n2392;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = n2385 & n2395;
  assign n2397 = ~n2385 & ~n2395;
  assign n2398 = ~n2396 & ~n2397;
  assign n2399 = n2379 & ~n2398;
  assign n2400 = ~n2379 & n2398;
  assign n2401 = ~n2399 & ~n2400;
  assign n2402 = ~n2230 & ~n2234;
  assign n2403 = ~n2269 & ~n2272;
  assign n2404 = n2402 & n2403;
  assign n2405 = ~n2402 & ~n2403;
  assign n2406 = ~n2404 & ~n2405;
  assign n2407 = ~n2186 & ~n2202;
  assign n2408 = ~n2406 & n2407;
  assign n2409 = n2406 & ~n2407;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = ~n2237 & ~n2240;
  assign n2412 = ~n2410 & n2411;
  assign n2413 = n2410 & ~n2411;
  assign n2414 = ~n2412 & ~n2413;
  assign n2415 = n2401 & n2414;
  assign n2416 = ~n2401 & ~n2414;
  assign n2417 = ~n2415 & ~n2416;
  assign n2418 = n2378 & n2417;
  assign n2419 = ~n2378 & ~n2417;
  assign n2420 = ~n2418 & ~n2419;
  assign n2421 = ~n2295 & n2420;
  assign n2422 = n2295 & ~n2420;
  assign n2423 = ~n2421 & ~n2422;
  assign n2424 = ~n2288 & ~n2293;
  assign n2425 = n2423 & ~n2424;
  assign n2426 = ~n2423 & n2424;
  assign po33  = ~n2425 & ~n2426;
  assign n2428 = n2336 & n2348;
  assign n2429 = ~n2336 & ~n2348;
  assign n2430 = ~n2428 & ~n2429;
  assign n2431 = n2363 & ~n2430;
  assign n2432 = ~n2363 & n2430;
  assign n2433 = ~n2431 & ~n2432;
  assign n2434 = n2305 & n2318;
  assign n2435 = ~n2305 & ~n2318;
  assign n2436 = ~n2434 & ~n2435;
  assign n2437 = pi2  & pi31 ;
  assign n2438 = pi22  & pi33 ;
  assign n2439 = n434 & n2438;
  assign n2440 = pi0  & pi33 ;
  assign n2441 = pi11  & pi22 ;
  assign n2442 = ~n2440 & ~n2441;
  assign n2443 = n2437 & ~n2439;
  assign n2444 = ~n2442 & n2443;
  assign n2445 = n2437 & ~n2444;
  assign n2446 = ~n2439 & ~n2444;
  assign n2447 = ~n2442 & n2446;
  assign n2448 = ~n2445 & ~n2447;
  assign n2449 = n2436 & ~n2448;
  assign n2450 = n2436 & ~n2449;
  assign n2451 = ~n2448 & ~n2449;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = ~n2433 & n2452;
  assign n2454 = n2433 & ~n2452;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = pi4  & pi29 ;
  assign n2457 = pi9  & pi24 ;
  assign n2458 = ~n2456 & ~n2457;
  assign n2459 = n2456 & n2457;
  assign n2460 = pi3  & pi30 ;
  assign n2461 = ~n2458 & n2460;
  assign n2462 = ~n2459 & n2461;
  assign n2463 = ~n2459 & ~n2462;
  assign n2464 = ~n2458 & n2463;
  assign n2465 = n2460 & ~n2462;
  assign n2466 = ~n2464 & ~n2465;
  assign n2467 = pi5  & pi28 ;
  assign n2468 = pi25  & pi27 ;
  assign n2469 = n305 & n2468;
  assign n2470 = pi8  & pi25 ;
  assign n2471 = pi6  & pi27 ;
  assign n2472 = ~n2470 & ~n2471;
  assign n2473 = n2467 & ~n2469;
  assign n2474 = ~n2472 & n2473;
  assign n2475 = n2467 & ~n2474;
  assign n2476 = ~n2469 & ~n2474;
  assign n2477 = ~n2472 & n2476;
  assign n2478 = ~n2475 & ~n2477;
  assign n2479 = ~n2466 & ~n2478;
  assign n2480 = ~n2466 & ~n2479;
  assign n2481 = ~n2478 & ~n2479;
  assign n2482 = ~n2480 & ~n2481;
  assign n2483 = pi7  & pi26 ;
  assign n2484 = n840 & n1199;
  assign n2485 = pi15  & pi18 ;
  assign n2486 = ~n989 & ~n2485;
  assign n2487 = n2483 & ~n2484;
  assign n2488 = ~n2486 & n2487;
  assign n2489 = n2483 & ~n2488;
  assign n2490 = ~n2484 & ~n2488;
  assign n2491 = ~n2486 & n2490;
  assign n2492 = ~n2489 & ~n2491;
  assign n2493 = ~n2482 & ~n2492;
  assign n2494 = ~n2482 & ~n2493;
  assign n2495 = ~n2492 & ~n2493;
  assign n2496 = ~n2494 & ~n2495;
  assign n2497 = n2455 & n2496;
  assign n2498 = ~n2455 & ~n2496;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = ~n2381 & ~n2384;
  assign n2501 = ~n2351 & ~n2366;
  assign n2502 = n2500 & n2501;
  assign n2503 = ~n2500 & ~n2501;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = ~n2321 & ~n2327;
  assign n2506 = ~n2504 & n2505;
  assign n2507 = n2504 & ~n2505;
  assign n2508 = ~n2506 & ~n2507;
  assign n2509 = ~n2371 & ~n2373;
  assign n2510 = n2508 & ~n2509;
  assign n2511 = ~n2508 & n2509;
  assign n2512 = ~n2510 & ~n2511;
  assign n2513 = ~n2499 & n2512;
  assign n2514 = n2499 & ~n2512;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = pi10  & pi23 ;
  assign n2517 = ~n2388 & ~n2516;
  assign n2518 = n2388 & n2516;
  assign n2519 = pi1  & pi32 ;
  assign n2520 = pi17  & ~n2519;
  assign n2521 = ~pi17  & n2519;
  assign n2522 = ~n2520 & ~n2521;
  assign n2523 = ~n2517 & ~n2518;
  assign n2524 = ~n2522 & n2523;
  assign n2525 = ~n2518 & ~n2524;
  assign n2526 = ~n2517 & n2525;
  assign n2527 = ~n2522 & ~n2524;
  assign n2528 = ~n2526 & ~n2527;
  assign n2529 = pi12  & pi21 ;
  assign n2530 = n706 & n1407;
  assign n2531 = pi13  & pi20 ;
  assign n2532 = pi14  & pi19 ;
  assign n2533 = ~n2531 & ~n2532;
  assign n2534 = n2529 & ~n2530;
  assign n2535 = ~n2533 & n2534;
  assign n2536 = n2529 & ~n2535;
  assign n2537 = ~n2530 & ~n2535;
  assign n2538 = ~n2533 & n2537;
  assign n2539 = ~n2536 & ~n2538;
  assign n2540 = ~n2528 & ~n2539;
  assign n2541 = ~n2528 & ~n2540;
  assign n2542 = ~n2539 & ~n2540;
  assign n2543 = ~n2541 & ~n2542;
  assign n2544 = ~n2391 & ~n2393;
  assign n2545 = n2543 & n2544;
  assign n2546 = ~n2543 & ~n2544;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = ~n2405 & ~n2409;
  assign n2549 = ~n2547 & n2548;
  assign n2550 = n2547 & ~n2548;
  assign n2551 = ~n2549 & ~n2550;
  assign n2552 = ~n2396 & ~n2400;
  assign n2553 = ~n2551 & n2552;
  assign n2554 = n2551 & ~n2552;
  assign n2555 = ~n2553 & ~n2554;
  assign n2556 = ~n2413 & ~n2415;
  assign n2557 = n2555 & ~n2556;
  assign n2558 = ~n2555 & n2556;
  assign n2559 = ~n2557 & ~n2558;
  assign n2560 = n2515 & n2559;
  assign n2561 = ~n2515 & ~n2559;
  assign n2562 = ~n2560 & ~n2561;
  assign n2563 = ~n2376 & ~n2418;
  assign n2564 = ~n2562 & n2563;
  assign n2565 = n2562 & ~n2563;
  assign n2566 = ~n2564 & ~n2565;
  assign n2567 = ~n2421 & ~n2425;
  assign n2568 = ~n2566 & n2567;
  assign n2569 = n2566 & ~n2567;
  assign po34  = ~n2568 & ~n2569;
  assign n2571 = ~n2557 & ~n2560;
  assign n2572 = n2446 & n2463;
  assign n2573 = ~n2446 & ~n2463;
  assign n2574 = ~n2572 & ~n2573;
  assign n2575 = n2476 & ~n2574;
  assign n2576 = ~n2476 & n2574;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = ~n2479 & ~n2493;
  assign n2579 = pi17  & n2519;
  assign n2580 = pi16  & pi18 ;
  assign n2581 = pi1  & pi33 ;
  assign n2582 = n2580 & n2581;
  assign n2583 = ~n2580 & ~n2581;
  assign n2584 = ~n2582 & ~n2583;
  assign n2585 = n2579 & n2584;
  assign n2586 = ~n2579 & ~n2584;
  assign n2587 = ~n2585 & ~n2586;
  assign n2588 = ~n2490 & n2587;
  assign n2589 = n2490 & ~n2587;
  assign n2590 = ~n2588 & ~n2589;
  assign n2591 = ~n2578 & n2590;
  assign n2592 = n2578 & ~n2590;
  assign n2593 = ~n2591 & ~n2592;
  assign n2594 = n2577 & n2593;
  assign n2595 = ~n2577 & ~n2593;
  assign n2596 = ~n2594 & ~n2595;
  assign n2597 = n2525 & n2537;
  assign n2598 = ~n2525 & ~n2537;
  assign n2599 = ~n2597 & ~n2598;
  assign n2600 = pi2  & pi32 ;
  assign n2601 = n579 & n1806;
  assign n2602 = pi11  & pi23 ;
  assign n2603 = pi12  & pi22 ;
  assign n2604 = ~n2602 & ~n2603;
  assign n2605 = n2600 & ~n2601;
  assign n2606 = ~n2604 & n2605;
  assign n2607 = n2600 & ~n2606;
  assign n2608 = ~n2601 & ~n2606;
  assign n2609 = ~n2604 & n2608;
  assign n2610 = ~n2607 & ~n2609;
  assign n2611 = n2599 & ~n2610;
  assign n2612 = n2599 & ~n2611;
  assign n2613 = ~n2610 & ~n2611;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = ~n2540 & ~n2546;
  assign n2616 = n2614 & n2615;
  assign n2617 = ~n2614 & ~n2615;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = pi5  & pi29 ;
  assign n2620 = pi9  & pi25 ;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = n2619 & n2620;
  assign n2623 = pi10  & pi24 ;
  assign n2624 = ~n2621 & n2623;
  assign n2625 = ~n2622 & n2624;
  assign n2626 = ~n2622 & ~n2625;
  assign n2627 = ~n2621 & n2626;
  assign n2628 = n2623 & ~n2625;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = pi13  & pi21 ;
  assign n2631 = n1041 & n1407;
  assign n2632 = pi14  & pi20 ;
  assign n2633 = pi15  & pi19 ;
  assign n2634 = ~n2632 & ~n2633;
  assign n2635 = n2630 & ~n2631;
  assign n2636 = ~n2634 & n2635;
  assign n2637 = n2630 & ~n2636;
  assign n2638 = ~n2631 & ~n2636;
  assign n2639 = ~n2634 & n2638;
  assign n2640 = ~n2637 & ~n2639;
  assign n2641 = ~n2629 & ~n2640;
  assign n2642 = ~n2629 & ~n2641;
  assign n2643 = ~n2640 & ~n2641;
  assign n2644 = ~n2642 & ~n2643;
  assign n2645 = pi6  & pi28 ;
  assign n2646 = pi26  & pi27 ;
  assign n2647 = n521 & n2646;
  assign n2648 = pi7  & pi27 ;
  assign n2649 = pi8  & pi26 ;
  assign n2650 = ~n2648 & ~n2649;
  assign n2651 = n2645 & ~n2647;
  assign n2652 = ~n2650 & n2651;
  assign n2653 = n2645 & ~n2652;
  assign n2654 = ~n2647 & ~n2652;
  assign n2655 = ~n2650 & n2654;
  assign n2656 = ~n2653 & ~n2655;
  assign n2657 = ~n2644 & ~n2656;
  assign n2658 = ~n2644 & ~n2657;
  assign n2659 = ~n2656 & ~n2657;
  assign n2660 = ~n2658 & ~n2659;
  assign n2661 = n2618 & ~n2660;
  assign n2662 = ~n2618 & n2660;
  assign n2663 = ~n2661 & ~n2662;
  assign n2664 = n2596 & n2663;
  assign n2665 = n2596 & ~n2664;
  assign n2666 = n2663 & ~n2664;
  assign n2667 = ~n2665 & ~n2666;
  assign n2668 = ~n2550 & ~n2554;
  assign n2669 = n2667 & n2668;
  assign n2670 = ~n2667 & ~n2668;
  assign n2671 = ~n2669 & ~n2670;
  assign n2672 = ~n2510 & ~n2513;
  assign n2673 = ~n2503 & ~n2507;
  assign n2674 = ~n2453 & ~n2497;
  assign n2675 = n2673 & ~n2674;
  assign n2676 = ~n2673 & n2674;
  assign n2677 = ~n2675 & ~n2676;
  assign n2678 = ~n2435 & ~n2449;
  assign n2679 = ~n2429 & ~n2432;
  assign n2680 = pi30  & pi31 ;
  assign n2681 = n209 & n2680;
  assign n2682 = pi3  & pi31 ;
  assign n2683 = pi4  & pi30 ;
  assign n2684 = ~n2682 & ~n2683;
  assign n2685 = ~n2681 & ~n2684;
  assign n2686 = pi0  & pi34 ;
  assign n2687 = ~n2685 & ~n2686;
  assign n2688 = n2685 & n2686;
  assign n2689 = ~n2687 & ~n2688;
  assign n2690 = ~n2679 & n2689;
  assign n2691 = n2679 & ~n2689;
  assign n2692 = ~n2690 & ~n2691;
  assign n2693 = ~n2678 & n2692;
  assign n2694 = n2678 & ~n2692;
  assign n2695 = ~n2693 & ~n2694;
  assign n2696 = n2677 & n2695;
  assign n2697 = ~n2677 & ~n2695;
  assign n2698 = ~n2696 & ~n2697;
  assign n2699 = n2672 & ~n2698;
  assign n2700 = ~n2672 & n2698;
  assign n2701 = ~n2699 & ~n2700;
  assign n2702 = n2671 & n2701;
  assign n2703 = ~n2671 & ~n2701;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = ~n2571 & n2704;
  assign n2706 = n2571 & ~n2704;
  assign n2707 = ~n2705 & ~n2706;
  assign n2708 = ~n2565 & ~n2569;
  assign n2709 = ~n2707 & n2708;
  assign n2710 = ~n2706 & ~n2708;
  assign n2711 = ~n2705 & n2710;
  assign po35  = ~n2709 & ~n2711;
  assign n2713 = ~n2705 & ~n2710;
  assign n2714 = ~n2700 & ~n2702;
  assign n2715 = ~n2664 & ~n2670;
  assign n2716 = ~n2573 & ~n2576;
  assign n2717 = ~n2585 & ~n2588;
  assign n2718 = n2716 & n2717;
  assign n2719 = ~n2716 & ~n2717;
  assign n2720 = ~n2718 & ~n2719;
  assign n2721 = ~n2598 & ~n2611;
  assign n2722 = ~n2720 & n2721;
  assign n2723 = n2720 & ~n2721;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = ~n2591 & ~n2594;
  assign n2726 = ~n2724 & n2725;
  assign n2727 = n2724 & ~n2725;
  assign n2728 = ~n2726 & ~n2727;
  assign n2729 = ~n2617 & ~n2661;
  assign n2730 = n2728 & ~n2729;
  assign n2731 = ~n2728 & n2729;
  assign n2732 = ~n2730 & ~n2731;
  assign n2733 = n2715 & ~n2732;
  assign n2734 = ~n2715 & n2732;
  assign n2735 = ~n2733 & ~n2734;
  assign n2736 = ~n2676 & ~n2696;
  assign n2737 = n2608 & n2638;
  assign n2738 = ~n2608 & ~n2638;
  assign n2739 = ~n2737 & ~n2738;
  assign n2740 = ~n2681 & ~n2688;
  assign n2741 = ~n2739 & n2740;
  assign n2742 = n2739 & ~n2740;
  assign n2743 = ~n2741 & ~n2742;
  assign n2744 = ~n2641 & ~n2657;
  assign n2745 = pi34  & n922;
  assign n2746 = pi1  & pi34 ;
  assign n2747 = ~pi18  & ~n2746;
  assign n2748 = ~n2745 & ~n2747;
  assign n2749 = n2654 & ~n2748;
  assign n2750 = ~n2654 & n2748;
  assign n2751 = ~n2749 & ~n2750;
  assign n2752 = ~n2626 & n2751;
  assign n2753 = n2626 & ~n2751;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = ~n2744 & n2754;
  assign n2756 = n2744 & ~n2754;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = n2743 & n2757;
  assign n2759 = ~n2743 & ~n2757;
  assign n2760 = ~n2758 & ~n2759;
  assign n2761 = ~n2736 & n2760;
  assign n2762 = n2736 & ~n2760;
  assign n2763 = ~n2761 & ~n2762;
  assign n2764 = pi8  & pi27 ;
  assign n2765 = pi6  & pi29 ;
  assign n2766 = ~n2764 & ~n2765;
  assign n2767 = n305 & n1923;
  assign n2768 = pi5  & pi30 ;
  assign n2769 = ~n2766 & n2768;
  assign n2770 = ~n2767 & n2769;
  assign n2771 = ~n2767 & ~n2770;
  assign n2772 = ~n2766 & n2771;
  assign n2773 = n2768 & ~n2770;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = pi7  & pi28 ;
  assign n2776 = pi16  & pi19 ;
  assign n2777 = n1199 & n2776;
  assign n2778 = ~n1199 & ~n2776;
  assign n2779 = n2775 & ~n2777;
  assign n2780 = ~n2778 & n2779;
  assign n2781 = n2775 & ~n2780;
  assign n2782 = ~n2777 & ~n2780;
  assign n2783 = ~n2778 & n2782;
  assign n2784 = ~n2781 & ~n2783;
  assign n2785 = ~n2774 & ~n2784;
  assign n2786 = ~n2774 & ~n2785;
  assign n2787 = ~n2784 & ~n2785;
  assign n2788 = ~n2786 & ~n2787;
  assign n2789 = pi4  & pi31 ;
  assign n2790 = n591 & n2310;
  assign n2791 = pi9  & pi26 ;
  assign n2792 = pi10  & pi25 ;
  assign n2793 = ~n2791 & ~n2792;
  assign n2794 = n2789 & ~n2790;
  assign n2795 = ~n2793 & n2794;
  assign n2796 = n2789 & ~n2795;
  assign n2797 = ~n2790 & ~n2795;
  assign n2798 = ~n2793 & n2797;
  assign n2799 = ~n2796 & ~n2798;
  assign n2800 = ~n2788 & ~n2799;
  assign n2801 = ~n2788 & ~n2800;
  assign n2802 = ~n2799 & ~n2800;
  assign n2803 = ~n2801 & ~n2802;
  assign n2804 = ~n2690 & ~n2693;
  assign n2805 = n2803 & n2804;
  assign n2806 = ~n2803 & ~n2804;
  assign n2807 = ~n2805 & ~n2806;
  assign n2808 = pi0  & pi35 ;
  assign n2809 = pi2  & pi33 ;
  assign n2810 = ~n2808 & ~n2809;
  assign n2811 = pi33  & pi35 ;
  assign n2812 = n196 & n2811;
  assign n2813 = n2582 & ~n2810;
  assign n2814 = ~n2812 & n2813;
  assign n2815 = ~n2812 & ~n2814;
  assign n2816 = ~n2810 & n2815;
  assign n2817 = n2582 & ~n2814;
  assign n2818 = ~n2816 & ~n2817;
  assign n2819 = pi3  & pi32 ;
  assign n2820 = n579 & n2110;
  assign n2821 = pi11  & pi24 ;
  assign n2822 = pi12  & pi23 ;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = n2819 & ~n2820;
  assign n2825 = ~n2823 & n2824;
  assign n2826 = n2819 & ~n2825;
  assign n2827 = ~n2820 & ~n2825;
  assign n2828 = ~n2823 & n2827;
  assign n2829 = ~n2826 & ~n2828;
  assign n2830 = ~n2818 & ~n2829;
  assign n2831 = ~n2818 & ~n2830;
  assign n2832 = ~n2829 & ~n2830;
  assign n2833 = ~n2831 & ~n2832;
  assign n2834 = pi13  & pi22 ;
  assign n2835 = n1041 & n1593;
  assign n2836 = pi14  & pi21 ;
  assign n2837 = pi15  & pi20 ;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = n2834 & ~n2835;
  assign n2840 = ~n2838 & n2839;
  assign n2841 = n2834 & ~n2840;
  assign n2842 = ~n2835 & ~n2840;
  assign n2843 = ~n2838 & n2842;
  assign n2844 = ~n2841 & ~n2843;
  assign n2845 = ~n2833 & ~n2844;
  assign n2846 = ~n2833 & ~n2845;
  assign n2847 = ~n2844 & ~n2845;
  assign n2848 = ~n2846 & ~n2847;
  assign n2849 = n2807 & ~n2848;
  assign n2850 = ~n2807 & n2848;
  assign n2851 = ~n2849 & ~n2850;
  assign n2852 = n2763 & n2851;
  assign n2853 = n2763 & ~n2852;
  assign n2854 = n2851 & ~n2852;
  assign n2855 = ~n2853 & ~n2854;
  assign n2856 = ~n2735 & n2855;
  assign n2857 = n2735 & ~n2855;
  assign n2858 = ~n2856 & ~n2857;
  assign n2859 = n2714 & ~n2858;
  assign n2860 = ~n2714 & n2858;
  assign n2861 = ~n2859 & ~n2860;
  assign n2862 = ~n2713 & ~n2861;
  assign n2863 = n2713 & n2861;
  assign po36  = n2862 | n2863;
  assign n2865 = ~n2734 & ~n2857;
  assign n2866 = ~n2761 & ~n2852;
  assign n2867 = ~n2738 & ~n2742;
  assign n2868 = ~n2750 & ~n2752;
  assign n2869 = n2867 & n2868;
  assign n2870 = ~n2867 & ~n2868;
  assign n2871 = ~n2869 & ~n2870;
  assign n2872 = ~n2830 & ~n2845;
  assign n2873 = ~n2871 & n2872;
  assign n2874 = n2871 & ~n2872;
  assign n2875 = ~n2873 & ~n2874;
  assign n2876 = ~n2755 & ~n2758;
  assign n2877 = ~n2875 & n2876;
  assign n2878 = n2875 & ~n2876;
  assign n2879 = ~n2877 & ~n2878;
  assign n2880 = ~n2806 & ~n2849;
  assign n2881 = n2879 & ~n2880;
  assign n2882 = ~n2879 & n2880;
  assign n2883 = ~n2881 & ~n2882;
  assign n2884 = ~n2866 & n2883;
  assign n2885 = n2866 & ~n2883;
  assign n2886 = ~n2884 & ~n2885;
  assign n2887 = pi12  & pi24 ;
  assign n2888 = pi13  & pi23 ;
  assign n2889 = ~n2887 & ~n2888;
  assign n2890 = n952 & n2110;
  assign n2891 = pi2  & pi34 ;
  assign n2892 = ~n2889 & n2891;
  assign n2893 = ~n2890 & n2892;
  assign n2894 = ~n2890 & ~n2893;
  assign n2895 = ~n2889 & n2894;
  assign n2896 = n2891 & ~n2893;
  assign n2897 = ~n2895 & ~n2896;
  assign n2898 = pi10  & pi26 ;
  assign n2899 = pi9  & pi31 ;
  assign n2900 = n2298 & n2899;
  assign n2901 = pi5  & pi31 ;
  assign n2902 = pi9  & pi27 ;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = n2898 & ~n2900;
  assign n2905 = ~n2903 & n2904;
  assign n2906 = n2898 & ~n2905;
  assign n2907 = ~n2900 & ~n2905;
  assign n2908 = ~n2903 & n2907;
  assign n2909 = ~n2906 & ~n2908;
  assign n2910 = ~n2897 & ~n2909;
  assign n2911 = ~n2897 & ~n2910;
  assign n2912 = ~n2909 & ~n2910;
  assign n2913 = ~n2911 & ~n2912;
  assign n2914 = pi6  & pi30 ;
  assign n2915 = pi28  & pi29 ;
  assign n2916 = n521 & n2915;
  assign n2917 = pi7  & pi29 ;
  assign n2918 = pi8  & pi28 ;
  assign n2919 = ~n2917 & ~n2918;
  assign n2920 = n2914 & ~n2916;
  assign n2921 = ~n2919 & n2920;
  assign n2922 = n2914 & ~n2921;
  assign n2923 = ~n2916 & ~n2921;
  assign n2924 = ~n2919 & n2923;
  assign n2925 = ~n2922 & ~n2924;
  assign n2926 = ~n2913 & ~n2925;
  assign n2927 = ~n2913 & ~n2926;
  assign n2928 = ~n2925 & ~n2926;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = ~n2719 & ~n2723;
  assign n2931 = pi0  & pi36 ;
  assign n2932 = n2745 & n2931;
  assign n2933 = n2745 & ~n2932;
  assign n2934 = ~n2745 & n2931;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = pi1  & pi35 ;
  assign n2937 = pi17  & pi19 ;
  assign n2938 = n2936 & n2937;
  assign n2939 = n2936 & ~n2938;
  assign n2940 = n2937 & ~n2938;
  assign n2941 = ~n2939 & ~n2940;
  assign n2942 = ~n2935 & ~n2941;
  assign n2943 = ~n2935 & ~n2942;
  assign n2944 = ~n2941 & ~n2942;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = pi11  & pi25 ;
  assign n2947 = pi4  & pi32 ;
  assign n2948 = ~n2946 & ~n2947;
  assign n2949 = n2946 & n2947;
  assign n2950 = pi3  & pi33 ;
  assign n2951 = ~n2948 & n2950;
  assign n2952 = ~n2949 & n2951;
  assign n2953 = ~n2949 & ~n2952;
  assign n2954 = ~n2948 & n2953;
  assign n2955 = n2950 & ~n2952;
  assign n2956 = ~n2954 & ~n2955;
  assign n2957 = pi14  & pi22 ;
  assign n2958 = n840 & n1593;
  assign n2959 = pi15  & pi21 ;
  assign n2960 = pi16  & pi20 ;
  assign n2961 = ~n2959 & ~n2960;
  assign n2962 = n2957 & ~n2958;
  assign n2963 = ~n2961 & n2962;
  assign n2964 = n2957 & ~n2963;
  assign n2965 = ~n2958 & ~n2963;
  assign n2966 = ~n2961 & n2965;
  assign n2967 = ~n2964 & ~n2966;
  assign n2968 = ~n2956 & ~n2967;
  assign n2969 = ~n2956 & ~n2968;
  assign n2970 = ~n2967 & ~n2968;
  assign n2971 = ~n2969 & ~n2970;
  assign n2972 = ~n2945 & n2971;
  assign n2973 = n2945 & ~n2971;
  assign n2974 = ~n2972 & ~n2973;
  assign n2975 = ~n2930 & ~n2974;
  assign n2976 = ~n2930 & ~n2975;
  assign n2977 = ~n2974 & ~n2975;
  assign n2978 = ~n2976 & ~n2977;
  assign n2979 = ~n2929 & ~n2978;
  assign n2980 = ~n2929 & ~n2979;
  assign n2981 = ~n2978 & ~n2979;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = ~n2727 & ~n2730;
  assign n2984 = n2771 & n2797;
  assign n2985 = ~n2771 & ~n2797;
  assign n2986 = ~n2984 & ~n2985;
  assign n2987 = n2782 & ~n2986;
  assign n2988 = ~n2782 & n2986;
  assign n2989 = ~n2987 & ~n2988;
  assign n2990 = n2827 & n2842;
  assign n2991 = ~n2827 & ~n2842;
  assign n2992 = ~n2990 & ~n2991;
  assign n2993 = n2815 & ~n2992;
  assign n2994 = ~n2815 & n2992;
  assign n2995 = ~n2993 & ~n2994;
  assign n2996 = ~n2785 & ~n2800;
  assign n2997 = ~n2995 & n2996;
  assign n2998 = n2995 & ~n2996;
  assign n2999 = ~n2997 & ~n2998;
  assign n3000 = n2989 & n2999;
  assign n3001 = ~n2989 & ~n2999;
  assign n3002 = ~n3000 & ~n3001;
  assign n3003 = ~n2983 & n3002;
  assign n3004 = ~n2983 & ~n3003;
  assign n3005 = n3002 & ~n3003;
  assign n3006 = ~n3004 & ~n3005;
  assign n3007 = ~n2982 & ~n3006;
  assign n3008 = n2982 & n3006;
  assign n3009 = ~n3007 & ~n3008;
  assign n3010 = n2886 & n3009;
  assign n3011 = ~n2886 & ~n3009;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = n2865 & ~n3012;
  assign n3014 = ~n2865 & n3012;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = ~n2713 & ~n2859;
  assign n3017 = ~n2860 & ~n3016;
  assign n3018 = ~n3015 & n3017;
  assign n3019 = n3015 & ~n3017;
  assign po37  = ~n3018 & ~n3019;
  assign n3021 = ~n2884 & ~n3010;
  assign n3022 = ~n2878 & ~n2881;
  assign n3023 = ~n2932 & ~n2942;
  assign n3024 = n2907 & n3023;
  assign n3025 = ~n2907 & ~n3023;
  assign n3026 = ~n3024 & ~n3025;
  assign n3027 = pi13  & pi24 ;
  assign n3028 = n1041 & n1806;
  assign n3029 = pi14  & pi23 ;
  assign n3030 = pi15  & pi22 ;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = n3027 & ~n3028;
  assign n3033 = ~n3031 & n3032;
  assign n3034 = n3027 & ~n3033;
  assign n3035 = ~n3028 & ~n3033;
  assign n3036 = ~n3031 & n3035;
  assign n3037 = ~n3034 & ~n3036;
  assign n3038 = n3026 & ~n3037;
  assign n3039 = n3026 & ~n3038;
  assign n3040 = ~n3037 & ~n3038;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042 = n2953 & n2965;
  assign n3043 = ~n2953 & ~n2965;
  assign n3044 = ~n3042 & ~n3043;
  assign n3045 = n2894 & ~n3044;
  assign n3046 = ~n2894 & n3044;
  assign n3047 = ~n3045 & ~n3046;
  assign n3048 = ~n2945 & ~n2971;
  assign n3049 = ~n2968 & ~n3048;
  assign n3050 = n3047 & ~n3049;
  assign n3051 = ~n3047 & n3049;
  assign n3052 = ~n3050 & ~n3051;
  assign n3053 = n3041 & n3052;
  assign n3054 = ~n3041 & ~n3052;
  assign n3055 = ~n3053 & ~n3054;
  assign n3056 = ~n3022 & ~n3055;
  assign n3057 = n3022 & n3055;
  assign n3058 = ~n3056 & ~n3057;
  assign n3059 = pi5  & pi32 ;
  assign n3060 = pi10  & pi27 ;
  assign n3061 = ~n3059 & ~n3060;
  assign n3062 = pi10  & pi32 ;
  assign n3063 = n2298 & n3062;
  assign n3064 = pi11  & pi26 ;
  assign n3065 = ~n3061 & n3064;
  assign n3066 = ~n3063 & n3065;
  assign n3067 = ~n3063 & ~n3066;
  assign n3068 = ~n3061 & n3067;
  assign n3069 = n3064 & ~n3066;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = pi8  & pi29 ;
  assign n3072 = n1199 & n1407;
  assign n3073 = pi17  & pi20 ;
  assign n3074 = ~n1085 & ~n3073;
  assign n3075 = n3071 & ~n3072;
  assign n3076 = ~n3074 & n3075;
  assign n3077 = n3071 & ~n3076;
  assign n3078 = ~n3072 & ~n3076;
  assign n3079 = ~n3074 & n3078;
  assign n3080 = ~n3077 & ~n3079;
  assign n3081 = ~n3070 & ~n3080;
  assign n3082 = ~n3070 & ~n3081;
  assign n3083 = ~n3080 & ~n3081;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = ~n2991 & ~n2994;
  assign n3086 = n3084 & n3085;
  assign n3087 = ~n3084 & ~n3085;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = ~n2870 & ~n2874;
  assign n3090 = ~n3088 & n3089;
  assign n3091 = n3088 & ~n3089;
  assign n3092 = ~n3090 & ~n3091;
  assign n3093 = pi4  & pi33 ;
  assign n3094 = pi12  & pi25 ;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = pi25  & pi33 ;
  assign n3097 = n705 & n3096;
  assign n3098 = pi0  & pi37 ;
  assign n3099 = ~n3095 & n3098;
  assign n3100 = ~n3097 & n3099;
  assign n3101 = ~n3097 & ~n3100;
  assign n3102 = ~n3095 & n3101;
  assign n3103 = n3098 & ~n3100;
  assign n3104 = ~n3102 & ~n3103;
  assign n3105 = pi16  & pi21 ;
  assign n3106 = pi34  & pi35 ;
  assign n3107 = n218 & n3106;
  assign n3108 = pi2  & pi35 ;
  assign n3109 = pi3  & pi34 ;
  assign n3110 = ~n3108 & ~n3109;
  assign n3111 = n3105 & ~n3107;
  assign n3112 = ~n3110 & n3111;
  assign n3113 = n3105 & ~n3112;
  assign n3114 = ~n3107 & ~n3112;
  assign n3115 = ~n3110 & n3114;
  assign n3116 = ~n3113 & ~n3115;
  assign n3117 = ~n3104 & ~n3116;
  assign n3118 = ~n3104 & ~n3117;
  assign n3119 = ~n3116 & ~n3117;
  assign n3120 = ~n3118 & ~n3119;
  assign n3121 = pi9  & pi28 ;
  assign n3122 = n432 & n2680;
  assign n3123 = pi6  & pi31 ;
  assign n3124 = pi7  & pi30 ;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = n3121 & ~n3122;
  assign n3127 = ~n3125 & n3126;
  assign n3128 = n3121 & ~n3127;
  assign n3129 = ~n3122 & ~n3127;
  assign n3130 = ~n3125 & n3129;
  assign n3131 = ~n3128 & ~n3130;
  assign n3132 = ~n3120 & ~n3131;
  assign n3133 = ~n3120 & ~n3132;
  assign n3134 = ~n3131 & ~n3132;
  assign n3135 = ~n3133 & ~n3134;
  assign n3136 = ~n3092 & n3135;
  assign n3137 = n3092 & ~n3135;
  assign n3138 = ~n3136 & ~n3137;
  assign n3139 = n3058 & n3138;
  assign n3140 = ~n3058 & ~n3138;
  assign n3141 = ~n3139 & ~n3140;
  assign n3142 = ~n3003 & ~n3007;
  assign n3143 = ~n2975 & ~n2979;
  assign n3144 = ~n2998 & ~n3000;
  assign n3145 = ~n2910 & ~n2926;
  assign n3146 = ~n2985 & ~n2988;
  assign n3147 = pi36  & n1013;
  assign n3148 = pi1  & pi36 ;
  assign n3149 = ~pi19  & ~n3148;
  assign n3150 = ~n3147 & ~n3149;
  assign n3151 = n2938 & n3150;
  assign n3152 = n2938 & ~n3151;
  assign n3153 = n3150 & ~n3151;
  assign n3154 = ~n3152 & ~n3153;
  assign n3155 = ~n2923 & ~n3154;
  assign n3156 = n2923 & ~n3152;
  assign n3157 = ~n3153 & n3156;
  assign n3158 = ~n3155 & ~n3157;
  assign n3159 = ~n3146 & n3158;
  assign n3160 = n3146 & ~n3158;
  assign n3161 = ~n3159 & ~n3160;
  assign n3162 = ~n3145 & n3161;
  assign n3163 = n3145 & ~n3161;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = ~n3144 & n3164;
  assign n3166 = n3144 & ~n3164;
  assign n3167 = ~n3165 & ~n3166;
  assign n3168 = ~n3143 & n3167;
  assign n3169 = n3143 & ~n3167;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = ~n3142 & n3170;
  assign n3172 = ~n3142 & ~n3171;
  assign n3173 = n3170 & ~n3171;
  assign n3174 = ~n3172 & ~n3173;
  assign n3175 = n3141 & ~n3174;
  assign n3176 = ~n3141 & n3174;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = ~n3021 & n3177;
  assign n3179 = n3021 & ~n3177;
  assign n3180 = ~n3178 & ~n3179;
  assign n3181 = ~n3014 & ~n3019;
  assign n3182 = ~n3180 & n3181;
  assign n3183 = n3180 & ~n3181;
  assign po38  = ~n3182 & ~n3183;
  assign n3185 = ~n3171 & ~n3175;
  assign n3186 = ~n3091 & ~n3137;
  assign n3187 = ~n3051 & ~n3053;
  assign n3188 = ~n3186 & n3187;
  assign n3189 = ~n3186 & ~n3188;
  assign n3190 = n3187 & ~n3188;
  assign n3191 = ~n3189 & ~n3190;
  assign n3192 = n3101 & n3114;
  assign n3193 = ~n3101 & ~n3114;
  assign n3194 = ~n3192 & ~n3193;
  assign n3195 = n3035 & ~n3194;
  assign n3196 = ~n3035 & n3194;
  assign n3197 = ~n3195 & ~n3196;
  assign n3198 = ~n3081 & ~n3087;
  assign n3199 = ~n3197 & n3198;
  assign n3200 = n3197 & ~n3198;
  assign n3201 = ~n3199 & ~n3200;
  assign n3202 = pi6  & pi32 ;
  assign n3203 = pi10  & pi28 ;
  assign n3204 = ~n3202 & ~n3203;
  assign n3205 = n3202 & n3203;
  assign n3206 = pi5  & pi33 ;
  assign n3207 = ~n3204 & n3206;
  assign n3208 = ~n3205 & n3207;
  assign n3209 = ~n3205 & ~n3208;
  assign n3210 = ~n3204 & n3209;
  assign n3211 = n3206 & ~n3208;
  assign n3212 = ~n3210 & ~n3211;
  assign n3213 = pi15  & pi23 ;
  assign n3214 = n989 & n1481;
  assign n3215 = pi16  & pi22 ;
  assign n3216 = pi17  & pi21 ;
  assign n3217 = ~n3215 & ~n3216;
  assign n3218 = n3213 & ~n3214;
  assign n3219 = ~n3217 & n3218;
  assign n3220 = n3213 & ~n3219;
  assign n3221 = ~n3214 & ~n3219;
  assign n3222 = ~n3217 & n3221;
  assign n3223 = ~n3220 & ~n3222;
  assign n3224 = ~n3212 & ~n3223;
  assign n3225 = ~n3212 & ~n3224;
  assign n3226 = ~n3223 & ~n3224;
  assign n3227 = ~n3225 & ~n3226;
  assign n3228 = pi9  & pi29 ;
  assign n3229 = n521 & n2680;
  assign n3230 = pi7  & pi31 ;
  assign n3231 = pi8  & pi30 ;
  assign n3232 = ~n3230 & ~n3231;
  assign n3233 = n3228 & ~n3229;
  assign n3234 = ~n3232 & n3233;
  assign n3235 = n3228 & ~n3234;
  assign n3236 = ~n3229 & ~n3234;
  assign n3237 = ~n3232 & n3236;
  assign n3238 = ~n3235 & ~n3237;
  assign n3239 = ~n3227 & ~n3238;
  assign n3240 = ~n3227 & ~n3239;
  assign n3241 = ~n3238 & ~n3239;
  assign n3242 = ~n3240 & ~n3241;
  assign n3243 = n3201 & ~n3242;
  assign n3244 = ~n3201 & n3242;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = ~n3191 & n3245;
  assign n3247 = ~n3191 & ~n3246;
  assign n3248 = n3245 & ~n3246;
  assign n3249 = ~n3247 & ~n3248;
  assign n3250 = ~n3056 & ~n3139;
  assign n3251 = n3249 & n3250;
  assign n3252 = ~n3249 & ~n3250;
  assign n3253 = ~n3251 & ~n3252;
  assign n3254 = ~n3165 & ~n3168;
  assign n3255 = ~n3025 & ~n3038;
  assign n3256 = ~n3117 & ~n3132;
  assign n3257 = n3255 & n3256;
  assign n3258 = ~n3255 & ~n3256;
  assign n3259 = ~n3257 & ~n3258;
  assign n3260 = pi1  & pi37 ;
  assign n3261 = n1257 & n3260;
  assign n3262 = ~n1257 & ~n3260;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = n3078 & ~n3263;
  assign n3265 = ~n3078 & n3263;
  assign n3266 = ~n3264 & ~n3265;
  assign n3267 = ~n3129 & n3266;
  assign n3268 = n3129 & ~n3266;
  assign n3269 = ~n3267 & ~n3268;
  assign n3270 = n3259 & n3269;
  assign n3271 = ~n3259 & ~n3269;
  assign n3272 = ~n3270 & ~n3271;
  assign n3273 = n3254 & ~n3272;
  assign n3274 = ~n3254 & n3272;
  assign n3275 = ~n3273 & ~n3274;
  assign n3276 = ~n3151 & ~n3155;
  assign n3277 = pi12  & pi26 ;
  assign n3278 = pi27  & pi34 ;
  assign n3279 = n619 & n3278;
  assign n3280 = pi4  & pi34 ;
  assign n3281 = pi11  & pi27 ;
  assign n3282 = ~n3280 & ~n3281;
  assign n3283 = n3277 & ~n3279;
  assign n3284 = ~n3282 & n3283;
  assign n3285 = n3277 & ~n3284;
  assign n3286 = ~n3279 & ~n3284;
  assign n3287 = ~n3282 & n3286;
  assign n3288 = ~n3285 & ~n3287;
  assign n3289 = ~n3276 & ~n3288;
  assign n3290 = ~n3276 & ~n3289;
  assign n3291 = ~n3288 & ~n3289;
  assign n3292 = ~n3290 & ~n3291;
  assign n3293 = ~n3043 & ~n3046;
  assign n3294 = n3292 & n3293;
  assign n3295 = ~n3292 & ~n3293;
  assign n3296 = ~n3294 & ~n3295;
  assign n3297 = ~n3159 & ~n3162;
  assign n3298 = pi0  & pi38 ;
  assign n3299 = pi2  & pi36 ;
  assign n3300 = ~n3298 & ~n3299;
  assign n3301 = pi36  & pi38 ;
  assign n3302 = n196 & n3301;
  assign n3303 = n3147 & ~n3300;
  assign n3304 = ~n3302 & n3303;
  assign n3305 = ~n3302 & ~n3304;
  assign n3306 = ~n3300 & n3305;
  assign n3307 = n3147 & ~n3304;
  assign n3308 = ~n3306 & ~n3307;
  assign n3309 = n3067 & ~n3308;
  assign n3310 = ~n3067 & n3308;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = pi3  & pi35 ;
  assign n3313 = n706 & n1789;
  assign n3314 = pi13  & pi25 ;
  assign n3315 = pi14  & pi24 ;
  assign n3316 = ~n3314 & ~n3315;
  assign n3317 = n3312 & ~n3313;
  assign n3318 = ~n3316 & n3317;
  assign n3319 = n3312 & ~n3318;
  assign n3320 = ~n3313 & ~n3318;
  assign n3321 = ~n3316 & n3320;
  assign n3322 = ~n3319 & ~n3321;
  assign n3323 = ~n3311 & ~n3322;
  assign n3324 = n3311 & n3322;
  assign n3325 = ~n3323 & ~n3324;
  assign n3326 = n3297 & ~n3325;
  assign n3327 = ~n3297 & n3325;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = n3296 & n3328;
  assign n3330 = ~n3296 & ~n3328;
  assign n3331 = ~n3329 & ~n3330;
  assign n3332 = n3275 & n3331;
  assign n3333 = ~n3275 & ~n3331;
  assign n3334 = ~n3332 & ~n3333;
  assign n3335 = ~n3253 & ~n3334;
  assign n3336 = n3253 & n3334;
  assign n3337 = ~n3335 & ~n3336;
  assign n3338 = ~n3185 & n3337;
  assign n3339 = n3185 & ~n3337;
  assign n3340 = ~n3338 & ~n3339;
  assign n3341 = ~n3178 & ~n3183;
  assign n3342 = ~n3340 & n3341;
  assign n3343 = n3340 & ~n3341;
  assign po39  = ~n3342 & ~n3343;
  assign n3345 = ~n3252 & ~n3336;
  assign n3346 = ~n3274 & ~n3332;
  assign n3347 = ~n3327 & ~n3329;
  assign n3348 = pi0  & pi39 ;
  assign n3349 = n3261 & n3348;
  assign n3350 = n3261 & ~n3349;
  assign n3351 = ~n3261 & n3348;
  assign n3352 = ~n3350 & ~n3351;
  assign n3353 = pi38  & n1132;
  assign n3354 = pi20  & ~n3353;
  assign n3355 = pi1  & pi38 ;
  assign n3356 = ~n3353 & n3355;
  assign n3357 = ~n3354 & ~n3356;
  assign n3358 = ~n3352 & ~n3357;
  assign n3359 = ~n3352 & ~n3358;
  assign n3360 = ~n3357 & ~n3358;
  assign n3361 = ~n3359 & ~n3360;
  assign n3362 = ~n3265 & ~n3267;
  assign n3363 = n3361 & n3362;
  assign n3364 = ~n3361 & ~n3362;
  assign n3365 = ~n3363 & ~n3364;
  assign n3366 = ~n3193 & ~n3196;
  assign n3367 = ~n3365 & n3366;
  assign n3368 = n3365 & ~n3366;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = n3305 & n3320;
  assign n3371 = ~n3305 & ~n3320;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = n3221 & ~n3372;
  assign n3374 = ~n3221 & n3372;
  assign n3375 = ~n3373 & ~n3374;
  assign n3376 = ~n3224 & ~n3239;
  assign n3377 = ~n3067 & ~n3308;
  assign n3378 = ~n3323 & ~n3377;
  assign n3379 = n3376 & n3378;
  assign n3380 = ~n3376 & ~n3378;
  assign n3381 = ~n3379 & ~n3380;
  assign n3382 = n3375 & n3381;
  assign n3383 = ~n3375 & ~n3381;
  assign n3384 = ~n3382 & ~n3383;
  assign n3385 = n3369 & n3384;
  assign n3386 = ~n3369 & ~n3384;
  assign n3387 = ~n3385 & ~n3386;
  assign n3388 = ~n3347 & n3387;
  assign n3389 = n3347 & ~n3387;
  assign n3390 = ~n3388 & ~n3389;
  assign n3391 = n3346 & ~n3390;
  assign n3392 = ~n3346 & n3390;
  assign n3393 = ~n3391 & ~n3392;
  assign n3394 = ~n3188 & ~n3246;
  assign n3395 = n3236 & n3286;
  assign n3396 = ~n3236 & ~n3286;
  assign n3397 = ~n3395 & ~n3396;
  assign n3398 = n3209 & ~n3397;
  assign n3399 = ~n3209 & n3397;
  assign n3400 = ~n3398 & ~n3399;
  assign n3401 = ~n3289 & ~n3295;
  assign n3402 = ~n3400 & n3401;
  assign n3403 = n3400 & ~n3401;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = pi4  & pi35 ;
  assign n3406 = pi12  & pi27 ;
  assign n3407 = ~n3405 & ~n3406;
  assign n3408 = n3405 & n3406;
  assign n3409 = pi17  & pi22 ;
  assign n3410 = ~n3407 & n3409;
  assign n3411 = ~n3408 & n3410;
  assign n3412 = ~n3408 & ~n3411;
  assign n3413 = ~n3407 & n3412;
  assign n3414 = n3409 & ~n3411;
  assign n3415 = ~n3413 & ~n3414;
  assign n3416 = pi8  & pi31 ;
  assign n3417 = n1085 & n1593;
  assign n3418 = pi18  & pi21 ;
  assign n3419 = ~n1407 & ~n3418;
  assign n3420 = n3416 & ~n3417;
  assign n3421 = ~n3419 & n3420;
  assign n3422 = n3416 & ~n3421;
  assign n3423 = ~n3417 & ~n3421;
  assign n3424 = ~n3419 & n3423;
  assign n3425 = ~n3422 & ~n3424;
  assign n3426 = ~n3415 & ~n3425;
  assign n3427 = ~n3415 & ~n3426;
  assign n3428 = ~n3425 & ~n3426;
  assign n3429 = ~n3427 & ~n3428;
  assign n3430 = pi11  & pi28 ;
  assign n3431 = pi29  & pi34 ;
  assign n3432 = n653 & n3431;
  assign n3433 = pi5  & pi34 ;
  assign n3434 = pi10  & pi29 ;
  assign n3435 = ~n3433 & ~n3434;
  assign n3436 = n3430 & ~n3432;
  assign n3437 = ~n3435 & n3436;
  assign n3438 = n3430 & ~n3437;
  assign n3439 = ~n3432 & ~n3437;
  assign n3440 = ~n3435 & n3439;
  assign n3441 = ~n3438 & ~n3440;
  assign n3442 = ~n3429 & ~n3441;
  assign n3443 = ~n3429 & ~n3442;
  assign n3444 = ~n3441 & ~n3442;
  assign n3445 = ~n3443 & ~n3444;
  assign n3446 = n3404 & ~n3445;
  assign n3447 = ~n3404 & n3445;
  assign n3448 = ~n3446 & ~n3447;
  assign n3449 = ~n3394 & n3448;
  assign n3450 = ~n3394 & ~n3449;
  assign n3451 = n3448 & ~n3449;
  assign n3452 = ~n3450 & ~n3451;
  assign n3453 = pi3  & pi36 ;
  assign n3454 = pi13  & pi26 ;
  assign n3455 = ~n3453 & ~n3454;
  assign n3456 = n3453 & n3454;
  assign n3457 = pi2  & pi37 ;
  assign n3458 = ~n3455 & n3457;
  assign n3459 = ~n3456 & n3458;
  assign n3460 = ~n3456 & ~n3459;
  assign n3461 = ~n3455 & n3460;
  assign n3462 = n3457 & ~n3459;
  assign n3463 = ~n3461 & ~n3462;
  assign n3464 = pi14  & pi25 ;
  assign n3465 = n840 & n2110;
  assign n3466 = pi15  & pi24 ;
  assign n3467 = pi16  & pi23 ;
  assign n3468 = ~n3466 & ~n3467;
  assign n3469 = n3464 & ~n3465;
  assign n3470 = ~n3468 & n3469;
  assign n3471 = n3464 & ~n3470;
  assign n3472 = ~n3465 & ~n3470;
  assign n3473 = ~n3468 & n3472;
  assign n3474 = ~n3471 & ~n3473;
  assign n3475 = ~n3463 & ~n3474;
  assign n3476 = ~n3463 & ~n3475;
  assign n3477 = ~n3474 & ~n3475;
  assign n3478 = ~n3476 & ~n3477;
  assign n3479 = pi6  & pi33 ;
  assign n3480 = n722 & n2332;
  assign n3481 = pi9  & pi30 ;
  assign n3482 = pi7  & pi32 ;
  assign n3483 = ~n3481 & ~n3482;
  assign n3484 = n3479 & ~n3480;
  assign n3485 = ~n3483 & n3484;
  assign n3486 = n3479 & ~n3485;
  assign n3487 = ~n3480 & ~n3485;
  assign n3488 = ~n3483 & n3487;
  assign n3489 = ~n3486 & ~n3488;
  assign n3490 = ~n3478 & ~n3489;
  assign n3491 = ~n3478 & ~n3490;
  assign n3492 = ~n3489 & ~n3490;
  assign n3493 = ~n3491 & ~n3492;
  assign n3494 = ~n3258 & ~n3270;
  assign n3495 = n3493 & n3494;
  assign n3496 = ~n3493 & ~n3494;
  assign n3497 = ~n3495 & ~n3496;
  assign n3498 = ~n3200 & ~n3243;
  assign n3499 = n3497 & ~n3498;
  assign n3500 = ~n3497 & n3498;
  assign n3501 = ~n3499 & ~n3500;
  assign n3502 = n3452 & n3501;
  assign n3503 = ~n3452 & ~n3501;
  assign n3504 = ~n3502 & ~n3503;
  assign n3505 = n3393 & ~n3504;
  assign n3506 = ~n3393 & n3504;
  assign n3507 = ~n3505 & ~n3506;
  assign n3508 = ~n3345 & n3507;
  assign n3509 = n3345 & ~n3507;
  assign n3510 = ~n3508 & ~n3509;
  assign n3511 = ~n3338 & ~n3343;
  assign n3512 = ~n3510 & n3511;
  assign n3513 = n3510 & ~n3511;
  assign po40  = ~n3512 & ~n3513;
  assign n3515 = ~n3392 & ~n3505;
  assign n3516 = ~n3496 & ~n3499;
  assign n3517 = ~n3403 & ~n3446;
  assign n3518 = n3439 & n3460;
  assign n3519 = ~n3439 & ~n3460;
  assign n3520 = ~n3518 & ~n3519;
  assign n3521 = n3412 & ~n3520;
  assign n3522 = ~n3412 & n3520;
  assign n3523 = ~n3521 & ~n3522;
  assign n3524 = ~n3426 & ~n3442;
  assign n3525 = ~n3475 & ~n3490;
  assign n3526 = n3524 & n3525;
  assign n3527 = ~n3524 & ~n3525;
  assign n3528 = ~n3526 & ~n3527;
  assign n3529 = n3523 & n3528;
  assign n3530 = ~n3523 & ~n3528;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = ~n3517 & n3531;
  assign n3533 = n3517 & ~n3531;
  assign n3534 = ~n3532 & ~n3533;
  assign n3535 = ~n3516 & n3534;
  assign n3536 = n3516 & ~n3534;
  assign n3537 = ~n3535 & ~n3536;
  assign n3538 = ~n3452 & n3501;
  assign n3539 = ~n3449 & ~n3538;
  assign n3540 = n3537 & ~n3539;
  assign n3541 = n3537 & ~n3540;
  assign n3542 = ~n3539 & ~n3540;
  assign n3543 = ~n3541 & ~n3542;
  assign n3544 = n3472 & n3487;
  assign n3545 = ~n3472 & ~n3487;
  assign n3546 = ~n3544 & ~n3545;
  assign n3547 = ~n3349 & ~n3358;
  assign n3548 = ~n3546 & n3547;
  assign n3549 = n3546 & ~n3547;
  assign n3550 = ~n3548 & ~n3549;
  assign n3551 = ~n3364 & ~n3368;
  assign n3552 = ~n3550 & n3551;
  assign n3553 = n3550 & ~n3551;
  assign n3554 = ~n3552 & ~n3553;
  assign n3555 = pi0  & pi40 ;
  assign n3556 = pi2  & pi38 ;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = pi38  & pi40 ;
  assign n3559 = n196 & n3558;
  assign n3560 = n1387 & ~n3557;
  assign n3561 = ~n3559 & n3560;
  assign n3562 = ~n3559 & ~n3561;
  assign n3563 = ~n3557 & n3562;
  assign n3564 = n1387 & ~n3561;
  assign n3565 = ~n3563 & ~n3564;
  assign n3566 = pi7  & pi33 ;
  assign n3567 = pi31  & pi32 ;
  assign n3568 = n414 & n3567;
  assign n3569 = pi8  & pi32 ;
  assign n3570 = ~n2899 & ~n3569;
  assign n3571 = n3566 & ~n3568;
  assign n3572 = ~n3570 & n3571;
  assign n3573 = n3566 & ~n3572;
  assign n3574 = ~n3568 & ~n3572;
  assign n3575 = ~n3570 & n3574;
  assign n3576 = ~n3573 & ~n3575;
  assign n3577 = ~n3565 & ~n3576;
  assign n3578 = ~n3565 & ~n3577;
  assign n3579 = ~n3576 & ~n3577;
  assign n3580 = ~n3578 & ~n3579;
  assign n3581 = pi4  & pi36 ;
  assign n3582 = pi5  & pi35 ;
  assign n3583 = pi12  & pi28 ;
  assign n3584 = n3582 & n3583;
  assign n3585 = ~n3582 & ~n3583;
  assign n3586 = n3581 & ~n3584;
  assign n3587 = ~n3585 & n3586;
  assign n3588 = n3581 & ~n3587;
  assign n3589 = ~n3584 & ~n3587;
  assign n3590 = ~n3585 & n3589;
  assign n3591 = ~n3588 & ~n3590;
  assign n3592 = ~n3580 & ~n3591;
  assign n3593 = ~n3580 & ~n3592;
  assign n3594 = ~n3591 & ~n3592;
  assign n3595 = ~n3593 & ~n3594;
  assign n3596 = ~n3554 & n3595;
  assign n3597 = n3554 & ~n3595;
  assign n3598 = ~n3596 & ~n3597;
  assign n3599 = ~n3385 & ~n3388;
  assign n3600 = n3598 & ~n3599;
  assign n3601 = ~n3598 & n3599;
  assign n3602 = ~n3600 & ~n3601;
  assign n3603 = pi13  & pi27 ;
  assign n3604 = pi14  & pi26 ;
  assign n3605 = ~n3603 & ~n3604;
  assign n3606 = n706 & n2646;
  assign n3607 = pi3  & pi37 ;
  assign n3608 = ~n3605 & n3607;
  assign n3609 = ~n3606 & n3608;
  assign n3610 = ~n3606 & ~n3609;
  assign n3611 = ~n3605 & n3610;
  assign n3612 = n3607 & ~n3609;
  assign n3613 = ~n3611 & ~n3612;
  assign n3614 = pi15  & pi25 ;
  assign n3615 = n989 & n2110;
  assign n3616 = pi17  & pi23 ;
  assign n3617 = pi16  & pi24 ;
  assign n3618 = ~n3616 & ~n3617;
  assign n3619 = n3614 & ~n3615;
  assign n3620 = ~n3618 & n3619;
  assign n3621 = n3614 & ~n3620;
  assign n3622 = ~n3615 & ~n3620;
  assign n3623 = ~n3618 & n3622;
  assign n3624 = ~n3621 & ~n3623;
  assign n3625 = ~n3613 & ~n3624;
  assign n3626 = ~n3613 & ~n3625;
  assign n3627 = ~n3624 & ~n3625;
  assign n3628 = ~n3626 & ~n3627;
  assign n3629 = pi11  & pi29 ;
  assign n3630 = pi6  & pi34 ;
  assign n3631 = pi10  & pi30 ;
  assign n3632 = n3630 & n3631;
  assign n3633 = ~n3630 & ~n3631;
  assign n3634 = n3629 & ~n3632;
  assign n3635 = ~n3633 & n3634;
  assign n3636 = n3629 & ~n3635;
  assign n3637 = ~n3632 & ~n3635;
  assign n3638 = ~n3633 & n3637;
  assign n3639 = ~n3636 & ~n3638;
  assign n3640 = ~n3628 & ~n3639;
  assign n3641 = ~n3628 & ~n3640;
  assign n3642 = ~n3639 & ~n3640;
  assign n3643 = ~n3641 & ~n3642;
  assign n3644 = ~n3380 & ~n3382;
  assign n3645 = ~n3643 & ~n3644;
  assign n3646 = n3643 & n3644;
  assign n3647 = ~n3645 & ~n3646;
  assign n3648 = ~n3396 & ~n3399;
  assign n3649 = ~n3371 & ~n3374;
  assign n3650 = n3648 & n3649;
  assign n3651 = ~n3648 & ~n3649;
  assign n3652 = ~n3650 & ~n3651;
  assign n3653 = pi19  & pi21 ;
  assign n3654 = pi1  & pi39 ;
  assign n3655 = n3653 & n3654;
  assign n3656 = ~n3653 & ~n3654;
  assign n3657 = ~n3655 & ~n3656;
  assign n3658 = n3353 & n3657;
  assign n3659 = ~n3353 & ~n3657;
  assign n3660 = ~n3658 & ~n3659;
  assign n3661 = ~n3423 & n3660;
  assign n3662 = n3423 & ~n3660;
  assign n3663 = ~n3661 & ~n3662;
  assign n3664 = n3652 & n3663;
  assign n3665 = ~n3652 & ~n3663;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = n3647 & n3666;
  assign n3668 = ~n3647 & ~n3666;
  assign n3669 = ~n3667 & ~n3668;
  assign n3670 = n3602 & n3669;
  assign n3671 = ~n3602 & ~n3669;
  assign n3672 = ~n3670 & ~n3671;
  assign n3673 = ~n3543 & n3672;
  assign n3674 = n3543 & ~n3672;
  assign n3675 = ~n3673 & ~n3674;
  assign n3676 = ~n3515 & n3675;
  assign n3677 = n3515 & ~n3675;
  assign n3678 = ~n3676 & ~n3677;
  assign n3679 = ~n3508 & ~n3513;
  assign n3680 = ~n3678 & n3679;
  assign n3681 = ~n3677 & ~n3679;
  assign n3682 = ~n3676 & n3681;
  assign po41  = ~n3680 & ~n3682;
  assign n3684 = ~n3540 & ~n3673;
  assign n3685 = ~n3645 & ~n3667;
  assign n3686 = ~n3553 & ~n3597;
  assign n3687 = n3562 & n3622;
  assign n3688 = ~n3562 & ~n3622;
  assign n3689 = ~n3687 & ~n3688;
  assign n3690 = n3610 & ~n3689;
  assign n3691 = ~n3610 & n3689;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = ~n3577 & ~n3592;
  assign n3694 = ~n3692 & n3693;
  assign n3695 = n3692 & ~n3693;
  assign n3696 = ~n3694 & ~n3695;
  assign n3697 = pi40  & n1220;
  assign n3698 = pi1  & pi40 ;
  assign n3699 = ~pi21  & ~n3698;
  assign n3700 = ~n3697 & ~n3699;
  assign n3701 = n3574 & ~n3700;
  assign n3702 = ~n3574 & n3700;
  assign n3703 = ~n3701 & ~n3702;
  assign n3704 = ~n3637 & n3703;
  assign n3705 = n3637 & ~n3703;
  assign n3706 = ~n3704 & ~n3705;
  assign n3707 = n3696 & n3706;
  assign n3708 = ~n3696 & ~n3706;
  assign n3709 = ~n3707 & ~n3708;
  assign n3710 = ~n3686 & n3709;
  assign n3711 = n3686 & ~n3709;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = n3685 & ~n3712;
  assign n3714 = ~n3685 & n3712;
  assign n3715 = ~n3713 & ~n3714;
  assign n3716 = ~n3600 & ~n3670;
  assign n3717 = ~n3715 & n3716;
  assign n3718 = n3715 & ~n3716;
  assign n3719 = ~n3717 & ~n3718;
  assign n3720 = ~n3545 & ~n3549;
  assign n3721 = ~n3519 & ~n3522;
  assign n3722 = n3720 & n3721;
  assign n3723 = ~n3720 & ~n3721;
  assign n3724 = ~n3722 & ~n3723;
  assign n3725 = ~n3625 & ~n3640;
  assign n3726 = ~n3724 & n3725;
  assign n3727 = n3724 & ~n3725;
  assign n3728 = ~n3726 & ~n3727;
  assign n3729 = pi39  & pi41 ;
  assign n3730 = n196 & n3729;
  assign n3731 = pi0  & pi41 ;
  assign n3732 = pi2  & pi39 ;
  assign n3733 = ~n3731 & ~n3732;
  assign n3734 = ~n3730 & ~n3733;
  assign n3735 = n3655 & n3734;
  assign n3736 = ~n3655 & ~n3734;
  assign n3737 = ~n3735 & ~n3736;
  assign n3738 = ~n3589 & n3737;
  assign n3739 = n3589 & ~n3737;
  assign n3740 = ~n3738 & ~n3739;
  assign n3741 = pi3  & pi38 ;
  assign n3742 = pi26  & pi28 ;
  assign n3743 = n777 & n3742;
  assign n3744 = pi13  & pi28 ;
  assign n3745 = pi15  & pi26 ;
  assign n3746 = ~n3744 & ~n3745;
  assign n3747 = n3741 & ~n3743;
  assign n3748 = ~n3746 & n3747;
  assign n3749 = n3741 & ~n3748;
  assign n3750 = ~n3743 & ~n3748;
  assign n3751 = ~n3746 & n3750;
  assign n3752 = ~n3749 & ~n3751;
  assign n3753 = n3740 & ~n3752;
  assign n3754 = n3740 & ~n3753;
  assign n3755 = ~n3752 & ~n3753;
  assign n3756 = ~n3754 & ~n3755;
  assign n3757 = ~n3527 & ~n3529;
  assign n3758 = ~n3756 & ~n3757;
  assign n3759 = ~n3756 & ~n3758;
  assign n3760 = ~n3757 & ~n3758;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = ~n3728 & n3761;
  assign n3763 = n3728 & ~n3761;
  assign n3764 = ~n3762 & ~n3763;
  assign n3765 = ~n3532 & ~n3535;
  assign n3766 = pi6  & pi35 ;
  assign n3767 = pi11  & pi30 ;
  assign n3768 = ~n3766 & ~n3767;
  assign n3769 = pi30  & pi35 ;
  assign n3770 = n776 & n3769;
  assign n3771 = pi5  & pi36 ;
  assign n3772 = ~n3768 & n3771;
  assign n3773 = ~n3770 & n3772;
  assign n3774 = ~n3770 & ~n3773;
  assign n3775 = ~n3768 & n3774;
  assign n3776 = n3771 & ~n3773;
  assign n3777 = ~n3775 & ~n3776;
  assign n3778 = pi8  & pi33 ;
  assign n3779 = pi19  & pi22 ;
  assign n3780 = n1593 & n3779;
  assign n3781 = ~n1593 & ~n3779;
  assign n3782 = n3778 & ~n3780;
  assign n3783 = ~n3781 & n3782;
  assign n3784 = n3778 & ~n3783;
  assign n3785 = ~n3780 & ~n3783;
  assign n3786 = ~n3781 & n3785;
  assign n3787 = ~n3784 & ~n3786;
  assign n3788 = ~n3777 & ~n3787;
  assign n3789 = ~n3777 & ~n3788;
  assign n3790 = ~n3787 & ~n3788;
  assign n3791 = ~n3789 & ~n3790;
  assign n3792 = ~n3658 & ~n3661;
  assign n3793 = n3791 & n3792;
  assign n3794 = ~n3791 & ~n3792;
  assign n3795 = ~n3793 & ~n3794;
  assign n3796 = ~n3651 & ~n3664;
  assign n3797 = ~n3795 & n3796;
  assign n3798 = n3795 & ~n3796;
  assign n3799 = ~n3797 & ~n3798;
  assign n3800 = pi4  & pi37 ;
  assign n3801 = pi12  & pi29 ;
  assign n3802 = ~n3800 & ~n3801;
  assign n3803 = n3800 & n3801;
  assign n3804 = pi14  & pi27 ;
  assign n3805 = ~n3802 & n3804;
  assign n3806 = ~n3803 & n3805;
  assign n3807 = ~n3803 & ~n3806;
  assign n3808 = ~n3802 & n3807;
  assign n3809 = n3804 & ~n3806;
  assign n3810 = ~n3808 & ~n3809;
  assign n3811 = pi16  & pi25 ;
  assign n3812 = n1199 & n2110;
  assign n3813 = pi17  & pi24 ;
  assign n3814 = pi18  & pi23 ;
  assign n3815 = ~n3813 & ~n3814;
  assign n3816 = n3811 & ~n3812;
  assign n3817 = ~n3815 & n3816;
  assign n3818 = n3811 & ~n3817;
  assign n3819 = ~n3812 & ~n3817;
  assign n3820 = ~n3815 & n3819;
  assign n3821 = ~n3818 & ~n3820;
  assign n3822 = ~n3810 & ~n3821;
  assign n3823 = ~n3810 & ~n3822;
  assign n3824 = ~n3821 & ~n3822;
  assign n3825 = ~n3823 & ~n3824;
  assign n3826 = pi10  & pi31 ;
  assign n3827 = pi32  & pi34 ;
  assign n3828 = n722 & n3827;
  assign n3829 = pi7  & pi34 ;
  assign n3830 = pi9  & pi32 ;
  assign n3831 = ~n3829 & ~n3830;
  assign n3832 = n3826 & ~n3828;
  assign n3833 = ~n3831 & n3832;
  assign n3834 = n3826 & ~n3833;
  assign n3835 = ~n3828 & ~n3833;
  assign n3836 = ~n3831 & n3835;
  assign n3837 = ~n3834 & ~n3836;
  assign n3838 = ~n3825 & ~n3837;
  assign n3839 = ~n3825 & ~n3838;
  assign n3840 = ~n3837 & ~n3838;
  assign n3841 = ~n3839 & ~n3840;
  assign n3842 = ~n3799 & n3841;
  assign n3843 = n3799 & ~n3841;
  assign n3844 = ~n3842 & ~n3843;
  assign n3845 = ~n3765 & n3844;
  assign n3846 = ~n3765 & ~n3845;
  assign n3847 = n3844 & ~n3845;
  assign n3848 = ~n3846 & ~n3847;
  assign n3849 = n3764 & ~n3848;
  assign n3850 = ~n3764 & n3848;
  assign n3851 = ~n3849 & ~n3850;
  assign n3852 = n3719 & n3851;
  assign n3853 = ~n3719 & ~n3851;
  assign n3854 = ~n3852 & ~n3853;
  assign n3855 = n3684 & ~n3854;
  assign n3856 = ~n3684 & n3854;
  assign n3857 = ~n3855 & ~n3856;
  assign n3858 = ~n3676 & ~n3681;
  assign n3859 = ~n3857 & n3858;
  assign n3860 = n3857 & ~n3858;
  assign po42  = ~n3859 & ~n3860;
  assign n3862 = ~n3718 & ~n3852;
  assign n3863 = ~n3845 & ~n3849;
  assign n3864 = ~n3758 & ~n3763;
  assign n3865 = ~n3688 & ~n3691;
  assign n3866 = ~n3738 & ~n3753;
  assign n3867 = n3865 & n3866;
  assign n3868 = ~n3865 & ~n3866;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = ~n3822 & ~n3838;
  assign n3871 = ~n3869 & n3870;
  assign n3872 = n3869 & ~n3870;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = ~n3798 & ~n3843;
  assign n3875 = n3873 & ~n3874;
  assign n3876 = ~n3873 & n3874;
  assign n3877 = ~n3875 & ~n3876;
  assign n3878 = ~n3864 & n3877;
  assign n3879 = n3864 & ~n3877;
  assign n3880 = ~n3878 & ~n3879;
  assign n3881 = ~n3863 & n3880;
  assign n3882 = n3863 & ~n3880;
  assign n3883 = ~n3881 & ~n3882;
  assign n3884 = ~n3710 & ~n3714;
  assign n3885 = ~n3723 & ~n3727;
  assign n3886 = pi6  & pi36 ;
  assign n3887 = pi7  & pi35 ;
  assign n3888 = pi11  & pi31 ;
  assign n3889 = n3887 & n3888;
  assign n3890 = ~n3887 & ~n3888;
  assign n3891 = n3886 & ~n3889;
  assign n3892 = ~n3890 & n3891;
  assign n3893 = n3886 & ~n3892;
  assign n3894 = ~n3889 & ~n3892;
  assign n3895 = ~n3890 & n3894;
  assign n3896 = ~n3893 & ~n3895;
  assign n3897 = n3835 & ~n3896;
  assign n3898 = ~n3835 & n3896;
  assign n3899 = ~n3897 & ~n3898;
  assign n3900 = pi33  & pi34 ;
  assign n3901 = n414 & n3900;
  assign n3902 = pi8  & pi34 ;
  assign n3903 = pi9  & pi33 ;
  assign n3904 = ~n3902 & ~n3903;
  assign n3905 = n3062 & ~n3901;
  assign n3906 = ~n3904 & n3905;
  assign n3907 = n3062 & ~n3906;
  assign n3908 = ~n3901 & ~n3906;
  assign n3909 = ~n3904 & n3908;
  assign n3910 = ~n3907 & ~n3909;
  assign n3911 = ~n3899 & ~n3910;
  assign n3912 = n3899 & n3910;
  assign n3913 = ~n3911 & ~n3912;
  assign n3914 = n3885 & ~n3913;
  assign n3915 = ~n3885 & n3913;
  assign n3916 = ~n3914 & ~n3915;
  assign n3917 = pi3  & pi39 ;
  assign n3918 = pi16  & pi26 ;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = n3917 & n3918;
  assign n3921 = pi2  & pi40 ;
  assign n3922 = ~n3919 & n3921;
  assign n3923 = ~n3920 & n3922;
  assign n3924 = ~n3920 & ~n3923;
  assign n3925 = ~n3919 & n3924;
  assign n3926 = n3921 & ~n3923;
  assign n3927 = ~n3925 & ~n3926;
  assign n3928 = pi17  & pi25 ;
  assign n3929 = n1085 & n2110;
  assign n3930 = pi18  & pi24 ;
  assign n3931 = pi19  & pi23 ;
  assign n3932 = ~n3930 & ~n3931;
  assign n3933 = n3928 & ~n3929;
  assign n3934 = ~n3932 & n3933;
  assign n3935 = n3928 & ~n3934;
  assign n3936 = ~n3929 & ~n3934;
  assign n3937 = ~n3932 & n3936;
  assign n3938 = ~n3935 & ~n3937;
  assign n3939 = ~n3927 & ~n3938;
  assign n3940 = ~n3927 & ~n3939;
  assign n3941 = ~n3938 & ~n3939;
  assign n3942 = ~n3940 & ~n3941;
  assign n3943 = pi15  & pi27 ;
  assign n3944 = pi14  & pi38 ;
  assign n3945 = n2299 & n3944;
  assign n3946 = pi4  & pi38 ;
  assign n3947 = pi14  & pi28 ;
  assign n3948 = ~n3946 & ~n3947;
  assign n3949 = n3943 & ~n3945;
  assign n3950 = ~n3948 & n3949;
  assign n3951 = n3943 & ~n3950;
  assign n3952 = ~n3945 & ~n3950;
  assign n3953 = ~n3948 & n3952;
  assign n3954 = ~n3951 & ~n3953;
  assign n3955 = ~n3942 & ~n3954;
  assign n3956 = ~n3942 & ~n3955;
  assign n3957 = ~n3954 & ~n3955;
  assign n3958 = ~n3956 & ~n3957;
  assign n3959 = n3916 & ~n3958;
  assign n3960 = ~n3916 & n3958;
  assign n3961 = ~n3959 & ~n3960;
  assign n3962 = ~n3884 & n3961;
  assign n3963 = ~n3884 & ~n3962;
  assign n3964 = n3961 & ~n3962;
  assign n3965 = ~n3963 & ~n3964;
  assign n3966 = pi0  & pi42 ;
  assign n3967 = n3697 & n3966;
  assign n3968 = n3697 & ~n3967;
  assign n3969 = ~n3697 & n3966;
  assign n3970 = ~n3968 & ~n3969;
  assign n3971 = pi1  & pi41 ;
  assign n3972 = pi20  & pi22 ;
  assign n3973 = n3971 & n3972;
  assign n3974 = n3971 & ~n3973;
  assign n3975 = n3972 & ~n3973;
  assign n3976 = ~n3974 & ~n3975;
  assign n3977 = ~n3970 & ~n3976;
  assign n3978 = ~n3970 & ~n3977;
  assign n3979 = ~n3976 & ~n3977;
  assign n3980 = ~n3978 & ~n3979;
  assign n3981 = pi13  & pi29 ;
  assign n3982 = pi5  & pi37 ;
  assign n3983 = pi12  & pi30 ;
  assign n3984 = n3982 & n3983;
  assign n3985 = ~n3982 & ~n3983;
  assign n3986 = n3981 & ~n3984;
  assign n3987 = ~n3985 & n3986;
  assign n3988 = n3981 & ~n3987;
  assign n3989 = ~n3984 & ~n3987;
  assign n3990 = ~n3985 & n3989;
  assign n3991 = ~n3988 & ~n3990;
  assign n3992 = ~n3980 & ~n3991;
  assign n3993 = ~n3980 & ~n3992;
  assign n3994 = ~n3991 & ~n3992;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = ~n3702 & ~n3704;
  assign n3997 = n3995 & n3996;
  assign n3998 = ~n3995 & ~n3996;
  assign n3999 = ~n3997 & ~n3998;
  assign n4000 = ~n3695 & ~n3707;
  assign n4001 = ~n3999 & n4000;
  assign n4002 = n3999 & ~n4000;
  assign n4003 = ~n4001 & ~n4002;
  assign n4004 = n3785 & n3807;
  assign n4005 = ~n3785 & ~n3807;
  assign n4006 = ~n4004 & ~n4005;
  assign n4007 = n3774 & ~n4006;
  assign n4008 = ~n3774 & n4006;
  assign n4009 = ~n4007 & ~n4008;
  assign n4010 = ~n3788 & ~n3794;
  assign n4011 = ~n4009 & n4010;
  assign n4012 = n4009 & ~n4010;
  assign n4013 = ~n4011 & ~n4012;
  assign n4014 = n3750 & n3819;
  assign n4015 = ~n3750 & ~n3819;
  assign n4016 = ~n4014 & ~n4015;
  assign n4017 = ~n3730 & ~n3735;
  assign n4018 = ~n4016 & n4017;
  assign n4019 = n4016 & ~n4017;
  assign n4020 = ~n4018 & ~n4019;
  assign n4021 = n4013 & n4020;
  assign n4022 = ~n4013 & ~n4020;
  assign n4023 = ~n4021 & ~n4022;
  assign n4024 = n4003 & n4023;
  assign n4025 = ~n4003 & ~n4023;
  assign n4026 = ~n4024 & ~n4025;
  assign n4027 = n3965 & n4026;
  assign n4028 = ~n3965 & ~n4026;
  assign n4029 = ~n4027 & ~n4028;
  assign n4030 = n3883 & ~n4029;
  assign n4031 = n3883 & ~n4030;
  assign n4032 = ~n4029 & ~n4030;
  assign n4033 = ~n4031 & ~n4032;
  assign n4034 = ~n3862 & ~n4033;
  assign n4035 = n3862 & n4033;
  assign n4036 = ~n4034 & ~n4035;
  assign n4037 = ~n3856 & ~n3860;
  assign n4038 = n4036 & ~n4037;
  assign n4039 = ~n4036 & n4037;
  assign po43  = ~n4038 & ~n4039;
  assign n4041 = ~n3881 & ~n4030;
  assign n4042 = ~n3965 & n4026;
  assign n4043 = ~n3962 & ~n4042;
  assign n4044 = ~n4002 & ~n4024;
  assign n4045 = ~n3915 & ~n3959;
  assign n4046 = ~n3939 & ~n3955;
  assign n4047 = ~n3835 & ~n3896;
  assign n4048 = ~n3911 & ~n4047;
  assign n4049 = pi42  & n1324;
  assign n4050 = pi1  & pi42 ;
  assign n4051 = ~pi22  & ~n4050;
  assign n4052 = ~n4049 & ~n4051;
  assign n4053 = n3973 & n4052;
  assign n4054 = ~n3973 & ~n4052;
  assign n4055 = ~n4053 & ~n4054;
  assign n4056 = ~n3908 & n4055;
  assign n4057 = n3908 & ~n4055;
  assign n4058 = ~n4056 & ~n4057;
  assign n4059 = ~n4048 & n4058;
  assign n4060 = ~n4048 & ~n4059;
  assign n4061 = n4058 & ~n4059;
  assign n4062 = ~n4060 & ~n4061;
  assign n4063 = ~n4046 & ~n4062;
  assign n4064 = n4046 & n4062;
  assign n4065 = ~n4063 & ~n4064;
  assign n4066 = ~n4045 & n4065;
  assign n4067 = n4045 & ~n4065;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = ~n4044 & n4068;
  assign n4070 = n4044 & ~n4068;
  assign n4071 = ~n4069 & ~n4070;
  assign n4072 = ~n4043 & n4071;
  assign n4073 = ~n4043 & ~n4072;
  assign n4074 = n4071 & ~n4072;
  assign n4075 = ~n4073 & ~n4074;
  assign n4076 = ~n3875 & ~n3878;
  assign n4077 = ~n3868 & ~n3872;
  assign n4078 = pi0  & pi43 ;
  assign n4079 = pi3  & pi40 ;
  assign n4080 = ~n4078 & ~n4079;
  assign n4081 = n4078 & n4079;
  assign n4082 = pi4  & pi39 ;
  assign n4083 = ~n4080 & n4082;
  assign n4084 = ~n4081 & n4083;
  assign n4085 = ~n4081 & ~n4084;
  assign n4086 = ~n4080 & n4085;
  assign n4087 = n4082 & ~n4084;
  assign n4088 = ~n4086 & ~n4087;
  assign n4089 = pi14  & pi29 ;
  assign n4090 = n840 & n2191;
  assign n4091 = pi15  & pi28 ;
  assign n4092 = pi16  & pi27 ;
  assign n4093 = ~n4091 & ~n4092;
  assign n4094 = n4089 & ~n4090;
  assign n4095 = ~n4093 & n4094;
  assign n4096 = n4089 & ~n4095;
  assign n4097 = ~n4090 & ~n4095;
  assign n4098 = ~n4093 & n4097;
  assign n4099 = ~n4096 & ~n4098;
  assign n4100 = ~n4088 & ~n4099;
  assign n4101 = ~n4088 & ~n4100;
  assign n4102 = ~n4099 & ~n4100;
  assign n4103 = ~n4101 & ~n4102;
  assign n4104 = pi17  & pi26 ;
  assign n4105 = n1085 & n1789;
  assign n4106 = pi19  & pi24 ;
  assign n4107 = pi18  & pi25 ;
  assign n4108 = ~n4106 & ~n4107;
  assign n4109 = n4104 & ~n4105;
  assign n4110 = ~n4108 & n4109;
  assign n4111 = n4104 & ~n4110;
  assign n4112 = ~n4105 & ~n4110;
  assign n4113 = ~n4108 & n4112;
  assign n4114 = ~n4111 & ~n4113;
  assign n4115 = ~n4103 & ~n4114;
  assign n4116 = ~n4103 & ~n4115;
  assign n4117 = ~n4114 & ~n4115;
  assign n4118 = ~n4116 & ~n4117;
  assign n4119 = pi8  & pi35 ;
  assign n4120 = pi10  & pi33 ;
  assign n4121 = ~n4119 & ~n4120;
  assign n4122 = n855 & n2811;
  assign n4123 = pi7  & pi36 ;
  assign n4124 = ~n4121 & n4123;
  assign n4125 = ~n4122 & n4124;
  assign n4126 = ~n4122 & ~n4125;
  assign n4127 = ~n4121 & n4126;
  assign n4128 = n4123 & ~n4125;
  assign n4129 = ~n4127 & ~n4128;
  assign n4130 = pi9  & pi34 ;
  assign n4131 = n1593 & n1806;
  assign n4132 = pi20  & pi23 ;
  assign n4133 = ~n1481 & ~n4132;
  assign n4134 = n4130 & ~n4131;
  assign n4135 = ~n4133 & n4134;
  assign n4136 = n4130 & ~n4135;
  assign n4137 = ~n4131 & ~n4135;
  assign n4138 = ~n4133 & n4137;
  assign n4139 = ~n4136 & ~n4138;
  assign n4140 = ~n4129 & ~n4139;
  assign n4141 = ~n4129 & ~n4140;
  assign n4142 = ~n4139 & ~n4140;
  assign n4143 = ~n4141 & ~n4142;
  assign n4144 = pi2  & pi41 ;
  assign n4145 = pi5  & pi38 ;
  assign n4146 = pi13  & pi30 ;
  assign n4147 = n4145 & n4146;
  assign n4148 = ~n4145 & ~n4146;
  assign n4149 = n4144 & ~n4147;
  assign n4150 = ~n4148 & n4149;
  assign n4151 = n4144 & ~n4150;
  assign n4152 = ~n4147 & ~n4150;
  assign n4153 = ~n4148 & n4152;
  assign n4154 = ~n4151 & ~n4153;
  assign n4155 = ~n4143 & ~n4154;
  assign n4156 = ~n4143 & ~n4155;
  assign n4157 = ~n4154 & ~n4155;
  assign n4158 = ~n4156 & ~n4157;
  assign n4159 = ~n4118 & n4158;
  assign n4160 = n4118 & ~n4158;
  assign n4161 = ~n4159 & ~n4160;
  assign n4162 = ~n4077 & ~n4161;
  assign n4163 = n4077 & n4161;
  assign n4164 = ~n4162 & ~n4163;
  assign n4165 = ~n4076 & n4164;
  assign n4166 = n4076 & ~n4164;
  assign n4167 = ~n4165 & ~n4166;
  assign n4168 = ~n3992 & ~n3998;
  assign n4169 = n3894 & n3952;
  assign n4170 = ~n3894 & ~n3952;
  assign n4171 = ~n4169 & ~n4170;
  assign n4172 = n3936 & ~n4171;
  assign n4173 = ~n3936 & n4171;
  assign n4174 = ~n4172 & ~n4173;
  assign n4175 = n3924 & n3989;
  assign n4176 = ~n3924 & ~n3989;
  assign n4177 = ~n4175 & ~n4176;
  assign n4178 = ~n3967 & ~n3977;
  assign n4179 = ~n4177 & n4178;
  assign n4180 = n4177 & ~n4178;
  assign n4181 = ~n4179 & ~n4180;
  assign n4182 = ~n4174 & ~n4181;
  assign n4183 = n4174 & n4181;
  assign n4184 = ~n4182 & ~n4183;
  assign n4185 = ~n4168 & n4184;
  assign n4186 = n4168 & ~n4184;
  assign n4187 = ~n4185 & ~n4186;
  assign n4188 = ~n4005 & ~n4008;
  assign n4189 = pi12  & pi31 ;
  assign n4190 = pi6  & pi37 ;
  assign n4191 = pi11  & pi32 ;
  assign n4192 = n4190 & n4191;
  assign n4193 = ~n4190 & ~n4191;
  assign n4194 = n4189 & ~n4192;
  assign n4195 = ~n4193 & n4194;
  assign n4196 = n4189 & ~n4195;
  assign n4197 = ~n4192 & ~n4195;
  assign n4198 = ~n4193 & n4197;
  assign n4199 = ~n4196 & ~n4198;
  assign n4200 = ~n4188 & ~n4199;
  assign n4201 = ~n4188 & ~n4200;
  assign n4202 = ~n4199 & ~n4200;
  assign n4203 = ~n4201 & ~n4202;
  assign n4204 = ~n4015 & ~n4019;
  assign n4205 = n4203 & n4204;
  assign n4206 = ~n4203 & ~n4204;
  assign n4207 = ~n4205 & ~n4206;
  assign n4208 = ~n4012 & ~n4021;
  assign n4209 = n4207 & ~n4208;
  assign n4210 = ~n4207 & n4208;
  assign n4211 = ~n4209 & ~n4210;
  assign n4212 = n4187 & n4211;
  assign n4213 = ~n4187 & ~n4211;
  assign n4214 = ~n4212 & ~n4213;
  assign n4215 = n4167 & n4214;
  assign n4216 = ~n4167 & ~n4214;
  assign n4217 = ~n4215 & ~n4216;
  assign n4218 = ~n4075 & n4217;
  assign n4219 = n4075 & ~n4217;
  assign n4220 = ~n4218 & ~n4219;
  assign n4221 = ~n4041 & n4220;
  assign n4222 = n4041 & ~n4220;
  assign n4223 = ~n4221 & ~n4222;
  assign n4224 = ~n4034 & ~n4038;
  assign n4225 = ~n4223 & n4224;
  assign n4226 = n4223 & ~n4224;
  assign po44  = ~n4225 & ~n4226;
  assign n4228 = ~n4072 & ~n4218;
  assign n4229 = ~n4066 & ~n4069;
  assign n4230 = ~n4059 & ~n4063;
  assign n4231 = pi15  & pi29 ;
  assign n4232 = pi17  & pi27 ;
  assign n4233 = ~n4231 & ~n4232;
  assign n4234 = n942 & n1923;
  assign n4235 = pi3  & pi41 ;
  assign n4236 = ~n4233 & n4235;
  assign n4237 = ~n4234 & n4236;
  assign n4238 = ~n4234 & ~n4237;
  assign n4239 = ~n4233 & n4238;
  assign n4240 = n4235 & ~n4237;
  assign n4241 = ~n4239 & ~n4240;
  assign n4242 = pi18  & pi26 ;
  assign n4243 = n1407 & n1789;
  assign n4244 = pi19  & pi25 ;
  assign n4245 = pi20  & pi24 ;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = n4242 & ~n4243;
  assign n4248 = ~n4246 & n4247;
  assign n4249 = n4242 & ~n4248;
  assign n4250 = ~n4243 & ~n4248;
  assign n4251 = ~n4246 & n4250;
  assign n4252 = ~n4249 & ~n4251;
  assign n4253 = ~n4241 & ~n4252;
  assign n4254 = ~n4241 & ~n4253;
  assign n4255 = ~n4252 & ~n4253;
  assign n4256 = ~n4254 & ~n4255;
  assign n4257 = pi6  & pi38 ;
  assign n4258 = pi11  & pi37 ;
  assign n4259 = n3566 & n4258;
  assign n4260 = pi7  & pi37 ;
  assign n4261 = pi11  & pi33 ;
  assign n4262 = ~n4260 & ~n4261;
  assign n4263 = n4257 & ~n4259;
  assign n4264 = ~n4262 & n4263;
  assign n4265 = n4257 & ~n4264;
  assign n4266 = ~n4259 & ~n4264;
  assign n4267 = ~n4262 & n4266;
  assign n4268 = ~n4265 & ~n4267;
  assign n4269 = ~n4256 & ~n4268;
  assign n4270 = ~n4256 & ~n4269;
  assign n4271 = ~n4268 & ~n4269;
  assign n4272 = ~n4270 & ~n4271;
  assign n4273 = pi4  & pi40 ;
  assign n4274 = pi14  & pi30 ;
  assign n4275 = ~n4273 & ~n4274;
  assign n4276 = n4273 & n4274;
  assign n4277 = pi16  & pi28 ;
  assign n4278 = ~n4275 & n4277;
  assign n4279 = ~n4276 & n4278;
  assign n4280 = ~n4276 & ~n4279;
  assign n4281 = ~n4275 & n4280;
  assign n4282 = n4277 & ~n4279;
  assign n4283 = ~n4281 & ~n4282;
  assign n4284 = pi8  & pi36 ;
  assign n4285 = n591 & n3106;
  assign n4286 = pi9  & pi35 ;
  assign n4287 = pi10  & pi34 ;
  assign n4288 = ~n4286 & ~n4287;
  assign n4289 = n4284 & ~n4285;
  assign n4290 = ~n4288 & n4289;
  assign n4291 = n4284 & ~n4290;
  assign n4292 = ~n4285 & ~n4290;
  assign n4293 = ~n4288 & n4292;
  assign n4294 = ~n4291 & ~n4293;
  assign n4295 = ~n4283 & ~n4294;
  assign n4296 = ~n4283 & ~n4295;
  assign n4297 = ~n4294 & ~n4295;
  assign n4298 = ~n4296 & ~n4297;
  assign n4299 = pi5  & pi39 ;
  assign n4300 = n952 & n3567;
  assign n4301 = pi12  & pi32 ;
  assign n4302 = pi13  & pi31 ;
  assign n4303 = ~n4301 & ~n4302;
  assign n4304 = n4299 & ~n4300;
  assign n4305 = ~n4303 & n4304;
  assign n4306 = n4299 & ~n4305;
  assign n4307 = ~n4300 & ~n4305;
  assign n4308 = ~n4303 & n4307;
  assign n4309 = ~n4306 & ~n4308;
  assign n4310 = ~n4298 & ~n4309;
  assign n4311 = ~n4298 & ~n4310;
  assign n4312 = ~n4309 & ~n4310;
  assign n4313 = ~n4311 & ~n4312;
  assign n4314 = n4272 & n4313;
  assign n4315 = ~n4272 & ~n4313;
  assign n4316 = ~n4314 & ~n4315;
  assign n4317 = ~n4230 & n4316;
  assign n4318 = n4230 & ~n4316;
  assign n4319 = ~n4317 & ~n4318;
  assign n4320 = n4229 & ~n4319;
  assign n4321 = ~n4229 & n4319;
  assign n4322 = ~n4320 & ~n4321;
  assign n4323 = n4097 & n4197;
  assign n4324 = ~n4097 & ~n4197;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = pi0  & pi44 ;
  assign n4327 = pi2  & pi42 ;
  assign n4328 = ~n4326 & ~n4327;
  assign n4329 = pi42  & pi44 ;
  assign n4330 = n196 & n4329;
  assign n4331 = n4049 & ~n4328;
  assign n4332 = ~n4330 & n4331;
  assign n4333 = n4049 & ~n4332;
  assign n4334 = ~n4330 & ~n4332;
  assign n4335 = ~n4328 & n4334;
  assign n4336 = ~n4333 & ~n4335;
  assign n4337 = n4325 & ~n4336;
  assign n4338 = n4325 & ~n4337;
  assign n4339 = ~n4336 & ~n4337;
  assign n4340 = ~n4338 & ~n4339;
  assign n4341 = pi1  & pi43 ;
  assign n4342 = ~n1287 & ~n4341;
  assign n4343 = n1287 & n4341;
  assign n4344 = ~n4342 & ~n4343;
  assign n4345 = n4137 & ~n4344;
  assign n4346 = ~n4137 & n4344;
  assign n4347 = ~n4345 & ~n4346;
  assign n4348 = ~n4126 & n4347;
  assign n4349 = n4126 & ~n4347;
  assign n4350 = ~n4348 & ~n4349;
  assign n4351 = ~n4340 & n4350;
  assign n4352 = ~n4340 & ~n4351;
  assign n4353 = n4350 & ~n4351;
  assign n4354 = ~n4352 & ~n4353;
  assign n4355 = ~n4200 & ~n4206;
  assign n4356 = n4354 & n4355;
  assign n4357 = ~n4354 & ~n4355;
  assign n4358 = ~n4356 & ~n4357;
  assign n4359 = ~n4183 & ~n4185;
  assign n4360 = ~n4176 & ~n4180;
  assign n4361 = ~n4053 & ~n4056;
  assign n4362 = n4360 & n4361;
  assign n4363 = ~n4360 & ~n4361;
  assign n4364 = ~n4362 & ~n4363;
  assign n4365 = ~n4170 & ~n4173;
  assign n4366 = ~n4364 & n4365;
  assign n4367 = n4364 & ~n4365;
  assign n4368 = ~n4366 & ~n4367;
  assign n4369 = ~n4359 & n4368;
  assign n4370 = n4359 & ~n4368;
  assign n4371 = ~n4369 & ~n4370;
  assign n4372 = ~n4358 & ~n4371;
  assign n4373 = n4358 & n4371;
  assign n4374 = ~n4372 & ~n4373;
  assign n4375 = n4322 & n4374;
  assign n4376 = n4322 & ~n4375;
  assign n4377 = n4374 & ~n4375;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = ~n4165 & ~n4215;
  assign n4380 = ~n4209 & ~n4212;
  assign n4381 = ~n4118 & ~n4158;
  assign n4382 = ~n4162 & ~n4381;
  assign n4383 = n4085 & n4152;
  assign n4384 = ~n4085 & ~n4152;
  assign n4385 = ~n4383 & ~n4384;
  assign n4386 = n4112 & ~n4385;
  assign n4387 = ~n4112 & n4385;
  assign n4388 = ~n4386 & ~n4387;
  assign n4389 = ~n4140 & ~n4155;
  assign n4390 = ~n4100 & ~n4115;
  assign n4391 = n4389 & n4390;
  assign n4392 = ~n4389 & ~n4390;
  assign n4393 = ~n4391 & ~n4392;
  assign n4394 = n4388 & n4393;
  assign n4395 = ~n4388 & ~n4393;
  assign n4396 = ~n4394 & ~n4395;
  assign n4397 = ~n4382 & n4396;
  assign n4398 = n4382 & ~n4396;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = ~n4380 & n4399;
  assign n4401 = n4380 & ~n4399;
  assign n4402 = ~n4400 & ~n4401;
  assign n4403 = ~n4379 & n4402;
  assign n4404 = n4379 & ~n4402;
  assign n4405 = ~n4403 & ~n4404;
  assign n4406 = ~n4378 & ~n4405;
  assign n4407 = n4378 & n4405;
  assign n4408 = ~n4406 & ~n4407;
  assign n4409 = ~n4228 & ~n4408;
  assign n4410 = n4228 & n4408;
  assign n4411 = ~n4409 & ~n4410;
  assign n4412 = ~n4221 & ~n4226;
  assign n4413 = ~n4411 & n4412;
  assign n4414 = n4411 & ~n4412;
  assign po45  = ~n4413 & ~n4414;
  assign n4416 = ~n4315 & ~n4317;
  assign n4417 = ~n4369 & ~n4373;
  assign n4418 = ~n4416 & n4417;
  assign n4419 = n4416 & ~n4417;
  assign n4420 = ~n4418 & ~n4419;
  assign n4421 = n4238 & n4334;
  assign n4422 = ~n4238 & ~n4334;
  assign n4423 = ~n4421 & ~n4422;
  assign n4424 = n4250 & ~n4423;
  assign n4425 = ~n4250 & n4423;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = ~n4363 & ~n4367;
  assign n4428 = ~n4426 & n4427;
  assign n4429 = n4426 & ~n4427;
  assign n4430 = ~n4428 & ~n4429;
  assign n4431 = pi11  & pi34 ;
  assign n4432 = pi6  & pi39 ;
  assign n4433 = ~n4431 & ~n4432;
  assign n4434 = pi34  & pi39 ;
  assign n4435 = n776 & n4434;
  assign n4436 = pi12  & pi33 ;
  assign n4437 = ~n4433 & n4436;
  assign n4438 = ~n4435 & n4437;
  assign n4439 = ~n4435 & ~n4438;
  assign n4440 = ~n4433 & n4439;
  assign n4441 = n4436 & ~n4438;
  assign n4442 = ~n4440 & ~n4441;
  assign n4443 = pi15  & pi30 ;
  assign n4444 = n989 & n2915;
  assign n4445 = pi16  & pi29 ;
  assign n4446 = pi17  & pi28 ;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = n4443 & ~n4444;
  assign n4449 = ~n4447 & n4448;
  assign n4450 = n4443 & ~n4449;
  assign n4451 = ~n4444 & ~n4449;
  assign n4452 = ~n4447 & n4451;
  assign n4453 = ~n4450 & ~n4452;
  assign n4454 = ~n4442 & ~n4453;
  assign n4455 = ~n4442 & ~n4454;
  assign n4456 = ~n4453 & ~n4454;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = pi44  & n1376;
  assign n4459 = pi1  & pi44 ;
  assign n4460 = ~n4458 & n4459;
  assign n4461 = pi23  & ~n4458;
  assign n4462 = ~n4460 & ~n4461;
  assign n4463 = pi3  & pi42 ;
  assign n4464 = ~n4343 & ~n4463;
  assign n4465 = n4343 & n4463;
  assign n4466 = ~n4464 & ~n4465;
  assign n4467 = ~n4462 & n4466;
  assign n4468 = ~n4462 & ~n4467;
  assign n4469 = ~n4465 & ~n4467;
  assign n4470 = ~n4464 & n4469;
  assign n4471 = ~n4468 & ~n4470;
  assign n4472 = ~n4457 & ~n4471;
  assign n4473 = ~n4457 & ~n4472;
  assign n4474 = ~n4471 & ~n4472;
  assign n4475 = ~n4473 & ~n4474;
  assign n4476 = n4430 & ~n4475;
  assign n4477 = ~n4430 & n4475;
  assign n4478 = ~n4476 & ~n4477;
  assign n4479 = ~n4420 & n4478;
  assign n4480 = ~n4420 & ~n4479;
  assign n4481 = n4478 & ~n4479;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = ~n4321 & ~n4375;
  assign n4484 = n4482 & n4483;
  assign n4485 = ~n4482 & ~n4483;
  assign n4486 = ~n4484 & ~n4485;
  assign n4487 = pi2  & pi43 ;
  assign n4488 = pi4  & pi41 ;
  assign n4489 = ~n4487 & ~n4488;
  assign n4490 = pi41  & pi43 ;
  assign n4491 = n249 & n4490;
  assign n4492 = pi0  & pi45 ;
  assign n4493 = ~n4489 & n4492;
  assign n4494 = ~n4491 & n4493;
  assign n4495 = ~n4491 & ~n4494;
  assign n4496 = ~n4489 & n4495;
  assign n4497 = n4492 & ~n4494;
  assign n4498 = ~n4496 & ~n4497;
  assign n4499 = pi7  & pi38 ;
  assign n4500 = pi36  & pi37 ;
  assign n4501 = n414 & n4500;
  assign n4502 = pi8  & pi37 ;
  assign n4503 = pi9  & pi36 ;
  assign n4504 = ~n4502 & ~n4503;
  assign n4505 = n4499 & ~n4501;
  assign n4506 = ~n4504 & n4505;
  assign n4507 = n4499 & ~n4506;
  assign n4508 = ~n4501 & ~n4506;
  assign n4509 = ~n4504 & n4508;
  assign n4510 = ~n4507 & ~n4509;
  assign n4511 = ~n4498 & ~n4510;
  assign n4512 = ~n4498 & ~n4511;
  assign n4513 = ~n4510 & ~n4511;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = pi10  & pi35 ;
  assign n4516 = n1481 & n2110;
  assign n4517 = pi21  & pi24 ;
  assign n4518 = ~n1806 & ~n4517;
  assign n4519 = n4515 & ~n4516;
  assign n4520 = ~n4518 & n4519;
  assign n4521 = n4515 & ~n4520;
  assign n4522 = ~n4516 & ~n4520;
  assign n4523 = ~n4518 & n4522;
  assign n4524 = ~n4521 & ~n4523;
  assign n4525 = ~n4514 & ~n4524;
  assign n4526 = ~n4514 & ~n4525;
  assign n4527 = ~n4524 & ~n4525;
  assign n4528 = ~n4526 & ~n4527;
  assign n4529 = pi5  & pi40 ;
  assign n4530 = pi13  & pi32 ;
  assign n4531 = ~n4529 & ~n4530;
  assign n4532 = n4529 & n4530;
  assign n4533 = pi14  & pi31 ;
  assign n4534 = ~n4531 & n4533;
  assign n4535 = ~n4532 & n4534;
  assign n4536 = ~n4532 & ~n4535;
  assign n4537 = ~n4531 & n4536;
  assign n4538 = n4533 & ~n4535;
  assign n4539 = ~n4537 & ~n4538;
  assign n4540 = pi18  & pi27 ;
  assign n4541 = n1407 & n2310;
  assign n4542 = pi19  & pi26 ;
  assign n4543 = ~n1733 & ~n4542;
  assign n4544 = n4540 & ~n4541;
  assign n4545 = ~n4543 & n4544;
  assign n4546 = n4540 & ~n4545;
  assign n4547 = ~n4541 & ~n4545;
  assign n4548 = ~n4543 & n4547;
  assign n4549 = ~n4546 & ~n4548;
  assign n4550 = ~n4292 & ~n4549;
  assign n4551 = ~n4292 & ~n4550;
  assign n4552 = ~n4549 & ~n4550;
  assign n4553 = ~n4551 & ~n4552;
  assign n4554 = ~n4539 & ~n4553;
  assign n4555 = ~n4539 & ~n4554;
  assign n4556 = ~n4553 & ~n4554;
  assign n4557 = ~n4555 & ~n4556;
  assign n4558 = ~n4528 & ~n4557;
  assign n4559 = ~n4528 & ~n4558;
  assign n4560 = ~n4557 & ~n4558;
  assign n4561 = ~n4559 & ~n4560;
  assign n4562 = ~n4392 & ~n4394;
  assign n4563 = ~n4561 & ~n4562;
  assign n4564 = ~n4561 & ~n4563;
  assign n4565 = ~n4562 & ~n4563;
  assign n4566 = ~n4564 & ~n4565;
  assign n4567 = ~n4397 & ~n4400;
  assign n4568 = n4566 & n4567;
  assign n4569 = ~n4566 & ~n4567;
  assign n4570 = ~n4568 & ~n4569;
  assign n4571 = ~n4324 & ~n4337;
  assign n4572 = ~n4384 & ~n4387;
  assign n4573 = n4571 & n4572;
  assign n4574 = ~n4571 & ~n4572;
  assign n4575 = ~n4573 & ~n4574;
  assign n4576 = ~n4346 & ~n4348;
  assign n4577 = ~n4575 & n4576;
  assign n4578 = n4575 & ~n4576;
  assign n4579 = ~n4577 & ~n4578;
  assign n4580 = ~n4351 & ~n4357;
  assign n4581 = ~n4579 & n4580;
  assign n4582 = n4579 & ~n4580;
  assign n4583 = ~n4581 & ~n4582;
  assign n4584 = n4266 & n4280;
  assign n4585 = ~n4266 & ~n4280;
  assign n4586 = ~n4584 & ~n4585;
  assign n4587 = n4307 & ~n4586;
  assign n4588 = ~n4307 & n4586;
  assign n4589 = ~n4587 & ~n4588;
  assign n4590 = ~n4295 & ~n4310;
  assign n4591 = ~n4253 & ~n4269;
  assign n4592 = n4590 & n4591;
  assign n4593 = ~n4590 & ~n4591;
  assign n4594 = ~n4592 & ~n4593;
  assign n4595 = n4589 & n4594;
  assign n4596 = ~n4589 & ~n4594;
  assign n4597 = ~n4595 & ~n4596;
  assign n4598 = n4583 & n4597;
  assign n4599 = ~n4583 & ~n4597;
  assign n4600 = ~n4598 & ~n4599;
  assign n4601 = n4570 & n4600;
  assign n4602 = ~n4570 & ~n4600;
  assign n4603 = ~n4601 & ~n4602;
  assign n4604 = n4486 & n4603;
  assign n4605 = n4486 & ~n4604;
  assign n4606 = n4603 & ~n4604;
  assign n4607 = ~n4605 & ~n4606;
  assign n4608 = ~n4404 & ~n4407;
  assign n4609 = ~n4607 & n4608;
  assign n4610 = n4607 & ~n4608;
  assign n4611 = ~n4609 & ~n4610;
  assign n4612 = ~n4409 & ~n4414;
  assign n4613 = ~n4611 & n4612;
  assign n4614 = n4611 & ~n4612;
  assign po46  = ~n4613 & ~n4614;
  assign n4616 = ~n4485 & ~n4604;
  assign n4617 = ~n4569 & ~n4601;
  assign n4618 = ~n4582 & ~n4598;
  assign n4619 = ~n4558 & ~n4563;
  assign n4620 = n4618 & n4619;
  assign n4621 = ~n4618 & ~n4619;
  assign n4622 = ~n4620 & ~n4621;
  assign n4623 = pi5  & pi41 ;
  assign n4624 = pi15  & pi31 ;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = pi31  & pi41 ;
  assign n4627 = n1043 & n4626;
  assign n4628 = pi2  & pi44 ;
  assign n4629 = ~n4625 & n4628;
  assign n4630 = ~n4627 & n4629;
  assign n4631 = ~n4627 & ~n4630;
  assign n4632 = ~n4625 & n4631;
  assign n4633 = n4628 & ~n4630;
  assign n4634 = ~n4632 & ~n4633;
  assign n4635 = pi14  & pi32 ;
  assign n4636 = pi6  & pi40 ;
  assign n4637 = pi13  & pi33 ;
  assign n4638 = n4636 & n4637;
  assign n4639 = ~n4636 & ~n4637;
  assign n4640 = n4635 & ~n4638;
  assign n4641 = ~n4639 & n4640;
  assign n4642 = n4635 & ~n4641;
  assign n4643 = ~n4638 & ~n4641;
  assign n4644 = ~n4639 & n4643;
  assign n4645 = ~n4642 & ~n4644;
  assign n4646 = ~n4634 & ~n4645;
  assign n4647 = ~n4634 & ~n4646;
  assign n4648 = ~n4645 & ~n4646;
  assign n4649 = ~n4647 & ~n4648;
  assign n4650 = ~n4585 & ~n4588;
  assign n4651 = n4649 & n4650;
  assign n4652 = ~n4649 & ~n4650;
  assign n4653 = ~n4651 & ~n4652;
  assign n4654 = n4451 & n4547;
  assign n4655 = ~n4451 & ~n4547;
  assign n4656 = ~n4654 & ~n4655;
  assign n4657 = n4439 & ~n4656;
  assign n4658 = ~n4439 & n4656;
  assign n4659 = ~n4657 & ~n4658;
  assign n4660 = ~n4574 & ~n4578;
  assign n4661 = ~n4659 & n4660;
  assign n4662 = n4659 & ~n4660;
  assign n4663 = ~n4661 & ~n4662;
  assign n4664 = n4653 & n4663;
  assign n4665 = ~n4653 & ~n4663;
  assign n4666 = ~n4664 & ~n4665;
  assign n4667 = n4622 & n4666;
  assign n4668 = ~n4622 & ~n4666;
  assign n4669 = ~n4667 & ~n4668;
  assign n4670 = ~n4617 & n4669;
  assign n4671 = n4617 & ~n4669;
  assign n4672 = ~n4670 & ~n4671;
  assign n4673 = n4616 & ~n4672;
  assign n4674 = ~n4616 & n4672;
  assign n4675 = ~n4673 & ~n4674;
  assign n4676 = ~n4416 & ~n4417;
  assign n4677 = ~n4479 & ~n4676;
  assign n4678 = ~n4593 & ~n4595;
  assign n4679 = pi0  & pi46 ;
  assign n4680 = pi4  & pi42 ;
  assign n4681 = ~n4679 & ~n4680;
  assign n4682 = n4679 & n4680;
  assign n4683 = pi3  & pi43 ;
  assign n4684 = ~n4681 & n4683;
  assign n4685 = ~n4682 & n4684;
  assign n4686 = ~n4682 & ~n4685;
  assign n4687 = ~n4681 & n4686;
  assign n4688 = n4683 & ~n4685;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = pi9  & pi37 ;
  assign n4691 = pi35  & pi36 ;
  assign n4692 = n1111 & n4691;
  assign n4693 = pi10  & pi36 ;
  assign n4694 = pi11  & pi35 ;
  assign n4695 = ~n4693 & ~n4694;
  assign n4696 = n4690 & ~n4692;
  assign n4697 = ~n4695 & n4696;
  assign n4698 = n4690 & ~n4697;
  assign n4699 = ~n4692 & ~n4697;
  assign n4700 = ~n4695 & n4699;
  assign n4701 = ~n4698 & ~n4700;
  assign n4702 = ~n4689 & ~n4701;
  assign n4703 = ~n4689 & ~n4702;
  assign n4704 = ~n4701 & ~n4702;
  assign n4705 = ~n4703 & ~n4704;
  assign n4706 = pi19  & pi27 ;
  assign n4707 = n1593 & n2310;
  assign n4708 = pi20  & pi26 ;
  assign n4709 = pi21  & pi25 ;
  assign n4710 = ~n4708 & ~n4709;
  assign n4711 = n4706 & ~n4707;
  assign n4712 = ~n4710 & n4711;
  assign n4713 = n4706 & ~n4712;
  assign n4714 = ~n4707 & ~n4712;
  assign n4715 = ~n4710 & n4714;
  assign n4716 = ~n4713 & ~n4715;
  assign n4717 = ~n4705 & ~n4716;
  assign n4718 = ~n4705 & ~n4717;
  assign n4719 = ~n4716 & ~n4717;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = pi16  & pi30 ;
  assign n4722 = n1199 & n2915;
  assign n4723 = pi17  & pi29 ;
  assign n4724 = pi18  & pi28 ;
  assign n4725 = ~n4723 & ~n4724;
  assign n4726 = n4721 & ~n4722;
  assign n4727 = ~n4725 & n4726;
  assign n4728 = n4721 & ~n4727;
  assign n4729 = ~n4722 & ~n4727;
  assign n4730 = ~n4725 & n4729;
  assign n4731 = ~n4728 & ~n4730;
  assign n4732 = n4469 & ~n4731;
  assign n4733 = ~n4469 & n4731;
  assign n4734 = ~n4732 & ~n4733;
  assign n4735 = pi12  & pi34 ;
  assign n4736 = pi38  & pi39 ;
  assign n4737 = n521 & n4736;
  assign n4738 = pi7  & pi39 ;
  assign n4739 = pi8  & pi38 ;
  assign n4740 = ~n4738 & ~n4739;
  assign n4741 = n4735 & ~n4737;
  assign n4742 = ~n4740 & n4741;
  assign n4743 = n4735 & ~n4742;
  assign n4744 = ~n4737 & ~n4742;
  assign n4745 = ~n4740 & n4744;
  assign n4746 = ~n4743 & ~n4745;
  assign n4747 = ~n4734 & ~n4746;
  assign n4748 = n4734 & n4746;
  assign n4749 = ~n4747 & ~n4748;
  assign n4750 = ~n4720 & ~n4749;
  assign n4751 = n4720 & n4749;
  assign n4752 = ~n4750 & ~n4751;
  assign n4753 = ~n4678 & ~n4752;
  assign n4754 = n4678 & n4752;
  assign n4755 = ~n4753 & ~n4754;
  assign n4756 = ~n4677 & n4755;
  assign n4757 = n4677 & ~n4755;
  assign n4758 = ~n4756 & ~n4757;
  assign n4759 = ~n4550 & ~n4554;
  assign n4760 = ~n4511 & ~n4525;
  assign n4761 = n4759 & n4760;
  assign n4762 = ~n4759 & ~n4760;
  assign n4763 = ~n4761 & ~n4762;
  assign n4764 = ~n4454 & ~n4472;
  assign n4765 = ~n4763 & n4764;
  assign n4766 = n4763 & ~n4764;
  assign n4767 = ~n4765 & ~n4766;
  assign n4768 = ~n4429 & ~n4476;
  assign n4769 = n4495 & n4536;
  assign n4770 = ~n4495 & ~n4536;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = n4508 & ~n4771;
  assign n4773 = ~n4508 & n4771;
  assign n4774 = ~n4772 & ~n4773;
  assign n4775 = ~n4422 & ~n4425;
  assign n4776 = pi1  & pi45 ;
  assign n4777 = n1990 & n4776;
  assign n4778 = ~n1990 & ~n4776;
  assign n4779 = ~n4777 & ~n4778;
  assign n4780 = n4458 & n4779;
  assign n4781 = n4458 & ~n4780;
  assign n4782 = ~n4458 & n4779;
  assign n4783 = ~n4781 & ~n4782;
  assign n4784 = ~n4522 & ~n4783;
  assign n4785 = n4522 & n4783;
  assign n4786 = ~n4784 & ~n4785;
  assign n4787 = ~n4775 & n4786;
  assign n4788 = n4775 & ~n4786;
  assign n4789 = ~n4787 & ~n4788;
  assign n4790 = n4774 & n4789;
  assign n4791 = ~n4774 & ~n4789;
  assign n4792 = ~n4790 & ~n4791;
  assign n4793 = ~n4768 & n4792;
  assign n4794 = n4768 & ~n4792;
  assign n4795 = ~n4793 & ~n4794;
  assign n4796 = n4767 & n4795;
  assign n4797 = ~n4767 & ~n4795;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = n4758 & n4798;
  assign n4800 = ~n4758 & ~n4798;
  assign n4801 = ~n4799 & ~n4800;
  assign n4802 = ~n4675 & ~n4801;
  assign n4803 = n4675 & n4801;
  assign n4804 = ~n4802 & ~n4803;
  assign n4805 = ~n4609 & ~n4614;
  assign n4806 = ~n4804 & n4805;
  assign n4807 = n4804 & ~n4805;
  assign po47  = ~n4806 & ~n4807;
  assign n4809 = ~n4670 & ~n4674;
  assign n4810 = ~n4621 & ~n4667;
  assign n4811 = ~n4793 & ~n4796;
  assign n4812 = n4810 & n4811;
  assign n4813 = ~n4810 & ~n4811;
  assign n4814 = ~n4812 & ~n4813;
  assign n4815 = n4631 & n4714;
  assign n4816 = ~n4631 & ~n4714;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = n4686 & ~n4817;
  assign n4819 = ~n4686 & n4817;
  assign n4820 = ~n4818 & ~n4819;
  assign n4821 = ~n4702 & ~n4717;
  assign n4822 = ~n4820 & n4821;
  assign n4823 = n4820 & ~n4821;
  assign n4824 = ~n4822 & ~n4823;
  assign n4825 = ~n4646 & ~n4652;
  assign n4826 = ~n4824 & n4825;
  assign n4827 = n4824 & ~n4825;
  assign n4828 = ~n4826 & ~n4827;
  assign n4829 = ~n4720 & n4749;
  assign n4830 = ~n4753 & ~n4829;
  assign n4831 = ~n4662 & ~n4664;
  assign n4832 = ~n4830 & ~n4831;
  assign n4833 = ~n4830 & ~n4832;
  assign n4834 = ~n4831 & ~n4832;
  assign n4835 = ~n4833 & ~n4834;
  assign n4836 = n4828 & ~n4835;
  assign n4837 = ~n4828 & n4835;
  assign n4838 = ~n4836 & ~n4837;
  assign n4839 = n4814 & n4838;
  assign n4840 = n4814 & ~n4839;
  assign n4841 = n4838 & ~n4839;
  assign n4842 = ~n4840 & ~n4841;
  assign n4843 = ~n4756 & ~n4799;
  assign n4844 = ~n4780 & ~n4784;
  assign n4845 = pi13  & pi34 ;
  assign n4846 = pi12  & pi40 ;
  assign n4847 = n3887 & n4846;
  assign n4848 = pi7  & pi40 ;
  assign n4849 = pi12  & pi35 ;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = n4845 & ~n4847;
  assign n4852 = ~n4850 & n4851;
  assign n4853 = n4845 & ~n4852;
  assign n4854 = ~n4847 & ~n4852;
  assign n4855 = ~n4850 & n4854;
  assign n4856 = ~n4853 & ~n4855;
  assign n4857 = ~n4844 & ~n4856;
  assign n4858 = ~n4844 & ~n4857;
  assign n4859 = ~n4856 & ~n4857;
  assign n4860 = ~n4858 & ~n4859;
  assign n4861 = ~n4655 & ~n4658;
  assign n4862 = n4860 & n4861;
  assign n4863 = ~n4860 & ~n4861;
  assign n4864 = ~n4862 & ~n4863;
  assign n4865 = ~n4787 & ~n4790;
  assign n4866 = ~n4864 & n4865;
  assign n4867 = n4864 & ~n4865;
  assign n4868 = ~n4866 & ~n4867;
  assign n4869 = ~n4762 & ~n4766;
  assign n4870 = ~n4868 & n4869;
  assign n4871 = n4868 & ~n4869;
  assign n4872 = ~n4870 & ~n4871;
  assign n4873 = ~n4469 & ~n4731;
  assign n4874 = ~n4747 & ~n4873;
  assign n4875 = ~n4770 & ~n4773;
  assign n4876 = n4874 & n4875;
  assign n4877 = ~n4874 & ~n4875;
  assign n4878 = ~n4876 & ~n4877;
  assign n4879 = pi1  & pi46 ;
  assign n4880 = ~pi24  & ~n4879;
  assign n4881 = pi24  & pi46 ;
  assign n4882 = pi1  & n4881;
  assign n4883 = ~n4880 & ~n4882;
  assign n4884 = ~n4699 & n4883;
  assign n4885 = ~n4699 & ~n4884;
  assign n4886 = n4883 & ~n4884;
  assign n4887 = ~n4885 & ~n4886;
  assign n4888 = ~n4744 & ~n4887;
  assign n4889 = ~n4744 & ~n4888;
  assign n4890 = ~n4887 & ~n4888;
  assign n4891 = ~n4889 & ~n4890;
  assign n4892 = n4878 & ~n4891;
  assign n4893 = n4878 & ~n4892;
  assign n4894 = ~n4891 & ~n4892;
  assign n4895 = ~n4893 & ~n4894;
  assign n4896 = pi0  & pi47 ;
  assign n4897 = pi2  & pi45 ;
  assign n4898 = ~n4896 & ~n4897;
  assign n4899 = pi45  & pi47 ;
  assign n4900 = n196 & n4899;
  assign n4901 = n4777 & ~n4898;
  assign n4902 = ~n4900 & n4901;
  assign n4903 = ~n4900 & ~n4902;
  assign n4904 = ~n4898 & n4903;
  assign n4905 = n4777 & ~n4902;
  assign n4906 = ~n4904 & ~n4905;
  assign n4907 = pi16  & pi31 ;
  assign n4908 = pi29  & pi30 ;
  assign n4909 = n1199 & n4908;
  assign n4910 = pi17  & pi30 ;
  assign n4911 = pi18  & pi29 ;
  assign n4912 = ~n4910 & ~n4911;
  assign n4913 = n4907 & ~n4909;
  assign n4914 = ~n4912 & n4913;
  assign n4915 = n4907 & ~n4914;
  assign n4916 = ~n4909 & ~n4914;
  assign n4917 = ~n4912 & n4916;
  assign n4918 = ~n4915 & ~n4917;
  assign n4919 = ~n4906 & ~n4918;
  assign n4920 = ~n4906 & ~n4919;
  assign n4921 = ~n4918 & ~n4919;
  assign n4922 = ~n4920 & ~n4921;
  assign n4923 = pi19  & pi28 ;
  assign n4924 = n1593 & n2646;
  assign n4925 = pi20  & pi27 ;
  assign n4926 = ~n1965 & ~n4925;
  assign n4927 = n4923 & ~n4924;
  assign n4928 = ~n4926 & n4927;
  assign n4929 = n4923 & ~n4928;
  assign n4930 = ~n4924 & ~n4928;
  assign n4931 = ~n4926 & n4930;
  assign n4932 = ~n4929 & ~n4931;
  assign n4933 = ~n4922 & ~n4932;
  assign n4934 = ~n4922 & ~n4933;
  assign n4935 = ~n4932 & ~n4933;
  assign n4936 = ~n4934 & ~n4935;
  assign n4937 = n4643 & n4729;
  assign n4938 = ~n4643 & ~n4729;
  assign n4939 = ~n4937 & ~n4938;
  assign n4940 = pi3  & pi44 ;
  assign n4941 = pi32  & pi43 ;
  assign n4942 = n940 & n4941;
  assign n4943 = pi4  & pi43 ;
  assign n4944 = pi15  & pi32 ;
  assign n4945 = ~n4943 & ~n4944;
  assign n4946 = n4940 & ~n4942;
  assign n4947 = ~n4945 & n4946;
  assign n4948 = n4940 & ~n4947;
  assign n4949 = ~n4942 & ~n4947;
  assign n4950 = ~n4945 & n4949;
  assign n4951 = ~n4948 & ~n4950;
  assign n4952 = n4939 & ~n4951;
  assign n4953 = n4939 & ~n4952;
  assign n4954 = ~n4951 & ~n4952;
  assign n4955 = ~n4953 & ~n4954;
  assign n4956 = pi9  & pi38 ;
  assign n4957 = pi11  & pi36 ;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = n1012 & n3301;
  assign n4960 = pi8  & pi39 ;
  assign n4961 = ~n4958 & n4960;
  assign n4962 = ~n4959 & n4961;
  assign n4963 = ~n4959 & ~n4962;
  assign n4964 = ~n4958 & n4963;
  assign n4965 = n4960 & ~n4962;
  assign n4966 = ~n4964 & ~n4965;
  assign n4967 = pi10  & pi37 ;
  assign n4968 = n1789 & n1806;
  assign n4969 = pi22  & pi25 ;
  assign n4970 = ~n2110 & ~n4969;
  assign n4971 = n4967 & ~n4968;
  assign n4972 = ~n4970 & n4971;
  assign n4973 = n4967 & ~n4972;
  assign n4974 = ~n4968 & ~n4972;
  assign n4975 = ~n4970 & n4974;
  assign n4976 = ~n4973 & ~n4975;
  assign n4977 = ~n4966 & ~n4976;
  assign n4978 = ~n4966 & ~n4977;
  assign n4979 = ~n4976 & ~n4977;
  assign n4980 = ~n4978 & ~n4979;
  assign n4981 = pi5  & pi42 ;
  assign n4982 = pi33  & pi41 ;
  assign n4983 = n1044 & n4982;
  assign n4984 = pi6  & pi41 ;
  assign n4985 = pi14  & pi33 ;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = n4981 & ~n4983;
  assign n4988 = ~n4986 & n4987;
  assign n4989 = n4981 & ~n4988;
  assign n4990 = ~n4983 & ~n4988;
  assign n4991 = ~n4986 & n4990;
  assign n4992 = ~n4989 & ~n4991;
  assign n4993 = ~n4980 & ~n4992;
  assign n4994 = ~n4980 & ~n4993;
  assign n4995 = ~n4992 & ~n4993;
  assign n4996 = ~n4994 & ~n4995;
  assign n4997 = ~n4955 & n4996;
  assign n4998 = n4955 & ~n4996;
  assign n4999 = ~n4997 & ~n4998;
  assign n5000 = ~n4936 & ~n4999;
  assign n5001 = n4936 & n4999;
  assign n5002 = ~n5000 & ~n5001;
  assign n5003 = ~n4895 & n5002;
  assign n5004 = ~n4895 & ~n5003;
  assign n5005 = n5002 & ~n5003;
  assign n5006 = ~n5004 & ~n5005;
  assign n5007 = n4872 & ~n5006;
  assign n5008 = ~n4872 & n5006;
  assign n5009 = ~n5007 & ~n5008;
  assign n5010 = ~n4843 & n5009;
  assign n5011 = ~n4843 & ~n5010;
  assign n5012 = n5009 & ~n5010;
  assign n5013 = ~n5011 & ~n5012;
  assign n5014 = ~n4842 & ~n5013;
  assign n5015 = n4842 & n5013;
  assign n5016 = ~n5014 & ~n5015;
  assign n5017 = ~n4809 & n5016;
  assign n5018 = n4809 & ~n5016;
  assign n5019 = ~n5017 & ~n5018;
  assign n5020 = ~n4803 & ~n4807;
  assign n5021 = ~n5019 & n5020;
  assign n5022 = n5019 & ~n5020;
  assign po48  = ~n5021 & ~n5022;
  assign n5024 = ~n5010 & ~n5014;
  assign n5025 = ~n4813 & ~n4839;
  assign n5026 = ~n4832 & ~n4836;
  assign n5027 = ~n4867 & ~n4871;
  assign n5028 = pi6  & pi42 ;
  assign n5029 = pi13  & pi35 ;
  assign n5030 = ~n5028 & ~n5029;
  assign n5031 = n5028 & n5029;
  assign n5032 = pi14  & pi34 ;
  assign n5033 = ~n5030 & n5032;
  assign n5034 = ~n5031 & n5033;
  assign n5035 = ~n5031 & ~n5034;
  assign n5036 = ~n5030 & n5035;
  assign n5037 = n5032 & ~n5034;
  assign n5038 = ~n5036 & ~n5037;
  assign n5039 = pi7  & pi41 ;
  assign n5040 = n4284 & n4846;
  assign n5041 = pi12  & pi36 ;
  assign n5042 = pi8  & pi40 ;
  assign n5043 = ~n5041 & ~n5042;
  assign n5044 = n5039 & ~n5040;
  assign n5045 = ~n5043 & n5044;
  assign n5046 = n5039 & ~n5045;
  assign n5047 = ~n5040 & ~n5045;
  assign n5048 = ~n5043 & n5047;
  assign n5049 = ~n5046 & ~n5048;
  assign n5050 = ~n5038 & ~n5049;
  assign n5051 = ~n5038 & ~n5050;
  assign n5052 = ~n5049 & ~n5050;
  assign n5053 = ~n5051 & ~n5052;
  assign n5054 = pi9  & pi39 ;
  assign n5055 = pi37  & pi38 ;
  assign n5056 = n1111 & n5055;
  assign n5057 = pi10  & pi38 ;
  assign n5058 = ~n4258 & ~n5057;
  assign n5059 = n5054 & ~n5056;
  assign n5060 = ~n5058 & n5059;
  assign n5061 = n5054 & ~n5060;
  assign n5062 = ~n5056 & ~n5060;
  assign n5063 = ~n5058 & n5062;
  assign n5064 = ~n5061 & ~n5063;
  assign n5065 = ~n5053 & ~n5064;
  assign n5066 = ~n5053 & ~n5065;
  assign n5067 = ~n5064 & ~n5065;
  assign n5068 = ~n5066 & ~n5067;
  assign n5069 = ~n4857 & ~n4863;
  assign n5070 = n5068 & n5069;
  assign n5071 = ~n5068 & ~n5069;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = pi5  & pi43 ;
  assign n5074 = pi15  & pi33 ;
  assign n5075 = ~n5073 & ~n5074;
  assign n5076 = pi33  & pi43 ;
  assign n5077 = n1043 & n5076;
  assign n5078 = pi4  & pi44 ;
  assign n5079 = ~n5075 & n5078;
  assign n5080 = ~n5077 & n5079;
  assign n5081 = ~n5077 & ~n5080;
  assign n5082 = ~n5075 & n5081;
  assign n5083 = n5078 & ~n5080;
  assign n5084 = ~n5082 & ~n5083;
  assign n5085 = pi20  & pi28 ;
  assign n5086 = n1481 & n2646;
  assign n5087 = pi21  & pi27 ;
  assign n5088 = pi22  & pi26 ;
  assign n5089 = ~n5087 & ~n5088;
  assign n5090 = n5085 & ~n5086;
  assign n5091 = ~n5089 & n5090;
  assign n5092 = n5085 & ~n5091;
  assign n5093 = ~n5086 & ~n5091;
  assign n5094 = ~n5089 & n5093;
  assign n5095 = ~n5092 & ~n5094;
  assign n5096 = ~n5084 & ~n5095;
  assign n5097 = ~n5084 & ~n5096;
  assign n5098 = ~n5095 & ~n5096;
  assign n5099 = ~n5097 & ~n5098;
  assign n5100 = pi17  & pi31 ;
  assign n5101 = n1085 & n4908;
  assign n5102 = pi18  & pi30 ;
  assign n5103 = pi19  & pi29 ;
  assign n5104 = ~n5102 & ~n5103;
  assign n5105 = n5100 & ~n5101;
  assign n5106 = ~n5104 & n5105;
  assign n5107 = n5100 & ~n5106;
  assign n5108 = ~n5101 & ~n5106;
  assign n5109 = ~n5104 & n5108;
  assign n5110 = ~n5107 & ~n5109;
  assign n5111 = ~n5099 & ~n5110;
  assign n5112 = ~n5099 & ~n5111;
  assign n5113 = ~n5110 & ~n5111;
  assign n5114 = ~n5112 & ~n5113;
  assign n5115 = ~n5072 & n5114;
  assign n5116 = n5072 & ~n5114;
  assign n5117 = ~n5115 & ~n5116;
  assign n5118 = ~n5027 & n5117;
  assign n5119 = n5027 & ~n5117;
  assign n5120 = ~n5118 & ~n5119;
  assign n5121 = ~n5026 & n5120;
  assign n5122 = n5026 & ~n5120;
  assign n5123 = ~n5121 & ~n5122;
  assign n5124 = n5025 & ~n5123;
  assign n5125 = ~n5025 & n5123;
  assign n5126 = ~n5124 & ~n5125;
  assign n5127 = ~n5003 & ~n5007;
  assign n5128 = ~n4823 & ~n4827;
  assign n5129 = ~n4877 & ~n4892;
  assign n5130 = n5128 & n5129;
  assign n5131 = ~n5128 & ~n5129;
  assign n5132 = ~n5130 & ~n5131;
  assign n5133 = pi0  & pi48 ;
  assign n5134 = n4882 & n5133;
  assign n5135 = n4882 & ~n5134;
  assign n5136 = ~n4882 & n5133;
  assign n5137 = ~n5135 & ~n5136;
  assign n5138 = pi1  & pi47 ;
  assign n5139 = n1457 & n5138;
  assign n5140 = n5138 & ~n5139;
  assign n5141 = n1457 & ~n5139;
  assign n5142 = ~n5140 & ~n5141;
  assign n5143 = ~n5137 & ~n5142;
  assign n5144 = ~n5137 & ~n5143;
  assign n5145 = ~n5142 & ~n5143;
  assign n5146 = ~n5144 & ~n5145;
  assign n5147 = ~n4816 & ~n4819;
  assign n5148 = n5146 & n5147;
  assign n5149 = ~n5146 & ~n5147;
  assign n5150 = ~n5148 & ~n5149;
  assign n5151 = ~n4938 & ~n4952;
  assign n5152 = ~n5150 & n5151;
  assign n5153 = n5150 & ~n5151;
  assign n5154 = ~n5152 & ~n5153;
  assign n5155 = n5132 & n5154;
  assign n5156 = ~n5132 & ~n5154;
  assign n5157 = ~n5155 & ~n5156;
  assign n5158 = ~n5127 & n5157;
  assign n5159 = ~n5127 & ~n5158;
  assign n5160 = n5157 & ~n5158;
  assign n5161 = ~n5159 & ~n5160;
  assign n5162 = n4930 & n4963;
  assign n5163 = ~n4930 & ~n4963;
  assign n5164 = ~n5162 & ~n5163;
  assign n5165 = n4990 & ~n5164;
  assign n5166 = ~n4990 & n5164;
  assign n5167 = ~n5165 & ~n5166;
  assign n5168 = ~n4977 & ~n4993;
  assign n5169 = ~n5167 & n5168;
  assign n5170 = n5167 & ~n5168;
  assign n5171 = ~n5169 & ~n5170;
  assign n5172 = n4854 & n4974;
  assign n5173 = ~n4854 & ~n4974;
  assign n5174 = ~n5172 & ~n5173;
  assign n5175 = pi2  & pi46 ;
  assign n5176 = pi3  & pi45 ;
  assign n5177 = pi16  & pi32 ;
  assign n5178 = n5176 & n5177;
  assign n5179 = ~n5176 & ~n5177;
  assign n5180 = n5175 & ~n5178;
  assign n5181 = ~n5179 & n5180;
  assign n5182 = n5175 & ~n5181;
  assign n5183 = ~n5178 & ~n5181;
  assign n5184 = ~n5179 & n5183;
  assign n5185 = ~n5182 & ~n5184;
  assign n5186 = n5174 & ~n5185;
  assign n5187 = n5174 & ~n5186;
  assign n5188 = ~n5185 & ~n5186;
  assign n5189 = ~n5187 & ~n5188;
  assign n5190 = ~n5171 & n5189;
  assign n5191 = n5171 & ~n5189;
  assign n5192 = ~n5190 & ~n5191;
  assign n5193 = ~n4955 & ~n4996;
  assign n5194 = ~n5000 & ~n5193;
  assign n5195 = n5192 & ~n5194;
  assign n5196 = ~n5192 & n5194;
  assign n5197 = ~n5195 & ~n5196;
  assign n5198 = n4916 & n4949;
  assign n5199 = ~n4916 & ~n4949;
  assign n5200 = ~n5198 & ~n5199;
  assign n5201 = n4903 & ~n5200;
  assign n5202 = ~n4903 & n5200;
  assign n5203 = ~n5201 & ~n5202;
  assign n5204 = ~n4884 & ~n4888;
  assign n5205 = ~n4919 & ~n4933;
  assign n5206 = n5204 & n5205;
  assign n5207 = ~n5204 & ~n5205;
  assign n5208 = ~n5206 & ~n5207;
  assign n5209 = n5203 & n5208;
  assign n5210 = ~n5203 & ~n5208;
  assign n5211 = ~n5209 & ~n5210;
  assign n5212 = n5197 & n5211;
  assign n5213 = ~n5197 & ~n5211;
  assign n5214 = ~n5212 & ~n5213;
  assign n5215 = ~n5161 & n5214;
  assign n5216 = n5161 & ~n5214;
  assign n5217 = ~n5215 & ~n5216;
  assign n5218 = n5126 & n5217;
  assign n5219 = ~n5126 & ~n5217;
  assign n5220 = ~n5218 & ~n5219;
  assign n5221 = n5024 & ~n5220;
  assign n5222 = ~n5024 & n5220;
  assign n5223 = ~n5221 & ~n5222;
  assign n5224 = ~n5017 & ~n5022;
  assign n5225 = ~n5223 & n5224;
  assign n5226 = ~n5221 & ~n5224;
  assign n5227 = ~n5222 & n5226;
  assign po49  = ~n5225 & ~n5227;
  assign n5229 = ~n5158 & ~n5215;
  assign n5230 = ~n5195 & ~n5212;
  assign n5231 = ~n5131 & ~n5155;
  assign n5232 = pi7  & pi42 ;
  assign n5233 = pi8  & pi41 ;
  assign n5234 = ~n5232 & ~n5233;
  assign n5235 = pi41  & pi42 ;
  assign n5236 = n521 & n5235;
  assign n5237 = pi13  & pi36 ;
  assign n5238 = ~n5234 & n5237;
  assign n5239 = ~n5236 & n5238;
  assign n5240 = ~n5236 & ~n5239;
  assign n5241 = ~n5234 & n5240;
  assign n5242 = n5237 & ~n5239;
  assign n5243 = ~n5241 & ~n5242;
  assign n5244 = pi11  & pi38 ;
  assign n5245 = pi23  & pi26 ;
  assign n5246 = n1789 & n5245;
  assign n5247 = ~n1789 & ~n5245;
  assign n5248 = n5244 & ~n5246;
  assign n5249 = ~n5247 & n5248;
  assign n5250 = n5244 & ~n5249;
  assign n5251 = ~n5246 & ~n5249;
  assign n5252 = ~n5247 & n5251;
  assign n5253 = ~n5250 & ~n5252;
  assign n5254 = ~n5243 & ~n5253;
  assign n5255 = ~n5243 & ~n5254;
  assign n5256 = ~n5253 & ~n5254;
  assign n5257 = ~n5255 & ~n5256;
  assign n5258 = pi15  & pi34 ;
  assign n5259 = pi35  & pi43 ;
  assign n5260 = n1044 & n5259;
  assign n5261 = pi6  & pi43 ;
  assign n5262 = pi14  & pi35 ;
  assign n5263 = ~n5261 & ~n5262;
  assign n5264 = n5258 & ~n5260;
  assign n5265 = ~n5263 & n5264;
  assign n5266 = n5258 & ~n5265;
  assign n5267 = ~n5260 & ~n5265;
  assign n5268 = ~n5263 & n5267;
  assign n5269 = ~n5266 & ~n5268;
  assign n5270 = ~n5257 & ~n5269;
  assign n5271 = ~n5257 & ~n5270;
  assign n5272 = ~n5269 & ~n5270;
  assign n5273 = ~n5271 & ~n5272;
  assign n5274 = pi3  & pi46 ;
  assign n5275 = pi2  & pi47 ;
  assign n5276 = ~n5274 & ~n5275;
  assign n5277 = pi46  & pi47 ;
  assign n5278 = n218 & n5277;
  assign n5279 = pi22  & pi27 ;
  assign n5280 = ~n5276 & n5279;
  assign n5281 = ~n5278 & n5280;
  assign n5282 = ~n5278 & ~n5281;
  assign n5283 = ~n5276 & n5282;
  assign n5284 = n5279 & ~n5281;
  assign n5285 = ~n5283 & ~n5284;
  assign n5286 = pi19  & pi30 ;
  assign n5287 = n1593 & n2915;
  assign n5288 = pi20  & pi29 ;
  assign n5289 = pi21  & pi28 ;
  assign n5290 = ~n5288 & ~n5289;
  assign n5291 = n5286 & ~n5287;
  assign n5292 = ~n5290 & n5291;
  assign n5293 = n5286 & ~n5292;
  assign n5294 = ~n5287 & ~n5292;
  assign n5295 = ~n5290 & n5294;
  assign n5296 = ~n5293 & ~n5295;
  assign n5297 = ~n5285 & ~n5296;
  assign n5298 = ~n5285 & ~n5297;
  assign n5299 = ~n5296 & ~n5297;
  assign n5300 = ~n5298 & ~n5299;
  assign n5301 = pi9  & pi40 ;
  assign n5302 = pi37  & pi39 ;
  assign n5303 = n460 & n5302;
  assign n5304 = pi12  & pi37 ;
  assign n5305 = pi10  & pi39 ;
  assign n5306 = ~n5304 & ~n5305;
  assign n5307 = n5301 & ~n5303;
  assign n5308 = ~n5306 & n5307;
  assign n5309 = n5301 & ~n5308;
  assign n5310 = ~n5303 & ~n5308;
  assign n5311 = ~n5306 & n5310;
  assign n5312 = ~n5309 & ~n5311;
  assign n5313 = ~n5300 & ~n5312;
  assign n5314 = ~n5300 & ~n5313;
  assign n5315 = ~n5312 & ~n5313;
  assign n5316 = ~n5314 & ~n5315;
  assign n5317 = pi0  & pi49 ;
  assign n5318 = pi44  & pi45 ;
  assign n5319 = n226 & n5318;
  assign n5320 = pi4  & pi45 ;
  assign n5321 = pi5  & pi44 ;
  assign n5322 = ~n5320 & ~n5321;
  assign n5323 = n5317 & ~n5319;
  assign n5324 = ~n5322 & n5323;
  assign n5325 = n5317 & ~n5324;
  assign n5326 = ~n5319 & ~n5324;
  assign n5327 = ~n5322 & n5326;
  assign n5328 = ~n5325 & ~n5327;
  assign n5329 = ~n5134 & ~n5143;
  assign n5330 = ~n5328 & n5329;
  assign n5331 = n5328 & ~n5329;
  assign n5332 = ~n5330 & ~n5331;
  assign n5333 = pi16  & pi33 ;
  assign n5334 = n1199 & n3567;
  assign n5335 = pi17  & pi32 ;
  assign n5336 = pi18  & pi31 ;
  assign n5337 = ~n5335 & ~n5336;
  assign n5338 = n5333 & ~n5334;
  assign n5339 = ~n5337 & n5338;
  assign n5340 = n5333 & ~n5339;
  assign n5341 = ~n5334 & ~n5339;
  assign n5342 = ~n5337 & n5341;
  assign n5343 = ~n5340 & ~n5342;
  assign n5344 = ~n5332 & ~n5343;
  assign n5345 = n5332 & n5343;
  assign n5346 = ~n5344 & ~n5345;
  assign n5347 = n5316 & n5346;
  assign n5348 = ~n5316 & ~n5346;
  assign n5349 = ~n5347 & ~n5348;
  assign n5350 = ~n5273 & ~n5349;
  assign n5351 = n5273 & n5349;
  assign n5352 = ~n5350 & ~n5351;
  assign n5353 = ~n5231 & n5352;
  assign n5354 = n5231 & ~n5352;
  assign n5355 = ~n5353 & ~n5354;
  assign n5356 = ~n5230 & n5355;
  assign n5357 = n5230 & ~n5355;
  assign n5358 = ~n5356 & ~n5357;
  assign n5359 = ~n5229 & n5358;
  assign n5360 = n5229 & ~n5358;
  assign n5361 = ~n5359 & ~n5360;
  assign n5362 = ~n5118 & ~n5121;
  assign n5363 = ~n5163 & ~n5166;
  assign n5364 = ~n5173 & ~n5186;
  assign n5365 = n5363 & n5364;
  assign n5366 = ~n5363 & ~n5364;
  assign n5367 = ~n5365 & ~n5366;
  assign n5368 = ~n5199 & ~n5202;
  assign n5369 = ~n5367 & n5368;
  assign n5370 = n5367 & ~n5368;
  assign n5371 = ~n5369 & ~n5370;
  assign n5372 = ~n5170 & ~n5191;
  assign n5373 = ~n5207 & ~n5209;
  assign n5374 = ~n5372 & ~n5373;
  assign n5375 = ~n5372 & ~n5374;
  assign n5376 = ~n5373 & ~n5374;
  assign n5377 = ~n5375 & ~n5376;
  assign n5378 = ~n5371 & n5377;
  assign n5379 = n5371 & ~n5377;
  assign n5380 = ~n5378 & ~n5379;
  assign n5381 = ~n5362 & n5380;
  assign n5382 = ~n5362 & ~n5381;
  assign n5383 = n5380 & ~n5381;
  assign n5384 = ~n5382 & ~n5383;
  assign n5385 = n5035 & n5108;
  assign n5386 = ~n5035 & ~n5108;
  assign n5387 = ~n5385 & ~n5386;
  assign n5388 = n5047 & ~n5387;
  assign n5389 = ~n5047 & n5387;
  assign n5390 = ~n5388 & ~n5389;
  assign n5391 = ~n5096 & ~n5111;
  assign n5392 = ~n5390 & n5391;
  assign n5393 = n5390 & ~n5391;
  assign n5394 = ~n5392 & ~n5393;
  assign n5395 = ~n5149 & ~n5153;
  assign n5396 = ~n5394 & n5395;
  assign n5397 = n5394 & ~n5395;
  assign n5398 = ~n5396 & ~n5397;
  assign n5399 = ~n5071 & ~n5116;
  assign n5400 = n5398 & ~n5399;
  assign n5401 = ~n5398 & n5399;
  assign n5402 = ~n5400 & ~n5401;
  assign n5403 = n5081 & n5183;
  assign n5404 = ~n5081 & ~n5183;
  assign n5405 = ~n5403 & ~n5404;
  assign n5406 = n5093 & ~n5405;
  assign n5407 = ~n5093 & n5405;
  assign n5408 = ~n5406 & ~n5407;
  assign n5409 = ~n5050 & ~n5065;
  assign n5410 = pi48  & n1645;
  assign n5411 = pi1  & pi48 ;
  assign n5412 = ~pi25  & ~n5411;
  assign n5413 = ~n5410 & ~n5412;
  assign n5414 = n5139 & n5413;
  assign n5415 = ~n5139 & ~n5413;
  assign n5416 = ~n5414 & ~n5415;
  assign n5417 = ~n5062 & n5416;
  assign n5418 = n5062 & ~n5416;
  assign n5419 = ~n5417 & ~n5418;
  assign n5420 = ~n5409 & n5419;
  assign n5421 = n5409 & ~n5419;
  assign n5422 = ~n5420 & ~n5421;
  assign n5423 = n5408 & n5422;
  assign n5424 = ~n5408 & ~n5422;
  assign n5425 = ~n5423 & ~n5424;
  assign n5426 = n5402 & n5425;
  assign n5427 = ~n5402 & ~n5425;
  assign n5428 = ~n5426 & ~n5427;
  assign n5429 = ~n5384 & n5428;
  assign n5430 = n5384 & ~n5428;
  assign n5431 = ~n5429 & ~n5430;
  assign n5432 = n5361 & n5431;
  assign n5433 = ~n5361 & ~n5431;
  assign n5434 = ~n5432 & ~n5433;
  assign n5435 = ~n5125 & ~n5218;
  assign n5436 = ~n5434 & n5435;
  assign n5437 = n5434 & ~n5435;
  assign n5438 = ~n5436 & ~n5437;
  assign n5439 = ~n5222 & ~n5226;
  assign n5440 = ~n5438 & n5439;
  assign n5441 = n5438 & ~n5439;
  assign po50  = ~n5440 & ~n5441;
  assign n5443 = ~n5359 & ~n5432;
  assign n5444 = ~n5381 & ~n5429;
  assign n5445 = ~n5400 & ~n5426;
  assign n5446 = ~n5374 & ~n5379;
  assign n5447 = pi5  & pi45 ;
  assign n5448 = pi15  & pi35 ;
  assign n5449 = ~n5447 & ~n5448;
  assign n5450 = pi35  & pi45 ;
  assign n5451 = n1043 & n5450;
  assign n5452 = pi16  & pi34 ;
  assign n5453 = ~n5449 & n5452;
  assign n5454 = ~n5451 & n5453;
  assign n5455 = ~n5451 & ~n5454;
  assign n5456 = ~n5449 & n5455;
  assign n5457 = n5452 & ~n5454;
  assign n5458 = ~n5456 & ~n5457;
  assign n5459 = pi22  & pi28 ;
  assign n5460 = pi18  & pi32 ;
  assign n5461 = pi23  & pi27 ;
  assign n5462 = n5460 & n5461;
  assign n5463 = ~n5460 & ~n5461;
  assign n5464 = n5459 & ~n5462;
  assign n5465 = ~n5463 & n5464;
  assign n5466 = n5459 & ~n5465;
  assign n5467 = ~n5462 & ~n5465;
  assign n5468 = ~n5463 & n5467;
  assign n5469 = ~n5466 & ~n5468;
  assign n5470 = ~n5458 & ~n5469;
  assign n5471 = ~n5458 & ~n5470;
  assign n5472 = ~n5469 & ~n5470;
  assign n5473 = ~n5471 & ~n5472;
  assign n5474 = ~n5414 & ~n5417;
  assign n5475 = n5473 & n5474;
  assign n5476 = ~n5473 & ~n5474;
  assign n5477 = ~n5475 & ~n5476;
  assign n5478 = pi0  & pi50 ;
  assign n5479 = pi2  & pi48 ;
  assign n5480 = ~n5478 & ~n5479;
  assign n5481 = pi48  & pi50 ;
  assign n5482 = n196 & n5481;
  assign n5483 = n5410 & ~n5480;
  assign n5484 = ~n5482 & n5483;
  assign n5485 = ~n5482 & ~n5484;
  assign n5486 = ~n5480 & n5485;
  assign n5487 = n5410 & ~n5484;
  assign n5488 = ~n5486 & ~n5487;
  assign n5489 = pi3  & pi47 ;
  assign n5490 = pi33  & pi46 ;
  assign n5491 = n1109 & n5490;
  assign n5492 = pi4  & pi46 ;
  assign n5493 = pi17  & pi33 ;
  assign n5494 = ~n5492 & ~n5493;
  assign n5495 = n5489 & ~n5491;
  assign n5496 = ~n5494 & n5495;
  assign n5497 = n5489 & ~n5496;
  assign n5498 = ~n5491 & ~n5496;
  assign n5499 = ~n5494 & n5498;
  assign n5500 = ~n5497 & ~n5499;
  assign n5501 = ~n5488 & ~n5500;
  assign n5502 = ~n5488 & ~n5501;
  assign n5503 = ~n5500 & ~n5501;
  assign n5504 = ~n5502 & ~n5503;
  assign n5505 = pi19  & pi31 ;
  assign n5506 = n1593 & n4908;
  assign n5507 = pi20  & pi30 ;
  assign n5508 = pi21  & pi29 ;
  assign n5509 = ~n5507 & ~n5508;
  assign n5510 = n5505 & ~n5506;
  assign n5511 = ~n5509 & n5510;
  assign n5512 = n5505 & ~n5511;
  assign n5513 = ~n5506 & ~n5511;
  assign n5514 = ~n5509 & n5513;
  assign n5515 = ~n5512 & ~n5514;
  assign n5516 = ~n5504 & ~n5515;
  assign n5517 = ~n5504 & ~n5516;
  assign n5518 = ~n5515 & ~n5516;
  assign n5519 = ~n5517 & ~n5518;
  assign n5520 = pi7  & pi43 ;
  assign n5521 = pi14  & pi36 ;
  assign n5522 = ~n5520 & ~n5521;
  assign n5523 = n5520 & n5521;
  assign n5524 = pi6  & pi44 ;
  assign n5525 = ~n5522 & n5524;
  assign n5526 = ~n5523 & n5525;
  assign n5527 = ~n5523 & ~n5526;
  assign n5528 = ~n5522 & n5527;
  assign n5529 = n5524 & ~n5526;
  assign n5530 = ~n5528 & ~n5529;
  assign n5531 = pi8  & pi42 ;
  assign n5532 = pi37  & pi41 ;
  assign n5533 = n506 & n5532;
  assign n5534 = pi13  & pi37 ;
  assign n5535 = pi9  & pi41 ;
  assign n5536 = ~n5534 & ~n5535;
  assign n5537 = n5531 & ~n5533;
  assign n5538 = ~n5536 & n5537;
  assign n5539 = n5531 & ~n5538;
  assign n5540 = ~n5533 & ~n5538;
  assign n5541 = ~n5536 & n5540;
  assign n5542 = ~n5539 & ~n5541;
  assign n5543 = ~n5530 & ~n5542;
  assign n5544 = ~n5530 & ~n5543;
  assign n5545 = ~n5542 & ~n5543;
  assign n5546 = ~n5544 & ~n5545;
  assign n5547 = pi12  & pi38 ;
  assign n5548 = pi39  & pi40 ;
  assign n5549 = n1111 & n5548;
  assign n5550 = pi11  & pi39 ;
  assign n5551 = pi10  & pi40 ;
  assign n5552 = ~n5550 & ~n5551;
  assign n5553 = n5547 & ~n5549;
  assign n5554 = ~n5552 & n5553;
  assign n5555 = n5547 & ~n5554;
  assign n5556 = ~n5549 & ~n5554;
  assign n5557 = ~n5552 & n5556;
  assign n5558 = ~n5555 & ~n5557;
  assign n5559 = ~n5546 & ~n5558;
  assign n5560 = ~n5546 & ~n5559;
  assign n5561 = ~n5558 & ~n5559;
  assign n5562 = ~n5560 & ~n5561;
  assign n5563 = ~n5519 & n5562;
  assign n5564 = n5519 & ~n5562;
  assign n5565 = ~n5563 & ~n5564;
  assign n5566 = n5477 & ~n5565;
  assign n5567 = ~n5477 & n5565;
  assign n5568 = ~n5566 & ~n5567;
  assign n5569 = ~n5446 & n5568;
  assign n5570 = ~n5446 & ~n5569;
  assign n5571 = n5568 & ~n5569;
  assign n5572 = ~n5570 & ~n5571;
  assign n5573 = ~n5445 & ~n5572;
  assign n5574 = n5445 & n5572;
  assign n5575 = ~n5573 & ~n5574;
  assign n5576 = ~n5444 & n5575;
  assign n5577 = n5444 & ~n5575;
  assign n5578 = ~n5576 & ~n5577;
  assign n5579 = ~n5353 & ~n5356;
  assign n5580 = ~n5393 & ~n5397;
  assign n5581 = ~n5420 & ~n5423;
  assign n5582 = n5580 & n5581;
  assign n5583 = ~n5580 & ~n5581;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = ~n5386 & ~n5389;
  assign n5586 = ~n5404 & ~n5407;
  assign n5587 = n5585 & n5586;
  assign n5588 = ~n5585 & ~n5586;
  assign n5589 = ~n5587 & ~n5588;
  assign n5590 = n5282 & n5326;
  assign n5591 = ~n5282 & ~n5326;
  assign n5592 = ~n5590 & ~n5591;
  assign n5593 = n5267 & ~n5592;
  assign n5594 = ~n5267 & n5592;
  assign n5595 = ~n5593 & ~n5594;
  assign n5596 = n5589 & n5595;
  assign n5597 = ~n5589 & ~n5595;
  assign n5598 = ~n5596 & ~n5597;
  assign n5599 = n5584 & n5598;
  assign n5600 = ~n5584 & ~n5598;
  assign n5601 = ~n5599 & ~n5600;
  assign n5602 = n5579 & ~n5601;
  assign n5603 = ~n5579 & n5601;
  assign n5604 = ~n5602 & ~n5603;
  assign n5605 = ~n5297 & ~n5313;
  assign n5606 = ~n5328 & ~n5329;
  assign n5607 = ~n5344 & ~n5606;
  assign n5608 = n5605 & n5607;
  assign n5609 = ~n5605 & ~n5607;
  assign n5610 = ~n5608 & ~n5609;
  assign n5611 = pi1  & pi49 ;
  assign n5612 = n2167 & n5611;
  assign n5613 = ~n2167 & ~n5611;
  assign n5614 = ~n5612 & ~n5613;
  assign n5615 = n5251 & ~n5614;
  assign n5616 = ~n5251 & n5614;
  assign n5617 = ~n5615 & ~n5616;
  assign n5618 = ~n5310 & n5617;
  assign n5619 = n5310 & ~n5617;
  assign n5620 = ~n5618 & ~n5619;
  assign n5621 = n5610 & n5620;
  assign n5622 = ~n5610 & ~n5620;
  assign n5623 = ~n5621 & ~n5622;
  assign n5624 = n5294 & n5341;
  assign n5625 = ~n5294 & ~n5341;
  assign n5626 = ~n5624 & ~n5625;
  assign n5627 = n5240 & ~n5626;
  assign n5628 = ~n5240 & n5626;
  assign n5629 = ~n5627 & ~n5628;
  assign n5630 = ~n5254 & ~n5270;
  assign n5631 = ~n5629 & n5630;
  assign n5632 = n5629 & ~n5630;
  assign n5633 = ~n5631 & ~n5632;
  assign n5634 = ~n5366 & ~n5370;
  assign n5635 = ~n5633 & n5634;
  assign n5636 = n5633 & ~n5634;
  assign n5637 = ~n5635 & ~n5636;
  assign n5638 = ~n5316 & n5346;
  assign n5639 = ~n5350 & ~n5638;
  assign n5640 = n5637 & ~n5639;
  assign n5641 = ~n5637 & n5639;
  assign n5642 = ~n5640 & ~n5641;
  assign n5643 = n5623 & n5642;
  assign n5644 = ~n5623 & ~n5642;
  assign n5645 = ~n5643 & ~n5644;
  assign n5646 = n5604 & n5645;
  assign n5647 = ~n5604 & ~n5645;
  assign n5648 = ~n5646 & ~n5647;
  assign n5649 = n5578 & n5648;
  assign n5650 = ~n5578 & ~n5648;
  assign n5651 = ~n5649 & ~n5650;
  assign n5652 = n5443 & ~n5651;
  assign n5653 = ~n5443 & n5651;
  assign n5654 = ~n5652 & ~n5653;
  assign n5655 = ~n5437 & ~n5441;
  assign n5656 = ~n5654 & n5655;
  assign n5657 = ~n5652 & ~n5655;
  assign n5658 = ~n5653 & n5657;
  assign po51  = ~n5656 & ~n5658;
  assign n5660 = ~n5653 & ~n5657;
  assign n5661 = ~n5576 & ~n5649;
  assign n5662 = ~n5603 & ~n5646;
  assign n5663 = ~n5640 & ~n5643;
  assign n5664 = ~n5583 & ~n5599;
  assign n5665 = pi0  & pi51 ;
  assign n5666 = n5612 & n5665;
  assign n5667 = n5612 & ~n5666;
  assign n5668 = ~n5612 & n5665;
  assign n5669 = ~n5667 & ~n5668;
  assign n5670 = pi1  & pi50 ;
  assign n5671 = pi26  & n5670;
  assign n5672 = pi26  & ~n5671;
  assign n5673 = n5670 & ~n5671;
  assign n5674 = ~n5672 & ~n5673;
  assign n5675 = ~n5669 & ~n5674;
  assign n5676 = ~n5669 & ~n5675;
  assign n5677 = ~n5674 & ~n5675;
  assign n5678 = ~n5676 & ~n5677;
  assign n5679 = pi17  & pi34 ;
  assign n5680 = pi20  & pi31 ;
  assign n5681 = pi19  & pi32 ;
  assign n5682 = ~n5680 & ~n5681;
  assign n5683 = n1407 & n3567;
  assign n5684 = n5679 & ~n5682;
  assign n5685 = ~n5683 & n5684;
  assign n5686 = n5679 & ~n5685;
  assign n5687 = ~n5683 & ~n5685;
  assign n5688 = ~n5682 & n5687;
  assign n5689 = ~n5686 & ~n5688;
  assign n5690 = ~n5678 & ~n5689;
  assign n5691 = ~n5678 & ~n5690;
  assign n5692 = ~n5689 & ~n5690;
  assign n5693 = ~n5691 & ~n5692;
  assign n5694 = ~n5625 & ~n5628;
  assign n5695 = n5693 & n5694;
  assign n5696 = ~n5693 & ~n5694;
  assign n5697 = ~n5695 & ~n5696;
  assign n5698 = pi5  & pi46 ;
  assign n5699 = pi16  & pi35 ;
  assign n5700 = ~n5698 & ~n5699;
  assign n5701 = n5698 & n5699;
  assign n5702 = pi18  & pi33 ;
  assign n5703 = ~n5700 & n5702;
  assign n5704 = ~n5701 & n5703;
  assign n5705 = ~n5701 & ~n5704;
  assign n5706 = ~n5700 & n5705;
  assign n5707 = n5702 & ~n5704;
  assign n5708 = ~n5706 & ~n5707;
  assign n5709 = pi21  & pi30 ;
  assign n5710 = n1806 & n2915;
  assign n5711 = pi22  & pi29 ;
  assign n5712 = pi23  & pi28 ;
  assign n5713 = ~n5711 & ~n5712;
  assign n5714 = n5709 & ~n5710;
  assign n5715 = ~n5713 & n5714;
  assign n5716 = n5709 & ~n5715;
  assign n5717 = ~n5710 & ~n5715;
  assign n5718 = ~n5713 & n5717;
  assign n5719 = ~n5716 & ~n5718;
  assign n5720 = ~n5708 & ~n5719;
  assign n5721 = ~n5708 & ~n5720;
  assign n5722 = ~n5719 & ~n5720;
  assign n5723 = ~n5721 & ~n5722;
  assign n5724 = pi15  & pi36 ;
  assign n5725 = pi37  & pi45 ;
  assign n5726 = n1044 & n5725;
  assign n5727 = pi6  & pi45 ;
  assign n5728 = pi14  & pi37 ;
  assign n5729 = ~n5727 & ~n5728;
  assign n5730 = n5724 & ~n5726;
  assign n5731 = ~n5729 & n5730;
  assign n5732 = n5724 & ~n5731;
  assign n5733 = ~n5726 & ~n5731;
  assign n5734 = ~n5729 & n5733;
  assign n5735 = ~n5732 & ~n5734;
  assign n5736 = ~n5723 & ~n5735;
  assign n5737 = ~n5723 & ~n5736;
  assign n5738 = ~n5735 & ~n5736;
  assign n5739 = ~n5737 & ~n5738;
  assign n5740 = pi8  & pi43 ;
  assign n5741 = pi13  & pi38 ;
  assign n5742 = ~n5740 & ~n5741;
  assign n5743 = pi13  & pi43 ;
  assign n5744 = n4739 & n5743;
  assign n5745 = pi7  & pi44 ;
  assign n5746 = ~n5742 & n5745;
  assign n5747 = ~n5744 & n5746;
  assign n5748 = ~n5744 & ~n5747;
  assign n5749 = ~n5742 & n5748;
  assign n5750 = n5745 & ~n5747;
  assign n5751 = ~n5749 & ~n5750;
  assign n5752 = pi9  & pi42 ;
  assign n5753 = n460 & n3729;
  assign n5754 = pi12  & pi39 ;
  assign n5755 = pi10  & pi41 ;
  assign n5756 = ~n5754 & ~n5755;
  assign n5757 = n5752 & ~n5753;
  assign n5758 = ~n5756 & n5757;
  assign n5759 = n5752 & ~n5758;
  assign n5760 = ~n5753 & ~n5758;
  assign n5761 = ~n5756 & n5760;
  assign n5762 = ~n5759 & ~n5761;
  assign n5763 = ~n5751 & ~n5762;
  assign n5764 = ~n5751 & ~n5763;
  assign n5765 = ~n5762 & ~n5763;
  assign n5766 = ~n5764 & ~n5765;
  assign n5767 = pi11  & pi40 ;
  assign n5768 = n1789 & n2646;
  assign n5769 = pi24  & pi27 ;
  assign n5770 = ~n2310 & ~n5769;
  assign n5771 = n5767 & ~n5768;
  assign n5772 = ~n5770 & n5771;
  assign n5773 = n5767 & ~n5772;
  assign n5774 = ~n5768 & ~n5772;
  assign n5775 = ~n5770 & n5774;
  assign n5776 = ~n5773 & ~n5775;
  assign n5777 = ~n5766 & ~n5776;
  assign n5778 = ~n5766 & ~n5777;
  assign n5779 = ~n5776 & ~n5777;
  assign n5780 = ~n5778 & ~n5779;
  assign n5781 = ~n5739 & n5780;
  assign n5782 = n5739 & ~n5780;
  assign n5783 = ~n5781 & ~n5782;
  assign n5784 = n5697 & ~n5783;
  assign n5785 = ~n5697 & n5783;
  assign n5786 = ~n5784 & ~n5785;
  assign n5787 = ~n5664 & n5786;
  assign n5788 = n5664 & ~n5786;
  assign n5789 = ~n5787 & ~n5788;
  assign n5790 = ~n5663 & n5789;
  assign n5791 = n5663 & ~n5789;
  assign n5792 = ~n5790 & ~n5791;
  assign n5793 = ~n5662 & n5792;
  assign n5794 = n5662 & ~n5792;
  assign n5795 = ~n5793 & ~n5794;
  assign n5796 = ~n5569 & ~n5573;
  assign n5797 = ~n5632 & ~n5636;
  assign n5798 = ~n5609 & ~n5621;
  assign n5799 = n5797 & n5798;
  assign n5800 = ~n5797 & ~n5798;
  assign n5801 = ~n5799 & ~n5800;
  assign n5802 = ~n5591 & ~n5594;
  assign n5803 = ~n5616 & ~n5618;
  assign n5804 = n5802 & n5803;
  assign n5805 = ~n5802 & ~n5803;
  assign n5806 = ~n5804 & ~n5805;
  assign n5807 = ~n5501 & ~n5516;
  assign n5808 = ~n5806 & n5807;
  assign n5809 = n5806 & ~n5807;
  assign n5810 = ~n5808 & ~n5809;
  assign n5811 = n5801 & n5810;
  assign n5812 = ~n5801 & ~n5810;
  assign n5813 = ~n5811 & ~n5812;
  assign n5814 = ~n5796 & n5813;
  assign n5815 = n5796 & ~n5813;
  assign n5816 = ~n5814 & ~n5815;
  assign n5817 = ~n5519 & ~n5562;
  assign n5818 = ~n5566 & ~n5817;
  assign n5819 = n5455 & n5556;
  assign n5820 = ~n5455 & ~n5556;
  assign n5821 = ~n5819 & ~n5820;
  assign n5822 = pi2  & pi49 ;
  assign n5823 = pi47  & pi48 ;
  assign n5824 = n209 & n5823;
  assign n5825 = pi3  & pi48 ;
  assign n5826 = pi4  & pi47 ;
  assign n5827 = ~n5825 & ~n5826;
  assign n5828 = n5822 & ~n5824;
  assign n5829 = ~n5827 & n5828;
  assign n5830 = n5822 & ~n5829;
  assign n5831 = ~n5824 & ~n5829;
  assign n5832 = ~n5827 & n5831;
  assign n5833 = ~n5830 & ~n5832;
  assign n5834 = n5821 & ~n5833;
  assign n5835 = n5821 & ~n5834;
  assign n5836 = ~n5833 & ~n5834;
  assign n5837 = ~n5835 & ~n5836;
  assign n5838 = ~n5470 & ~n5476;
  assign n5839 = n5837 & n5838;
  assign n5840 = ~n5837 & ~n5838;
  assign n5841 = ~n5839 & ~n5840;
  assign n5842 = ~n5588 & ~n5596;
  assign n5843 = n5841 & ~n5842;
  assign n5844 = ~n5841 & n5842;
  assign n5845 = ~n5843 & ~n5844;
  assign n5846 = ~n5818 & n5845;
  assign n5847 = n5818 & ~n5845;
  assign n5848 = ~n5846 & ~n5847;
  assign n5849 = n5527 & n5540;
  assign n5850 = ~n5527 & ~n5540;
  assign n5851 = ~n5849 & ~n5850;
  assign n5852 = n5467 & ~n5851;
  assign n5853 = ~n5467 & n5851;
  assign n5854 = ~n5852 & ~n5853;
  assign n5855 = ~n5543 & ~n5559;
  assign n5856 = ~n5854 & n5855;
  assign n5857 = n5854 & ~n5855;
  assign n5858 = ~n5856 & ~n5857;
  assign n5859 = n5498 & n5513;
  assign n5860 = ~n5498 & ~n5513;
  assign n5861 = ~n5859 & ~n5860;
  assign n5862 = n5485 & ~n5861;
  assign n5863 = ~n5485 & n5861;
  assign n5864 = ~n5862 & ~n5863;
  assign n5865 = n5858 & n5864;
  assign n5866 = ~n5858 & ~n5864;
  assign n5867 = ~n5865 & ~n5866;
  assign n5868 = n5848 & n5867;
  assign n5869 = ~n5848 & ~n5867;
  assign n5870 = ~n5868 & ~n5869;
  assign n5871 = n5816 & n5870;
  assign n5872 = ~n5816 & ~n5870;
  assign n5873 = ~n5871 & ~n5872;
  assign n5874 = n5795 & n5873;
  assign n5875 = ~n5795 & ~n5873;
  assign n5876 = ~n5874 & ~n5875;
  assign n5877 = ~n5661 & n5876;
  assign n5878 = n5661 & ~n5876;
  assign n5879 = ~n5877 & ~n5878;
  assign n5880 = ~n5660 & ~n5879;
  assign n5881 = n5660 & n5879;
  assign po52  = n5880 | n5881;
  assign n5883 = ~n5660 & ~n5878;
  assign n5884 = ~n5877 & ~n5883;
  assign n5885 = ~n5793 & ~n5874;
  assign n5886 = ~n5787 & ~n5790;
  assign n5887 = ~n5860 & ~n5863;
  assign n5888 = pi19  & pi33 ;
  assign n5889 = pi49  & pi50 ;
  assign n5890 = n218 & n5889;
  assign n5891 = pi2  & pi50 ;
  assign n5892 = pi3  & pi49 ;
  assign n5893 = ~n5891 & ~n5892;
  assign n5894 = n5888 & ~n5890;
  assign n5895 = ~n5893 & n5894;
  assign n5896 = n5888 & ~n5895;
  assign n5897 = ~n5890 & ~n5895;
  assign n5898 = ~n5893 & n5897;
  assign n5899 = ~n5896 & ~n5898;
  assign n5900 = ~n5887 & ~n5899;
  assign n5901 = ~n5887 & ~n5900;
  assign n5902 = ~n5899 & ~n5900;
  assign n5903 = ~n5901 & ~n5902;
  assign n5904 = ~n5850 & ~n5853;
  assign n5905 = n5903 & n5904;
  assign n5906 = ~n5903 & ~n5904;
  assign n5907 = ~n5905 & ~n5906;
  assign n5908 = ~n5840 & ~n5843;
  assign n5909 = ~n5907 & n5908;
  assign n5910 = n5907 & ~n5908;
  assign n5911 = ~n5909 & ~n5910;
  assign n5912 = ~n5763 & ~n5777;
  assign n5913 = ~n5820 & ~n5834;
  assign n5914 = pi1  & pi51 ;
  assign n5915 = ~n2468 & ~n5914;
  assign n5916 = n2468 & n5914;
  assign n5917 = ~n5915 & ~n5916;
  assign n5918 = n5671 & n5917;
  assign n5919 = ~n5671 & ~n5917;
  assign n5920 = ~n5918 & ~n5919;
  assign n5921 = ~n5774 & n5920;
  assign n5922 = n5774 & ~n5920;
  assign n5923 = ~n5921 & ~n5922;
  assign n5924 = ~n5913 & n5923;
  assign n5925 = n5913 & ~n5923;
  assign n5926 = ~n5924 & ~n5925;
  assign n5927 = ~n5912 & n5926;
  assign n5928 = n5912 & ~n5926;
  assign n5929 = ~n5927 & ~n5928;
  assign n5930 = n5911 & n5929;
  assign n5931 = ~n5911 & ~n5929;
  assign n5932 = ~n5930 & ~n5931;
  assign n5933 = n5886 & ~n5932;
  assign n5934 = ~n5886 & n5932;
  assign n5935 = ~n5933 & ~n5934;
  assign n5936 = ~n5666 & ~n5675;
  assign n5937 = n5760 & n5936;
  assign n5938 = ~n5760 & ~n5936;
  assign n5939 = ~n5937 & ~n5938;
  assign n5940 = pi0  & pi52 ;
  assign n5941 = pi4  & pi48 ;
  assign n5942 = pi17  & pi35 ;
  assign n5943 = n5941 & n5942;
  assign n5944 = ~n5941 & ~n5942;
  assign n5945 = n5940 & ~n5943;
  assign n5946 = ~n5944 & n5945;
  assign n5947 = n5940 & ~n5946;
  assign n5948 = ~n5943 & ~n5946;
  assign n5949 = ~n5944 & n5948;
  assign n5950 = ~n5947 & ~n5949;
  assign n5951 = n5939 & ~n5950;
  assign n5952 = n5939 & ~n5951;
  assign n5953 = ~n5950 & ~n5951;
  assign n5954 = ~n5952 & ~n5953;
  assign n5955 = ~n5690 & ~n5696;
  assign n5956 = n5954 & n5955;
  assign n5957 = ~n5954 & ~n5955;
  assign n5958 = ~n5956 & ~n5957;
  assign n5959 = ~n5805 & ~n5809;
  assign n5960 = ~n5958 & n5959;
  assign n5961 = n5958 & ~n5959;
  assign n5962 = ~n5960 & ~n5961;
  assign n5963 = ~n5739 & ~n5780;
  assign n5964 = ~n5784 & ~n5963;
  assign n5965 = n5705 & n5748;
  assign n5966 = ~n5705 & ~n5748;
  assign n5967 = ~n5965 & ~n5966;
  assign n5968 = n5717 & ~n5967;
  assign n5969 = ~n5717 & n5967;
  assign n5970 = ~n5968 & ~n5969;
  assign n5971 = n5687 & n5831;
  assign n5972 = ~n5687 & ~n5831;
  assign n5973 = ~n5971 & ~n5972;
  assign n5974 = n5733 & ~n5973;
  assign n5975 = ~n5733 & n5973;
  assign n5976 = ~n5974 & ~n5975;
  assign n5977 = ~n5720 & ~n5736;
  assign n5978 = ~n5976 & n5977;
  assign n5979 = n5976 & ~n5977;
  assign n5980 = ~n5978 & ~n5979;
  assign n5981 = n5970 & n5980;
  assign n5982 = ~n5970 & ~n5980;
  assign n5983 = ~n5981 & ~n5982;
  assign n5984 = ~n5964 & n5983;
  assign n5985 = ~n5964 & ~n5984;
  assign n5986 = n5983 & ~n5984;
  assign n5987 = ~n5985 & ~n5986;
  assign n5988 = n5962 & ~n5987;
  assign n5989 = n5962 & ~n5988;
  assign n5990 = ~n5987 & ~n5988;
  assign n5991 = ~n5989 & ~n5990;
  assign n5992 = n5935 & ~n5991;
  assign n5993 = n5935 & ~n5992;
  assign n5994 = ~n5991 & ~n5992;
  assign n5995 = ~n5993 & ~n5994;
  assign n5996 = ~n5846 & ~n5868;
  assign n5997 = ~n5800 & ~n5811;
  assign n5998 = ~n5857 & ~n5865;
  assign n5999 = pi16  & pi36 ;
  assign n6000 = pi6  & pi46 ;
  assign n6001 = ~n5999 & ~n6000;
  assign n6002 = pi36  & pi46 ;
  assign n6003 = n685 & n6002;
  assign n6004 = pi5  & pi47 ;
  assign n6005 = ~n6001 & n6004;
  assign n6006 = ~n6003 & n6005;
  assign n6007 = ~n6003 & ~n6006;
  assign n6008 = ~n6001 & n6007;
  assign n6009 = n6004 & ~n6006;
  assign n6010 = ~n6008 & ~n6009;
  assign n6011 = pi10  & pi42 ;
  assign n6012 = pi40  & pi41 ;
  assign n6013 = n579 & n6012;
  assign n6014 = pi11  & pi41 ;
  assign n6015 = ~n4846 & ~n6014;
  assign n6016 = n6011 & ~n6013;
  assign n6017 = ~n6015 & n6016;
  assign n6018 = n6011 & ~n6017;
  assign n6019 = ~n6013 & ~n6017;
  assign n6020 = ~n6015 & n6019;
  assign n6021 = ~n6018 & ~n6020;
  assign n6022 = ~n6010 & ~n6021;
  assign n6023 = ~n6010 & ~n6022;
  assign n6024 = ~n6021 & ~n6022;
  assign n6025 = ~n6023 & ~n6024;
  assign n6026 = pi15  & pi37 ;
  assign n6027 = n521 & n5318;
  assign n6028 = pi7  & pi45 ;
  assign n6029 = pi8  & pi44 ;
  assign n6030 = ~n6028 & ~n6029;
  assign n6031 = n6026 & ~n6027;
  assign n6032 = ~n6030 & n6031;
  assign n6033 = n6026 & ~n6032;
  assign n6034 = ~n6027 & ~n6032;
  assign n6035 = ~n6030 & n6034;
  assign n6036 = ~n6033 & ~n6035;
  assign n6037 = ~n6025 & ~n6036;
  assign n6038 = ~n6025 & ~n6037;
  assign n6039 = ~n6036 & ~n6037;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = pi20  & pi32 ;
  assign n6042 = pi21  & pi31 ;
  assign n6043 = ~n6041 & ~n6042;
  assign n6044 = n1593 & n3567;
  assign n6045 = pi18  & pi34 ;
  assign n6046 = ~n6043 & n6045;
  assign n6047 = ~n6044 & n6046;
  assign n6048 = ~n6044 & ~n6047;
  assign n6049 = ~n6043 & n6048;
  assign n6050 = n6045 & ~n6047;
  assign n6051 = ~n6049 & ~n6050;
  assign n6052 = pi22  & pi30 ;
  assign n6053 = n2110 & n2915;
  assign n6054 = pi23  & pi29 ;
  assign n6055 = pi24  & pi28 ;
  assign n6056 = ~n6054 & ~n6055;
  assign n6057 = n6052 & ~n6053;
  assign n6058 = ~n6056 & n6057;
  assign n6059 = n6052 & ~n6058;
  assign n6060 = ~n6053 & ~n6058;
  assign n6061 = ~n6056 & n6060;
  assign n6062 = ~n6059 & ~n6061;
  assign n6063 = ~n6051 & ~n6062;
  assign n6064 = ~n6051 & ~n6063;
  assign n6065 = ~n6062 & ~n6063;
  assign n6066 = ~n6064 & ~n6065;
  assign n6067 = n5054 & n5743;
  assign n6068 = pi9  & pi43 ;
  assign n6069 = pi13  & pi39 ;
  assign n6070 = ~n6068 & ~n6069;
  assign n6071 = n3944 & ~n6067;
  assign n6072 = ~n6070 & n6071;
  assign n6073 = n3944 & ~n6072;
  assign n6074 = ~n6067 & ~n6072;
  assign n6075 = ~n6070 & n6074;
  assign n6076 = ~n6073 & ~n6075;
  assign n6077 = ~n6066 & ~n6076;
  assign n6078 = ~n6066 & ~n6077;
  assign n6079 = ~n6076 & ~n6077;
  assign n6080 = ~n6078 & ~n6079;
  assign n6081 = n6040 & n6080;
  assign n6082 = ~n6040 & ~n6080;
  assign n6083 = ~n6081 & ~n6082;
  assign n6084 = ~n5998 & n6083;
  assign n6085 = n5998 & ~n6083;
  assign n6086 = ~n6084 & ~n6085;
  assign n6087 = ~n5997 & n6086;
  assign n6088 = n5997 & ~n6086;
  assign n6089 = ~n6087 & ~n6088;
  assign n6090 = n5996 & ~n6089;
  assign n6091 = ~n5996 & n6089;
  assign n6092 = ~n6090 & ~n6091;
  assign n6093 = ~n5814 & ~n5871;
  assign n6094 = n6092 & ~n6093;
  assign n6095 = ~n6092 & n6093;
  assign n6096 = ~n6094 & ~n6095;
  assign n6097 = ~n5995 & n6096;
  assign n6098 = n5995 & ~n6096;
  assign n6099 = ~n6097 & ~n6098;
  assign n6100 = n5885 & ~n6099;
  assign n6101 = ~n5885 & n6099;
  assign n6102 = ~n6100 & ~n6101;
  assign n6103 = n5884 & ~n6102;
  assign n6104 = ~n5884 & ~n6100;
  assign n6105 = ~n6101 & n6104;
  assign po53  = ~n6103 & ~n6105;
  assign n6107 = ~n6101 & ~n6104;
  assign n6108 = ~n6094 & ~n6097;
  assign n6109 = ~n5934 & ~n5992;
  assign n6110 = ~n5984 & ~n5988;
  assign n6111 = pi2  & pi51 ;
  assign n6112 = pi3  & pi50 ;
  assign n6113 = ~n6111 & ~n6112;
  assign n6114 = pi50  & pi51 ;
  assign n6115 = n218 & n6114;
  assign n6116 = n5916 & ~n6113;
  assign n6117 = ~n6115 & n6116;
  assign n6118 = ~n6115 & ~n6117;
  assign n6119 = ~n6113 & n6118;
  assign n6120 = n5916 & ~n6117;
  assign n6121 = ~n6119 & ~n6120;
  assign n6122 = pi4  & pi49 ;
  assign n6123 = n1199 & n4691;
  assign n6124 = pi17  & pi36 ;
  assign n6125 = pi18  & pi35 ;
  assign n6126 = ~n6124 & ~n6125;
  assign n6127 = n6122 & ~n6123;
  assign n6128 = ~n6126 & n6127;
  assign n6129 = n6122 & ~n6128;
  assign n6130 = ~n6123 & ~n6128;
  assign n6131 = ~n6126 & n6130;
  assign n6132 = ~n6129 & ~n6131;
  assign n6133 = ~n6121 & ~n6132;
  assign n6134 = ~n6121 & ~n6133;
  assign n6135 = ~n6132 & ~n6133;
  assign n6136 = ~n6134 & ~n6135;
  assign n6137 = pi19  & pi34 ;
  assign n6138 = pi32  & pi33 ;
  assign n6139 = n1593 & n6138;
  assign n6140 = pi20  & pi33 ;
  assign n6141 = pi21  & pi32 ;
  assign n6142 = ~n6140 & ~n6141;
  assign n6143 = n6137 & ~n6139;
  assign n6144 = ~n6142 & n6143;
  assign n6145 = n6137 & ~n6144;
  assign n6146 = ~n6139 & ~n6144;
  assign n6147 = ~n6142 & n6146;
  assign n6148 = ~n6145 & ~n6147;
  assign n6149 = ~n6136 & ~n6148;
  assign n6150 = ~n6136 & ~n6149;
  assign n6151 = ~n6148 & ~n6149;
  assign n6152 = ~n6150 & ~n6151;
  assign n6153 = ~n5900 & ~n5906;
  assign n6154 = n6152 & n6153;
  assign n6155 = ~n6152 & ~n6153;
  assign n6156 = ~n6154 & ~n6155;
  assign n6157 = pi15  & pi38 ;
  assign n6158 = pi7  & pi46 ;
  assign n6159 = ~n6157 & ~n6158;
  assign n6160 = n6157 & n6158;
  assign n6161 = pi6  & pi47 ;
  assign n6162 = ~n6159 & n6161;
  assign n6163 = ~n6160 & n6162;
  assign n6164 = ~n6160 & ~n6163;
  assign n6165 = ~n6159 & n6164;
  assign n6166 = n6161 & ~n6163;
  assign n6167 = ~n6165 & ~n6166;
  assign n6168 = pi14  & pi39 ;
  assign n6169 = pi9  & pi44 ;
  assign n6170 = ~n6168 & ~n6169;
  assign n6171 = pi14  & pi44 ;
  assign n6172 = n5054 & n6171;
  assign n6173 = pi8  & pi45 ;
  assign n6174 = ~n6170 & n6173;
  assign n6175 = ~n6172 & n6174;
  assign n6176 = ~n6172 & ~n6175;
  assign n6177 = ~n6170 & n6176;
  assign n6178 = n6173 & ~n6175;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = ~n6167 & ~n6179;
  assign n6181 = ~n6167 & ~n6180;
  assign n6182 = ~n6179 & ~n6180;
  assign n6183 = ~n6181 & ~n6182;
  assign n6184 = pi0  & pi53 ;
  assign n6185 = pi16  & pi48 ;
  assign n6186 = n3982 & n6185;
  assign n6187 = pi5  & pi48 ;
  assign n6188 = pi16  & pi37 ;
  assign n6189 = ~n6187 & ~n6188;
  assign n6190 = n6184 & ~n6186;
  assign n6191 = ~n6189 & n6190;
  assign n6192 = n6184 & ~n6191;
  assign n6193 = ~n6186 & ~n6191;
  assign n6194 = ~n6189 & n6193;
  assign n6195 = ~n6192 & ~n6194;
  assign n6196 = ~n6183 & ~n6195;
  assign n6197 = ~n6183 & ~n6196;
  assign n6198 = ~n6195 & ~n6196;
  assign n6199 = ~n6197 & ~n6198;
  assign n6200 = ~n6156 & n6199;
  assign n6201 = n6156 & ~n6199;
  assign n6202 = ~n6200 & ~n6201;
  assign n6203 = pi10  & pi43 ;
  assign n6204 = pi12  & pi41 ;
  assign n6205 = ~n6203 & ~n6204;
  assign n6206 = n460 & n4490;
  assign n6207 = pi13  & pi40 ;
  assign n6208 = ~n6205 & n6207;
  assign n6209 = ~n6206 & n6208;
  assign n6210 = ~n6206 & ~n6209;
  assign n6211 = ~n6205 & n6210;
  assign n6212 = n6207 & ~n6209;
  assign n6213 = ~n6211 & ~n6212;
  assign n6214 = n2110 & n4908;
  assign n6215 = pi23  & pi30 ;
  assign n6216 = pi24  & pi29 ;
  assign n6217 = ~n6215 & ~n6216;
  assign n6218 = n2209 & ~n6214;
  assign n6219 = ~n6217 & n6218;
  assign n6220 = n2209 & ~n6219;
  assign n6221 = ~n6214 & ~n6219;
  assign n6222 = ~n6217 & n6221;
  assign n6223 = ~n6220 & ~n6222;
  assign n6224 = ~n6213 & ~n6223;
  assign n6225 = ~n6213 & ~n6224;
  assign n6226 = ~n6223 & ~n6224;
  assign n6227 = ~n6225 & ~n6226;
  assign n6228 = pi11  & pi42 ;
  assign n6229 = n2191 & n2310;
  assign n6230 = pi25  & pi28 ;
  assign n6231 = ~n2646 & ~n6230;
  assign n6232 = n6228 & ~n6229;
  assign n6233 = ~n6231 & n6232;
  assign n6234 = n6228 & ~n6233;
  assign n6235 = ~n6229 & ~n6233;
  assign n6236 = ~n6231 & n6235;
  assign n6237 = ~n6234 & ~n6236;
  assign n6238 = ~n6227 & ~n6237;
  assign n6239 = ~n6227 & ~n6238;
  assign n6240 = ~n6237 & ~n6238;
  assign n6241 = ~n6239 & ~n6240;
  assign n6242 = ~n5924 & ~n5927;
  assign n6243 = n6241 & n6242;
  assign n6244 = ~n6241 & ~n6242;
  assign n6245 = ~n6243 & ~n6244;
  assign n6246 = ~n5979 & ~n5981;
  assign n6247 = n6245 & ~n6246;
  assign n6248 = ~n6245 & n6246;
  assign n6249 = ~n6247 & ~n6248;
  assign n6250 = n6202 & n6249;
  assign n6251 = ~n6202 & ~n6249;
  assign n6252 = ~n6250 & ~n6251;
  assign n6253 = ~n6110 & n6252;
  assign n6254 = n6110 & ~n6252;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~n6109 & n6255;
  assign n6257 = n6109 & ~n6255;
  assign n6258 = ~n6256 & ~n6257;
  assign n6259 = n5897 & n5948;
  assign n6260 = ~n5897 & ~n5948;
  assign n6261 = ~n6259 & ~n6260;
  assign n6262 = n6060 & ~n6261;
  assign n6263 = ~n6060 & n6261;
  assign n6264 = ~n6262 & ~n6263;
  assign n6265 = ~n6063 & ~n6077;
  assign n6266 = ~n5938 & ~n5951;
  assign n6267 = n6265 & n6266;
  assign n6268 = ~n6265 & ~n6266;
  assign n6269 = ~n6267 & ~n6268;
  assign n6270 = n6264 & n6269;
  assign n6271 = ~n6264 & ~n6269;
  assign n6272 = ~n6270 & ~n6271;
  assign n6273 = n6007 & n6048;
  assign n6274 = ~n6007 & ~n6048;
  assign n6275 = ~n6273 & ~n6274;
  assign n6276 = n6034 & ~n6275;
  assign n6277 = ~n6034 & n6275;
  assign n6278 = ~n6276 & ~n6277;
  assign n6279 = ~n6022 & ~n6037;
  assign n6280 = pi52  & n1826;
  assign n6281 = pi1  & pi52 ;
  assign n6282 = ~pi27  & ~n6281;
  assign n6283 = ~n6280 & ~n6282;
  assign n6284 = n6019 & ~n6283;
  assign n6285 = ~n6019 & n6283;
  assign n6286 = ~n6284 & ~n6285;
  assign n6287 = ~n6074 & n6286;
  assign n6288 = n6074 & ~n6286;
  assign n6289 = ~n6287 & ~n6288;
  assign n6290 = ~n6279 & n6289;
  assign n6291 = ~n6279 & ~n6290;
  assign n6292 = n6289 & ~n6290;
  assign n6293 = ~n6291 & ~n6292;
  assign n6294 = n6278 & ~n6293;
  assign n6295 = n6278 & ~n6294;
  assign n6296 = ~n6293 & ~n6294;
  assign n6297 = ~n6295 & ~n6296;
  assign n6298 = n6272 & ~n6297;
  assign n6299 = n6272 & ~n6298;
  assign n6300 = ~n6297 & ~n6298;
  assign n6301 = ~n6299 & ~n6300;
  assign n6302 = ~n5910 & ~n5930;
  assign n6303 = n6301 & n6302;
  assign n6304 = ~n6301 & ~n6302;
  assign n6305 = ~n6303 & ~n6304;
  assign n6306 = ~n6082 & ~n6084;
  assign n6307 = ~n5966 & ~n5969;
  assign n6308 = ~n5918 & ~n5921;
  assign n6309 = n6307 & n6308;
  assign n6310 = ~n6307 & ~n6308;
  assign n6311 = ~n6309 & ~n6310;
  assign n6312 = ~n5972 & ~n5975;
  assign n6313 = ~n6311 & n6312;
  assign n6314 = n6311 & ~n6312;
  assign n6315 = ~n6313 & ~n6314;
  assign n6316 = ~n5957 & ~n5961;
  assign n6317 = ~n6315 & n6316;
  assign n6318 = n6315 & ~n6316;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = ~n6306 & n6319;
  assign n6321 = n6306 & ~n6319;
  assign n6322 = ~n6320 & ~n6321;
  assign n6323 = ~n6087 & ~n6091;
  assign n6324 = ~n6322 & n6323;
  assign n6325 = n6322 & ~n6323;
  assign n6326 = ~n6324 & ~n6325;
  assign n6327 = n6305 & n6326;
  assign n6328 = ~n6305 & ~n6326;
  assign n6329 = ~n6327 & ~n6328;
  assign n6330 = n6258 & n6329;
  assign n6331 = ~n6258 & ~n6329;
  assign n6332 = ~n6330 & ~n6331;
  assign n6333 = ~n6108 & n6332;
  assign n6334 = n6108 & ~n6332;
  assign n6335 = ~n6333 & ~n6334;
  assign n6336 = ~n6107 & ~n6335;
  assign n6337 = n6107 & n6335;
  assign po54  = n6336 | n6337;
  assign n6339 = ~n6256 & ~n6330;
  assign n6340 = ~n6298 & ~n6304;
  assign n6341 = ~n6318 & ~n6320;
  assign n6342 = n6340 & n6341;
  assign n6343 = ~n6340 & ~n6341;
  assign n6344 = ~n6342 & ~n6343;
  assign n6345 = ~n6290 & ~n6294;
  assign n6346 = ~n6268 & ~n6270;
  assign n6347 = pi0  & pi54 ;
  assign n6348 = n6280 & n6347;
  assign n6349 = n6280 & ~n6348;
  assign n6350 = ~n6280 & n6347;
  assign n6351 = ~n6349 & ~n6350;
  assign n6352 = pi1  & pi53 ;
  assign n6353 = n3742 & n6352;
  assign n6354 = n6352 & ~n6353;
  assign n6355 = n3742 & ~n6353;
  assign n6356 = ~n6354 & ~n6355;
  assign n6357 = ~n6351 & ~n6356;
  assign n6358 = ~n6351 & ~n6357;
  assign n6359 = ~n6356 & ~n6357;
  assign n6360 = ~n6358 & ~n6359;
  assign n6361 = pi21  & pi33 ;
  assign n6362 = pi22  & pi32 ;
  assign n6363 = ~n6361 & ~n6362;
  assign n6364 = n1481 & n6138;
  assign n6365 = pi19  & pi35 ;
  assign n6366 = ~n6363 & n6365;
  assign n6367 = ~n6364 & n6366;
  assign n6368 = ~n6364 & ~n6367;
  assign n6369 = ~n6363 & n6368;
  assign n6370 = n6365 & ~n6367;
  assign n6371 = ~n6369 & ~n6370;
  assign n6372 = pi23  & pi31 ;
  assign n6373 = n1789 & n4908;
  assign n6374 = pi24  & pi30 ;
  assign n6375 = pi25  & pi29 ;
  assign n6376 = ~n6374 & ~n6375;
  assign n6377 = n6372 & ~n6373;
  assign n6378 = ~n6376 & n6377;
  assign n6379 = n6372 & ~n6378;
  assign n6380 = ~n6373 & ~n6378;
  assign n6381 = ~n6376 & n6380;
  assign n6382 = ~n6379 & ~n6381;
  assign n6383 = ~n6371 & ~n6382;
  assign n6384 = ~n6371 & ~n6383;
  assign n6385 = ~n6382 & ~n6383;
  assign n6386 = ~n6384 & ~n6385;
  assign n6387 = ~n6360 & n6386;
  assign n6388 = n6360 & ~n6386;
  assign n6389 = ~n6387 & ~n6388;
  assign n6390 = ~n6346 & ~n6389;
  assign n6391 = ~n6346 & ~n6390;
  assign n6392 = ~n6389 & ~n6390;
  assign n6393 = ~n6391 & ~n6392;
  assign n6394 = ~n6345 & ~n6393;
  assign n6395 = ~n6345 & ~n6394;
  assign n6396 = ~n6393 & ~n6394;
  assign n6397 = ~n6395 & ~n6396;
  assign n6398 = n6344 & ~n6397;
  assign n6399 = n6344 & ~n6398;
  assign n6400 = ~n6397 & ~n6398;
  assign n6401 = ~n6399 & ~n6400;
  assign n6402 = ~n6325 & ~n6327;
  assign n6403 = ~n6401 & ~n6402;
  assign n6404 = ~n6401 & ~n6403;
  assign n6405 = ~n6402 & ~n6403;
  assign n6406 = ~n6404 & ~n6405;
  assign n6407 = ~n6250 & ~n6253;
  assign n6408 = ~n6274 & ~n6277;
  assign n6409 = ~n6260 & ~n6263;
  assign n6410 = n6408 & n6409;
  assign n6411 = ~n6408 & ~n6409;
  assign n6412 = ~n6410 & ~n6411;
  assign n6413 = ~n6285 & ~n6287;
  assign n6414 = ~n6412 & n6413;
  assign n6415 = n6412 & ~n6413;
  assign n6416 = ~n6414 & ~n6415;
  assign n6417 = ~n6155 & ~n6201;
  assign n6418 = n6416 & ~n6417;
  assign n6419 = ~n6416 & n6417;
  assign n6420 = ~n6418 & ~n6419;
  assign n6421 = n6164 & n6193;
  assign n6422 = ~n6164 & ~n6193;
  assign n6423 = ~n6421 & ~n6422;
  assign n6424 = n6235 & ~n6423;
  assign n6425 = ~n6235 & n6423;
  assign n6426 = ~n6424 & ~n6425;
  assign n6427 = n6130 & n6146;
  assign n6428 = ~n6130 & ~n6146;
  assign n6429 = ~n6427 & ~n6428;
  assign n6430 = n6221 & ~n6429;
  assign n6431 = ~n6221 & n6429;
  assign n6432 = ~n6430 & ~n6431;
  assign n6433 = ~n6180 & ~n6196;
  assign n6434 = ~n6432 & n6433;
  assign n6435 = n6432 & ~n6433;
  assign n6436 = ~n6434 & ~n6435;
  assign n6437 = n6426 & n6436;
  assign n6438 = ~n6426 & ~n6436;
  assign n6439 = ~n6437 & ~n6438;
  assign n6440 = n6420 & n6439;
  assign n6441 = ~n6420 & ~n6439;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = n6407 & ~n6442;
  assign n6444 = ~n6407 & n6442;
  assign n6445 = ~n6443 & ~n6444;
  assign n6446 = pi5  & pi49 ;
  assign n6447 = pi18  & pi36 ;
  assign n6448 = ~n6446 & ~n6447;
  assign n6449 = n6446 & n6447;
  assign n6450 = pi20  & pi34 ;
  assign n6451 = ~n6448 & n6450;
  assign n6452 = ~n6449 & n6451;
  assign n6453 = ~n6449 & ~n6452;
  assign n6454 = ~n6448 & n6453;
  assign n6455 = n6450 & ~n6452;
  assign n6456 = ~n6454 & ~n6455;
  assign n6457 = pi13  & pi41 ;
  assign n6458 = pi42  & pi43 ;
  assign n6459 = n579 & n6458;
  assign n6460 = pi11  & pi43 ;
  assign n6461 = pi12  & pi42 ;
  assign n6462 = ~n6460 & ~n6461;
  assign n6463 = n6457 & ~n6459;
  assign n6464 = ~n6462 & n6463;
  assign n6465 = n6457 & ~n6464;
  assign n6466 = ~n6459 & ~n6464;
  assign n6467 = ~n6462 & n6466;
  assign n6468 = ~n6465 & ~n6467;
  assign n6469 = ~n6456 & ~n6468;
  assign n6470 = ~n6456 & ~n6469;
  assign n6471 = ~n6468 & ~n6469;
  assign n6472 = ~n6470 & ~n6471;
  assign n6473 = pi17  & pi37 ;
  assign n6474 = pi38  & pi48 ;
  assign n6475 = n685 & n6474;
  assign n6476 = pi6  & pi48 ;
  assign n6477 = pi16  & pi38 ;
  assign n6478 = ~n6476 & ~n6477;
  assign n6479 = n6473 & ~n6475;
  assign n6480 = ~n6478 & n6479;
  assign n6481 = n6473 & ~n6480;
  assign n6482 = ~n6475 & ~n6480;
  assign n6483 = ~n6478 & n6482;
  assign n6484 = ~n6481 & ~n6483;
  assign n6485 = ~n6472 & ~n6484;
  assign n6486 = ~n6472 & ~n6485;
  assign n6487 = ~n6484 & ~n6485;
  assign n6488 = ~n6486 & ~n6487;
  assign n6489 = ~n6310 & ~n6314;
  assign n6490 = n6488 & n6489;
  assign n6491 = ~n6488 & ~n6489;
  assign n6492 = ~n6490 & ~n6491;
  assign n6493 = pi3  & pi51 ;
  assign n6494 = pi4  & pi50 ;
  assign n6495 = ~n6493 & ~n6494;
  assign n6496 = n209 & n6114;
  assign n6497 = pi2  & pi52 ;
  assign n6498 = ~n6495 & n6497;
  assign n6499 = ~n6496 & n6498;
  assign n6500 = ~n6496 & ~n6499;
  assign n6501 = ~n6495 & n6500;
  assign n6502 = n6497 & ~n6499;
  assign n6503 = ~n6501 & ~n6502;
  assign n6504 = pi7  & pi47 ;
  assign n6505 = pi15  & pi39 ;
  assign n6506 = pi8  & pi46 ;
  assign n6507 = n6505 & n6506;
  assign n6508 = ~n6505 & ~n6506;
  assign n6509 = n6504 & ~n6507;
  assign n6510 = ~n6508 & n6509;
  assign n6511 = n6504 & ~n6510;
  assign n6512 = ~n6507 & ~n6510;
  assign n6513 = ~n6508 & n6512;
  assign n6514 = ~n6511 & ~n6513;
  assign n6515 = ~n6503 & ~n6514;
  assign n6516 = ~n6503 & ~n6515;
  assign n6517 = ~n6514 & ~n6515;
  assign n6518 = ~n6516 & ~n6517;
  assign n6519 = pi9  & pi45 ;
  assign n6520 = n5551 & n6171;
  assign n6521 = pi14  & pi40 ;
  assign n6522 = pi10  & pi44 ;
  assign n6523 = ~n6521 & ~n6522;
  assign n6524 = n6519 & ~n6520;
  assign n6525 = ~n6523 & n6524;
  assign n6526 = n6519 & ~n6525;
  assign n6527 = ~n6520 & ~n6525;
  assign n6528 = ~n6523 & n6527;
  assign n6529 = ~n6526 & ~n6528;
  assign n6530 = ~n6518 & ~n6529;
  assign n6531 = ~n6518 & ~n6530;
  assign n6532 = ~n6529 & ~n6530;
  assign n6533 = ~n6531 & ~n6532;
  assign n6534 = ~n6492 & n6533;
  assign n6535 = n6492 & ~n6533;
  assign n6536 = ~n6534 & ~n6535;
  assign n6537 = ~n6244 & ~n6247;
  assign n6538 = n6118 & n6176;
  assign n6539 = ~n6118 & ~n6176;
  assign n6540 = ~n6538 & ~n6539;
  assign n6541 = n6210 & ~n6540;
  assign n6542 = ~n6210 & n6540;
  assign n6543 = ~n6541 & ~n6542;
  assign n6544 = ~n6224 & ~n6238;
  assign n6545 = ~n6133 & ~n6149;
  assign n6546 = n6544 & n6545;
  assign n6547 = ~n6544 & ~n6545;
  assign n6548 = ~n6546 & ~n6547;
  assign n6549 = n6543 & n6548;
  assign n6550 = ~n6543 & ~n6548;
  assign n6551 = ~n6549 & ~n6550;
  assign n6552 = ~n6537 & n6551;
  assign n6553 = ~n6537 & ~n6552;
  assign n6554 = n6551 & ~n6552;
  assign n6555 = ~n6553 & ~n6554;
  assign n6556 = n6536 & ~n6555;
  assign n6557 = n6536 & ~n6556;
  assign n6558 = ~n6555 & ~n6556;
  assign n6559 = ~n6557 & ~n6558;
  assign n6560 = n6445 & ~n6559;
  assign n6561 = n6445 & ~n6560;
  assign n6562 = ~n6559 & ~n6560;
  assign n6563 = ~n6561 & ~n6562;
  assign n6564 = ~n6406 & n6563;
  assign n6565 = n6406 & ~n6563;
  assign n6566 = ~n6564 & ~n6565;
  assign n6567 = ~n6339 & ~n6566;
  assign n6568 = n6339 & n6566;
  assign n6569 = ~n6567 & ~n6568;
  assign n6570 = ~n6107 & ~n6334;
  assign n6571 = ~n6333 & ~n6570;
  assign n6572 = ~n6569 & n6571;
  assign n6573 = n6569 & ~n6571;
  assign po55  = ~n6572 & ~n6573;
  assign n6575 = ~n6406 & ~n6563;
  assign n6576 = ~n6403 & ~n6575;
  assign n6577 = ~n6444 & ~n6560;
  assign n6578 = ~n6552 & ~n6556;
  assign n6579 = ~n6418 & ~n6440;
  assign n6580 = ~n6435 & ~n6437;
  assign n6581 = pi6  & pi49 ;
  assign n6582 = pi17  & pi38 ;
  assign n6583 = ~n6581 & ~n6582;
  assign n6584 = pi17  & pi49 ;
  assign n6585 = n4257 & n6584;
  assign n6586 = pi3  & pi52 ;
  assign n6587 = ~n6583 & n6586;
  assign n6588 = ~n6585 & n6587;
  assign n6589 = ~n6585 & ~n6588;
  assign n6590 = ~n6583 & n6589;
  assign n6591 = n6586 & ~n6588;
  assign n6592 = ~n6590 & ~n6591;
  assign n6593 = pi15  & pi40 ;
  assign n6594 = pi9  & pi46 ;
  assign n6595 = pi14  & pi41 ;
  assign n6596 = n6594 & n6595;
  assign n6597 = ~n6594 & ~n6595;
  assign n6598 = n6593 & ~n6596;
  assign n6599 = ~n6597 & n6598;
  assign n6600 = n6593 & ~n6599;
  assign n6601 = ~n6596 & ~n6599;
  assign n6602 = ~n6597 & n6601;
  assign n6603 = ~n6600 & ~n6602;
  assign n6604 = ~n6592 & ~n6603;
  assign n6605 = ~n6592 & ~n6604;
  assign n6606 = ~n6603 & ~n6604;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = ~n6428 & ~n6431;
  assign n6609 = n6607 & n6608;
  assign n6610 = ~n6607 & ~n6608;
  assign n6611 = ~n6609 & ~n6610;
  assign n6612 = ~n6547 & ~n6549;
  assign n6613 = n6611 & ~n6612;
  assign n6614 = ~n6611 & n6612;
  assign n6615 = ~n6613 & ~n6614;
  assign n6616 = ~n6580 & n6615;
  assign n6617 = n6580 & ~n6615;
  assign n6618 = ~n6616 & ~n6617;
  assign n6619 = ~n6579 & n6618;
  assign n6620 = ~n6579 & ~n6619;
  assign n6621 = n6618 & ~n6619;
  assign n6622 = ~n6620 & ~n6621;
  assign n6623 = ~n6578 & ~n6622;
  assign n6624 = ~n6578 & ~n6623;
  assign n6625 = ~n6622 & ~n6623;
  assign n6626 = ~n6624 & ~n6625;
  assign n6627 = ~n6577 & ~n6626;
  assign n6628 = ~n6577 & ~n6627;
  assign n6629 = ~n6626 & ~n6627;
  assign n6630 = ~n6628 & ~n6629;
  assign n6631 = ~n6422 & ~n6425;
  assign n6632 = ~n6539 & ~n6542;
  assign n6633 = n6631 & n6632;
  assign n6634 = ~n6631 & ~n6632;
  assign n6635 = ~n6633 & ~n6634;
  assign n6636 = pi28  & pi54 ;
  assign n6637 = pi1  & n6636;
  assign n6638 = pi1  & pi54 ;
  assign n6639 = ~pi28  & ~n6638;
  assign n6640 = ~n6637 & ~n6639;
  assign n6641 = n6353 & n6640;
  assign n6642 = n6353 & ~n6641;
  assign n6643 = n6640 & ~n6641;
  assign n6644 = ~n6642 & ~n6643;
  assign n6645 = ~n6466 & ~n6644;
  assign n6646 = ~n6466 & ~n6645;
  assign n6647 = ~n6644 & ~n6645;
  assign n6648 = ~n6646 & ~n6647;
  assign n6649 = n6635 & ~n6648;
  assign n6650 = n6635 & ~n6649;
  assign n6651 = ~n6648 & ~n6649;
  assign n6652 = ~n6650 & ~n6651;
  assign n6653 = ~n6491 & ~n6535;
  assign n6654 = ~n6652 & ~n6653;
  assign n6655 = ~n6652 & ~n6654;
  assign n6656 = ~n6653 & ~n6654;
  assign n6657 = ~n6655 & ~n6656;
  assign n6658 = ~n6348 & ~n6357;
  assign n6659 = n6512 & n6658;
  assign n6660 = ~n6512 & ~n6658;
  assign n6661 = ~n6659 & ~n6660;
  assign n6662 = pi5  & pi50 ;
  assign n6663 = n1085 & n4500;
  assign n6664 = pi18  & pi37 ;
  assign n6665 = pi19  & pi36 ;
  assign n6666 = ~n6664 & ~n6665;
  assign n6667 = n6662 & ~n6663;
  assign n6668 = ~n6666 & n6667;
  assign n6669 = n6662 & ~n6668;
  assign n6670 = ~n6663 & ~n6668;
  assign n6671 = ~n6666 & n6670;
  assign n6672 = ~n6669 & ~n6671;
  assign n6673 = n6661 & ~n6672;
  assign n6674 = n6661 & ~n6673;
  assign n6675 = ~n6672 & ~n6673;
  assign n6676 = ~n6674 & ~n6675;
  assign n6677 = n6500 & n6527;
  assign n6678 = ~n6500 & ~n6527;
  assign n6679 = ~n6677 & ~n6678;
  assign n6680 = n6453 & ~n6679;
  assign n6681 = ~n6453 & n6679;
  assign n6682 = ~n6680 & ~n6681;
  assign n6683 = ~n6360 & ~n6386;
  assign n6684 = ~n6383 & ~n6683;
  assign n6685 = n6682 & ~n6684;
  assign n6686 = ~n6682 & n6684;
  assign n6687 = ~n6685 & ~n6686;
  assign n6688 = ~n6676 & n6687;
  assign n6689 = ~n6676 & ~n6688;
  assign n6690 = n6687 & ~n6688;
  assign n6691 = ~n6689 & ~n6690;
  assign n6692 = ~n6657 & ~n6691;
  assign n6693 = ~n6657 & ~n6692;
  assign n6694 = ~n6691 & ~n6692;
  assign n6695 = ~n6693 & ~n6694;
  assign n6696 = ~n6343 & ~n6398;
  assign n6697 = n6695 & n6696;
  assign n6698 = ~n6695 & ~n6696;
  assign n6699 = ~n6697 & ~n6698;
  assign n6700 = ~n6390 & ~n6394;
  assign n6701 = n6368 & n6380;
  assign n6702 = ~n6368 & ~n6380;
  assign n6703 = ~n6701 & ~n6702;
  assign n6704 = n6482 & ~n6703;
  assign n6705 = ~n6482 & n6703;
  assign n6706 = ~n6704 & ~n6705;
  assign n6707 = ~n6469 & ~n6485;
  assign n6708 = ~n6515 & ~n6530;
  assign n6709 = n6707 & n6708;
  assign n6710 = ~n6707 & ~n6708;
  assign n6711 = ~n6709 & ~n6710;
  assign n6712 = n6706 & n6711;
  assign n6713 = ~n6706 & ~n6711;
  assign n6714 = ~n6712 & ~n6713;
  assign n6715 = ~n6700 & n6714;
  assign n6716 = n6700 & ~n6714;
  assign n6717 = ~n6715 & ~n6716;
  assign n6718 = pi13  & pi42 ;
  assign n6719 = pi11  & pi44 ;
  assign n6720 = ~n6718 & ~n6719;
  assign n6721 = n1377 & n4329;
  assign n6722 = pi10  & pi45 ;
  assign n6723 = ~n6720 & n6722;
  assign n6724 = ~n6721 & n6723;
  assign n6725 = ~n6721 & ~n6724;
  assign n6726 = ~n6720 & n6725;
  assign n6727 = n6722 & ~n6724;
  assign n6728 = ~n6726 & ~n6727;
  assign n6729 = pi12  & pi43 ;
  assign n6730 = pi26  & pi29 ;
  assign n6731 = n2191 & n6730;
  assign n6732 = ~n2191 & ~n6730;
  assign n6733 = n6729 & ~n6731;
  assign n6734 = ~n6732 & n6733;
  assign n6735 = n6729 & ~n6734;
  assign n6736 = ~n6731 & ~n6734;
  assign n6737 = ~n6732 & n6736;
  assign n6738 = ~n6735 & ~n6737;
  assign n6739 = ~n6728 & ~n6738;
  assign n6740 = ~n6728 & ~n6739;
  assign n6741 = ~n6738 & ~n6739;
  assign n6742 = ~n6740 & ~n6741;
  assign n6743 = pi16  & pi39 ;
  assign n6744 = n521 & n5823;
  assign n6745 = pi7  & pi48 ;
  assign n6746 = pi8  & pi47 ;
  assign n6747 = ~n6745 & ~n6746;
  assign n6748 = n6743 & ~n6744;
  assign n6749 = ~n6747 & n6748;
  assign n6750 = n6743 & ~n6749;
  assign n6751 = ~n6744 & ~n6749;
  assign n6752 = ~n6747 & n6751;
  assign n6753 = ~n6750 & ~n6752;
  assign n6754 = ~n6742 & ~n6753;
  assign n6755 = ~n6742 & ~n6754;
  assign n6756 = ~n6753 & ~n6754;
  assign n6757 = ~n6755 & ~n6756;
  assign n6758 = ~n6411 & ~n6415;
  assign n6759 = n6757 & n6758;
  assign n6760 = ~n6757 & ~n6758;
  assign n6761 = ~n6759 & ~n6760;
  assign n6762 = pi2  & pi53 ;
  assign n6763 = pi4  & pi51 ;
  assign n6764 = ~n6762 & ~n6763;
  assign n6765 = pi51  & pi53 ;
  assign n6766 = n249 & n6765;
  assign n6767 = pi0  & pi55 ;
  assign n6768 = ~n6764 & n6767;
  assign n6769 = ~n6766 & n6768;
  assign n6770 = ~n6766 & ~n6769;
  assign n6771 = ~n6764 & n6770;
  assign n6772 = n6767 & ~n6769;
  assign n6773 = ~n6771 & ~n6772;
  assign n6774 = pi20  & pi35 ;
  assign n6775 = n1481 & n3900;
  assign n6776 = pi21  & pi34 ;
  assign n6777 = ~n2438 & ~n6776;
  assign n6778 = n6774 & ~n6775;
  assign n6779 = ~n6777 & n6778;
  assign n6780 = n6774 & ~n6779;
  assign n6781 = ~n6775 & ~n6779;
  assign n6782 = ~n6777 & n6781;
  assign n6783 = ~n6780 & ~n6782;
  assign n6784 = ~n6773 & ~n6783;
  assign n6785 = ~n6773 & ~n6784;
  assign n6786 = ~n6783 & ~n6784;
  assign n6787 = ~n6785 & ~n6786;
  assign n6788 = pi23  & pi32 ;
  assign n6789 = n1789 & n2680;
  assign n6790 = pi24  & pi31 ;
  assign n6791 = pi25  & pi30 ;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = n6788 & ~n6789;
  assign n6794 = ~n6792 & n6793;
  assign n6795 = n6788 & ~n6794;
  assign n6796 = ~n6789 & ~n6794;
  assign n6797 = ~n6792 & n6796;
  assign n6798 = ~n6795 & ~n6797;
  assign n6799 = ~n6787 & ~n6798;
  assign n6800 = ~n6787 & ~n6799;
  assign n6801 = ~n6798 & ~n6799;
  assign n6802 = ~n6800 & ~n6801;
  assign n6803 = n6761 & ~n6802;
  assign n6804 = ~n6761 & n6802;
  assign n6805 = ~n6803 & ~n6804;
  assign n6806 = n6717 & n6805;
  assign n6807 = n6717 & ~n6806;
  assign n6808 = n6805 & ~n6806;
  assign n6809 = ~n6807 & ~n6808;
  assign n6810 = ~n6699 & n6809;
  assign n6811 = n6699 & ~n6809;
  assign n6812 = ~n6810 & ~n6811;
  assign n6813 = ~n6630 & n6812;
  assign n6814 = n6630 & ~n6812;
  assign n6815 = ~n6813 & ~n6814;
  assign n6816 = ~n6576 & n6815;
  assign n6817 = n6576 & ~n6815;
  assign n6818 = ~n6816 & ~n6817;
  assign n6819 = ~n6567 & ~n6573;
  assign n6820 = ~n6818 & n6819;
  assign n6821 = n6818 & ~n6819;
  assign po56  = ~n6820 & ~n6821;
  assign n6823 = ~n6627 & ~n6813;
  assign n6824 = pi7  & pi49 ;
  assign n6825 = pi17  & pi39 ;
  assign n6826 = ~n6824 & ~n6825;
  assign n6827 = n6824 & n6825;
  assign n6828 = pi6  & pi50 ;
  assign n6829 = ~n6826 & n6828;
  assign n6830 = ~n6827 & n6829;
  assign n6831 = ~n6827 & ~n6830;
  assign n6832 = ~n6826 & n6831;
  assign n6833 = n6828 & ~n6830;
  assign n6834 = ~n6832 & ~n6833;
  assign n6835 = pi11  & pi45 ;
  assign n6836 = pi43  & pi44 ;
  assign n6837 = n952 & n6836;
  assign n6838 = pi12  & pi44 ;
  assign n6839 = ~n5743 & ~n6838;
  assign n6840 = n6835 & ~n6837;
  assign n6841 = ~n6839 & n6840;
  assign n6842 = n6835 & ~n6841;
  assign n6843 = ~n6837 & ~n6841;
  assign n6844 = ~n6839 & n6843;
  assign n6845 = ~n6842 & ~n6844;
  assign n6846 = ~n6834 & ~n6845;
  assign n6847 = ~n6834 & ~n6846;
  assign n6848 = ~n6845 & ~n6846;
  assign n6849 = ~n6847 & ~n6848;
  assign n6850 = pi16  & pi40 ;
  assign n6851 = pi15  & pi48 ;
  assign n6852 = n5233 & n6851;
  assign n6853 = pi8  & pi48 ;
  assign n6854 = pi15  & pi41 ;
  assign n6855 = ~n6853 & ~n6854;
  assign n6856 = n6850 & ~n6852;
  assign n6857 = ~n6855 & n6856;
  assign n6858 = n6850 & ~n6857;
  assign n6859 = ~n6852 & ~n6857;
  assign n6860 = ~n6855 & n6859;
  assign n6861 = ~n6858 & ~n6860;
  assign n6862 = ~n6849 & ~n6861;
  assign n6863 = ~n6849 & ~n6862;
  assign n6864 = ~n6861 & ~n6862;
  assign n6865 = ~n6863 & ~n6864;
  assign n6866 = pi22  & pi34 ;
  assign n6867 = pi23  & pi33 ;
  assign n6868 = ~n6866 & ~n6867;
  assign n6869 = n1806 & n3900;
  assign n6870 = pi20  & pi36 ;
  assign n6871 = ~n6868 & n6870;
  assign n6872 = ~n6869 & n6871;
  assign n6873 = ~n6869 & ~n6872;
  assign n6874 = ~n6868 & n6873;
  assign n6875 = n6870 & ~n6872;
  assign n6876 = ~n6874 & ~n6875;
  assign n6877 = pi24  & pi32 ;
  assign n6878 = n2310 & n2680;
  assign n6879 = pi25  & pi31 ;
  assign n6880 = pi26  & pi30 ;
  assign n6881 = ~n6879 & ~n6880;
  assign n6882 = n6877 & ~n6878;
  assign n6883 = ~n6881 & n6882;
  assign n6884 = n6877 & ~n6883;
  assign n6885 = ~n6878 & ~n6883;
  assign n6886 = ~n6881 & n6885;
  assign n6887 = ~n6884 & ~n6886;
  assign n6888 = ~n6876 & ~n6887;
  assign n6889 = ~n6876 & ~n6888;
  assign n6890 = ~n6887 & ~n6888;
  assign n6891 = ~n6889 & ~n6890;
  assign n6892 = pi9  & pi47 ;
  assign n6893 = pi14  & pi46 ;
  assign n6894 = n6011 & n6893;
  assign n6895 = pi14  & pi42 ;
  assign n6896 = pi10  & pi46 ;
  assign n6897 = ~n6895 & ~n6896;
  assign n6898 = n6892 & ~n6894;
  assign n6899 = ~n6897 & n6898;
  assign n6900 = n6892 & ~n6899;
  assign n6901 = ~n6894 & ~n6899;
  assign n6902 = ~n6897 & n6901;
  assign n6903 = ~n6900 & ~n6902;
  assign n6904 = ~n6891 & ~n6903;
  assign n6905 = ~n6891 & ~n6904;
  assign n6906 = ~n6903 & ~n6904;
  assign n6907 = ~n6905 & ~n6906;
  assign n6908 = ~n6865 & n6907;
  assign n6909 = n6865 & ~n6907;
  assign n6910 = ~n6908 & ~n6909;
  assign n6911 = pi54  & pi56 ;
  assign n6912 = n196 & n6911;
  assign n6913 = pi0  & pi56 ;
  assign n6914 = pi2  & pi54 ;
  assign n6915 = ~n6913 & ~n6914;
  assign n6916 = ~n6912 & ~n6915;
  assign n6917 = n6637 & n6916;
  assign n6918 = ~n6637 & ~n6916;
  assign n6919 = ~n6917 & ~n6918;
  assign n6920 = ~n6751 & n6919;
  assign n6921 = n6751 & ~n6919;
  assign n6922 = ~n6920 & ~n6921;
  assign n6923 = pi3  & pi53 ;
  assign n6924 = pi4  & pi52 ;
  assign n6925 = pi19  & pi37 ;
  assign n6926 = n6924 & n6925;
  assign n6927 = ~n6924 & ~n6925;
  assign n6928 = n6923 & ~n6926;
  assign n6929 = ~n6927 & n6928;
  assign n6930 = n6923 & ~n6929;
  assign n6931 = ~n6926 & ~n6929;
  assign n6932 = ~n6927 & n6931;
  assign n6933 = ~n6930 & ~n6932;
  assign n6934 = n6922 & ~n6933;
  assign n6935 = n6922 & ~n6934;
  assign n6936 = ~n6933 & ~n6934;
  assign n6937 = ~n6935 & ~n6936;
  assign n6938 = n6910 & n6937;
  assign n6939 = ~n6910 & ~n6937;
  assign n6940 = ~n6938 & ~n6939;
  assign n6941 = ~n6613 & ~n6616;
  assign n6942 = n6781 & n6796;
  assign n6943 = ~n6781 & ~n6796;
  assign n6944 = ~n6942 & ~n6943;
  assign n6945 = n6589 & ~n6944;
  assign n6946 = ~n6589 & n6944;
  assign n6947 = ~n6945 & ~n6946;
  assign n6948 = ~n6739 & ~n6754;
  assign n6949 = pi1  & pi55 ;
  assign n6950 = ~n1923 & ~n6949;
  assign n6951 = n1923 & n6949;
  assign n6952 = ~n6950 & ~n6951;
  assign n6953 = ~n6736 & n6952;
  assign n6954 = ~n6736 & ~n6953;
  assign n6955 = n6952 & ~n6953;
  assign n6956 = ~n6954 & ~n6955;
  assign n6957 = ~n6725 & ~n6956;
  assign n6958 = n6725 & n6956;
  assign n6959 = ~n6957 & ~n6958;
  assign n6960 = ~n6948 & n6959;
  assign n6961 = n6948 & ~n6959;
  assign n6962 = ~n6960 & ~n6961;
  assign n6963 = n6947 & n6962;
  assign n6964 = ~n6947 & ~n6962;
  assign n6965 = ~n6963 & ~n6964;
  assign n6966 = ~n6941 & n6965;
  assign n6967 = ~n6941 & ~n6966;
  assign n6968 = n6965 & ~n6966;
  assign n6969 = ~n6967 & ~n6968;
  assign n6970 = n6940 & ~n6969;
  assign n6971 = n6940 & ~n6970;
  assign n6972 = ~n6969 & ~n6970;
  assign n6973 = ~n6971 & ~n6972;
  assign n6974 = ~n6619 & ~n6623;
  assign n6975 = n6670 & n6770;
  assign n6976 = ~n6670 & ~n6770;
  assign n6977 = ~n6975 & ~n6976;
  assign n6978 = n6601 & ~n6977;
  assign n6979 = ~n6601 & n6977;
  assign n6980 = ~n6978 & ~n6979;
  assign n6981 = ~n6604 & ~n6610;
  assign n6982 = ~n6980 & n6981;
  assign n6983 = n6980 & ~n6981;
  assign n6984 = ~n6982 & ~n6983;
  assign n6985 = ~n6634 & ~n6649;
  assign n6986 = ~n6984 & n6985;
  assign n6987 = n6984 & ~n6985;
  assign n6988 = ~n6986 & ~n6987;
  assign n6989 = ~n6702 & ~n6705;
  assign n6990 = ~n6660 & ~n6673;
  assign n6991 = n6989 & n6990;
  assign n6992 = ~n6989 & ~n6990;
  assign n6993 = ~n6991 & ~n6992;
  assign n6994 = ~n6784 & ~n6799;
  assign n6995 = ~n6993 & n6994;
  assign n6996 = n6993 & ~n6994;
  assign n6997 = ~n6995 & ~n6996;
  assign n6998 = ~n6760 & ~n6803;
  assign n6999 = n6997 & ~n6998;
  assign n7000 = n6997 & ~n6999;
  assign n7001 = ~n6998 & ~n6999;
  assign n7002 = ~n7000 & ~n7001;
  assign n7003 = n6988 & ~n7002;
  assign n7004 = ~n6988 & n7002;
  assign n7005 = ~n7003 & ~n7004;
  assign n7006 = ~n6974 & n7005;
  assign n7007 = ~n6974 & ~n7006;
  assign n7008 = n7005 & ~n7006;
  assign n7009 = ~n7007 & ~n7008;
  assign n7010 = ~n6973 & ~n7009;
  assign n7011 = ~n6973 & ~n7010;
  assign n7012 = ~n7009 & ~n7010;
  assign n7013 = ~n7011 & ~n7012;
  assign n7014 = ~n6685 & ~n6688;
  assign n7015 = ~n6641 & ~n6645;
  assign n7016 = pi21  & pi35 ;
  assign n7017 = pi38  & pi51 ;
  assign n7018 = n1255 & n7017;
  assign n7019 = pi5  & pi51 ;
  assign n7020 = pi18  & pi38 ;
  assign n7021 = ~n7019 & ~n7020;
  assign n7022 = n7016 & ~n7018;
  assign n7023 = ~n7021 & n7022;
  assign n7024 = n7016 & ~n7023;
  assign n7025 = ~n7018 & ~n7023;
  assign n7026 = ~n7021 & n7025;
  assign n7027 = ~n7024 & ~n7026;
  assign n7028 = ~n7015 & ~n7027;
  assign n7029 = ~n7015 & ~n7028;
  assign n7030 = ~n7027 & ~n7028;
  assign n7031 = ~n7029 & ~n7030;
  assign n7032 = ~n6678 & ~n6681;
  assign n7033 = n7031 & n7032;
  assign n7034 = ~n7031 & ~n7032;
  assign n7035 = ~n7033 & ~n7034;
  assign n7036 = ~n6710 & ~n6712;
  assign n7037 = n7035 & ~n7036;
  assign n7038 = ~n7035 & n7036;
  assign n7039 = ~n7037 & ~n7038;
  assign n7040 = n7014 & ~n7039;
  assign n7041 = ~n7014 & n7039;
  assign n7042 = ~n7040 & ~n7041;
  assign n7043 = ~n6654 & ~n6692;
  assign n7044 = ~n7042 & n7043;
  assign n7045 = n7042 & ~n7043;
  assign n7046 = ~n7044 & ~n7045;
  assign n7047 = ~n6715 & ~n6806;
  assign n7048 = ~n7046 & n7047;
  assign n7049 = n7046 & ~n7047;
  assign n7050 = ~n7048 & ~n7049;
  assign n7051 = ~n6698 & ~n6811;
  assign n7052 = n7050 & ~n7051;
  assign n7053 = n7050 & ~n7052;
  assign n7054 = ~n7051 & ~n7052;
  assign n7055 = ~n7053 & ~n7054;
  assign n7056 = ~n7013 & ~n7055;
  assign n7057 = n7013 & n7055;
  assign n7058 = ~n7056 & ~n7057;
  assign n7059 = ~n6823 & n7058;
  assign n7060 = n6823 & ~n7058;
  assign n7061 = ~n7059 & ~n7060;
  assign n7062 = ~n6816 & ~n6821;
  assign n7063 = ~n7061 & n7062;
  assign n7064 = n7061 & ~n7062;
  assign po57  = ~n7063 & ~n7064;
  assign n7066 = ~n7052 & ~n7056;
  assign n7067 = ~n7045 & ~n7049;
  assign n7068 = ~n6953 & ~n6957;
  assign n7069 = ~n6920 & ~n6934;
  assign n7070 = n7068 & n7069;
  assign n7071 = ~n7068 & ~n7069;
  assign n7072 = ~n7070 & ~n7071;
  assign n7073 = ~n6888 & ~n6904;
  assign n7074 = ~n7072 & n7073;
  assign n7075 = n7072 & ~n7073;
  assign n7076 = ~n7074 & ~n7075;
  assign n7077 = ~n6865 & ~n6907;
  assign n7078 = ~n6939 & ~n7077;
  assign n7079 = n7076 & ~n7078;
  assign n7080 = ~n7076 & n7078;
  assign n7081 = ~n7079 & ~n7080;
  assign n7082 = ~n6846 & ~n6862;
  assign n7083 = n6859 & n6885;
  assign n7084 = ~n6859 & ~n6885;
  assign n7085 = ~n7083 & ~n7084;
  assign n7086 = n6831 & ~n7085;
  assign n7087 = ~n6831 & n7085;
  assign n7088 = ~n7086 & ~n7087;
  assign n7089 = n6873 & n6931;
  assign n7090 = ~n6873 & ~n6931;
  assign n7091 = ~n7089 & ~n7090;
  assign n7092 = ~n6912 & ~n6917;
  assign n7093 = ~n7091 & n7092;
  assign n7094 = n7091 & ~n7092;
  assign n7095 = ~n7093 & ~n7094;
  assign n7096 = n7088 & n7095;
  assign n7097 = ~n7088 & ~n7095;
  assign n7098 = ~n7096 & ~n7097;
  assign n7099 = ~n7082 & n7098;
  assign n7100 = n7082 & ~n7098;
  assign n7101 = ~n7099 & ~n7100;
  assign n7102 = n7081 & n7101;
  assign n7103 = ~n7081 & ~n7101;
  assign n7104 = ~n7102 & ~n7103;
  assign n7105 = n7067 & ~n7104;
  assign n7106 = ~n7067 & n7104;
  assign n7107 = ~n7105 & ~n7106;
  assign n7108 = ~n7037 & ~n7041;
  assign n7109 = n6901 & n7025;
  assign n7110 = ~n6901 & ~n7025;
  assign n7111 = ~n7109 & ~n7110;
  assign n7112 = n6843 & ~n7111;
  assign n7113 = ~n6843 & n7111;
  assign n7114 = ~n7112 & ~n7113;
  assign n7115 = ~n7028 & ~n7034;
  assign n7116 = ~n7114 & n7115;
  assign n7117 = n7114 & ~n7115;
  assign n7118 = ~n7116 & ~n7117;
  assign n7119 = pi8  & pi49 ;
  assign n7120 = pi16  & pi41 ;
  assign n7121 = ~n7119 & ~n7120;
  assign n7122 = pi16  & pi49 ;
  assign n7123 = n5233 & n7122;
  assign n7124 = pi7  & pi50 ;
  assign n7125 = ~n7121 & n7124;
  assign n7126 = ~n7123 & n7125;
  assign n7127 = ~n7123 & ~n7126;
  assign n7128 = ~n7121 & n7127;
  assign n7129 = n7124 & ~n7126;
  assign n7130 = ~n7128 & ~n7129;
  assign n7131 = pi21  & pi36 ;
  assign n7132 = n1806 & n3106;
  assign n7133 = pi22  & pi35 ;
  assign n7134 = pi23  & pi34 ;
  assign n7135 = ~n7133 & ~n7134;
  assign n7136 = n7131 & ~n7132;
  assign n7137 = ~n7135 & n7136;
  assign n7138 = n7131 & ~n7137;
  assign n7139 = ~n7132 & ~n7137;
  assign n7140 = ~n7135 & n7139;
  assign n7141 = ~n7138 & ~n7140;
  assign n7142 = ~n7130 & ~n7141;
  assign n7143 = ~n7130 & ~n7142;
  assign n7144 = ~n7141 & ~n7142;
  assign n7145 = ~n7143 & ~n7144;
  assign n7146 = pi24  & pi33 ;
  assign n7147 = n2310 & n3567;
  assign n7148 = pi25  & pi32 ;
  assign n7149 = pi26  & pi31 ;
  assign n7150 = ~n7148 & ~n7149;
  assign n7151 = n7146 & ~n7147;
  assign n7152 = ~n7150 & n7151;
  assign n7153 = n7146 & ~n7152;
  assign n7154 = ~n7147 & ~n7152;
  assign n7155 = ~n7150 & n7154;
  assign n7156 = ~n7153 & ~n7155;
  assign n7157 = ~n7145 & ~n7156;
  assign n7158 = ~n7145 & ~n7157;
  assign n7159 = ~n7156 & ~n7157;
  assign n7160 = ~n7158 & ~n7159;
  assign n7161 = n7118 & ~n7160;
  assign n7162 = ~n7118 & n7160;
  assign n7163 = ~n7161 & ~n7162;
  assign n7164 = ~n7108 & n7163;
  assign n7165 = ~n7108 & ~n7164;
  assign n7166 = n7163 & ~n7164;
  assign n7167 = ~n7165 & ~n7166;
  assign n7168 = ~n6992 & ~n6996;
  assign n7169 = pi2  & pi55 ;
  assign n7170 = pi4  & pi53 ;
  assign n7171 = ~n7169 & ~n7170;
  assign n7172 = pi53  & pi55 ;
  assign n7173 = n249 & n7172;
  assign n7174 = pi3  & pi54 ;
  assign n7175 = ~n7171 & n7174;
  assign n7176 = ~n7173 & n7175;
  assign n7177 = ~n7173 & ~n7176;
  assign n7178 = ~n7171 & n7177;
  assign n7179 = n7174 & ~n7176;
  assign n7180 = ~n7178 & ~n7179;
  assign n7181 = pi5  & pi52 ;
  assign n7182 = n1407 & n5055;
  assign n7183 = pi19  & pi38 ;
  assign n7184 = pi20  & pi37 ;
  assign n7185 = ~n7183 & ~n7184;
  assign n7186 = n7181 & ~n7182;
  assign n7187 = ~n7185 & n7186;
  assign n7188 = n7181 & ~n7187;
  assign n7189 = ~n7182 & ~n7187;
  assign n7190 = ~n7185 & n7189;
  assign n7191 = ~n7188 & ~n7190;
  assign n7192 = ~n7180 & ~n7191;
  assign n7193 = ~n7180 & ~n7192;
  assign n7194 = ~n7191 & ~n7192;
  assign n7195 = ~n7193 & ~n7194;
  assign n7196 = pi15  & pi42 ;
  assign n7197 = n591 & n5823;
  assign n7198 = pi9  & pi48 ;
  assign n7199 = pi10  & pi47 ;
  assign n7200 = ~n7198 & ~n7199;
  assign n7201 = n7196 & ~n7197;
  assign n7202 = ~n7200 & n7201;
  assign n7203 = n7196 & ~n7202;
  assign n7204 = ~n7197 & ~n7202;
  assign n7205 = ~n7200 & n7204;
  assign n7206 = ~n7203 & ~n7205;
  assign n7207 = ~n7195 & ~n7206;
  assign n7208 = ~n7195 & ~n7207;
  assign n7209 = ~n7206 & ~n7207;
  assign n7210 = ~n7208 & ~n7209;
  assign n7211 = pi13  & pi44 ;
  assign n7212 = pi11  & pi46 ;
  assign n7213 = ~n7211 & ~n7212;
  assign n7214 = pi44  & pi46 ;
  assign n7215 = n1377 & n7214;
  assign n7216 = pi14  & pi43 ;
  assign n7217 = ~n7213 & n7216;
  assign n7218 = ~n7215 & n7217;
  assign n7219 = ~n7215 & ~n7218;
  assign n7220 = ~n7213 & n7219;
  assign n7221 = n7216 & ~n7218;
  assign n7222 = ~n7220 & ~n7221;
  assign n7223 = pi12  & pi45 ;
  assign n7224 = n2191 & n4908;
  assign n7225 = pi27  & pi30 ;
  assign n7226 = ~n2915 & ~n7225;
  assign n7227 = n7223 & ~n7224;
  assign n7228 = ~n7226 & n7227;
  assign n7229 = n7223 & ~n7228;
  assign n7230 = ~n7224 & ~n7228;
  assign n7231 = ~n7226 & n7230;
  assign n7232 = ~n7229 & ~n7231;
  assign n7233 = ~n7222 & ~n7232;
  assign n7234 = ~n7222 & ~n7233;
  assign n7235 = ~n7232 & ~n7233;
  assign n7236 = ~n7234 & ~n7235;
  assign n7237 = pi18  & pi39 ;
  assign n7238 = pi17  & pi51 ;
  assign n7239 = n4636 & n7238;
  assign n7240 = pi6  & pi51 ;
  assign n7241 = pi17  & pi40 ;
  assign n7242 = ~n7240 & ~n7241;
  assign n7243 = n7237 & ~n7239;
  assign n7244 = ~n7242 & n7243;
  assign n7245 = n7237 & ~n7244;
  assign n7246 = ~n7239 & ~n7244;
  assign n7247 = ~n7242 & n7246;
  assign n7248 = ~n7245 & ~n7247;
  assign n7249 = ~n7236 & ~n7248;
  assign n7250 = ~n7236 & ~n7249;
  assign n7251 = ~n7248 & ~n7249;
  assign n7252 = ~n7250 & ~n7251;
  assign n7253 = n7210 & n7252;
  assign n7254 = ~n7210 & ~n7252;
  assign n7255 = ~n7253 & ~n7254;
  assign n7256 = ~n7168 & n7255;
  assign n7257 = n7168 & ~n7255;
  assign n7258 = ~n7256 & ~n7257;
  assign n7259 = n7167 & n7258;
  assign n7260 = ~n7167 & ~n7258;
  assign n7261 = ~n7259 & ~n7260;
  assign n7262 = n7107 & ~n7261;
  assign n7263 = n7107 & ~n7262;
  assign n7264 = ~n7261 & ~n7262;
  assign n7265 = ~n7263 & ~n7264;
  assign n7266 = ~n7006 & ~n7010;
  assign n7267 = ~n6966 & ~n6970;
  assign n7268 = ~n6999 & ~n7003;
  assign n7269 = ~n6983 & ~n6987;
  assign n7270 = ~n6960 & ~n6963;
  assign n7271 = n7269 & n7270;
  assign n7272 = ~n7269 & ~n7270;
  assign n7273 = ~n7271 & ~n7272;
  assign n7274 = pi0  & pi57 ;
  assign n7275 = n6951 & n7274;
  assign n7276 = n6951 & ~n7275;
  assign n7277 = ~n6951 & n7274;
  assign n7278 = ~n7276 & ~n7277;
  assign n7279 = pi1  & pi56 ;
  assign n7280 = pi29  & n7279;
  assign n7281 = pi29  & ~n7280;
  assign n7282 = n7279 & ~n7280;
  assign n7283 = ~n7281 & ~n7282;
  assign n7284 = ~n7278 & ~n7283;
  assign n7285 = ~n7278 & ~n7284;
  assign n7286 = ~n7283 & ~n7284;
  assign n7287 = ~n7285 & ~n7286;
  assign n7288 = ~n6943 & ~n6946;
  assign n7289 = n7287 & n7288;
  assign n7290 = ~n7287 & ~n7288;
  assign n7291 = ~n7289 & ~n7290;
  assign n7292 = ~n6976 & ~n6979;
  assign n7293 = ~n7291 & n7292;
  assign n7294 = n7291 & ~n7292;
  assign n7295 = ~n7293 & ~n7294;
  assign n7296 = n7273 & n7295;
  assign n7297 = ~n7273 & ~n7295;
  assign n7298 = ~n7296 & ~n7297;
  assign n7299 = ~n7268 & n7298;
  assign n7300 = n7268 & ~n7298;
  assign n7301 = ~n7299 & ~n7300;
  assign n7302 = ~n7267 & n7301;
  assign n7303 = n7267 & ~n7301;
  assign n7304 = ~n7302 & ~n7303;
  assign n7305 = ~n7266 & n7304;
  assign n7306 = ~n7266 & ~n7305;
  assign n7307 = n7304 & ~n7305;
  assign n7308 = ~n7306 & ~n7307;
  assign n7309 = ~n7265 & ~n7308;
  assign n7310 = n7265 & n7308;
  assign n7311 = ~n7309 & ~n7310;
  assign n7312 = ~n7066 & n7311;
  assign n7313 = n7066 & ~n7311;
  assign n7314 = ~n7312 & ~n7313;
  assign n7315 = ~n7059 & ~n7064;
  assign n7316 = ~n7314 & n7315;
  assign n7317 = n7314 & ~n7315;
  assign po58  = ~n7316 & ~n7317;
  assign n7319 = ~n7305 & ~n7309;
  assign n7320 = ~n7106 & ~n7262;
  assign n7321 = ~n7079 & ~n7102;
  assign n7322 = ~n7117 & ~n7161;
  assign n7323 = ~n7110 & ~n7113;
  assign n7324 = ~n7090 & ~n7094;
  assign n7325 = n7323 & n7324;
  assign n7326 = ~n7323 & ~n7324;
  assign n7327 = ~n7325 & ~n7326;
  assign n7328 = ~n7084 & ~n7087;
  assign n7329 = ~n7327 & n7328;
  assign n7330 = n7327 & ~n7328;
  assign n7331 = ~n7329 & ~n7330;
  assign n7332 = ~n7096 & ~n7099;
  assign n7333 = n7331 & ~n7332;
  assign n7334 = ~n7331 & n7332;
  assign n7335 = ~n7333 & ~n7334;
  assign n7336 = ~n7322 & n7335;
  assign n7337 = n7322 & ~n7335;
  assign n7338 = ~n7336 & ~n7337;
  assign n7339 = n7321 & ~n7338;
  assign n7340 = ~n7321 & n7338;
  assign n7341 = ~n7339 & ~n7340;
  assign n7342 = ~n7167 & n7258;
  assign n7343 = ~n7164 & ~n7342;
  assign n7344 = n7341 & ~n7343;
  assign n7345 = ~n7341 & n7343;
  assign n7346 = ~n7344 & ~n7345;
  assign n7347 = n7320 & ~n7346;
  assign n7348 = ~n7320 & n7346;
  assign n7349 = ~n7347 & ~n7348;
  assign n7350 = ~n7299 & ~n7302;
  assign n7351 = ~n7254 & ~n7256;
  assign n7352 = ~n7233 & ~n7249;
  assign n7353 = ~n7192 & ~n7207;
  assign n7354 = pi28  & pi30 ;
  assign n7355 = pi1  & pi57 ;
  assign n7356 = n7354 & n7355;
  assign n7357 = ~n7354 & ~n7355;
  assign n7358 = ~n7356 & ~n7357;
  assign n7359 = ~n7280 & ~n7358;
  assign n7360 = n7280 & n7358;
  assign n7361 = ~n7359 & ~n7360;
  assign n7362 = ~n7230 & n7361;
  assign n7363 = n7230 & ~n7361;
  assign n7364 = ~n7362 & ~n7363;
  assign n7365 = ~n7353 & n7364;
  assign n7366 = ~n7353 & ~n7365;
  assign n7367 = n7364 & ~n7365;
  assign n7368 = ~n7366 & ~n7367;
  assign n7369 = ~n7352 & ~n7368;
  assign n7370 = n7352 & n7368;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = ~n7351 & n7371;
  assign n7373 = n7351 & ~n7371;
  assign n7374 = ~n7372 & ~n7373;
  assign n7375 = ~n7142 & ~n7157;
  assign n7376 = n7154 & n7204;
  assign n7377 = ~n7154 & ~n7204;
  assign n7378 = ~n7376 & ~n7377;
  assign n7379 = n7139 & ~n7378;
  assign n7380 = ~n7139 & n7378;
  assign n7381 = ~n7379 & ~n7380;
  assign n7382 = n7177 & n7189;
  assign n7383 = ~n7177 & ~n7189;
  assign n7384 = ~n7382 & ~n7383;
  assign n7385 = n7219 & ~n7384;
  assign n7386 = ~n7219 & n7384;
  assign n7387 = ~n7385 & ~n7386;
  assign n7388 = n7381 & n7387;
  assign n7389 = ~n7381 & ~n7387;
  assign n7390 = ~n7388 & ~n7389;
  assign n7391 = ~n7375 & n7390;
  assign n7392 = n7375 & ~n7390;
  assign n7393 = ~n7391 & ~n7392;
  assign n7394 = n7374 & n7393;
  assign n7395 = ~n7374 & ~n7393;
  assign n7396 = ~n7394 & ~n7395;
  assign n7397 = n7350 & ~n7396;
  assign n7398 = ~n7350 & n7396;
  assign n7399 = ~n7397 & ~n7398;
  assign n7400 = pi0  & pi58 ;
  assign n7401 = pi4  & pi54 ;
  assign n7402 = ~n7400 & ~n7401;
  assign n7403 = n7400 & n7401;
  assign n7404 = pi2  & pi56 ;
  assign n7405 = ~n7402 & n7404;
  assign n7406 = ~n7403 & n7405;
  assign n7407 = ~n7403 & ~n7406;
  assign n7408 = ~n7402 & n7407;
  assign n7409 = n7404 & ~n7406;
  assign n7410 = ~n7408 & ~n7409;
  assign n7411 = pi5  & pi53 ;
  assign n7412 = n1593 & n5055;
  assign n7413 = pi20  & pi38 ;
  assign n7414 = pi21  & pi37 ;
  assign n7415 = ~n7413 & ~n7414;
  assign n7416 = n7411 & ~n7412;
  assign n7417 = ~n7415 & n7416;
  assign n7418 = n7411 & ~n7417;
  assign n7419 = ~n7412 & ~n7417;
  assign n7420 = ~n7415 & n7419;
  assign n7421 = ~n7418 & ~n7420;
  assign n7422 = ~n7410 & ~n7421;
  assign n7423 = ~n7410 & ~n7422;
  assign n7424 = ~n7421 & ~n7422;
  assign n7425 = ~n7423 & ~n7424;
  assign n7426 = pi17  & pi41 ;
  assign n7427 = pi42  & pi49 ;
  assign n7428 = n803 & n7427;
  assign n7429 = pi9  & pi49 ;
  assign n7430 = pi16  & pi42 ;
  assign n7431 = ~n7429 & ~n7430;
  assign n7432 = n7426 & ~n7428;
  assign n7433 = ~n7431 & n7432;
  assign n7434 = n7426 & ~n7433;
  assign n7435 = ~n7428 & ~n7433;
  assign n7436 = ~n7431 & n7435;
  assign n7437 = ~n7434 & ~n7436;
  assign n7438 = ~n7425 & ~n7437;
  assign n7439 = ~n7425 & ~n7438;
  assign n7440 = ~n7437 & ~n7438;
  assign n7441 = ~n7439 & ~n7440;
  assign n7442 = pi7  & pi51 ;
  assign n7443 = pi8  & pi50 ;
  assign n7444 = ~n7442 & ~n7443;
  assign n7445 = n521 & n6114;
  assign n7446 = pi18  & pi40 ;
  assign n7447 = ~n7444 & n7446;
  assign n7448 = ~n7445 & n7447;
  assign n7449 = ~n7445 & ~n7448;
  assign n7450 = ~n7444 & n7449;
  assign n7451 = n7446 & ~n7448;
  assign n7452 = ~n7450 & ~n7451;
  assign n7453 = pi22  & pi36 ;
  assign n7454 = n2110 & n3106;
  assign n7455 = pi23  & pi35 ;
  assign n7456 = pi24  & pi34 ;
  assign n7457 = ~n7455 & ~n7456;
  assign n7458 = n7453 & ~n7454;
  assign n7459 = ~n7457 & n7458;
  assign n7460 = n7453 & ~n7459;
  assign n7461 = ~n7454 & ~n7459;
  assign n7462 = ~n7457 & n7461;
  assign n7463 = ~n7460 & ~n7462;
  assign n7464 = ~n7452 & ~n7463;
  assign n7465 = ~n7452 & ~n7464;
  assign n7466 = ~n7463 & ~n7464;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = n2646 & n3567;
  assign n7469 = pi26  & pi32 ;
  assign n7470 = pi27  & pi31 ;
  assign n7471 = ~n7469 & ~n7470;
  assign n7472 = n3096 & ~n7468;
  assign n7473 = ~n7471 & n7472;
  assign n7474 = n3096 & ~n7473;
  assign n7475 = ~n7468 & ~n7473;
  assign n7476 = ~n7471 & n7475;
  assign n7477 = ~n7474 & ~n7476;
  assign n7478 = ~n7467 & ~n7477;
  assign n7479 = ~n7467 & ~n7478;
  assign n7480 = ~n7477 & ~n7478;
  assign n7481 = ~n7479 & ~n7480;
  assign n7482 = ~n7441 & n7481;
  assign n7483 = n7441 & ~n7481;
  assign n7484 = ~n7482 & ~n7483;
  assign n7485 = ~n7071 & ~n7075;
  assign n7486 = n7484 & n7485;
  assign n7487 = ~n7484 & ~n7485;
  assign n7488 = ~n7486 & ~n7487;
  assign n7489 = ~n7272 & ~n7296;
  assign n7490 = n7127 & n7246;
  assign n7491 = ~n7127 & ~n7246;
  assign n7492 = ~n7490 & ~n7491;
  assign n7493 = ~n7275 & ~n7284;
  assign n7494 = ~n7492 & n7493;
  assign n7495 = n7492 & ~n7493;
  assign n7496 = ~n7494 & ~n7495;
  assign n7497 = ~n7290 & ~n7294;
  assign n7498 = ~n7496 & n7497;
  assign n7499 = n7496 & ~n7497;
  assign n7500 = ~n7498 & ~n7499;
  assign n7501 = pi15  & pi43 ;
  assign n7502 = pi11  & pi47 ;
  assign n7503 = ~n7501 & ~n7502;
  assign n7504 = pi43  & pi47 ;
  assign n7505 = n1579 & n7504;
  assign n7506 = pi10  & pi48 ;
  assign n7507 = ~n7503 & n7506;
  assign n7508 = ~n7505 & n7507;
  assign n7509 = ~n7505 & ~n7508;
  assign n7510 = ~n7503 & n7509;
  assign n7511 = n7506 & ~n7508;
  assign n7512 = ~n7510 & ~n7511;
  assign n7513 = pi45  & pi46 ;
  assign n7514 = n952 & n7513;
  assign n7515 = pi13  & pi45 ;
  assign n7516 = pi12  & pi46 ;
  assign n7517 = ~n7515 & ~n7516;
  assign n7518 = n6171 & ~n7514;
  assign n7519 = ~n7517 & n7518;
  assign n7520 = n6171 & ~n7519;
  assign n7521 = ~n7514 & ~n7519;
  assign n7522 = ~n7517 & n7521;
  assign n7523 = ~n7520 & ~n7522;
  assign n7524 = ~n7512 & ~n7523;
  assign n7525 = ~n7512 & ~n7524;
  assign n7526 = ~n7523 & ~n7524;
  assign n7527 = ~n7525 & ~n7526;
  assign n7528 = pi3  & pi55 ;
  assign n7529 = pi6  & pi52 ;
  assign n7530 = pi19  & pi39 ;
  assign n7531 = n7529 & n7530;
  assign n7532 = ~n7529 & ~n7530;
  assign n7533 = n7528 & ~n7531;
  assign n7534 = ~n7532 & n7533;
  assign n7535 = n7528 & ~n7534;
  assign n7536 = ~n7531 & ~n7534;
  assign n7537 = ~n7532 & n7536;
  assign n7538 = ~n7535 & ~n7537;
  assign n7539 = ~n7527 & ~n7538;
  assign n7540 = ~n7527 & ~n7539;
  assign n7541 = ~n7538 & ~n7539;
  assign n7542 = ~n7540 & ~n7541;
  assign n7543 = ~n7500 & n7542;
  assign n7544 = n7500 & ~n7542;
  assign n7545 = ~n7543 & ~n7544;
  assign n7546 = ~n7489 & n7545;
  assign n7547 = ~n7489 & ~n7546;
  assign n7548 = n7545 & ~n7546;
  assign n7549 = ~n7547 & ~n7548;
  assign n7550 = n7488 & ~n7549;
  assign n7551 = n7488 & ~n7550;
  assign n7552 = ~n7549 & ~n7550;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = n7399 & ~n7553;
  assign n7555 = n7399 & ~n7554;
  assign n7556 = ~n7553 & ~n7554;
  assign n7557 = ~n7555 & ~n7556;
  assign n7558 = ~n7349 & n7557;
  assign n7559 = n7349 & ~n7557;
  assign n7560 = ~n7558 & ~n7559;
  assign n7561 = ~n7319 & n7560;
  assign n7562 = n7319 & ~n7560;
  assign n7563 = ~n7561 & ~n7562;
  assign n7564 = ~n7312 & ~n7317;
  assign n7565 = ~n7563 & n7564;
  assign n7566 = ~n7562 & ~n7564;
  assign n7567 = ~n7561 & n7566;
  assign po59  = ~n7565 & ~n7567;
  assign n7569 = ~n7398 & ~n7554;
  assign n7570 = ~n7546 & ~n7550;
  assign n7571 = ~n7372 & ~n7394;
  assign n7572 = ~n7499 & ~n7544;
  assign n7573 = ~n7491 & ~n7495;
  assign n7574 = ~n7383 & ~n7386;
  assign n7575 = n7573 & n7574;
  assign n7576 = ~n7573 & ~n7574;
  assign n7577 = ~n7575 & ~n7576;
  assign n7578 = ~n7377 & ~n7380;
  assign n7579 = ~n7577 & n7578;
  assign n7580 = n7577 & ~n7578;
  assign n7581 = ~n7579 & ~n7580;
  assign n7582 = ~n7388 & ~n7391;
  assign n7583 = n7581 & ~n7582;
  assign n7584 = ~n7581 & n7582;
  assign n7585 = ~n7583 & ~n7584;
  assign n7586 = ~n7572 & n7585;
  assign n7587 = n7572 & ~n7585;
  assign n7588 = ~n7586 & ~n7587;
  assign n7589 = ~n7571 & n7588;
  assign n7590 = n7571 & ~n7588;
  assign n7591 = ~n7589 & ~n7590;
  assign n7592 = ~n7570 & n7591;
  assign n7593 = n7570 & ~n7591;
  assign n7594 = ~n7592 & ~n7593;
  assign n7595 = n7569 & ~n7594;
  assign n7596 = ~n7569 & n7594;
  assign n7597 = ~n7595 & ~n7596;
  assign n7598 = ~n7333 & ~n7336;
  assign n7599 = ~n7365 & ~n7369;
  assign n7600 = pi12  & pi47 ;
  assign n7601 = pi14  & pi45 ;
  assign n7602 = ~n7600 & ~n7601;
  assign n7603 = n1644 & n4899;
  assign n7604 = pi11  & pi48 ;
  assign n7605 = ~n7602 & n7604;
  assign n7606 = ~n7603 & n7605;
  assign n7607 = ~n7603 & ~n7606;
  assign n7608 = ~n7602 & n7607;
  assign n7609 = n7604 & ~n7606;
  assign n7610 = ~n7608 & ~n7609;
  assign n7611 = pi13  & pi46 ;
  assign n7612 = pi28  & pi31 ;
  assign n7613 = n4908 & n7612;
  assign n7614 = ~n4908 & ~n7612;
  assign n7615 = n7611 & ~n7613;
  assign n7616 = ~n7614 & n7615;
  assign n7617 = n7611 & ~n7616;
  assign n7618 = ~n7613 & ~n7616;
  assign n7619 = ~n7614 & n7618;
  assign n7620 = ~n7617 & ~n7619;
  assign n7621 = ~n7610 & ~n7620;
  assign n7622 = ~n7610 & ~n7621;
  assign n7623 = ~n7620 & ~n7621;
  assign n7624 = ~n7622 & ~n7623;
  assign n7625 = pi8  & pi51 ;
  assign n7626 = n989 & n6458;
  assign n7627 = pi16  & pi43 ;
  assign n7628 = pi17  & pi42 ;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = n7625 & ~n7626;
  assign n7631 = ~n7629 & n7630;
  assign n7632 = n7625 & ~n7631;
  assign n7633 = ~n7626 & ~n7631;
  assign n7634 = ~n7629 & n7633;
  assign n7635 = ~n7632 & ~n7634;
  assign n7636 = ~n7624 & ~n7635;
  assign n7637 = ~n7624 & ~n7636;
  assign n7638 = ~n7635 & ~n7636;
  assign n7639 = ~n7637 & ~n7638;
  assign n7640 = pi2  & pi57 ;
  assign n7641 = pi3  & pi56 ;
  assign n7642 = ~n7640 & ~n7641;
  assign n7643 = pi56  & pi57 ;
  assign n7644 = n218 & n7643;
  assign n7645 = n7356 & ~n7642;
  assign n7646 = ~n7644 & n7645;
  assign n7647 = ~n7644 & ~n7646;
  assign n7648 = ~n7642 & n7647;
  assign n7649 = n7356 & ~n7646;
  assign n7650 = ~n7648 & ~n7649;
  assign n7651 = n7475 & ~n7650;
  assign n7652 = ~n7475 & n7650;
  assign n7653 = ~n7651 & ~n7652;
  assign n7654 = pi4  & pi55 ;
  assign n7655 = pi5  & pi54 ;
  assign n7656 = pi19  & pi40 ;
  assign n7657 = n7655 & n7656;
  assign n7658 = ~n7655 & ~n7656;
  assign n7659 = n7654 & ~n7657;
  assign n7660 = ~n7658 & n7659;
  assign n7661 = n7654 & ~n7660;
  assign n7662 = ~n7657 & ~n7660;
  assign n7663 = ~n7658 & n7662;
  assign n7664 = ~n7661 & ~n7663;
  assign n7665 = ~n7653 & ~n7664;
  assign n7666 = n7653 & n7664;
  assign n7667 = ~n7665 & ~n7666;
  assign n7668 = n7639 & ~n7667;
  assign n7669 = ~n7639 & n7667;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = ~n7599 & n7670;
  assign n7672 = n7599 & ~n7670;
  assign n7673 = ~n7671 & ~n7672;
  assign n7674 = n7598 & ~n7673;
  assign n7675 = ~n7598 & n7673;
  assign n7676 = ~n7674 & ~n7675;
  assign n7677 = pi7  & pi52 ;
  assign n7678 = pi18  & pi41 ;
  assign n7679 = ~n7677 & ~n7678;
  assign n7680 = pi18  & pi52 ;
  assign n7681 = n5039 & n7680;
  assign n7682 = pi6  & pi53 ;
  assign n7683 = ~n7679 & n7682;
  assign n7684 = ~n7681 & n7683;
  assign n7685 = ~n7681 & ~n7684;
  assign n7686 = ~n7679 & n7685;
  assign n7687 = n7682 & ~n7684;
  assign n7688 = ~n7686 & ~n7687;
  assign n7689 = pi9  & pi50 ;
  assign n7690 = pi44  & pi49 ;
  assign n7691 = n1459 & n7690;
  assign n7692 = pi15  & pi44 ;
  assign n7693 = pi10  & pi49 ;
  assign n7694 = ~n7692 & ~n7693;
  assign n7695 = n7689 & ~n7691;
  assign n7696 = ~n7694 & n7695;
  assign n7697 = n7689 & ~n7696;
  assign n7698 = ~n7691 & ~n7696;
  assign n7699 = ~n7694 & n7698;
  assign n7700 = ~n7697 & ~n7699;
  assign n7701 = ~n7688 & ~n7700;
  assign n7702 = ~n7688 & ~n7701;
  assign n7703 = ~n7700 & ~n7701;
  assign n7704 = ~n7702 & ~n7703;
  assign n7705 = ~n7360 & ~n7362;
  assign n7706 = n7704 & n7705;
  assign n7707 = ~n7704 & ~n7705;
  assign n7708 = ~n7706 & ~n7707;
  assign n7709 = ~n7326 & ~n7330;
  assign n7710 = ~n7708 & n7709;
  assign n7711 = n7708 & ~n7709;
  assign n7712 = ~n7710 & ~n7711;
  assign n7713 = pi21  & pi38 ;
  assign n7714 = pi22  & pi37 ;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = n1481 & n5055;
  assign n7717 = pi20  & pi39 ;
  assign n7718 = ~n7715 & n7717;
  assign n7719 = ~n7716 & n7718;
  assign n7720 = ~n7716 & ~n7719;
  assign n7721 = ~n7715 & n7720;
  assign n7722 = n7717 & ~n7719;
  assign n7723 = ~n7721 & ~n7722;
  assign n7724 = pi23  & pi36 ;
  assign n7725 = n1789 & n3106;
  assign n7726 = pi24  & pi35 ;
  assign n7727 = pi25  & pi34 ;
  assign n7728 = ~n7726 & ~n7727;
  assign n7729 = n7724 & ~n7725;
  assign n7730 = ~n7728 & n7729;
  assign n7731 = n7724 & ~n7730;
  assign n7732 = ~n7725 & ~n7730;
  assign n7733 = ~n7728 & n7732;
  assign n7734 = ~n7731 & ~n7733;
  assign n7735 = ~n7723 & ~n7734;
  assign n7736 = ~n7723 & ~n7735;
  assign n7737 = ~n7734 & ~n7735;
  assign n7738 = ~n7736 & ~n7737;
  assign n7739 = pi26  & pi33 ;
  assign n7740 = pi32  & pi59 ;
  assign n7741 = n1701 & n7740;
  assign n7742 = pi0  & pi59 ;
  assign n7743 = pi27  & pi32 ;
  assign n7744 = ~n7742 & ~n7743;
  assign n7745 = n7739 & ~n7741;
  assign n7746 = ~n7744 & n7745;
  assign n7747 = n7739 & ~n7746;
  assign n7748 = ~n7741 & ~n7746;
  assign n7749 = ~n7744 & n7748;
  assign n7750 = ~n7747 & ~n7749;
  assign n7751 = ~n7738 & ~n7750;
  assign n7752 = ~n7738 & ~n7751;
  assign n7753 = ~n7750 & ~n7751;
  assign n7754 = ~n7752 & ~n7753;
  assign n7755 = n7712 & ~n7754;
  assign n7756 = ~n7712 & n7754;
  assign n7757 = ~n7755 & ~n7756;
  assign n7758 = n7676 & n7757;
  assign n7759 = n7676 & ~n7758;
  assign n7760 = n7757 & ~n7758;
  assign n7761 = ~n7759 & ~n7760;
  assign n7762 = ~n7340 & ~n7344;
  assign n7763 = ~n7524 & ~n7539;
  assign n7764 = ~n7464 & ~n7478;
  assign n7765 = n7763 & n7764;
  assign n7766 = ~n7763 & ~n7764;
  assign n7767 = ~n7765 & ~n7766;
  assign n7768 = ~n7422 & ~n7438;
  assign n7769 = ~n7767 & n7768;
  assign n7770 = n7767 & ~n7768;
  assign n7771 = ~n7769 & ~n7770;
  assign n7772 = ~n7441 & ~n7481;
  assign n7773 = ~n7487 & ~n7772;
  assign n7774 = n7407 & n7536;
  assign n7775 = ~n7407 & ~n7536;
  assign n7776 = ~n7774 & ~n7775;
  assign n7777 = n7435 & ~n7776;
  assign n7778 = ~n7435 & n7776;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = n7419 & n7461;
  assign n7781 = ~n7419 & ~n7461;
  assign n7782 = ~n7780 & ~n7781;
  assign n7783 = n7449 & ~n7782;
  assign n7784 = ~n7449 & n7782;
  assign n7785 = ~n7783 & ~n7784;
  assign n7786 = pi58  & n2252;
  assign n7787 = pi1  & pi58 ;
  assign n7788 = ~pi30  & ~n7787;
  assign n7789 = ~n7786 & ~n7788;
  assign n7790 = n7521 & ~n7789;
  assign n7791 = ~n7521 & n7789;
  assign n7792 = ~n7790 & ~n7791;
  assign n7793 = ~n7509 & n7792;
  assign n7794 = n7509 & ~n7792;
  assign n7795 = ~n7793 & ~n7794;
  assign n7796 = n7785 & n7795;
  assign n7797 = n7785 & ~n7796;
  assign n7798 = n7795 & ~n7796;
  assign n7799 = ~n7797 & ~n7798;
  assign n7800 = n7779 & ~n7799;
  assign n7801 = ~n7779 & n7799;
  assign n7802 = ~n7800 & ~n7801;
  assign n7803 = ~n7773 & n7802;
  assign n7804 = ~n7773 & ~n7803;
  assign n7805 = n7802 & ~n7803;
  assign n7806 = ~n7804 & ~n7805;
  assign n7807 = n7771 & ~n7806;
  assign n7808 = ~n7771 & n7806;
  assign n7809 = ~n7807 & ~n7808;
  assign n7810 = ~n7762 & n7809;
  assign n7811 = n7762 & ~n7809;
  assign n7812 = ~n7810 & ~n7811;
  assign n7813 = ~n7761 & n7812;
  assign n7814 = n7761 & ~n7812;
  assign n7815 = ~n7813 & ~n7814;
  assign n7816 = n7597 & n7815;
  assign n7817 = ~n7597 & ~n7815;
  assign n7818 = ~n7816 & ~n7817;
  assign n7819 = ~n7348 & ~n7559;
  assign n7820 = ~n7818 & n7819;
  assign n7821 = n7818 & ~n7819;
  assign n7822 = ~n7820 & ~n7821;
  assign n7823 = ~n7561 & ~n7566;
  assign n7824 = ~n7822 & n7823;
  assign n7825 = n7822 & ~n7823;
  assign po60  = ~n7824 & ~n7825;
  assign n7827 = ~n7596 & ~n7816;
  assign n7828 = ~n7810 & ~n7813;
  assign n7829 = ~n7675 & ~n7758;
  assign n7830 = ~n7803 & ~n7807;
  assign n7831 = ~n7781 & ~n7784;
  assign n7832 = ~n7775 & ~n7778;
  assign n7833 = n7831 & n7832;
  assign n7834 = ~n7831 & ~n7832;
  assign n7835 = ~n7833 & ~n7834;
  assign n7836 = ~n7475 & ~n7650;
  assign n7837 = ~n7665 & ~n7836;
  assign n7838 = ~n7835 & n7837;
  assign n7839 = n7835 & ~n7837;
  assign n7840 = ~n7838 & ~n7839;
  assign n7841 = ~n7766 & ~n7770;
  assign n7842 = ~n7840 & n7841;
  assign n7843 = n7840 & ~n7841;
  assign n7844 = ~n7842 & ~n7843;
  assign n7845 = ~n7711 & ~n7755;
  assign n7846 = n7844 & ~n7845;
  assign n7847 = ~n7844 & n7845;
  assign n7848 = ~n7846 & ~n7847;
  assign n7849 = ~n7830 & n7848;
  assign n7850 = n7830 & ~n7848;
  assign n7851 = ~n7849 & ~n7850;
  assign n7852 = ~n7829 & n7851;
  assign n7853 = n7829 & ~n7851;
  assign n7854 = ~n7852 & ~n7853;
  assign n7855 = n7828 & ~n7854;
  assign n7856 = ~n7828 & n7854;
  assign n7857 = ~n7855 & ~n7856;
  assign n7858 = ~n7796 & ~n7800;
  assign n7859 = pi0  & pi60 ;
  assign n7860 = n7786 & n7859;
  assign n7861 = n7786 & ~n7860;
  assign n7862 = ~n7786 & n7859;
  assign n7863 = ~n7861 & ~n7862;
  assign n7864 = pi1  & pi59 ;
  assign n7865 = pi29  & pi31 ;
  assign n7866 = n7864 & n7865;
  assign n7867 = n7864 & ~n7866;
  assign n7868 = n7865 & ~n7866;
  assign n7869 = ~n7867 & ~n7868;
  assign n7870 = ~n7863 & ~n7869;
  assign n7871 = ~n7863 & ~n7870;
  assign n7872 = ~n7869 & ~n7870;
  assign n7873 = ~n7871 & ~n7872;
  assign n7874 = pi27  & pi33 ;
  assign n7875 = pi28  & pi32 ;
  assign n7876 = pi23  & pi37 ;
  assign n7877 = n7875 & n7876;
  assign n7878 = ~n7875 & ~n7876;
  assign n7879 = n7874 & ~n7877;
  assign n7880 = ~n7878 & n7879;
  assign n7881 = n7874 & ~n7880;
  assign n7882 = ~n7877 & ~n7880;
  assign n7883 = ~n7878 & n7882;
  assign n7884 = ~n7881 & ~n7883;
  assign n7885 = ~n7873 & ~n7884;
  assign n7886 = ~n7873 & ~n7885;
  assign n7887 = ~n7884 & ~n7885;
  assign n7888 = ~n7886 & ~n7887;
  assign n7889 = ~n7791 & ~n7793;
  assign n7890 = n7888 & n7889;
  assign n7891 = ~n7888 & ~n7889;
  assign n7892 = ~n7890 & ~n7891;
  assign n7893 = pi8  & pi52 ;
  assign n7894 = pi18  & pi42 ;
  assign n7895 = ~n7893 & ~n7894;
  assign n7896 = n7893 & n7894;
  assign n7897 = pi7  & pi53 ;
  assign n7898 = ~n7895 & n7897;
  assign n7899 = ~n7896 & n7898;
  assign n7900 = ~n7896 & ~n7899;
  assign n7901 = ~n7895 & n7900;
  assign n7902 = n7897 & ~n7899;
  assign n7903 = ~n7901 & ~n7902;
  assign n7904 = n952 & n5823;
  assign n7905 = pi12  & pi48 ;
  assign n7906 = pi13  & pi47 ;
  assign n7907 = ~n7905 & ~n7906;
  assign n7908 = n6893 & ~n7904;
  assign n7909 = ~n7907 & n7908;
  assign n7910 = n6893 & ~n7909;
  assign n7911 = ~n7904 & ~n7909;
  assign n7912 = ~n7907 & n7911;
  assign n7913 = ~n7910 & ~n7912;
  assign n7914 = ~n7903 & ~n7913;
  assign n7915 = ~n7903 & ~n7914;
  assign n7916 = ~n7913 & ~n7914;
  assign n7917 = ~n7915 & ~n7916;
  assign n7918 = pi5  & pi55 ;
  assign n7919 = pi6  & pi54 ;
  assign n7920 = pi19  & pi41 ;
  assign n7921 = n7919 & n7920;
  assign n7922 = ~n7919 & ~n7920;
  assign n7923 = n7918 & ~n7921;
  assign n7924 = ~n7922 & n7923;
  assign n7925 = n7918 & ~n7924;
  assign n7926 = ~n7921 & ~n7924;
  assign n7927 = ~n7922 & n7926;
  assign n7928 = ~n7925 & ~n7927;
  assign n7929 = ~n7917 & ~n7928;
  assign n7930 = ~n7917 & ~n7929;
  assign n7931 = ~n7928 & ~n7929;
  assign n7932 = ~n7930 & ~n7931;
  assign n7933 = ~n7892 & n7932;
  assign n7934 = n7892 & ~n7932;
  assign n7935 = ~n7933 & ~n7934;
  assign n7936 = ~n7858 & n7935;
  assign n7937 = n7858 & ~n7935;
  assign n7938 = ~n7936 & ~n7937;
  assign n7939 = ~n7583 & ~n7586;
  assign n7940 = pi3  & pi57 ;
  assign n7941 = pi4  & pi56 ;
  assign n7942 = ~n7940 & ~n7941;
  assign n7943 = n209 & n7643;
  assign n7944 = pi2  & pi58 ;
  assign n7945 = ~n7942 & n7944;
  assign n7946 = ~n7943 & n7945;
  assign n7947 = ~n7943 & ~n7946;
  assign n7948 = ~n7942 & n7947;
  assign n7949 = n7944 & ~n7946;
  assign n7950 = ~n7948 & ~n7949;
  assign n7951 = pi20  & pi40 ;
  assign n7952 = n1481 & n4736;
  assign n7953 = pi21  & pi39 ;
  assign n7954 = pi22  & pi38 ;
  assign n7955 = ~n7953 & ~n7954;
  assign n7956 = n7951 & ~n7952;
  assign n7957 = ~n7955 & n7956;
  assign n7958 = n7951 & ~n7957;
  assign n7959 = ~n7952 & ~n7957;
  assign n7960 = ~n7955 & n7959;
  assign n7961 = ~n7958 & ~n7960;
  assign n7962 = ~n7950 & ~n7961;
  assign n7963 = ~n7950 & ~n7962;
  assign n7964 = ~n7961 & ~n7962;
  assign n7965 = ~n7963 & ~n7964;
  assign n7966 = pi24  & pi36 ;
  assign n7967 = n2310 & n3106;
  assign n7968 = pi25  & pi35 ;
  assign n7969 = pi26  & pi34 ;
  assign n7970 = ~n7968 & ~n7969;
  assign n7971 = n7966 & ~n7967;
  assign n7972 = ~n7970 & n7971;
  assign n7973 = n7966 & ~n7972;
  assign n7974 = ~n7967 & ~n7972;
  assign n7975 = ~n7970 & n7974;
  assign n7976 = ~n7973 & ~n7975;
  assign n7977 = ~n7965 & ~n7976;
  assign n7978 = ~n7965 & ~n7977;
  assign n7979 = ~n7976 & ~n7977;
  assign n7980 = ~n7978 & ~n7979;
  assign n7981 = ~n7576 & ~n7580;
  assign n7982 = n7980 & n7981;
  assign n7983 = ~n7980 & ~n7981;
  assign n7984 = ~n7982 & ~n7983;
  assign n7985 = pi17  & pi43 ;
  assign n7986 = pi44  & pi51 ;
  assign n7987 = n803 & n7986;
  assign n7988 = pi9  & pi51 ;
  assign n7989 = pi16  & pi44 ;
  assign n7990 = ~n7988 & ~n7989;
  assign n7991 = n7985 & ~n7987;
  assign n7992 = ~n7990 & n7991;
  assign n7993 = n7985 & ~n7992;
  assign n7994 = ~n7987 & ~n7992;
  assign n7995 = ~n7990 & n7994;
  assign n7996 = ~n7993 & ~n7995;
  assign n7997 = n7607 & ~n7996;
  assign n7998 = ~n7607 & n7996;
  assign n7999 = ~n7997 & ~n7998;
  assign n8000 = pi10  & pi50 ;
  assign n8001 = pi45  & pi49 ;
  assign n8002 = n1579 & n8001;
  assign n8003 = pi11  & pi49 ;
  assign n8004 = pi15  & pi45 ;
  assign n8005 = ~n8003 & ~n8004;
  assign n8006 = n8000 & ~n8002;
  assign n8007 = ~n8005 & n8006;
  assign n8008 = n8000 & ~n8007;
  assign n8009 = ~n8002 & ~n8007;
  assign n8010 = ~n8005 & n8009;
  assign n8011 = ~n8008 & ~n8010;
  assign n8012 = ~n7999 & ~n8011;
  assign n8013 = n7999 & n8011;
  assign n8014 = ~n8012 & ~n8013;
  assign n8015 = ~n7984 & ~n8014;
  assign n8016 = n7984 & n8014;
  assign n8017 = ~n8015 & ~n8016;
  assign n8018 = ~n7939 & n8017;
  assign n8019 = ~n7939 & ~n8018;
  assign n8020 = n8017 & ~n8018;
  assign n8021 = ~n8019 & ~n8020;
  assign n8022 = n7938 & ~n8021;
  assign n8023 = n7938 & ~n8022;
  assign n8024 = ~n8021 & ~n8022;
  assign n8025 = ~n8023 & ~n8024;
  assign n8026 = ~n7589 & ~n7592;
  assign n8027 = n7633 & n7685;
  assign n8028 = ~n7633 & ~n7685;
  assign n8029 = ~n8027 & ~n8028;
  assign n8030 = n7618 & ~n8029;
  assign n8031 = ~n7618 & n8029;
  assign n8032 = ~n8030 & ~n8031;
  assign n8033 = ~n7735 & ~n7751;
  assign n8034 = ~n8032 & n8033;
  assign n8035 = n8032 & ~n8033;
  assign n8036 = ~n8034 & ~n8035;
  assign n8037 = ~n7621 & ~n7636;
  assign n8038 = ~n8036 & n8037;
  assign n8039 = n8036 & ~n8037;
  assign n8040 = ~n8038 & ~n8039;
  assign n8041 = ~n7669 & ~n7671;
  assign n8042 = ~n7701 & ~n7707;
  assign n8043 = n7662 & n7720;
  assign n8044 = ~n7662 & ~n7720;
  assign n8045 = ~n8043 & ~n8044;
  assign n8046 = n7732 & ~n8045;
  assign n8047 = ~n7732 & n8045;
  assign n8048 = ~n8046 & ~n8047;
  assign n8049 = n7647 & n7748;
  assign n8050 = ~n7647 & ~n7748;
  assign n8051 = ~n8049 & ~n8050;
  assign n8052 = n7698 & ~n8051;
  assign n8053 = ~n7698 & n8051;
  assign n8054 = ~n8052 & ~n8053;
  assign n8055 = n8048 & n8054;
  assign n8056 = ~n8048 & ~n8054;
  assign n8057 = ~n8055 & ~n8056;
  assign n8058 = ~n8042 & n8057;
  assign n8059 = n8042 & ~n8057;
  assign n8060 = ~n8058 & ~n8059;
  assign n8061 = ~n8041 & n8060;
  assign n8062 = ~n8041 & ~n8061;
  assign n8063 = n8060 & ~n8061;
  assign n8064 = ~n8062 & ~n8063;
  assign n8065 = n8040 & ~n8064;
  assign n8066 = ~n8040 & n8064;
  assign n8067 = ~n8065 & ~n8066;
  assign n8068 = ~n8026 & n8067;
  assign n8069 = ~n8026 & ~n8068;
  assign n8070 = n8067 & ~n8068;
  assign n8071 = ~n8069 & ~n8070;
  assign n8072 = ~n8025 & ~n8071;
  assign n8073 = n8025 & n8071;
  assign n8074 = ~n8072 & ~n8073;
  assign n8075 = n7857 & n8074;
  assign n8076 = ~n7857 & ~n8074;
  assign n8077 = ~n8075 & ~n8076;
  assign n8078 = n7827 & ~n8077;
  assign n8079 = ~n7827 & n8077;
  assign n8080 = ~n8078 & ~n8079;
  assign n8081 = ~n7821 & ~n7825;
  assign n8082 = ~n8080 & n8081;
  assign n8083 = n8080 & ~n8081;
  assign po61  = ~n8082 & ~n8083;
  assign n8085 = ~n7856 & ~n8075;
  assign n8086 = ~n8068 & ~n8072;
  assign n8087 = ~n8018 & ~n8022;
  assign n8088 = ~n8035 & ~n8039;
  assign n8089 = pi7  & pi54 ;
  assign n8090 = pi8  & pi53 ;
  assign n8091 = ~n8089 & ~n8090;
  assign n8092 = pi53  & pi54 ;
  assign n8093 = n521 & n8092;
  assign n8094 = pi19  & pi42 ;
  assign n8095 = ~n8091 & n8094;
  assign n8096 = ~n8093 & n8095;
  assign n8097 = ~n8093 & ~n8096;
  assign n8098 = ~n8091 & n8097;
  assign n8099 = n8094 & ~n8096;
  assign n8100 = ~n8098 & ~n8099;
  assign n8101 = pi18  & pi43 ;
  assign n8102 = pi44  & pi52 ;
  assign n8103 = n1577 & n8102;
  assign n8104 = pi9  & pi52 ;
  assign n8105 = pi17  & pi44 ;
  assign n8106 = ~n8104 & ~n8105;
  assign n8107 = n8101 & ~n8103;
  assign n8108 = ~n8106 & n8107;
  assign n8109 = n8101 & ~n8108;
  assign n8110 = ~n8103 & ~n8108;
  assign n8111 = ~n8106 & n8110;
  assign n8112 = ~n8109 & ~n8111;
  assign n8113 = ~n8100 & ~n8112;
  assign n8114 = ~n8100 & ~n8113;
  assign n8115 = ~n8112 & ~n8113;
  assign n8116 = ~n8114 & ~n8115;
  assign n8117 = pi26  & pi35 ;
  assign n8118 = n2191 & n3900;
  assign n8119 = pi28  & pi33 ;
  assign n8120 = ~n3278 & ~n8119;
  assign n8121 = n8117 & ~n8118;
  assign n8122 = ~n8120 & n8121;
  assign n8123 = n8117 & ~n8122;
  assign n8124 = ~n8118 & ~n8122;
  assign n8125 = ~n8120 & n8124;
  assign n8126 = ~n8123 & ~n8125;
  assign n8127 = ~n8116 & ~n8126;
  assign n8128 = ~n8116 & ~n8127;
  assign n8129 = ~n8126 & ~n8127;
  assign n8130 = ~n8128 & ~n8129;
  assign n8131 = ~n8055 & ~n8058;
  assign n8132 = ~n8130 & ~n8131;
  assign n8133 = ~n8130 & ~n8132;
  assign n8134 = ~n8131 & ~n8132;
  assign n8135 = ~n8133 & ~n8134;
  assign n8136 = ~n8088 & ~n8135;
  assign n8137 = ~n8088 & ~n8136;
  assign n8138 = ~n8135 & ~n8136;
  assign n8139 = ~n8137 & ~n8138;
  assign n8140 = ~n7983 & ~n8016;
  assign n8141 = ~n8050 & ~n8053;
  assign n8142 = ~n8028 & ~n8031;
  assign n8143 = pi23  & pi38 ;
  assign n8144 = pi57  & pi58 ;
  assign n8145 = n209 & n8144;
  assign n8146 = pi3  & pi58 ;
  assign n8147 = pi4  & pi57 ;
  assign n8148 = ~n8146 & ~n8147;
  assign n8149 = n8143 & ~n8145;
  assign n8150 = ~n8148 & n8149;
  assign n8151 = n8143 & ~n8150;
  assign n8152 = ~n8145 & ~n8150;
  assign n8153 = ~n8148 & n8152;
  assign n8154 = ~n8151 & ~n8153;
  assign n8155 = ~n8142 & ~n8154;
  assign n8156 = ~n8142 & ~n8155;
  assign n8157 = ~n8154 & ~n8155;
  assign n8158 = ~n8156 & ~n8157;
  assign n8159 = ~n8141 & ~n8158;
  assign n8160 = ~n8141 & ~n8159;
  assign n8161 = ~n8158 & ~n8159;
  assign n8162 = ~n8160 & ~n8161;
  assign n8163 = ~n7607 & ~n7996;
  assign n8164 = ~n8012 & ~n8163;
  assign n8165 = ~n8044 & ~n8047;
  assign n8166 = pi1  & pi60 ;
  assign n8167 = pi31  & n8166;
  assign n8168 = ~pi31  & ~n8166;
  assign n8169 = ~n8167 & ~n8168;
  assign n8170 = n7866 & n8169;
  assign n8171 = ~n7866 & ~n8169;
  assign n8172 = ~n8170 & ~n8171;
  assign n8173 = ~n7911 & n8172;
  assign n8174 = n7911 & ~n8172;
  assign n8175 = ~n8173 & ~n8174;
  assign n8176 = ~n8165 & n8175;
  assign n8177 = n8165 & ~n8175;
  assign n8178 = ~n8176 & ~n8177;
  assign n8179 = ~n8164 & n8178;
  assign n8180 = n8164 & ~n8178;
  assign n8181 = ~n8179 & ~n8180;
  assign n8182 = ~n8162 & n8181;
  assign n8183 = ~n8162 & ~n8182;
  assign n8184 = n8181 & ~n8182;
  assign n8185 = ~n8183 & ~n8184;
  assign n8186 = ~n8140 & ~n8185;
  assign n8187 = n8140 & n8185;
  assign n8188 = ~n8186 & ~n8187;
  assign n8189 = ~n8139 & n8188;
  assign n8190 = ~n8139 & ~n8189;
  assign n8191 = n8188 & ~n8189;
  assign n8192 = ~n8190 & ~n8191;
  assign n8193 = ~n8087 & ~n8192;
  assign n8194 = n8087 & n8192;
  assign n8195 = ~n8193 & ~n8194;
  assign n8196 = ~n8086 & n8195;
  assign n8197 = ~n8086 & ~n8196;
  assign n8198 = n8195 & ~n8196;
  assign n8199 = ~n8197 & ~n8198;
  assign n8200 = ~n7934 & ~n7936;
  assign n8201 = n7900 & n7994;
  assign n8202 = ~n7900 & ~n7994;
  assign n8203 = ~n8201 & ~n8202;
  assign n8204 = ~n7860 & ~n7870;
  assign n8205 = ~n8203 & n8204;
  assign n8206 = n8203 & ~n8204;
  assign n8207 = ~n8205 & ~n8206;
  assign n8208 = ~n7914 & ~n7929;
  assign n8209 = ~n8207 & n8208;
  assign n8210 = n8207 & ~n8208;
  assign n8211 = ~n8209 & ~n8210;
  assign n8212 = ~n7885 & ~n7891;
  assign n8213 = ~n8211 & n8212;
  assign n8214 = n8211 & ~n8212;
  assign n8215 = ~n8213 & ~n8214;
  assign n8216 = ~n7962 & ~n7977;
  assign n8217 = n7882 & n7974;
  assign n8218 = ~n7882 & ~n7974;
  assign n8219 = ~n8217 & ~n8218;
  assign n8220 = n7959 & ~n8219;
  assign n8221 = ~n7959 & n8219;
  assign n8222 = ~n8220 & ~n8221;
  assign n8223 = n7926 & n7947;
  assign n8224 = ~n7926 & ~n7947;
  assign n8225 = ~n8223 & ~n8224;
  assign n8226 = n8009 & ~n8225;
  assign n8227 = ~n8009 & n8225;
  assign n8228 = ~n8226 & ~n8227;
  assign n8229 = ~n8222 & ~n8228;
  assign n8230 = n8222 & n8228;
  assign n8231 = ~n8229 & ~n8230;
  assign n8232 = ~n8216 & n8231;
  assign n8233 = n8216 & ~n8231;
  assign n8234 = ~n8232 & ~n8233;
  assign n8235 = ~n8215 & ~n8234;
  assign n8236 = n8215 & n8234;
  assign n8237 = ~n8200 & ~n8235;
  assign n8238 = ~n8236 & n8237;
  assign n8239 = ~n8200 & ~n8238;
  assign n8240 = ~n8236 & ~n8238;
  assign n8241 = ~n8235 & n8240;
  assign n8242 = ~n8239 & ~n8241;
  assign n8243 = ~n7849 & ~n7852;
  assign n8244 = n8242 & n8243;
  assign n8245 = ~n8242 & ~n8243;
  assign n8246 = ~n8244 & ~n8245;
  assign n8247 = ~n8061 & ~n8065;
  assign n8248 = ~n7843 & ~n7846;
  assign n8249 = pi10  & pi51 ;
  assign n8250 = pi15  & pi46 ;
  assign n8251 = ~n8249 & ~n8250;
  assign n8252 = pi46  & pi51 ;
  assign n8253 = n1459 & n8252;
  assign n8254 = pi16  & pi45 ;
  assign n8255 = ~n8251 & n8254;
  assign n8256 = ~n8253 & n8255;
  assign n8257 = ~n8253 & ~n8256;
  assign n8258 = ~n8251 & n8257;
  assign n8259 = n8254 & ~n8256;
  assign n8260 = ~n8258 & ~n8259;
  assign n8261 = pi11  & pi50 ;
  assign n8262 = pi47  & pi49 ;
  assign n8263 = n1644 & n8262;
  assign n8264 = pi14  & pi47 ;
  assign n8265 = pi12  & pi49 ;
  assign n8266 = ~n8264 & ~n8265;
  assign n8267 = n8261 & ~n8263;
  assign n8268 = ~n8266 & n8267;
  assign n8269 = n8261 & ~n8268;
  assign n8270 = ~n8263 & ~n8268;
  assign n8271 = ~n8266 & n8270;
  assign n8272 = ~n8269 & ~n8271;
  assign n8273 = ~n8260 & ~n8272;
  assign n8274 = ~n8260 & ~n8273;
  assign n8275 = ~n8272 & ~n8273;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = pi13  & pi48 ;
  assign n8278 = n3567 & n4908;
  assign n8279 = pi29  & pi32 ;
  assign n8280 = ~n2680 & ~n8279;
  assign n8281 = n8277 & ~n8278;
  assign n8282 = ~n8280 & n8281;
  assign n8283 = n8277 & ~n8282;
  assign n8284 = ~n8278 & ~n8282;
  assign n8285 = ~n8280 & n8284;
  assign n8286 = ~n8283 & ~n8285;
  assign n8287 = ~n8276 & ~n8286;
  assign n8288 = ~n8276 & ~n8287;
  assign n8289 = ~n8286 & ~n8287;
  assign n8290 = ~n8288 & ~n8289;
  assign n8291 = ~n7834 & ~n7839;
  assign n8292 = n8290 & n8291;
  assign n8293 = ~n8290 & ~n8291;
  assign n8294 = ~n8292 & ~n8293;
  assign n8295 = pi2  & pi59 ;
  assign n8296 = pi5  & pi56 ;
  assign n8297 = ~n8295 & ~n8296;
  assign n8298 = pi5  & pi59 ;
  assign n8299 = n7404 & n8298;
  assign n8300 = pi0  & pi61 ;
  assign n8301 = ~n8297 & n8300;
  assign n8302 = ~n8299 & n8301;
  assign n8303 = ~n8299 & ~n8302;
  assign n8304 = ~n8297 & n8303;
  assign n8305 = n8300 & ~n8302;
  assign n8306 = ~n8304 & ~n8305;
  assign n8307 = pi6  & pi55 ;
  assign n8308 = n1593 & n6012;
  assign n8309 = pi20  & pi41 ;
  assign n8310 = pi21  & pi40 ;
  assign n8311 = ~n8309 & ~n8310;
  assign n8312 = n8307 & ~n8308;
  assign n8313 = ~n8311 & n8312;
  assign n8314 = n8307 & ~n8313;
  assign n8315 = ~n8308 & ~n8313;
  assign n8316 = ~n8311 & n8315;
  assign n8317 = ~n8314 & ~n8316;
  assign n8318 = ~n8306 & ~n8317;
  assign n8319 = ~n8306 & ~n8318;
  assign n8320 = ~n8317 & ~n8318;
  assign n8321 = ~n8319 & ~n8320;
  assign n8322 = pi22  & pi39 ;
  assign n8323 = n1789 & n4500;
  assign n8324 = pi24  & pi37 ;
  assign n8325 = pi25  & pi36 ;
  assign n8326 = ~n8324 & ~n8325;
  assign n8327 = n8322 & ~n8323;
  assign n8328 = ~n8326 & n8327;
  assign n8329 = n8322 & ~n8328;
  assign n8330 = ~n8323 & ~n8328;
  assign n8331 = ~n8326 & n8330;
  assign n8332 = ~n8329 & ~n8331;
  assign n8333 = ~n8321 & ~n8332;
  assign n8334 = ~n8321 & ~n8333;
  assign n8335 = ~n8332 & ~n8333;
  assign n8336 = ~n8334 & ~n8335;
  assign n8337 = ~n8294 & n8336;
  assign n8338 = n8294 & ~n8336;
  assign n8339 = ~n8337 & ~n8338;
  assign n8340 = ~n8248 & n8339;
  assign n8341 = n8248 & ~n8339;
  assign n8342 = ~n8340 & ~n8341;
  assign n8343 = ~n8247 & n8342;
  assign n8344 = n8247 & ~n8342;
  assign n8345 = ~n8343 & ~n8344;
  assign n8346 = n8246 & n8345;
  assign n8347 = ~n8246 & ~n8345;
  assign n8348 = ~n8346 & ~n8347;
  assign n8349 = ~n8199 & n8348;
  assign n8350 = n8199 & ~n8348;
  assign n8351 = ~n8349 & ~n8350;
  assign n8352 = ~n8085 & n8351;
  assign n8353 = n8085 & ~n8351;
  assign n8354 = ~n8352 & ~n8353;
  assign n8355 = ~n8079 & ~n8083;
  assign n8356 = ~n8354 & n8355;
  assign n8357 = n8354 & ~n8355;
  assign po62  = ~n8356 & ~n8357;
  assign n8359 = ~n8196 & ~n8349;
  assign n8360 = ~n8189 & ~n8193;
  assign n8361 = n8110 & n8257;
  assign n8362 = ~n8110 & ~n8257;
  assign n8363 = ~n8361 & ~n8362;
  assign n8364 = pi3  & pi59 ;
  assign n8365 = n226 & n8144;
  assign n8366 = pi4  & pi58 ;
  assign n8367 = pi5  & pi57 ;
  assign n8368 = ~n8366 & ~n8367;
  assign n8369 = n8364 & ~n8365;
  assign n8370 = ~n8368 & n8369;
  assign n8371 = n8364 & ~n8370;
  assign n8372 = ~n8365 & ~n8370;
  assign n8373 = ~n8368 & n8372;
  assign n8374 = ~n8371 & ~n8373;
  assign n8375 = n8363 & ~n8374;
  assign n8376 = n8363 & ~n8375;
  assign n8377 = ~n8374 & ~n8375;
  assign n8378 = ~n8376 & ~n8377;
  assign n8379 = ~n8113 & ~n8127;
  assign n8380 = n8378 & n8379;
  assign n8381 = ~n8378 & ~n8379;
  assign n8382 = ~n8380 & ~n8381;
  assign n8383 = ~n8155 & ~n8159;
  assign n8384 = ~n8382 & n8383;
  assign n8385 = n8382 & ~n8383;
  assign n8386 = ~n8384 & ~n8385;
  assign n8387 = ~n8202 & ~n8206;
  assign n8388 = ~n8170 & ~n8173;
  assign n8389 = n8387 & n8388;
  assign n8390 = ~n8387 & ~n8388;
  assign n8391 = ~n8389 & ~n8390;
  assign n8392 = ~n8218 & ~n8221;
  assign n8393 = ~n8391 & n8392;
  assign n8394 = n8391 & ~n8392;
  assign n8395 = ~n8393 & ~n8394;
  assign n8396 = ~n8293 & ~n8338;
  assign n8397 = n8395 & ~n8396;
  assign n8398 = n8395 & ~n8397;
  assign n8399 = ~n8396 & ~n8397;
  assign n8400 = ~n8398 & ~n8399;
  assign n8401 = n8386 & ~n8400;
  assign n8402 = ~n8386 & n8400;
  assign n8403 = ~n8401 & ~n8402;
  assign n8404 = ~n8360 & n8403;
  assign n8405 = n8360 & ~n8403;
  assign n8406 = ~n8404 & ~n8405;
  assign n8407 = ~n8182 & ~n8186;
  assign n8408 = pi8  & pi54 ;
  assign n8409 = pi18  & pi44 ;
  assign n8410 = ~n8408 & ~n8409;
  assign n8411 = pi18  & pi54 ;
  assign n8412 = n6029 & n8411;
  assign n8413 = pi19  & pi43 ;
  assign n8414 = ~n8410 & n8413;
  assign n8415 = ~n8412 & n8414;
  assign n8416 = ~n8412 & ~n8415;
  assign n8417 = ~n8410 & n8416;
  assign n8418 = n8413 & ~n8415;
  assign n8419 = ~n8417 & ~n8418;
  assign n8420 = pi27  & pi35 ;
  assign n8421 = n2915 & n3900;
  assign n8422 = pi28  & pi34 ;
  assign n8423 = pi29  & pi33 ;
  assign n8424 = ~n8422 & ~n8423;
  assign n8425 = n8420 & ~n8421;
  assign n8426 = ~n8424 & n8425;
  assign n8427 = n8420 & ~n8426;
  assign n8428 = ~n8421 & ~n8426;
  assign n8429 = ~n8424 & n8428;
  assign n8430 = ~n8427 & ~n8429;
  assign n8431 = ~n8419 & ~n8430;
  assign n8432 = ~n8419 & ~n8431;
  assign n8433 = ~n8430 & ~n8431;
  assign n8434 = ~n8432 & ~n8433;
  assign n8435 = pi22  & pi40 ;
  assign n8436 = n2110 & n4736;
  assign n8437 = pi23  & pi39 ;
  assign n8438 = pi24  & pi38 ;
  assign n8439 = ~n8437 & ~n8438;
  assign n8440 = n8435 & ~n8436;
  assign n8441 = ~n8439 & n8440;
  assign n8442 = n8435 & ~n8441;
  assign n8443 = ~n8436 & ~n8441;
  assign n8444 = ~n8439 & n8443;
  assign n8445 = ~n8442 & ~n8444;
  assign n8446 = ~n8434 & ~n8445;
  assign n8447 = ~n8434 & ~n8446;
  assign n8448 = ~n8445 & ~n8446;
  assign n8449 = ~n8447 & ~n8448;
  assign n8450 = pi0  & pi62 ;
  assign n8451 = pi2  & pi60 ;
  assign n8452 = ~n8450 & ~n8451;
  assign n8453 = pi60  & pi62 ;
  assign n8454 = n196 & n8453;
  assign n8455 = n8167 & ~n8452;
  assign n8456 = ~n8454 & n8455;
  assign n8457 = ~n8454 & ~n8456;
  assign n8458 = ~n8452 & n8457;
  assign n8459 = n8167 & ~n8456;
  assign n8460 = ~n8458 & ~n8459;
  assign n8461 = pi21  & pi41 ;
  assign n8462 = n2310 & n4500;
  assign n8463 = pi25  & pi37 ;
  assign n8464 = pi26  & pi36 ;
  assign n8465 = ~n8463 & ~n8464;
  assign n8466 = n8461 & ~n8462;
  assign n8467 = ~n8465 & n8466;
  assign n8468 = n8461 & ~n8467;
  assign n8469 = ~n8462 & ~n8467;
  assign n8470 = ~n8465 & n8469;
  assign n8471 = ~n8468 & ~n8470;
  assign n8472 = ~n8460 & ~n8471;
  assign n8473 = ~n8460 & ~n8472;
  assign n8474 = ~n8471 & ~n8472;
  assign n8475 = ~n8473 & ~n8474;
  assign n8476 = pi9  & pi53 ;
  assign n8477 = pi45  & pi52 ;
  assign n8478 = n1747 & n8477;
  assign n8479 = pi10  & pi52 ;
  assign n8480 = pi17  & pi45 ;
  assign n8481 = ~n8479 & ~n8480;
  assign n8482 = n8476 & ~n8478;
  assign n8483 = ~n8481 & n8482;
  assign n8484 = n8476 & ~n8483;
  assign n8485 = ~n8478 & ~n8483;
  assign n8486 = ~n8481 & n8485;
  assign n8487 = ~n8484 & ~n8486;
  assign n8488 = ~n8475 & ~n8487;
  assign n8489 = ~n8475 & ~n8488;
  assign n8490 = ~n8487 & ~n8488;
  assign n8491 = ~n8489 & ~n8490;
  assign n8492 = pi11  & pi51 ;
  assign n8493 = pi15  & pi47 ;
  assign n8494 = ~n8492 & ~n8493;
  assign n8495 = pi47  & pi51 ;
  assign n8496 = n1579 & n8495;
  assign n8497 = pi16  & pi46 ;
  assign n8498 = ~n8494 & n8497;
  assign n8499 = ~n8496 & n8498;
  assign n8500 = ~n8496 & ~n8499;
  assign n8501 = ~n8494 & n8500;
  assign n8502 = n8497 & ~n8499;
  assign n8503 = ~n8501 & ~n8502;
  assign n8504 = pi12  & pi50 ;
  assign n8505 = pi48  & pi49 ;
  assign n8506 = n706 & n8505;
  assign n8507 = pi13  & pi49 ;
  assign n8508 = pi14  & pi48 ;
  assign n8509 = ~n8507 & ~n8508;
  assign n8510 = n8504 & ~n8506;
  assign n8511 = ~n8509 & n8510;
  assign n8512 = n8504 & ~n8511;
  assign n8513 = ~n8506 & ~n8511;
  assign n8514 = ~n8509 & n8513;
  assign n8515 = ~n8512 & ~n8514;
  assign n8516 = ~n8503 & ~n8515;
  assign n8517 = ~n8503 & ~n8516;
  assign n8518 = ~n8515 & ~n8516;
  assign n8519 = ~n8517 & ~n8518;
  assign n8520 = pi20  & pi42 ;
  assign n8521 = pi55  & pi56 ;
  assign n8522 = n432 & n8521;
  assign n8523 = pi6  & pi56 ;
  assign n8524 = pi7  & pi55 ;
  assign n8525 = ~n8523 & ~n8524;
  assign n8526 = n8520 & ~n8522;
  assign n8527 = ~n8525 & n8526;
  assign n8528 = n8520 & ~n8527;
  assign n8529 = ~n8522 & ~n8527;
  assign n8530 = ~n8525 & n8529;
  assign n8531 = ~n8528 & ~n8530;
  assign n8532 = ~n8519 & ~n8531;
  assign n8533 = ~n8519 & ~n8532;
  assign n8534 = ~n8531 & ~n8532;
  assign n8535 = ~n8533 & ~n8534;
  assign n8536 = ~n8491 & n8535;
  assign n8537 = n8491 & ~n8535;
  assign n8538 = ~n8536 & ~n8537;
  assign n8539 = ~n8449 & ~n8538;
  assign n8540 = n8449 & n8538;
  assign n8541 = ~n8539 & ~n8540;
  assign n8542 = ~n8407 & n8541;
  assign n8543 = ~n8407 & ~n8542;
  assign n8544 = n8541 & ~n8542;
  assign n8545 = ~n8543 & ~n8544;
  assign n8546 = ~n8240 & ~n8545;
  assign n8547 = ~n8240 & ~n8546;
  assign n8548 = ~n8545 & ~n8546;
  assign n8549 = ~n8547 & ~n8548;
  assign n8550 = ~n8406 & n8549;
  assign n8551 = n8406 & ~n8549;
  assign n8552 = ~n8550 & ~n8551;
  assign n8553 = ~n8245 & ~n8346;
  assign n8554 = ~n8224 & ~n8227;
  assign n8555 = ~n8318 & ~n8333;
  assign n8556 = n8554 & n8555;
  assign n8557 = ~n8554 & ~n8555;
  assign n8558 = ~n8556 & ~n8557;
  assign n8559 = ~n8273 & ~n8287;
  assign n8560 = ~n8558 & n8559;
  assign n8561 = n8558 & ~n8559;
  assign n8562 = ~n8560 & ~n8561;
  assign n8563 = n8303 & n8315;
  assign n8564 = ~n8303 & ~n8315;
  assign n8565 = ~n8563 & ~n8564;
  assign n8566 = n8097 & ~n8565;
  assign n8567 = ~n8097 & n8565;
  assign n8568 = ~n8566 & ~n8567;
  assign n8569 = n8124 & n8152;
  assign n8570 = ~n8124 & ~n8152;
  assign n8571 = ~n8569 & ~n8570;
  assign n8572 = n8330 & ~n8571;
  assign n8573 = ~n8330 & n8571;
  assign n8574 = ~n8572 & ~n8573;
  assign n8575 = pi1  & pi61 ;
  assign n8576 = n2332 & n8575;
  assign n8577 = ~n2332 & ~n8575;
  assign n8578 = ~n8576 & ~n8577;
  assign n8579 = n8284 & ~n8578;
  assign n8580 = ~n8284 & n8578;
  assign n8581 = ~n8579 & ~n8580;
  assign n8582 = ~n8270 & n8581;
  assign n8583 = n8270 & ~n8581;
  assign n8584 = ~n8582 & ~n8583;
  assign n8585 = n8574 & n8584;
  assign n8586 = n8574 & ~n8585;
  assign n8587 = n8584 & ~n8585;
  assign n8588 = ~n8586 & ~n8587;
  assign n8589 = n8568 & ~n8588;
  assign n8590 = n8568 & ~n8589;
  assign n8591 = ~n8588 & ~n8589;
  assign n8592 = ~n8590 & ~n8591;
  assign n8593 = n8562 & ~n8592;
  assign n8594 = n8562 & ~n8593;
  assign n8595 = ~n8592 & ~n8593;
  assign n8596 = ~n8594 & ~n8595;
  assign n8597 = ~n8132 & ~n8136;
  assign n8598 = n8596 & n8597;
  assign n8599 = ~n8596 & ~n8597;
  assign n8600 = ~n8598 & ~n8599;
  assign n8601 = ~n8230 & ~n8232;
  assign n8602 = ~n8176 & ~n8179;
  assign n8603 = n8601 & n8602;
  assign n8604 = ~n8601 & ~n8602;
  assign n8605 = ~n8603 & ~n8604;
  assign n8606 = ~n8210 & ~n8214;
  assign n8607 = ~n8605 & n8606;
  assign n8608 = n8605 & ~n8606;
  assign n8609 = ~n8607 & ~n8608;
  assign n8610 = ~n8340 & ~n8343;
  assign n8611 = ~n8609 & n8610;
  assign n8612 = n8609 & ~n8610;
  assign n8613 = ~n8611 & ~n8612;
  assign n8614 = n8600 & n8613;
  assign n8615 = ~n8600 & ~n8613;
  assign n8616 = ~n8614 & ~n8615;
  assign n8617 = ~n8553 & n8616;
  assign n8618 = ~n8553 & ~n8617;
  assign n8619 = n8616 & ~n8617;
  assign n8620 = ~n8618 & ~n8619;
  assign n8621 = n8552 & ~n8620;
  assign n8622 = ~n8552 & n8620;
  assign n8623 = ~n8621 & ~n8622;
  assign n8624 = ~n8359 & n8623;
  assign n8625 = n8359 & ~n8623;
  assign n8626 = ~n8624 & ~n8625;
  assign n8627 = ~n8352 & ~n8357;
  assign n8628 = ~n8626 & n8627;
  assign n8629 = ~n8625 & ~n8627;
  assign n8630 = ~n8624 & n8629;
  assign po63  = ~n8628 & ~n8630;
  assign n8632 = ~n8624 & ~n8629;
  assign n8633 = ~n8617 & ~n8621;
  assign n8634 = ~n8542 & ~n8546;
  assign n8635 = ~n8585 & ~n8589;
  assign n8636 = ~n8557 & ~n8561;
  assign n8637 = n8635 & n8636;
  assign n8638 = ~n8635 & ~n8636;
  assign n8639 = ~n8637 & ~n8638;
  assign n8640 = ~n8381 & ~n8385;
  assign n8641 = ~n8639 & n8640;
  assign n8642 = n8639 & ~n8640;
  assign n8643 = ~n8641 & ~n8642;
  assign n8644 = ~n8362 & ~n8375;
  assign n8645 = ~n8570 & ~n8573;
  assign n8646 = n8644 & n8645;
  assign n8647 = ~n8644 & ~n8645;
  assign n8648 = ~n8646 & ~n8647;
  assign n8649 = ~n8580 & ~n8582;
  assign n8650 = ~n8648 & n8649;
  assign n8651 = n8648 & ~n8649;
  assign n8652 = ~n8650 & ~n8651;
  assign n8653 = ~n8491 & ~n8535;
  assign n8654 = ~n8539 & ~n8653;
  assign n8655 = n8652 & ~n8654;
  assign n8656 = ~n8652 & n8654;
  assign n8657 = ~n8655 & ~n8656;
  assign n8658 = n8443 & n8529;
  assign n8659 = ~n8443 & ~n8529;
  assign n8660 = ~n8658 & ~n8659;
  assign n8661 = n8513 & ~n8660;
  assign n8662 = ~n8513 & n8660;
  assign n8663 = ~n8661 & ~n8662;
  assign n8664 = n8372 & n8469;
  assign n8665 = ~n8372 & ~n8469;
  assign n8666 = ~n8664 & ~n8665;
  assign n8667 = n8457 & ~n8666;
  assign n8668 = ~n8457 & n8666;
  assign n8669 = ~n8667 & ~n8668;
  assign n8670 = ~n8564 & ~n8567;
  assign n8671 = ~n8669 & n8670;
  assign n8672 = n8669 & ~n8670;
  assign n8673 = ~n8671 & ~n8672;
  assign n8674 = n8663 & n8673;
  assign n8675 = ~n8663 & ~n8673;
  assign n8676 = ~n8674 & ~n8675;
  assign n8677 = n8657 & n8676;
  assign n8678 = ~n8657 & ~n8676;
  assign n8679 = ~n8677 & ~n8678;
  assign n8680 = n8643 & n8679;
  assign n8681 = ~n8643 & ~n8679;
  assign n8682 = ~n8680 & ~n8681;
  assign n8683 = ~n8634 & n8682;
  assign n8684 = ~n8634 & ~n8683;
  assign n8685 = ~n8680 & ~n8683;
  assign n8686 = ~n8681 & n8685;
  assign n8687 = ~n8684 & ~n8686;
  assign n8688 = ~n8404 & ~n8551;
  assign n8689 = n8687 & n8688;
  assign n8690 = ~n8687 & ~n8688;
  assign n8691 = ~n8689 & ~n8690;
  assign n8692 = ~n8612 & ~n8614;
  assign n8693 = ~n8604 & ~n8608;
  assign n8694 = n8428 & n8485;
  assign n8695 = ~n8428 & ~n8485;
  assign n8696 = ~n8694 & ~n8695;
  assign n8697 = n8416 & ~n8696;
  assign n8698 = ~n8416 & n8696;
  assign n8699 = ~n8697 & ~n8698;
  assign n8700 = ~n8431 & ~n8446;
  assign n8701 = ~n8699 & n8700;
  assign n8702 = n8699 & ~n8700;
  assign n8703 = ~n8701 & ~n8702;
  assign n8704 = ~n8516 & ~n8532;
  assign n8705 = ~n8703 & n8704;
  assign n8706 = n8703 & ~n8704;
  assign n8707 = ~n8705 & ~n8706;
  assign n8708 = ~n8390 & ~n8394;
  assign n8709 = ~n8472 & ~n8488;
  assign n8710 = n8708 & n8709;
  assign n8711 = ~n8708 & ~n8709;
  assign n8712 = ~n8710 & ~n8711;
  assign n8713 = pi0  & pi63 ;
  assign n8714 = n8576 & n8713;
  assign n8715 = n8576 & ~n8714;
  assign n8716 = ~n8576 & n8713;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = pi62  & n2519;
  assign n8719 = pi32  & ~n8718;
  assign n8720 = pi1  & ~n8718;
  assign n8721 = pi62  & n8720;
  assign n8722 = ~n8719 & ~n8721;
  assign n8723 = ~n8717 & ~n8722;
  assign n8724 = ~n8717 & ~n8723;
  assign n8725 = ~n8722 & ~n8723;
  assign n8726 = ~n8724 & ~n8725;
  assign n8727 = pi25  & pi38 ;
  assign n8728 = pi26  & pi37 ;
  assign n8729 = ~n8727 & ~n8728;
  assign n8730 = n2310 & n5055;
  assign n8731 = pi24  & pi39 ;
  assign n8732 = ~n8729 & n8731;
  assign n8733 = ~n8730 & n8732;
  assign n8734 = ~n8730 & ~n8733;
  assign n8735 = ~n8729 & n8734;
  assign n8736 = n8731 & ~n8733;
  assign n8737 = ~n8735 & ~n8736;
  assign n8738 = pi27  & pi36 ;
  assign n8739 = n2915 & n3106;
  assign n8740 = pi28  & pi35 ;
  assign n8741 = ~n3431 & ~n8740;
  assign n8742 = n8738 & ~n8739;
  assign n8743 = ~n8741 & n8742;
  assign n8744 = n8738 & ~n8743;
  assign n8745 = ~n8739 & ~n8743;
  assign n8746 = ~n8741 & n8745;
  assign n8747 = ~n8744 & ~n8746;
  assign n8748 = ~n8737 & ~n8747;
  assign n8749 = ~n8737 & ~n8748;
  assign n8750 = ~n8747 & ~n8748;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = ~n8726 & n8751;
  assign n8753 = n8726 & ~n8751;
  assign n8754 = ~n8752 & ~n8753;
  assign n8755 = n8712 & ~n8754;
  assign n8756 = n8712 & ~n8755;
  assign n8757 = ~n8754 & ~n8755;
  assign n8758 = ~n8756 & ~n8757;
  assign n8759 = ~n8707 & n8758;
  assign n8760 = n8707 & ~n8758;
  assign n8761 = ~n8759 & ~n8760;
  assign n8762 = ~n8693 & n8761;
  assign n8763 = n8693 & ~n8761;
  assign n8764 = ~n8762 & ~n8763;
  assign n8765 = ~n8692 & n8764;
  assign n8766 = n8692 & ~n8764;
  assign n8767 = ~n8765 & ~n8766;
  assign n8768 = ~n8593 & ~n8599;
  assign n8769 = ~n8397 & ~n8401;
  assign n8770 = pi9  & pi54 ;
  assign n8771 = pi17  & pi46 ;
  assign n8772 = ~n8770 & ~n8771;
  assign n8773 = pi46  & pi54 ;
  assign n8774 = n1577 & n8773;
  assign n8775 = pi18  & pi45 ;
  assign n8776 = ~n8772 & n8775;
  assign n8777 = ~n8774 & n8776;
  assign n8778 = ~n8774 & ~n8777;
  assign n8779 = ~n8772 & n8778;
  assign n8780 = n8775 & ~n8777;
  assign n8781 = ~n8779 & ~n8780;
  assign n8782 = pi10  & pi53 ;
  assign n8783 = pi47  & pi52 ;
  assign n8784 = n1732 & n8783;
  assign n8785 = pi11  & pi52 ;
  assign n8786 = pi16  & pi47 ;
  assign n8787 = ~n8785 & ~n8786;
  assign n8788 = n8782 & ~n8784;
  assign n8789 = ~n8787 & n8788;
  assign n8790 = n8782 & ~n8789;
  assign n8791 = ~n8784 & ~n8789;
  assign n8792 = ~n8787 & n8791;
  assign n8793 = ~n8790 & ~n8792;
  assign n8794 = ~n8781 & ~n8793;
  assign n8795 = ~n8781 & ~n8794;
  assign n8796 = ~n8793 & ~n8794;
  assign n8797 = ~n8795 & ~n8796;
  assign n8798 = n952 & n6114;
  assign n8799 = pi12  & pi51 ;
  assign n8800 = pi13  & pi50 ;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = n6851 & ~n8798;
  assign n8803 = ~n8801 & n8802;
  assign n8804 = n6851 & ~n8803;
  assign n8805 = ~n8798 & ~n8803;
  assign n8806 = ~n8801 & n8805;
  assign n8807 = ~n8804 & ~n8806;
  assign n8808 = ~n8797 & ~n8807;
  assign n8809 = ~n8797 & ~n8808;
  assign n8810 = ~n8807 & ~n8808;
  assign n8811 = ~n8809 & ~n8810;
  assign n8812 = pi6  & pi57 ;
  assign n8813 = pi20  & pi43 ;
  assign n8814 = ~n8812 & ~n8813;
  assign n8815 = n8812 & n8813;
  assign n8816 = pi23  & pi40 ;
  assign n8817 = ~n8814 & n8816;
  assign n8818 = ~n8815 & n8817;
  assign n8819 = ~n8815 & ~n8818;
  assign n8820 = ~n8814 & n8819;
  assign n8821 = n8816 & ~n8818;
  assign n8822 = ~n8820 & ~n8821;
  assign n8823 = pi14  & pi49 ;
  assign n8824 = pi30  & pi33 ;
  assign n8825 = n3567 & n8824;
  assign n8826 = ~n3567 & ~n8824;
  assign n8827 = n8823 & ~n8825;
  assign n8828 = ~n8826 & n8827;
  assign n8829 = n8823 & ~n8828;
  assign n8830 = ~n8825 & ~n8828;
  assign n8831 = ~n8826 & n8830;
  assign n8832 = ~n8829 & ~n8831;
  assign n8833 = ~n8822 & ~n8832;
  assign n8834 = ~n8822 & ~n8833;
  assign n8835 = ~n8832 & ~n8833;
  assign n8836 = ~n8834 & ~n8835;
  assign n8837 = pi7  & pi56 ;
  assign n8838 = pi44  & pi55 ;
  assign n8839 = n1745 & n8838;
  assign n8840 = pi8  & pi55 ;
  assign n8841 = pi19  & pi44 ;
  assign n8842 = ~n8840 & ~n8841;
  assign n8843 = n8837 & ~n8839;
  assign n8844 = ~n8842 & n8843;
  assign n8845 = n8837 & ~n8844;
  assign n8846 = ~n8839 & ~n8844;
  assign n8847 = ~n8842 & n8846;
  assign n8848 = ~n8845 & ~n8847;
  assign n8849 = ~n8836 & ~n8848;
  assign n8850 = ~n8836 & ~n8849;
  assign n8851 = ~n8848 & ~n8849;
  assign n8852 = ~n8850 & ~n8851;
  assign n8853 = pi2  & pi61 ;
  assign n8854 = pi59  & pi60 ;
  assign n8855 = n209 & n8854;
  assign n8856 = pi3  & pi60 ;
  assign n8857 = pi4  & pi59 ;
  assign n8858 = ~n8856 & ~n8857;
  assign n8859 = n8853 & ~n8855;
  assign n8860 = ~n8858 & n8859;
  assign n8861 = n8853 & ~n8860;
  assign n8862 = ~n8855 & ~n8860;
  assign n8863 = ~n8858 & n8862;
  assign n8864 = ~n8861 & ~n8863;
  assign n8865 = n8500 & ~n8864;
  assign n8866 = ~n8500 & n8864;
  assign n8867 = ~n8865 & ~n8866;
  assign n8868 = pi5  & pi58 ;
  assign n8869 = n1481 & n5235;
  assign n8870 = pi21  & pi42 ;
  assign n8871 = pi22  & pi41 ;
  assign n8872 = ~n8870 & ~n8871;
  assign n8873 = n8868 & ~n8869;
  assign n8874 = ~n8872 & n8873;
  assign n8875 = n8868 & ~n8874;
  assign n8876 = ~n8869 & ~n8874;
  assign n8877 = ~n8872 & n8876;
  assign n8878 = ~n8875 & ~n8877;
  assign n8879 = ~n8867 & ~n8878;
  assign n8880 = n8867 & n8878;
  assign n8881 = ~n8879 & ~n8880;
  assign n8882 = n8852 & n8881;
  assign n8883 = ~n8852 & ~n8881;
  assign n8884 = ~n8882 & ~n8883;
  assign n8885 = ~n8811 & ~n8884;
  assign n8886 = n8811 & n8884;
  assign n8887 = ~n8885 & ~n8886;
  assign n8888 = ~n8769 & n8887;
  assign n8889 = ~n8769 & ~n8888;
  assign n8890 = n8887 & ~n8888;
  assign n8891 = ~n8889 & ~n8890;
  assign n8892 = ~n8768 & ~n8891;
  assign n8893 = ~n8768 & ~n8892;
  assign n8894 = ~n8891 & ~n8892;
  assign n8895 = ~n8893 & ~n8894;
  assign n8896 = n8767 & ~n8895;
  assign n8897 = n8767 & ~n8896;
  assign n8898 = ~n8895 & ~n8896;
  assign n8899 = ~n8897 & ~n8898;
  assign n8900 = ~n8691 & n8899;
  assign n8901 = n8691 & ~n8899;
  assign n8902 = ~n8900 & ~n8901;
  assign n8903 = n8633 & ~n8902;
  assign n8904 = ~n8633 & n8902;
  assign n8905 = ~n8903 & ~n8904;
  assign n8906 = ~n8632 & ~n8905;
  assign n8907 = n8632 & n8905;
  assign po64  = n8906 | n8907;
  assign n8909 = ~n8632 & ~n8903;
  assign n8910 = ~n8904 & ~n8909;
  assign n8911 = ~n8765 & ~n8896;
  assign n8912 = ~n8888 & ~n8892;
  assign n8913 = ~n8760 & ~n8762;
  assign n8914 = ~n8852 & n8881;
  assign n8915 = ~n8885 & ~n8914;
  assign n8916 = ~n8711 & ~n8755;
  assign n8917 = n8915 & n8916;
  assign n8918 = ~n8915 & ~n8916;
  assign n8919 = ~n8917 & ~n8918;
  assign n8920 = ~n8726 & ~n8751;
  assign n8921 = ~n8748 & ~n8920;
  assign n8922 = n8778 & n8819;
  assign n8923 = ~n8778 & ~n8819;
  assign n8924 = ~n8922 & ~n8923;
  assign n8925 = n8745 & ~n8924;
  assign n8926 = ~n8745 & n8924;
  assign n8927 = ~n8925 & ~n8926;
  assign n8928 = n8862 & n8876;
  assign n8929 = ~n8862 & ~n8876;
  assign n8930 = ~n8928 & ~n8929;
  assign n8931 = n8846 & ~n8930;
  assign n8932 = ~n8846 & n8930;
  assign n8933 = ~n8931 & ~n8932;
  assign n8934 = ~n8927 & ~n8933;
  assign n8935 = n8927 & n8933;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = ~n8921 & n8936;
  assign n8938 = n8921 & ~n8936;
  assign n8939 = ~n8937 & ~n8938;
  assign n8940 = ~n8919 & ~n8939;
  assign n8941 = n8919 & n8939;
  assign n8942 = ~n8940 & ~n8941;
  assign n8943 = ~n8913 & n8942;
  assign n8944 = ~n8913 & ~n8943;
  assign n8945 = n8942 & ~n8943;
  assign n8946 = ~n8944 & ~n8945;
  assign n8947 = ~n8912 & ~n8946;
  assign n8948 = ~n8912 & ~n8947;
  assign n8949 = ~n8946 & ~n8947;
  assign n8950 = ~n8948 & ~n8949;
  assign n8951 = ~n8911 & ~n8950;
  assign n8952 = ~n8911 & ~n8951;
  assign n8953 = ~n8950 & ~n8951;
  assign n8954 = ~n8952 & ~n8953;
  assign n8955 = ~n8655 & ~n8677;
  assign n8956 = pi17  & pi47 ;
  assign n8957 = pi7  & pi57 ;
  assign n8958 = ~n8956 & ~n8957;
  assign n8959 = pi17  & pi57 ;
  assign n8960 = n6504 & n8959;
  assign n8961 = pi6  & pi58 ;
  assign n8962 = ~n8958 & n8961;
  assign n8963 = ~n8960 & n8962;
  assign n8964 = ~n8960 & ~n8963;
  assign n8965 = ~n8958 & n8964;
  assign n8966 = n8961 & ~n8963;
  assign n8967 = ~n8965 & ~n8966;
  assign n8968 = pi20  & pi44 ;
  assign n8969 = n1481 & n6458;
  assign n8970 = pi21  & pi43 ;
  assign n8971 = pi22  & pi42 ;
  assign n8972 = ~n8970 & ~n8971;
  assign n8973 = n8968 & ~n8969;
  assign n8974 = ~n8972 & n8973;
  assign n8975 = n8968 & ~n8974;
  assign n8976 = ~n8969 & ~n8974;
  assign n8977 = ~n8972 & n8976;
  assign n8978 = ~n8975 & ~n8977;
  assign n8979 = ~n8967 & ~n8978;
  assign n8980 = ~n8967 & ~n8979;
  assign n8981 = ~n8978 & ~n8979;
  assign n8982 = ~n8980 & ~n8981;
  assign n8983 = pi23  & pi41 ;
  assign n8984 = n1789 & n5548;
  assign n8985 = pi24  & pi40 ;
  assign n8986 = pi25  & pi39 ;
  assign n8987 = ~n8985 & ~n8986;
  assign n8988 = n8983 & ~n8984;
  assign n8989 = ~n8987 & n8988;
  assign n8990 = n8983 & ~n8989;
  assign n8991 = ~n8984 & ~n8989;
  assign n8992 = ~n8987 & n8991;
  assign n8993 = ~n8990 & ~n8992;
  assign n8994 = ~n8982 & ~n8993;
  assign n8995 = ~n8982 & ~n8994;
  assign n8996 = ~n8993 & ~n8994;
  assign n8997 = ~n8995 & ~n8996;
  assign n8998 = pi8  & pi56 ;
  assign n8999 = ~n6185 & ~n8998;
  assign n9000 = pi48  & pi56 ;
  assign n9001 = n1421 & n9000;
  assign n9002 = pi26  & pi38 ;
  assign n9003 = ~n8999 & n9002;
  assign n9004 = ~n9001 & n9003;
  assign n9005 = ~n9001 & ~n9004;
  assign n9006 = ~n8999 & n9005;
  assign n9007 = n9002 & ~n9004;
  assign n9008 = ~n9006 & ~n9007;
  assign n9009 = pi27  & pi37 ;
  assign n9010 = n2915 & n4691;
  assign n9011 = pi28  & pi36 ;
  assign n9012 = pi29  & pi35 ;
  assign n9013 = ~n9011 & ~n9012;
  assign n9014 = n9009 & ~n9010;
  assign n9015 = ~n9013 & n9014;
  assign n9016 = n9009 & ~n9015;
  assign n9017 = ~n9010 & ~n9015;
  assign n9018 = ~n9013 & n9017;
  assign n9019 = ~n9016 & ~n9018;
  assign n9020 = ~n9008 & ~n9019;
  assign n9021 = ~n9008 & ~n9020;
  assign n9022 = ~n9019 & ~n9020;
  assign n9023 = ~n9021 & ~n9022;
  assign n9024 = pi14  & pi50 ;
  assign n9025 = n2680 & n3900;
  assign n9026 = pi31  & pi33 ;
  assign n9027 = pi30  & pi34 ;
  assign n9028 = ~n9026 & ~n9027;
  assign n9029 = n9024 & ~n9025;
  assign n9030 = ~n9028 & n9029;
  assign n9031 = n9024 & ~n9030;
  assign n9032 = ~n9025 & ~n9030;
  assign n9033 = ~n9028 & n9032;
  assign n9034 = ~n9031 & ~n9033;
  assign n9035 = ~n9023 & ~n9034;
  assign n9036 = ~n9023 & ~n9035;
  assign n9037 = ~n9034 & ~n9035;
  assign n9038 = ~n9036 & ~n9037;
  assign n9039 = pi18  & pi46 ;
  assign n9040 = pi19  & pi45 ;
  assign n9041 = ~n9039 & ~n9040;
  assign n9042 = n1085 & n7513;
  assign n9043 = n8298 & ~n9041;
  assign n9044 = ~n9042 & n9043;
  assign n9045 = n8298 & ~n9044;
  assign n9046 = ~n9042 & ~n9044;
  assign n9047 = ~n9041 & n9046;
  assign n9048 = ~n9045 & ~n9047;
  assign n9049 = ~n8714 & ~n8723;
  assign n9050 = ~n9048 & n9049;
  assign n9051 = n9048 & ~n9049;
  assign n9052 = ~n9050 & ~n9051;
  assign n9053 = pi2  & pi62 ;
  assign n9054 = pi60  & pi61 ;
  assign n9055 = n209 & n9054;
  assign n9056 = pi3  & pi61 ;
  assign n9057 = pi4  & pi60 ;
  assign n9058 = ~n9056 & ~n9057;
  assign n9059 = n9053 & ~n9055;
  assign n9060 = ~n9058 & n9059;
  assign n9061 = n9053 & ~n9060;
  assign n9062 = ~n9055 & ~n9060;
  assign n9063 = ~n9058 & n9062;
  assign n9064 = ~n9061 & ~n9063;
  assign n9065 = ~n9052 & ~n9064;
  assign n9066 = n9052 & n9064;
  assign n9067 = ~n9065 & ~n9066;
  assign n9068 = n9038 & n9067;
  assign n9069 = ~n9038 & ~n9067;
  assign n9070 = ~n9068 & ~n9069;
  assign n9071 = ~n8997 & ~n9070;
  assign n9072 = n8997 & n9070;
  assign n9073 = ~n9071 & ~n9072;
  assign n9074 = ~n8955 & n9073;
  assign n9075 = n8955 & ~n9073;
  assign n9076 = ~n9074 & ~n9075;
  assign n9077 = ~n8659 & ~n8662;
  assign n9078 = ~n8695 & ~n8698;
  assign n9079 = n9077 & n9078;
  assign n9080 = ~n9077 & ~n9078;
  assign n9081 = ~n9079 & ~n9080;
  assign n9082 = ~n8665 & ~n8668;
  assign n9083 = ~n9081 & n9082;
  assign n9084 = n9081 & ~n9082;
  assign n9085 = ~n9083 & ~n9084;
  assign n9086 = ~n8702 & ~n8706;
  assign n9087 = ~n8672 & ~n8674;
  assign n9088 = ~n9086 & ~n9087;
  assign n9089 = ~n9086 & ~n9088;
  assign n9090 = ~n9087 & ~n9088;
  assign n9091 = ~n9089 & ~n9090;
  assign n9092 = n9085 & ~n9091;
  assign n9093 = ~n9085 & n9091;
  assign n9094 = ~n9092 & ~n9093;
  assign n9095 = n9076 & n9094;
  assign n9096 = n9076 & ~n9095;
  assign n9097 = n9094 & ~n9095;
  assign n9098 = ~n9096 & ~n9097;
  assign n9099 = n8734 & n8805;
  assign n9100 = ~n8734 & ~n8805;
  assign n9101 = ~n9099 & ~n9100;
  assign n9102 = n8791 & ~n9101;
  assign n9103 = ~n8791 & n9101;
  assign n9104 = ~n9102 & ~n9103;
  assign n9105 = ~n8833 & ~n8849;
  assign n9106 = ~n9104 & n9105;
  assign n9107 = n9104 & ~n9105;
  assign n9108 = ~n9106 & ~n9107;
  assign n9109 = ~n8794 & ~n8808;
  assign n9110 = ~n9108 & n9109;
  assign n9111 = n9108 & ~n9109;
  assign n9112 = ~n9110 & ~n9111;
  assign n9113 = ~n8638 & ~n8642;
  assign n9114 = ~n9112 & n9113;
  assign n9115 = n9112 & ~n9113;
  assign n9116 = ~n9114 & ~n9115;
  assign n9117 = ~n8647 & ~n8651;
  assign n9118 = ~n8500 & ~n8864;
  assign n9119 = ~n8879 & ~n9118;
  assign n9120 = n9117 & n9119;
  assign n9121 = ~n9117 & ~n9119;
  assign n9122 = ~n9120 & ~n9121;
  assign n9123 = pi62  & pi63 ;
  assign n9124 = n2519 & n9123;
  assign n9125 = n8718 & ~n9124;
  assign n9126 = pi63  & n8720;
  assign n9127 = ~n9125 & ~n9126;
  assign n9128 = ~n8830 & ~n9127;
  assign n9129 = ~n8830 & ~n9128;
  assign n9130 = ~n9127 & ~n9128;
  assign n9131 = ~n9129 & ~n9130;
  assign n9132 = pi10  & pi54 ;
  assign n9133 = pi15  & pi49 ;
  assign n9134 = ~n9132 & ~n9133;
  assign n9135 = n9132 & n9133;
  assign n9136 = pi9  & pi55 ;
  assign n9137 = ~n9134 & n9136;
  assign n9138 = ~n9135 & n9137;
  assign n9139 = ~n9135 & ~n9138;
  assign n9140 = ~n9134 & n9139;
  assign n9141 = n9136 & ~n9138;
  assign n9142 = ~n9140 & ~n9141;
  assign n9143 = pi13  & pi51 ;
  assign n9144 = pi52  & pi53 ;
  assign n9145 = n579 & n9144;
  assign n9146 = pi11  & pi53 ;
  assign n9147 = pi12  & pi52 ;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = n9143 & ~n9145;
  assign n9150 = ~n9148 & n9149;
  assign n9151 = n9143 & ~n9150;
  assign n9152 = ~n9145 & ~n9150;
  assign n9153 = ~n9148 & n9152;
  assign n9154 = ~n9151 & ~n9153;
  assign n9155 = ~n9142 & ~n9154;
  assign n9156 = ~n9142 & ~n9155;
  assign n9157 = ~n9154 & ~n9155;
  assign n9158 = ~n9156 & ~n9157;
  assign n9159 = ~n9131 & n9158;
  assign n9160 = n9131 & ~n9158;
  assign n9161 = ~n9159 & ~n9160;
  assign n9162 = n9122 & ~n9161;
  assign n9163 = n9122 & ~n9162;
  assign n9164 = ~n9161 & ~n9162;
  assign n9165 = ~n9163 & ~n9164;
  assign n9166 = ~n9116 & n9165;
  assign n9167 = n9116 & ~n9165;
  assign n9168 = ~n9166 & ~n9167;
  assign n9169 = ~n8685 & n9168;
  assign n9170 = n8685 & ~n9168;
  assign n9171 = ~n9169 & ~n9170;
  assign n9172 = ~n9098 & n9171;
  assign n9173 = n9098 & ~n9171;
  assign n9174 = ~n9172 & ~n9173;
  assign n9175 = ~n8954 & n9174;
  assign n9176 = n8954 & ~n9174;
  assign n9177 = ~n9175 & ~n9176;
  assign n9178 = ~n8690 & ~n8901;
  assign n9179 = ~n9177 & n9178;
  assign n9180 = n9177 & ~n9178;
  assign n9181 = ~n9179 & ~n9180;
  assign n9182 = n8910 & ~n9181;
  assign n9183 = ~n8910 & ~n9179;
  assign n9184 = ~n9180 & n9183;
  assign po65  = ~n9182 & ~n9184;
  assign n9186 = ~n9180 & ~n9183;
  assign n9187 = ~n8951 & ~n9175;
  assign n9188 = ~n9169 & ~n9172;
  assign n9189 = ~n9074 & ~n9095;
  assign n9190 = ~n9115 & ~n9167;
  assign n9191 = ~n9038 & n9067;
  assign n9192 = ~n9071 & ~n9191;
  assign n9193 = ~n9121 & ~n9162;
  assign n9194 = n9192 & n9193;
  assign n9195 = ~n9192 & ~n9193;
  assign n9196 = ~n9194 & ~n9195;
  assign n9197 = ~n9131 & ~n9158;
  assign n9198 = ~n9155 & ~n9197;
  assign n9199 = n8991 & n9139;
  assign n9200 = ~n8991 & ~n9139;
  assign n9201 = ~n9199 & ~n9200;
  assign n9202 = n8964 & ~n9201;
  assign n9203 = ~n8964 & n9201;
  assign n9204 = ~n9202 & ~n9203;
  assign n9205 = n9046 & n9062;
  assign n9206 = ~n9046 & ~n9062;
  assign n9207 = ~n9205 & ~n9206;
  assign n9208 = n9005 & ~n9207;
  assign n9209 = ~n9005 & n9207;
  assign n9210 = ~n9208 & ~n9209;
  assign n9211 = ~n9204 & ~n9210;
  assign n9212 = n9204 & n9210;
  assign n9213 = ~n9211 & ~n9212;
  assign n9214 = ~n9198 & n9213;
  assign n9215 = n9198 & ~n9213;
  assign n9216 = ~n9214 & ~n9215;
  assign n9217 = ~n9196 & ~n9216;
  assign n9218 = n9196 & n9216;
  assign n9219 = ~n9217 & ~n9218;
  assign n9220 = ~n9190 & n9219;
  assign n9221 = n9190 & ~n9219;
  assign n9222 = ~n9220 & ~n9221;
  assign n9223 = ~n9189 & n9222;
  assign n9224 = n9189 & ~n9222;
  assign n9225 = ~n9223 & ~n9224;
  assign n9226 = n9188 & ~n9225;
  assign n9227 = ~n9188 & n9225;
  assign n9228 = ~n9226 & ~n9227;
  assign n9229 = ~n8943 & ~n8947;
  assign n9230 = ~n9080 & ~n9084;
  assign n9231 = ~n9048 & ~n9049;
  assign n9232 = ~n9065 & ~n9231;
  assign n9233 = n9230 & n9232;
  assign n9234 = ~n9230 & ~n9232;
  assign n9235 = ~n9233 & ~n9234;
  assign n9236 = pi61  & pi63 ;
  assign n9237 = n249 & n9236;
  assign n9238 = pi4  & pi61 ;
  assign n9239 = ~n9237 & n9238;
  assign n9240 = pi2  & pi63 ;
  assign n9241 = ~n9237 & n9240;
  assign n9242 = ~n9239 & ~n9241;
  assign n9243 = ~n9032 & ~n9242;
  assign n9244 = ~n9032 & ~n9243;
  assign n9245 = ~n9242 & ~n9243;
  assign n9246 = ~n9244 & ~n9245;
  assign n9247 = pi13  & pi52 ;
  assign n9248 = pi18  & pi47 ;
  assign n9249 = ~n9247 & ~n9248;
  assign n9250 = n9247 & n9248;
  assign n9251 = pi12  & pi53 ;
  assign n9252 = ~n9249 & n9251;
  assign n9253 = ~n9250 & n9252;
  assign n9254 = ~n9250 & ~n9253;
  assign n9255 = ~n9249 & n9254;
  assign n9256 = n9251 & ~n9253;
  assign n9257 = ~n9255 & ~n9256;
  assign n9258 = n1041 & n6114;
  assign n9259 = pi14  & pi51 ;
  assign n9260 = pi15  & pi50 ;
  assign n9261 = ~n9259 & ~n9260;
  assign n9262 = n7122 & ~n9258;
  assign n9263 = ~n9261 & n9262;
  assign n9264 = n7122 & ~n9263;
  assign n9265 = ~n9258 & ~n9263;
  assign n9266 = ~n9261 & n9265;
  assign n9267 = ~n9264 & ~n9266;
  assign n9268 = ~n9257 & ~n9267;
  assign n9269 = ~n9257 & ~n9268;
  assign n9270 = ~n9267 & ~n9268;
  assign n9271 = ~n9269 & ~n9270;
  assign n9272 = ~n9246 & n9271;
  assign n9273 = n9246 & ~n9271;
  assign n9274 = ~n9272 & ~n9273;
  assign n9275 = n9235 & ~n9274;
  assign n9276 = n9235 & ~n9275;
  assign n9277 = ~n9274 & ~n9275;
  assign n9278 = ~n9276 & ~n9277;
  assign n9279 = n8976 & n9017;
  assign n9280 = ~n8976 & ~n9017;
  assign n9281 = ~n9279 & ~n9280;
  assign n9282 = n9152 & ~n9281;
  assign n9283 = ~n9152 & n9281;
  assign n9284 = ~n9282 & ~n9283;
  assign n9285 = ~n9020 & ~n9035;
  assign n9286 = ~n9284 & n9285;
  assign n9287 = n9284 & ~n9285;
  assign n9288 = ~n9286 & ~n9287;
  assign n9289 = ~n8979 & ~n8994;
  assign n9290 = ~n9288 & n9289;
  assign n9291 = n9288 & ~n9289;
  assign n9292 = ~n9290 & ~n9291;
  assign n9293 = ~n9088 & ~n9092;
  assign n9294 = n9292 & ~n9293;
  assign n9295 = n9292 & ~n9294;
  assign n9296 = ~n9293 & ~n9294;
  assign n9297 = ~n9295 & ~n9296;
  assign n9298 = ~n9278 & ~n9297;
  assign n9299 = ~n9278 & ~n9298;
  assign n9300 = ~n9297 & ~n9298;
  assign n9301 = ~n9299 & ~n9300;
  assign n9302 = ~n9229 & ~n9301;
  assign n9303 = ~n9229 & ~n9302;
  assign n9304 = ~n9301 & ~n9302;
  assign n9305 = ~n9303 & ~n9304;
  assign n9306 = ~n8918 & ~n8941;
  assign n9307 = pi10  & pi55 ;
  assign n9308 = pi20  & pi45 ;
  assign n9309 = ~n9307 & ~n9308;
  assign n9310 = n9307 & n9308;
  assign n9311 = pi9  & pi56 ;
  assign n9312 = ~n9309 & n9311;
  assign n9313 = ~n9310 & n9312;
  assign n9314 = ~n9310 & ~n9313;
  assign n9315 = ~n9309 & n9314;
  assign n9316 = n9311 & ~n9313;
  assign n9317 = ~n9315 & ~n9316;
  assign n9318 = pi23  & pi42 ;
  assign n9319 = n1789 & n6012;
  assign n9320 = pi24  & pi41 ;
  assign n9321 = pi25  & pi40 ;
  assign n9322 = ~n9320 & ~n9321;
  assign n9323 = n9318 & ~n9319;
  assign n9324 = ~n9322 & n9323;
  assign n9325 = n9318 & ~n9324;
  assign n9326 = ~n9319 & ~n9324;
  assign n9327 = ~n9322 & n9326;
  assign n9328 = ~n9325 & ~n9327;
  assign n9329 = ~n9317 & ~n9328;
  assign n9330 = ~n9317 & ~n9329;
  assign n9331 = ~n9328 & ~n9329;
  assign n9332 = ~n9330 & ~n9331;
  assign n9333 = pi26  & pi39 ;
  assign n9334 = n2191 & n5055;
  assign n9335 = pi27  & pi38 ;
  assign n9336 = pi28  & pi37 ;
  assign n9337 = ~n9335 & ~n9336;
  assign n9338 = n9333 & ~n9334;
  assign n9339 = ~n9337 & n9338;
  assign n9340 = n9333 & ~n9339;
  assign n9341 = ~n9334 & ~n9339;
  assign n9342 = ~n9337 & n9341;
  assign n9343 = ~n9340 & ~n9342;
  assign n9344 = ~n9332 & ~n9343;
  assign n9345 = ~n9332 & ~n9344;
  assign n9346 = ~n9343 & ~n9344;
  assign n9347 = ~n9345 & ~n9346;
  assign n9348 = pi11  & pi54 ;
  assign n9349 = pi19  & pi46 ;
  assign n9350 = ~n9348 & ~n9349;
  assign n9351 = n9348 & n9349;
  assign n9352 = pi29  & pi36 ;
  assign n9353 = ~n9350 & n9352;
  assign n9354 = ~n9351 & n9353;
  assign n9355 = ~n9351 & ~n9354;
  assign n9356 = ~n9350 & n9355;
  assign n9357 = n9352 & ~n9354;
  assign n9358 = ~n9356 & ~n9357;
  assign n9359 = n3567 & n3900;
  assign n9360 = pi31  & pi34 ;
  assign n9361 = ~n6138 & ~n9360;
  assign n9362 = n3769 & ~n9359;
  assign n9363 = ~n9361 & n9362;
  assign n9364 = n3769 & ~n9363;
  assign n9365 = ~n9359 & ~n9363;
  assign n9366 = ~n9361 & n9365;
  assign n9367 = ~n9364 & ~n9366;
  assign n9368 = ~n9358 & ~n9367;
  assign n9369 = ~n9358 & ~n9368;
  assign n9370 = ~n9367 & ~n9368;
  assign n9371 = ~n9369 & ~n9370;
  assign n9372 = pi17  & pi48 ;
  assign n9373 = pi3  & pi62 ;
  assign n9374 = pi33  & n9373;
  assign n9375 = ~pi33  & ~n9373;
  assign n9376 = n9372 & ~n9374;
  assign n9377 = ~n9375 & n9376;
  assign n9378 = n9372 & ~n9377;
  assign n9379 = ~n9374 & ~n9377;
  assign n9380 = ~n9375 & n9379;
  assign n9381 = ~n9378 & ~n9380;
  assign n9382 = ~n9371 & ~n9381;
  assign n9383 = ~n9371 & ~n9382;
  assign n9384 = ~n9381 & ~n9382;
  assign n9385 = ~n9383 & ~n9384;
  assign n9386 = pi8  & pi57 ;
  assign n9387 = n1481 & n6836;
  assign n9388 = pi21  & pi44 ;
  assign n9389 = pi22  & pi43 ;
  assign n9390 = ~n9388 & ~n9389;
  assign n9391 = n9386 & ~n9387;
  assign n9392 = ~n9390 & n9391;
  assign n9393 = n9386 & ~n9392;
  assign n9394 = ~n9387 & ~n9392;
  assign n9395 = ~n9390 & n9394;
  assign n9396 = ~n9393 & ~n9395;
  assign n9397 = ~n9124 & ~n9128;
  assign n9398 = ~n9396 & n9397;
  assign n9399 = n9396 & ~n9397;
  assign n9400 = ~n9398 & ~n9399;
  assign n9401 = pi5  & pi60 ;
  assign n9402 = pi58  & pi59 ;
  assign n9403 = n432 & n9402;
  assign n9404 = pi6  & pi59 ;
  assign n9405 = pi7  & pi58 ;
  assign n9406 = ~n9404 & ~n9405;
  assign n9407 = n9401 & ~n9403;
  assign n9408 = ~n9406 & n9407;
  assign n9409 = n9401 & ~n9408;
  assign n9410 = ~n9403 & ~n9408;
  assign n9411 = ~n9406 & n9410;
  assign n9412 = ~n9409 & ~n9411;
  assign n9413 = ~n9400 & ~n9412;
  assign n9414 = n9400 & n9412;
  assign n9415 = ~n9413 & ~n9414;
  assign n9416 = n9385 & n9415;
  assign n9417 = ~n9385 & ~n9415;
  assign n9418 = ~n9416 & ~n9417;
  assign n9419 = ~n9347 & ~n9418;
  assign n9420 = ~n9347 & ~n9419;
  assign n9421 = ~n9418 & ~n9419;
  assign n9422 = ~n9420 & ~n9421;
  assign n9423 = ~n9306 & ~n9422;
  assign n9424 = ~n9306 & ~n9423;
  assign n9425 = ~n9422 & ~n9423;
  assign n9426 = ~n9424 & ~n9425;
  assign n9427 = ~n9100 & ~n9103;
  assign n9428 = ~n8923 & ~n8926;
  assign n9429 = n9427 & n9428;
  assign n9430 = ~n9427 & ~n9428;
  assign n9431 = ~n9429 & ~n9430;
  assign n9432 = ~n8929 & ~n8932;
  assign n9433 = ~n9431 & n9432;
  assign n9434 = n9431 & ~n9432;
  assign n9435 = ~n9433 & ~n9434;
  assign n9436 = ~n8935 & ~n8937;
  assign n9437 = ~n9107 & ~n9111;
  assign n9438 = ~n9436 & n9437;
  assign n9439 = n9436 & ~n9437;
  assign n9440 = ~n9438 & ~n9439;
  assign n9441 = n9435 & ~n9440;
  assign n9442 = ~n9435 & n9440;
  assign n9443 = ~n9441 & ~n9442;
  assign n9444 = ~n9426 & n9443;
  assign n9445 = ~n9426 & ~n9444;
  assign n9446 = n9443 & ~n9444;
  assign n9447 = ~n9445 & ~n9446;
  assign n9448 = ~n9305 & n9447;
  assign n9449 = n9305 & ~n9447;
  assign n9450 = ~n9448 & ~n9449;
  assign n9451 = n9228 & ~n9450;
  assign n9452 = ~n9228 & n9450;
  assign n9453 = ~n9451 & ~n9452;
  assign n9454 = ~n9187 & n9453;
  assign n9455 = n9187 & ~n9453;
  assign n9456 = ~n9454 & ~n9455;
  assign n9457 = ~n9186 & ~n9456;
  assign n9458 = n9186 & n9456;
  assign po66  = n9457 | n9458;
  assign n9460 = ~n9186 & ~n9455;
  assign n9461 = ~n9454 & ~n9460;
  assign n9462 = ~n9227 & ~n9451;
  assign n9463 = ~n9305 & ~n9447;
  assign n9464 = ~n9302 & ~n9463;
  assign n9465 = ~n9436 & ~n9437;
  assign n9466 = ~n9441 & ~n9465;
  assign n9467 = ~n9237 & ~n9243;
  assign n9468 = n9341 & n9467;
  assign n9469 = ~n9341 & ~n9467;
  assign n9470 = ~n9468 & ~n9469;
  assign n9471 = pi6  & pi60 ;
  assign n9472 = n521 & n9402;
  assign n9473 = pi7  & pi59 ;
  assign n9474 = pi8  & pi58 ;
  assign n9475 = ~n9473 & ~n9474;
  assign n9476 = n9471 & ~n9472;
  assign n9477 = ~n9475 & n9476;
  assign n9478 = n9471 & ~n9477;
  assign n9479 = ~n9472 & ~n9477;
  assign n9480 = ~n9475 & n9479;
  assign n9481 = ~n9478 & ~n9480;
  assign n9482 = n9470 & ~n9481;
  assign n9483 = n9470 & ~n9482;
  assign n9484 = ~n9481 & ~n9482;
  assign n9485 = ~n9483 & ~n9484;
  assign n9486 = ~n9246 & ~n9271;
  assign n9487 = ~n9268 & ~n9486;
  assign n9488 = ~n9485 & ~n9487;
  assign n9489 = ~n9485 & ~n9488;
  assign n9490 = ~n9487 & ~n9488;
  assign n9491 = ~n9489 & ~n9490;
  assign n9492 = ~n9430 & ~n9434;
  assign n9493 = n9491 & n9492;
  assign n9494 = ~n9491 & ~n9492;
  assign n9495 = ~n9493 & ~n9494;
  assign n9496 = n9365 & n9379;
  assign n9497 = ~n9365 & ~n9379;
  assign n9498 = ~n9496 & ~n9497;
  assign n9499 = n9265 & ~n9498;
  assign n9500 = ~n9265 & n9498;
  assign n9501 = ~n9499 & ~n9500;
  assign n9502 = n9394 & n9410;
  assign n9503 = ~n9394 & ~n9410;
  assign n9504 = ~n9502 & ~n9503;
  assign n9505 = n9355 & ~n9504;
  assign n9506 = ~n9355 & n9504;
  assign n9507 = ~n9505 & ~n9506;
  assign n9508 = ~n9368 & ~n9382;
  assign n9509 = ~n9507 & n9508;
  assign n9510 = n9507 & ~n9508;
  assign n9511 = ~n9509 & ~n9510;
  assign n9512 = n9501 & n9511;
  assign n9513 = ~n9501 & ~n9511;
  assign n9514 = ~n9512 & ~n9513;
  assign n9515 = n9495 & n9514;
  assign n9516 = ~n9495 & ~n9514;
  assign n9517 = ~n9515 & ~n9516;
  assign n9518 = ~n9466 & n9517;
  assign n9519 = n9466 & ~n9517;
  assign n9520 = ~n9518 & ~n9519;
  assign n9521 = ~n9294 & ~n9298;
  assign n9522 = n9254 & n9314;
  assign n9523 = ~n9254 & ~n9314;
  assign n9524 = ~n9522 & ~n9523;
  assign n9525 = n9326 & ~n9524;
  assign n9526 = ~n9326 & n9524;
  assign n9527 = ~n9525 & ~n9526;
  assign n9528 = ~n9396 & ~n9397;
  assign n9529 = ~n9413 & ~n9528;
  assign n9530 = ~n9527 & n9529;
  assign n9531 = n9527 & ~n9529;
  assign n9532 = ~n9530 & ~n9531;
  assign n9533 = ~n9329 & ~n9344;
  assign n9534 = ~n9532 & n9533;
  assign n9535 = n9532 & ~n9533;
  assign n9536 = ~n9534 & ~n9535;
  assign n9537 = ~n9385 & n9415;
  assign n9538 = ~n9419 & ~n9537;
  assign n9539 = ~n9234 & ~n9275;
  assign n9540 = n9538 & n9539;
  assign n9541 = ~n9538 & ~n9539;
  assign n9542 = ~n9540 & ~n9541;
  assign n9543 = n9536 & n9542;
  assign n9544 = ~n9536 & ~n9542;
  assign n9545 = ~n9543 & ~n9544;
  assign n9546 = ~n9521 & n9545;
  assign n9547 = ~n9521 & ~n9546;
  assign n9548 = n9545 & ~n9546;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = n9520 & ~n9549;
  assign n9551 = n9520 & ~n9550;
  assign n9552 = ~n9549 & ~n9550;
  assign n9553 = ~n9551 & ~n9552;
  assign n9554 = ~n9464 & ~n9553;
  assign n9555 = ~n9464 & ~n9554;
  assign n9556 = ~n9553 & ~n9554;
  assign n9557 = ~n9555 & ~n9556;
  assign n9558 = ~n9220 & ~n9223;
  assign n9559 = ~n9423 & ~n9444;
  assign n9560 = n9558 & n9559;
  assign n9561 = ~n9558 & ~n9559;
  assign n9562 = ~n9560 & ~n9561;
  assign n9563 = ~n9195 & ~n9218;
  assign n9564 = pi5  & pi61 ;
  assign n9565 = pi4  & pi62 ;
  assign n9566 = ~n9564 & ~n9565;
  assign n9567 = pi61  & pi62 ;
  assign n9568 = n226 & n9567;
  assign n9569 = pi3  & pi63 ;
  assign n9570 = ~n9566 & n9569;
  assign n9571 = ~n9568 & n9570;
  assign n9572 = ~n9568 & ~n9571;
  assign n9573 = ~n9566 & n9572;
  assign n9574 = n9569 & ~n9571;
  assign n9575 = ~n9573 & ~n9574;
  assign n9576 = pi27  & pi39 ;
  assign n9577 = n2915 & n5055;
  assign n9578 = pi28  & pi38 ;
  assign n9579 = pi29  & pi37 ;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = n9576 & ~n9577;
  assign n9582 = ~n9580 & n9581;
  assign n9583 = n9576 & ~n9582;
  assign n9584 = ~n9577 & ~n9582;
  assign n9585 = ~n9580 & n9584;
  assign n9586 = ~n9583 & ~n9585;
  assign n9587 = ~n9575 & ~n9586;
  assign n9588 = ~n9575 & ~n9587;
  assign n9589 = ~n9586 & ~n9587;
  assign n9590 = ~n9588 & ~n9589;
  assign n9591 = pi11  & pi55 ;
  assign n9592 = pi19  & pi47 ;
  assign n9593 = pi12  & pi54 ;
  assign n9594 = n9592 & n9593;
  assign n9595 = ~n9592 & ~n9593;
  assign n9596 = n9591 & ~n9594;
  assign n9597 = ~n9595 & n9596;
  assign n9598 = n9591 & ~n9597;
  assign n9599 = ~n9594 & ~n9597;
  assign n9600 = ~n9595 & n9599;
  assign n9601 = ~n9598 & ~n9600;
  assign n9602 = ~n9590 & ~n9601;
  assign n9603 = ~n9590 & ~n9602;
  assign n9604 = ~n9601 & ~n9602;
  assign n9605 = ~n9603 & ~n9604;
  assign n9606 = pi9  & pi57 ;
  assign n9607 = pi24  & pi42 ;
  assign n9608 = ~n9606 & ~n9607;
  assign n9609 = pi24  & pi57 ;
  assign n9610 = n5752 & n9609;
  assign n9611 = pi23  & pi43 ;
  assign n9612 = ~n9608 & n9611;
  assign n9613 = ~n9610 & n9612;
  assign n9614 = ~n9610 & ~n9613;
  assign n9615 = ~n9608 & n9614;
  assign n9616 = n9611 & ~n9613;
  assign n9617 = ~n9615 & ~n9616;
  assign n9618 = pi20  & pi46 ;
  assign n9619 = n1481 & n5318;
  assign n9620 = pi21  & pi45 ;
  assign n9621 = pi22  & pi44 ;
  assign n9622 = ~n9620 & ~n9621;
  assign n9623 = n9618 & ~n9619;
  assign n9624 = ~n9622 & n9623;
  assign n9625 = n9618 & ~n9624;
  assign n9626 = ~n9619 & ~n9624;
  assign n9627 = ~n9622 & n9626;
  assign n9628 = ~n9625 & ~n9627;
  assign n9629 = ~n9617 & ~n9628;
  assign n9630 = ~n9617 & ~n9629;
  assign n9631 = ~n9628 & ~n9629;
  assign n9632 = ~n9630 & ~n9631;
  assign n9633 = pi10  & pi56 ;
  assign n9634 = n2310 & n6012;
  assign n9635 = pi25  & pi41 ;
  assign n9636 = pi26  & pi40 ;
  assign n9637 = ~n9635 & ~n9636;
  assign n9638 = n9633 & ~n9634;
  assign n9639 = ~n9637 & n9638;
  assign n9640 = n9633 & ~n9639;
  assign n9641 = ~n9634 & ~n9639;
  assign n9642 = ~n9637 & n9641;
  assign n9643 = ~n9640 & ~n9642;
  assign n9644 = ~n9632 & ~n9643;
  assign n9645 = ~n9632 & ~n9644;
  assign n9646 = ~n9643 & ~n9644;
  assign n9647 = ~n9645 & ~n9646;
  assign n9648 = pi13  & pi53 ;
  assign n9649 = pi15  & pi51 ;
  assign n9650 = ~n9648 & ~n9649;
  assign n9651 = n777 & n6765;
  assign n9652 = pi18  & pi48 ;
  assign n9653 = ~n9650 & n9652;
  assign n9654 = ~n9651 & n9653;
  assign n9655 = ~n9651 & ~n9654;
  assign n9656 = ~n9650 & n9655;
  assign n9657 = n9652 & ~n9654;
  assign n9658 = ~n9656 & ~n9657;
  assign n9659 = pi14  & pi52 ;
  assign n9660 = n2680 & n4691;
  assign n9661 = pi30  & pi36 ;
  assign n9662 = pi31  & pi35 ;
  assign n9663 = ~n9661 & ~n9662;
  assign n9664 = n9659 & ~n9660;
  assign n9665 = ~n9663 & n9664;
  assign n9666 = n9659 & ~n9665;
  assign n9667 = ~n9660 & ~n9665;
  assign n9668 = ~n9663 & n9667;
  assign n9669 = ~n9666 & ~n9668;
  assign n9670 = ~n9658 & ~n9669;
  assign n9671 = ~n9658 & ~n9670;
  assign n9672 = ~n9669 & ~n9670;
  assign n9673 = ~n9671 & ~n9672;
  assign n9674 = n989 & n5889;
  assign n9675 = pi16  & pi50 ;
  assign n9676 = ~n6584 & ~n9675;
  assign n9677 = n3827 & ~n9674;
  assign n9678 = ~n9676 & n9677;
  assign n9679 = n3827 & ~n9678;
  assign n9680 = ~n9674 & ~n9678;
  assign n9681 = ~n9676 & n9680;
  assign n9682 = ~n9679 & ~n9681;
  assign n9683 = ~n9673 & ~n9682;
  assign n9684 = ~n9673 & ~n9683;
  assign n9685 = ~n9682 & ~n9683;
  assign n9686 = ~n9684 & ~n9685;
  assign n9687 = ~n9647 & n9686;
  assign n9688 = n9647 & ~n9686;
  assign n9689 = ~n9687 & ~n9688;
  assign n9690 = ~n9605 & ~n9689;
  assign n9691 = n9605 & n9689;
  assign n9692 = ~n9690 & ~n9691;
  assign n9693 = ~n9563 & n9692;
  assign n9694 = n9563 & ~n9692;
  assign n9695 = ~n9693 & ~n9694;
  assign n9696 = ~n9200 & ~n9203;
  assign n9697 = ~n9206 & ~n9209;
  assign n9698 = n9696 & n9697;
  assign n9699 = ~n9696 & ~n9697;
  assign n9700 = ~n9698 & ~n9699;
  assign n9701 = ~n9280 & ~n9283;
  assign n9702 = ~n9700 & n9701;
  assign n9703 = n9700 & ~n9701;
  assign n9704 = ~n9702 & ~n9703;
  assign n9705 = ~n9212 & ~n9214;
  assign n9706 = ~n9287 & ~n9291;
  assign n9707 = ~n9705 & n9706;
  assign n9708 = n9705 & ~n9706;
  assign n9709 = ~n9707 & ~n9708;
  assign n9710 = n9704 & ~n9709;
  assign n9711 = ~n9704 & n9709;
  assign n9712 = ~n9710 & ~n9711;
  assign n9713 = n9695 & n9712;
  assign n9714 = ~n9695 & ~n9712;
  assign n9715 = ~n9713 & ~n9714;
  assign n9716 = n9562 & n9715;
  assign n9717 = ~n9562 & ~n9715;
  assign n9718 = ~n9716 & ~n9717;
  assign n9719 = ~n9557 & n9718;
  assign n9720 = ~n9557 & ~n9719;
  assign n9721 = n9718 & ~n9719;
  assign n9722 = ~n9720 & ~n9721;
  assign n9723 = ~n9462 & ~n9722;
  assign n9724 = n9462 & n9722;
  assign n9725 = ~n9723 & ~n9724;
  assign n9726 = ~n9461 & n9725;
  assign n9727 = n9461 & ~n9725;
  assign po67  = ~n9726 & ~n9727;
  assign n9729 = ~n9554 & ~n9719;
  assign n9730 = ~n9561 & ~n9716;
  assign n9731 = ~n9515 & ~n9518;
  assign n9732 = ~n9705 & ~n9706;
  assign n9733 = ~n9710 & ~n9732;
  assign n9734 = ~n9629 & ~n9644;
  assign n9735 = ~n9469 & ~n9482;
  assign n9736 = n9734 & n9735;
  assign n9737 = ~n9734 & ~n9735;
  assign n9738 = ~n9736 & ~n9737;
  assign n9739 = ~n9587 & ~n9602;
  assign n9740 = ~n9738 & n9739;
  assign n9741 = n9738 & ~n9739;
  assign n9742 = ~n9740 & ~n9741;
  assign n9743 = n9479 & n9572;
  assign n9744 = ~n9479 & ~n9572;
  assign n9745 = ~n9743 & ~n9744;
  assign n9746 = n9584 & ~n9745;
  assign n9747 = ~n9584 & n9745;
  assign n9748 = ~n9746 & ~n9747;
  assign n9749 = n9614 & n9641;
  assign n9750 = ~n9614 & ~n9641;
  assign n9751 = ~n9749 & ~n9750;
  assign n9752 = n9626 & ~n9751;
  assign n9753 = ~n9626 & n9751;
  assign n9754 = ~n9752 & ~n9753;
  assign n9755 = pi6  & pi61 ;
  assign n9756 = ~n9680 & n9755;
  assign n9757 = n9680 & ~n9755;
  assign n9758 = ~n9756 & ~n9757;
  assign n9759 = n9667 & ~n9758;
  assign n9760 = ~n9667 & n9758;
  assign n9761 = ~n9759 & ~n9760;
  assign n9762 = n9754 & n9761;
  assign n9763 = ~n9754 & ~n9761;
  assign n9764 = ~n9762 & ~n9763;
  assign n9765 = n9748 & n9764;
  assign n9766 = ~n9748 & ~n9764;
  assign n9767 = ~n9765 & ~n9766;
  assign n9768 = n9742 & n9767;
  assign n9769 = ~n9742 & ~n9767;
  assign n9770 = ~n9768 & ~n9769;
  assign n9771 = ~n9733 & n9770;
  assign n9772 = n9733 & ~n9770;
  assign n9773 = ~n9771 & ~n9772;
  assign n9774 = n9731 & ~n9773;
  assign n9775 = ~n9731 & n9773;
  assign n9776 = ~n9774 & ~n9775;
  assign n9777 = n9599 & n9655;
  assign n9778 = ~n9599 & ~n9655;
  assign n9779 = ~n9777 & ~n9778;
  assign n9780 = pi10  & pi57 ;
  assign n9781 = pi20  & pi56 ;
  assign n9782 = n7502 & n9781;
  assign n9783 = pi11  & pi56 ;
  assign n9784 = pi20  & pi47 ;
  assign n9785 = ~n9783 & ~n9784;
  assign n9786 = n9780 & ~n9782;
  assign n9787 = ~n9785 & n9786;
  assign n9788 = n9780 & ~n9787;
  assign n9789 = ~n9782 & ~n9787;
  assign n9790 = ~n9785 & n9789;
  assign n9791 = ~n9788 & ~n9790;
  assign n9792 = n9779 & ~n9791;
  assign n9793 = n9779 & ~n9792;
  assign n9794 = ~n9791 & ~n9792;
  assign n9795 = ~n9793 & ~n9794;
  assign n9796 = ~n9670 & ~n9683;
  assign n9797 = n9795 & n9796;
  assign n9798 = ~n9795 & ~n9796;
  assign n9799 = ~n9797 & ~n9798;
  assign n9800 = ~n9699 & ~n9703;
  assign n9801 = ~n9799 & n9800;
  assign n9802 = n9799 & ~n9800;
  assign n9803 = ~n9801 & ~n9802;
  assign n9804 = ~n9647 & ~n9686;
  assign n9805 = ~n9690 & ~n9804;
  assign n9806 = ~n9488 & ~n9494;
  assign n9807 = n9805 & n9806;
  assign n9808 = ~n9805 & ~n9806;
  assign n9809 = ~n9807 & ~n9808;
  assign n9810 = n9803 & n9809;
  assign n9811 = ~n9803 & ~n9809;
  assign n9812 = ~n9810 & ~n9811;
  assign n9813 = n9776 & n9812;
  assign n9814 = ~n9776 & ~n9812;
  assign n9815 = ~n9813 & ~n9814;
  assign n9816 = ~n9730 & n9815;
  assign n9817 = n9730 & ~n9815;
  assign n9818 = ~n9816 & ~n9817;
  assign n9819 = ~n9546 & ~n9550;
  assign n9820 = ~n9693 & ~n9713;
  assign n9821 = n9819 & n9820;
  assign n9822 = ~n9819 & ~n9820;
  assign n9823 = ~n9821 & ~n9822;
  assign n9824 = ~n9541 & ~n9543;
  assign n9825 = pi17  & pi50 ;
  assign n9826 = pi14  & pi53 ;
  assign n9827 = ~n9825 & ~n9826;
  assign n9828 = n9825 & n9826;
  assign n9829 = pi19  & pi48 ;
  assign n9830 = ~n9827 & n9829;
  assign n9831 = ~n9828 & n9830;
  assign n9832 = ~n9828 & ~n9831;
  assign n9833 = ~n9827 & n9832;
  assign n9834 = n9829 & ~n9831;
  assign n9835 = ~n9833 & ~n9834;
  assign n9836 = pi25  & pi42 ;
  assign n9837 = pi21  & pi46 ;
  assign n9838 = pi26  & pi41 ;
  assign n9839 = n9837 & n9838;
  assign n9840 = ~n9837 & ~n9838;
  assign n9841 = n9836 & ~n9839;
  assign n9842 = ~n9840 & n9841;
  assign n9843 = n9836 & ~n9842;
  assign n9844 = ~n9839 & ~n9842;
  assign n9845 = ~n9840 & n9844;
  assign n9846 = ~n9843 & ~n9845;
  assign n9847 = ~n9835 & ~n9846;
  assign n9848 = ~n9835 & ~n9847;
  assign n9849 = ~n9846 & ~n9847;
  assign n9850 = ~n9848 & ~n9849;
  assign n9851 = pi4  & pi63 ;
  assign n9852 = n2191 & n5548;
  assign n9853 = pi27  & pi40 ;
  assign n9854 = pi28  & pi39 ;
  assign n9855 = ~n9853 & ~n9854;
  assign n9856 = n9851 & ~n9852;
  assign n9857 = ~n9855 & n9856;
  assign n9858 = n9851 & ~n9857;
  assign n9859 = ~n9852 & ~n9857;
  assign n9860 = ~n9855 & n9859;
  assign n9861 = ~n9858 & ~n9860;
  assign n9862 = ~n9850 & ~n9861;
  assign n9863 = ~n9850 & ~n9862;
  assign n9864 = ~n9861 & ~n9862;
  assign n9865 = ~n9863 & ~n9864;
  assign n9866 = pi5  & pi62 ;
  assign n9867 = ~pi34  & ~n9866;
  assign n9868 = pi62  & n3433;
  assign n9869 = pi18  & pi49 ;
  assign n9870 = ~n9867 & n9869;
  assign n9871 = ~n9868 & n9870;
  assign n9872 = ~n9868 & ~n9871;
  assign n9873 = ~n9867 & n9872;
  assign n9874 = n9869 & ~n9871;
  assign n9875 = ~n9873 & ~n9874;
  assign n9876 = pi31  & pi36 ;
  assign n9877 = n3106 & n6138;
  assign n9878 = pi32  & pi35 ;
  assign n9879 = ~n3900 & ~n9878;
  assign n9880 = n9876 & ~n9877;
  assign n9881 = ~n9879 & n9880;
  assign n9882 = n9876 & ~n9881;
  assign n9883 = ~n9877 & ~n9881;
  assign n9884 = ~n9879 & n9883;
  assign n9885 = ~n9882 & ~n9884;
  assign n9886 = ~n9875 & ~n9885;
  assign n9887 = ~n9875 & ~n9886;
  assign n9888 = ~n9885 & ~n9886;
  assign n9889 = ~n9887 & ~n9888;
  assign n9890 = pi29  & pi38 ;
  assign n9891 = pi54  & pi55 ;
  assign n9892 = n952 & n9891;
  assign n9893 = pi12  & pi55 ;
  assign n9894 = pi13  & pi54 ;
  assign n9895 = ~n9893 & ~n9894;
  assign n9896 = n9890 & ~n9892;
  assign n9897 = ~n9895 & n9896;
  assign n9898 = n9890 & ~n9897;
  assign n9899 = ~n9892 & ~n9897;
  assign n9900 = ~n9895 & n9899;
  assign n9901 = ~n9898 & ~n9900;
  assign n9902 = ~n9889 & ~n9901;
  assign n9903 = ~n9889 & ~n9902;
  assign n9904 = ~n9901 & ~n9902;
  assign n9905 = ~n9903 & ~n9904;
  assign n9906 = pi8  & pi59 ;
  assign n9907 = pi9  & pi58 ;
  assign n9908 = ~n9906 & ~n9907;
  assign n9909 = n414 & n9402;
  assign n9910 = pi7  & pi60 ;
  assign n9911 = ~n9908 & n9910;
  assign n9912 = ~n9909 & n9911;
  assign n9913 = ~n9909 & ~n9912;
  assign n9914 = ~n9908 & n9913;
  assign n9915 = n9910 & ~n9912;
  assign n9916 = ~n9914 & ~n9915;
  assign n9917 = pi22  & pi45 ;
  assign n9918 = n2110 & n6836;
  assign n9919 = pi23  & pi44 ;
  assign n9920 = pi24  & pi43 ;
  assign n9921 = ~n9919 & ~n9920;
  assign n9922 = n9917 & ~n9918;
  assign n9923 = ~n9921 & n9922;
  assign n9924 = n9917 & ~n9923;
  assign n9925 = ~n9918 & ~n9923;
  assign n9926 = ~n9921 & n9925;
  assign n9927 = ~n9924 & ~n9926;
  assign n9928 = ~n9916 & ~n9927;
  assign n9929 = ~n9916 & ~n9928;
  assign n9930 = ~n9927 & ~n9928;
  assign n9931 = ~n9929 & ~n9930;
  assign n9932 = pi15  & pi52 ;
  assign n9933 = pi16  & pi51 ;
  assign n9934 = pi30  & pi37 ;
  assign n9935 = n9933 & n9934;
  assign n9936 = ~n9933 & ~n9934;
  assign n9937 = n9932 & ~n9935;
  assign n9938 = ~n9936 & n9937;
  assign n9939 = n9932 & ~n9938;
  assign n9940 = ~n9935 & ~n9938;
  assign n9941 = ~n9936 & n9940;
  assign n9942 = ~n9939 & ~n9941;
  assign n9943 = ~n9931 & ~n9942;
  assign n9944 = ~n9931 & ~n9943;
  assign n9945 = ~n9942 & ~n9943;
  assign n9946 = ~n9944 & ~n9945;
  assign n9947 = ~n9905 & n9946;
  assign n9948 = n9905 & ~n9946;
  assign n9949 = ~n9947 & ~n9948;
  assign n9950 = ~n9865 & ~n9949;
  assign n9951 = n9865 & n9949;
  assign n9952 = ~n9950 & ~n9951;
  assign n9953 = ~n9824 & n9952;
  assign n9954 = n9824 & ~n9952;
  assign n9955 = ~n9953 & ~n9954;
  assign n9956 = ~n9503 & ~n9506;
  assign n9957 = ~n9523 & ~n9526;
  assign n9958 = n9956 & n9957;
  assign n9959 = ~n9956 & ~n9957;
  assign n9960 = ~n9958 & ~n9959;
  assign n9961 = ~n9497 & ~n9500;
  assign n9962 = ~n9960 & n9961;
  assign n9963 = n9960 & ~n9961;
  assign n9964 = ~n9962 & ~n9963;
  assign n9965 = ~n9510 & ~n9512;
  assign n9966 = ~n9531 & ~n9535;
  assign n9967 = n9965 & n9966;
  assign n9968 = ~n9965 & ~n9966;
  assign n9969 = ~n9967 & ~n9968;
  assign n9970 = n9964 & n9969;
  assign n9971 = ~n9964 & ~n9969;
  assign n9972 = ~n9970 & ~n9971;
  assign n9973 = n9955 & n9972;
  assign n9974 = ~n9955 & ~n9972;
  assign n9975 = ~n9973 & ~n9974;
  assign n9976 = n9823 & n9975;
  assign n9977 = ~n9823 & ~n9975;
  assign n9978 = ~n9976 & ~n9977;
  assign n9979 = n9818 & n9978;
  assign n9980 = n9818 & ~n9979;
  assign n9981 = n9978 & ~n9979;
  assign n9982 = ~n9980 & ~n9981;
  assign n9983 = ~n9729 & ~n9982;
  assign n9984 = n9729 & n9982;
  assign n9985 = ~n9983 & ~n9984;
  assign n9986 = ~n9723 & ~n9726;
  assign n9987 = ~n9985 & n9986;
  assign n9988 = n9985 & ~n9986;
  assign po68  = ~n9987 & ~n9988;
  assign n9990 = ~n9822 & ~n9976;
  assign n9991 = ~n9968 & ~n9970;
  assign n9992 = n9832 & n9844;
  assign n9993 = ~n9832 & ~n9844;
  assign n9994 = ~n9992 & ~n9993;
  assign n9995 = n9899 & ~n9994;
  assign n9996 = ~n9899 & n9994;
  assign n9997 = ~n9995 & ~n9996;
  assign n9998 = ~n9847 & ~n9862;
  assign n9999 = ~n9886 & ~n9902;
  assign n10000 = n9998 & n9999;
  assign n10001 = ~n9998 & ~n9999;
  assign n10002 = ~n10000 & ~n10001;
  assign n10003 = n9997 & n10002;
  assign n10004 = ~n9997 & ~n10002;
  assign n10005 = ~n10003 & ~n10004;
  assign n10006 = ~n9959 & ~n9963;
  assign n10007 = n9789 & n9925;
  assign n10008 = ~n9789 & ~n9925;
  assign n10009 = ~n10007 & ~n10008;
  assign n10010 = n9913 & ~n10009;
  assign n10011 = ~n9913 & n10009;
  assign n10012 = ~n10010 & ~n10011;
  assign n10013 = n9859 & n9883;
  assign n10014 = ~n9859 & ~n9883;
  assign n10015 = ~n10013 & ~n10014;
  assign n10016 = n9940 & ~n10015;
  assign n10017 = ~n9940 & n10015;
  assign n10018 = ~n10016 & ~n10017;
  assign n10019 = n10012 & n10018;
  assign n10020 = ~n10012 & ~n10018;
  assign n10021 = ~n10019 & ~n10020;
  assign n10022 = ~n10006 & n10021;
  assign n10023 = n10006 & ~n10021;
  assign n10024 = ~n10022 & ~n10023;
  assign n10025 = n10005 & n10024;
  assign n10026 = ~n10005 & ~n10024;
  assign n10027 = ~n10025 & ~n10026;
  assign n10028 = ~n9991 & n10027;
  assign n10029 = n9991 & ~n10027;
  assign n10030 = ~n10028 & ~n10029;
  assign n10031 = ~n9768 & ~n9771;
  assign n10032 = ~n9905 & ~n9946;
  assign n10033 = ~n9950 & ~n10032;
  assign n10034 = ~n9778 & ~n9792;
  assign n10035 = ~n9750 & ~n9753;
  assign n10036 = n10034 & n10035;
  assign n10037 = ~n10034 & ~n10035;
  assign n10038 = ~n10036 & ~n10037;
  assign n10039 = ~n9928 & ~n9943;
  assign n10040 = ~n10038 & n10039;
  assign n10041 = n10038 & ~n10039;
  assign n10042 = ~n10040 & ~n10041;
  assign n10043 = n521 & n9054;
  assign n10044 = pi8  & pi60 ;
  assign n10045 = ~n10043 & n10044;
  assign n10046 = pi7  & pi61 ;
  assign n10047 = ~n10043 & n10046;
  assign n10048 = ~n10045 & ~n10047;
  assign n10049 = ~n9872 & ~n10048;
  assign n10050 = ~n9872 & ~n10049;
  assign n10051 = ~n10048 & ~n10049;
  assign n10052 = ~n10050 & ~n10051;
  assign n10053 = ~n9756 & ~n9760;
  assign n10054 = n10052 & n10053;
  assign n10055 = ~n10052 & ~n10053;
  assign n10056 = ~n10054 & ~n10055;
  assign n10057 = ~n9744 & ~n9747;
  assign n10058 = ~n10056 & n10057;
  assign n10059 = n10056 & ~n10057;
  assign n10060 = ~n10058 & ~n10059;
  assign n10061 = n10042 & n10060;
  assign n10062 = ~n10042 & ~n10060;
  assign n10063 = ~n10061 & ~n10062;
  assign n10064 = ~n10033 & n10063;
  assign n10065 = n10033 & ~n10063;
  assign n10066 = ~n10064 & ~n10065;
  assign n10067 = ~n10031 & n10066;
  assign n10068 = ~n10031 & ~n10067;
  assign n10069 = n10066 & ~n10067;
  assign n10070 = ~n10068 & ~n10069;
  assign n10071 = n10030 & ~n10070;
  assign n10072 = n10030 & ~n10071;
  assign n10073 = ~n10070 & ~n10071;
  assign n10074 = ~n10072 & ~n10073;
  assign n10075 = ~n9990 & ~n10074;
  assign n10076 = ~n9990 & ~n10075;
  assign n10077 = ~n10074 & ~n10075;
  assign n10078 = ~n10076 & ~n10077;
  assign n10079 = ~n9775 & ~n9813;
  assign n10080 = ~n9953 & ~n9973;
  assign n10081 = ~n9808 & ~n9810;
  assign n10082 = ~n9762 & ~n9765;
  assign n10083 = ~n9737 & ~n9741;
  assign n10084 = n10082 & n10083;
  assign n10085 = ~n10082 & ~n10083;
  assign n10086 = ~n10084 & ~n10085;
  assign n10087 = ~n9798 & ~n9802;
  assign n10088 = ~n10086 & n10087;
  assign n10089 = n10086 & ~n10087;
  assign n10090 = ~n10088 & ~n10089;
  assign n10091 = pi10  & pi58 ;
  assign n10092 = pi11  & pi57 ;
  assign n10093 = ~n10091 & ~n10092;
  assign n10094 = n1111 & n8144;
  assign n10095 = pi9  & pi59 ;
  assign n10096 = ~n10093 & n10095;
  assign n10097 = ~n10094 & n10096;
  assign n10098 = ~n10094 & ~n10097;
  assign n10099 = ~n10093 & n10098;
  assign n10100 = n10095 & ~n10097;
  assign n10101 = ~n10099 & ~n10100;
  assign n10102 = pi27  & pi41 ;
  assign n10103 = n2915 & n5548;
  assign n10104 = pi28  & pi40 ;
  assign n10105 = pi29  & pi39 ;
  assign n10106 = ~n10104 & ~n10105;
  assign n10107 = n10102 & ~n10103;
  assign n10108 = ~n10106 & n10107;
  assign n10109 = n10102 & ~n10108;
  assign n10110 = ~n10103 & ~n10108;
  assign n10111 = ~n10106 & n10110;
  assign n10112 = ~n10109 & ~n10111;
  assign n10113 = ~n10101 & ~n10112;
  assign n10114 = ~n10101 & ~n10113;
  assign n10115 = ~n10112 & ~n10113;
  assign n10116 = ~n10114 & ~n10115;
  assign n10117 = pi21  & pi47 ;
  assign n10118 = n326 & n9123;
  assign n10119 = pi5  & pi63 ;
  assign n10120 = pi6  & pi62 ;
  assign n10121 = ~n10119 & ~n10120;
  assign n10122 = n10117 & ~n10118;
  assign n10123 = ~n10121 & n10122;
  assign n10124 = n10117 & ~n10123;
  assign n10125 = ~n10118 & ~n10123;
  assign n10126 = ~n10121 & n10125;
  assign n10127 = ~n10124 & ~n10126;
  assign n10128 = ~n10116 & ~n10127;
  assign n10129 = ~n10116 & ~n10128;
  assign n10130 = ~n10127 & ~n10128;
  assign n10131 = ~n10129 & ~n10130;
  assign n10132 = pi18  & pi50 ;
  assign n10133 = pi19  & pi49 ;
  assign n10134 = ~n10132 & ~n10133;
  assign n10135 = n1085 & n5889;
  assign n10136 = n2811 & ~n10134;
  assign n10137 = ~n10135 & n10136;
  assign n10138 = ~n10135 & ~n10137;
  assign n10139 = ~n10134 & n10138;
  assign n10140 = n2811 & ~n10137;
  assign n10141 = ~n10139 & ~n10140;
  assign n10142 = pi30  & pi38 ;
  assign n10143 = n3567 & n4500;
  assign n10144 = pi31  & pi37 ;
  assign n10145 = pi32  & pi36 ;
  assign n10146 = ~n10144 & ~n10145;
  assign n10147 = n10142 & ~n10143;
  assign n10148 = ~n10146 & n10147;
  assign n10149 = n10142 & ~n10148;
  assign n10150 = ~n10143 & ~n10148;
  assign n10151 = ~n10146 & n10150;
  assign n10152 = ~n10149 & ~n10151;
  assign n10153 = ~n10141 & ~n10152;
  assign n10154 = ~n10141 & ~n10153;
  assign n10155 = ~n10152 & ~n10153;
  assign n10156 = ~n10154 & ~n10155;
  assign n10157 = pi12  & pi56 ;
  assign n10158 = pi13  & pi55 ;
  assign n10159 = n7238 & n10158;
  assign n10160 = ~n7238 & ~n10158;
  assign n10161 = n10157 & ~n10159;
  assign n10162 = ~n10160 & n10161;
  assign n10163 = n10157 & ~n10162;
  assign n10164 = ~n10159 & ~n10162;
  assign n10165 = ~n10160 & n10164;
  assign n10166 = ~n10163 & ~n10165;
  assign n10167 = ~n10156 & ~n10166;
  assign n10168 = ~n10156 & ~n10167;
  assign n10169 = ~n10166 & ~n10167;
  assign n10170 = ~n10168 & ~n10169;
  assign n10171 = pi15  & pi53 ;
  assign n10172 = pi16  & pi52 ;
  assign n10173 = ~n10171 & ~n10172;
  assign n10174 = n840 & n9144;
  assign n10175 = pi14  & pi54 ;
  assign n10176 = ~n10173 & n10175;
  assign n10177 = ~n10174 & n10176;
  assign n10178 = ~n10174 & ~n10177;
  assign n10179 = ~n10173 & n10178;
  assign n10180 = n10175 & ~n10177;
  assign n10181 = ~n10179 & ~n10180;
  assign n10182 = pi20  & pi48 ;
  assign n10183 = pi23  & pi45 ;
  assign n10184 = pi22  & pi46 ;
  assign n10185 = ~n10183 & ~n10184;
  assign n10186 = n1806 & n7513;
  assign n10187 = n10182 & ~n10185;
  assign n10188 = ~n10186 & n10187;
  assign n10189 = n10182 & ~n10188;
  assign n10190 = ~n10186 & ~n10188;
  assign n10191 = ~n10185 & n10190;
  assign n10192 = ~n10189 & ~n10191;
  assign n10193 = ~n10181 & ~n10192;
  assign n10194 = ~n10181 & ~n10193;
  assign n10195 = ~n10192 & ~n10193;
  assign n10196 = ~n10194 & ~n10195;
  assign n10197 = pi24  & pi44 ;
  assign n10198 = n2310 & n6458;
  assign n10199 = pi25  & pi43 ;
  assign n10200 = pi26  & pi42 ;
  assign n10201 = ~n10199 & ~n10200;
  assign n10202 = n10197 & ~n10198;
  assign n10203 = ~n10201 & n10202;
  assign n10204 = n10197 & ~n10203;
  assign n10205 = ~n10198 & ~n10203;
  assign n10206 = ~n10201 & n10205;
  assign n10207 = ~n10204 & ~n10206;
  assign n10208 = ~n10196 & ~n10207;
  assign n10209 = ~n10196 & ~n10208;
  assign n10210 = ~n10207 & ~n10208;
  assign n10211 = ~n10209 & ~n10210;
  assign n10212 = ~n10170 & n10211;
  assign n10213 = n10170 & ~n10211;
  assign n10214 = ~n10212 & ~n10213;
  assign n10215 = ~n10131 & ~n10214;
  assign n10216 = n10131 & n10214;
  assign n10217 = ~n10215 & ~n10216;
  assign n10218 = n10090 & n10217;
  assign n10219 = ~n10090 & ~n10217;
  assign n10220 = ~n10218 & ~n10219;
  assign n10221 = ~n10081 & n10220;
  assign n10222 = n10081 & ~n10220;
  assign n10223 = ~n10221 & ~n10222;
  assign n10224 = ~n10080 & n10223;
  assign n10225 = n10080 & ~n10223;
  assign n10226 = ~n10224 & ~n10225;
  assign n10227 = ~n10079 & n10226;
  assign n10228 = n10079 & ~n10226;
  assign n10229 = ~n10227 & ~n10228;
  assign n10230 = ~n10078 & ~n10229;
  assign n10231 = n10078 & n10229;
  assign n10232 = ~n10230 & ~n10231;
  assign n10233 = ~n9816 & ~n9979;
  assign n10234 = n10232 & n10233;
  assign n10235 = ~n10232 & ~n10233;
  assign n10236 = ~n10234 & ~n10235;
  assign n10237 = ~n9983 & ~n9988;
  assign n10238 = ~n10236 & n10237;
  assign n10239 = n10236 & ~n10237;
  assign po69  = ~n10238 & ~n10239;
  assign n10241 = ~n10224 & ~n10227;
  assign n10242 = ~n10025 & ~n10028;
  assign n10243 = ~n10170 & ~n10211;
  assign n10244 = ~n10215 & ~n10243;
  assign n10245 = ~n10019 & ~n10022;
  assign n10246 = n10164 & n10205;
  assign n10247 = ~n10164 & ~n10205;
  assign n10248 = ~n10246 & ~n10247;
  assign n10249 = n10110 & ~n10248;
  assign n10250 = ~n10110 & n10248;
  assign n10251 = ~n10249 & ~n10250;
  assign n10252 = ~n10014 & ~n10017;
  assign n10253 = ~n9993 & ~n9996;
  assign n10254 = n10252 & n10253;
  assign n10255 = ~n10252 & ~n10253;
  assign n10256 = ~n10254 & ~n10255;
  assign n10257 = n10251 & n10256;
  assign n10258 = ~n10251 & ~n10256;
  assign n10259 = ~n10257 & ~n10258;
  assign n10260 = ~n10245 & n10259;
  assign n10261 = n10245 & ~n10259;
  assign n10262 = ~n10260 & ~n10261;
  assign n10263 = ~n10244 & n10262;
  assign n10264 = n10244 & ~n10262;
  assign n10265 = ~n10263 & ~n10264;
  assign n10266 = n10242 & ~n10265;
  assign n10267 = ~n10242 & n10265;
  assign n10268 = ~n10266 & ~n10267;
  assign n10269 = ~n10085 & ~n10089;
  assign n10270 = ~n10153 & ~n10167;
  assign n10271 = ~n10193 & ~n10208;
  assign n10272 = n10270 & n10271;
  assign n10273 = ~n10270 & ~n10271;
  assign n10274 = ~n10272 & ~n10273;
  assign n10275 = ~n10055 & ~n10059;
  assign n10276 = ~n10274 & n10275;
  assign n10277 = n10274 & ~n10275;
  assign n10278 = ~n10276 & ~n10277;
  assign n10279 = n10098 & n10125;
  assign n10280 = ~n10098 & ~n10125;
  assign n10281 = ~n10279 & ~n10280;
  assign n10282 = n10190 & ~n10281;
  assign n10283 = ~n10190 & n10281;
  assign n10284 = ~n10282 & ~n10283;
  assign n10285 = n10138 & n10150;
  assign n10286 = ~n10138 & ~n10150;
  assign n10287 = ~n10285 & ~n10286;
  assign n10288 = n10178 & ~n10287;
  assign n10289 = ~n10178 & n10287;
  assign n10290 = ~n10288 & ~n10289;
  assign n10291 = ~n10113 & ~n10128;
  assign n10292 = ~n10290 & n10291;
  assign n10293 = n10290 & ~n10291;
  assign n10294 = ~n10292 & ~n10293;
  assign n10295 = n10284 & n10294;
  assign n10296 = ~n10284 & ~n10294;
  assign n10297 = ~n10295 & ~n10296;
  assign n10298 = n10278 & n10297;
  assign n10299 = ~n10278 & ~n10297;
  assign n10300 = ~n10298 & ~n10299;
  assign n10301 = n10269 & ~n10300;
  assign n10302 = ~n10269 & n10300;
  assign n10303 = ~n10301 & ~n10302;
  assign n10304 = n10268 & n10303;
  assign n10305 = ~n10268 & ~n10303;
  assign n10306 = ~n10304 & ~n10305;
  assign n10307 = ~n10241 & n10306;
  assign n10308 = n10241 & ~n10306;
  assign n10309 = ~n10307 & ~n10308;
  assign n10310 = ~n10067 & ~n10071;
  assign n10311 = ~n10218 & ~n10221;
  assign n10312 = n10310 & n10311;
  assign n10313 = ~n10310 & ~n10311;
  assign n10314 = ~n10312 & ~n10313;
  assign n10315 = ~n10001 & ~n10003;
  assign n10316 = pi17  & pi52 ;
  assign n10317 = pi18  & pi51 ;
  assign n10318 = ~n10316 & ~n10317;
  assign n10319 = pi51  & pi52 ;
  assign n10320 = n1199 & n10319;
  assign n10321 = pi19  & pi50 ;
  assign n10322 = ~n10318 & n10321;
  assign n10323 = ~n10320 & n10322;
  assign n10324 = ~n10320 & ~n10323;
  assign n10325 = ~n10318 & n10324;
  assign n10326 = n10321 & ~n10323;
  assign n10327 = ~n10325 & ~n10326;
  assign n10328 = pi28  & pi41 ;
  assign n10329 = n4908 & n5548;
  assign n10330 = pi29  & pi40 ;
  assign n10331 = pi30  & pi39 ;
  assign n10332 = ~n10330 & ~n10331;
  assign n10333 = n10328 & ~n10329;
  assign n10334 = ~n10332 & n10333;
  assign n10335 = n10328 & ~n10334;
  assign n10336 = ~n10329 & ~n10334;
  assign n10337 = ~n10332 & n10336;
  assign n10338 = ~n10335 & ~n10337;
  assign n10339 = ~n10327 & ~n10338;
  assign n10340 = ~n10327 & ~n10339;
  assign n10341 = ~n10338 & ~n10339;
  assign n10342 = ~n10340 & ~n10341;
  assign n10343 = ~n10008 & ~n10011;
  assign n10344 = n10342 & n10343;
  assign n10345 = ~n10342 & ~n10343;
  assign n10346 = ~n10344 & ~n10345;
  assign n10347 = pi62  & n3887;
  assign n10348 = n3106 & ~n10347;
  assign n10349 = ~n10347 & ~n10348;
  assign n10350 = pi7  & pi62 ;
  assign n10351 = ~pi35  & ~n10350;
  assign n10352 = n10349 & ~n10351;
  assign n10353 = n3106 & ~n10348;
  assign n10354 = ~n10352 & ~n10353;
  assign n10355 = pi31  & pi38 ;
  assign n10356 = n4500 & n6138;
  assign n10357 = pi33  & pi36 ;
  assign n10358 = pi32  & pi37 ;
  assign n10359 = ~n10357 & ~n10358;
  assign n10360 = n10355 & ~n10356;
  assign n10361 = ~n10359 & n10360;
  assign n10362 = n10355 & ~n10361;
  assign n10363 = ~n10356 & ~n10361;
  assign n10364 = ~n10359 & n10363;
  assign n10365 = ~n10362 & ~n10364;
  assign n10366 = ~n10354 & ~n10365;
  assign n10367 = ~n10354 & ~n10366;
  assign n10368 = ~n10365 & ~n10366;
  assign n10369 = ~n10367 & ~n10368;
  assign n10370 = pi15  & pi54 ;
  assign n10371 = pi20  & pi49 ;
  assign n10372 = pi16  & pi53 ;
  assign n10373 = n10371 & n10372;
  assign n10374 = ~n10371 & ~n10372;
  assign n10375 = n10370 & ~n10373;
  assign n10376 = ~n10374 & n10375;
  assign n10377 = n10370 & ~n10376;
  assign n10378 = ~n10373 & ~n10376;
  assign n10379 = ~n10374 & n10378;
  assign n10380 = ~n10377 & ~n10379;
  assign n10381 = ~n10369 & ~n10380;
  assign n10382 = ~n10369 & ~n10381;
  assign n10383 = ~n10380 & ~n10381;
  assign n10384 = ~n10382 & ~n10383;
  assign n10385 = n10346 & ~n10384;
  assign n10386 = ~n10346 & n10384;
  assign n10387 = ~n10385 & ~n10386;
  assign n10388 = ~n10315 & n10387;
  assign n10389 = ~n10315 & ~n10388;
  assign n10390 = ~n10385 & ~n10388;
  assign n10391 = ~n10386 & n10390;
  assign n10392 = ~n10389 & ~n10391;
  assign n10393 = ~n10061 & ~n10064;
  assign n10394 = ~n10392 & ~n10393;
  assign n10395 = ~n10392 & ~n10394;
  assign n10396 = ~n10393 & ~n10394;
  assign n10397 = ~n10395 & ~n10396;
  assign n10398 = pi9  & pi60 ;
  assign n10399 = pi10  & pi59 ;
  assign n10400 = ~n10398 & ~n10399;
  assign n10401 = n591 & n8854;
  assign n10402 = pi8  & pi61 ;
  assign n10403 = ~n10400 & n10402;
  assign n10404 = ~n10401 & n10403;
  assign n10405 = ~n10401 & ~n10404;
  assign n10406 = ~n10400 & n10405;
  assign n10407 = n10402 & ~n10404;
  assign n10408 = ~n10406 & ~n10407;
  assign n10409 = pi23  & pi46 ;
  assign n10410 = n1789 & n5318;
  assign n10411 = pi24  & pi45 ;
  assign n10412 = pi25  & pi44 ;
  assign n10413 = ~n10411 & ~n10412;
  assign n10414 = n10409 & ~n10410;
  assign n10415 = ~n10413 & n10414;
  assign n10416 = n10409 & ~n10415;
  assign n10417 = ~n10410 & ~n10415;
  assign n10418 = ~n10413 & n10417;
  assign n10419 = ~n10416 & ~n10418;
  assign n10420 = ~n10408 & ~n10419;
  assign n10421 = ~n10408 & ~n10420;
  assign n10422 = ~n10419 & ~n10420;
  assign n10423 = ~n10421 & ~n10422;
  assign n10424 = pi6  & pi63 ;
  assign n10425 = n2646 & n6458;
  assign n10426 = pi26  & pi43 ;
  assign n10427 = pi27  & pi42 ;
  assign n10428 = ~n10426 & ~n10427;
  assign n10429 = n10424 & ~n10425;
  assign n10430 = ~n10428 & n10429;
  assign n10431 = n10424 & ~n10430;
  assign n10432 = ~n10425 & ~n10430;
  assign n10433 = ~n10428 & n10432;
  assign n10434 = ~n10431 & ~n10433;
  assign n10435 = ~n10423 & ~n10434;
  assign n10436 = ~n10423 & ~n10435;
  assign n10437 = ~n10434 & ~n10435;
  assign n10438 = ~n10436 & ~n10437;
  assign n10439 = ~n10037 & ~n10041;
  assign n10440 = n10438 & n10439;
  assign n10441 = ~n10438 & ~n10439;
  assign n10442 = ~n10440 & ~n10441;
  assign n10443 = pi11  & pi58 ;
  assign n10444 = n952 & n7643;
  assign n10445 = pi12  & pi57 ;
  assign n10446 = pi13  & pi56 ;
  assign n10447 = ~n10445 & ~n10446;
  assign n10448 = n10443 & ~n10444;
  assign n10449 = ~n10447 & n10448;
  assign n10450 = n10443 & ~n10449;
  assign n10451 = ~n10444 & ~n10449;
  assign n10452 = ~n10447 & n10451;
  assign n10453 = ~n10450 & ~n10452;
  assign n10454 = ~n10043 & ~n10049;
  assign n10455 = ~n10453 & n10454;
  assign n10456 = n10453 & ~n10454;
  assign n10457 = ~n10455 & ~n10456;
  assign n10458 = pi14  & pi55 ;
  assign n10459 = n1481 & n5823;
  assign n10460 = pi21  & pi48 ;
  assign n10461 = pi22  & pi47 ;
  assign n10462 = ~n10460 & ~n10461;
  assign n10463 = n10458 & ~n10459;
  assign n10464 = ~n10462 & n10463;
  assign n10465 = n10458 & ~n10464;
  assign n10466 = ~n10459 & ~n10464;
  assign n10467 = ~n10462 & n10466;
  assign n10468 = ~n10465 & ~n10467;
  assign n10469 = ~n10457 & ~n10468;
  assign n10470 = n10457 & n10468;
  assign n10471 = ~n10469 & ~n10470;
  assign n10472 = n10442 & n10471;
  assign n10473 = ~n10442 & ~n10471;
  assign n10474 = ~n10472 & ~n10473;
  assign n10475 = ~n10397 & n10474;
  assign n10476 = ~n10397 & ~n10475;
  assign n10477 = n10474 & ~n10475;
  assign n10478 = ~n10476 & ~n10477;
  assign n10479 = n10314 & ~n10478;
  assign n10480 = ~n10314 & n10478;
  assign n10481 = ~n10479 & ~n10480;
  assign n10482 = n10309 & n10481;
  assign n10483 = n10309 & ~n10482;
  assign n10484 = n10481 & ~n10482;
  assign n10485 = ~n10483 & ~n10484;
  assign n10486 = ~n10078 & n10229;
  assign n10487 = ~n10075 & ~n10486;
  assign n10488 = ~n10485 & ~n10487;
  assign n10489 = n10485 & n10487;
  assign n10490 = ~n10488 & ~n10489;
  assign n10491 = ~n10235 & ~n10239;
  assign n10492 = ~n10490 & n10491;
  assign n10493 = n10490 & ~n10491;
  assign po70  = ~n10492 & ~n10493;
  assign n10495 = ~n10307 & ~n10482;
  assign n10496 = ~n10267 & ~n10304;
  assign n10497 = n10336 & n10432;
  assign n10498 = ~n10336 & ~n10432;
  assign n10499 = ~n10497 & ~n10498;
  assign n10500 = n10417 & ~n10499;
  assign n10501 = ~n10417 & n10499;
  assign n10502 = ~n10500 & ~n10501;
  assign n10503 = pi8  & pi62 ;
  assign n10504 = ~n10349 & n10503;
  assign n10505 = n10349 & ~n10503;
  assign n10506 = ~n10363 & ~n10504;
  assign n10507 = ~n10505 & n10506;
  assign n10508 = ~n10363 & ~n10507;
  assign n10509 = ~n10504 & ~n10507;
  assign n10510 = ~n10505 & n10509;
  assign n10511 = ~n10508 & ~n10510;
  assign n10512 = n10502 & ~n10511;
  assign n10513 = n10502 & ~n10512;
  assign n10514 = ~n10511 & ~n10512;
  assign n10515 = ~n10513 & ~n10514;
  assign n10516 = ~n10339 & ~n10345;
  assign n10517 = n10515 & n10516;
  assign n10518 = ~n10515 & ~n10516;
  assign n10519 = ~n10517 & ~n10518;
  assign n10520 = ~n10420 & ~n10435;
  assign n10521 = ~n10453 & ~n10454;
  assign n10522 = ~n10469 & ~n10521;
  assign n10523 = n10520 & n10522;
  assign n10524 = ~n10520 & ~n10522;
  assign n10525 = ~n10523 & ~n10524;
  assign n10526 = ~n10366 & ~n10381;
  assign n10527 = ~n10525 & n10526;
  assign n10528 = n10525 & ~n10526;
  assign n10529 = ~n10527 & ~n10528;
  assign n10530 = ~n10390 & n10529;
  assign n10531 = n10390 & ~n10529;
  assign n10532 = ~n10530 & ~n10531;
  assign n10533 = ~n10519 & ~n10532;
  assign n10534 = n10519 & n10532;
  assign n10535 = ~n10533 & ~n10534;
  assign n10536 = ~n10496 & n10535;
  assign n10537 = ~n10496 & ~n10536;
  assign n10538 = n10535 & ~n10536;
  assign n10539 = ~n10537 & ~n10538;
  assign n10540 = ~n10293 & ~n10295;
  assign n10541 = pi7  & pi63 ;
  assign n10542 = pi23  & pi47 ;
  assign n10543 = ~n10541 & ~n10542;
  assign n10544 = n10541 & n10542;
  assign n10545 = pi28  & pi42 ;
  assign n10546 = ~n10543 & n10545;
  assign n10547 = ~n10544 & n10546;
  assign n10548 = ~n10544 & ~n10547;
  assign n10549 = ~n10543 & n10548;
  assign n10550 = n10545 & ~n10547;
  assign n10551 = ~n10549 & ~n10550;
  assign n10552 = pi29  & pi41 ;
  assign n10553 = n2680 & n5548;
  assign n10554 = pi30  & pi40 ;
  assign n10555 = pi31  & pi39 ;
  assign n10556 = ~n10554 & ~n10555;
  assign n10557 = n10552 & ~n10553;
  assign n10558 = ~n10556 & n10557;
  assign n10559 = n10552 & ~n10558;
  assign n10560 = ~n10553 & ~n10558;
  assign n10561 = ~n10556 & n10560;
  assign n10562 = ~n10559 & ~n10561;
  assign n10563 = ~n10551 & ~n10562;
  assign n10564 = ~n10551 & ~n10563;
  assign n10565 = ~n10562 & ~n10563;
  assign n10566 = ~n10564 & ~n10565;
  assign n10567 = ~n10286 & ~n10289;
  assign n10568 = n10566 & n10567;
  assign n10569 = ~n10566 & ~n10567;
  assign n10570 = ~n10568 & ~n10569;
  assign n10571 = pi14  & pi56 ;
  assign n10572 = pi15  & pi55 ;
  assign n10573 = ~n10571 & ~n10572;
  assign n10574 = n1041 & n8521;
  assign n10575 = pi22  & pi48 ;
  assign n10576 = ~n10573 & n10575;
  assign n10577 = ~n10574 & n10576;
  assign n10578 = ~n10574 & ~n10577;
  assign n10579 = ~n10573 & n10578;
  assign n10580 = n10575 & ~n10577;
  assign n10581 = ~n10579 & ~n10580;
  assign n10582 = pi25  & pi45 ;
  assign n10583 = n2646 & n6836;
  assign n10584 = pi26  & pi44 ;
  assign n10585 = pi27  & pi43 ;
  assign n10586 = ~n10584 & ~n10585;
  assign n10587 = n10582 & ~n10583;
  assign n10588 = ~n10586 & n10587;
  assign n10589 = n10582 & ~n10588;
  assign n10590 = ~n10583 & ~n10588;
  assign n10591 = ~n10586 & n10590;
  assign n10592 = ~n10589 & ~n10591;
  assign n10593 = ~n10581 & ~n10592;
  assign n10594 = ~n10581 & ~n10593;
  assign n10595 = ~n10592 & ~n10593;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = pi21  & pi49 ;
  assign n10598 = n1407 & n6114;
  assign n10599 = pi19  & pi51 ;
  assign n10600 = pi20  & pi50 ;
  assign n10601 = ~n10599 & ~n10600;
  assign n10602 = n10597 & ~n10598;
  assign n10603 = ~n10601 & n10602;
  assign n10604 = n10597 & ~n10603;
  assign n10605 = ~n10598 & ~n10603;
  assign n10606 = ~n10601 & n10605;
  assign n10607 = ~n10604 & ~n10606;
  assign n10608 = ~n10596 & ~n10607;
  assign n10609 = ~n10596 & ~n10608;
  assign n10610 = ~n10607 & ~n10608;
  assign n10611 = ~n10609 & ~n10610;
  assign n10612 = n10570 & ~n10611;
  assign n10613 = ~n10570 & n10611;
  assign n10614 = ~n10612 & ~n10613;
  assign n10615 = ~n10540 & n10614;
  assign n10616 = ~n10540 & ~n10615;
  assign n10617 = ~n10612 & ~n10615;
  assign n10618 = ~n10613 & n10617;
  assign n10619 = ~n10616 & ~n10618;
  assign n10620 = ~n10260 & ~n10263;
  assign n10621 = pi10  & pi60 ;
  assign n10622 = pi11  & pi59 ;
  assign n10623 = ~n10621 & ~n10622;
  assign n10624 = n1111 & n8854;
  assign n10625 = pi9  & pi61 ;
  assign n10626 = ~n10623 & n10625;
  assign n10627 = ~n10624 & n10626;
  assign n10628 = ~n10624 & ~n10627;
  assign n10629 = ~n10623 & n10628;
  assign n10630 = n10625 & ~n10627;
  assign n10631 = ~n10629 & ~n10630;
  assign n10632 = n989 & n8092;
  assign n10633 = pi17  & pi53 ;
  assign n10634 = pi16  & pi54 ;
  assign n10635 = ~n10633 & ~n10634;
  assign n10636 = n7680 & ~n10632;
  assign n10637 = ~n10635 & n10636;
  assign n10638 = n7680 & ~n10637;
  assign n10639 = ~n10632 & ~n10637;
  assign n10640 = ~n10635 & n10639;
  assign n10641 = ~n10638 & ~n10640;
  assign n10642 = ~n10631 & ~n10641;
  assign n10643 = ~n10631 & ~n10642;
  assign n10644 = ~n10641 & ~n10642;
  assign n10645 = ~n10643 & ~n10644;
  assign n10646 = pi12  & pi58 ;
  assign n10647 = n7611 & n9609;
  assign n10648 = pi13  & pi57 ;
  assign n10649 = ~n4881 & ~n10648;
  assign n10650 = n10646 & ~n10647;
  assign n10651 = ~n10649 & n10650;
  assign n10652 = n10646 & ~n10651;
  assign n10653 = ~n10647 & ~n10651;
  assign n10654 = ~n10649 & n10653;
  assign n10655 = ~n10652 & ~n10654;
  assign n10656 = ~n10645 & ~n10655;
  assign n10657 = ~n10645 & ~n10656;
  assign n10658 = ~n10655 & ~n10656;
  assign n10659 = ~n10657 & ~n10658;
  assign n10660 = n10324 & n10378;
  assign n10661 = ~n10324 & ~n10378;
  assign n10662 = ~n10660 & ~n10661;
  assign n10663 = pi32  & pi38 ;
  assign n10664 = n3900 & n4500;
  assign n10665 = pi34  & pi36 ;
  assign n10666 = pi33  & pi37 ;
  assign n10667 = ~n10665 & ~n10666;
  assign n10668 = n10663 & ~n10664;
  assign n10669 = ~n10667 & n10668;
  assign n10670 = n10663 & ~n10669;
  assign n10671 = ~n10664 & ~n10669;
  assign n10672 = ~n10667 & n10671;
  assign n10673 = ~n10670 & ~n10672;
  assign n10674 = n10662 & ~n10673;
  assign n10675 = n10662 & ~n10674;
  assign n10676 = ~n10673 & ~n10674;
  assign n10677 = ~n10675 & ~n10676;
  assign n10678 = ~n10255 & ~n10257;
  assign n10679 = ~n10677 & ~n10678;
  assign n10680 = n10677 & n10678;
  assign n10681 = ~n10679 & ~n10680;
  assign n10682 = ~n10659 & n10681;
  assign n10683 = n10659 & ~n10681;
  assign n10684 = ~n10682 & ~n10683;
  assign n10685 = ~n10620 & n10684;
  assign n10686 = n10620 & ~n10684;
  assign n10687 = ~n10685 & ~n10686;
  assign n10688 = ~n10619 & n10687;
  assign n10689 = ~n10619 & ~n10688;
  assign n10690 = n10687 & ~n10688;
  assign n10691 = ~n10689 & ~n10690;
  assign n10692 = ~n10539 & ~n10691;
  assign n10693 = ~n10539 & ~n10692;
  assign n10694 = ~n10691 & ~n10692;
  assign n10695 = ~n10693 & ~n10694;
  assign n10696 = ~n10298 & ~n10302;
  assign n10697 = ~n10441 & ~n10472;
  assign n10698 = ~n10273 & ~n10277;
  assign n10699 = n10405 & n10451;
  assign n10700 = ~n10405 & ~n10451;
  assign n10701 = ~n10699 & ~n10700;
  assign n10702 = n10466 & ~n10701;
  assign n10703 = ~n10466 & n10701;
  assign n10704 = ~n10702 & ~n10703;
  assign n10705 = ~n10280 & ~n10283;
  assign n10706 = ~n10247 & ~n10250;
  assign n10707 = n10705 & n10706;
  assign n10708 = ~n10705 & ~n10706;
  assign n10709 = ~n10707 & ~n10708;
  assign n10710 = n10704 & n10709;
  assign n10711 = ~n10704 & ~n10709;
  assign n10712 = ~n10710 & ~n10711;
  assign n10713 = ~n10698 & n10712;
  assign n10714 = ~n10698 & ~n10713;
  assign n10715 = n10712 & ~n10713;
  assign n10716 = ~n10714 & ~n10715;
  assign n10717 = ~n10697 & ~n10716;
  assign n10718 = ~n10697 & ~n10717;
  assign n10719 = ~n10716 & ~n10717;
  assign n10720 = ~n10718 & ~n10719;
  assign n10721 = ~n10696 & ~n10720;
  assign n10722 = ~n10696 & ~n10721;
  assign n10723 = ~n10720 & ~n10721;
  assign n10724 = ~n10722 & ~n10723;
  assign n10725 = ~n10394 & ~n10475;
  assign n10726 = n10724 & n10725;
  assign n10727 = ~n10724 & ~n10725;
  assign n10728 = ~n10726 & ~n10727;
  assign n10729 = ~n10313 & ~n10479;
  assign n10730 = n10728 & ~n10729;
  assign n10731 = n10728 & ~n10730;
  assign n10732 = ~n10729 & ~n10730;
  assign n10733 = ~n10731 & ~n10732;
  assign n10734 = ~n10695 & ~n10733;
  assign n10735 = n10695 & n10733;
  assign n10736 = ~n10734 & ~n10735;
  assign n10737 = n10495 & ~n10736;
  assign n10738 = ~n10495 & n10736;
  assign n10739 = ~n10737 & ~n10738;
  assign n10740 = ~n10488 & ~n10493;
  assign n10741 = ~n10739 & n10740;
  assign n10742 = ~n10737 & ~n10740;
  assign n10743 = ~n10738 & n10742;
  assign po71  = ~n10741 & ~n10743;
  assign n10745 = ~n10738 & ~n10742;
  assign n10746 = ~n10730 & ~n10734;
  assign n10747 = ~n10685 & ~n10688;
  assign n10748 = ~n10661 & ~n10674;
  assign n10749 = n10509 & n10748;
  assign n10750 = ~n10509 & ~n10748;
  assign n10751 = ~n10749 & ~n10750;
  assign n10752 = ~n10498 & ~n10501;
  assign n10753 = ~n10751 & n10752;
  assign n10754 = n10751 & ~n10752;
  assign n10755 = ~n10753 & ~n10754;
  assign n10756 = ~n10512 & ~n10518;
  assign n10757 = ~n10755 & n10756;
  assign n10758 = n10755 & ~n10756;
  assign n10759 = ~n10757 & ~n10758;
  assign n10760 = ~n10679 & ~n10682;
  assign n10761 = ~n10759 & n10760;
  assign n10762 = n10759 & ~n10760;
  assign n10763 = ~n10761 & ~n10762;
  assign n10764 = ~n10530 & ~n10534;
  assign n10765 = n10763 & ~n10764;
  assign n10766 = ~n10763 & n10764;
  assign n10767 = ~n10765 & ~n10766;
  assign n10768 = n10747 & ~n10767;
  assign n10769 = ~n10747 & n10767;
  assign n10770 = ~n10768 & ~n10769;
  assign n10771 = ~n10536 & ~n10692;
  assign n10772 = ~n10770 & n10771;
  assign n10773 = n10770 & ~n10771;
  assign n10774 = ~n10772 & ~n10773;
  assign n10775 = ~n10721 & ~n10727;
  assign n10776 = ~n10642 & ~n10656;
  assign n10777 = ~n10700 & ~n10703;
  assign n10778 = n10776 & n10777;
  assign n10779 = ~n10776 & ~n10777;
  assign n10780 = ~n10778 & ~n10779;
  assign n10781 = ~n10593 & ~n10608;
  assign n10782 = ~n10780 & n10781;
  assign n10783 = n10780 & ~n10781;
  assign n10784 = ~n10782 & ~n10783;
  assign n10785 = ~n10617 & n10784;
  assign n10786 = n10617 & ~n10784;
  assign n10787 = ~n10785 & ~n10786;
  assign n10788 = ~n10563 & ~n10569;
  assign n10789 = n10628 & n10653;
  assign n10790 = ~n10628 & ~n10653;
  assign n10791 = ~n10789 & ~n10790;
  assign n10792 = n10590 & ~n10791;
  assign n10793 = ~n10590 & n10791;
  assign n10794 = ~n10792 & ~n10793;
  assign n10795 = n10560 & n10578;
  assign n10796 = ~n10560 & ~n10578;
  assign n10797 = ~n10795 & ~n10796;
  assign n10798 = n10548 & ~n10797;
  assign n10799 = ~n10548 & n10797;
  assign n10800 = ~n10798 & ~n10799;
  assign n10801 = ~n10794 & ~n10800;
  assign n10802 = n10794 & n10800;
  assign n10803 = ~n10801 & ~n10802;
  assign n10804 = ~n10788 & n10803;
  assign n10805 = n10788 & ~n10803;
  assign n10806 = ~n10804 & ~n10805;
  assign n10807 = n10787 & n10806;
  assign n10808 = ~n10787 & ~n10806;
  assign n10809 = ~n10807 & ~n10808;
  assign n10810 = ~n10775 & n10809;
  assign n10811 = n10775 & ~n10809;
  assign n10812 = ~n10810 & ~n10811;
  assign n10813 = ~n10713 & ~n10717;
  assign n10814 = pi9  & pi62 ;
  assign n10815 = ~pi36  & ~n10814;
  assign n10816 = pi36  & pi62 ;
  assign n10817 = pi9  & n10816;
  assign n10818 = pi22  & pi49 ;
  assign n10819 = ~n10815 & n10818;
  assign n10820 = ~n10817 & n10819;
  assign n10821 = ~n10817 & ~n10820;
  assign n10822 = ~n10815 & n10821;
  assign n10823 = n10818 & ~n10820;
  assign n10824 = ~n10822 & ~n10823;
  assign n10825 = pi21  & pi50 ;
  assign n10826 = n1407 & n10319;
  assign n10827 = pi19  & pi52 ;
  assign n10828 = pi20  & pi51 ;
  assign n10829 = ~n10827 & ~n10828;
  assign n10830 = n10825 & ~n10826;
  assign n10831 = ~n10829 & n10830;
  assign n10832 = n10825 & ~n10831;
  assign n10833 = ~n10826 & ~n10831;
  assign n10834 = ~n10829 & n10833;
  assign n10835 = ~n10832 & ~n10834;
  assign n10836 = ~n10824 & ~n10835;
  assign n10837 = ~n10824 & ~n10836;
  assign n10838 = ~n10835 & ~n10836;
  assign n10839 = ~n10837 & ~n10838;
  assign n10840 = pi33  & pi38 ;
  assign n10841 = pi34  & pi37 ;
  assign n10842 = n4691 & n10841;
  assign n10843 = ~n4691 & ~n10841;
  assign n10844 = n10840 & ~n10842;
  assign n10845 = ~n10843 & n10844;
  assign n10846 = n10840 & ~n10845;
  assign n10847 = ~n10842 & ~n10845;
  assign n10848 = ~n10843 & n10847;
  assign n10849 = ~n10846 & ~n10848;
  assign n10850 = ~n10839 & ~n10849;
  assign n10851 = ~n10839 & ~n10850;
  assign n10852 = ~n10849 & ~n10850;
  assign n10853 = ~n10851 & ~n10852;
  assign n10854 = n10639 & n10671;
  assign n10855 = ~n10639 & ~n10671;
  assign n10856 = ~n10854 & ~n10855;
  assign n10857 = pi11  & pi60 ;
  assign n10858 = n855 & n9236;
  assign n10859 = pi8  & pi63 ;
  assign n10860 = pi10  & pi61 ;
  assign n10861 = ~n10859 & ~n10860;
  assign n10862 = n10857 & ~n10858;
  assign n10863 = ~n10861 & n10862;
  assign n10864 = n10857 & ~n10863;
  assign n10865 = ~n10858 & ~n10863;
  assign n10866 = ~n10861 & n10865;
  assign n10867 = ~n10864 & ~n10866;
  assign n10868 = n10856 & ~n10867;
  assign n10869 = n10856 & ~n10868;
  assign n10870 = ~n10867 & ~n10868;
  assign n10871 = ~n10869 & ~n10870;
  assign n10872 = ~n10708 & ~n10710;
  assign n10873 = ~n10871 & ~n10872;
  assign n10874 = n10871 & n10872;
  assign n10875 = ~n10873 & ~n10874;
  assign n10876 = ~n10853 & n10875;
  assign n10877 = n10853 & ~n10875;
  assign n10878 = ~n10876 & ~n10877;
  assign n10879 = ~n10813 & n10878;
  assign n10880 = n10813 & ~n10878;
  assign n10881 = ~n10879 & ~n10880;
  assign n10882 = ~n10524 & ~n10528;
  assign n10883 = pi28  & pi43 ;
  assign n10884 = pi29  & pi42 ;
  assign n10885 = ~n10883 & ~n10884;
  assign n10886 = n2915 & n6458;
  assign n10887 = pi27  & pi44 ;
  assign n10888 = ~n10885 & n10887;
  assign n10889 = ~n10886 & n10888;
  assign n10890 = ~n10886 & ~n10889;
  assign n10891 = ~n10885 & n10890;
  assign n10892 = n10887 & ~n10889;
  assign n10893 = ~n10891 & ~n10892;
  assign n10894 = pi30  & pi41 ;
  assign n10895 = n3567 & n5548;
  assign n10896 = pi31  & pi40 ;
  assign n10897 = pi32  & pi39 ;
  assign n10898 = ~n10896 & ~n10897;
  assign n10899 = n10894 & ~n10895;
  assign n10900 = ~n10898 & n10899;
  assign n10901 = n10894 & ~n10900;
  assign n10902 = ~n10895 & ~n10900;
  assign n10903 = ~n10898 & n10902;
  assign n10904 = ~n10901 & ~n10903;
  assign n10905 = ~n10893 & ~n10904;
  assign n10906 = ~n10893 & ~n10905;
  assign n10907 = ~n10904 & ~n10905;
  assign n10908 = ~n10906 & ~n10907;
  assign n10909 = pi23  & pi48 ;
  assign n10910 = n1199 & n8092;
  assign n10911 = pi18  & pi53 ;
  assign n10912 = pi17  & pi54 ;
  assign n10913 = ~n10911 & ~n10912;
  assign n10914 = n10909 & ~n10910;
  assign n10915 = ~n10913 & n10914;
  assign n10916 = n10909 & ~n10915;
  assign n10917 = ~n10910 & ~n10915;
  assign n10918 = ~n10913 & n10917;
  assign n10919 = ~n10916 & ~n10918;
  assign n10920 = ~n10908 & ~n10919;
  assign n10921 = ~n10908 & ~n10920;
  assign n10922 = ~n10919 & ~n10920;
  assign n10923 = ~n10921 & ~n10922;
  assign n10924 = n952 & n9402;
  assign n10925 = pi13  & pi58 ;
  assign n10926 = ~n10924 & n10925;
  assign n10927 = pi12  & pi59 ;
  assign n10928 = ~n10924 & n10927;
  assign n10929 = ~n10926 & ~n10928;
  assign n10930 = ~n10605 & ~n10929;
  assign n10931 = ~n10605 & ~n10930;
  assign n10932 = ~n10929 & ~n10930;
  assign n10933 = ~n10931 & ~n10932;
  assign n10934 = pi15  & pi56 ;
  assign n10935 = pi16  & pi55 ;
  assign n10936 = ~n10934 & ~n10935;
  assign n10937 = n840 & n8521;
  assign n10938 = pi14  & pi57 ;
  assign n10939 = ~n10936 & n10938;
  assign n10940 = ~n10937 & n10939;
  assign n10941 = ~n10937 & ~n10940;
  assign n10942 = ~n10936 & n10941;
  assign n10943 = n10938 & ~n10940;
  assign n10944 = ~n10942 & ~n10943;
  assign n10945 = pi24  & pi47 ;
  assign n10946 = n2310 & n7513;
  assign n10947 = pi25  & pi46 ;
  assign n10948 = pi26  & pi45 ;
  assign n10949 = ~n10947 & ~n10948;
  assign n10950 = n10945 & ~n10946;
  assign n10951 = ~n10949 & n10950;
  assign n10952 = n10945 & ~n10951;
  assign n10953 = ~n10946 & ~n10951;
  assign n10954 = ~n10949 & n10953;
  assign n10955 = ~n10952 & ~n10954;
  assign n10956 = ~n10944 & ~n10955;
  assign n10957 = ~n10944 & ~n10956;
  assign n10958 = ~n10955 & ~n10956;
  assign n10959 = ~n10957 & ~n10958;
  assign n10960 = ~n10933 & n10959;
  assign n10961 = n10933 & ~n10959;
  assign n10962 = ~n10960 & ~n10961;
  assign n10963 = ~n10923 & ~n10962;
  assign n10964 = n10923 & n10962;
  assign n10965 = ~n10963 & ~n10964;
  assign n10966 = ~n10882 & n10965;
  assign n10967 = n10882 & ~n10965;
  assign n10968 = ~n10966 & ~n10967;
  assign n10969 = n10881 & n10968;
  assign n10970 = ~n10881 & ~n10968;
  assign n10971 = ~n10969 & ~n10970;
  assign n10972 = n10812 & n10971;
  assign n10973 = ~n10812 & ~n10971;
  assign n10974 = ~n10972 & ~n10973;
  assign n10975 = ~n10774 & ~n10974;
  assign n10976 = n10774 & n10974;
  assign n10977 = ~n10975 & ~n10976;
  assign n10978 = n10746 & ~n10977;
  assign n10979 = ~n10746 & n10977;
  assign n10980 = ~n10978 & ~n10979;
  assign n10981 = ~n10745 & ~n10980;
  assign n10982 = n10745 & n10980;
  assign po72  = n10981 | n10982;
  assign n10984 = ~n10745 & ~n10978;
  assign n10985 = ~n10979 & ~n10984;
  assign n10986 = ~n10879 & ~n10969;
  assign n10987 = ~n10802 & ~n10804;
  assign n10988 = ~n10855 & ~n10868;
  assign n10989 = pi29  & pi43 ;
  assign n10990 = n2680 & n5235;
  assign n10991 = pi30  & pi42 ;
  assign n10992 = ~n4626 & ~n10991;
  assign n10993 = n10989 & ~n10990;
  assign n10994 = ~n10992 & n10993;
  assign n10995 = n10989 & ~n10994;
  assign n10996 = ~n10990 & ~n10994;
  assign n10997 = ~n10992 & n10996;
  assign n10998 = ~n10995 & ~n10997;
  assign n10999 = ~n10988 & ~n10998;
  assign n11000 = ~n10988 & ~n10999;
  assign n11001 = ~n10998 & ~n10999;
  assign n11002 = ~n11000 & ~n11001;
  assign n11003 = ~n10796 & ~n10799;
  assign n11004 = n11002 & n11003;
  assign n11005 = ~n11002 & ~n11003;
  assign n11006 = ~n11004 & ~n11005;
  assign n11007 = ~n10987 & n11006;
  assign n11008 = n10987 & ~n11006;
  assign n11009 = ~n11007 & ~n11008;
  assign n11010 = ~n10873 & ~n10876;
  assign n11011 = ~n11009 & n11010;
  assign n11012 = n11009 & ~n11010;
  assign n11013 = ~n11011 & ~n11012;
  assign n11014 = ~n10785 & ~n10807;
  assign n11015 = n11013 & ~n11014;
  assign n11016 = ~n11013 & n11014;
  assign n11017 = ~n11015 & ~n11016;
  assign n11018 = n10986 & ~n11017;
  assign n11019 = ~n10986 & n11017;
  assign n11020 = ~n11018 & ~n11019;
  assign n11021 = ~n10810 & ~n10972;
  assign n11022 = ~n11020 & n11021;
  assign n11023 = n11020 & ~n11021;
  assign n11024 = ~n11022 & ~n11023;
  assign n11025 = ~n10765 & ~n10769;
  assign n11026 = ~n10905 & ~n10920;
  assign n11027 = ~n10790 & ~n10793;
  assign n11028 = n11026 & n11027;
  assign n11029 = ~n11026 & ~n11027;
  assign n11030 = ~n11028 & ~n11029;
  assign n11031 = ~n10836 & ~n10850;
  assign n11032 = ~n11030 & n11031;
  assign n11033 = n11030 & ~n11031;
  assign n11034 = ~n11032 & ~n11033;
  assign n11035 = ~n10963 & ~n10966;
  assign n11036 = ~n11034 & n11035;
  assign n11037 = n11034 & ~n11035;
  assign n11038 = ~n11036 & ~n11037;
  assign n11039 = ~n10933 & ~n10959;
  assign n11040 = ~n10956 & ~n11039;
  assign n11041 = n10890 & n10917;
  assign n11042 = ~n10890 & ~n10917;
  assign n11043 = ~n11041 & ~n11042;
  assign n11044 = n10902 & ~n11043;
  assign n11045 = ~n10902 & n11043;
  assign n11046 = ~n11044 & ~n11045;
  assign n11047 = n10821 & n10847;
  assign n11048 = ~n10821 & ~n10847;
  assign n11049 = ~n11047 & ~n11048;
  assign n11050 = n10833 & ~n11049;
  assign n11051 = ~n10833 & n11049;
  assign n11052 = ~n11050 & ~n11051;
  assign n11053 = n11046 & n11052;
  assign n11054 = ~n11046 & ~n11052;
  assign n11055 = ~n11053 & ~n11054;
  assign n11056 = ~n11040 & n11055;
  assign n11057 = n11040 & ~n11055;
  assign n11058 = ~n11056 & ~n11057;
  assign n11059 = n11038 & n11058;
  assign n11060 = ~n11038 & ~n11058;
  assign n11061 = ~n11059 & ~n11060;
  assign n11062 = n11025 & ~n11061;
  assign n11063 = ~n11025 & n11061;
  assign n11064 = ~n11062 & ~n11063;
  assign n11065 = ~n10779 & ~n10783;
  assign n11066 = pi16  & pi56 ;
  assign n11067 = pi23  & pi49 ;
  assign n11068 = ~n11066 & ~n11067;
  assign n11069 = n11066 & n11067;
  assign n11070 = pi32  & pi40 ;
  assign n11071 = ~n11068 & n11070;
  assign n11072 = ~n11069 & n11071;
  assign n11073 = ~n11069 & ~n11072;
  assign n11074 = ~n11068 & n11073;
  assign n11075 = n11070 & ~n11072;
  assign n11076 = ~n11074 & ~n11075;
  assign n11077 = pi35  & pi37 ;
  assign n11078 = n1481 & n6114;
  assign n11079 = pi21  & pi51 ;
  assign n11080 = pi22  & pi50 ;
  assign n11081 = ~n11079 & ~n11080;
  assign n11082 = n11077 & ~n11078;
  assign n11083 = ~n11081 & n11082;
  assign n11084 = n11077 & ~n11083;
  assign n11085 = ~n11078 & ~n11083;
  assign n11086 = ~n11081 & n11085;
  assign n11087 = ~n11084 & ~n11086;
  assign n11088 = ~n11076 & ~n11087;
  assign n11089 = ~n11076 & ~n11088;
  assign n11090 = ~n11087 & ~n11088;
  assign n11091 = ~n11089 & ~n11090;
  assign n11092 = pi17  & pi55 ;
  assign n11093 = pi52  & pi54 ;
  assign n11094 = n1257 & n11093;
  assign n11095 = pi20  & pi52 ;
  assign n11096 = ~n8411 & ~n11095;
  assign n11097 = n11092 & ~n11094;
  assign n11098 = ~n11096 & n11097;
  assign n11099 = n11092 & ~n11098;
  assign n11100 = ~n11094 & ~n11098;
  assign n11101 = ~n11096 & n11100;
  assign n11102 = ~n11099 & ~n11101;
  assign n11103 = ~n11091 & ~n11102;
  assign n11104 = ~n11091 & ~n11103;
  assign n11105 = ~n11102 & ~n11103;
  assign n11106 = ~n11104 & ~n11105;
  assign n11107 = pi10  & pi62 ;
  assign n11108 = pi11  & pi61 ;
  assign n11109 = ~n11107 & ~n11108;
  assign n11110 = n1111 & n9567;
  assign n11111 = pi9  & pi63 ;
  assign n11112 = ~n11109 & n11111;
  assign n11113 = ~n11110 & n11112;
  assign n11114 = ~n11110 & ~n11113;
  assign n11115 = ~n11109 & n11114;
  assign n11116 = n11111 & ~n11113;
  assign n11117 = ~n11115 & ~n11116;
  assign n11118 = ~n10924 & ~n10930;
  assign n11119 = pi12  & pi60 ;
  assign n11120 = n1789 & n5823;
  assign n11121 = pi24  & pi48 ;
  assign n11122 = pi25  & pi47 ;
  assign n11123 = ~n11121 & ~n11122;
  assign n11124 = n11119 & ~n11120;
  assign n11125 = ~n11123 & n11124;
  assign n11126 = n11119 & ~n11125;
  assign n11127 = ~n11120 & ~n11125;
  assign n11128 = ~n11123 & n11127;
  assign n11129 = ~n11126 & ~n11128;
  assign n11130 = ~n11118 & ~n11129;
  assign n11131 = ~n11118 & ~n11130;
  assign n11132 = ~n11129 & ~n11130;
  assign n11133 = ~n11131 & ~n11132;
  assign n11134 = ~n11117 & ~n11133;
  assign n11135 = n11117 & n11133;
  assign n11136 = ~n11134 & ~n11135;
  assign n11137 = ~n11106 & n11136;
  assign n11138 = n11106 & ~n11136;
  assign n11139 = ~n11137 & ~n11138;
  assign n11140 = ~n11065 & n11139;
  assign n11141 = n11065 & ~n11139;
  assign n11142 = ~n11140 & ~n11141;
  assign n11143 = ~n10758 & ~n10762;
  assign n11144 = n10941 & n10953;
  assign n11145 = ~n10941 & ~n10953;
  assign n11146 = ~n11144 & ~n11145;
  assign n11147 = n10865 & ~n11146;
  assign n11148 = ~n10865 & n11146;
  assign n11149 = ~n11147 & ~n11148;
  assign n11150 = ~n10750 & ~n10754;
  assign n11151 = ~n11149 & n11150;
  assign n11152 = n11149 & ~n11150;
  assign n11153 = ~n11151 & ~n11152;
  assign n11154 = pi14  & pi58 ;
  assign n11155 = pi15  & pi57 ;
  assign n11156 = ~n11154 & ~n11155;
  assign n11157 = n1041 & n8144;
  assign n11158 = pi13  & pi59 ;
  assign n11159 = ~n11156 & n11158;
  assign n11160 = ~n11157 & n11159;
  assign n11161 = ~n11157 & ~n11160;
  assign n11162 = ~n11156 & n11161;
  assign n11163 = n11158 & ~n11160;
  assign n11164 = ~n11162 & ~n11163;
  assign n11165 = pi26  & pi46 ;
  assign n11166 = n2191 & n5318;
  assign n11167 = pi27  & pi45 ;
  assign n11168 = pi28  & pi44 ;
  assign n11169 = ~n11167 & ~n11168;
  assign n11170 = n11165 & ~n11166;
  assign n11171 = ~n11169 & n11170;
  assign n11172 = n11165 & ~n11171;
  assign n11173 = ~n11166 & ~n11171;
  assign n11174 = ~n11169 & n11173;
  assign n11175 = ~n11172 & ~n11174;
  assign n11176 = ~n11164 & ~n11175;
  assign n11177 = ~n11164 & ~n11176;
  assign n11178 = ~n11175 & ~n11176;
  assign n11179 = ~n11177 & ~n11178;
  assign n11180 = pi19  & pi53 ;
  assign n11181 = n3900 & n4736;
  assign n11182 = pi34  & pi38 ;
  assign n11183 = pi33  & pi39 ;
  assign n11184 = ~n11182 & ~n11183;
  assign n11185 = n11180 & ~n11181;
  assign n11186 = ~n11184 & n11185;
  assign n11187 = n11180 & ~n11186;
  assign n11188 = ~n11181 & ~n11186;
  assign n11189 = ~n11184 & n11188;
  assign n11190 = ~n11187 & ~n11189;
  assign n11191 = ~n11179 & ~n11190;
  assign n11192 = ~n11179 & ~n11191;
  assign n11193 = ~n11190 & ~n11191;
  assign n11194 = ~n11192 & ~n11193;
  assign n11195 = ~n11153 & n11194;
  assign n11196 = n11153 & ~n11194;
  assign n11197 = ~n11195 & ~n11196;
  assign n11198 = ~n11143 & n11197;
  assign n11199 = ~n11143 & ~n11198;
  assign n11200 = n11197 & ~n11198;
  assign n11201 = ~n11199 & ~n11200;
  assign n11202 = n11142 & ~n11201;
  assign n11203 = n11142 & ~n11202;
  assign n11204 = ~n11201 & ~n11202;
  assign n11205 = ~n11203 & ~n11204;
  assign n11206 = n11064 & ~n11205;
  assign n11207 = n11064 & ~n11206;
  assign n11208 = ~n11205 & ~n11206;
  assign n11209 = ~n11207 & ~n11208;
  assign n11210 = ~n11024 & n11209;
  assign n11211 = n11024 & ~n11209;
  assign n11212 = ~n11210 & ~n11211;
  assign n11213 = ~n10773 & ~n10976;
  assign n11214 = ~n11212 & n11213;
  assign n11215 = n11212 & ~n11213;
  assign n11216 = ~n11214 & ~n11215;
  assign n11217 = n10985 & ~n11216;
  assign n11218 = ~n10985 & ~n11214;
  assign n11219 = ~n11215 & n11218;
  assign po73  = ~n11217 & ~n11219;
  assign n11221 = ~n11215 & ~n11218;
  assign n11222 = ~n11023 & ~n11211;
  assign n11223 = ~n11063 & ~n11206;
  assign n11224 = ~n11198 & ~n11202;
  assign n11225 = ~n11037 & ~n11059;
  assign n11226 = ~n11152 & ~n11196;
  assign n11227 = ~n11145 & ~n11148;
  assign n11228 = pi31  & pi42 ;
  assign n11229 = n6012 & n6138;
  assign n11230 = pi32  & pi41 ;
  assign n11231 = pi33  & pi40 ;
  assign n11232 = ~n11230 & ~n11231;
  assign n11233 = n11228 & ~n11229;
  assign n11234 = ~n11232 & n11233;
  assign n11235 = n11228 & ~n11234;
  assign n11236 = ~n11229 & ~n11234;
  assign n11237 = ~n11232 & n11236;
  assign n11238 = ~n11235 & ~n11237;
  assign n11239 = ~n11227 & ~n11238;
  assign n11240 = ~n11227 & ~n11239;
  assign n11241 = ~n11238 & ~n11239;
  assign n11242 = ~n11240 & ~n11241;
  assign n11243 = ~n11042 & ~n11045;
  assign n11244 = n11242 & n11243;
  assign n11245 = ~n11242 & ~n11243;
  assign n11246 = ~n11244 & ~n11245;
  assign n11247 = ~n11053 & ~n11056;
  assign n11248 = n11246 & ~n11247;
  assign n11249 = ~n11246 & n11247;
  assign n11250 = ~n11248 & ~n11249;
  assign n11251 = ~n11226 & n11250;
  assign n11252 = n11226 & ~n11250;
  assign n11253 = ~n11251 & ~n11252;
  assign n11254 = ~n11225 & n11253;
  assign n11255 = n11225 & ~n11253;
  assign n11256 = ~n11254 & ~n11255;
  assign n11257 = ~n11224 & n11256;
  assign n11258 = n11224 & ~n11256;
  assign n11259 = ~n11257 & ~n11258;
  assign n11260 = n11223 & ~n11259;
  assign n11261 = ~n11223 & n11259;
  assign n11262 = ~n11260 & ~n11261;
  assign n11263 = ~n11015 & ~n11019;
  assign n11264 = ~n11130 & ~n11134;
  assign n11265 = ~n11048 & ~n11051;
  assign n11266 = n11264 & n11265;
  assign n11267 = ~n11264 & ~n11265;
  assign n11268 = ~n11266 & ~n11267;
  assign n11269 = ~n11176 & ~n11191;
  assign n11270 = ~n11268 & n11269;
  assign n11271 = n11268 & ~n11269;
  assign n11272 = ~n11270 & ~n11271;
  assign n11273 = ~n11137 & ~n11140;
  assign n11274 = ~n11272 & n11273;
  assign n11275 = n11272 & ~n11273;
  assign n11276 = ~n11274 & ~n11275;
  assign n11277 = ~n11088 & ~n11103;
  assign n11278 = pi13  & pi60 ;
  assign n11279 = ~n11085 & n11278;
  assign n11280 = n11085 & ~n11278;
  assign n11281 = ~n11279 & ~n11280;
  assign n11282 = n11188 & ~n11281;
  assign n11283 = ~n11188 & n11281;
  assign n11284 = ~n11282 & ~n11283;
  assign n11285 = n11114 & n11127;
  assign n11286 = ~n11114 & ~n11127;
  assign n11287 = ~n11285 & ~n11286;
  assign n11288 = n11100 & ~n11287;
  assign n11289 = ~n11100 & n11287;
  assign n11290 = ~n11288 & ~n11289;
  assign n11291 = n11284 & n11290;
  assign n11292 = ~n11284 & ~n11290;
  assign n11293 = ~n11291 & ~n11292;
  assign n11294 = ~n11277 & n11293;
  assign n11295 = n11277 & ~n11293;
  assign n11296 = ~n11294 & ~n11295;
  assign n11297 = n11276 & n11296;
  assign n11298 = ~n11276 & ~n11296;
  assign n11299 = ~n11297 & ~n11298;
  assign n11300 = n11263 & ~n11299;
  assign n11301 = ~n11263 & n11299;
  assign n11302 = ~n11300 & ~n11301;
  assign n11303 = pi11  & pi62 ;
  assign n11304 = ~pi37  & ~n11303;
  assign n11305 = pi62  & n4258;
  assign n11306 = pi23  & pi50 ;
  assign n11307 = ~n11304 & n11306;
  assign n11308 = ~n11305 & n11307;
  assign n11309 = ~n11305 & ~n11308;
  assign n11310 = ~n11304 & n11309;
  assign n11311 = n11306 & ~n11308;
  assign n11312 = ~n11310 & ~n11311;
  assign n11313 = pi18  & pi55 ;
  assign n11314 = pi49  & pi54 ;
  assign n11315 = n4106 & n11314;
  assign n11316 = pi19  & pi54 ;
  assign n11317 = pi24  & pi49 ;
  assign n11318 = ~n11316 & ~n11317;
  assign n11319 = n11313 & ~n11315;
  assign n11320 = ~n11318 & n11319;
  assign n11321 = n11313 & ~n11320;
  assign n11322 = ~n11315 & ~n11320;
  assign n11323 = ~n11318 & n11322;
  assign n11324 = ~n11321 & ~n11323;
  assign n11325 = ~n11312 & ~n11324;
  assign n11326 = ~n11312 & ~n11325;
  assign n11327 = ~n11324 & ~n11325;
  assign n11328 = ~n11326 & ~n11327;
  assign n11329 = pi22  & pi51 ;
  assign n11330 = n1593 & n9144;
  assign n11331 = pi20  & pi53 ;
  assign n11332 = pi21  & pi52 ;
  assign n11333 = ~n11331 & ~n11332;
  assign n11334 = n11329 & ~n11330;
  assign n11335 = ~n11333 & n11334;
  assign n11336 = n11329 & ~n11335;
  assign n11337 = ~n11330 & ~n11335;
  assign n11338 = ~n11333 & n11337;
  assign n11339 = ~n11336 & ~n11338;
  assign n11340 = ~n11328 & ~n11339;
  assign n11341 = ~n11328 & ~n11340;
  assign n11342 = ~n11339 & ~n11340;
  assign n11343 = ~n11341 & ~n11342;
  assign n11344 = pi15  & pi58 ;
  assign n11345 = pi16  & pi57 ;
  assign n11346 = ~n11344 & ~n11345;
  assign n11347 = n840 & n8144;
  assign n11348 = pi14  & pi59 ;
  assign n11349 = ~n11346 & n11348;
  assign n11350 = ~n11347 & n11349;
  assign n11351 = ~n11347 & ~n11350;
  assign n11352 = ~n11346 & n11351;
  assign n11353 = n11348 & ~n11350;
  assign n11354 = ~n11352 & ~n11353;
  assign n11355 = pi17  & pi56 ;
  assign n11356 = n2646 & n5277;
  assign n11357 = pi26  & pi47 ;
  assign n11358 = pi27  & pi46 ;
  assign n11359 = ~n11357 & ~n11358;
  assign n11360 = n11355 & ~n11356;
  assign n11361 = ~n11359 & n11360;
  assign n11362 = n11355 & ~n11361;
  assign n11363 = ~n11356 & ~n11361;
  assign n11364 = ~n11359 & n11363;
  assign n11365 = ~n11362 & ~n11364;
  assign n11366 = ~n11073 & ~n11365;
  assign n11367 = n11073 & n11365;
  assign n11368 = ~n11366 & ~n11367;
  assign n11369 = ~n11354 & n11368;
  assign n11370 = ~n11354 & ~n11369;
  assign n11371 = n11368 & ~n11369;
  assign n11372 = ~n11370 & ~n11371;
  assign n11373 = ~n11343 & ~n11372;
  assign n11374 = ~n11343 & ~n11373;
  assign n11375 = ~n11372 & ~n11373;
  assign n11376 = ~n11374 & ~n11375;
  assign n11377 = ~n11029 & ~n11033;
  assign n11378 = n11376 & n11377;
  assign n11379 = ~n11376 & ~n11377;
  assign n11380 = ~n11378 & ~n11379;
  assign n11381 = ~n11007 & ~n11012;
  assign n11382 = n11161 & n11173;
  assign n11383 = ~n11161 & ~n11173;
  assign n11384 = ~n11382 & ~n11383;
  assign n11385 = n10996 & ~n11384;
  assign n11386 = ~n10996 & n11384;
  assign n11387 = ~n11385 & ~n11386;
  assign n11388 = ~n10999 & ~n11005;
  assign n11389 = ~n11387 & n11388;
  assign n11390 = n11387 & ~n11388;
  assign n11391 = ~n11389 & ~n11390;
  assign n11392 = pi10  & pi63 ;
  assign n11393 = pi12  & pi61 ;
  assign n11394 = ~n11392 & ~n11393;
  assign n11395 = n460 & n9236;
  assign n11396 = pi25  & pi48 ;
  assign n11397 = ~n11394 & n11396;
  assign n11398 = ~n11395 & n11397;
  assign n11399 = ~n11395 & ~n11398;
  assign n11400 = ~n11394 & n11399;
  assign n11401 = n11396 & ~n11398;
  assign n11402 = ~n11400 & ~n11401;
  assign n11403 = pi28  & pi45 ;
  assign n11404 = n4908 & n6836;
  assign n11405 = pi29  & pi44 ;
  assign n11406 = pi30  & pi43 ;
  assign n11407 = ~n11405 & ~n11406;
  assign n11408 = n11403 & ~n11404;
  assign n11409 = ~n11407 & n11408;
  assign n11410 = n11403 & ~n11409;
  assign n11411 = ~n11404 & ~n11409;
  assign n11412 = ~n11407 & n11411;
  assign n11413 = ~n11410 & ~n11412;
  assign n11414 = ~n11402 & ~n11413;
  assign n11415 = ~n11402 & ~n11414;
  assign n11416 = ~n11413 & ~n11414;
  assign n11417 = ~n11415 & ~n11416;
  assign n11418 = n4691 & n5055;
  assign n11419 = pi35  & pi38 ;
  assign n11420 = ~n4500 & ~n11419;
  assign n11421 = n4434 & ~n11418;
  assign n11422 = ~n11420 & n11421;
  assign n11423 = n4434 & ~n11422;
  assign n11424 = ~n11418 & ~n11422;
  assign n11425 = ~n11420 & n11424;
  assign n11426 = ~n11423 & ~n11425;
  assign n11427 = ~n11417 & ~n11426;
  assign n11428 = ~n11417 & ~n11427;
  assign n11429 = ~n11426 & ~n11427;
  assign n11430 = ~n11428 & ~n11429;
  assign n11431 = ~n11391 & n11430;
  assign n11432 = n11391 & ~n11430;
  assign n11433 = ~n11431 & ~n11432;
  assign n11434 = ~n11381 & n11433;
  assign n11435 = ~n11381 & ~n11434;
  assign n11436 = n11433 & ~n11434;
  assign n11437 = ~n11435 & ~n11436;
  assign n11438 = n11380 & ~n11437;
  assign n11439 = n11380 & ~n11438;
  assign n11440 = ~n11437 & ~n11438;
  assign n11441 = ~n11439 & ~n11440;
  assign n11442 = n11302 & ~n11441;
  assign n11443 = n11302 & ~n11442;
  assign n11444 = ~n11441 & ~n11442;
  assign n11445 = ~n11443 & ~n11444;
  assign n11446 = ~n11262 & n11445;
  assign n11447 = n11262 & ~n11445;
  assign n11448 = ~n11446 & ~n11447;
  assign n11449 = n11222 & ~n11448;
  assign n11450 = ~n11222 & n11448;
  assign n11451 = ~n11449 & ~n11450;
  assign n11452 = ~n11221 & ~n11451;
  assign n11453 = n11221 & n11451;
  assign po74  = n11452 | n11453;
  assign n11455 = ~n11261 & ~n11447;
  assign n11456 = ~n11254 & ~n11257;
  assign n11457 = n11236 & n11424;
  assign n11458 = ~n11236 & ~n11424;
  assign n11459 = ~n11457 & ~n11458;
  assign n11460 = pi14  & pi60 ;
  assign n11461 = n840 & n9402;
  assign n11462 = pi15  & pi59 ;
  assign n11463 = pi16  & pi58 ;
  assign n11464 = ~n11462 & ~n11463;
  assign n11465 = n11460 & ~n11461;
  assign n11466 = ~n11464 & n11465;
  assign n11467 = n11460 & ~n11466;
  assign n11468 = ~n11461 & ~n11466;
  assign n11469 = ~n11464 & n11468;
  assign n11470 = ~n11467 & ~n11469;
  assign n11471 = n11459 & ~n11470;
  assign n11472 = n11459 & ~n11471;
  assign n11473 = ~n11470 & ~n11471;
  assign n11474 = ~n11472 & ~n11473;
  assign n11475 = ~n11325 & ~n11340;
  assign n11476 = n11474 & n11475;
  assign n11477 = ~n11474 & ~n11475;
  assign n11478 = ~n11476 & ~n11477;
  assign n11479 = ~n11239 & ~n11245;
  assign n11480 = ~n11478 & n11479;
  assign n11481 = n11478 & ~n11479;
  assign n11482 = ~n11480 & ~n11481;
  assign n11483 = ~n11373 & ~n11379;
  assign n11484 = ~n11390 & ~n11432;
  assign n11485 = ~n11483 & ~n11484;
  assign n11486 = ~n11483 & ~n11485;
  assign n11487 = ~n11484 & ~n11485;
  assign n11488 = ~n11486 & ~n11487;
  assign n11489 = n11482 & ~n11488;
  assign n11490 = ~n11482 & n11488;
  assign n11491 = ~n11489 & ~n11490;
  assign n11492 = ~n11456 & n11491;
  assign n11493 = ~n11456 & ~n11492;
  assign n11494 = n11491 & ~n11492;
  assign n11495 = ~n11493 & ~n11494;
  assign n11496 = ~n11248 & ~n11251;
  assign n11497 = n11363 & n11411;
  assign n11498 = ~n11363 & ~n11411;
  assign n11499 = ~n11497 & ~n11498;
  assign n11500 = n11351 & ~n11499;
  assign n11501 = ~n11351 & n11499;
  assign n11502 = ~n11500 & ~n11501;
  assign n11503 = n11322 & n11337;
  assign n11504 = ~n11322 & ~n11337;
  assign n11505 = ~n11503 & ~n11504;
  assign n11506 = n11399 & ~n11505;
  assign n11507 = ~n11399 & n11505;
  assign n11508 = ~n11506 & ~n11507;
  assign n11509 = ~n11414 & ~n11427;
  assign n11510 = ~n11508 & n11509;
  assign n11511 = n11508 & ~n11509;
  assign n11512 = ~n11510 & ~n11511;
  assign n11513 = n11502 & n11512;
  assign n11514 = ~n11502 & ~n11512;
  assign n11515 = ~n11513 & ~n11514;
  assign n11516 = ~n11496 & n11515;
  assign n11517 = n11496 & ~n11515;
  assign n11518 = ~n11516 & ~n11517;
  assign n11519 = n952 & n9567;
  assign n11520 = pi13  & pi61 ;
  assign n11521 = ~n11519 & n11520;
  assign n11522 = pi12  & pi62 ;
  assign n11523 = ~n11519 & n11522;
  assign n11524 = ~n11521 & ~n11523;
  assign n11525 = ~n11309 & ~n11524;
  assign n11526 = ~n11309 & ~n11525;
  assign n11527 = ~n11524 & ~n11525;
  assign n11528 = ~n11526 & ~n11527;
  assign n11529 = pi29  & pi45 ;
  assign n11530 = pi30  & pi44 ;
  assign n11531 = n8959 & n11530;
  assign n11532 = ~n8959 & ~n11530;
  assign n11533 = n11529 & ~n11531;
  assign n11534 = ~n11532 & n11533;
  assign n11535 = n11529 & ~n11534;
  assign n11536 = ~n11531 & ~n11534;
  assign n11537 = ~n11532 & n11536;
  assign n11538 = ~n11535 & ~n11537;
  assign n11539 = ~n11528 & ~n11538;
  assign n11540 = ~n11528 & ~n11539;
  assign n11541 = ~n11538 & ~n11539;
  assign n11542 = ~n11540 & ~n11541;
  assign n11543 = ~n11383 & ~n11386;
  assign n11544 = n11542 & n11543;
  assign n11545 = ~n11542 & ~n11543;
  assign n11546 = ~n11544 & ~n11545;
  assign n11547 = pi31  & pi43 ;
  assign n11548 = pi32  & pi42 ;
  assign n11549 = ~n11547 & ~n11548;
  assign n11550 = n3567 & n6458;
  assign n11551 = pi11  & pi63 ;
  assign n11552 = ~n11549 & n11551;
  assign n11553 = ~n11550 & n11552;
  assign n11554 = ~n11550 & ~n11553;
  assign n11555 = ~n11549 & n11554;
  assign n11556 = n11551 & ~n11553;
  assign n11557 = ~n11555 & ~n11556;
  assign n11558 = pi25  & pi56 ;
  assign n11559 = n9869 & n11558;
  assign n11560 = pi18  & pi56 ;
  assign n11561 = pi25  & pi49 ;
  assign n11562 = ~n11560 & ~n11561;
  assign n11563 = n4982 & ~n11559;
  assign n11564 = ~n11562 & n11563;
  assign n11565 = n4982 & ~n11564;
  assign n11566 = ~n11559 & ~n11564;
  assign n11567 = ~n11562 & n11566;
  assign n11568 = ~n11565 & ~n11567;
  assign n11569 = ~n11557 & ~n11568;
  assign n11570 = ~n11557 & ~n11569;
  assign n11571 = ~n11568 & ~n11569;
  assign n11572 = ~n11570 & ~n11571;
  assign n11573 = pi26  & pi48 ;
  assign n11574 = n2191 & n5277;
  assign n11575 = pi27  & pi47 ;
  assign n11576 = pi28  & pi46 ;
  assign n11577 = ~n11575 & ~n11576;
  assign n11578 = n11573 & ~n11574;
  assign n11579 = ~n11577 & n11578;
  assign n11580 = n11573 & ~n11579;
  assign n11581 = ~n11574 & ~n11579;
  assign n11582 = ~n11577 & n11581;
  assign n11583 = ~n11580 & ~n11582;
  assign n11584 = ~n11572 & ~n11583;
  assign n11585 = ~n11572 & ~n11584;
  assign n11586 = ~n11583 & ~n11584;
  assign n11587 = ~n11585 & ~n11586;
  assign n11588 = pi19  & pi55 ;
  assign n11589 = pi21  & pi53 ;
  assign n11590 = ~n11588 & ~n11589;
  assign n11591 = n3653 & n7172;
  assign n11592 = pi22  & pi52 ;
  assign n11593 = ~n11590 & n11592;
  assign n11594 = ~n11591 & n11593;
  assign n11595 = ~n11591 & ~n11594;
  assign n11596 = ~n11590 & n11595;
  assign n11597 = n11592 & ~n11594;
  assign n11598 = ~n11596 & ~n11597;
  assign n11599 = pi20  & pi54 ;
  assign n11600 = n3106 & n5548;
  assign n11601 = pi34  & pi40 ;
  assign n11602 = pi35  & pi39 ;
  assign n11603 = ~n11601 & ~n11602;
  assign n11604 = n11599 & ~n11600;
  assign n11605 = ~n11603 & n11604;
  assign n11606 = n11599 & ~n11605;
  assign n11607 = ~n11600 & ~n11605;
  assign n11608 = ~n11603 & n11607;
  assign n11609 = ~n11606 & ~n11608;
  assign n11610 = ~n11598 & ~n11609;
  assign n11611 = ~n11598 & ~n11610;
  assign n11612 = ~n11609 & ~n11610;
  assign n11613 = ~n11611 & ~n11612;
  assign n11614 = n2110 & n6114;
  assign n11615 = pi23  & pi51 ;
  assign n11616 = pi24  & pi50 ;
  assign n11617 = ~n11615 & ~n11616;
  assign n11618 = n3301 & ~n11614;
  assign n11619 = ~n11617 & n11618;
  assign n11620 = n3301 & ~n11619;
  assign n11621 = ~n11614 & ~n11619;
  assign n11622 = ~n11617 & n11621;
  assign n11623 = ~n11620 & ~n11622;
  assign n11624 = ~n11613 & ~n11623;
  assign n11625 = ~n11613 & ~n11624;
  assign n11626 = ~n11623 & ~n11624;
  assign n11627 = ~n11625 & ~n11626;
  assign n11628 = ~n11587 & n11627;
  assign n11629 = n11587 & ~n11627;
  assign n11630 = ~n11628 & ~n11629;
  assign n11631 = n11546 & ~n11630;
  assign n11632 = n11546 & ~n11631;
  assign n11633 = ~n11630 & ~n11631;
  assign n11634 = ~n11632 & ~n11633;
  assign n11635 = n11518 & ~n11634;
  assign n11636 = n11518 & ~n11635;
  assign n11637 = ~n11634 & ~n11635;
  assign n11638 = ~n11636 & ~n11637;
  assign n11639 = ~n11495 & n11638;
  assign n11640 = n11495 & ~n11638;
  assign n11641 = ~n11639 & ~n11640;
  assign n11642 = ~n11301 & ~n11442;
  assign n11643 = ~n11434 & ~n11438;
  assign n11644 = ~n11275 & ~n11297;
  assign n11645 = ~n11286 & ~n11289;
  assign n11646 = ~n11279 & ~n11283;
  assign n11647 = n11645 & n11646;
  assign n11648 = ~n11645 & ~n11646;
  assign n11649 = ~n11647 & ~n11648;
  assign n11650 = ~n11366 & ~n11369;
  assign n11651 = ~n11649 & n11650;
  assign n11652 = n11649 & ~n11650;
  assign n11653 = ~n11651 & ~n11652;
  assign n11654 = ~n11291 & ~n11294;
  assign n11655 = ~n11267 & ~n11271;
  assign n11656 = n11654 & n11655;
  assign n11657 = ~n11654 & ~n11655;
  assign n11658 = ~n11656 & ~n11657;
  assign n11659 = n11653 & n11658;
  assign n11660 = ~n11653 & ~n11658;
  assign n11661 = ~n11659 & ~n11660;
  assign n11662 = ~n11644 & n11661;
  assign n11663 = n11644 & ~n11661;
  assign n11664 = ~n11662 & ~n11663;
  assign n11665 = ~n11643 & n11664;
  assign n11666 = n11643 & ~n11664;
  assign n11667 = ~n11665 & ~n11666;
  assign n11668 = ~n11642 & n11667;
  assign n11669 = n11642 & ~n11667;
  assign n11670 = ~n11668 & ~n11669;
  assign n11671 = ~n11641 & n11670;
  assign n11672 = n11641 & ~n11670;
  assign n11673 = ~n11671 & ~n11672;
  assign n11674 = n11455 & ~n11673;
  assign n11675 = ~n11455 & n11673;
  assign n11676 = ~n11674 & ~n11675;
  assign n11677 = ~n11221 & ~n11449;
  assign n11678 = ~n11450 & ~n11677;
  assign n11679 = ~n11676 & n11678;
  assign n11680 = n11676 & ~n11678;
  assign po75  = ~n11679 & ~n11680;
  assign n11682 = ~n11668 & ~n11671;
  assign n11683 = ~n11662 & ~n11665;
  assign n11684 = ~n11458 & ~n11471;
  assign n11685 = ~n11504 & ~n11507;
  assign n11686 = n11684 & n11685;
  assign n11687 = ~n11684 & ~n11685;
  assign n11688 = ~n11686 & ~n11687;
  assign n11689 = ~n11498 & ~n11501;
  assign n11690 = ~n11688 & n11689;
  assign n11691 = n11688 & ~n11689;
  assign n11692 = ~n11690 & ~n11691;
  assign n11693 = ~n11587 & ~n11627;
  assign n11694 = ~n11631 & ~n11693;
  assign n11695 = n11692 & ~n11694;
  assign n11696 = ~n11692 & n11694;
  assign n11697 = ~n11695 & ~n11696;
  assign n11698 = ~n11539 & ~n11545;
  assign n11699 = n11607 & n11621;
  assign n11700 = ~n11607 & ~n11621;
  assign n11701 = ~n11699 & ~n11700;
  assign n11702 = n11595 & ~n11701;
  assign n11703 = ~n11595 & n11701;
  assign n11704 = ~n11702 & ~n11703;
  assign n11705 = n11554 & n11566;
  assign n11706 = ~n11554 & ~n11566;
  assign n11707 = ~n11705 & ~n11706;
  assign n11708 = ~n11519 & ~n11525;
  assign n11709 = ~n11707 & n11708;
  assign n11710 = n11707 & ~n11708;
  assign n11711 = ~n11709 & ~n11710;
  assign n11712 = n11704 & n11711;
  assign n11713 = ~n11704 & ~n11711;
  assign n11714 = ~n11712 & ~n11713;
  assign n11715 = ~n11698 & n11714;
  assign n11716 = n11698 & ~n11714;
  assign n11717 = ~n11715 & ~n11716;
  assign n11718 = n11697 & n11717;
  assign n11719 = ~n11697 & ~n11717;
  assign n11720 = ~n11718 & ~n11719;
  assign n11721 = n11683 & ~n11720;
  assign n11722 = ~n11683 & n11720;
  assign n11723 = ~n11721 & ~n11722;
  assign n11724 = ~n11657 & ~n11659;
  assign n11725 = n11536 & n11581;
  assign n11726 = ~n11536 & ~n11581;
  assign n11727 = ~n11725 & ~n11726;
  assign n11728 = n11468 & ~n11727;
  assign n11729 = ~n11468 & n11727;
  assign n11730 = ~n11728 & ~n11729;
  assign n11731 = ~n11610 & ~n11624;
  assign n11732 = ~n11569 & ~n11584;
  assign n11733 = n11731 & n11732;
  assign n11734 = ~n11731 & ~n11732;
  assign n11735 = ~n11733 & ~n11734;
  assign n11736 = n11730 & n11735;
  assign n11737 = ~n11730 & ~n11735;
  assign n11738 = ~n11736 & ~n11737;
  assign n11739 = ~n11724 & n11738;
  assign n11740 = n11724 & ~n11738;
  assign n11741 = ~n11739 & ~n11740;
  assign n11742 = pi12  & pi63 ;
  assign n11743 = pi19  & pi56 ;
  assign n11744 = ~n11742 & ~n11743;
  assign n11745 = pi19  & pi63 ;
  assign n11746 = n10157 & n11745;
  assign n11747 = pi30  & pi45 ;
  assign n11748 = ~n11744 & n11747;
  assign n11749 = ~n11746 & n11748;
  assign n11750 = ~n11746 & ~n11749;
  assign n11751 = ~n11744 & n11750;
  assign n11752 = n11747 & ~n11749;
  assign n11753 = ~n11751 & ~n11752;
  assign n11754 = pi23  & pi52 ;
  assign n11755 = n4691 & n5548;
  assign n11756 = pi36  & pi39 ;
  assign n11757 = pi35  & pi40 ;
  assign n11758 = ~n11756 & ~n11757;
  assign n11759 = n11754 & ~n11755;
  assign n11760 = ~n11758 & n11759;
  assign n11761 = n11754 & ~n11760;
  assign n11762 = ~n11755 & ~n11760;
  assign n11763 = ~n11758 & n11762;
  assign n11764 = ~n11761 & ~n11763;
  assign n11765 = ~n11753 & ~n11764;
  assign n11766 = ~n11753 & ~n11765;
  assign n11767 = ~n11764 & ~n11765;
  assign n11768 = ~n11766 & ~n11767;
  assign n11769 = pi38  & pi62 ;
  assign n11770 = pi13  & n11769;
  assign n11771 = n5055 & ~n11770;
  assign n11772 = n5055 & ~n11771;
  assign n11773 = ~n11770 & ~n11771;
  assign n11774 = pi13  & pi62 ;
  assign n11775 = ~pi38  & ~n11774;
  assign n11776 = n11773 & ~n11775;
  assign n11777 = ~n11772 & ~n11776;
  assign n11778 = ~n11768 & ~n11777;
  assign n11779 = ~n11768 & ~n11778;
  assign n11780 = ~n11777 & ~n11778;
  assign n11781 = ~n11779 & ~n11780;
  assign n11782 = ~n11648 & ~n11652;
  assign n11783 = n11781 & n11782;
  assign n11784 = ~n11781 & ~n11782;
  assign n11785 = ~n11783 & ~n11784;
  assign n11786 = pi15  & pi60 ;
  assign n11787 = pi16  & pi59 ;
  assign n11788 = ~n11786 & ~n11787;
  assign n11789 = n840 & n8854;
  assign n11790 = pi14  & pi61 ;
  assign n11791 = ~n11788 & n11790;
  assign n11792 = ~n11789 & n11791;
  assign n11793 = ~n11789 & ~n11792;
  assign n11794 = ~n11788 & n11793;
  assign n11795 = n11790 & ~n11792;
  assign n11796 = ~n11794 & ~n11795;
  assign n11797 = pi17  & pi58 ;
  assign n11798 = pi49  & pi57 ;
  assign n11799 = n4242 & n11798;
  assign n11800 = pi18  & pi57 ;
  assign n11801 = pi26  & pi49 ;
  assign n11802 = ~n11800 & ~n11801;
  assign n11803 = n11797 & ~n11799;
  assign n11804 = ~n11802 & n11803;
  assign n11805 = n11797 & ~n11804;
  assign n11806 = ~n11799 & ~n11804;
  assign n11807 = ~n11802 & n11806;
  assign n11808 = ~n11805 & ~n11807;
  assign n11809 = ~n11796 & ~n11808;
  assign n11810 = ~n11796 & ~n11809;
  assign n11811 = ~n11808 & ~n11809;
  assign n11812 = ~n11810 & ~n11811;
  assign n11813 = pi27  & pi48 ;
  assign n11814 = n2915 & n5277;
  assign n11815 = pi28  & pi47 ;
  assign n11816 = pi29  & pi46 ;
  assign n11817 = ~n11815 & ~n11816;
  assign n11818 = n11813 & ~n11814;
  assign n11819 = ~n11817 & n11818;
  assign n11820 = n11813 & ~n11819;
  assign n11821 = ~n11814 & ~n11819;
  assign n11822 = ~n11817 & n11821;
  assign n11823 = ~n11820 & ~n11822;
  assign n11824 = ~n11812 & ~n11823;
  assign n11825 = ~n11812 & ~n11824;
  assign n11826 = ~n11823 & ~n11824;
  assign n11827 = ~n11825 & ~n11826;
  assign n11828 = n11785 & ~n11827;
  assign n11829 = ~n11785 & n11827;
  assign n11830 = ~n11828 & ~n11829;
  assign n11831 = n11741 & n11830;
  assign n11832 = n11741 & ~n11831;
  assign n11833 = n11830 & ~n11831;
  assign n11834 = ~n11832 & ~n11833;
  assign n11835 = ~n11723 & n11834;
  assign n11836 = n11723 & ~n11834;
  assign n11837 = ~n11835 & ~n11836;
  assign n11838 = ~n11477 & ~n11481;
  assign n11839 = pi20  & pi55 ;
  assign n11840 = pi25  & pi50 ;
  assign n11841 = ~n11839 & ~n11840;
  assign n11842 = n11839 & n11840;
  assign n11843 = pi34  & pi41 ;
  assign n11844 = ~n11841 & n11843;
  assign n11845 = ~n11842 & n11844;
  assign n11846 = ~n11842 & ~n11845;
  assign n11847 = ~n11841 & n11846;
  assign n11848 = n11843 & ~n11845;
  assign n11849 = ~n11847 & ~n11848;
  assign n11850 = pi31  & pi44 ;
  assign n11851 = n6138 & n6458;
  assign n11852 = pi33  & pi42 ;
  assign n11853 = ~n4941 & ~n11852;
  assign n11854 = n11850 & ~n11851;
  assign n11855 = ~n11853 & n11854;
  assign n11856 = n11850 & ~n11855;
  assign n11857 = ~n11851 & ~n11855;
  assign n11858 = ~n11853 & n11857;
  assign n11859 = ~n11856 & ~n11858;
  assign n11860 = ~n11849 & ~n11859;
  assign n11861 = ~n11849 & ~n11860;
  assign n11862 = ~n11859 & ~n11860;
  assign n11863 = ~n11861 & ~n11862;
  assign n11864 = pi21  & pi54 ;
  assign n11865 = n1990 & n6765;
  assign n11866 = pi22  & pi53 ;
  assign n11867 = pi24  & pi51 ;
  assign n11868 = ~n11866 & ~n11867;
  assign n11869 = n11864 & ~n11865;
  assign n11870 = ~n11868 & n11869;
  assign n11871 = n11864 & ~n11870;
  assign n11872 = ~n11865 & ~n11870;
  assign n11873 = ~n11868 & n11872;
  assign n11874 = ~n11871 & ~n11873;
  assign n11875 = ~n11863 & ~n11874;
  assign n11876 = ~n11863 & ~n11875;
  assign n11877 = ~n11874 & ~n11875;
  assign n11878 = ~n11876 & ~n11877;
  assign n11879 = ~n11511 & ~n11513;
  assign n11880 = ~n11878 & ~n11879;
  assign n11881 = ~n11878 & ~n11880;
  assign n11882 = ~n11879 & ~n11880;
  assign n11883 = ~n11881 & ~n11882;
  assign n11884 = ~n11838 & ~n11883;
  assign n11885 = ~n11838 & ~n11884;
  assign n11886 = ~n11883 & ~n11884;
  assign n11887 = ~n11885 & ~n11886;
  assign n11888 = ~n11485 & ~n11489;
  assign n11889 = ~n11887 & ~n11888;
  assign n11890 = ~n11887 & ~n11889;
  assign n11891 = ~n11888 & ~n11889;
  assign n11892 = ~n11890 & ~n11891;
  assign n11893 = ~n11516 & ~n11635;
  assign n11894 = n11892 & n11893;
  assign n11895 = ~n11892 & ~n11893;
  assign n11896 = ~n11894 & ~n11895;
  assign n11897 = ~n11495 & ~n11638;
  assign n11898 = ~n11492 & ~n11897;
  assign n11899 = n11896 & ~n11898;
  assign n11900 = ~n11896 & n11898;
  assign n11901 = ~n11899 & ~n11900;
  assign n11902 = n11837 & n11901;
  assign n11903 = ~n11837 & ~n11901;
  assign n11904 = ~n11902 & ~n11903;
  assign n11905 = ~n11682 & n11904;
  assign n11906 = n11682 & ~n11904;
  assign n11907 = ~n11905 & ~n11906;
  assign n11908 = ~n11675 & ~n11680;
  assign n11909 = ~n11907 & n11908;
  assign n11910 = n11907 & ~n11908;
  assign po76  = ~n11909 & ~n11910;
  assign n11912 = ~n11899 & ~n11902;
  assign n11913 = ~n11722 & ~n11836;
  assign n11914 = ~n11739 & ~n11831;
  assign n11915 = ~n11695 & ~n11718;
  assign n11916 = ~n11712 & ~n11715;
  assign n11917 = pi31  & pi45 ;
  assign n11918 = pi32  & pi44 ;
  assign n11919 = ~n11917 & ~n11918;
  assign n11920 = n3567 & n5318;
  assign n11921 = pi13  & pi63 ;
  assign n11922 = ~n11919 & n11921;
  assign n11923 = ~n11920 & n11922;
  assign n11924 = ~n11920 & ~n11923;
  assign n11925 = ~n11919 & n11924;
  assign n11926 = n11921 & ~n11923;
  assign n11927 = ~n11925 & ~n11926;
  assign n11928 = pi19  & pi57 ;
  assign n11929 = pi23  & pi53 ;
  assign n11930 = n11928 & n11929;
  assign n11931 = ~n11928 & ~n11929;
  assign n11932 = n5076 & ~n11930;
  assign n11933 = ~n11931 & n11932;
  assign n11934 = n5076 & ~n11933;
  assign n11935 = ~n11930 & ~n11933;
  assign n11936 = ~n11931 & n11935;
  assign n11937 = ~n11934 & ~n11936;
  assign n11938 = ~n11927 & ~n11937;
  assign n11939 = ~n11927 & ~n11938;
  assign n11940 = ~n11937 & ~n11938;
  assign n11941 = ~n11939 & ~n11940;
  assign n11942 = n1481 & n9891;
  assign n11943 = pi21  & pi55 ;
  assign n11944 = pi22  & pi54 ;
  assign n11945 = ~n11943 & ~n11944;
  assign n11946 = n9781 & ~n11942;
  assign n11947 = ~n11945 & n11946;
  assign n11948 = n9781 & ~n11947;
  assign n11949 = ~n11942 & ~n11947;
  assign n11950 = ~n11945 & n11949;
  assign n11951 = ~n11948 & ~n11950;
  assign n11952 = ~n11941 & ~n11951;
  assign n11953 = ~n11941 & ~n11952;
  assign n11954 = ~n11951 & ~n11952;
  assign n11955 = ~n11953 & ~n11954;
  assign n11956 = ~n11734 & ~n11736;
  assign n11957 = ~n11955 & ~n11956;
  assign n11958 = n11955 & n11956;
  assign n11959 = ~n11957 & ~n11958;
  assign n11960 = ~n11916 & n11959;
  assign n11961 = n11916 & ~n11959;
  assign n11962 = ~n11960 & ~n11961;
  assign n11963 = ~n11915 & n11962;
  assign n11964 = n11915 & ~n11962;
  assign n11965 = ~n11963 & ~n11964;
  assign n11966 = ~n11914 & n11965;
  assign n11967 = n11914 & ~n11965;
  assign n11968 = ~n11966 & ~n11967;
  assign n11969 = ~n11913 & n11968;
  assign n11970 = n11913 & ~n11968;
  assign n11971 = ~n11969 & ~n11970;
  assign n11972 = ~n11706 & ~n11710;
  assign n11973 = ~n11726 & ~n11729;
  assign n11974 = n11972 & n11973;
  assign n11975 = ~n11972 & ~n11973;
  assign n11976 = ~n11974 & ~n11975;
  assign n11977 = ~n11700 & ~n11703;
  assign n11978 = ~n11976 & n11977;
  assign n11979 = n11976 & ~n11977;
  assign n11980 = ~n11978 & ~n11979;
  assign n11981 = ~n11784 & ~n11828;
  assign n11982 = n11980 & ~n11981;
  assign n11983 = ~n11980 & n11981;
  assign n11984 = ~n11982 & ~n11983;
  assign n11985 = n11821 & n11846;
  assign n11986 = ~n11821 & ~n11846;
  assign n11987 = ~n11985 & ~n11986;
  assign n11988 = n11750 & ~n11987;
  assign n11989 = ~n11750 & n11987;
  assign n11990 = ~n11988 & ~n11989;
  assign n11991 = ~n11860 & ~n11875;
  assign n11992 = pi14  & pi62 ;
  assign n11993 = n11773 & ~n11992;
  assign n11994 = ~n11773 & n11992;
  assign n11995 = ~n11762 & ~n11993;
  assign n11996 = ~n11994 & n11995;
  assign n11997 = ~n11994 & ~n11996;
  assign n11998 = ~n11993 & n11997;
  assign n11999 = ~n11762 & ~n11996;
  assign n12000 = ~n11998 & ~n11999;
  assign n12001 = ~n11991 & ~n12000;
  assign n12002 = ~n11991 & ~n12001;
  assign n12003 = ~n12000 & ~n12001;
  assign n12004 = ~n12002 & ~n12003;
  assign n12005 = n11990 & ~n12004;
  assign n12006 = n11990 & ~n12005;
  assign n12007 = ~n12004 & ~n12005;
  assign n12008 = ~n12006 & ~n12007;
  assign n12009 = n11984 & ~n12008;
  assign n12010 = n11984 & ~n12009;
  assign n12011 = ~n12008 & ~n12009;
  assign n12012 = ~n12010 & ~n12011;
  assign n12013 = ~n11889 & ~n11895;
  assign n12014 = n12012 & n12013;
  assign n12015 = ~n12012 & ~n12013;
  assign n12016 = ~n12014 & ~n12015;
  assign n12017 = ~n11880 & ~n11884;
  assign n12018 = n11793 & n11806;
  assign n12019 = ~n11793 & ~n11806;
  assign n12020 = ~n12018 & ~n12019;
  assign n12021 = n11857 & ~n12020;
  assign n12022 = ~n11857 & n12020;
  assign n12023 = ~n12021 & ~n12022;
  assign n12024 = ~n11809 & ~n11824;
  assign n12025 = ~n11765 & ~n11778;
  assign n12026 = n12024 & n12025;
  assign n12027 = ~n12024 & ~n12025;
  assign n12028 = ~n12026 & ~n12027;
  assign n12029 = n12023 & n12028;
  assign n12030 = ~n12023 & ~n12028;
  assign n12031 = ~n12029 & ~n12030;
  assign n12032 = n12017 & ~n12031;
  assign n12033 = ~n12017 & n12031;
  assign n12034 = ~n12032 & ~n12033;
  assign n12035 = pi29  & pi47 ;
  assign n12036 = pi30  & pi46 ;
  assign n12037 = ~n12035 & ~n12036;
  assign n12038 = n4908 & n5277;
  assign n12039 = pi28  & pi48 ;
  assign n12040 = ~n12037 & n12039;
  assign n12041 = ~n12038 & n12040;
  assign n12042 = ~n12038 & ~n12041;
  assign n12043 = ~n12037 & n12042;
  assign n12044 = n12039 & ~n12041;
  assign n12045 = ~n12043 & ~n12044;
  assign n12046 = pi34  & pi42 ;
  assign n12047 = n4691 & n6012;
  assign n12048 = pi35  & pi41 ;
  assign n12049 = pi36  & pi40 ;
  assign n12050 = ~n12048 & ~n12049;
  assign n12051 = n12046 & ~n12047;
  assign n12052 = ~n12050 & n12051;
  assign n12053 = n12046 & ~n12052;
  assign n12054 = ~n12047 & ~n12052;
  assign n12055 = ~n12050 & n12054;
  assign n12056 = ~n12053 & ~n12055;
  assign n12057 = ~n12045 & ~n12056;
  assign n12058 = ~n12045 & ~n12057;
  assign n12059 = ~n12056 & ~n12057;
  assign n12060 = ~n12058 & ~n12059;
  assign n12061 = n1789 & n10319;
  assign n12062 = pi24  & pi52 ;
  assign n12063 = pi25  & pi51 ;
  assign n12064 = ~n12062 & ~n12063;
  assign n12065 = n5302 & ~n12061;
  assign n12066 = ~n12064 & n12065;
  assign n12067 = n5302 & ~n12066;
  assign n12068 = ~n12061 & ~n12066;
  assign n12069 = ~n12064 & n12068;
  assign n12070 = ~n12067 & ~n12069;
  assign n12071 = ~n12060 & ~n12070;
  assign n12072 = ~n12060 & ~n12071;
  assign n12073 = ~n12070 & ~n12071;
  assign n12074 = ~n12072 & ~n12073;
  assign n12075 = ~n11687 & ~n11691;
  assign n12076 = n12074 & n12075;
  assign n12077 = ~n12074 & ~n12075;
  assign n12078 = ~n12076 & ~n12077;
  assign n12079 = pi15  & pi61 ;
  assign n12080 = n989 & n8854;
  assign n12081 = pi16  & pi60 ;
  assign n12082 = pi17  & pi59 ;
  assign n12083 = ~n12081 & ~n12082;
  assign n12084 = n12079 & ~n12080;
  assign n12085 = ~n12083 & n12084;
  assign n12086 = n12079 & ~n12085;
  assign n12087 = ~n12080 & ~n12085;
  assign n12088 = ~n12083 & n12087;
  assign n12089 = ~n12086 & ~n12088;
  assign n12090 = n11872 & ~n12089;
  assign n12091 = ~n11872 & n12089;
  assign n12092 = ~n12090 & ~n12091;
  assign n12093 = pi18  & pi58 ;
  assign n12094 = n2646 & n5889;
  assign n12095 = pi26  & pi50 ;
  assign n12096 = pi27  & pi49 ;
  assign n12097 = ~n12095 & ~n12096;
  assign n12098 = n12093 & ~n12094;
  assign n12099 = ~n12097 & n12098;
  assign n12100 = n12093 & ~n12099;
  assign n12101 = ~n12094 & ~n12099;
  assign n12102 = ~n12097 & n12101;
  assign n12103 = ~n12100 & ~n12102;
  assign n12104 = ~n12092 & ~n12103;
  assign n12105 = n12092 & n12103;
  assign n12106 = ~n12104 & ~n12105;
  assign n12107 = n12078 & n12106;
  assign n12108 = ~n12078 & ~n12106;
  assign n12109 = ~n12107 & ~n12108;
  assign n12110 = n12034 & n12109;
  assign n12111 = n12034 & ~n12110;
  assign n12112 = n12109 & ~n12110;
  assign n12113 = ~n12111 & ~n12112;
  assign n12114 = n12016 & ~n12113;
  assign n12115 = ~n12016 & n12113;
  assign n12116 = ~n12114 & ~n12115;
  assign n12117 = n11971 & n12116;
  assign n12118 = n11971 & ~n12117;
  assign n12119 = n12116 & ~n12117;
  assign n12120 = ~n12118 & ~n12119;
  assign n12121 = ~n11912 & ~n12120;
  assign n12122 = n11912 & n12120;
  assign n12123 = ~n12121 & ~n12122;
  assign n12124 = ~n11905 & ~n11910;
  assign n12125 = n12123 & ~n12124;
  assign n12126 = ~n12123 & n12124;
  assign po77  = ~n12125 & ~n12126;
  assign n12128 = ~n11969 & ~n12117;
  assign n12129 = ~n12015 & ~n12114;
  assign n12130 = ~n12033 & ~n12110;
  assign n12131 = ~n11982 & ~n12009;
  assign n12132 = ~n12001 & ~n12005;
  assign n12133 = pi22  & pi55 ;
  assign n12134 = pi26  & pi51 ;
  assign n12135 = ~n12133 & ~n12134;
  assign n12136 = n12133 & n12134;
  assign n12137 = pi34  & pi43 ;
  assign n12138 = ~n12135 & n12137;
  assign n12139 = ~n12136 & n12138;
  assign n12140 = ~n12136 & ~n12139;
  assign n12141 = ~n12135 & n12140;
  assign n12142 = n12137 & ~n12139;
  assign n12143 = ~n12141 & ~n12142;
  assign n12144 = pi25  & pi52 ;
  assign n12145 = n2110 & n8092;
  assign n12146 = pi23  & pi54 ;
  assign n12147 = pi24  & pi53 ;
  assign n12148 = ~n12146 & ~n12147;
  assign n12149 = n12144 & ~n12145;
  assign n12150 = ~n12148 & n12149;
  assign n12151 = n12144 & ~n12150;
  assign n12152 = ~n12145 & ~n12150;
  assign n12153 = ~n12148 & n12152;
  assign n12154 = ~n12151 & ~n12153;
  assign n12155 = ~n12143 & ~n12154;
  assign n12156 = ~n12143 & ~n12155;
  assign n12157 = ~n12154 & ~n12155;
  assign n12158 = ~n12156 & ~n12157;
  assign n12159 = pi16  & pi61 ;
  assign n12160 = n5318 & n6138;
  assign n12161 = pi33  & pi44 ;
  assign n12162 = pi32  & pi45 ;
  assign n12163 = ~n12161 & ~n12162;
  assign n12164 = n12159 & ~n12160;
  assign n12165 = ~n12163 & n12164;
  assign n12166 = n12159 & ~n12165;
  assign n12167 = ~n12160 & ~n12165;
  assign n12168 = ~n12163 & n12167;
  assign n12169 = ~n12166 & ~n12168;
  assign n12170 = ~n12158 & ~n12169;
  assign n12171 = ~n12158 & ~n12170;
  assign n12172 = ~n12169 & ~n12170;
  assign n12173 = ~n12171 & ~n12172;
  assign n12174 = ~n12027 & ~n12029;
  assign n12175 = ~n12173 & ~n12174;
  assign n12176 = ~n12173 & ~n12175;
  assign n12177 = ~n12174 & ~n12175;
  assign n12178 = ~n12176 & ~n12177;
  assign n12179 = ~n12132 & ~n12178;
  assign n12180 = n12132 & n12178;
  assign n12181 = ~n12179 & ~n12180;
  assign n12182 = ~n12131 & n12181;
  assign n12183 = n12131 & ~n12181;
  assign n12184 = ~n12182 & ~n12183;
  assign n12185 = ~n12130 & n12184;
  assign n12186 = n12130 & ~n12184;
  assign n12187 = ~n12185 & ~n12186;
  assign n12188 = ~n12129 & n12187;
  assign n12189 = n12129 & ~n12187;
  assign n12190 = ~n12188 & ~n12189;
  assign n12191 = ~n11963 & ~n11966;
  assign n12192 = n1199 & n8854;
  assign n12193 = pi18  & pi59 ;
  assign n12194 = ~n12192 & n12193;
  assign n12195 = pi17  & pi60 ;
  assign n12196 = ~n12192 & n12195;
  assign n12197 = ~n12194 & ~n12196;
  assign n12198 = ~n12068 & ~n12197;
  assign n12199 = ~n12068 & ~n12198;
  assign n12200 = ~n12197 & ~n12198;
  assign n12201 = ~n12199 & ~n12200;
  assign n12202 = ~n12019 & ~n12022;
  assign n12203 = n12201 & n12202;
  assign n12204 = ~n12201 & ~n12202;
  assign n12205 = ~n12203 & ~n12204;
  assign n12206 = ~n11986 & ~n11989;
  assign n12207 = ~n12205 & n12206;
  assign n12208 = n12205 & ~n12206;
  assign n12209 = ~n12207 & ~n12208;
  assign n12210 = ~n12077 & ~n12107;
  assign n12211 = n12209 & ~n12210;
  assign n12212 = ~n12209 & n12210;
  assign n12213 = ~n12211 & ~n12212;
  assign n12214 = n11949 & n12042;
  assign n12215 = ~n11949 & ~n12042;
  assign n12216 = ~n12214 & ~n12215;
  assign n12217 = n11924 & ~n12216;
  assign n12218 = ~n11924 & n12216;
  assign n12219 = ~n12217 & ~n12218;
  assign n12220 = n12087 & n12101;
  assign n12221 = ~n12087 & ~n12101;
  assign n12222 = ~n12220 & ~n12221;
  assign n12223 = n11935 & ~n12222;
  assign n12224 = ~n11935 & n12222;
  assign n12225 = ~n12223 & ~n12224;
  assign n12226 = ~n11938 & ~n11952;
  assign n12227 = ~n12225 & n12226;
  assign n12228 = n12225 & ~n12226;
  assign n12229 = ~n12227 & ~n12228;
  assign n12230 = n12219 & n12229;
  assign n12231 = ~n12219 & ~n12229;
  assign n12232 = ~n12230 & ~n12231;
  assign n12233 = n12213 & n12232;
  assign n12234 = ~n12213 & ~n12232;
  assign n12235 = ~n12233 & ~n12234;
  assign n12236 = n12191 & ~n12235;
  assign n12237 = ~n12191 & n12235;
  assign n12238 = ~n12236 & ~n12237;
  assign n12239 = ~n11872 & ~n12089;
  assign n12240 = ~n12104 & ~n12239;
  assign n12241 = n11997 & n12240;
  assign n12242 = ~n11997 & ~n12240;
  assign n12243 = ~n12241 & ~n12242;
  assign n12244 = ~n12057 & ~n12071;
  assign n12245 = ~n12243 & n12244;
  assign n12246 = n12243 & ~n12244;
  assign n12247 = ~n12245 & ~n12246;
  assign n12248 = ~n11957 & ~n11960;
  assign n12249 = ~n12247 & n12248;
  assign n12250 = n12247 & ~n12248;
  assign n12251 = ~n12249 & ~n12250;
  assign n12252 = pi14  & pi63 ;
  assign n12253 = pi31  & pi46 ;
  assign n12254 = ~n12252 & ~n12253;
  assign n12255 = pi31  & pi63 ;
  assign n12256 = n6893 & n12255;
  assign n12257 = pi30  & pi47 ;
  assign n12258 = ~n12254 & n12257;
  assign n12259 = ~n12256 & n12258;
  assign n12260 = ~n12256 & ~n12259;
  assign n12261 = ~n12254 & n12260;
  assign n12262 = n12257 & ~n12259;
  assign n12263 = ~n12261 & ~n12262;
  assign n12264 = pi35  & pi42 ;
  assign n12265 = n4500 & n6012;
  assign n12266 = pi37  & pi40 ;
  assign n12267 = pi36  & pi41 ;
  assign n12268 = ~n12266 & ~n12267;
  assign n12269 = n12264 & ~n12265;
  assign n12270 = ~n12268 & n12269;
  assign n12271 = n12264 & ~n12270;
  assign n12272 = ~n12265 & ~n12270;
  assign n12273 = ~n12268 & n12272;
  assign n12274 = ~n12271 & ~n12273;
  assign n12275 = ~n12263 & ~n12274;
  assign n12276 = ~n12263 & ~n12275;
  assign n12277 = ~n12274 & ~n12275;
  assign n12278 = ~n12276 & ~n12277;
  assign n12279 = pi62  & n6505;
  assign n12280 = n4736 & ~n12279;
  assign n12281 = n4736 & ~n12280;
  assign n12282 = ~n12279 & ~n12280;
  assign n12283 = pi15  & pi62 ;
  assign n12284 = ~pi39  & ~n12283;
  assign n12285 = n12282 & ~n12284;
  assign n12286 = ~n12281 & ~n12285;
  assign n12287 = ~n12278 & ~n12286;
  assign n12288 = ~n12278 & ~n12287;
  assign n12289 = ~n12286 & ~n12287;
  assign n12290 = ~n12288 & ~n12289;
  assign n12291 = ~n11975 & ~n11979;
  assign n12292 = n12290 & n12291;
  assign n12293 = ~n12290 & ~n12291;
  assign n12294 = ~n12292 & ~n12293;
  assign n12295 = pi19  & pi58 ;
  assign n12296 = n1593 & n7643;
  assign n12297 = pi20  & pi57 ;
  assign n12298 = pi21  & pi56 ;
  assign n12299 = ~n12297 & ~n12298;
  assign n12300 = n12295 & ~n12296;
  assign n12301 = ~n12299 & n12300;
  assign n12302 = n12295 & ~n12301;
  assign n12303 = ~n12296 & ~n12301;
  assign n12304 = ~n12299 & n12303;
  assign n12305 = ~n12302 & ~n12304;
  assign n12306 = n12054 & ~n12305;
  assign n12307 = ~n12054 & n12305;
  assign n12308 = ~n12306 & ~n12307;
  assign n12309 = pi27  & pi50 ;
  assign n12310 = n2915 & n8505;
  assign n12311 = pi28  & pi49 ;
  assign n12312 = pi29  & pi48 ;
  assign n12313 = ~n12311 & ~n12312;
  assign n12314 = n12309 & ~n12310;
  assign n12315 = ~n12313 & n12314;
  assign n12316 = n12309 & ~n12315;
  assign n12317 = ~n12310 & ~n12315;
  assign n12318 = ~n12313 & n12317;
  assign n12319 = ~n12316 & ~n12318;
  assign n12320 = ~n12308 & ~n12319;
  assign n12321 = n12308 & n12319;
  assign n12322 = ~n12320 & ~n12321;
  assign n12323 = n12294 & n12322;
  assign n12324 = ~n12294 & ~n12322;
  assign n12325 = ~n12323 & ~n12324;
  assign n12326 = n12251 & n12325;
  assign n12327 = n12251 & ~n12326;
  assign n12328 = n12325 & ~n12326;
  assign n12329 = ~n12327 & ~n12328;
  assign n12330 = n12238 & ~n12329;
  assign n12331 = ~n12238 & n12329;
  assign n12332 = ~n12330 & ~n12331;
  assign n12333 = n12190 & n12332;
  assign n12334 = n12190 & ~n12333;
  assign n12335 = n12332 & ~n12333;
  assign n12336 = ~n12334 & ~n12335;
  assign n12337 = ~n12128 & ~n12336;
  assign n12338 = n12128 & n12336;
  assign n12339 = ~n12337 & ~n12338;
  assign n12340 = ~n12121 & ~n12125;
  assign n12341 = ~n12339 & n12340;
  assign n12342 = n12339 & ~n12340;
  assign po78  = ~n12341 & ~n12342;
  assign n12344 = ~n12188 & ~n12333;
  assign n12345 = ~n12250 & ~n12326;
  assign n12346 = ~n12211 & ~n12233;
  assign n12347 = ~n12242 & ~n12246;
  assign n12348 = pi19  & pi59 ;
  assign n12349 = pi21  & pi57 ;
  assign n12350 = ~n12348 & ~n12349;
  assign n12351 = pi57  & pi59 ;
  assign n12352 = n3653 & n12351;
  assign n12353 = pi18  & pi60 ;
  assign n12354 = ~n12350 & n12353;
  assign n12355 = ~n12352 & n12354;
  assign n12356 = ~n12352 & ~n12355;
  assign n12357 = ~n12350 & n12356;
  assign n12358 = n12353 & ~n12355;
  assign n12359 = ~n12357 & ~n12358;
  assign n12360 = pi27  & pi51 ;
  assign n12361 = n2915 & n5889;
  assign n12362 = pi28  & pi50 ;
  assign n12363 = pi29  & pi49 ;
  assign n12364 = ~n12362 & ~n12363;
  assign n12365 = n12360 & ~n12361;
  assign n12366 = ~n12364 & n12365;
  assign n12367 = n12360 & ~n12366;
  assign n12368 = ~n12361 & ~n12366;
  assign n12369 = ~n12364 & n12368;
  assign n12370 = ~n12367 & ~n12369;
  assign n12371 = ~n12359 & ~n12370;
  assign n12372 = ~n12359 & ~n12371;
  assign n12373 = ~n12370 & ~n12371;
  assign n12374 = ~n12372 & ~n12373;
  assign n12375 = pi15  & pi63 ;
  assign n12376 = n989 & n9567;
  assign n12377 = pi16  & pi62 ;
  assign n12378 = pi17  & pi61 ;
  assign n12379 = ~n12377 & ~n12378;
  assign n12380 = n12375 & ~n12376;
  assign n12381 = ~n12379 & n12380;
  assign n12382 = n12375 & ~n12381;
  assign n12383 = ~n12376 & ~n12381;
  assign n12384 = ~n12379 & n12383;
  assign n12385 = ~n12382 & ~n12384;
  assign n12386 = ~n12374 & ~n12385;
  assign n12387 = ~n12374 & ~n12386;
  assign n12388 = ~n12385 & ~n12386;
  assign n12389 = ~n12387 & ~n12388;
  assign n12390 = pi30  & pi48 ;
  assign n12391 = pi31  & pi47 ;
  assign n12392 = ~n12390 & ~n12391;
  assign n12393 = n2680 & n5823;
  assign n12394 = pi20  & pi58 ;
  assign n12395 = ~n12392 & n12394;
  assign n12396 = ~n12393 & n12395;
  assign n12397 = ~n12393 & ~n12396;
  assign n12398 = ~n12392 & n12397;
  assign n12399 = n12394 & ~n12396;
  assign n12400 = ~n12398 & ~n12399;
  assign n12401 = pi33  & pi45 ;
  assign n12402 = pi34  & pi44 ;
  assign n12403 = ~n12401 & ~n12402;
  assign n12404 = n3900 & n5318;
  assign n12405 = pi32  & pi46 ;
  assign n12406 = ~n12403 & n12405;
  assign n12407 = ~n12404 & n12406;
  assign n12408 = ~n12404 & ~n12407;
  assign n12409 = ~n12403 & n12408;
  assign n12410 = n12405 & ~n12407;
  assign n12411 = ~n12409 & ~n12410;
  assign n12412 = ~n12400 & ~n12411;
  assign n12413 = ~n12400 & ~n12412;
  assign n12414 = ~n12411 & ~n12412;
  assign n12415 = ~n12413 & ~n12414;
  assign n12416 = pi25  & pi53 ;
  assign n12417 = n1990 & n6911;
  assign n12418 = pi24  & pi54 ;
  assign n12419 = pi22  & pi56 ;
  assign n12420 = ~n12418 & ~n12419;
  assign n12421 = n12416 & ~n12417;
  assign n12422 = ~n12420 & n12421;
  assign n12423 = n12416 & ~n12422;
  assign n12424 = ~n12417 & ~n12422;
  assign n12425 = ~n12420 & n12424;
  assign n12426 = ~n12423 & ~n12425;
  assign n12427 = ~n12415 & ~n12426;
  assign n12428 = ~n12415 & ~n12427;
  assign n12429 = ~n12426 & ~n12427;
  assign n12430 = ~n12428 & ~n12429;
  assign n12431 = ~n12389 & n12430;
  assign n12432 = n12389 & ~n12430;
  assign n12433 = ~n12431 & ~n12432;
  assign n12434 = ~n12347 & ~n12433;
  assign n12435 = n12347 & n12433;
  assign n12436 = ~n12434 & ~n12435;
  assign n12437 = ~n12346 & n12436;
  assign n12438 = n12346 & ~n12436;
  assign n12439 = ~n12437 & ~n12438;
  assign n12440 = n12345 & ~n12439;
  assign n12441 = ~n12345 & n12439;
  assign n12442 = ~n12440 & ~n12441;
  assign n12443 = ~n12237 & ~n12330;
  assign n12444 = n12442 & ~n12443;
  assign n12445 = ~n12442 & n12443;
  assign n12446 = ~n12444 & ~n12445;
  assign n12447 = ~n12182 & ~n12185;
  assign n12448 = ~n12054 & ~n12305;
  assign n12449 = ~n12320 & ~n12448;
  assign n12450 = ~n12275 & ~n12287;
  assign n12451 = n12449 & n12450;
  assign n12452 = ~n12449 & ~n12450;
  assign n12453 = ~n12451 & ~n12452;
  assign n12454 = ~n12155 & ~n12170;
  assign n12455 = ~n12453 & n12454;
  assign n12456 = n12453 & ~n12454;
  assign n12457 = ~n12455 & ~n12456;
  assign n12458 = ~n12228 & ~n12230;
  assign n12459 = n12457 & ~n12458;
  assign n12460 = ~n12457 & n12458;
  assign n12461 = ~n12459 & ~n12460;
  assign n12462 = n12272 & n12282;
  assign n12463 = ~n12272 & ~n12282;
  assign n12464 = ~n12462 & ~n12463;
  assign n12465 = n12152 & ~n12464;
  assign n12466 = ~n12152 & n12464;
  assign n12467 = ~n12465 & ~n12466;
  assign n12468 = n12260 & n12317;
  assign n12469 = ~n12260 & ~n12317;
  assign n12470 = ~n12468 & ~n12469;
  assign n12471 = n12167 & ~n12470;
  assign n12472 = ~n12167 & n12470;
  assign n12473 = ~n12471 & ~n12472;
  assign n12474 = ~n12221 & ~n12224;
  assign n12475 = ~n12473 & n12474;
  assign n12476 = n12473 & ~n12474;
  assign n12477 = ~n12475 & ~n12476;
  assign n12478 = n12467 & n12477;
  assign n12479 = ~n12467 & ~n12477;
  assign n12480 = ~n12478 & ~n12479;
  assign n12481 = n12461 & n12480;
  assign n12482 = ~n12461 & ~n12480;
  assign n12483 = ~n12481 & ~n12482;
  assign n12484 = n12447 & ~n12483;
  assign n12485 = ~n12447 & n12483;
  assign n12486 = ~n12484 & ~n12485;
  assign n12487 = ~n12175 & ~n12179;
  assign n12488 = ~n12293 & ~n12323;
  assign n12489 = ~n12487 & ~n12488;
  assign n12490 = ~n12487 & ~n12489;
  assign n12491 = ~n12488 & ~n12489;
  assign n12492 = ~n12490 & ~n12491;
  assign n12493 = pi36  & pi42 ;
  assign n12494 = ~n5259 & ~n12493;
  assign n12495 = n4691 & n6458;
  assign n12496 = pi23  & pi55 ;
  assign n12497 = ~n12494 & n12496;
  assign n12498 = ~n12495 & n12497;
  assign n12499 = ~n12495 & ~n12498;
  assign n12500 = ~n12494 & n12499;
  assign n12501 = n12496 & ~n12498;
  assign n12502 = ~n12500 & ~n12501;
  assign n12503 = pi26  & pi52 ;
  assign n12504 = n3558 & n12503;
  assign n12505 = ~n3558 & ~n12503;
  assign n12506 = n5532 & ~n12504;
  assign n12507 = ~n12505 & n12506;
  assign n12508 = n5532 & ~n12507;
  assign n12509 = ~n12504 & ~n12507;
  assign n12510 = ~n12505 & n12509;
  assign n12511 = ~n12508 & ~n12510;
  assign n12512 = ~n12502 & ~n12511;
  assign n12513 = ~n12502 & ~n12512;
  assign n12514 = ~n12511 & ~n12512;
  assign n12515 = ~n12513 & ~n12514;
  assign n12516 = ~n12215 & ~n12218;
  assign n12517 = n12515 & n12516;
  assign n12518 = ~n12515 & ~n12516;
  assign n12519 = ~n12517 & ~n12518;
  assign n12520 = n12140 & n12303;
  assign n12521 = ~n12140 & ~n12303;
  assign n12522 = ~n12520 & ~n12521;
  assign n12523 = ~n12192 & ~n12198;
  assign n12524 = ~n12522 & n12523;
  assign n12525 = n12522 & ~n12523;
  assign n12526 = ~n12524 & ~n12525;
  assign n12527 = ~n12204 & ~n12208;
  assign n12528 = ~n12526 & n12527;
  assign n12529 = n12526 & ~n12527;
  assign n12530 = ~n12528 & ~n12529;
  assign n12531 = n12519 & n12530;
  assign n12532 = ~n12519 & ~n12530;
  assign n12533 = ~n12531 & ~n12532;
  assign n12534 = ~n12492 & n12533;
  assign n12535 = ~n12492 & ~n12534;
  assign n12536 = n12533 & ~n12534;
  assign n12537 = ~n12535 & ~n12536;
  assign n12538 = n12486 & ~n12537;
  assign n12539 = ~n12486 & n12537;
  assign n12540 = ~n12538 & ~n12539;
  assign n12541 = n12446 & n12540;
  assign n12542 = n12446 & ~n12541;
  assign n12543 = n12540 & ~n12541;
  assign n12544 = ~n12542 & ~n12543;
  assign n12545 = ~n12344 & ~n12544;
  assign n12546 = n12344 & n12544;
  assign n12547 = ~n12545 & ~n12546;
  assign n12548 = ~n12337 & ~n12342;
  assign n12549 = n12547 & ~n12548;
  assign n12550 = ~n12547 & n12548;
  assign po79  = ~n12549 & ~n12550;
  assign n12552 = ~n12444 & ~n12541;
  assign n12553 = ~n12489 & ~n12534;
  assign n12554 = ~n12389 & ~n12430;
  assign n12555 = ~n12434 & ~n12554;
  assign n12556 = n12356 & n12368;
  assign n12557 = ~n12356 & ~n12368;
  assign n12558 = ~n12556 & ~n12557;
  assign n12559 = n12424 & ~n12558;
  assign n12560 = ~n12424 & n12558;
  assign n12561 = ~n12559 & ~n12560;
  assign n12562 = ~n12512 & ~n12518;
  assign n12563 = ~n12561 & n12562;
  assign n12564 = n12561 & ~n12562;
  assign n12565 = ~n12563 & ~n12564;
  assign n12566 = pi34  & pi45 ;
  assign n12567 = pi35  & pi44 ;
  assign n12568 = ~n12566 & ~n12567;
  assign n12569 = n3106 & n5318;
  assign n12570 = pi16  & pi63 ;
  assign n12571 = ~n12568 & n12570;
  assign n12572 = ~n12569 & n12571;
  assign n12573 = ~n12569 & ~n12572;
  assign n12574 = ~n12568 & n12573;
  assign n12575 = n12570 & ~n12572;
  assign n12576 = ~n12574 & ~n12575;
  assign n12577 = pi36  & pi43 ;
  assign n12578 = pi27  & pi56 ;
  assign n12579 = n11754 & n12578;
  assign n12580 = pi23  & pi56 ;
  assign n12581 = pi27  & pi52 ;
  assign n12582 = ~n12580 & ~n12581;
  assign n12583 = n12577 & ~n12579;
  assign n12584 = ~n12582 & n12583;
  assign n12585 = n12577 & ~n12584;
  assign n12586 = ~n12579 & ~n12584;
  assign n12587 = ~n12582 & n12586;
  assign n12588 = ~n12585 & ~n12587;
  assign n12589 = ~n12576 & ~n12588;
  assign n12590 = ~n12576 & ~n12589;
  assign n12591 = ~n12588 & ~n12589;
  assign n12592 = ~n12590 & ~n12591;
  assign n12593 = ~n12521 & ~n12525;
  assign n12594 = n12592 & n12593;
  assign n12595 = ~n12592 & ~n12593;
  assign n12596 = ~n12594 & ~n12595;
  assign n12597 = n12565 & n12596;
  assign n12598 = ~n12565 & ~n12596;
  assign n12599 = ~n12597 & ~n12598;
  assign n12600 = n12555 & ~n12599;
  assign n12601 = ~n12555 & n12599;
  assign n12602 = ~n12600 & ~n12601;
  assign n12603 = ~n12412 & ~n12427;
  assign n12604 = pi18  & pi61 ;
  assign n12605 = ~n12509 & n12604;
  assign n12606 = n12509 & ~n12604;
  assign n12607 = ~n12605 & ~n12606;
  assign n12608 = n12499 & ~n12607;
  assign n12609 = ~n12499 & n12607;
  assign n12610 = ~n12608 & ~n12609;
  assign n12611 = n12383 & n12397;
  assign n12612 = ~n12383 & ~n12397;
  assign n12613 = ~n12611 & ~n12612;
  assign n12614 = n12408 & ~n12613;
  assign n12615 = ~n12408 & n12613;
  assign n12616 = ~n12614 & ~n12615;
  assign n12617 = n12610 & n12616;
  assign n12618 = ~n12610 & ~n12616;
  assign n12619 = ~n12617 & ~n12618;
  assign n12620 = ~n12603 & n12619;
  assign n12621 = n12603 & ~n12619;
  assign n12622 = ~n12620 & ~n12621;
  assign n12623 = n12602 & n12622;
  assign n12624 = ~n12602 & ~n12622;
  assign n12625 = ~n12623 & ~n12624;
  assign n12626 = n12553 & ~n12625;
  assign n12627 = ~n12553 & n12625;
  assign n12628 = ~n12626 & ~n12627;
  assign n12629 = ~n12437 & ~n12441;
  assign n12630 = ~n12628 & n12629;
  assign n12631 = n12628 & ~n12629;
  assign n12632 = ~n12630 & ~n12631;
  assign n12633 = ~n12459 & ~n12481;
  assign n12634 = ~n12476 & ~n12478;
  assign n12635 = pi25  & pi54 ;
  assign n12636 = pi26  & pi53 ;
  assign n12637 = ~n12635 & ~n12636;
  assign n12638 = n2310 & n8092;
  assign n12639 = pi24  & pi55 ;
  assign n12640 = ~n12637 & n12639;
  assign n12641 = ~n12638 & n12640;
  assign n12642 = ~n12638 & ~n12641;
  assign n12643 = ~n12637 & n12642;
  assign n12644 = n12639 & ~n12641;
  assign n12645 = ~n12643 & ~n12644;
  assign n12646 = pi37  & pi42 ;
  assign n12647 = n4736 & n6012;
  assign n12648 = pi38  & pi41 ;
  assign n12649 = ~n5548 & ~n12648;
  assign n12650 = n12646 & ~n12647;
  assign n12651 = ~n12649 & n12650;
  assign n12652 = n12646 & ~n12651;
  assign n12653 = ~n12647 & ~n12651;
  assign n12654 = ~n12649 & n12653;
  assign n12655 = ~n12652 & ~n12654;
  assign n12656 = ~n12645 & ~n12655;
  assign n12657 = ~n12645 & ~n12656;
  assign n12658 = ~n12655 & ~n12656;
  assign n12659 = ~n12657 & ~n12658;
  assign n12660 = pi28  & pi51 ;
  assign n12661 = pi40  & pi62 ;
  assign n12662 = pi17  & n12661;
  assign n12663 = pi17  & pi62 ;
  assign n12664 = ~pi40  & ~n12663;
  assign n12665 = n12660 & ~n12662;
  assign n12666 = ~n12664 & n12665;
  assign n12667 = n12660 & ~n12666;
  assign n12668 = ~n12662 & ~n12666;
  assign n12669 = ~n12664 & n12668;
  assign n12670 = ~n12667 & ~n12669;
  assign n12671 = ~n12659 & ~n12670;
  assign n12672 = ~n12659 & ~n12671;
  assign n12673 = ~n12670 & ~n12671;
  assign n12674 = ~n12672 & ~n12673;
  assign n12675 = pi20  & pi59 ;
  assign n12676 = pi21  & pi58 ;
  assign n12677 = ~n12675 & ~n12676;
  assign n12678 = n1593 & n9402;
  assign n12679 = pi19  & pi60 ;
  assign n12680 = ~n12677 & n12679;
  assign n12681 = ~n12678 & n12680;
  assign n12682 = ~n12678 & ~n12681;
  assign n12683 = ~n12677 & n12682;
  assign n12684 = n12679 & ~n12681;
  assign n12685 = ~n12683 & ~n12684;
  assign n12686 = pi22  & pi57 ;
  assign n12687 = n4908 & n5889;
  assign n12688 = pi29  & pi50 ;
  assign n12689 = pi30  & pi49 ;
  assign n12690 = ~n12688 & ~n12689;
  assign n12691 = n12686 & ~n12687;
  assign n12692 = ~n12690 & n12691;
  assign n12693 = n12686 & ~n12692;
  assign n12694 = ~n12687 & ~n12692;
  assign n12695 = ~n12690 & n12694;
  assign n12696 = ~n12693 & ~n12695;
  assign n12697 = ~n12685 & ~n12696;
  assign n12698 = ~n12685 & ~n12697;
  assign n12699 = ~n12696 & ~n12697;
  assign n12700 = ~n12698 & ~n12699;
  assign n12701 = pi31  & pi48 ;
  assign n12702 = n5277 & n6138;
  assign n12703 = pi32  & pi47 ;
  assign n12704 = ~n5490 & ~n12703;
  assign n12705 = n12701 & ~n12702;
  assign n12706 = ~n12704 & n12705;
  assign n12707 = n12701 & ~n12706;
  assign n12708 = ~n12702 & ~n12706;
  assign n12709 = ~n12704 & n12708;
  assign n12710 = ~n12707 & ~n12709;
  assign n12711 = ~n12700 & ~n12710;
  assign n12712 = ~n12700 & ~n12711;
  assign n12713 = ~n12710 & ~n12711;
  assign n12714 = ~n12712 & ~n12713;
  assign n12715 = n12674 & n12714;
  assign n12716 = ~n12674 & ~n12714;
  assign n12717 = ~n12715 & ~n12716;
  assign n12718 = ~n12634 & n12717;
  assign n12719 = n12634 & ~n12717;
  assign n12720 = ~n12718 & ~n12719;
  assign n12721 = n12633 & ~n12720;
  assign n12722 = ~n12633 & n12720;
  assign n12723 = ~n12721 & ~n12722;
  assign n12724 = ~n12469 & ~n12472;
  assign n12725 = ~n12463 & ~n12466;
  assign n12726 = n12724 & n12725;
  assign n12727 = ~n12724 & ~n12725;
  assign n12728 = ~n12726 & ~n12727;
  assign n12729 = ~n12371 & ~n12386;
  assign n12730 = ~n12728 & n12729;
  assign n12731 = n12728 & ~n12729;
  assign n12732 = ~n12730 & ~n12731;
  assign n12733 = ~n12452 & ~n12456;
  assign n12734 = ~n12732 & n12733;
  assign n12735 = n12732 & ~n12733;
  assign n12736 = ~n12734 & ~n12735;
  assign n12737 = ~n12529 & ~n12531;
  assign n12738 = n12736 & ~n12737;
  assign n12739 = ~n12736 & n12737;
  assign n12740 = ~n12738 & ~n12739;
  assign n12741 = n12723 & n12740;
  assign n12742 = ~n12723 & ~n12740;
  assign n12743 = ~n12741 & ~n12742;
  assign n12744 = ~n12485 & ~n12538;
  assign n12745 = n12743 & ~n12744;
  assign n12746 = n12743 & ~n12745;
  assign n12747 = ~n12744 & ~n12745;
  assign n12748 = ~n12746 & ~n12747;
  assign n12749 = n12632 & ~n12748;
  assign n12750 = ~n12632 & n12748;
  assign n12751 = ~n12749 & ~n12750;
  assign n12752 = ~n12552 & n12751;
  assign n12753 = n12552 & ~n12751;
  assign n12754 = ~n12752 & ~n12753;
  assign n12755 = ~n12545 & ~n12549;
  assign n12756 = ~n12754 & n12755;
  assign n12757 = n12754 & ~n12755;
  assign po80  = ~n12756 & ~n12757;
  assign n12759 = ~n12745 & ~n12749;
  assign n12760 = ~n12627 & ~n12631;
  assign n12761 = ~n12601 & ~n12623;
  assign n12762 = ~n12735 & ~n12738;
  assign n12763 = pi17  & pi63 ;
  assign n12764 = pi29  & pi51 ;
  assign n12765 = ~n12763 & ~n12764;
  assign n12766 = pi29  & pi63 ;
  assign n12767 = n7238 & n12766;
  assign n12768 = pi33  & pi47 ;
  assign n12769 = ~n12765 & n12768;
  assign n12770 = ~n12767 & n12769;
  assign n12771 = ~n12767 & ~n12770;
  assign n12772 = ~n12765 & n12771;
  assign n12773 = n12768 & ~n12770;
  assign n12774 = ~n12772 & ~n12773;
  assign n12775 = pi34  & pi46 ;
  assign n12776 = n4691 & n5318;
  assign n12777 = pi36  & pi44 ;
  assign n12778 = ~n5450 & ~n12777;
  assign n12779 = n12775 & ~n12776;
  assign n12780 = ~n12778 & n12779;
  assign n12781 = n12775 & ~n12780;
  assign n12782 = ~n12776 & ~n12780;
  assign n12783 = ~n12778 & n12782;
  assign n12784 = ~n12781 & ~n12783;
  assign n12785 = ~n12774 & ~n12784;
  assign n12786 = ~n12774 & ~n12785;
  assign n12787 = ~n12784 & ~n12785;
  assign n12788 = ~n12786 & ~n12787;
  assign n12789 = n1085 & n9567;
  assign n12790 = pi19  & pi61 ;
  assign n12791 = ~n12789 & n12790;
  assign n12792 = pi18  & pi62 ;
  assign n12793 = ~n12789 & n12792;
  assign n12794 = ~n12791 & ~n12793;
  assign n12795 = ~n12668 & ~n12794;
  assign n12796 = ~n12668 & ~n12795;
  assign n12797 = ~n12794 & ~n12795;
  assign n12798 = ~n12796 & ~n12797;
  assign n12799 = ~n12788 & n12798;
  assign n12800 = n12788 & ~n12798;
  assign n12801 = ~n12799 & ~n12800;
  assign n12802 = n1481 & n9402;
  assign n12803 = pi21  & pi59 ;
  assign n12804 = pi22  & pi58 ;
  assign n12805 = ~n12803 & ~n12804;
  assign n12806 = ~n12802 & ~n12805;
  assign n12807 = pi20  & pi60 ;
  assign n12808 = ~n12806 & ~n12807;
  assign n12809 = n12806 & n12807;
  assign n12810 = ~n12808 & ~n12809;
  assign n12811 = ~n12653 & n12810;
  assign n12812 = n12653 & ~n12810;
  assign n12813 = ~n12811 & ~n12812;
  assign n12814 = pi30  & pi50 ;
  assign n12815 = n3567 & n8505;
  assign n12816 = pi31  & pi49 ;
  assign n12817 = pi32  & pi48 ;
  assign n12818 = ~n12816 & ~n12817;
  assign n12819 = n12814 & ~n12815;
  assign n12820 = ~n12818 & n12819;
  assign n12821 = n12814 & ~n12820;
  assign n12822 = ~n12815 & ~n12820;
  assign n12823 = ~n12818 & n12822;
  assign n12824 = ~n12821 & ~n12823;
  assign n12825 = n12813 & ~n12824;
  assign n12826 = n12813 & ~n12825;
  assign n12827 = ~n12824 & ~n12825;
  assign n12828 = ~n12826 & ~n12827;
  assign n12829 = pi24  & pi56 ;
  assign n12830 = pi26  & pi54 ;
  assign n12831 = ~n12829 & ~n12830;
  assign n12832 = n2167 & n6911;
  assign n12833 = pi23  & pi57 ;
  assign n12834 = ~n12831 & n12833;
  assign n12835 = ~n12832 & n12834;
  assign n12836 = ~n12832 & ~n12835;
  assign n12837 = ~n12831 & n12836;
  assign n12838 = n12833 & ~n12835;
  assign n12839 = ~n12837 & ~n12838;
  assign n12840 = pi25  & pi55 ;
  assign n12841 = n5055 & n6458;
  assign n12842 = pi37  & pi43 ;
  assign n12843 = pi38  & pi42 ;
  assign n12844 = ~n12842 & ~n12843;
  assign n12845 = n12840 & ~n12841;
  assign n12846 = ~n12844 & n12845;
  assign n12847 = n12840 & ~n12846;
  assign n12848 = ~n12841 & ~n12846;
  assign n12849 = ~n12844 & n12848;
  assign n12850 = ~n12847 & ~n12849;
  assign n12851 = ~n12839 & ~n12850;
  assign n12852 = ~n12839 & ~n12851;
  assign n12853 = ~n12850 & ~n12851;
  assign n12854 = ~n12852 & ~n12853;
  assign n12855 = n2191 & n9144;
  assign n12856 = pi27  & pi53 ;
  assign n12857 = pi28  & pi52 ;
  assign n12858 = ~n12856 & ~n12857;
  assign n12859 = n3729 & ~n12855;
  assign n12860 = ~n12858 & n12859;
  assign n12861 = n3729 & ~n12860;
  assign n12862 = ~n12855 & ~n12860;
  assign n12863 = ~n12858 & n12862;
  assign n12864 = ~n12861 & ~n12863;
  assign n12865 = ~n12854 & ~n12864;
  assign n12866 = ~n12854 & ~n12865;
  assign n12867 = ~n12864 & ~n12865;
  assign n12868 = ~n12866 & ~n12867;
  assign n12869 = ~n12828 & n12868;
  assign n12870 = n12828 & ~n12868;
  assign n12871 = ~n12869 & ~n12870;
  assign n12872 = ~n12801 & ~n12871;
  assign n12873 = n12801 & n12871;
  assign n12874 = ~n12872 & ~n12873;
  assign n12875 = ~n12762 & n12874;
  assign n12876 = n12762 & ~n12874;
  assign n12877 = ~n12875 & ~n12876;
  assign n12878 = ~n12761 & n12877;
  assign n12879 = n12761 & ~n12877;
  assign n12880 = ~n12878 & ~n12879;
  assign n12881 = n12760 & ~n12880;
  assign n12882 = ~n12760 & n12880;
  assign n12883 = ~n12881 & ~n12882;
  assign n12884 = ~n12722 & ~n12741;
  assign n12885 = ~n12716 & ~n12718;
  assign n12886 = n12573 & n12642;
  assign n12887 = ~n12573 & ~n12642;
  assign n12888 = ~n12886 & ~n12887;
  assign n12889 = n12586 & ~n12888;
  assign n12890 = ~n12586 & n12888;
  assign n12891 = ~n12889 & ~n12890;
  assign n12892 = ~n12589 & ~n12595;
  assign n12893 = ~n12891 & n12892;
  assign n12894 = n12891 & ~n12892;
  assign n12895 = ~n12893 & ~n12894;
  assign n12896 = ~n12727 & ~n12731;
  assign n12897 = ~n12895 & n12896;
  assign n12898 = n12895 & ~n12896;
  assign n12899 = ~n12897 & ~n12898;
  assign n12900 = ~n12885 & n12899;
  assign n12901 = n12885 & ~n12899;
  assign n12902 = ~n12900 & ~n12901;
  assign n12903 = n12682 & n12694;
  assign n12904 = ~n12682 & ~n12694;
  assign n12905 = ~n12903 & ~n12904;
  assign n12906 = n12708 & ~n12905;
  assign n12907 = ~n12708 & n12905;
  assign n12908 = ~n12906 & ~n12907;
  assign n12909 = ~n12656 & ~n12671;
  assign n12910 = ~n12697 & ~n12711;
  assign n12911 = n12909 & n12910;
  assign n12912 = ~n12909 & ~n12910;
  assign n12913 = ~n12911 & ~n12912;
  assign n12914 = n12908 & n12913;
  assign n12915 = ~n12908 & ~n12913;
  assign n12916 = ~n12914 & ~n12915;
  assign n12917 = n12902 & n12916;
  assign n12918 = ~n12902 & ~n12916;
  assign n12919 = ~n12917 & ~n12918;
  assign n12920 = ~n12557 & ~n12560;
  assign n12921 = ~n12612 & ~n12615;
  assign n12922 = n12920 & n12921;
  assign n12923 = ~n12920 & ~n12921;
  assign n12924 = ~n12922 & ~n12923;
  assign n12925 = ~n12605 & ~n12609;
  assign n12926 = ~n12924 & n12925;
  assign n12927 = n12924 & ~n12925;
  assign n12928 = ~n12926 & ~n12927;
  assign n12929 = ~n12564 & ~n12597;
  assign n12930 = ~n12617 & ~n12620;
  assign n12931 = ~n12929 & ~n12930;
  assign n12932 = ~n12929 & ~n12931;
  assign n12933 = ~n12930 & ~n12931;
  assign n12934 = ~n12932 & ~n12933;
  assign n12935 = ~n12928 & n12934;
  assign n12936 = n12928 & ~n12934;
  assign n12937 = ~n12935 & ~n12936;
  assign n12938 = n12919 & n12937;
  assign n12939 = n12919 & ~n12938;
  assign n12940 = n12937 & ~n12938;
  assign n12941 = ~n12939 & ~n12940;
  assign n12942 = ~n12884 & ~n12941;
  assign n12943 = n12884 & n12941;
  assign n12944 = ~n12942 & ~n12943;
  assign n12945 = n12883 & n12944;
  assign n12946 = ~n12883 & ~n12944;
  assign n12947 = ~n12945 & ~n12946;
  assign n12948 = n12759 & ~n12947;
  assign n12949 = ~n12759 & n12947;
  assign n12950 = ~n12948 & ~n12949;
  assign n12951 = ~n12752 & ~n12757;
  assign n12952 = ~n12950 & n12951;
  assign n12953 = ~n12948 & ~n12951;
  assign n12954 = ~n12949 & n12953;
  assign po81  = ~n12952 & ~n12954;
  assign n12956 = ~n12949 & ~n12953;
  assign n12957 = ~n12938 & ~n12942;
  assign n12958 = ~n12900 & ~n12917;
  assign n12959 = ~n12931 & ~n12936;
  assign n12960 = pi41  & pi62 ;
  assign n12961 = pi19  & n12960;
  assign n12962 = n6012 & ~n12961;
  assign n12963 = ~n12961 & ~n12962;
  assign n12964 = pi19  & pi62 ;
  assign n12965 = ~pi41  & ~n12964;
  assign n12966 = n12963 & ~n12965;
  assign n12967 = n6012 & ~n12962;
  assign n12968 = ~n12966 & ~n12967;
  assign n12969 = pi22  & pi59 ;
  assign n12970 = pi56  & pi58 ;
  assign n12971 = n1457 & n12970;
  assign n12972 = pi23  & pi58 ;
  assign n12973 = ~n11558 & ~n12972;
  assign n12974 = n12969 & ~n12971;
  assign n12975 = ~n12973 & n12974;
  assign n12976 = n12969 & ~n12975;
  assign n12977 = ~n12971 & ~n12975;
  assign n12978 = ~n12973 & n12977;
  assign n12979 = ~n12976 & ~n12978;
  assign n12980 = ~n12968 & ~n12979;
  assign n12981 = ~n12968 & ~n12980;
  assign n12982 = ~n12979 & ~n12980;
  assign n12983 = ~n12981 & ~n12982;
  assign n12984 = n3900 & n5823;
  assign n12985 = pi33  & pi48 ;
  assign n12986 = pi34  & pi47 ;
  assign n12987 = ~n12985 & ~n12986;
  assign n12988 = n9609 & ~n12984;
  assign n12989 = ~n12987 & n12988;
  assign n12990 = n9609 & ~n12989;
  assign n12991 = ~n12984 & ~n12989;
  assign n12992 = ~n12987 & n12991;
  assign n12993 = ~n12990 & ~n12992;
  assign n12994 = ~n12983 & ~n12993;
  assign n12995 = ~n12983 & ~n12994;
  assign n12996 = ~n12993 & ~n12994;
  assign n12997 = ~n12995 & ~n12996;
  assign n12998 = ~n12923 & ~n12927;
  assign n12999 = n12997 & n12998;
  assign n13000 = ~n12997 & ~n12998;
  assign n13001 = ~n12999 & ~n13000;
  assign n13002 = pi20  & pi61 ;
  assign n13003 = pi21  & pi60 ;
  assign n13004 = ~n13002 & ~n13003;
  assign n13005 = n1593 & n9054;
  assign n13006 = pi18  & pi63 ;
  assign n13007 = ~n13004 & n13006;
  assign n13008 = ~n13005 & n13007;
  assign n13009 = ~n13005 & ~n13008;
  assign n13010 = ~n13004 & n13009;
  assign n13011 = n13006 & ~n13008;
  assign n13012 = ~n13010 & ~n13011;
  assign n13013 = pi35  & pi46 ;
  assign n13014 = n4500 & n5318;
  assign n13015 = pi37  & pi44 ;
  assign n13016 = pi36  & pi45 ;
  assign n13017 = ~n13015 & ~n13016;
  assign n13018 = n13013 & ~n13014;
  assign n13019 = ~n13017 & n13018;
  assign n13020 = n13013 & ~n13019;
  assign n13021 = ~n13014 & ~n13019;
  assign n13022 = ~n13017 & n13021;
  assign n13023 = ~n13020 & ~n13022;
  assign n13024 = ~n13012 & ~n13023;
  assign n13025 = ~n13012 & ~n13024;
  assign n13026 = ~n13023 & ~n13024;
  assign n13027 = ~n13025 & ~n13026;
  assign n13028 = pi26  & pi55 ;
  assign n13029 = n2915 & n9144;
  assign n13030 = pi28  & pi53 ;
  assign n13031 = pi29  & pi52 ;
  assign n13032 = ~n13030 & ~n13031;
  assign n13033 = n13028 & ~n13029;
  assign n13034 = ~n13032 & n13033;
  assign n13035 = n13028 & ~n13034;
  assign n13036 = ~n13029 & ~n13034;
  assign n13037 = ~n13032 & n13036;
  assign n13038 = ~n13035 & ~n13037;
  assign n13039 = ~n13027 & ~n13038;
  assign n13040 = ~n13027 & ~n13039;
  assign n13041 = ~n13038 & ~n13039;
  assign n13042 = ~n13040 & ~n13041;
  assign n13043 = ~n13001 & n13042;
  assign n13044 = n13001 & ~n13042;
  assign n13045 = ~n13043 & ~n13044;
  assign n13046 = ~n12959 & n13045;
  assign n13047 = ~n12959 & ~n13046;
  assign n13048 = n13045 & ~n13046;
  assign n13049 = ~n13047 & ~n13048;
  assign n13050 = ~n12958 & ~n13049;
  assign n13051 = ~n12958 & ~n13050;
  assign n13052 = ~n13049 & ~n13050;
  assign n13053 = ~n13051 & ~n13052;
  assign n13054 = ~n12957 & ~n13053;
  assign n13055 = ~n12957 & ~n13054;
  assign n13056 = ~n13053 & ~n13054;
  assign n13057 = ~n13055 & ~n13056;
  assign n13058 = ~n12875 & ~n12878;
  assign n13059 = ~n12904 & ~n12907;
  assign n13060 = pi27  & pi54 ;
  assign n13061 = n4736 & n6458;
  assign n13062 = pi38  & pi43 ;
  assign n13063 = pi39  & pi42 ;
  assign n13064 = ~n13062 & ~n13063;
  assign n13065 = n13060 & ~n13061;
  assign n13066 = ~n13064 & n13065;
  assign n13067 = n13060 & ~n13066;
  assign n13068 = ~n13061 & ~n13066;
  assign n13069 = ~n13064 & n13068;
  assign n13070 = ~n13067 & ~n13069;
  assign n13071 = ~n13059 & ~n13070;
  assign n13072 = ~n13059 & ~n13071;
  assign n13073 = ~n13070 & ~n13071;
  assign n13074 = ~n13072 & ~n13073;
  assign n13075 = ~n12887 & ~n12890;
  assign n13076 = n13074 & n13075;
  assign n13077 = ~n13074 & ~n13075;
  assign n13078 = ~n13076 & ~n13077;
  assign n13079 = ~n12894 & ~n12898;
  assign n13080 = ~n12912 & ~n12914;
  assign n13081 = ~n13079 & ~n13080;
  assign n13082 = ~n13079 & ~n13081;
  assign n13083 = ~n13080 & ~n13081;
  assign n13084 = ~n13082 & ~n13083;
  assign n13085 = n13078 & ~n13084;
  assign n13086 = ~n13078 & n13084;
  assign n13087 = ~n13085 & ~n13086;
  assign n13088 = ~n13058 & n13087;
  assign n13089 = ~n13058 & ~n13088;
  assign n13090 = n13087 & ~n13088;
  assign n13091 = ~n13089 & ~n13090;
  assign n13092 = ~n12789 & ~n12795;
  assign n13093 = n12782 & n13092;
  assign n13094 = ~n12782 & ~n13092;
  assign n13095 = ~n13093 & ~n13094;
  assign n13096 = pi30  & pi51 ;
  assign n13097 = n3567 & n5889;
  assign n13098 = pi31  & pi50 ;
  assign n13099 = pi32  & pi49 ;
  assign n13100 = ~n13098 & ~n13099;
  assign n13101 = n13096 & ~n13097;
  assign n13102 = ~n13100 & n13101;
  assign n13103 = n13096 & ~n13102;
  assign n13104 = ~n13097 & ~n13102;
  assign n13105 = ~n13100 & n13104;
  assign n13106 = ~n13103 & ~n13105;
  assign n13107 = n13095 & ~n13106;
  assign n13108 = n13095 & ~n13107;
  assign n13109 = ~n13106 & ~n13107;
  assign n13110 = ~n13108 & ~n13109;
  assign n13111 = n12771 & n12822;
  assign n13112 = ~n12771 & ~n12822;
  assign n13113 = ~n13111 & ~n13112;
  assign n13114 = ~n12802 & ~n12809;
  assign n13115 = ~n13113 & n13114;
  assign n13116 = n13113 & ~n13114;
  assign n13117 = ~n13115 & ~n13116;
  assign n13118 = ~n12788 & ~n12798;
  assign n13119 = ~n12785 & ~n13118;
  assign n13120 = n13117 & ~n13119;
  assign n13121 = ~n13117 & n13119;
  assign n13122 = ~n13120 & ~n13121;
  assign n13123 = n13110 & n13122;
  assign n13124 = ~n13110 & ~n13122;
  assign n13125 = ~n13123 & ~n13124;
  assign n13126 = ~n12828 & ~n12868;
  assign n13127 = ~n12872 & ~n13126;
  assign n13128 = n13125 & n13127;
  assign n13129 = ~n13125 & ~n13127;
  assign n13130 = ~n13128 & ~n13129;
  assign n13131 = n12848 & n12862;
  assign n13132 = ~n12848 & ~n12862;
  assign n13133 = ~n13131 & ~n13132;
  assign n13134 = n12836 & ~n13133;
  assign n13135 = ~n12836 & n13133;
  assign n13136 = ~n13134 & ~n13135;
  assign n13137 = ~n12851 & ~n12865;
  assign n13138 = ~n12811 & ~n12825;
  assign n13139 = n13137 & n13138;
  assign n13140 = ~n13137 & ~n13138;
  assign n13141 = ~n13139 & ~n13140;
  assign n13142 = n13136 & n13141;
  assign n13143 = ~n13136 & ~n13141;
  assign n13144 = ~n13142 & ~n13143;
  assign n13145 = n13130 & n13144;
  assign n13146 = ~n13130 & ~n13144;
  assign n13147 = ~n13145 & ~n13146;
  assign n13148 = ~n13091 & ~n13147;
  assign n13149 = n13091 & n13147;
  assign n13150 = ~n13148 & ~n13149;
  assign n13151 = ~n13057 & ~n13150;
  assign n13152 = ~n13057 & ~n13151;
  assign n13153 = ~n13150 & ~n13151;
  assign n13154 = ~n13152 & ~n13153;
  assign n13155 = ~n12882 & ~n12945;
  assign n13156 = ~n13154 & ~n13155;
  assign n13157 = n13154 & n13155;
  assign n13158 = ~n13156 & ~n13157;
  assign n13159 = ~n12956 & ~n13158;
  assign n13160 = n12956 & n13158;
  assign po82  = n13159 | n13160;
  assign n13162 = ~n12956 & ~n13157;
  assign n13163 = ~n13156 & ~n13162;
  assign n13164 = ~n13054 & ~n13151;
  assign n13165 = ~n13091 & n13147;
  assign n13166 = ~n13088 & ~n13165;
  assign n13167 = ~n13129 & ~n13145;
  assign n13168 = ~n13081 & ~n13085;
  assign n13169 = pi31  & pi51 ;
  assign n13170 = pi21  & pi61 ;
  assign n13171 = ~n13169 & ~n13170;
  assign n13172 = n13169 & n13170;
  assign n13173 = pi20  & pi62 ;
  assign n13174 = ~n13171 & n13173;
  assign n13175 = ~n13172 & n13174;
  assign n13176 = ~n13172 & ~n13175;
  assign n13177 = ~n13171 & n13176;
  assign n13178 = n13173 & ~n13175;
  assign n13179 = ~n13177 & ~n13178;
  assign n13180 = pi32  & pi50 ;
  assign n13181 = n3900 & n8505;
  assign n13182 = pi33  & pi49 ;
  assign n13183 = pi34  & pi48 ;
  assign n13184 = ~n13182 & ~n13183;
  assign n13185 = n13180 & ~n13181;
  assign n13186 = ~n13184 & n13185;
  assign n13187 = n13180 & ~n13186;
  assign n13188 = ~n13181 & ~n13186;
  assign n13189 = ~n13184 & n13188;
  assign n13190 = ~n13187 & ~n13189;
  assign n13191 = ~n13179 & ~n13190;
  assign n13192 = ~n13179 & ~n13191;
  assign n13193 = ~n13190 & ~n13191;
  assign n13194 = ~n13192 & ~n13193;
  assign n13195 = pi22  & pi60 ;
  assign n13196 = n2110 & n9402;
  assign n13197 = pi24  & pi58 ;
  assign n13198 = pi23  & pi59 ;
  assign n13199 = ~n13197 & ~n13198;
  assign n13200 = n13195 & ~n13196;
  assign n13201 = ~n13199 & n13200;
  assign n13202 = n13195 & ~n13201;
  assign n13203 = ~n13196 & ~n13201;
  assign n13204 = ~n13199 & n13203;
  assign n13205 = ~n13202 & ~n13204;
  assign n13206 = ~n13194 & ~n13205;
  assign n13207 = ~n13194 & ~n13206;
  assign n13208 = ~n13205 & ~n13206;
  assign n13209 = ~n13207 & ~n13208;
  assign n13210 = ~n13071 & ~n13077;
  assign n13211 = n13209 & n13210;
  assign n13212 = ~n13209 & ~n13210;
  assign n13213 = ~n13211 & ~n13212;
  assign n13214 = pi38  & pi44 ;
  assign n13215 = pi39  & pi43 ;
  assign n13216 = ~n13214 & ~n13215;
  assign n13217 = n4736 & n6836;
  assign n13218 = pi26  & pi56 ;
  assign n13219 = ~n13216 & n13218;
  assign n13220 = ~n13217 & n13219;
  assign n13221 = ~n13217 & ~n13220;
  assign n13222 = ~n13216 & n13221;
  assign n13223 = n13218 & ~n13220;
  assign n13224 = ~n13222 & ~n13223;
  assign n13225 = pi40  & pi42 ;
  assign n13226 = n4908 & n9144;
  assign n13227 = pi29  & pi53 ;
  assign n13228 = pi30  & pi52 ;
  assign n13229 = ~n13227 & ~n13228;
  assign n13230 = n13225 & ~n13226;
  assign n13231 = ~n13229 & n13230;
  assign n13232 = n13225 & ~n13231;
  assign n13233 = ~n13226 & ~n13231;
  assign n13234 = ~n13229 & n13233;
  assign n13235 = ~n13232 & ~n13234;
  assign n13236 = ~n13224 & ~n13235;
  assign n13237 = ~n13224 & ~n13236;
  assign n13238 = ~n13235 & ~n13236;
  assign n13239 = ~n13237 & ~n13238;
  assign n13240 = pi35  & pi47 ;
  assign n13241 = n4500 & n7513;
  assign n13242 = ~n5725 & ~n6002;
  assign n13243 = n13240 & ~n13241;
  assign n13244 = ~n13242 & n13243;
  assign n13245 = n13240 & ~n13244;
  assign n13246 = ~n13241 & ~n13244;
  assign n13247 = ~n13242 & n13246;
  assign n13248 = ~n13245 & ~n13247;
  assign n13249 = ~n13239 & ~n13248;
  assign n13250 = ~n13239 & ~n13249;
  assign n13251 = ~n13248 & ~n13249;
  assign n13252 = ~n13250 & ~n13251;
  assign n13253 = ~n13213 & n13252;
  assign n13254 = n13213 & ~n13252;
  assign n13255 = ~n13253 & ~n13254;
  assign n13256 = ~n13168 & n13255;
  assign n13257 = ~n13168 & ~n13256;
  assign n13258 = n13255 & ~n13256;
  assign n13259 = ~n13257 & ~n13258;
  assign n13260 = ~n13167 & ~n13259;
  assign n13261 = ~n13167 & ~n13260;
  assign n13262 = ~n13259 & ~n13260;
  assign n13263 = ~n13261 & ~n13262;
  assign n13264 = ~n13166 & ~n13263;
  assign n13265 = ~n13166 & ~n13264;
  assign n13266 = ~n13263 & ~n13264;
  assign n13267 = ~n13265 & ~n13266;
  assign n13268 = ~n13046 & ~n13050;
  assign n13269 = ~n13112 & ~n13116;
  assign n13270 = pi55  & pi57 ;
  assign n13271 = n2468 & n13270;
  assign n13272 = pi25  & pi57 ;
  assign n13273 = pi27  & pi55 ;
  assign n13274 = ~n13272 & ~n13273;
  assign n13275 = n6636 & ~n13271;
  assign n13276 = ~n13274 & n13275;
  assign n13277 = n6636 & ~n13276;
  assign n13278 = ~n13271 & ~n13276;
  assign n13279 = ~n13274 & n13278;
  assign n13280 = ~n13277 & ~n13279;
  assign n13281 = ~n13269 & ~n13280;
  assign n13282 = ~n13269 & ~n13281;
  assign n13283 = ~n13280 & ~n13281;
  assign n13284 = ~n13282 & ~n13283;
  assign n13285 = ~n13132 & ~n13135;
  assign n13286 = n13284 & n13285;
  assign n13287 = ~n13284 & ~n13285;
  assign n13288 = ~n13286 & ~n13287;
  assign n13289 = ~n13121 & ~n13123;
  assign n13290 = ~n13140 & ~n13142;
  assign n13291 = n13289 & ~n13290;
  assign n13292 = n13289 & ~n13291;
  assign n13293 = ~n13290 & ~n13291;
  assign n13294 = ~n13292 & ~n13293;
  assign n13295 = n13288 & ~n13294;
  assign n13296 = ~n13288 & n13294;
  assign n13297 = ~n13295 & ~n13296;
  assign n13298 = ~n13268 & n13297;
  assign n13299 = ~n13268 & ~n13298;
  assign n13300 = n13297 & ~n13298;
  assign n13301 = ~n13299 & ~n13300;
  assign n13302 = ~n13000 & ~n13044;
  assign n13303 = n12991 & n13104;
  assign n13304 = ~n12991 & ~n13104;
  assign n13305 = ~n13303 & ~n13304;
  assign n13306 = n13036 & ~n13305;
  assign n13307 = ~n13036 & n13305;
  assign n13308 = ~n13306 & ~n13307;
  assign n13309 = n12977 & n13009;
  assign n13310 = ~n12977 & ~n13009;
  assign n13311 = ~n13309 & ~n13310;
  assign n13312 = n13021 & ~n13311;
  assign n13313 = ~n13021 & n13311;
  assign n13314 = ~n13312 & ~n13313;
  assign n13315 = ~n13024 & ~n13039;
  assign n13316 = ~n13314 & n13315;
  assign n13317 = n13314 & ~n13315;
  assign n13318 = ~n13316 & ~n13317;
  assign n13319 = n13308 & n13318;
  assign n13320 = ~n13308 & ~n13318;
  assign n13321 = ~n13319 & ~n13320;
  assign n13322 = n13302 & ~n13321;
  assign n13323 = ~n13302 & n13321;
  assign n13324 = ~n13322 & ~n13323;
  assign n13325 = ~n13094 & ~n13107;
  assign n13326 = ~n12980 & ~n12994;
  assign n13327 = n13325 & n13326;
  assign n13328 = ~n13325 & ~n13326;
  assign n13329 = ~n13327 & ~n13328;
  assign n13330 = n11745 & ~n12963;
  assign n13331 = ~n11745 & n12963;
  assign n13332 = ~n13330 & ~n13331;
  assign n13333 = n13068 & ~n13332;
  assign n13334 = ~n13068 & n13332;
  assign n13335 = ~n13333 & ~n13334;
  assign n13336 = n13329 & n13335;
  assign n13337 = ~n13329 & ~n13335;
  assign n13338 = ~n13336 & ~n13337;
  assign n13339 = n13324 & n13338;
  assign n13340 = ~n13324 & ~n13338;
  assign n13341 = ~n13339 & ~n13340;
  assign n13342 = ~n13301 & ~n13341;
  assign n13343 = n13301 & n13341;
  assign n13344 = ~n13342 & ~n13343;
  assign n13345 = ~n13267 & ~n13344;
  assign n13346 = ~n13267 & ~n13345;
  assign n13347 = ~n13344 & ~n13345;
  assign n13348 = ~n13346 & ~n13347;
  assign n13349 = ~n13164 & ~n13348;
  assign n13350 = n13164 & n13348;
  assign n13351 = ~n13349 & ~n13350;
  assign n13352 = ~n13163 & n13351;
  assign n13353 = n13163 & ~n13351;
  assign po83  = ~n13352 & ~n13353;
  assign n13355 = ~n13264 & ~n13345;
  assign n13356 = ~n13301 & n13341;
  assign n13357 = ~n13298 & ~n13356;
  assign n13358 = ~n13323 & ~n13339;
  assign n13359 = ~n13291 & ~n13295;
  assign n13360 = pi42  & pi62 ;
  assign n13361 = pi21  & n13360;
  assign n13362 = n5235 & ~n13361;
  assign n13363 = ~n13361 & ~n13362;
  assign n13364 = pi21  & pi62 ;
  assign n13365 = ~pi42  & ~n13364;
  assign n13366 = n13363 & ~n13365;
  assign n13367 = n5235 & ~n13362;
  assign n13368 = ~n13366 & ~n13367;
  assign n13369 = pi29  & pi54 ;
  assign n13370 = n5548 & n6836;
  assign n13371 = pi39  & pi44 ;
  assign n13372 = pi40  & pi43 ;
  assign n13373 = ~n13371 & ~n13372;
  assign n13374 = n13369 & ~n13370;
  assign n13375 = ~n13373 & n13374;
  assign n13376 = n13369 & ~n13375;
  assign n13377 = ~n13370 & ~n13375;
  assign n13378 = ~n13373 & n13377;
  assign n13379 = ~n13376 & ~n13378;
  assign n13380 = ~n13368 & ~n13379;
  assign n13381 = ~n13368 & ~n13380;
  assign n13382 = ~n13379 & ~n13380;
  assign n13383 = ~n13381 & ~n13382;
  assign n13384 = pi33  & pi50 ;
  assign n13385 = n3106 & n8505;
  assign n13386 = pi34  & pi49 ;
  assign n13387 = pi35  & pi48 ;
  assign n13388 = ~n13386 & ~n13387;
  assign n13389 = n13384 & ~n13385;
  assign n13390 = ~n13388 & n13389;
  assign n13391 = n13384 & ~n13390;
  assign n13392 = ~n13385 & ~n13390;
  assign n13393 = ~n13388 & n13392;
  assign n13394 = ~n13391 & ~n13393;
  assign n13395 = ~n13383 & ~n13394;
  assign n13396 = ~n13383 & ~n13395;
  assign n13397 = ~n13394 & ~n13395;
  assign n13398 = ~n13396 & ~n13397;
  assign n13399 = ~n13281 & ~n13287;
  assign n13400 = n13398 & n13399;
  assign n13401 = ~n13398 & ~n13399;
  assign n13402 = ~n13400 & ~n13401;
  assign n13403 = pi26  & pi57 ;
  assign n13404 = pi32  & pi51 ;
  assign n13405 = ~n13403 & ~n13404;
  assign n13406 = pi51  & pi57 ;
  assign n13407 = n7469 & n13406;
  assign n13408 = pi25  & pi58 ;
  assign n13409 = ~n13405 & n13408;
  assign n13410 = ~n13407 & n13409;
  assign n13411 = ~n13407 & ~n13410;
  assign n13412 = ~n13405 & n13411;
  assign n13413 = n13408 & ~n13410;
  assign n13414 = ~n13412 & ~n13413;
  assign n13415 = pi36  & pi47 ;
  assign n13416 = n5055 & n7513;
  assign n13417 = pi37  & pi46 ;
  assign n13418 = pi38  & pi45 ;
  assign n13419 = ~n13417 & ~n13418;
  assign n13420 = n13415 & ~n13416;
  assign n13421 = ~n13419 & n13420;
  assign n13422 = n13415 & ~n13421;
  assign n13423 = ~n13416 & ~n13421;
  assign n13424 = ~n13419 & n13423;
  assign n13425 = ~n13422 & ~n13424;
  assign n13426 = ~n13414 & ~n13425;
  assign n13427 = ~n13414 & ~n13426;
  assign n13428 = ~n13425 & ~n13426;
  assign n13429 = ~n13427 & ~n13428;
  assign n13430 = n3972 & n9236;
  assign n13431 = pi20  & pi63 ;
  assign n13432 = pi22  & pi61 ;
  assign n13433 = ~n13431 & ~n13432;
  assign n13434 = n12578 & ~n13430;
  assign n13435 = ~n13433 & n13434;
  assign n13436 = n12578 & ~n13435;
  assign n13437 = ~n13430 & ~n13435;
  assign n13438 = ~n13433 & n13437;
  assign n13439 = ~n13436 & ~n13438;
  assign n13440 = ~n13429 & ~n13439;
  assign n13441 = ~n13429 & ~n13440;
  assign n13442 = ~n13439 & ~n13440;
  assign n13443 = ~n13441 & ~n13442;
  assign n13444 = ~n13402 & n13443;
  assign n13445 = n13402 & ~n13443;
  assign n13446 = ~n13444 & ~n13445;
  assign n13447 = ~n13359 & n13446;
  assign n13448 = n13359 & ~n13446;
  assign n13449 = ~n13447 & ~n13448;
  assign n13450 = ~n13358 & n13449;
  assign n13451 = n13358 & ~n13449;
  assign n13452 = ~n13450 & ~n13451;
  assign n13453 = ~n13357 & n13452;
  assign n13454 = n13357 & ~n13452;
  assign n13455 = ~n13453 & ~n13454;
  assign n13456 = ~n13212 & ~n13254;
  assign n13457 = ~n13317 & ~n13319;
  assign n13458 = ~n13456 & ~n13457;
  assign n13459 = ~n13456 & ~n13458;
  assign n13460 = ~n13457 & ~n13458;
  assign n13461 = ~n13459 & ~n13460;
  assign n13462 = n13203 & n13246;
  assign n13463 = ~n13203 & ~n13246;
  assign n13464 = ~n13462 & ~n13463;
  assign n13465 = n13221 & ~n13464;
  assign n13466 = ~n13221 & n13464;
  assign n13467 = ~n13465 & ~n13466;
  assign n13468 = n13176 & n13188;
  assign n13469 = ~n13176 & ~n13188;
  assign n13470 = ~n13468 & ~n13469;
  assign n13471 = n13278 & ~n13470;
  assign n13472 = ~n13278 & n13470;
  assign n13473 = ~n13471 & ~n13472;
  assign n13474 = ~n13236 & ~n13249;
  assign n13475 = ~n13473 & n13474;
  assign n13476 = n13473 & ~n13474;
  assign n13477 = ~n13475 & ~n13476;
  assign n13478 = n13467 & n13477;
  assign n13479 = ~n13467 & ~n13477;
  assign n13480 = ~n13478 & ~n13479;
  assign n13481 = ~n13461 & n13480;
  assign n13482 = ~n13461 & ~n13481;
  assign n13483 = n13480 & ~n13481;
  assign n13484 = ~n13482 & ~n13483;
  assign n13485 = ~n13256 & ~n13260;
  assign n13486 = ~n13304 & ~n13307;
  assign n13487 = ~n13310 & ~n13313;
  assign n13488 = n13486 & n13487;
  assign n13489 = ~n13486 & ~n13487;
  assign n13490 = ~n13488 & ~n13489;
  assign n13491 = ~n13191 & ~n13206;
  assign n13492 = ~n13490 & n13491;
  assign n13493 = n13490 & ~n13491;
  assign n13494 = ~n13492 & ~n13493;
  assign n13495 = n2110 & n8854;
  assign n13496 = pi24  & pi59 ;
  assign n13497 = ~n13495 & n13496;
  assign n13498 = pi23  & pi60 ;
  assign n13499 = ~n13495 & n13498;
  assign n13500 = ~n13497 & ~n13499;
  assign n13501 = ~n13233 & ~n13500;
  assign n13502 = ~n13233 & ~n13501;
  assign n13503 = ~n13500 & ~n13501;
  assign n13504 = ~n13502 & ~n13503;
  assign n13505 = pi31  & pi52 ;
  assign n13506 = n7172 & n7354;
  assign n13507 = pi28  & pi55 ;
  assign n13508 = pi30  & pi53 ;
  assign n13509 = ~n13507 & ~n13508;
  assign n13510 = n13505 & ~n13506;
  assign n13511 = ~n13509 & n13510;
  assign n13512 = n13505 & ~n13511;
  assign n13513 = ~n13506 & ~n13511;
  assign n13514 = ~n13509 & n13513;
  assign n13515 = ~n13512 & ~n13514;
  assign n13516 = ~n13504 & ~n13515;
  assign n13517 = ~n13504 & ~n13516;
  assign n13518 = ~n13515 & ~n13516;
  assign n13519 = ~n13517 & ~n13518;
  assign n13520 = ~n13330 & ~n13334;
  assign n13521 = n13519 & n13520;
  assign n13522 = ~n13519 & ~n13520;
  assign n13523 = ~n13521 & ~n13522;
  assign n13524 = ~n13328 & ~n13336;
  assign n13525 = n13523 & ~n13524;
  assign n13526 = ~n13523 & n13524;
  assign n13527 = ~n13525 & ~n13526;
  assign n13528 = n13494 & n13527;
  assign n13529 = ~n13494 & ~n13527;
  assign n13530 = ~n13528 & ~n13529;
  assign n13531 = ~n13485 & n13530;
  assign n13532 = n13485 & ~n13530;
  assign n13533 = ~n13531 & ~n13532;
  assign n13534 = n13484 & n13533;
  assign n13535 = ~n13484 & ~n13533;
  assign n13536 = ~n13534 & ~n13535;
  assign n13537 = n13455 & ~n13536;
  assign n13538 = n13455 & ~n13537;
  assign n13539 = ~n13536 & ~n13537;
  assign n13540 = ~n13538 & ~n13539;
  assign n13541 = ~n13355 & ~n13540;
  assign n13542 = n13355 & n13540;
  assign n13543 = ~n13541 & ~n13542;
  assign n13544 = ~n13349 & ~n13352;
  assign n13545 = ~n13543 & n13544;
  assign n13546 = n13543 & ~n13544;
  assign po84  = ~n13545 & ~n13546;
  assign n13548 = ~n13453 & ~n13537;
  assign n13549 = ~n13532 & ~n13534;
  assign n13550 = ~n13495 & ~n13501;
  assign n13551 = n13437 & n13550;
  assign n13552 = ~n13437 & ~n13550;
  assign n13553 = ~n13551 & ~n13552;
  assign n13554 = pi26  & pi58 ;
  assign n13555 = n3567 & n9144;
  assign n13556 = pi31  & pi53 ;
  assign n13557 = pi32  & pi52 ;
  assign n13558 = ~n13556 & ~n13557;
  assign n13559 = n13554 & ~n13555;
  assign n13560 = ~n13558 & n13559;
  assign n13561 = n13554 & ~n13560;
  assign n13562 = ~n13555 & ~n13560;
  assign n13563 = ~n13558 & n13562;
  assign n13564 = ~n13561 & ~n13563;
  assign n13565 = n13553 & ~n13564;
  assign n13566 = n13553 & ~n13565;
  assign n13567 = ~n13564 & ~n13565;
  assign n13568 = ~n13566 & ~n13567;
  assign n13569 = ~n13516 & ~n13522;
  assign n13570 = n13568 & n13569;
  assign n13571 = ~n13568 & ~n13569;
  assign n13572 = ~n13570 & ~n13571;
  assign n13573 = ~n13489 & ~n13493;
  assign n13574 = ~n13572 & n13573;
  assign n13575 = n13572 & ~n13573;
  assign n13576 = ~n13574 & ~n13575;
  assign n13577 = ~n13525 & ~n13528;
  assign n13578 = ~n13576 & n13577;
  assign n13579 = n13576 & ~n13577;
  assign n13580 = ~n13578 & ~n13579;
  assign n13581 = pi22  & pi62 ;
  assign n13582 = pi23  & pi61 ;
  assign n13583 = ~n13581 & ~n13582;
  assign n13584 = n1806 & n9567;
  assign n13585 = pi21  & pi63 ;
  assign n13586 = ~n13583 & n13585;
  assign n13587 = ~n13584 & n13586;
  assign n13588 = ~n13584 & ~n13587;
  assign n13589 = ~n13583 & n13588;
  assign n13590 = n13585 & ~n13587;
  assign n13591 = ~n13589 & ~n13590;
  assign n13592 = pi33  & pi51 ;
  assign n13593 = n1789 & n8854;
  assign n13594 = pi24  & pi60 ;
  assign n13595 = pi25  & pi59 ;
  assign n13596 = ~n13594 & ~n13595;
  assign n13597 = n13592 & ~n13593;
  assign n13598 = ~n13596 & n13597;
  assign n13599 = n13592 & ~n13598;
  assign n13600 = ~n13593 & ~n13598;
  assign n13601 = ~n13596 & n13600;
  assign n13602 = ~n13599 & ~n13601;
  assign n13603 = ~n13591 & ~n13602;
  assign n13604 = ~n13591 & ~n13603;
  assign n13605 = ~n13602 & ~n13603;
  assign n13606 = ~n13604 & ~n13605;
  assign n13607 = pi34  & pi50 ;
  assign n13608 = n4691 & n8505;
  assign n13609 = pi35  & pi49 ;
  assign n13610 = pi36  & pi48 ;
  assign n13611 = ~n13609 & ~n13610;
  assign n13612 = n13607 & ~n13608;
  assign n13613 = ~n13611 & n13612;
  assign n13614 = n13607 & ~n13613;
  assign n13615 = ~n13608 & ~n13613;
  assign n13616 = ~n13611 & n13615;
  assign n13617 = ~n13614 & ~n13616;
  assign n13618 = ~n13606 & ~n13617;
  assign n13619 = ~n13606 & ~n13618;
  assign n13620 = ~n13617 & ~n13618;
  assign n13621 = ~n13619 & ~n13620;
  assign n13622 = pi29  & pi55 ;
  assign n13623 = pi38  & pi46 ;
  assign n13624 = ~n13622 & ~n13623;
  assign n13625 = n13622 & n13623;
  assign n13626 = pi28  & pi56 ;
  assign n13627 = ~n13624 & n13626;
  assign n13628 = ~n13625 & n13627;
  assign n13629 = ~n13625 & ~n13628;
  assign n13630 = ~n13624 & n13629;
  assign n13631 = n13626 & ~n13628;
  assign n13632 = ~n13630 & ~n13631;
  assign n13633 = pi39  & pi45 ;
  assign n13634 = n6012 & n6836;
  assign n13635 = pi40  & pi44 ;
  assign n13636 = ~n4490 & ~n13635;
  assign n13637 = n13633 & ~n13634;
  assign n13638 = ~n13636 & n13637;
  assign n13639 = n13633 & ~n13638;
  assign n13640 = ~n13634 & ~n13638;
  assign n13641 = ~n13636 & n13640;
  assign n13642 = ~n13639 & ~n13641;
  assign n13643 = ~n13632 & ~n13642;
  assign n13644 = ~n13632 & ~n13643;
  assign n13645 = ~n13642 & ~n13643;
  assign n13646 = ~n13644 & ~n13645;
  assign n13647 = pi37  & pi47 ;
  assign n13648 = pi30  & pi57 ;
  assign n13649 = n13060 & n13648;
  assign n13650 = pi27  & pi57 ;
  assign n13651 = pi30  & pi54 ;
  assign n13652 = ~n13650 & ~n13651;
  assign n13653 = n13647 & ~n13649;
  assign n13654 = ~n13652 & n13653;
  assign n13655 = n13647 & ~n13654;
  assign n13656 = ~n13649 & ~n13654;
  assign n13657 = ~n13652 & n13656;
  assign n13658 = ~n13655 & ~n13657;
  assign n13659 = ~n13646 & ~n13658;
  assign n13660 = ~n13646 & ~n13659;
  assign n13661 = ~n13658 & ~n13659;
  assign n13662 = ~n13660 & ~n13661;
  assign n13663 = ~n13621 & n13662;
  assign n13664 = n13621 & ~n13662;
  assign n13665 = ~n13663 & ~n13664;
  assign n13666 = n13392 & n13423;
  assign n13667 = ~n13392 & ~n13423;
  assign n13668 = ~n13666 & ~n13667;
  assign n13669 = n13411 & ~n13668;
  assign n13670 = ~n13411 & n13668;
  assign n13671 = ~n13669 & ~n13670;
  assign n13672 = ~n13463 & ~n13466;
  assign n13673 = ~n13469 & ~n13472;
  assign n13674 = n13672 & n13673;
  assign n13675 = ~n13672 & ~n13673;
  assign n13676 = ~n13674 & ~n13675;
  assign n13677 = n13671 & n13676;
  assign n13678 = ~n13671 & ~n13676;
  assign n13679 = ~n13677 & ~n13678;
  assign n13680 = ~n13665 & n13679;
  assign n13681 = ~n13665 & ~n13680;
  assign n13682 = n13679 & ~n13680;
  assign n13683 = ~n13681 & ~n13682;
  assign n13684 = n13580 & ~n13683;
  assign n13685 = ~n13580 & n13683;
  assign n13686 = ~n13684 & ~n13685;
  assign n13687 = n13549 & n13686;
  assign n13688 = n13549 & ~n13687;
  assign n13689 = n13686 & ~n13687;
  assign n13690 = ~n13688 & ~n13689;
  assign n13691 = ~n13447 & ~n13450;
  assign n13692 = ~n13458 & ~n13481;
  assign n13693 = n13691 & n13692;
  assign n13694 = ~n13691 & ~n13692;
  assign n13695 = ~n13693 & ~n13694;
  assign n13696 = ~n13401 & ~n13445;
  assign n13697 = ~n13476 & ~n13478;
  assign n13698 = ~n13696 & ~n13697;
  assign n13699 = ~n13696 & ~n13698;
  assign n13700 = ~n13697 & ~n13698;
  assign n13701 = ~n13699 & ~n13700;
  assign n13702 = n13363 & n13377;
  assign n13703 = ~n13363 & ~n13377;
  assign n13704 = ~n13702 & ~n13703;
  assign n13705 = n13513 & ~n13704;
  assign n13706 = ~n13513 & n13704;
  assign n13707 = ~n13705 & ~n13706;
  assign n13708 = ~n13426 & ~n13440;
  assign n13709 = ~n13380 & ~n13395;
  assign n13710 = n13708 & n13709;
  assign n13711 = ~n13708 & ~n13709;
  assign n13712 = ~n13710 & ~n13711;
  assign n13713 = n13707 & n13712;
  assign n13714 = ~n13707 & ~n13712;
  assign n13715 = ~n13713 & ~n13714;
  assign n13716 = ~n13701 & n13715;
  assign n13717 = ~n13701 & ~n13716;
  assign n13718 = n13715 & ~n13716;
  assign n13719 = ~n13717 & ~n13718;
  assign n13720 = n13695 & ~n13719;
  assign n13721 = ~n13695 & n13719;
  assign n13722 = ~n13720 & ~n13721;
  assign n13723 = ~n13690 & n13722;
  assign n13724 = ~n13690 & ~n13723;
  assign n13725 = n13722 & ~n13723;
  assign n13726 = ~n13724 & ~n13725;
  assign n13727 = ~n13548 & ~n13726;
  assign n13728 = n13548 & n13726;
  assign n13729 = ~n13727 & ~n13728;
  assign n13730 = ~n13541 & ~n13546;
  assign n13731 = n13729 & ~n13730;
  assign n13732 = ~n13729 & n13730;
  assign po85  = ~n13731 & ~n13732;
  assign n13734 = ~n13687 & ~n13723;
  assign n13735 = ~n13694 & ~n13720;
  assign n13736 = pi22  & pi63 ;
  assign n13737 = pi28  & pi57 ;
  assign n13738 = ~n13736 & ~n13737;
  assign n13739 = n13736 & n13737;
  assign n13740 = pi35  & pi50 ;
  assign n13741 = ~n13738 & n13740;
  assign n13742 = ~n13739 & n13741;
  assign n13743 = ~n13739 & ~n13742;
  assign n13744 = ~n13738 & n13743;
  assign n13745 = n13740 & ~n13742;
  assign n13746 = ~n13744 & ~n13745;
  assign n13747 = pi32  & pi53 ;
  assign n13748 = n3900 & n10319;
  assign n13749 = pi33  & pi52 ;
  assign n13750 = pi34  & pi51 ;
  assign n13751 = ~n13749 & ~n13750;
  assign n13752 = n13747 & ~n13748;
  assign n13753 = ~n13751 & n13752;
  assign n13754 = n13747 & ~n13753;
  assign n13755 = ~n13748 & ~n13753;
  assign n13756 = ~n13751 & n13755;
  assign n13757 = ~n13754 & ~n13756;
  assign n13758 = ~n13746 & ~n13757;
  assign n13759 = ~n13746 & ~n13758;
  assign n13760 = ~n13757 & ~n13758;
  assign n13761 = ~n13759 & ~n13760;
  assign n13762 = pi39  & pi46 ;
  assign n13763 = n5318 & n6012;
  assign n13764 = pi40  & pi45 ;
  assign n13765 = pi41  & pi44 ;
  assign n13766 = ~n13764 & ~n13765;
  assign n13767 = n13762 & ~n13763;
  assign n13768 = ~n13766 & n13767;
  assign n13769 = n13762 & ~n13768;
  assign n13770 = ~n13763 & ~n13768;
  assign n13771 = ~n13766 & n13770;
  assign n13772 = ~n13769 & ~n13771;
  assign n13773 = ~n13761 & ~n13772;
  assign n13774 = ~n13761 & ~n13773;
  assign n13775 = ~n13772 & ~n13773;
  assign n13776 = ~n13774 & ~n13775;
  assign n13777 = pi43  & pi62 ;
  assign n13778 = pi23  & n13777;
  assign n13779 = n6458 & ~n13778;
  assign n13780 = ~n13778 & ~n13779;
  assign n13781 = pi23  & pi62 ;
  assign n13782 = ~pi43  & ~n13781;
  assign n13783 = n13780 & ~n13782;
  assign n13784 = n6458 & ~n13779;
  assign n13785 = ~n13783 & ~n13784;
  assign n13786 = pi36  & pi49 ;
  assign n13787 = n5055 & n5823;
  assign n13788 = pi37  & pi48 ;
  assign n13789 = pi38  & pi47 ;
  assign n13790 = ~n13788 & ~n13789;
  assign n13791 = n13786 & ~n13787;
  assign n13792 = ~n13790 & n13791;
  assign n13793 = n13786 & ~n13792;
  assign n13794 = ~n13787 & ~n13792;
  assign n13795 = ~n13790 & n13794;
  assign n13796 = ~n13793 & ~n13795;
  assign n13797 = ~n13785 & ~n13796;
  assign n13798 = ~n13785 & ~n13797;
  assign n13799 = ~n13796 & ~n13797;
  assign n13800 = ~n13798 & ~n13799;
  assign n13801 = pi29  & pi56 ;
  assign n13802 = n2680 & n9891;
  assign n13803 = pi30  & pi55 ;
  assign n13804 = pi31  & pi54 ;
  assign n13805 = ~n13803 & ~n13804;
  assign n13806 = n13801 & ~n13802;
  assign n13807 = ~n13805 & n13806;
  assign n13808 = n13801 & ~n13807;
  assign n13809 = ~n13802 & ~n13807;
  assign n13810 = ~n13805 & n13809;
  assign n13811 = ~n13808 & ~n13810;
  assign n13812 = ~n13800 & ~n13811;
  assign n13813 = ~n13800 & ~n13812;
  assign n13814 = ~n13811 & ~n13812;
  assign n13815 = ~n13813 & ~n13814;
  assign n13816 = ~n13776 & n13815;
  assign n13817 = n13776 & ~n13815;
  assign n13818 = ~n13816 & ~n13817;
  assign n13819 = ~n13711 & ~n13713;
  assign n13820 = n13818 & n13819;
  assign n13821 = ~n13818 & ~n13819;
  assign n13822 = ~n13820 & ~n13821;
  assign n13823 = ~n13675 & ~n13677;
  assign n13824 = pi24  & pi61 ;
  assign n13825 = ~n13640 & n13824;
  assign n13826 = n13640 & ~n13824;
  assign n13827 = ~n13825 & ~n13826;
  assign n13828 = n13629 & ~n13827;
  assign n13829 = ~n13629 & n13827;
  assign n13830 = ~n13828 & ~n13829;
  assign n13831 = n13562 & n13656;
  assign n13832 = ~n13562 & ~n13656;
  assign n13833 = ~n13831 & ~n13832;
  assign n13834 = pi25  & pi60 ;
  assign n13835 = n2646 & n9402;
  assign n13836 = pi26  & pi59 ;
  assign n13837 = pi27  & pi58 ;
  assign n13838 = ~n13836 & ~n13837;
  assign n13839 = n13834 & ~n13835;
  assign n13840 = ~n13838 & n13839;
  assign n13841 = n13834 & ~n13840;
  assign n13842 = ~n13835 & ~n13840;
  assign n13843 = ~n13838 & n13842;
  assign n13844 = ~n13841 & ~n13843;
  assign n13845 = n13833 & ~n13844;
  assign n13846 = n13833 & ~n13845;
  assign n13847 = ~n13844 & ~n13845;
  assign n13848 = ~n13846 & ~n13847;
  assign n13849 = n13830 & ~n13848;
  assign n13850 = ~n13830 & n13848;
  assign n13851 = ~n13849 & ~n13850;
  assign n13852 = ~n13823 & n13851;
  assign n13853 = ~n13823 & ~n13852;
  assign n13854 = ~n13849 & ~n13852;
  assign n13855 = ~n13850 & n13854;
  assign n13856 = ~n13853 & ~n13855;
  assign n13857 = n13588 & n13615;
  assign n13858 = ~n13588 & ~n13615;
  assign n13859 = ~n13857 & ~n13858;
  assign n13860 = n13600 & ~n13859;
  assign n13861 = ~n13600 & n13859;
  assign n13862 = ~n13860 & ~n13861;
  assign n13863 = ~n13643 & ~n13659;
  assign n13864 = ~n13603 & ~n13618;
  assign n13865 = n13863 & n13864;
  assign n13866 = ~n13863 & ~n13864;
  assign n13867 = ~n13865 & ~n13866;
  assign n13868 = n13862 & n13867;
  assign n13869 = ~n13862 & ~n13867;
  assign n13870 = ~n13868 & ~n13869;
  assign n13871 = ~n13856 & n13870;
  assign n13872 = ~n13856 & ~n13871;
  assign n13873 = n13870 & ~n13871;
  assign n13874 = ~n13872 & ~n13873;
  assign n13875 = n13822 & ~n13874;
  assign n13876 = n13822 & ~n13875;
  assign n13877 = ~n13874 & ~n13875;
  assign n13878 = ~n13876 & ~n13877;
  assign n13879 = ~n13735 & ~n13878;
  assign n13880 = ~n13735 & ~n13879;
  assign n13881 = ~n13878 & ~n13879;
  assign n13882 = ~n13880 & ~n13881;
  assign n13883 = ~n13698 & ~n13716;
  assign n13884 = ~n13667 & ~n13670;
  assign n13885 = ~n13703 & ~n13706;
  assign n13886 = n13884 & n13885;
  assign n13887 = ~n13884 & ~n13885;
  assign n13888 = ~n13886 & ~n13887;
  assign n13889 = ~n13552 & ~n13565;
  assign n13890 = ~n13888 & n13889;
  assign n13891 = n13888 & ~n13889;
  assign n13892 = ~n13890 & ~n13891;
  assign n13893 = ~n13571 & ~n13575;
  assign n13894 = ~n13892 & n13893;
  assign n13895 = n13892 & ~n13893;
  assign n13896 = ~n13894 & ~n13895;
  assign n13897 = ~n13621 & ~n13662;
  assign n13898 = ~n13680 & ~n13897;
  assign n13899 = n13896 & ~n13898;
  assign n13900 = ~n13896 & n13898;
  assign n13901 = ~n13899 & ~n13900;
  assign n13902 = n13883 & ~n13901;
  assign n13903 = ~n13883 & n13901;
  assign n13904 = ~n13902 & ~n13903;
  assign n13905 = ~n13579 & ~n13684;
  assign n13906 = n13904 & ~n13905;
  assign n13907 = ~n13904 & n13905;
  assign n13908 = ~n13906 & ~n13907;
  assign n13909 = ~n13882 & ~n13908;
  assign n13910 = n13882 & n13908;
  assign n13911 = ~n13909 & ~n13910;
  assign n13912 = ~n13734 & ~n13911;
  assign n13913 = n13734 & n13911;
  assign n13914 = ~n13912 & ~n13913;
  assign n13915 = ~n13727 & ~n13731;
  assign n13916 = ~n13914 & ~n13915;
  assign n13917 = n13914 & n13915;
  assign po86  = n13916 | n13917;
  assign n13919 = ~n13913 & ~n13915;
  assign n13920 = ~n13912 & ~n13919;
  assign n13921 = ~n13882 & n13908;
  assign n13922 = ~n13879 & ~n13921;
  assign n13923 = ~n13903 & ~n13906;
  assign n13924 = ~n13832 & ~n13845;
  assign n13925 = ~n13758 & ~n13773;
  assign n13926 = n13924 & n13925;
  assign n13927 = ~n13924 & ~n13925;
  assign n13928 = ~n13926 & ~n13927;
  assign n13929 = ~n13797 & ~n13812;
  assign n13930 = ~n13928 & n13929;
  assign n13931 = n13928 & ~n13929;
  assign n13932 = ~n13930 & ~n13931;
  assign n13933 = ~n13887 & ~n13891;
  assign n13934 = n13770 & n13809;
  assign n13935 = ~n13770 & ~n13809;
  assign n13936 = ~n13934 & ~n13935;
  assign n13937 = n13794 & ~n13936;
  assign n13938 = ~n13794 & n13936;
  assign n13939 = ~n13937 & ~n13938;
  assign n13940 = n13755 & n13842;
  assign n13941 = ~n13755 & ~n13842;
  assign n13942 = ~n13940 & ~n13941;
  assign n13943 = n13743 & ~n13942;
  assign n13944 = ~n13743 & n13942;
  assign n13945 = ~n13943 & ~n13944;
  assign n13946 = n13939 & n13945;
  assign n13947 = ~n13939 & ~n13945;
  assign n13948 = ~n13946 & ~n13947;
  assign n13949 = ~n13933 & n13948;
  assign n13950 = n13933 & ~n13948;
  assign n13951 = ~n13949 & ~n13950;
  assign n13952 = n13932 & n13951;
  assign n13953 = ~n13932 & ~n13951;
  assign n13954 = ~n13952 & ~n13953;
  assign n13955 = ~n13866 & ~n13868;
  assign n13956 = pi36  & pi50 ;
  assign n13957 = pi37  & pi49 ;
  assign n13958 = ~n13956 & ~n13957;
  assign n13959 = n4500 & n5889;
  assign n13960 = pi23  & pi63 ;
  assign n13961 = ~n13958 & n13960;
  assign n13962 = ~n13959 & n13961;
  assign n13963 = ~n13959 & ~n13962;
  assign n13964 = ~n13958 & n13963;
  assign n13965 = n13960 & ~n13962;
  assign n13966 = ~n13964 & ~n13965;
  assign n13967 = pi33  & pi53 ;
  assign n13968 = n3106 & n10319;
  assign n13969 = pi34  & pi52 ;
  assign n13970 = pi35  & pi51 ;
  assign n13971 = ~n13969 & ~n13970;
  assign n13972 = n13967 & ~n13968;
  assign n13973 = ~n13971 & n13972;
  assign n13974 = n13967 & ~n13973;
  assign n13975 = ~n13968 & ~n13973;
  assign n13976 = ~n13971 & n13975;
  assign n13977 = ~n13974 & ~n13976;
  assign n13978 = ~n13966 & ~n13977;
  assign n13979 = ~n13966 & ~n13978;
  assign n13980 = ~n13977 & ~n13978;
  assign n13981 = ~n13979 & ~n13980;
  assign n13982 = n7865 & n13270;
  assign n13983 = pi29  & pi57 ;
  assign n13984 = pi31  & pi55 ;
  assign n13985 = ~n13983 & ~n13984;
  assign n13986 = n6474 & ~n13982;
  assign n13987 = ~n13985 & n13986;
  assign n13988 = n6474 & ~n13987;
  assign n13989 = ~n13982 & ~n13987;
  assign n13990 = ~n13985 & n13989;
  assign n13991 = ~n13988 & ~n13990;
  assign n13992 = ~n13981 & ~n13991;
  assign n13993 = ~n13981 & ~n13992;
  assign n13994 = ~n13991 & ~n13992;
  assign n13995 = ~n13993 & ~n13994;
  assign n13996 = pi27  & pi59 ;
  assign n13997 = pi28  & pi58 ;
  assign n13998 = ~n13996 & ~n13997;
  assign n13999 = n2191 & n9402;
  assign n14000 = pi26  & pi60 ;
  assign n14001 = ~n13998 & n14000;
  assign n14002 = ~n13999 & n14001;
  assign n14003 = ~n13999 & ~n14002;
  assign n14004 = ~n13998 & n14003;
  assign n14005 = n14000 & ~n14002;
  assign n14006 = ~n14004 & ~n14005;
  assign n14007 = pi41  & pi45 ;
  assign n14008 = pi32  & pi54 ;
  assign n14009 = n4329 & n14008;
  assign n14010 = ~n4329 & ~n14008;
  assign n14011 = n14007 & ~n14009;
  assign n14012 = ~n14010 & n14011;
  assign n14013 = n14007 & ~n14012;
  assign n14014 = ~n14009 & ~n14012;
  assign n14015 = ~n14010 & n14014;
  assign n14016 = ~n14013 & ~n14015;
  assign n14017 = ~n14006 & ~n14016;
  assign n14018 = ~n14006 & ~n14017;
  assign n14019 = ~n14016 & ~n14017;
  assign n14020 = ~n14018 & ~n14019;
  assign n14021 = pi30  & pi56 ;
  assign n14022 = n5277 & n5548;
  assign n14023 = pi40  & pi46 ;
  assign n14024 = pi39  & pi47 ;
  assign n14025 = ~n14023 & ~n14024;
  assign n14026 = n14021 & ~n14022;
  assign n14027 = ~n14025 & n14026;
  assign n14028 = n14021 & ~n14027;
  assign n14029 = ~n14022 & ~n14027;
  assign n14030 = ~n14025 & n14029;
  assign n14031 = ~n14028 & ~n14030;
  assign n14032 = ~n14020 & ~n14031;
  assign n14033 = ~n14020 & ~n14032;
  assign n14034 = ~n14031 & ~n14032;
  assign n14035 = ~n14033 & ~n14034;
  assign n14036 = n13995 & n14035;
  assign n14037 = ~n13995 & ~n14035;
  assign n14038 = ~n14036 & ~n14037;
  assign n14039 = ~n13955 & n14038;
  assign n14040 = n13955 & ~n14038;
  assign n14041 = ~n14039 & ~n14040;
  assign n14042 = n13954 & n14041;
  assign n14043 = ~n13954 & ~n14041;
  assign n14044 = ~n14042 & ~n14043;
  assign n14045 = ~n13923 & n14044;
  assign n14046 = ~n13923 & ~n14045;
  assign n14047 = n14044 & ~n14045;
  assign n14048 = ~n14046 & ~n14047;
  assign n14049 = ~n13871 & ~n13875;
  assign n14050 = ~n13895 & ~n13899;
  assign n14051 = n14049 & n14050;
  assign n14052 = ~n14049 & ~n14050;
  assign n14053 = ~n14051 & ~n14052;
  assign n14054 = n1789 & n9567;
  assign n14055 = pi25  & pi61 ;
  assign n14056 = ~n14054 & n14055;
  assign n14057 = pi24  & pi62 ;
  assign n14058 = ~n14054 & n14057;
  assign n14059 = ~n14056 & ~n14058;
  assign n14060 = ~n13780 & ~n14059;
  assign n14061 = ~n13780 & ~n14060;
  assign n14062 = ~n14059 & ~n14060;
  assign n14063 = ~n14061 & ~n14062;
  assign n14064 = ~n13825 & ~n13829;
  assign n14065 = n14063 & n14064;
  assign n14066 = ~n14063 & ~n14064;
  assign n14067 = ~n14065 & ~n14066;
  assign n14068 = ~n13858 & ~n13861;
  assign n14069 = ~n14067 & n14068;
  assign n14070 = n14067 & ~n14068;
  assign n14071 = ~n14069 & ~n14070;
  assign n14072 = ~n13854 & n14071;
  assign n14073 = n13854 & ~n14071;
  assign n14074 = ~n14072 & ~n14073;
  assign n14075 = ~n13776 & ~n13815;
  assign n14076 = ~n13821 & ~n14075;
  assign n14077 = n14074 & ~n14076;
  assign n14078 = ~n14074 & n14076;
  assign n14079 = ~n14077 & ~n14078;
  assign n14080 = n14053 & n14079;
  assign n14081 = ~n14053 & ~n14079;
  assign n14082 = ~n14080 & ~n14081;
  assign n14083 = ~n14048 & n14082;
  assign n14084 = n14048 & ~n14082;
  assign n14085 = ~n14083 & ~n14084;
  assign n14086 = n13922 & ~n14085;
  assign n14087 = ~n13922 & n14085;
  assign n14088 = ~n14086 & ~n14087;
  assign n14089 = n13920 & ~n14088;
  assign n14090 = ~n13920 & ~n14086;
  assign n14091 = ~n14087 & n14090;
  assign po87  = ~n14089 & ~n14091;
  assign n14093 = ~n14087 & ~n14090;
  assign n14094 = ~n14045 & ~n14083;
  assign n14095 = ~n14037 & ~n14039;
  assign n14096 = ~n13935 & ~n13938;
  assign n14097 = ~n13978 & ~n13992;
  assign n14098 = n14096 & n14097;
  assign n14099 = ~n14096 & ~n14097;
  assign n14100 = ~n14098 & ~n14099;
  assign n14101 = ~n14017 & ~n14032;
  assign n14102 = ~n14100 & n14101;
  assign n14103 = n14100 & ~n14101;
  assign n14104 = ~n14102 & ~n14103;
  assign n14105 = ~n14095 & n14104;
  assign n14106 = n14095 & ~n14104;
  assign n14107 = ~n14105 & ~n14106;
  assign n14108 = ~n14072 & ~n14077;
  assign n14109 = ~n14107 & n14108;
  assign n14110 = n14107 & ~n14108;
  assign n14111 = ~n14109 & ~n14110;
  assign n14112 = ~n14052 & ~n14080;
  assign n14113 = ~n14111 & n14112;
  assign n14114 = n14111 & ~n14112;
  assign n14115 = ~n14113 & ~n14114;
  assign n14116 = ~n13952 & ~n14042;
  assign n14117 = pi44  & pi62 ;
  assign n14118 = pi25  & n14117;
  assign n14119 = n6836 & ~n14118;
  assign n14120 = ~n14118 & ~n14119;
  assign n14121 = pi25  & pi62 ;
  assign n14122 = ~pi44  & ~n14121;
  assign n14123 = n14120 & ~n14122;
  assign n14124 = n6836 & ~n14119;
  assign n14125 = ~n14123 & ~n14124;
  assign n14126 = pi40  & pi47 ;
  assign n14127 = n6911 & n9026;
  assign n14128 = pi31  & pi56 ;
  assign n14129 = pi33  & pi54 ;
  assign n14130 = ~n14128 & ~n14129;
  assign n14131 = n14126 & ~n14127;
  assign n14132 = ~n14130 & n14131;
  assign n14133 = n14126 & ~n14132;
  assign n14134 = ~n14127 & ~n14132;
  assign n14135 = ~n14130 & n14134;
  assign n14136 = ~n14133 & ~n14135;
  assign n14137 = ~n14125 & ~n14136;
  assign n14138 = ~n14125 & ~n14137;
  assign n14139 = ~n14136 & ~n14137;
  assign n14140 = ~n14138 & ~n14139;
  assign n14141 = ~n13941 & ~n13944;
  assign n14142 = n14140 & n14141;
  assign n14143 = ~n14140 & ~n14141;
  assign n14144 = ~n14142 & ~n14143;
  assign n14145 = pi26  & pi61 ;
  assign n14146 = pi27  & pi60 ;
  assign n14147 = ~n14145 & ~n14146;
  assign n14148 = n2646 & n9054;
  assign n14149 = pi24  & pi63 ;
  assign n14150 = ~n14147 & n14149;
  assign n14151 = ~n14148 & n14150;
  assign n14152 = ~n14148 & ~n14151;
  assign n14153 = ~n14147 & n14152;
  assign n14154 = n14149 & ~n14151;
  assign n14155 = ~n14153 & ~n14154;
  assign n14156 = pi37  & pi50 ;
  assign n14157 = n4736 & n8505;
  assign n14158 = pi38  & pi49 ;
  assign n14159 = pi39  & pi48 ;
  assign n14160 = ~n14158 & ~n14159;
  assign n14161 = n14156 & ~n14157;
  assign n14162 = ~n14160 & n14161;
  assign n14163 = n14156 & ~n14162;
  assign n14164 = ~n14157 & ~n14162;
  assign n14165 = ~n14160 & n14164;
  assign n14166 = ~n14163 & ~n14165;
  assign n14167 = ~n14155 & ~n14166;
  assign n14168 = ~n14155 & ~n14167;
  assign n14169 = ~n14166 & ~n14167;
  assign n14170 = ~n14168 & ~n14169;
  assign n14171 = pi32  & pi55 ;
  assign n14172 = n5235 & n7513;
  assign n14173 = pi41  & pi46 ;
  assign n14174 = pi42  & pi45 ;
  assign n14175 = ~n14173 & ~n14174;
  assign n14176 = n14171 & ~n14172;
  assign n14177 = ~n14175 & n14176;
  assign n14178 = n14171 & ~n14177;
  assign n14179 = ~n14172 & ~n14177;
  assign n14180 = ~n14175 & n14179;
  assign n14181 = ~n14178 & ~n14180;
  assign n14182 = ~n14170 & ~n14181;
  assign n14183 = ~n14170 & ~n14182;
  assign n14184 = ~n14181 & ~n14182;
  assign n14185 = ~n14183 & ~n14184;
  assign n14186 = ~n14144 & n14185;
  assign n14187 = n14144 & ~n14185;
  assign n14188 = ~n14186 & ~n14187;
  assign n14189 = pi28  & pi59 ;
  assign n14190 = pi34  & pi53 ;
  assign n14191 = n13648 & n14190;
  assign n14192 = ~n13648 & ~n14190;
  assign n14193 = n14189 & ~n14191;
  assign n14194 = ~n14192 & n14193;
  assign n14195 = n14189 & ~n14194;
  assign n14196 = ~n14191 & ~n14194;
  assign n14197 = ~n14192 & n14196;
  assign n14198 = ~n14195 & ~n14197;
  assign n14199 = ~n14054 & ~n14060;
  assign n14200 = ~n14198 & n14199;
  assign n14201 = n14198 & ~n14199;
  assign n14202 = ~n14200 & ~n14201;
  assign n14203 = pi35  & pi52 ;
  assign n14204 = pi29  & pi58 ;
  assign n14205 = pi36  & pi51 ;
  assign n14206 = n14204 & n14205;
  assign n14207 = ~n14204 & ~n14205;
  assign n14208 = n14203 & ~n14206;
  assign n14209 = ~n14207 & n14208;
  assign n14210 = n14203 & ~n14209;
  assign n14211 = ~n14206 & ~n14209;
  assign n14212 = ~n14207 & n14211;
  assign n14213 = ~n14210 & ~n14212;
  assign n14214 = ~n14202 & ~n14213;
  assign n14215 = n14202 & n14213;
  assign n14216 = ~n14214 & ~n14215;
  assign n14217 = n14188 & n14216;
  assign n14218 = ~n14188 & ~n14216;
  assign n14219 = ~n14217 & ~n14218;
  assign n14220 = ~n14116 & n14219;
  assign n14221 = n14116 & ~n14219;
  assign n14222 = ~n14220 & ~n14221;
  assign n14223 = ~n13946 & ~n13949;
  assign n14224 = ~n13927 & ~n13931;
  assign n14225 = n14223 & n14224;
  assign n14226 = ~n14223 & ~n14224;
  assign n14227 = ~n14225 & ~n14226;
  assign n14228 = ~n14066 & ~n14070;
  assign n14229 = n14014 & n14029;
  assign n14230 = ~n14014 & ~n14029;
  assign n14231 = ~n14229 & ~n14230;
  assign n14232 = n13989 & ~n14231;
  assign n14233 = ~n13989 & n14231;
  assign n14234 = ~n14232 & ~n14233;
  assign n14235 = n13975 & n14003;
  assign n14236 = ~n13975 & ~n14003;
  assign n14237 = ~n14235 & ~n14236;
  assign n14238 = n13963 & ~n14237;
  assign n14239 = ~n13963 & n14237;
  assign n14240 = ~n14238 & ~n14239;
  assign n14241 = ~n14234 & ~n14240;
  assign n14242 = n14234 & n14240;
  assign n14243 = ~n14241 & ~n14242;
  assign n14244 = ~n14228 & n14243;
  assign n14245 = n14228 & ~n14243;
  assign n14246 = ~n14244 & ~n14245;
  assign n14247 = n14227 & n14246;
  assign n14248 = ~n14227 & ~n14246;
  assign n14249 = ~n14247 & ~n14248;
  assign n14250 = n14222 & n14249;
  assign n14251 = n14222 & ~n14250;
  assign n14252 = n14249 & ~n14250;
  assign n14253 = ~n14251 & ~n14252;
  assign n14254 = ~n14115 & n14253;
  assign n14255 = n14115 & ~n14253;
  assign n14256 = ~n14254 & ~n14255;
  assign n14257 = n14094 & ~n14256;
  assign n14258 = ~n14094 & n14256;
  assign n14259 = ~n14257 & ~n14258;
  assign n14260 = ~n14093 & ~n14259;
  assign n14261 = n14093 & n14259;
  assign po88  = n14260 | n14261;
  assign n14263 = ~n14114 & ~n14255;
  assign n14264 = ~n14220 & ~n14250;
  assign n14265 = ~n14226 & ~n14247;
  assign n14266 = ~n14236 & ~n14239;
  assign n14267 = ~n14198 & ~n14199;
  assign n14268 = ~n14214 & ~n14267;
  assign n14269 = n14266 & n14268;
  assign n14270 = ~n14266 & ~n14268;
  assign n14271 = ~n14269 & ~n14270;
  assign n14272 = ~n14167 & ~n14182;
  assign n14273 = ~n14271 & n14272;
  assign n14274 = n14271 & ~n14272;
  assign n14275 = ~n14273 & ~n14274;
  assign n14276 = ~n14187 & ~n14217;
  assign n14277 = n14275 & ~n14276;
  assign n14278 = ~n14275 & n14276;
  assign n14279 = ~n14277 & ~n14278;
  assign n14280 = ~n14265 & n14279;
  assign n14281 = n14265 & ~n14279;
  assign n14282 = ~n14280 & ~n14281;
  assign n14283 = ~n14264 & n14282;
  assign n14284 = n14264 & ~n14282;
  assign n14285 = ~n14283 & ~n14284;
  assign n14286 = ~n14105 & ~n14110;
  assign n14287 = pi27  & pi61 ;
  assign n14288 = pi28  & pi60 ;
  assign n14289 = ~n14287 & ~n14288;
  assign n14290 = n2191 & n9054;
  assign n14291 = pi26  & pi62 ;
  assign n14292 = ~n14289 & n14291;
  assign n14293 = ~n14290 & n14292;
  assign n14294 = ~n14290 & ~n14293;
  assign n14295 = ~n14289 & n14294;
  assign n14296 = n14291 & ~n14293;
  assign n14297 = ~n14295 & ~n14296;
  assign n14298 = pi31  & pi57 ;
  assign n14299 = n5235 & n5277;
  assign n14300 = pi42  & pi46 ;
  assign n14301 = pi41  & pi47 ;
  assign n14302 = ~n14300 & ~n14301;
  assign n14303 = n14298 & ~n14299;
  assign n14304 = ~n14302 & n14303;
  assign n14305 = n14298 & ~n14304;
  assign n14306 = ~n14299 & ~n14304;
  assign n14307 = ~n14302 & n14306;
  assign n14308 = ~n14305 & ~n14307;
  assign n14309 = ~n14297 & ~n14308;
  assign n14310 = ~n14297 & ~n14309;
  assign n14311 = ~n14308 & ~n14309;
  assign n14312 = ~n14310 & ~n14311;
  assign n14313 = pi35  & pi53 ;
  assign n14314 = n4500 & n10319;
  assign n14315 = pi37  & pi51 ;
  assign n14316 = pi36  & pi52 ;
  assign n14317 = ~n14315 & ~n14316;
  assign n14318 = n14313 & ~n14314;
  assign n14319 = ~n14317 & n14318;
  assign n14320 = n14313 & ~n14319;
  assign n14321 = ~n14314 & ~n14319;
  assign n14322 = ~n14317 & n14321;
  assign n14323 = ~n14320 & ~n14322;
  assign n14324 = ~n14312 & ~n14323;
  assign n14325 = ~n14312 & ~n14324;
  assign n14326 = ~n14323 & ~n14324;
  assign n14327 = ~n14325 & ~n14326;
  assign n14328 = pi38  & pi50 ;
  assign n14329 = pi39  & pi49 ;
  assign n14330 = ~n14328 & ~n14329;
  assign n14331 = n4736 & n5889;
  assign n14332 = pi29  & pi59 ;
  assign n14333 = ~n14330 & n14332;
  assign n14334 = ~n14331 & n14333;
  assign n14335 = ~n14331 & ~n14334;
  assign n14336 = ~n14330 & n14335;
  assign n14337 = n14332 & ~n14334;
  assign n14338 = ~n14336 & ~n14337;
  assign n14339 = pi40  & pi48 ;
  assign n14340 = n2332 & n12970;
  assign n14341 = pi30  & pi58 ;
  assign n14342 = pi32  & pi56 ;
  assign n14343 = ~n14341 & ~n14342;
  assign n14344 = n14339 & ~n14340;
  assign n14345 = ~n14343 & n14344;
  assign n14346 = n14339 & ~n14345;
  assign n14347 = ~n14340 & ~n14345;
  assign n14348 = ~n14343 & n14347;
  assign n14349 = ~n14346 & ~n14348;
  assign n14350 = ~n14338 & ~n14349;
  assign n14351 = ~n14338 & ~n14350;
  assign n14352 = ~n14349 & ~n14350;
  assign n14353 = ~n14351 & ~n14352;
  assign n14354 = ~n14230 & ~n14233;
  assign n14355 = n14353 & n14354;
  assign n14356 = ~n14353 & ~n14354;
  assign n14357 = ~n14355 & ~n14356;
  assign n14358 = pi25  & pi63 ;
  assign n14359 = ~n14120 & n14358;
  assign n14360 = n14120 & ~n14358;
  assign n14361 = ~n14359 & ~n14360;
  assign n14362 = n14179 & ~n14361;
  assign n14363 = ~n14179 & n14361;
  assign n14364 = ~n14362 & ~n14363;
  assign n14365 = n14357 & n14364;
  assign n14366 = ~n14357 & ~n14364;
  assign n14367 = ~n14365 & ~n14366;
  assign n14368 = ~n14327 & n14367;
  assign n14369 = ~n14327 & ~n14368;
  assign n14370 = n14367 & ~n14368;
  assign n14371 = ~n14369 & ~n14370;
  assign n14372 = ~n14286 & ~n14371;
  assign n14373 = ~n14286 & ~n14372;
  assign n14374 = ~n14371 & ~n14372;
  assign n14375 = ~n14373 & ~n14374;
  assign n14376 = ~n14242 & ~n14244;
  assign n14377 = ~n14099 & ~n14103;
  assign n14378 = n14376 & n14377;
  assign n14379 = ~n14376 & ~n14377;
  assign n14380 = ~n14378 & ~n14379;
  assign n14381 = n14152 & n14196;
  assign n14382 = ~n14152 & ~n14196;
  assign n14383 = ~n14381 & ~n14382;
  assign n14384 = n14164 & ~n14383;
  assign n14385 = ~n14164 & n14383;
  assign n14386 = ~n14384 & ~n14385;
  assign n14387 = n14134 & n14211;
  assign n14388 = ~n14134 & ~n14211;
  assign n14389 = ~n14387 & ~n14388;
  assign n14390 = pi43  & pi45 ;
  assign n14391 = n3900 & n9891;
  assign n14392 = pi33  & pi55 ;
  assign n14393 = pi34  & pi54 ;
  assign n14394 = ~n14392 & ~n14393;
  assign n14395 = n14390 & ~n14391;
  assign n14396 = ~n14394 & n14395;
  assign n14397 = n14390 & ~n14396;
  assign n14398 = ~n14391 & ~n14396;
  assign n14399 = ~n14394 & n14398;
  assign n14400 = ~n14397 & ~n14399;
  assign n14401 = n14389 & ~n14400;
  assign n14402 = n14389 & ~n14401;
  assign n14403 = ~n14400 & ~n14401;
  assign n14404 = ~n14402 & ~n14403;
  assign n14405 = ~n14137 & ~n14143;
  assign n14406 = n14404 & n14405;
  assign n14407 = ~n14404 & ~n14405;
  assign n14408 = ~n14406 & ~n14407;
  assign n14409 = n14386 & n14408;
  assign n14410 = ~n14386 & ~n14408;
  assign n14411 = ~n14409 & ~n14410;
  assign n14412 = n14380 & n14411;
  assign n14413 = ~n14380 & ~n14411;
  assign n14414 = ~n14412 & ~n14413;
  assign n14415 = ~n14375 & ~n14414;
  assign n14416 = n14375 & n14414;
  assign n14417 = ~n14415 & ~n14416;
  assign n14418 = n14285 & ~n14417;
  assign n14419 = n14285 & ~n14418;
  assign n14420 = ~n14417 & ~n14418;
  assign n14421 = ~n14419 & ~n14420;
  assign n14422 = n14263 & n14421;
  assign n14423 = ~n14263 & ~n14421;
  assign n14424 = ~n14422 & ~n14423;
  assign n14425 = ~n14093 & ~n14257;
  assign n14426 = ~n14258 & ~n14425;
  assign n14427 = ~n14424 & n14426;
  assign n14428 = n14424 & ~n14426;
  assign po89  = ~n14427 & ~n14428;
  assign n14430 = ~n14283 & ~n14418;
  assign n14431 = ~n14277 & ~n14280;
  assign n14432 = pi33  & pi56 ;
  assign n14433 = pi35  & pi54 ;
  assign n14434 = ~n14432 & ~n14433;
  assign n14435 = n2811 & n6911;
  assign n14436 = pi41  & pi48 ;
  assign n14437 = ~n14434 & n14436;
  assign n14438 = ~n14435 & n14437;
  assign n14439 = ~n14435 & ~n14438;
  assign n14440 = ~n14434 & n14439;
  assign n14441 = n14436 & ~n14438;
  assign n14442 = ~n14440 & ~n14441;
  assign n14443 = pi36  & pi53 ;
  assign n14444 = n5055 & n10319;
  assign n14445 = pi37  & pi52 ;
  assign n14446 = ~n7017 & ~n14445;
  assign n14447 = n14443 & ~n14444;
  assign n14448 = ~n14446 & n14447;
  assign n14449 = n14443 & ~n14448;
  assign n14450 = ~n14444 & ~n14448;
  assign n14451 = ~n14446 & n14450;
  assign n14452 = ~n14449 & ~n14451;
  assign n14453 = ~n14442 & ~n14452;
  assign n14454 = ~n14442 & ~n14453;
  assign n14455 = ~n14452 & ~n14453;
  assign n14456 = ~n14454 & ~n14455;
  assign n14457 = pi30  & pi59 ;
  assign n14458 = n3567 & n8144;
  assign n14459 = pi31  & pi58 ;
  assign n14460 = pi32  & pi57 ;
  assign n14461 = ~n14459 & ~n14460;
  assign n14462 = n14457 & ~n14458;
  assign n14463 = ~n14461 & n14462;
  assign n14464 = n14457 & ~n14463;
  assign n14465 = ~n14458 & ~n14463;
  assign n14466 = ~n14461 & n14465;
  assign n14467 = ~n14464 & ~n14466;
  assign n14468 = ~n14456 & ~n14467;
  assign n14469 = ~n14456 & ~n14468;
  assign n14470 = ~n14467 & ~n14468;
  assign n14471 = ~n14469 & ~n14470;
  assign n14472 = n14294 & n14321;
  assign n14473 = ~n14294 & ~n14321;
  assign n14474 = ~n14472 & ~n14473;
  assign n14475 = n14347 & ~n14474;
  assign n14476 = ~n14347 & n14474;
  assign n14477 = ~n14475 & ~n14476;
  assign n14478 = pi45  & pi62 ;
  assign n14479 = pi27  & n14478;
  assign n14480 = n5318 & ~n14479;
  assign n14481 = ~n14479 & ~n14480;
  assign n14482 = pi27  & pi62 ;
  assign n14483 = ~pi45  & ~n14482;
  assign n14484 = n14481 & ~n14483;
  assign n14485 = n5318 & ~n14480;
  assign n14486 = ~n14484 & ~n14485;
  assign n14487 = pi34  & pi55 ;
  assign n14488 = n5277 & n6458;
  assign n14489 = pi42  & pi47 ;
  assign n14490 = pi43  & pi46 ;
  assign n14491 = ~n14489 & ~n14490;
  assign n14492 = n14487 & ~n14488;
  assign n14493 = ~n14491 & n14492;
  assign n14494 = n14487 & ~n14493;
  assign n14495 = ~n14488 & ~n14493;
  assign n14496 = ~n14491 & n14495;
  assign n14497 = ~n14494 & ~n14496;
  assign n14498 = ~n14486 & ~n14497;
  assign n14499 = ~n14486 & ~n14498;
  assign n14500 = ~n14497 & ~n14498;
  assign n14501 = ~n14499 & ~n14500;
  assign n14502 = n2915 & n9054;
  assign n14503 = pi29  & pi60 ;
  assign n14504 = ~n14502 & n14503;
  assign n14505 = pi28  & pi61 ;
  assign n14506 = ~n14502 & n14505;
  assign n14507 = ~n14504 & ~n14506;
  assign n14508 = ~n14398 & ~n14507;
  assign n14509 = ~n14398 & ~n14508;
  assign n14510 = ~n14507 & ~n14508;
  assign n14511 = ~n14509 & ~n14510;
  assign n14512 = ~n14501 & n14511;
  assign n14513 = n14501 & ~n14511;
  assign n14514 = ~n14512 & ~n14513;
  assign n14515 = n14477 & ~n14514;
  assign n14516 = n14477 & ~n14515;
  assign n14517 = ~n14514 & ~n14515;
  assign n14518 = ~n14516 & ~n14517;
  assign n14519 = ~n14471 & ~n14518;
  assign n14520 = ~n14471 & ~n14519;
  assign n14521 = ~n14518 & ~n14519;
  assign n14522 = ~n14520 & ~n14521;
  assign n14523 = ~n14431 & ~n14522;
  assign n14524 = ~n14431 & ~n14523;
  assign n14525 = ~n14522 & ~n14523;
  assign n14526 = ~n14524 & ~n14525;
  assign n14527 = ~n14382 & ~n14385;
  assign n14528 = ~n14359 & ~n14363;
  assign n14529 = n14527 & n14528;
  assign n14530 = ~n14527 & ~n14528;
  assign n14531 = ~n14529 & ~n14530;
  assign n14532 = ~n14388 & ~n14401;
  assign n14533 = ~n14531 & n14532;
  assign n14534 = n14531 & ~n14532;
  assign n14535 = ~n14533 & ~n14534;
  assign n14536 = ~n14270 & ~n14274;
  assign n14537 = ~n14535 & n14536;
  assign n14538 = n14535 & ~n14536;
  assign n14539 = ~n14537 & ~n14538;
  assign n14540 = ~n14407 & ~n14409;
  assign n14541 = n14539 & ~n14540;
  assign n14542 = ~n14539 & n14540;
  assign n14543 = ~n14541 & ~n14542;
  assign n14544 = ~n14526 & n14543;
  assign n14545 = ~n14526 & ~n14544;
  assign n14546 = n14543 & ~n14544;
  assign n14547 = ~n14545 & ~n14546;
  assign n14548 = ~n14379 & ~n14412;
  assign n14549 = ~n14365 & ~n14368;
  assign n14550 = ~n14350 & ~n14356;
  assign n14551 = ~n14309 & ~n14324;
  assign n14552 = n14550 & n14551;
  assign n14553 = ~n14550 & ~n14551;
  assign n14554 = ~n14552 & ~n14553;
  assign n14555 = n14306 & n14335;
  assign n14556 = ~n14306 & ~n14335;
  assign n14557 = ~n14555 & ~n14556;
  assign n14558 = pi26  & pi63 ;
  assign n14559 = n5548 & n5889;
  assign n14560 = pi39  & pi50 ;
  assign n14561 = pi40  & pi49 ;
  assign n14562 = ~n14560 & ~n14561;
  assign n14563 = n14558 & ~n14559;
  assign n14564 = ~n14562 & n14563;
  assign n14565 = n14558 & ~n14564;
  assign n14566 = ~n14559 & ~n14564;
  assign n14567 = ~n14562 & n14566;
  assign n14568 = ~n14565 & ~n14567;
  assign n14569 = n14557 & ~n14568;
  assign n14570 = n14557 & ~n14569;
  assign n14571 = ~n14568 & ~n14569;
  assign n14572 = ~n14570 & ~n14571;
  assign n14573 = ~n14554 & n14572;
  assign n14574 = n14554 & ~n14572;
  assign n14575 = ~n14573 & ~n14574;
  assign n14576 = ~n14549 & n14575;
  assign n14577 = n14549 & ~n14575;
  assign n14578 = ~n14576 & ~n14577;
  assign n14579 = ~n14548 & n14578;
  assign n14580 = n14548 & ~n14578;
  assign n14581 = ~n14579 & ~n14580;
  assign n14582 = ~n14375 & n14414;
  assign n14583 = ~n14372 & ~n14582;
  assign n14584 = n14581 & ~n14583;
  assign n14585 = n14581 & ~n14584;
  assign n14586 = ~n14583 & ~n14584;
  assign n14587 = ~n14585 & ~n14586;
  assign n14588 = ~n14547 & ~n14587;
  assign n14589 = n14547 & n14587;
  assign n14590 = ~n14588 & ~n14589;
  assign n14591 = ~n14430 & n14590;
  assign n14592 = n14430 & ~n14590;
  assign n14593 = ~n14591 & ~n14592;
  assign n14594 = ~n14423 & ~n14428;
  assign n14595 = ~n14593 & n14594;
  assign n14596 = n14593 & ~n14594;
  assign po90  = ~n14595 & ~n14596;
  assign n14598 = ~n14584 & ~n14588;
  assign n14599 = ~n14538 & ~n14541;
  assign n14600 = ~n14515 & ~n14519;
  assign n14601 = n14481 & n14495;
  assign n14602 = ~n14481 & ~n14495;
  assign n14603 = ~n14601 & ~n14602;
  assign n14604 = n14439 & ~n14603;
  assign n14605 = ~n14439 & n14603;
  assign n14606 = ~n14604 & ~n14605;
  assign n14607 = ~n14501 & ~n14511;
  assign n14608 = ~n14498 & ~n14607;
  assign n14609 = ~n14453 & ~n14468;
  assign n14610 = n14608 & n14609;
  assign n14611 = ~n14608 & ~n14609;
  assign n14612 = ~n14610 & ~n14611;
  assign n14613 = n14606 & n14612;
  assign n14614 = ~n14606 & ~n14612;
  assign n14615 = ~n14613 & ~n14614;
  assign n14616 = ~n14600 & n14615;
  assign n14617 = n14600 & ~n14615;
  assign n14618 = ~n14616 & ~n14617;
  assign n14619 = n14599 & ~n14618;
  assign n14620 = ~n14599 & n14618;
  assign n14621 = ~n14619 & ~n14620;
  assign n14622 = ~n14523 & ~n14544;
  assign n14623 = ~n14621 & n14622;
  assign n14624 = n14621 & ~n14622;
  assign n14625 = ~n14623 & ~n14624;
  assign n14626 = ~n14576 & ~n14579;
  assign n14627 = n14450 & n14465;
  assign n14628 = ~n14450 & ~n14465;
  assign n14629 = ~n14627 & ~n14628;
  assign n14630 = n14566 & ~n14629;
  assign n14631 = ~n14566 & n14629;
  assign n14632 = ~n14630 & ~n14631;
  assign n14633 = ~n14530 & ~n14534;
  assign n14634 = ~n14632 & n14633;
  assign n14635 = n14632 & ~n14633;
  assign n14636 = ~n14634 & ~n14635;
  assign n14637 = pi33  & pi57 ;
  assign n14638 = pi34  & pi56 ;
  assign n14639 = ~n14637 & ~n14638;
  assign n14640 = n3900 & n7643;
  assign n14641 = pi35  & pi55 ;
  assign n14642 = ~n14639 & n14641;
  assign n14643 = ~n14640 & n14642;
  assign n14644 = ~n14640 & ~n14643;
  assign n14645 = ~n14639 & n14644;
  assign n14646 = n14641 & ~n14643;
  assign n14647 = ~n14645 & ~n14646;
  assign n14648 = pi36  & pi54 ;
  assign n14649 = n5055 & n9144;
  assign n14650 = pi37  & pi53 ;
  assign n14651 = pi38  & pi52 ;
  assign n14652 = ~n14650 & ~n14651;
  assign n14653 = n14648 & ~n14649;
  assign n14654 = ~n14652 & n14653;
  assign n14655 = n14648 & ~n14654;
  assign n14656 = ~n14649 & ~n14654;
  assign n14657 = ~n14652 & n14656;
  assign n14658 = ~n14655 & ~n14657;
  assign n14659 = ~n14647 & ~n14658;
  assign n14660 = ~n14647 & ~n14659;
  assign n14661 = ~n14658 & ~n14659;
  assign n14662 = ~n14660 & ~n14661;
  assign n14663 = pi42  & pi48 ;
  assign n14664 = n5277 & n6836;
  assign n14665 = ~n7214 & ~n7504;
  assign n14666 = n14663 & ~n14664;
  assign n14667 = ~n14665 & n14666;
  assign n14668 = n14663 & ~n14667;
  assign n14669 = ~n14664 & ~n14667;
  assign n14670 = ~n14665 & n14669;
  assign n14671 = ~n14668 & ~n14670;
  assign n14672 = ~n14662 & ~n14671;
  assign n14673 = ~n14662 & ~n14672;
  assign n14674 = ~n14671 & ~n14672;
  assign n14675 = ~n14673 & ~n14674;
  assign n14676 = n14636 & ~n14675;
  assign n14677 = ~n14636 & n14675;
  assign n14678 = ~n14676 & ~n14677;
  assign n14679 = ~n14626 & n14678;
  assign n14680 = ~n14626 & ~n14679;
  assign n14681 = n14678 & ~n14679;
  assign n14682 = ~n14680 & ~n14681;
  assign n14683 = ~n14553 & ~n14574;
  assign n14684 = ~n14473 & ~n14476;
  assign n14685 = pi39  & pi51 ;
  assign n14686 = n5889 & n6012;
  assign n14687 = pi41  & pi49 ;
  assign n14688 = pi40  & pi50 ;
  assign n14689 = ~n14687 & ~n14688;
  assign n14690 = n14685 & ~n14686;
  assign n14691 = ~n14689 & n14690;
  assign n14692 = n14685 & ~n14691;
  assign n14693 = ~n14686 & ~n14691;
  assign n14694 = ~n14689 & n14693;
  assign n14695 = ~n14692 & ~n14694;
  assign n14696 = ~n14684 & ~n14695;
  assign n14697 = ~n14684 & ~n14696;
  assign n14698 = ~n14695 & ~n14696;
  assign n14699 = ~n14697 & ~n14698;
  assign n14700 = ~n14556 & ~n14569;
  assign n14701 = n14699 & n14700;
  assign n14702 = ~n14699 & ~n14700;
  assign n14703 = ~n14701 & ~n14702;
  assign n14704 = pi28  & pi62 ;
  assign n14705 = pi29  & pi61 ;
  assign n14706 = ~n14704 & ~n14705;
  assign n14707 = n2915 & n9567;
  assign n14708 = pi27  & pi63 ;
  assign n14709 = ~n14706 & n14708;
  assign n14710 = ~n14707 & n14709;
  assign n14711 = ~n14707 & ~n14710;
  assign n14712 = ~n14706 & n14711;
  assign n14713 = n14708 & ~n14710;
  assign n14714 = ~n14712 & ~n14713;
  assign n14715 = ~n14502 & ~n14508;
  assign n14716 = n3567 & n9402;
  assign n14717 = pi32  & pi58 ;
  assign n14718 = pi31  & pi59 ;
  assign n14719 = ~n14717 & ~n14718;
  assign n14720 = ~n14716 & ~n14719;
  assign n14721 = pi30  & pi60 ;
  assign n14722 = ~n14720 & ~n14721;
  assign n14723 = n14720 & n14721;
  assign n14724 = ~n14722 & ~n14723;
  assign n14725 = ~n14715 & n14724;
  assign n14726 = ~n14715 & ~n14725;
  assign n14727 = n14724 & ~n14725;
  assign n14728 = ~n14726 & ~n14727;
  assign n14729 = ~n14714 & ~n14728;
  assign n14730 = n14714 & n14728;
  assign n14731 = ~n14729 & ~n14730;
  assign n14732 = n14703 & n14731;
  assign n14733 = n14703 & ~n14732;
  assign n14734 = n14731 & ~n14732;
  assign n14735 = ~n14733 & ~n14734;
  assign n14736 = ~n14683 & ~n14735;
  assign n14737 = ~n14683 & ~n14736;
  assign n14738 = ~n14735 & ~n14736;
  assign n14739 = ~n14737 & ~n14738;
  assign n14740 = ~n14682 & ~n14739;
  assign n14741 = ~n14682 & ~n14740;
  assign n14742 = ~n14739 & ~n14740;
  assign n14743 = ~n14741 & ~n14742;
  assign n14744 = ~n14625 & n14743;
  assign n14745 = n14625 & ~n14743;
  assign n14746 = ~n14744 & ~n14745;
  assign n14747 = n14598 & ~n14746;
  assign n14748 = ~n14598 & n14746;
  assign n14749 = ~n14747 & ~n14748;
  assign n14750 = ~n14591 & ~n14596;
  assign n14751 = ~n14749 & n14750;
  assign n14752 = ~n14747 & ~n14750;
  assign n14753 = ~n14748 & n14752;
  assign po91  = ~n14751 & ~n14753;
  assign n14755 = ~n14748 & ~n14752;
  assign n14756 = ~n14624 & ~n14745;
  assign n14757 = n14656 & n14711;
  assign n14758 = ~n14656 & ~n14711;
  assign n14759 = ~n14757 & ~n14758;
  assign n14760 = ~n14716 & ~n14723;
  assign n14761 = ~n14759 & n14760;
  assign n14762 = n14759 & ~n14760;
  assign n14763 = ~n14761 & ~n14762;
  assign n14764 = ~n14696 & ~n14702;
  assign n14765 = ~n14763 & n14764;
  assign n14766 = n14763 & ~n14764;
  assign n14767 = ~n14765 & ~n14766;
  assign n14768 = pi40  & pi51 ;
  assign n14769 = pi41  & pi50 ;
  assign n14770 = ~n14768 & ~n14769;
  assign n14771 = n6012 & n6114;
  assign n14772 = pi28  & pi63 ;
  assign n14773 = ~n14770 & n14772;
  assign n14774 = ~n14771 & n14773;
  assign n14775 = ~n14771 & ~n14774;
  assign n14776 = ~n14770 & n14775;
  assign n14777 = n14772 & ~n14774;
  assign n14778 = ~n14776 & ~n14777;
  assign n14779 = pi35  & pi56 ;
  assign n14780 = n5823 & n6836;
  assign n14781 = pi43  & pi48 ;
  assign n14782 = pi44  & pi47 ;
  assign n14783 = ~n14781 & ~n14782;
  assign n14784 = n14779 & ~n14780;
  assign n14785 = ~n14783 & n14784;
  assign n14786 = n14779 & ~n14785;
  assign n14787 = ~n14780 & ~n14785;
  assign n14788 = ~n14783 & n14787;
  assign n14789 = ~n14786 & ~n14788;
  assign n14790 = ~n14778 & ~n14789;
  assign n14791 = ~n14778 & ~n14790;
  assign n14792 = ~n14789 & ~n14790;
  assign n14793 = ~n14791 & ~n14792;
  assign n14794 = pi46  & pi62 ;
  assign n14795 = pi29  & n14794;
  assign n14796 = n7513 & ~n14795;
  assign n14797 = n7513 & ~n14796;
  assign n14798 = ~n14795 & ~n14796;
  assign n14799 = pi29  & pi62 ;
  assign n14800 = ~pi46  & ~n14799;
  assign n14801 = n14798 & ~n14800;
  assign n14802 = ~n14797 & ~n14801;
  assign n14803 = ~n14793 & ~n14802;
  assign n14804 = ~n14793 & ~n14803;
  assign n14805 = ~n14802 & ~n14803;
  assign n14806 = ~n14804 & ~n14805;
  assign n14807 = ~n14767 & n14806;
  assign n14808 = n14767 & ~n14806;
  assign n14809 = ~n14807 & ~n14808;
  assign n14810 = ~n14616 & ~n14620;
  assign n14811 = n14809 & ~n14810;
  assign n14812 = ~n14809 & n14810;
  assign n14813 = ~n14811 & ~n14812;
  assign n14814 = ~n14602 & ~n14605;
  assign n14815 = n10665 & n13270;
  assign n14816 = pi34  & pi57 ;
  assign n14817 = pi36  & pi55 ;
  assign n14818 = ~n14816 & ~n14817;
  assign n14819 = n7427 & ~n14815;
  assign n14820 = ~n14818 & n14819;
  assign n14821 = n7427 & ~n14820;
  assign n14822 = ~n14815 & ~n14820;
  assign n14823 = ~n14818 & n14822;
  assign n14824 = ~n14821 & ~n14823;
  assign n14825 = ~n14814 & ~n14824;
  assign n14826 = ~n14814 & ~n14825;
  assign n14827 = ~n14824 & ~n14825;
  assign n14828 = ~n14826 & ~n14827;
  assign n14829 = ~n14628 & ~n14631;
  assign n14830 = n14828 & n14829;
  assign n14831 = ~n14828 & ~n14829;
  assign n14832 = ~n14830 & ~n14831;
  assign n14833 = ~n14611 & ~n14613;
  assign n14834 = pi33  & pi58 ;
  assign n14835 = ~n7740 & ~n14834;
  assign n14836 = n6138 & n9402;
  assign n14837 = pi31  & pi60 ;
  assign n14838 = ~n14835 & n14837;
  assign n14839 = ~n14836 & n14838;
  assign n14840 = ~n14836 & ~n14839;
  assign n14841 = ~n14835 & n14840;
  assign n14842 = n14837 & ~n14839;
  assign n14843 = ~n14841 & ~n14842;
  assign n14844 = pi37  & pi54 ;
  assign n14845 = n4736 & n9144;
  assign n14846 = pi38  & pi53 ;
  assign n14847 = pi39  & pi52 ;
  assign n14848 = ~n14846 & ~n14847;
  assign n14849 = n14844 & ~n14845;
  assign n14850 = ~n14848 & n14849;
  assign n14851 = n14844 & ~n14850;
  assign n14852 = ~n14845 & ~n14850;
  assign n14853 = ~n14848 & n14852;
  assign n14854 = ~n14851 & ~n14853;
  assign n14855 = ~n14693 & ~n14854;
  assign n14856 = ~n14693 & ~n14855;
  assign n14857 = ~n14854 & ~n14855;
  assign n14858 = ~n14856 & ~n14857;
  assign n14859 = ~n14843 & ~n14858;
  assign n14860 = ~n14843 & ~n14859;
  assign n14861 = ~n14858 & ~n14859;
  assign n14862 = ~n14860 & ~n14861;
  assign n14863 = ~n14833 & ~n14862;
  assign n14864 = ~n14833 & ~n14863;
  assign n14865 = ~n14862 & ~n14863;
  assign n14866 = ~n14864 & ~n14865;
  assign n14867 = n14832 & ~n14866;
  assign n14868 = ~n14832 & n14866;
  assign n14869 = ~n14867 & ~n14868;
  assign n14870 = n14813 & n14869;
  assign n14871 = n14813 & ~n14870;
  assign n14872 = n14869 & ~n14870;
  assign n14873 = ~n14871 & ~n14872;
  assign n14874 = ~n14679 & ~n14740;
  assign n14875 = ~n14732 & ~n14736;
  assign n14876 = ~n14635 & ~n14676;
  assign n14877 = pi30  & pi61 ;
  assign n14878 = ~n14669 & n14877;
  assign n14879 = n14669 & ~n14877;
  assign n14880 = ~n14878 & ~n14879;
  assign n14881 = n14644 & ~n14880;
  assign n14882 = ~n14644 & n14880;
  assign n14883 = ~n14881 & ~n14882;
  assign n14884 = ~n14725 & ~n14729;
  assign n14885 = ~n14659 & ~n14672;
  assign n14886 = n14884 & n14885;
  assign n14887 = ~n14884 & ~n14885;
  assign n14888 = ~n14886 & ~n14887;
  assign n14889 = n14883 & n14888;
  assign n14890 = ~n14883 & ~n14888;
  assign n14891 = ~n14889 & ~n14890;
  assign n14892 = ~n14876 & n14891;
  assign n14893 = ~n14876 & ~n14892;
  assign n14894 = n14891 & ~n14892;
  assign n14895 = ~n14893 & ~n14894;
  assign n14896 = ~n14875 & ~n14895;
  assign n14897 = ~n14875 & ~n14896;
  assign n14898 = ~n14895 & ~n14896;
  assign n14899 = ~n14897 & ~n14898;
  assign n14900 = ~n14874 & ~n14899;
  assign n14901 = ~n14874 & ~n14900;
  assign n14902 = ~n14899 & ~n14900;
  assign n14903 = ~n14901 & ~n14902;
  assign n14904 = ~n14873 & n14903;
  assign n14905 = n14873 & ~n14903;
  assign n14906 = ~n14904 & ~n14905;
  assign n14907 = ~n14756 & ~n14906;
  assign n14908 = n14756 & n14906;
  assign n14909 = ~n14907 & ~n14908;
  assign n14910 = ~n14755 & ~n14909;
  assign n14911 = n14755 & n14909;
  assign po92  = n14910 | n14911;
  assign n14913 = ~n14755 & ~n14908;
  assign n14914 = ~n14907 & ~n14913;
  assign n14915 = ~n14892 & ~n14896;
  assign n14916 = ~n14863 & ~n14867;
  assign n14917 = ~n14887 & ~n14889;
  assign n14918 = n2680 & n9567;
  assign n14919 = pi31  & pi61 ;
  assign n14920 = ~n14918 & n14919;
  assign n14921 = pi30  & pi62 ;
  assign n14922 = ~n14918 & n14921;
  assign n14923 = ~n14920 & ~n14922;
  assign n14924 = ~n14798 & ~n14923;
  assign n14925 = ~n14798 & ~n14924;
  assign n14926 = ~n14923 & ~n14924;
  assign n14927 = ~n14925 & ~n14926;
  assign n14928 = pi39  & pi53 ;
  assign n14929 = n6012 & n10319;
  assign n14930 = pi40  & pi52 ;
  assign n14931 = pi41  & pi51 ;
  assign n14932 = ~n14930 & ~n14931;
  assign n14933 = n14928 & ~n14929;
  assign n14934 = ~n14932 & n14933;
  assign n14935 = n14928 & ~n14934;
  assign n14936 = ~n14929 & ~n14934;
  assign n14937 = ~n14932 & n14936;
  assign n14938 = ~n14935 & ~n14937;
  assign n14939 = ~n14927 & ~n14938;
  assign n14940 = ~n14927 & ~n14939;
  assign n14941 = ~n14938 & ~n14939;
  assign n14942 = ~n14940 & ~n14941;
  assign n14943 = ~n14878 & ~n14882;
  assign n14944 = n14942 & n14943;
  assign n14945 = ~n14942 & ~n14943;
  assign n14946 = ~n14944 & ~n14945;
  assign n14947 = pi42  & pi50 ;
  assign n14948 = pi35  & pi57 ;
  assign n14949 = ~n14947 & ~n14948;
  assign n14950 = n14947 & n14948;
  assign n14951 = pi34  & pi58 ;
  assign n14952 = ~n14949 & n14951;
  assign n14953 = ~n14950 & n14952;
  assign n14954 = ~n14950 & ~n14953;
  assign n14955 = ~n14949 & n14954;
  assign n14956 = n14951 & ~n14953;
  assign n14957 = ~n14955 & ~n14956;
  assign n14958 = pi43  & pi49 ;
  assign n14959 = n5318 & n5823;
  assign n14960 = pi44  & pi48 ;
  assign n14961 = ~n4899 & ~n14960;
  assign n14962 = n14958 & ~n14959;
  assign n14963 = ~n14961 & n14962;
  assign n14964 = n14958 & ~n14963;
  assign n14965 = ~n14959 & ~n14963;
  assign n14966 = ~n14961 & n14965;
  assign n14967 = ~n14964 & ~n14966;
  assign n14968 = ~n14957 & ~n14967;
  assign n14969 = ~n14957 & ~n14968;
  assign n14970 = ~n14967 & ~n14968;
  assign n14971 = ~n14969 & ~n14970;
  assign n14972 = pi36  & pi56 ;
  assign n14973 = pi33  & pi59 ;
  assign n14974 = n12766 & n14973;
  assign n14975 = ~n12766 & ~n14973;
  assign n14976 = n14972 & ~n14974;
  assign n14977 = ~n14975 & n14976;
  assign n14978 = n14972 & ~n14977;
  assign n14979 = ~n14974 & ~n14977;
  assign n14980 = ~n14975 & n14979;
  assign n14981 = ~n14978 & ~n14980;
  assign n14982 = ~n14971 & ~n14981;
  assign n14983 = ~n14971 & ~n14982;
  assign n14984 = ~n14981 & ~n14982;
  assign n14985 = ~n14983 & ~n14984;
  assign n14986 = ~n14946 & n14985;
  assign n14987 = n14946 & ~n14985;
  assign n14988 = ~n14986 & ~n14987;
  assign n14989 = ~n14917 & n14988;
  assign n14990 = n14917 & ~n14988;
  assign n14991 = ~n14989 & ~n14990;
  assign n14992 = ~n14916 & n14991;
  assign n14993 = n14916 & ~n14991;
  assign n14994 = ~n14992 & ~n14993;
  assign n14995 = ~n14915 & n14994;
  assign n14996 = n14915 & ~n14994;
  assign n14997 = ~n14995 & ~n14996;
  assign n14998 = ~n14811 & ~n14870;
  assign n14999 = ~n14855 & ~n14859;
  assign n15000 = ~n14758 & ~n14762;
  assign n15001 = n14999 & n15000;
  assign n15002 = ~n14999 & ~n15000;
  assign n15003 = ~n15001 & ~n15002;
  assign n15004 = ~n14790 & ~n14803;
  assign n15005 = ~n15003 & n15004;
  assign n15006 = n15003 & ~n15004;
  assign n15007 = ~n15005 & ~n15006;
  assign n15008 = ~n14766 & ~n14808;
  assign n15009 = ~n14825 & ~n14831;
  assign n15010 = n14840 & n14852;
  assign n15011 = ~n14840 & ~n14852;
  assign n15012 = ~n15010 & ~n15011;
  assign n15013 = n14775 & ~n15012;
  assign n15014 = ~n14775 & n15012;
  assign n15015 = ~n15013 & ~n15014;
  assign n15016 = n14787 & n14822;
  assign n15017 = ~n14787 & ~n14822;
  assign n15018 = ~n15016 & ~n15017;
  assign n15019 = pi32  & pi60 ;
  assign n15020 = pi37  & pi55 ;
  assign n15021 = pi38  & pi54 ;
  assign n15022 = ~n15020 & ~n15021;
  assign n15023 = n5055 & n9891;
  assign n15024 = n15019 & ~n15022;
  assign n15025 = ~n15023 & n15024;
  assign n15026 = n15019 & ~n15025;
  assign n15027 = ~n15023 & ~n15025;
  assign n15028 = ~n15022 & n15027;
  assign n15029 = ~n15026 & ~n15028;
  assign n15030 = n15018 & ~n15029;
  assign n15031 = n15018 & ~n15030;
  assign n15032 = ~n15029 & ~n15030;
  assign n15033 = ~n15031 & ~n15032;
  assign n15034 = ~n15015 & n15033;
  assign n15035 = n15015 & ~n15033;
  assign n15036 = ~n15034 & ~n15035;
  assign n15037 = ~n15009 & n15036;
  assign n15038 = n15009 & ~n15036;
  assign n15039 = ~n15037 & ~n15038;
  assign n15040 = ~n15008 & n15039;
  assign n15041 = n15008 & ~n15039;
  assign n15042 = ~n15040 & ~n15041;
  assign n15043 = n15007 & n15042;
  assign n15044 = ~n15007 & ~n15042;
  assign n15045 = ~n15043 & ~n15044;
  assign n15046 = ~n14998 & n15045;
  assign n15047 = n14998 & ~n15045;
  assign n15048 = ~n15046 & ~n15047;
  assign n15049 = n14997 & n15048;
  assign n15050 = ~n14997 & ~n15048;
  assign n15051 = ~n15049 & ~n15050;
  assign n15052 = ~n14873 & ~n14903;
  assign n15053 = ~n14900 & ~n15052;
  assign n15054 = ~n15051 & n15053;
  assign n15055 = n15051 & ~n15053;
  assign n15056 = ~n15054 & ~n15055;
  assign n15057 = n14914 & ~n15056;
  assign n15058 = ~n14914 & ~n15054;
  assign n15059 = ~n15055 & n15058;
  assign po93  = ~n15057 & ~n15059;
  assign n15061 = ~n15055 & ~n15058;
  assign n15062 = ~n15046 & ~n15049;
  assign n15063 = ~n14992 & ~n14995;
  assign n15064 = ~n15017 & ~n15030;
  assign n15065 = ~n15011 & ~n15014;
  assign n15066 = n15064 & n15065;
  assign n15067 = ~n15064 & ~n15065;
  assign n15068 = ~n15066 & ~n15067;
  assign n15069 = ~n14968 & ~n14982;
  assign n15070 = ~n15068 & n15069;
  assign n15071 = n15068 & ~n15069;
  assign n15072 = ~n15070 & ~n15071;
  assign n15073 = ~n15035 & ~n15037;
  assign n15074 = n15072 & ~n15073;
  assign n15075 = ~n15072 & n15073;
  assign n15076 = ~n15074 & ~n15075;
  assign n15077 = ~n14939 & ~n14945;
  assign n15078 = n14954 & n14965;
  assign n15079 = ~n14954 & ~n14965;
  assign n15080 = ~n15078 & ~n15079;
  assign n15081 = n14936 & ~n15080;
  assign n15082 = ~n14936 & n15080;
  assign n15083 = ~n15081 & ~n15082;
  assign n15084 = n14979 & n15027;
  assign n15085 = ~n14979 & ~n15027;
  assign n15086 = ~n15084 & ~n15085;
  assign n15087 = ~n14918 & ~n14924;
  assign n15088 = ~n15086 & n15087;
  assign n15089 = n15086 & ~n15087;
  assign n15090 = ~n15088 & ~n15089;
  assign n15091 = n15083 & n15090;
  assign n15092 = ~n15083 & ~n15090;
  assign n15093 = ~n15091 & ~n15092;
  assign n15094 = ~n15077 & n15093;
  assign n15095 = n15077 & ~n15093;
  assign n15096 = ~n15094 & ~n15095;
  assign n15097 = n15076 & n15096;
  assign n15098 = ~n15076 & ~n15096;
  assign n15099 = ~n15097 & ~n15098;
  assign n15100 = n15063 & ~n15099;
  assign n15101 = ~n15063 & n15099;
  assign n15102 = ~n15100 & ~n15101;
  assign n15103 = ~n15040 & ~n15043;
  assign n15104 = ~n14987 & ~n14989;
  assign n15105 = ~n15002 & ~n15006;
  assign n15106 = pi32  & pi61 ;
  assign n15107 = pi33  & pi60 ;
  assign n15108 = ~n15106 & ~n15107;
  assign n15109 = n6138 & n9054;
  assign n15110 = pi30  & pi63 ;
  assign n15111 = ~n15108 & n15110;
  assign n15112 = ~n15109 & n15111;
  assign n15113 = ~n15109 & ~n15112;
  assign n15114 = ~n15108 & n15113;
  assign n15115 = n15110 & ~n15112;
  assign n15116 = ~n15114 & ~n15115;
  assign n15117 = pi35  & pi58 ;
  assign n15118 = pi54  & pi57 ;
  assign n15119 = n11756 & n15118;
  assign n15120 = pi39  & pi54 ;
  assign n15121 = pi36  & pi57 ;
  assign n15122 = ~n15120 & ~n15121;
  assign n15123 = n15117 & ~n15119;
  assign n15124 = ~n15122 & n15123;
  assign n15125 = n15117 & ~n15124;
  assign n15126 = ~n15119 & ~n15124;
  assign n15127 = ~n15122 & n15126;
  assign n15128 = ~n15125 & ~n15127;
  assign n15129 = ~n15116 & ~n15128;
  assign n15130 = ~n15116 & ~n15129;
  assign n15131 = ~n15128 & ~n15129;
  assign n15132 = ~n15130 & ~n15131;
  assign n15133 = pi34  & pi59 ;
  assign n15134 = n6012 & n9144;
  assign n15135 = pi40  & pi53 ;
  assign n15136 = pi41  & pi52 ;
  assign n15137 = ~n15135 & ~n15136;
  assign n15138 = n15133 & ~n15134;
  assign n15139 = ~n15137 & n15138;
  assign n15140 = n15133 & ~n15139;
  assign n15141 = ~n15134 & ~n15139;
  assign n15142 = ~n15137 & n15141;
  assign n15143 = ~n15140 & ~n15142;
  assign n15144 = ~n15132 & ~n15143;
  assign n15145 = ~n15132 & ~n15144;
  assign n15146 = ~n15143 & ~n15144;
  assign n15147 = ~n15145 & ~n15146;
  assign n15148 = pi45  & pi48 ;
  assign n15149 = pi38  & pi55 ;
  assign n15150 = ~n15148 & ~n15149;
  assign n15151 = pi45  & pi55 ;
  assign n15152 = n6474 & n15151;
  assign n15153 = pi37  & pi56 ;
  assign n15154 = ~n15150 & n15153;
  assign n15155 = ~n15152 & n15154;
  assign n15156 = ~n15152 & ~n15155;
  assign n15157 = ~n15150 & n15156;
  assign n15158 = n15153 & ~n15155;
  assign n15159 = ~n15157 & ~n15158;
  assign n15160 = pi42  & pi51 ;
  assign n15161 = n5889 & n6836;
  assign n15162 = pi43  & pi50 ;
  assign n15163 = ~n7690 & ~n15162;
  assign n15164 = n15160 & ~n15161;
  assign n15165 = ~n15163 & n15164;
  assign n15166 = n15160 & ~n15165;
  assign n15167 = ~n15161 & ~n15165;
  assign n15168 = ~n15163 & n15167;
  assign n15169 = ~n15166 & ~n15168;
  assign n15170 = ~n15159 & ~n15169;
  assign n15171 = ~n15159 & ~n15170;
  assign n15172 = ~n15169 & ~n15170;
  assign n15173 = ~n15171 & ~n15172;
  assign n15174 = pi47  & pi62 ;
  assign n15175 = pi31  & n15174;
  assign n15176 = n5277 & ~n15175;
  assign n15177 = n5277 & ~n15176;
  assign n15178 = ~n15175 & ~n15176;
  assign n15179 = pi31  & pi62 ;
  assign n15180 = ~pi47  & ~n15179;
  assign n15181 = n15178 & ~n15180;
  assign n15182 = ~n15177 & ~n15181;
  assign n15183 = ~n15173 & ~n15182;
  assign n15184 = ~n15173 & ~n15183;
  assign n15185 = ~n15182 & ~n15183;
  assign n15186 = ~n15184 & ~n15185;
  assign n15187 = n15147 & n15186;
  assign n15188 = ~n15147 & ~n15186;
  assign n15189 = ~n15187 & ~n15188;
  assign n15190 = ~n15105 & n15189;
  assign n15191 = n15105 & ~n15189;
  assign n15192 = ~n15190 & ~n15191;
  assign n15193 = ~n15104 & n15192;
  assign n15194 = n15104 & ~n15192;
  assign n15195 = ~n15193 & ~n15194;
  assign n15196 = n15103 & ~n15195;
  assign n15197 = ~n15103 & n15195;
  assign n15198 = ~n15196 & ~n15197;
  assign n15199 = n15102 & n15198;
  assign n15200 = ~n15102 & ~n15198;
  assign n15201 = ~n15199 & ~n15200;
  assign n15202 = ~n15062 & n15201;
  assign n15203 = n15062 & ~n15201;
  assign n15204 = ~n15202 & ~n15203;
  assign n15205 = ~n15061 & ~n15204;
  assign n15206 = n15061 & n15204;
  assign po94  = n15205 | n15206;
  assign n15208 = ~n15193 & ~n15197;
  assign n15209 = ~n15188 & ~n15190;
  assign n15210 = ~n15085 & ~n15089;
  assign n15211 = ~n15079 & ~n15082;
  assign n15212 = n15210 & n15211;
  assign n15213 = ~n15210 & ~n15211;
  assign n15214 = ~n15212 & ~n15213;
  assign n15215 = ~n15129 & ~n15144;
  assign n15216 = ~n15214 & n15215;
  assign n15217 = n15214 & ~n15215;
  assign n15218 = ~n15216 & ~n15217;
  assign n15219 = ~n15091 & ~n15094;
  assign n15220 = n15218 & ~n15219;
  assign n15221 = ~n15218 & n15219;
  assign n15222 = ~n15220 & ~n15221;
  assign n15223 = ~n15209 & n15222;
  assign n15224 = n15209 & ~n15222;
  assign n15225 = ~n15223 & ~n15224;
  assign n15226 = n15208 & ~n15225;
  assign n15227 = ~n15208 & n15225;
  assign n15228 = ~n15226 & ~n15227;
  assign n15229 = ~n15074 & ~n15097;
  assign n15230 = n12255 & ~n15178;
  assign n15231 = ~n12255 & n15178;
  assign n15232 = ~n15230 & ~n15231;
  assign n15233 = n15156 & ~n15232;
  assign n15234 = ~n15156 & n15232;
  assign n15235 = ~n15233 & ~n15234;
  assign n15236 = ~n15170 & ~n15183;
  assign n15237 = ~n15235 & n15236;
  assign n15238 = n15235 & ~n15236;
  assign n15239 = ~n15237 & ~n15238;
  assign n15240 = n15113 & n15126;
  assign n15241 = ~n15113 & ~n15126;
  assign n15242 = ~n15240 & ~n15241;
  assign n15243 = n15141 & ~n15242;
  assign n15244 = ~n15141 & n15242;
  assign n15245 = ~n15243 & ~n15244;
  assign n15246 = n15239 & n15245;
  assign n15247 = ~n15239 & ~n15245;
  assign n15248 = ~n15246 & ~n15247;
  assign n15249 = ~n15229 & n15248;
  assign n15250 = n15229 & ~n15248;
  assign n15251 = ~n15249 & ~n15250;
  assign n15252 = pi44  & pi50 ;
  assign n15253 = pi43  & pi51 ;
  assign n15254 = ~n15252 & ~n15253;
  assign n15255 = n6114 & n6836;
  assign n15256 = pi36  & pi58 ;
  assign n15257 = ~n15254 & n15256;
  assign n15258 = ~n15255 & n15257;
  assign n15259 = ~n15255 & ~n15258;
  assign n15260 = ~n15254 & n15259;
  assign n15261 = n15256 & ~n15258;
  assign n15262 = ~n15260 & ~n15261;
  assign n15263 = pi40  & pi54 ;
  assign n15264 = n5235 & n9144;
  assign n15265 = pi41  & pi53 ;
  assign n15266 = pi42  & pi52 ;
  assign n15267 = ~n15265 & ~n15266;
  assign n15268 = n15263 & ~n15264;
  assign n15269 = ~n15267 & n15268;
  assign n15270 = n15263 & ~n15269;
  assign n15271 = ~n15264 & ~n15269;
  assign n15272 = ~n15267 & n15271;
  assign n15273 = ~n15270 & ~n15272;
  assign n15274 = ~n15262 & ~n15273;
  assign n15275 = ~n15262 & ~n15274;
  assign n15276 = ~n15273 & ~n15274;
  assign n15277 = ~n15275 & ~n15276;
  assign n15278 = pi46  & pi48 ;
  assign n15279 = pi38  & pi56 ;
  assign n15280 = n15278 & n15279;
  assign n15281 = ~n15278 & ~n15279;
  assign n15282 = n8001 & ~n15280;
  assign n15283 = ~n15281 & n15282;
  assign n15284 = n8001 & ~n15283;
  assign n15285 = ~n15280 & ~n15283;
  assign n15286 = ~n15281 & n15285;
  assign n15287 = ~n15284 & ~n15286;
  assign n15288 = ~n15277 & ~n15287;
  assign n15289 = ~n15277 & ~n15288;
  assign n15290 = ~n15287 & ~n15288;
  assign n15291 = ~n15289 & ~n15290;
  assign n15292 = ~n15067 & ~n15071;
  assign n15293 = n15291 & n15292;
  assign n15294 = ~n15291 & ~n15292;
  assign n15295 = ~n15293 & ~n15294;
  assign n15296 = pi32  & pi62 ;
  assign n15297 = pi59  & pi61 ;
  assign n15298 = n2811 & n15297;
  assign n15299 = pi33  & pi61 ;
  assign n15300 = pi35  & pi59 ;
  assign n15301 = ~n15299 & ~n15300;
  assign n15302 = n15296 & ~n15298;
  assign n15303 = ~n15301 & n15302;
  assign n15304 = n15296 & ~n15303;
  assign n15305 = ~n15298 & ~n15303;
  assign n15306 = ~n15301 & n15305;
  assign n15307 = ~n15304 & ~n15306;
  assign n15308 = n15167 & ~n15307;
  assign n15309 = ~n15167 & n15307;
  assign n15310 = ~n15308 & ~n15309;
  assign n15311 = pi37  & pi57 ;
  assign n15312 = pi34  & pi60 ;
  assign n15313 = pi39  & pi55 ;
  assign n15314 = n15312 & n15313;
  assign n15315 = ~n15312 & ~n15313;
  assign n15316 = n15311 & ~n15314;
  assign n15317 = ~n15315 & n15316;
  assign n15318 = n15311 & ~n15317;
  assign n15319 = ~n15314 & ~n15317;
  assign n15320 = ~n15315 & n15319;
  assign n15321 = ~n15318 & ~n15320;
  assign n15322 = ~n15310 & ~n15321;
  assign n15323 = n15310 & n15321;
  assign n15324 = ~n15322 & ~n15323;
  assign n15325 = n15295 & n15324;
  assign n15326 = ~n15295 & ~n15324;
  assign n15327 = ~n15325 & ~n15326;
  assign n15328 = n15251 & n15327;
  assign n15329 = n15251 & ~n15328;
  assign n15330 = n15327 & ~n15328;
  assign n15331 = ~n15329 & ~n15330;
  assign n15332 = ~n15228 & n15331;
  assign n15333 = n15228 & ~n15331;
  assign n15334 = ~n15332 & ~n15333;
  assign n15335 = ~n15101 & ~n15199;
  assign n15336 = ~n15334 & n15335;
  assign n15337 = n15334 & ~n15335;
  assign n15338 = ~n15336 & ~n15337;
  assign n15339 = ~n15061 & ~n15203;
  assign n15340 = ~n15202 & ~n15339;
  assign n15341 = ~n15338 & n15340;
  assign n15342 = n15338 & ~n15340;
  assign po95  = ~n15341 & ~n15342;
  assign n15344 = ~n15249 & ~n15328;
  assign n15345 = ~n15294 & ~n15325;
  assign n15346 = n4691 & n8854;
  assign n15347 = pi36  & pi59 ;
  assign n15348 = ~n15346 & n15347;
  assign n15349 = pi35  & pi60 ;
  assign n15350 = ~n15346 & n15349;
  assign n15351 = ~n15348 & ~n15350;
  assign n15352 = ~n15285 & ~n15351;
  assign n15353 = ~n15285 & ~n15352;
  assign n15354 = ~n15351 & ~n15352;
  assign n15355 = ~n15353 & ~n15354;
  assign n15356 = ~n15230 & ~n15234;
  assign n15357 = n15355 & n15356;
  assign n15358 = ~n15355 & ~n15356;
  assign n15359 = ~n15357 & ~n15358;
  assign n15360 = ~n15241 & ~n15244;
  assign n15361 = ~n15359 & n15360;
  assign n15362 = n15359 & ~n15360;
  assign n15363 = ~n15361 & ~n15362;
  assign n15364 = ~n15238 & ~n15246;
  assign n15365 = n15363 & ~n15364;
  assign n15366 = ~n15363 & n15364;
  assign n15367 = ~n15365 & ~n15366;
  assign n15368 = ~n15345 & n15367;
  assign n15369 = n15345 & ~n15367;
  assign n15370 = ~n15368 & ~n15369;
  assign n15371 = n15344 & ~n15370;
  assign n15372 = ~n15344 & n15370;
  assign n15373 = ~n15371 & ~n15372;
  assign n15374 = pi48  & pi62 ;
  assign n15375 = pi33  & n15374;
  assign n15376 = n5823 & ~n15375;
  assign n15377 = ~n15375 & ~n15376;
  assign n15378 = pi33  & pi62 ;
  assign n15379 = ~pi48  & ~n15378;
  assign n15380 = n15377 & ~n15379;
  assign n15381 = n5823 & ~n15376;
  assign n15382 = ~n15380 & ~n15381;
  assign n15383 = pi39  & pi56 ;
  assign n15384 = pi45  & pi50 ;
  assign n15385 = pi46  & pi49 ;
  assign n15386 = ~n15384 & ~n15385;
  assign n15387 = n5889 & n7513;
  assign n15388 = n15383 & ~n15386;
  assign n15389 = ~n15387 & n15388;
  assign n15390 = n15383 & ~n15389;
  assign n15391 = ~n15387 & ~n15389;
  assign n15392 = ~n15386 & n15391;
  assign n15393 = ~n15390 & ~n15392;
  assign n15394 = ~n15382 & ~n15393;
  assign n15395 = ~n15382 & ~n15394;
  assign n15396 = ~n15393 & ~n15394;
  assign n15397 = ~n15395 & ~n15396;
  assign n15398 = pi42  & pi53 ;
  assign n15399 = n6836 & n10319;
  assign n15400 = pi43  & pi52 ;
  assign n15401 = ~n7986 & ~n15400;
  assign n15402 = n15398 & ~n15399;
  assign n15403 = ~n15401 & n15402;
  assign n15404 = n15398 & ~n15403;
  assign n15405 = ~n15399 & ~n15403;
  assign n15406 = ~n15401 & n15405;
  assign n15407 = ~n15404 & ~n15406;
  assign n15408 = ~n15397 & ~n15407;
  assign n15409 = ~n15397 & ~n15408;
  assign n15410 = ~n15407 & ~n15408;
  assign n15411 = ~n15409 & ~n15410;
  assign n15412 = ~n15213 & ~n15217;
  assign n15413 = n15411 & n15412;
  assign n15414 = ~n15411 & ~n15412;
  assign n15415 = ~n15413 & ~n15414;
  assign n15416 = pi32  & pi63 ;
  assign n15417 = pi34  & pi61 ;
  assign n15418 = ~n15416 & ~n15417;
  assign n15419 = n3827 & n9236;
  assign n15420 = pi41  & pi54 ;
  assign n15421 = ~n15418 & n15420;
  assign n15422 = ~n15419 & n15421;
  assign n15423 = ~n15419 & ~n15422;
  assign n15424 = ~n15418 & n15423;
  assign n15425 = n15420 & ~n15422;
  assign n15426 = ~n15424 & ~n15425;
  assign n15427 = pi37  & pi58 ;
  assign n15428 = n3558 & n13270;
  assign n15429 = pi38  & pi57 ;
  assign n15430 = pi40  & pi55 ;
  assign n15431 = ~n15429 & ~n15430;
  assign n15432 = n15427 & ~n15428;
  assign n15433 = ~n15431 & n15432;
  assign n15434 = n15427 & ~n15433;
  assign n15435 = ~n15428 & ~n15433;
  assign n15436 = ~n15431 & n15435;
  assign n15437 = ~n15434 & ~n15436;
  assign n15438 = ~n15259 & ~n15437;
  assign n15439 = ~n15259 & ~n15438;
  assign n15440 = ~n15437 & ~n15438;
  assign n15441 = ~n15439 & ~n15440;
  assign n15442 = ~n15426 & ~n15441;
  assign n15443 = ~n15426 & ~n15442;
  assign n15444 = ~n15441 & ~n15442;
  assign n15445 = ~n15443 & ~n15444;
  assign n15446 = n15415 & ~n15445;
  assign n15447 = n15415 & ~n15446;
  assign n15448 = ~n15445 & ~n15446;
  assign n15449 = ~n15447 & ~n15448;
  assign n15450 = ~n15220 & ~n15223;
  assign n15451 = n15305 & n15319;
  assign n15452 = ~n15305 & ~n15319;
  assign n15453 = ~n15451 & ~n15452;
  assign n15454 = n15271 & ~n15453;
  assign n15455 = ~n15271 & n15453;
  assign n15456 = ~n15454 & ~n15455;
  assign n15457 = ~n15274 & ~n15288;
  assign n15458 = ~n15167 & ~n15307;
  assign n15459 = ~n15322 & ~n15458;
  assign n15460 = n15457 & n15459;
  assign n15461 = ~n15457 & ~n15459;
  assign n15462 = ~n15460 & ~n15461;
  assign n15463 = n15456 & n15462;
  assign n15464 = ~n15456 & ~n15462;
  assign n15465 = ~n15463 & ~n15464;
  assign n15466 = ~n15450 & n15465;
  assign n15467 = n15450 & ~n15465;
  assign n15468 = ~n15466 & ~n15467;
  assign n15469 = n15449 & n15468;
  assign n15470 = ~n15449 & ~n15468;
  assign n15471 = ~n15469 & ~n15470;
  assign n15472 = n15373 & ~n15471;
  assign n15473 = n15373 & ~n15472;
  assign n15474 = ~n15471 & ~n15472;
  assign n15475 = ~n15473 & ~n15474;
  assign n15476 = ~n15227 & ~n15333;
  assign n15477 = ~n15475 & ~n15476;
  assign n15478 = n15475 & n15476;
  assign n15479 = ~n15477 & ~n15478;
  assign n15480 = ~n15337 & ~n15342;
  assign n15481 = ~n15479 & n15480;
  assign n15482 = n15479 & ~n15480;
  assign po96  = ~n15481 & ~n15482;
  assign n15484 = ~n15372 & ~n15472;
  assign n15485 = ~n15414 & ~n15446;
  assign n15486 = pi37  & pi59 ;
  assign n15487 = pi40  & pi56 ;
  assign n15488 = ~n15486 & ~n15487;
  assign n15489 = pi56  & pi59 ;
  assign n15490 = n12266 & n15489;
  assign n15491 = pi36  & pi60 ;
  assign n15492 = ~n15488 & n15491;
  assign n15493 = ~n15490 & n15492;
  assign n15494 = ~n15490 & ~n15493;
  assign n15495 = ~n15488 & n15494;
  assign n15496 = n15491 & ~n15493;
  assign n15497 = ~n15495 & ~n15496;
  assign n15498 = n4736 & n8144;
  assign n15499 = pi38  & pi58 ;
  assign n15500 = pi39  & pi57 ;
  assign n15501 = ~n15499 & ~n15500;
  assign n15502 = n8102 & ~n15498;
  assign n15503 = ~n15501 & n15502;
  assign n15504 = n8102 & ~n15503;
  assign n15505 = ~n15498 & ~n15503;
  assign n15506 = ~n15501 & n15505;
  assign n15507 = ~n15504 & ~n15506;
  assign n15508 = ~n15497 & ~n15507;
  assign n15509 = ~n15497 & ~n15508;
  assign n15510 = ~n15507 & ~n15508;
  assign n15511 = ~n15509 & ~n15510;
  assign n15512 = pi45  & pi51 ;
  assign n15513 = n5277 & n5889;
  assign n15514 = pi46  & pi50 ;
  assign n15515 = ~n8262 & ~n15514;
  assign n15516 = n15512 & ~n15513;
  assign n15517 = ~n15515 & n15516;
  assign n15518 = n15512 & ~n15517;
  assign n15519 = ~n15513 & ~n15517;
  assign n15520 = ~n15515 & n15519;
  assign n15521 = ~n15518 & ~n15520;
  assign n15522 = ~n15511 & ~n15521;
  assign n15523 = ~n15511 & ~n15522;
  assign n15524 = ~n15521 & ~n15522;
  assign n15525 = ~n15523 & ~n15524;
  assign n15526 = ~n15461 & ~n15463;
  assign n15527 = ~n15525 & ~n15526;
  assign n15528 = ~n15525 & ~n15527;
  assign n15529 = ~n15526 & ~n15527;
  assign n15530 = ~n15528 & ~n15529;
  assign n15531 = ~n15485 & ~n15530;
  assign n15532 = ~n15485 & ~n15531;
  assign n15533 = ~n15530 & ~n15531;
  assign n15534 = ~n15532 & ~n15533;
  assign n15535 = ~n15467 & ~n15469;
  assign n15536 = ~n15534 & n15535;
  assign n15537 = ~n15534 & ~n15536;
  assign n15538 = n15535 & ~n15536;
  assign n15539 = ~n15537 & ~n15538;
  assign n15540 = ~n15365 & ~n15368;
  assign n15541 = n15377 & n15391;
  assign n15542 = ~n15377 & ~n15391;
  assign n15543 = ~n15541 & ~n15542;
  assign n15544 = n15405 & ~n15543;
  assign n15545 = ~n15405 & n15543;
  assign n15546 = ~n15544 & ~n15545;
  assign n15547 = ~n15438 & ~n15442;
  assign n15548 = ~n15394 & ~n15408;
  assign n15549 = n15547 & n15548;
  assign n15550 = ~n15547 & ~n15548;
  assign n15551 = ~n15549 & ~n15550;
  assign n15552 = n15546 & n15551;
  assign n15553 = ~n15546 & ~n15551;
  assign n15554 = ~n15552 & ~n15553;
  assign n15555 = ~n15540 & n15554;
  assign n15556 = n15540 & ~n15554;
  assign n15557 = ~n15555 & ~n15556;
  assign n15558 = pi34  & pi62 ;
  assign n15559 = pi35  & pi61 ;
  assign n15560 = ~n15558 & ~n15559;
  assign n15561 = n3106 & n9567;
  assign n15562 = pi33  & pi63 ;
  assign n15563 = ~n15560 & n15562;
  assign n15564 = ~n15561 & n15563;
  assign n15565 = ~n15561 & ~n15564;
  assign n15566 = ~n15560 & n15565;
  assign n15567 = n15562 & ~n15564;
  assign n15568 = ~n15566 & ~n15567;
  assign n15569 = pi41  & pi55 ;
  assign n15570 = n6458 & n8092;
  assign n15571 = pi43  & pi53 ;
  assign n15572 = pi42  & pi54 ;
  assign n15573 = ~n15571 & ~n15572;
  assign n15574 = n15569 & ~n15570;
  assign n15575 = ~n15573 & n15574;
  assign n15576 = n15569 & ~n15575;
  assign n15577 = ~n15570 & ~n15575;
  assign n15578 = ~n15573 & n15577;
  assign n15579 = ~n15576 & ~n15578;
  assign n15580 = ~n15568 & ~n15579;
  assign n15581 = ~n15568 & ~n15580;
  assign n15582 = ~n15579 & ~n15580;
  assign n15583 = ~n15581 & ~n15582;
  assign n15584 = ~n15452 & ~n15455;
  assign n15585 = n15583 & n15584;
  assign n15586 = ~n15583 & ~n15584;
  assign n15587 = ~n15585 & ~n15586;
  assign n15588 = n15423 & n15435;
  assign n15589 = ~n15423 & ~n15435;
  assign n15590 = ~n15588 & ~n15589;
  assign n15591 = ~n15346 & ~n15352;
  assign n15592 = ~n15590 & n15591;
  assign n15593 = n15590 & ~n15591;
  assign n15594 = ~n15592 & ~n15593;
  assign n15595 = ~n15358 & ~n15362;
  assign n15596 = ~n15594 & n15595;
  assign n15597 = n15594 & ~n15595;
  assign n15598 = ~n15596 & ~n15597;
  assign n15599 = n15587 & n15598;
  assign n15600 = ~n15587 & ~n15598;
  assign n15601 = ~n15599 & ~n15600;
  assign n15602 = n15557 & n15601;
  assign n15603 = ~n15557 & ~n15601;
  assign n15604 = ~n15602 & ~n15603;
  assign n15605 = ~n15539 & n15604;
  assign n15606 = n15539 & ~n15604;
  assign n15607 = ~n15605 & ~n15606;
  assign n15608 = n15484 & ~n15607;
  assign n15609 = ~n15484 & n15607;
  assign n15610 = ~n15608 & ~n15609;
  assign n15611 = ~n15477 & ~n15482;
  assign n15612 = ~n15610 & n15611;
  assign n15613 = ~n15608 & ~n15611;
  assign n15614 = ~n15609 & n15613;
  assign po97  = ~n15612 & ~n15614;
  assign n15616 = ~n15609 & ~n15613;
  assign n15617 = ~n15536 & ~n15605;
  assign n15618 = ~n15527 & ~n15531;
  assign n15619 = pi36  & pi61 ;
  assign n15620 = ~n15519 & n15619;
  assign n15621 = n15519 & ~n15619;
  assign n15622 = ~n15620 & ~n15621;
  assign n15623 = n15505 & ~n15622;
  assign n15624 = ~n15505 & n15622;
  assign n15625 = ~n15623 & ~n15624;
  assign n15626 = ~n15508 & ~n15522;
  assign n15627 = ~n15589 & ~n15593;
  assign n15628 = n15626 & n15627;
  assign n15629 = ~n15626 & ~n15627;
  assign n15630 = ~n15628 & ~n15629;
  assign n15631 = n15625 & n15630;
  assign n15632 = ~n15625 & ~n15630;
  assign n15633 = ~n15631 & ~n15632;
  assign n15634 = pi49  & pi62 ;
  assign n15635 = pi35  & n15634;
  assign n15636 = n8505 & ~n15635;
  assign n15637 = ~n15635 & ~n15636;
  assign n15638 = pi35  & pi62 ;
  assign n15639 = ~pi49  & ~n15638;
  assign n15640 = n15637 & ~n15639;
  assign n15641 = n8505 & ~n15636;
  assign n15642 = ~n15640 & ~n15641;
  assign n15643 = pi40  & pi57 ;
  assign n15644 = n5277 & n6114;
  assign n15645 = pi47  & pi50 ;
  assign n15646 = ~n8252 & ~n15645;
  assign n15647 = n15643 & ~n15644;
  assign n15648 = ~n15646 & n15647;
  assign n15649 = n15643 & ~n15648;
  assign n15650 = ~n15644 & ~n15648;
  assign n15651 = ~n15646 & n15650;
  assign n15652 = ~n15649 & ~n15651;
  assign n15653 = ~n15642 & ~n15652;
  assign n15654 = ~n15642 & ~n15653;
  assign n15655 = ~n15652 & ~n15653;
  assign n15656 = ~n15654 & ~n15655;
  assign n15657 = ~n15542 & ~n15545;
  assign n15658 = n15656 & n15657;
  assign n15659 = ~n15656 & ~n15657;
  assign n15660 = ~n15658 & ~n15659;
  assign n15661 = n15494 & n15565;
  assign n15662 = ~n15494 & ~n15565;
  assign n15663 = ~n15661 & ~n15662;
  assign n15664 = n15577 & ~n15663;
  assign n15665 = ~n15577 & n15663;
  assign n15666 = ~n15664 & ~n15665;
  assign n15667 = ~n15580 & ~n15586;
  assign n15668 = ~n15666 & n15667;
  assign n15669 = n15666 & ~n15667;
  assign n15670 = ~n15668 & ~n15669;
  assign n15671 = n15660 & n15670;
  assign n15672 = ~n15660 & ~n15670;
  assign n15673 = ~n15671 & ~n15672;
  assign n15674 = n15633 & n15673;
  assign n15675 = ~n15633 & ~n15673;
  assign n15676 = ~n15674 & ~n15675;
  assign n15677 = n15618 & ~n15676;
  assign n15678 = ~n15618 & n15676;
  assign n15679 = ~n15677 & ~n15678;
  assign n15680 = ~n15597 & ~n15599;
  assign n15681 = pi34  & pi63 ;
  assign n15682 = pi42  & pi55 ;
  assign n15683 = ~n15681 & ~n15682;
  assign n15684 = n15681 & n15682;
  assign n15685 = pi41  & pi56 ;
  assign n15686 = ~n15683 & n15685;
  assign n15687 = ~n15684 & n15686;
  assign n15688 = ~n15684 & ~n15687;
  assign n15689 = ~n15683 & n15688;
  assign n15690 = n15685 & ~n15687;
  assign n15691 = ~n15689 & ~n15690;
  assign n15692 = pi37  & pi60 ;
  assign n15693 = n4736 & n9402;
  assign n15694 = pi38  & pi59 ;
  assign n15695 = pi39  & pi58 ;
  assign n15696 = ~n15694 & ~n15695;
  assign n15697 = n15692 & ~n15693;
  assign n15698 = ~n15696 & n15697;
  assign n15699 = n15692 & ~n15698;
  assign n15700 = ~n15693 & ~n15698;
  assign n15701 = ~n15696 & n15700;
  assign n15702 = ~n15699 & ~n15701;
  assign n15703 = ~n15691 & ~n15702;
  assign n15704 = ~n15691 & ~n15703;
  assign n15705 = ~n15702 & ~n15703;
  assign n15706 = ~n15704 & ~n15705;
  assign n15707 = pi43  & pi54 ;
  assign n15708 = n5318 & n9144;
  assign n15709 = pi44  & pi53 ;
  assign n15710 = ~n8477 & ~n15709;
  assign n15711 = n15707 & ~n15708;
  assign n15712 = ~n15710 & n15711;
  assign n15713 = n15707 & ~n15712;
  assign n15714 = ~n15708 & ~n15712;
  assign n15715 = ~n15710 & n15714;
  assign n15716 = ~n15713 & ~n15715;
  assign n15717 = ~n15706 & ~n15716;
  assign n15718 = ~n15706 & ~n15717;
  assign n15719 = ~n15716 & ~n15717;
  assign n15720 = ~n15718 & ~n15719;
  assign n15721 = ~n15550 & ~n15552;
  assign n15722 = ~n15720 & ~n15721;
  assign n15723 = ~n15720 & ~n15722;
  assign n15724 = ~n15721 & ~n15722;
  assign n15725 = ~n15723 & ~n15724;
  assign n15726 = ~n15680 & ~n15725;
  assign n15727 = ~n15680 & ~n15726;
  assign n15728 = ~n15725 & ~n15726;
  assign n15729 = ~n15727 & ~n15728;
  assign n15730 = ~n15555 & ~n15602;
  assign n15731 = n15729 & n15730;
  assign n15732 = ~n15729 & ~n15730;
  assign n15733 = ~n15731 & ~n15732;
  assign n15734 = n15679 & n15733;
  assign n15735 = ~n15679 & ~n15733;
  assign n15736 = ~n15734 & ~n15735;
  assign n15737 = ~n15617 & n15736;
  assign n15738 = n15617 & ~n15736;
  assign n15739 = ~n15737 & ~n15738;
  assign n15740 = ~n15616 & ~n15739;
  assign n15741 = n15616 & n15739;
  assign po98  = n15740 | n15741;
  assign n15743 = ~n15732 & ~n15734;
  assign n15744 = ~n15722 & ~n15726;
  assign n15745 = ~n15662 & ~n15665;
  assign n15746 = ~n15620 & ~n15624;
  assign n15747 = n15745 & n15746;
  assign n15748 = ~n15745 & ~n15746;
  assign n15749 = ~n15747 & ~n15748;
  assign n15750 = ~n15703 & ~n15717;
  assign n15751 = ~n15749 & n15750;
  assign n15752 = n15749 & ~n15750;
  assign n15753 = ~n15751 & ~n15752;
  assign n15754 = n15688 & n15700;
  assign n15755 = ~n15688 & ~n15700;
  assign n15756 = ~n15754 & ~n15755;
  assign n15757 = n15714 & ~n15756;
  assign n15758 = ~n15714 & n15756;
  assign n15759 = ~n15757 & ~n15758;
  assign n15760 = ~n15653 & ~n15659;
  assign n15761 = ~n15759 & n15760;
  assign n15762 = n15759 & ~n15760;
  assign n15763 = ~n15761 & ~n15762;
  assign n15764 = pi39  & pi59 ;
  assign n15765 = pi40  & pi58 ;
  assign n15766 = ~n15764 & ~n15765;
  assign n15767 = n5548 & n9402;
  assign n15768 = pi45  & pi53 ;
  assign n15769 = ~n15766 & n15768;
  assign n15770 = ~n15767 & n15769;
  assign n15771 = ~n15767 & ~n15770;
  assign n15772 = ~n15766 & n15771;
  assign n15773 = n15768 & ~n15770;
  assign n15774 = ~n15772 & ~n15773;
  assign n15775 = pi46  & pi52 ;
  assign n15776 = n5823 & n6114;
  assign n15777 = ~n5481 & ~n8495;
  assign n15778 = n15775 & ~n15776;
  assign n15779 = ~n15777 & n15778;
  assign n15780 = n15775 & ~n15779;
  assign n15781 = ~n15776 & ~n15779;
  assign n15782 = ~n15777 & n15781;
  assign n15783 = ~n15780 & ~n15782;
  assign n15784 = ~n15774 & ~n15783;
  assign n15785 = ~n15774 & ~n15784;
  assign n15786 = ~n15783 & ~n15784;
  assign n15787 = ~n15785 & ~n15786;
  assign n15788 = n4500 & n9567;
  assign n15789 = pi37  & pi61 ;
  assign n15790 = ~n10816 & ~n15789;
  assign n15791 = ~n15788 & ~n15790;
  assign n15792 = ~n15637 & n15791;
  assign n15793 = n15637 & ~n15791;
  assign n15794 = ~n15792 & ~n15793;
  assign n15795 = n15787 & n15794;
  assign n15796 = ~n15787 & ~n15794;
  assign n15797 = ~n15795 & ~n15796;
  assign n15798 = n15763 & ~n15797;
  assign n15799 = n15763 & ~n15798;
  assign n15800 = ~n15797 & ~n15798;
  assign n15801 = ~n15799 & ~n15800;
  assign n15802 = n15753 & ~n15801;
  assign n15803 = ~n15753 & n15801;
  assign n15804 = ~n15802 & ~n15803;
  assign n15805 = ~n15744 & n15804;
  assign n15806 = ~n15744 & ~n15805;
  assign n15807 = ~n15802 & ~n15805;
  assign n15808 = ~n15803 & n15807;
  assign n15809 = ~n15806 & ~n15808;
  assign n15810 = ~n15674 & ~n15678;
  assign n15811 = ~n15669 & ~n15671;
  assign n15812 = n6836 & n9891;
  assign n15813 = pi43  & pi55 ;
  assign n15814 = pi44  & pi54 ;
  assign n15815 = ~n15813 & ~n15814;
  assign n15816 = ~n15812 & ~n15815;
  assign n15817 = pi35  & pi63 ;
  assign n15818 = ~n15816 & ~n15817;
  assign n15819 = n15816 & n15817;
  assign n15820 = ~n15818 & ~n15819;
  assign n15821 = ~n15650 & n15820;
  assign n15822 = n15650 & ~n15820;
  assign n15823 = ~n15821 & ~n15822;
  assign n15824 = pi38  & pi60 ;
  assign n15825 = n5235 & n7643;
  assign n15826 = pi41  & pi57 ;
  assign n15827 = pi42  & pi56 ;
  assign n15828 = ~n15826 & ~n15827;
  assign n15829 = n15824 & ~n15825;
  assign n15830 = ~n15828 & n15829;
  assign n15831 = n15824 & ~n15830;
  assign n15832 = ~n15825 & ~n15830;
  assign n15833 = ~n15828 & n15832;
  assign n15834 = ~n15831 & ~n15833;
  assign n15835 = n15823 & ~n15834;
  assign n15836 = n15823 & ~n15835;
  assign n15837 = ~n15834 & ~n15835;
  assign n15838 = ~n15836 & ~n15837;
  assign n15839 = ~n15629 & ~n15631;
  assign n15840 = ~n15838 & ~n15839;
  assign n15841 = ~n15838 & ~n15840;
  assign n15842 = ~n15839 & ~n15840;
  assign n15843 = ~n15841 & ~n15842;
  assign n15844 = ~n15811 & ~n15843;
  assign n15845 = n15811 & n15843;
  assign n15846 = ~n15844 & ~n15845;
  assign n15847 = ~n15810 & n15846;
  assign n15848 = ~n15810 & ~n15847;
  assign n15849 = n15846 & ~n15847;
  assign n15850 = ~n15848 & ~n15849;
  assign n15851 = ~n15809 & ~n15850;
  assign n15852 = n15809 & n15850;
  assign n15853 = ~n15851 & ~n15852;
  assign n15854 = n15743 & ~n15853;
  assign n15855 = ~n15743 & n15853;
  assign n15856 = ~n15854 & ~n15855;
  assign n15857 = ~n15616 & ~n15738;
  assign n15858 = ~n15737 & ~n15857;
  assign n15859 = ~n15856 & n15858;
  assign n15860 = n15856 & ~n15858;
  assign po99  = ~n15859 & ~n15860;
  assign n15862 = ~n15847 & ~n15851;
  assign n15863 = ~n15840 & ~n15844;
  assign n15864 = ~n15755 & ~n15758;
  assign n15865 = pi50  & pi62 ;
  assign n15866 = pi37  & n15865;
  assign n15867 = n5889 & ~n15866;
  assign n15868 = n5889 & ~n15867;
  assign n15869 = ~n15866 & ~n15867;
  assign n15870 = pi37  & pi62 ;
  assign n15871 = ~pi50  & ~n15870;
  assign n15872 = n15869 & ~n15871;
  assign n15873 = ~n15868 & ~n15872;
  assign n15874 = ~n15864 & ~n15873;
  assign n15875 = ~n15864 & ~n15874;
  assign n15876 = ~n15873 & ~n15874;
  assign n15877 = ~n15875 & ~n15876;
  assign n15878 = ~n15821 & ~n15835;
  assign n15879 = n15877 & n15878;
  assign n15880 = ~n15877 & ~n15878;
  assign n15881 = ~n15879 & ~n15880;
  assign n15882 = ~n15788 & ~n15792;
  assign n15883 = n15832 & n15882;
  assign n15884 = ~n15832 & ~n15882;
  assign n15885 = ~n15883 & ~n15884;
  assign n15886 = pi36  & pi63 ;
  assign n15887 = n4736 & n9054;
  assign n15888 = pi38  & pi61 ;
  assign n15889 = pi39  & pi60 ;
  assign n15890 = ~n15888 & ~n15889;
  assign n15891 = n15886 & ~n15887;
  assign n15892 = ~n15890 & n15891;
  assign n15893 = n15886 & ~n15892;
  assign n15894 = ~n15887 & ~n15892;
  assign n15895 = ~n15890 & n15894;
  assign n15896 = ~n15893 & ~n15895;
  assign n15897 = n15885 & ~n15896;
  assign n15898 = n15885 & ~n15897;
  assign n15899 = ~n15896 & ~n15897;
  assign n15900 = ~n15898 & ~n15899;
  assign n15901 = n15771 & n15781;
  assign n15902 = ~n15771 & ~n15781;
  assign n15903 = ~n15901 & ~n15902;
  assign n15904 = ~n15812 & ~n15819;
  assign n15905 = ~n15903 & n15904;
  assign n15906 = n15903 & ~n15904;
  assign n15907 = ~n15905 & ~n15906;
  assign n15908 = ~n15787 & n15794;
  assign n15909 = ~n15784 & ~n15908;
  assign n15910 = n15907 & ~n15909;
  assign n15911 = ~n15907 & n15909;
  assign n15912 = ~n15910 & ~n15911;
  assign n15913 = ~n15900 & ~n15912;
  assign n15914 = n15900 & n15912;
  assign n15915 = ~n15913 & ~n15914;
  assign n15916 = n15881 & ~n15915;
  assign n15917 = ~n15881 & n15915;
  assign n15918 = ~n15916 & ~n15917;
  assign n15919 = ~n15863 & n15918;
  assign n15920 = n15863 & ~n15918;
  assign n15921 = ~n15919 & ~n15920;
  assign n15922 = pi41  & pi58 ;
  assign n15923 = ~n8838 & ~n15922;
  assign n15924 = n8838 & n15922;
  assign n15925 = pi40  & pi59 ;
  assign n15926 = ~n15923 & n15925;
  assign n15927 = ~n15924 & n15926;
  assign n15928 = ~n15924 & ~n15927;
  assign n15929 = ~n15923 & n15928;
  assign n15930 = n15925 & ~n15927;
  assign n15931 = ~n15929 & ~n15930;
  assign n15932 = pi45  & pi54 ;
  assign n15933 = n5277 & n9144;
  assign n15934 = pi46  & pi53 ;
  assign n15935 = ~n8783 & ~n15934;
  assign n15936 = n15932 & ~n15933;
  assign n15937 = ~n15935 & n15936;
  assign n15938 = n15932 & ~n15937;
  assign n15939 = ~n15933 & ~n15937;
  assign n15940 = ~n15935 & n15939;
  assign n15941 = ~n15938 & ~n15940;
  assign n15942 = ~n15931 & ~n15941;
  assign n15943 = ~n15931 & ~n15942;
  assign n15944 = ~n15941 & ~n15942;
  assign n15945 = ~n15943 & ~n15944;
  assign n15946 = pi48  & pi51 ;
  assign n15947 = n6458 & n7643;
  assign n15948 = pi42  & pi57 ;
  assign n15949 = pi43  & pi56 ;
  assign n15950 = ~n15948 & ~n15949;
  assign n15951 = n15946 & ~n15947;
  assign n15952 = ~n15950 & n15951;
  assign n15953 = n15946 & ~n15952;
  assign n15954 = ~n15947 & ~n15952;
  assign n15955 = ~n15950 & n15954;
  assign n15956 = ~n15953 & ~n15955;
  assign n15957 = ~n15945 & ~n15956;
  assign n15958 = ~n15945 & ~n15957;
  assign n15959 = ~n15956 & ~n15957;
  assign n15960 = ~n15958 & ~n15959;
  assign n15961 = ~n15748 & ~n15752;
  assign n15962 = n15960 & n15961;
  assign n15963 = ~n15960 & ~n15961;
  assign n15964 = ~n15962 & ~n15963;
  assign n15965 = ~n15762 & ~n15798;
  assign n15966 = ~n15964 & n15965;
  assign n15967 = n15964 & ~n15965;
  assign n15968 = ~n15966 & ~n15967;
  assign n15969 = ~n15807 & n15968;
  assign n15970 = n15968 & ~n15969;
  assign n15971 = ~n15807 & ~n15969;
  assign n15972 = ~n15970 & ~n15971;
  assign n15973 = n15921 & ~n15972;
  assign n15974 = ~n15921 & n15972;
  assign n15975 = ~n15973 & ~n15974;
  assign n15976 = ~n15862 & n15975;
  assign n15977 = n15862 & ~n15975;
  assign n15978 = ~n15976 & ~n15977;
  assign n15979 = ~n15855 & ~n15860;
  assign n15980 = ~n15978 & n15979;
  assign n15981 = n15978 & ~n15979;
  assign po100  = ~n15980 & ~n15981;
  assign n15983 = ~n15969 & ~n15973;
  assign n15984 = ~n15902 & ~n15906;
  assign n15985 = pi47  & pi53 ;
  assign n15986 = n8505 & n10319;
  assign n15987 = pi49  & pi51 ;
  assign n15988 = pi48  & pi52 ;
  assign n15989 = ~n15987 & ~n15988;
  assign n15990 = n15985 & ~n15986;
  assign n15991 = ~n15989 & n15990;
  assign n15992 = n15985 & ~n15991;
  assign n15993 = ~n15986 & ~n15991;
  assign n15994 = ~n15989 & n15993;
  assign n15995 = ~n15992 & ~n15994;
  assign n15996 = ~n15984 & ~n15995;
  assign n15997 = ~n15984 & ~n15996;
  assign n15998 = ~n15995 & ~n15996;
  assign n15999 = ~n15997 & ~n15998;
  assign n16000 = ~n15884 & ~n15897;
  assign n16001 = n15999 & n16000;
  assign n16002 = ~n15999 & ~n16000;
  assign n16003 = ~n16001 & ~n16002;
  assign n16004 = ~n15963 & ~n15967;
  assign n16005 = ~n16003 & n16004;
  assign n16006 = n16003 & ~n16004;
  assign n16007 = ~n16005 & ~n16006;
  assign n16008 = n15894 & n15939;
  assign n16009 = ~n15894 & ~n15939;
  assign n16010 = ~n16008 & ~n16009;
  assign n16011 = n15928 & ~n16010;
  assign n16012 = ~n15928 & n16010;
  assign n16013 = ~n16011 & ~n16012;
  assign n16014 = ~n15942 & ~n15957;
  assign n16015 = ~n16013 & n16014;
  assign n16016 = n16013 & ~n16014;
  assign n16017 = ~n16015 & ~n16016;
  assign n16018 = pi37  & pi63 ;
  assign n16019 = ~n15869 & n16018;
  assign n16020 = n15869 & ~n16018;
  assign n16021 = ~n16019 & ~n16020;
  assign n16022 = n15954 & ~n16021;
  assign n16023 = ~n15954 & n16021;
  assign n16024 = ~n16022 & ~n16023;
  assign n16025 = n16017 & n16024;
  assign n16026 = ~n16017 & ~n16024;
  assign n16027 = ~n16025 & ~n16026;
  assign n16028 = n16007 & n16027;
  assign n16029 = ~n16007 & ~n16027;
  assign n16030 = ~n16028 & ~n16029;
  assign n16031 = ~n15916 & ~n15919;
  assign n16032 = pi40  & pi60 ;
  assign n16033 = pi39  & pi61 ;
  assign n16034 = ~n16032 & ~n16033;
  assign n16035 = n5548 & n9054;
  assign n16036 = n11769 & ~n16034;
  assign n16037 = ~n16035 & n16036;
  assign n16038 = ~n16035 & ~n16037;
  assign n16039 = ~n16034 & n16038;
  assign n16040 = n11769 & ~n16037;
  assign n16041 = ~n16039 & ~n16040;
  assign n16042 = pi43  & pi57 ;
  assign n16043 = n5318 & n8521;
  assign n16044 = pi44  & pi56 ;
  assign n16045 = ~n15151 & ~n16044;
  assign n16046 = n16042 & ~n16043;
  assign n16047 = ~n16045 & n16046;
  assign n16048 = n16042 & ~n16047;
  assign n16049 = ~n16043 & ~n16047;
  assign n16050 = ~n16045 & n16049;
  assign n16051 = ~n16048 & ~n16050;
  assign n16052 = ~n16041 & ~n16051;
  assign n16053 = ~n16041 & ~n16052;
  assign n16054 = ~n16051 & ~n16052;
  assign n16055 = ~n16053 & ~n16054;
  assign n16056 = n5235 & n9402;
  assign n16057 = pi41  & pi59 ;
  assign n16058 = pi42  & pi58 ;
  assign n16059 = ~n16057 & ~n16058;
  assign n16060 = n8773 & ~n16056;
  assign n16061 = ~n16059 & n16060;
  assign n16062 = n8773 & ~n16061;
  assign n16063 = ~n16056 & ~n16061;
  assign n16064 = ~n16059 & n16063;
  assign n16065 = ~n16062 & ~n16064;
  assign n16066 = ~n16055 & ~n16065;
  assign n16067 = ~n16055 & ~n16066;
  assign n16068 = ~n16065 & ~n16066;
  assign n16069 = ~n16067 & ~n16068;
  assign n16070 = ~n15874 & ~n15880;
  assign n16071 = n16069 & n16070;
  assign n16072 = ~n16069 & ~n16070;
  assign n16073 = ~n16071 & ~n16072;
  assign n16074 = ~n15911 & ~n15914;
  assign n16075 = n16073 & n16074;
  assign n16076 = ~n16073 & ~n16074;
  assign n16077 = ~n16075 & ~n16076;
  assign n16078 = ~n16031 & n16077;
  assign n16079 = n16031 & ~n16077;
  assign n16080 = ~n16078 & ~n16079;
  assign n16081 = n16030 & n16080;
  assign n16082 = ~n16030 & ~n16080;
  assign n16083 = ~n16081 & ~n16082;
  assign n16084 = ~n15983 & n16083;
  assign n16085 = n15983 & ~n16083;
  assign n16086 = ~n16084 & ~n16085;
  assign n16087 = ~n15976 & ~n15981;
  assign n16088 = ~n16086 & n16087;
  assign n16089 = ~n16085 & ~n16087;
  assign n16090 = ~n16084 & n16089;
  assign po101  = ~n16088 & ~n16090;
  assign n16092 = ~n16084 & ~n16089;
  assign n16093 = ~n16078 & ~n16081;
  assign n16094 = ~n16006 & ~n16028;
  assign n16095 = pi46  & pi55 ;
  assign n16096 = pi47  & pi54 ;
  assign n16097 = ~n16095 & ~n16096;
  assign n16098 = n5277 & n9891;
  assign n16099 = pi38  & pi63 ;
  assign n16100 = ~n16097 & n16099;
  assign n16101 = ~n16098 & n16100;
  assign n16102 = ~n16098 & ~n16101;
  assign n16103 = ~n16097 & n16102;
  assign n16104 = n16099 & ~n16101;
  assign n16105 = ~n16103 & ~n16104;
  assign n16106 = pi42  & pi59 ;
  assign n16107 = n12970 & n14390;
  assign n16108 = pi43  & pi58 ;
  assign n16109 = pi45  & pi56 ;
  assign n16110 = ~n16108 & ~n16109;
  assign n16111 = n16106 & ~n16107;
  assign n16112 = ~n16110 & n16111;
  assign n16113 = n16106 & ~n16112;
  assign n16114 = ~n16107 & ~n16112;
  assign n16115 = ~n16110 & n16114;
  assign n16116 = ~n16113 & ~n16115;
  assign n16117 = ~n16105 & ~n16116;
  assign n16118 = ~n16105 & ~n16117;
  assign n16119 = ~n16116 & ~n16117;
  assign n16120 = ~n16118 & ~n16119;
  assign n16121 = pi48  & pi53 ;
  assign n16122 = n8102 & n11798;
  assign n16123 = pi44  & pi57 ;
  assign n16124 = pi49  & pi52 ;
  assign n16125 = ~n16123 & ~n16124;
  assign n16126 = n16121 & ~n16122;
  assign n16127 = ~n16125 & n16126;
  assign n16128 = n16121 & ~n16127;
  assign n16129 = ~n16122 & ~n16127;
  assign n16130 = ~n16125 & n16129;
  assign n16131 = ~n16128 & ~n16130;
  assign n16132 = ~n16120 & ~n16131;
  assign n16133 = ~n16120 & ~n16132;
  assign n16134 = ~n16131 & ~n16132;
  assign n16135 = ~n16133 & ~n16134;
  assign n16136 = ~n15996 & ~n16002;
  assign n16137 = n16135 & n16136;
  assign n16138 = ~n16135 & ~n16136;
  assign n16139 = ~n16137 & ~n16138;
  assign n16140 = ~n16019 & ~n16023;
  assign n16141 = n6012 & n9054;
  assign n16142 = pi41  & pi60 ;
  assign n16143 = ~n16141 & n16142;
  assign n16144 = pi40  & pi61 ;
  assign n16145 = ~n16141 & n16144;
  assign n16146 = ~n16143 & ~n16145;
  assign n16147 = ~n15993 & ~n16146;
  assign n16148 = ~n15993 & ~n16147;
  assign n16149 = ~n16146 & ~n16147;
  assign n16150 = ~n16148 & ~n16149;
  assign n16151 = pi62  & n14685;
  assign n16152 = n6114 & ~n16151;
  assign n16153 = ~n16151 & ~n16152;
  assign n16154 = pi39  & pi62 ;
  assign n16155 = ~pi51  & ~n16154;
  assign n16156 = n16153 & ~n16155;
  assign n16157 = n6114 & ~n16152;
  assign n16158 = ~n16156 & ~n16157;
  assign n16159 = ~n16150 & ~n16158;
  assign n16160 = ~n16150 & ~n16159;
  assign n16161 = ~n16158 & ~n16159;
  assign n16162 = ~n16160 & ~n16161;
  assign n16163 = ~n16140 & ~n16162;
  assign n16164 = ~n16140 & ~n16163;
  assign n16165 = ~n16162 & ~n16163;
  assign n16166 = ~n16164 & ~n16165;
  assign n16167 = n16139 & ~n16166;
  assign n16168 = ~n16139 & n16166;
  assign n16169 = ~n16167 & ~n16168;
  assign n16170 = ~n16094 & n16169;
  assign n16171 = ~n16094 & ~n16170;
  assign n16172 = n16169 & ~n16170;
  assign n16173 = ~n16171 & ~n16172;
  assign n16174 = ~n16072 & ~n16075;
  assign n16175 = ~n16016 & ~n16025;
  assign n16176 = ~n16174 & ~n16175;
  assign n16177 = ~n16174 & ~n16176;
  assign n16178 = ~n16175 & ~n16176;
  assign n16179 = ~n16177 & ~n16178;
  assign n16180 = n16038 & n16063;
  assign n16181 = ~n16038 & ~n16063;
  assign n16182 = ~n16180 & ~n16181;
  assign n16183 = n16049 & ~n16182;
  assign n16184 = ~n16049 & n16182;
  assign n16185 = ~n16183 & ~n16184;
  assign n16186 = ~n16052 & ~n16066;
  assign n16187 = ~n16009 & ~n16012;
  assign n16188 = n16186 & n16187;
  assign n16189 = ~n16186 & ~n16187;
  assign n16190 = ~n16188 & ~n16189;
  assign n16191 = n16185 & n16190;
  assign n16192 = ~n16185 & ~n16190;
  assign n16193 = ~n16191 & ~n16192;
  assign n16194 = ~n16179 & n16193;
  assign n16195 = ~n16179 & ~n16194;
  assign n16196 = n16193 & ~n16194;
  assign n16197 = ~n16195 & ~n16196;
  assign n16198 = ~n16173 & n16197;
  assign n16199 = n16173 & ~n16197;
  assign n16200 = ~n16198 & ~n16199;
  assign n16201 = ~n16093 & ~n16200;
  assign n16202 = n16093 & n16200;
  assign n16203 = ~n16201 & ~n16202;
  assign n16204 = ~n16092 & ~n16203;
  assign n16205 = n16092 & n16203;
  assign po102  = n16204 | n16205;
  assign n16207 = ~n16092 & ~n16202;
  assign n16208 = ~n16201 & ~n16207;
  assign n16209 = ~n16173 & ~n16197;
  assign n16210 = ~n16170 & ~n16209;
  assign n16211 = ~n16176 & ~n16194;
  assign n16212 = ~n16141 & ~n16147;
  assign n16213 = n16114 & n16212;
  assign n16214 = ~n16114 & ~n16212;
  assign n16215 = ~n16213 & ~n16214;
  assign n16216 = pi39  & pi63 ;
  assign n16217 = n5235 & n9054;
  assign n16218 = pi41  & pi61 ;
  assign n16219 = pi42  & pi60 ;
  assign n16220 = ~n16218 & ~n16219;
  assign n16221 = n16216 & ~n16217;
  assign n16222 = ~n16220 & n16221;
  assign n16223 = n16216 & ~n16222;
  assign n16224 = ~n16217 & ~n16222;
  assign n16225 = ~n16220 & n16224;
  assign n16226 = ~n16223 & ~n16225;
  assign n16227 = n16215 & ~n16226;
  assign n16228 = n16215 & ~n16227;
  assign n16229 = ~n16226 & ~n16227;
  assign n16230 = ~n16228 & ~n16229;
  assign n16231 = ~n16159 & ~n16163;
  assign n16232 = n16230 & n16231;
  assign n16233 = ~n16230 & ~n16231;
  assign n16234 = ~n16232 & ~n16233;
  assign n16235 = pi43  & pi59 ;
  assign n16236 = pi44  & pi58 ;
  assign n16237 = ~n16235 & ~n16236;
  assign n16238 = n6836 & n9402;
  assign n16239 = n12661 & ~n16237;
  assign n16240 = ~n16238 & n16239;
  assign n16241 = ~n16238 & ~n16240;
  assign n16242 = ~n16237 & n16241;
  assign n16243 = n12661 & ~n16240;
  assign n16244 = ~n16242 & ~n16243;
  assign n16245 = pi45  & pi57 ;
  assign n16246 = n5277 & n8521;
  assign n16247 = pi46  & pi56 ;
  assign n16248 = pi47  & pi55 ;
  assign n16249 = ~n16247 & ~n16248;
  assign n16250 = n16245 & ~n16246;
  assign n16251 = ~n16249 & n16250;
  assign n16252 = n16245 & ~n16251;
  assign n16253 = ~n16246 & ~n16251;
  assign n16254 = ~n16249 & n16253;
  assign n16255 = ~n16252 & ~n16254;
  assign n16256 = ~n16244 & ~n16255;
  assign n16257 = ~n16244 & ~n16256;
  assign n16258 = ~n16255 & ~n16256;
  assign n16259 = ~n16257 & ~n16258;
  assign n16260 = pi48  & pi54 ;
  assign n16261 = n5889 & n9144;
  assign n16262 = pi50  & pi52 ;
  assign n16263 = pi49  & pi53 ;
  assign n16264 = ~n16262 & ~n16263;
  assign n16265 = n16260 & ~n16261;
  assign n16266 = ~n16264 & n16265;
  assign n16267 = n16260 & ~n16266;
  assign n16268 = ~n16261 & ~n16266;
  assign n16269 = ~n16264 & n16268;
  assign n16270 = ~n16267 & ~n16269;
  assign n16271 = ~n16259 & ~n16270;
  assign n16272 = ~n16259 & ~n16271;
  assign n16273 = ~n16270 & ~n16271;
  assign n16274 = ~n16272 & ~n16273;
  assign n16275 = n16234 & ~n16274;
  assign n16276 = ~n16234 & n16274;
  assign n16277 = ~n16275 & ~n16276;
  assign n16278 = ~n16211 & n16277;
  assign n16279 = ~n16211 & ~n16278;
  assign n16280 = n16277 & ~n16278;
  assign n16281 = ~n16279 & ~n16280;
  assign n16282 = n16129 & n16153;
  assign n16283 = ~n16129 & ~n16153;
  assign n16284 = ~n16282 & ~n16283;
  assign n16285 = n16102 & ~n16284;
  assign n16286 = ~n16102 & n16284;
  assign n16287 = ~n16285 & ~n16286;
  assign n16288 = ~n16181 & ~n16184;
  assign n16289 = ~n16287 & n16288;
  assign n16290 = n16287 & ~n16288;
  assign n16291 = ~n16289 & ~n16290;
  assign n16292 = ~n16117 & ~n16132;
  assign n16293 = ~n16291 & n16292;
  assign n16294 = n16291 & ~n16292;
  assign n16295 = ~n16293 & ~n16294;
  assign n16296 = ~n16138 & ~n16167;
  assign n16297 = ~n16189 & ~n16191;
  assign n16298 = ~n16296 & ~n16297;
  assign n16299 = ~n16296 & ~n16298;
  assign n16300 = ~n16297 & ~n16298;
  assign n16301 = ~n16299 & ~n16300;
  assign n16302 = n16295 & ~n16301;
  assign n16303 = ~n16295 & n16301;
  assign n16304 = ~n16302 & ~n16303;
  assign n16305 = ~n16281 & n16304;
  assign n16306 = ~n16281 & ~n16305;
  assign n16307 = n16304 & ~n16305;
  assign n16308 = ~n16306 & ~n16307;
  assign n16309 = n16210 & n16308;
  assign n16310 = ~n16210 & ~n16308;
  assign n16311 = ~n16309 & ~n16310;
  assign n16312 = n16208 & ~n16311;
  assign n16313 = ~n16208 & ~n16309;
  assign n16314 = ~n16310 & n16313;
  assign po103  = ~n16312 & ~n16314;
  assign n16316 = ~n16310 & ~n16313;
  assign n16317 = ~n16298 & ~n16302;
  assign n16318 = pi46  & pi57 ;
  assign n16319 = pi47  & pi56 ;
  assign n16320 = ~n16318 & ~n16319;
  assign n16321 = n5277 & n7643;
  assign n16322 = pi43  & pi60 ;
  assign n16323 = ~n16320 & n16322;
  assign n16324 = ~n16321 & n16323;
  assign n16325 = ~n16321 & ~n16324;
  assign n16326 = ~n16320 & n16325;
  assign n16327 = n16322 & ~n16324;
  assign n16328 = ~n16326 & ~n16327;
  assign n16329 = pi48  & pi55 ;
  assign n16330 = n5889 & n8092;
  assign n16331 = pi50  & pi53 ;
  assign n16332 = ~n11314 & ~n16331;
  assign n16333 = n16329 & ~n16330;
  assign n16334 = ~n16332 & n16333;
  assign n16335 = n16329 & ~n16334;
  assign n16336 = ~n16330 & ~n16334;
  assign n16337 = ~n16332 & n16336;
  assign n16338 = ~n16335 & ~n16337;
  assign n16339 = ~n16328 & ~n16338;
  assign n16340 = ~n16328 & ~n16339;
  assign n16341 = ~n16338 & ~n16339;
  assign n16342 = ~n16340 & ~n16341;
  assign n16343 = pi52  & n12960;
  assign n16344 = n10319 & ~n16343;
  assign n16345 = n10319 & ~n16344;
  assign n16346 = ~n16343 & ~n16344;
  assign n16347 = ~pi52  & ~n12960;
  assign n16348 = n16346 & ~n16347;
  assign n16349 = ~n16345 & ~n16348;
  assign n16350 = ~n16342 & ~n16349;
  assign n16351 = ~n16342 & ~n16350;
  assign n16352 = ~n16349 & ~n16350;
  assign n16353 = ~n16351 & ~n16352;
  assign n16354 = pi40  & pi63 ;
  assign n16355 = ~n16268 & n16354;
  assign n16356 = n16268 & ~n16354;
  assign n16357 = ~n16355 & ~n16356;
  assign n16358 = n16253 & ~n16357;
  assign n16359 = ~n16253 & n16357;
  assign n16360 = ~n16358 & ~n16359;
  assign n16361 = n16224 & n16241;
  assign n16362 = ~n16224 & ~n16241;
  assign n16363 = ~n16361 & ~n16362;
  assign n16364 = pi42  & pi61 ;
  assign n16365 = n5318 & n9402;
  assign n16366 = pi44  & pi59 ;
  assign n16367 = pi45  & pi58 ;
  assign n16368 = ~n16366 & ~n16367;
  assign n16369 = n16364 & ~n16365;
  assign n16370 = ~n16368 & n16369;
  assign n16371 = n16364 & ~n16370;
  assign n16372 = ~n16365 & ~n16370;
  assign n16373 = ~n16368 & n16372;
  assign n16374 = ~n16371 & ~n16373;
  assign n16375 = n16363 & ~n16374;
  assign n16376 = n16363 & ~n16375;
  assign n16377 = ~n16374 & ~n16375;
  assign n16378 = ~n16376 & ~n16377;
  assign n16379 = ~n16360 & n16378;
  assign n16380 = n16360 & ~n16378;
  assign n16381 = ~n16379 & ~n16380;
  assign n16382 = ~n16353 & n16381;
  assign n16383 = ~n16353 & ~n16382;
  assign n16384 = n16381 & ~n16382;
  assign n16385 = ~n16383 & ~n16384;
  assign n16386 = ~n16317 & ~n16385;
  assign n16387 = ~n16317 & ~n16386;
  assign n16388 = ~n16385 & ~n16386;
  assign n16389 = ~n16387 & ~n16388;
  assign n16390 = ~n16214 & ~n16227;
  assign n16391 = ~n16283 & ~n16286;
  assign n16392 = n16390 & n16391;
  assign n16393 = ~n16390 & ~n16391;
  assign n16394 = ~n16392 & ~n16393;
  assign n16395 = ~n16256 & ~n16271;
  assign n16396 = ~n16394 & n16395;
  assign n16397 = n16394 & ~n16395;
  assign n16398 = ~n16396 & ~n16397;
  assign n16399 = ~n16233 & ~n16275;
  assign n16400 = ~n16290 & ~n16294;
  assign n16401 = n16399 & n16400;
  assign n16402 = ~n16399 & ~n16400;
  assign n16403 = ~n16401 & ~n16402;
  assign n16404 = n16398 & n16403;
  assign n16405 = ~n16398 & ~n16403;
  assign n16406 = ~n16404 & ~n16405;
  assign n16407 = ~n16389 & n16406;
  assign n16408 = ~n16389 & ~n16407;
  assign n16409 = n16406 & ~n16407;
  assign n16410 = ~n16408 & ~n16409;
  assign n16411 = ~n16278 & ~n16305;
  assign n16412 = ~n16410 & ~n16411;
  assign n16413 = n16410 & n16411;
  assign n16414 = ~n16412 & ~n16413;
  assign n16415 = ~n16316 & ~n16414;
  assign n16416 = n16316 & n16414;
  assign po104  = n16415 | n16416;
  assign n16418 = ~n16316 & ~n16413;
  assign n16419 = ~n16412 & ~n16418;
  assign n16420 = ~n16386 & ~n16407;
  assign n16421 = ~n16402 & ~n16404;
  assign n16422 = n16325 & n16336;
  assign n16423 = ~n16325 & ~n16336;
  assign n16424 = ~n16422 & ~n16423;
  assign n16425 = n16372 & ~n16424;
  assign n16426 = ~n16372 & n16424;
  assign n16427 = ~n16425 & ~n16426;
  assign n16428 = ~n16339 & ~n16350;
  assign n16429 = ~n16427 & n16428;
  assign n16430 = n16427 & ~n16428;
  assign n16431 = ~n16429 & ~n16430;
  assign n16432 = pi43  & pi61 ;
  assign n16433 = pi45  & pi59 ;
  assign n16434 = ~n16432 & ~n16433;
  assign n16435 = n14390 & n15297;
  assign n16436 = pi44  & pi60 ;
  assign n16437 = ~n16434 & n16436;
  assign n16438 = ~n16435 & n16437;
  assign n16439 = ~n16435 & ~n16438;
  assign n16440 = ~n16434 & n16439;
  assign n16441 = n16436 & ~n16438;
  assign n16442 = ~n16440 & ~n16441;
  assign n16443 = pi46  & pi58 ;
  assign n16444 = n5823 & n7643;
  assign n16445 = pi47  & pi57 ;
  assign n16446 = ~n9000 & ~n16445;
  assign n16447 = n16443 & ~n16444;
  assign n16448 = ~n16446 & n16447;
  assign n16449 = n16443 & ~n16448;
  assign n16450 = ~n16444 & ~n16448;
  assign n16451 = ~n16446 & n16450;
  assign n16452 = ~n16449 & ~n16451;
  assign n16453 = ~n16442 & ~n16452;
  assign n16454 = ~n16442 & ~n16453;
  assign n16455 = ~n16452 & ~n16453;
  assign n16456 = ~n16454 & ~n16455;
  assign n16457 = pi49  & pi55 ;
  assign n16458 = n6114 & n8092;
  assign n16459 = pi50  & pi54 ;
  assign n16460 = ~n6765 & ~n16459;
  assign n16461 = n16457 & ~n16458;
  assign n16462 = ~n16460 & n16461;
  assign n16463 = n16457 & ~n16462;
  assign n16464 = ~n16458 & ~n16462;
  assign n16465 = ~n16460 & n16464;
  assign n16466 = ~n16463 & ~n16465;
  assign n16467 = ~n16456 & ~n16466;
  assign n16468 = ~n16456 & ~n16467;
  assign n16469 = ~n16466 & ~n16467;
  assign n16470 = ~n16468 & ~n16469;
  assign n16471 = n16431 & ~n16470;
  assign n16472 = ~n16431 & n16470;
  assign n16473 = ~n16471 & ~n16472;
  assign n16474 = ~n16421 & n16473;
  assign n16475 = ~n16421 & ~n16474;
  assign n16476 = n16473 & ~n16474;
  assign n16477 = ~n16475 & ~n16476;
  assign n16478 = ~n16380 & ~n16382;
  assign n16479 = ~n16393 & ~n16397;
  assign n16480 = n16478 & n16479;
  assign n16481 = ~n16478 & ~n16479;
  assign n16482 = ~n16480 & ~n16481;
  assign n16483 = ~n16355 & ~n16359;
  assign n16484 = n5235 & n9123;
  assign n16485 = pi41  & pi63 ;
  assign n16486 = ~n13360 & ~n16485;
  assign n16487 = ~n16484 & ~n16486;
  assign n16488 = ~n16346 & n16487;
  assign n16489 = n16346 & ~n16487;
  assign n16490 = ~n16488 & ~n16489;
  assign n16491 = n16483 & ~n16490;
  assign n16492 = ~n16483 & n16490;
  assign n16493 = ~n16491 & ~n16492;
  assign n16494 = ~n16362 & ~n16375;
  assign n16495 = ~n16493 & n16494;
  assign n16496 = n16493 & ~n16494;
  assign n16497 = ~n16495 & ~n16496;
  assign n16498 = n16482 & n16497;
  assign n16499 = ~n16482 & ~n16497;
  assign n16500 = ~n16498 & ~n16499;
  assign n16501 = ~n16477 & n16500;
  assign n16502 = ~n16477 & ~n16501;
  assign n16503 = n16500 & ~n16501;
  assign n16504 = ~n16502 & ~n16503;
  assign n16505 = ~n16420 & ~n16504;
  assign n16506 = n16420 & n16504;
  assign n16507 = ~n16505 & ~n16506;
  assign n16508 = ~n16419 & n16507;
  assign n16509 = n16419 & ~n16507;
  assign po105  = ~n16508 & ~n16509;
  assign n16511 = n16450 & n16464;
  assign n16512 = ~n16450 & ~n16464;
  assign n16513 = ~n16511 & ~n16512;
  assign n16514 = n16439 & ~n16513;
  assign n16515 = ~n16439 & n16513;
  assign n16516 = ~n16514 & ~n16515;
  assign n16517 = ~n16453 & ~n16467;
  assign n16518 = ~n16516 & n16517;
  assign n16519 = n16516 & ~n16517;
  assign n16520 = ~n16518 & ~n16519;
  assign n16521 = ~n16492 & ~n16496;
  assign n16522 = ~n16520 & n16521;
  assign n16523 = n16520 & ~n16521;
  assign n16524 = ~n16522 & ~n16523;
  assign n16525 = ~n16481 & ~n16498;
  assign n16526 = n16524 & ~n16525;
  assign n16527 = ~n16524 & n16525;
  assign n16528 = ~n16526 & ~n16527;
  assign n16529 = ~n16430 & ~n16471;
  assign n16530 = pi62  & n15571;
  assign n16531 = n9144 & ~n16530;
  assign n16532 = ~n16530 & ~n16531;
  assign n16533 = ~pi53  & ~n13777;
  assign n16534 = n16532 & ~n16533;
  assign n16535 = n9144 & ~n16531;
  assign n16536 = ~n16534 & ~n16535;
  assign n16537 = pi49  & pi56 ;
  assign n16538 = n6114 & n9891;
  assign n16539 = pi51  & pi54 ;
  assign n16540 = pi50  & pi55 ;
  assign n16541 = ~n16539 & ~n16540;
  assign n16542 = n16537 & ~n16538;
  assign n16543 = ~n16541 & n16542;
  assign n16544 = n16537 & ~n16543;
  assign n16545 = ~n16538 & ~n16543;
  assign n16546 = ~n16541 & n16545;
  assign n16547 = ~n16544 & ~n16546;
  assign n16548 = ~n16536 & ~n16547;
  assign n16549 = ~n16536 & ~n16548;
  assign n16550 = ~n16547 & ~n16548;
  assign n16551 = ~n16549 & ~n16550;
  assign n16552 = ~n16423 & ~n16426;
  assign n16553 = n16551 & n16552;
  assign n16554 = ~n16551 & ~n16552;
  assign n16555 = ~n16553 & ~n16554;
  assign n16556 = pi42  & pi63 ;
  assign n16557 = n5318 & n9054;
  assign n16558 = pi44  & pi61 ;
  assign n16559 = pi45  & pi60 ;
  assign n16560 = ~n16558 & ~n16559;
  assign n16561 = n16556 & ~n16557;
  assign n16562 = ~n16560 & n16561;
  assign n16563 = n16556 & ~n16562;
  assign n16564 = ~n16557 & ~n16562;
  assign n16565 = ~n16560 & n16564;
  assign n16566 = ~n16563 & ~n16565;
  assign n16567 = ~n16484 & ~n16488;
  assign n16568 = ~n16566 & n16567;
  assign n16569 = n16566 & ~n16567;
  assign n16570 = ~n16568 & ~n16569;
  assign n16571 = pi46  & pi59 ;
  assign n16572 = n5823 & n8144;
  assign n16573 = pi47  & pi58 ;
  assign n16574 = pi48  & pi57 ;
  assign n16575 = ~n16573 & ~n16574;
  assign n16576 = n16571 & ~n16572;
  assign n16577 = ~n16575 & n16576;
  assign n16578 = n16571 & ~n16577;
  assign n16579 = ~n16572 & ~n16577;
  assign n16580 = ~n16575 & n16579;
  assign n16581 = ~n16578 & ~n16580;
  assign n16582 = ~n16570 & ~n16581;
  assign n16583 = n16570 & n16581;
  assign n16584 = ~n16582 & ~n16583;
  assign n16585 = ~n16555 & ~n16584;
  assign n16586 = n16555 & n16584;
  assign n16587 = ~n16585 & ~n16586;
  assign n16588 = ~n16529 & n16587;
  assign n16589 = n16529 & ~n16587;
  assign n16590 = ~n16588 & ~n16589;
  assign n16591 = n16528 & n16590;
  assign n16592 = ~n16528 & ~n16590;
  assign n16593 = ~n16591 & ~n16592;
  assign n16594 = ~n16474 & ~n16501;
  assign n16595 = ~n16593 & n16594;
  assign n16596 = n16593 & ~n16594;
  assign n16597 = ~n16595 & ~n16596;
  assign n16598 = ~n16505 & ~n16508;
  assign n16599 = ~n16597 & n16598;
  assign n16600 = n16597 & ~n16598;
  assign po106  = ~n16599 & ~n16600;
  assign n16602 = ~n16526 & ~n16591;
  assign n16603 = ~n16519 & ~n16523;
  assign n16604 = pi48  & pi58 ;
  assign n16605 = ~n11798 & ~n16604;
  assign n16606 = n8144 & n8505;
  assign n16607 = pi47  & pi59 ;
  assign n16608 = ~n16605 & n16607;
  assign n16609 = ~n16606 & n16608;
  assign n16610 = ~n16606 & ~n16609;
  assign n16611 = ~n16605 & n16610;
  assign n16612 = n16607 & ~n16609;
  assign n16613 = ~n16611 & ~n16612;
  assign n16614 = pi50  & pi56 ;
  assign n16615 = n9891 & n10319;
  assign n16616 = pi51  & pi55 ;
  assign n16617 = ~n11093 & ~n16616;
  assign n16618 = n16614 & ~n16615;
  assign n16619 = ~n16617 & n16618;
  assign n16620 = n16614 & ~n16619;
  assign n16621 = ~n16615 & ~n16619;
  assign n16622 = ~n16617 & n16621;
  assign n16623 = ~n16620 & ~n16622;
  assign n16624 = ~n16613 & ~n16623;
  assign n16625 = ~n16613 & ~n16624;
  assign n16626 = ~n16623 & ~n16624;
  assign n16627 = ~n16625 & ~n16626;
  assign n16628 = ~n16512 & ~n16515;
  assign n16629 = n16627 & n16628;
  assign n16630 = ~n16627 & ~n16628;
  assign n16631 = ~n16629 & ~n16630;
  assign n16632 = n16564 & n16579;
  assign n16633 = ~n16564 & ~n16579;
  assign n16634 = ~n16632 & ~n16633;
  assign n16635 = n7513 & n9054;
  assign n16636 = pi45  & pi61 ;
  assign n16637 = pi46  & pi60 ;
  assign n16638 = ~n16636 & ~n16637;
  assign n16639 = n14117 & ~n16635;
  assign n16640 = ~n16638 & n16639;
  assign n16641 = n14117 & ~n16640;
  assign n16642 = ~n16635 & ~n16640;
  assign n16643 = ~n16638 & n16642;
  assign n16644 = ~n16641 & ~n16643;
  assign n16645 = n16634 & ~n16644;
  assign n16646 = n16634 & ~n16645;
  assign n16647 = ~n16644 & ~n16645;
  assign n16648 = ~n16646 & ~n16647;
  assign n16649 = n16631 & ~n16648;
  assign n16650 = ~n16631 & n16648;
  assign n16651 = ~n16649 & ~n16650;
  assign n16652 = ~n16603 & n16651;
  assign n16653 = ~n16603 & ~n16652;
  assign n16654 = ~n16649 & ~n16652;
  assign n16655 = ~n16650 & n16654;
  assign n16656 = ~n16653 & ~n16655;
  assign n16657 = pi43  & pi63 ;
  assign n16658 = ~n16532 & n16657;
  assign n16659 = n16532 & ~n16657;
  assign n16660 = ~n16658 & ~n16659;
  assign n16661 = n16545 & ~n16660;
  assign n16662 = ~n16545 & n16660;
  assign n16663 = ~n16661 & ~n16662;
  assign n16664 = ~n16566 & ~n16567;
  assign n16665 = ~n16582 & ~n16664;
  assign n16666 = ~n16663 & n16665;
  assign n16667 = n16663 & ~n16665;
  assign n16668 = ~n16666 & ~n16667;
  assign n16669 = ~n16548 & ~n16554;
  assign n16670 = ~n16668 & n16669;
  assign n16671 = n16668 & ~n16669;
  assign n16672 = ~n16670 & ~n16671;
  assign n16673 = ~n16586 & ~n16588;
  assign n16674 = n16672 & ~n16673;
  assign n16675 = ~n16672 & n16673;
  assign n16676 = ~n16674 & ~n16675;
  assign n16677 = n16656 & n16676;
  assign n16678 = ~n16656 & ~n16676;
  assign n16679 = ~n16677 & ~n16678;
  assign n16680 = ~n16602 & ~n16679;
  assign n16681 = n16602 & n16679;
  assign n16682 = ~n16680 & ~n16681;
  assign n16683 = ~n16596 & ~n16600;
  assign n16684 = ~n16682 & n16683;
  assign n16685 = ~n16681 & ~n16683;
  assign n16686 = ~n16680 & n16685;
  assign po107  = ~n16684 & ~n16686;
  assign n16688 = ~n16680 & ~n16685;
  assign n16689 = ~n16667 & ~n16671;
  assign n16690 = n16610 & n16642;
  assign n16691 = ~n16610 & ~n16642;
  assign n16692 = ~n16690 & ~n16691;
  assign n16693 = pi48  & pi59 ;
  assign n16694 = pi58  & pi63 ;
  assign n16695 = n7690 & n16694;
  assign n16696 = pi44  & pi63 ;
  assign n16697 = pi49  & pi58 ;
  assign n16698 = ~n16696 & ~n16697;
  assign n16699 = n16693 & ~n16695;
  assign n16700 = ~n16698 & n16699;
  assign n16701 = n16693 & ~n16700;
  assign n16702 = ~n16695 & ~n16700;
  assign n16703 = ~n16698 & n16702;
  assign n16704 = ~n16701 & ~n16703;
  assign n16705 = n16692 & ~n16704;
  assign n16706 = n16692 & ~n16705;
  assign n16707 = ~n16704 & ~n16705;
  assign n16708 = ~n16706 & ~n16707;
  assign n16709 = pi54  & n14478;
  assign n16710 = n8092 & ~n16709;
  assign n16711 = ~n16709 & ~n16710;
  assign n16712 = ~pi54  & ~n14478;
  assign n16713 = n16711 & ~n16712;
  assign n16714 = n8092 & ~n16710;
  assign n16715 = ~n16713 & ~n16714;
  assign n16716 = pi50  & pi57 ;
  assign n16717 = n8521 & n10319;
  assign n16718 = pi52  & pi55 ;
  assign n16719 = pi51  & pi56 ;
  assign n16720 = ~n16718 & ~n16719;
  assign n16721 = n16716 & ~n16717;
  assign n16722 = ~n16720 & n16721;
  assign n16723 = n16716 & ~n16722;
  assign n16724 = ~n16717 & ~n16722;
  assign n16725 = ~n16720 & n16724;
  assign n16726 = ~n16723 & ~n16725;
  assign n16727 = ~n16715 & ~n16726;
  assign n16728 = ~n16715 & ~n16727;
  assign n16729 = ~n16726 & ~n16727;
  assign n16730 = ~n16728 & ~n16729;
  assign n16731 = n5277 & n9054;
  assign n16732 = pi47  & pi60 ;
  assign n16733 = ~n16731 & n16732;
  assign n16734 = pi46  & pi61 ;
  assign n16735 = ~n16731 & n16734;
  assign n16736 = ~n16733 & ~n16735;
  assign n16737 = ~n16621 & ~n16736;
  assign n16738 = ~n16621 & ~n16737;
  assign n16739 = ~n16736 & ~n16737;
  assign n16740 = ~n16738 & ~n16739;
  assign n16741 = ~n16730 & n16740;
  assign n16742 = n16730 & ~n16740;
  assign n16743 = ~n16741 & ~n16742;
  assign n16744 = ~n16708 & ~n16743;
  assign n16745 = n16708 & n16743;
  assign n16746 = ~n16744 & ~n16745;
  assign n16747 = n16689 & ~n16746;
  assign n16748 = ~n16689 & n16746;
  assign n16749 = ~n16747 & ~n16748;
  assign n16750 = ~n16633 & ~n16645;
  assign n16751 = ~n16658 & ~n16662;
  assign n16752 = n16750 & n16751;
  assign n16753 = ~n16750 & ~n16751;
  assign n16754 = ~n16752 & ~n16753;
  assign n16755 = ~n16624 & ~n16630;
  assign n16756 = ~n16754 & n16755;
  assign n16757 = n16754 & ~n16755;
  assign n16758 = ~n16756 & ~n16757;
  assign n16759 = ~n16654 & n16758;
  assign n16760 = n16654 & ~n16758;
  assign n16761 = ~n16759 & ~n16760;
  assign n16762 = n16749 & n16761;
  assign n16763 = ~n16749 & ~n16761;
  assign n16764 = ~n16762 & ~n16763;
  assign n16765 = ~n16675 & ~n16677;
  assign n16766 = ~n16764 & ~n16765;
  assign n16767 = n16764 & n16765;
  assign n16768 = ~n16766 & ~n16767;
  assign n16769 = ~n16688 & ~n16768;
  assign n16770 = n16688 & n16768;
  assign po108  = n16769 | n16770;
  assign n16772 = ~n16688 & ~n16766;
  assign n16773 = ~n16767 & ~n16772;
  assign n16774 = ~n16759 & ~n16762;
  assign n16775 = ~n16691 & ~n16705;
  assign n16776 = n8521 & n9144;
  assign n16777 = pi52  & pi56 ;
  assign n16778 = ~n7172 & ~n16777;
  assign n16779 = n13406 & ~n16776;
  assign n16780 = ~n16778 & n16779;
  assign n16781 = n13406 & ~n16780;
  assign n16782 = ~n16776 & ~n16780;
  assign n16783 = ~n16778 & n16782;
  assign n16784 = ~n16781 & ~n16783;
  assign n16785 = ~n16775 & ~n16784;
  assign n16786 = ~n16775 & ~n16785;
  assign n16787 = ~n16784 & ~n16785;
  assign n16788 = ~n16786 & ~n16787;
  assign n16789 = ~n16730 & ~n16740;
  assign n16790 = ~n16727 & ~n16789;
  assign n16791 = ~n16788 & ~n16790;
  assign n16792 = ~n16788 & ~n16791;
  assign n16793 = ~n16790 & ~n16791;
  assign n16794 = ~n16792 & ~n16793;
  assign n16795 = ~n16744 & ~n16748;
  assign n16796 = n16794 & n16795;
  assign n16797 = ~n16794 & ~n16795;
  assign n16798 = ~n16796 & ~n16797;
  assign n16799 = n16711 & n16724;
  assign n16800 = ~n16711 & ~n16724;
  assign n16801 = ~n16799 & ~n16800;
  assign n16802 = n16702 & ~n16801;
  assign n16803 = ~n16702 & n16801;
  assign n16804 = ~n16802 & ~n16803;
  assign n16805 = ~n16753 & ~n16757;
  assign n16806 = ~n16804 & n16805;
  assign n16807 = n16804 & ~n16805;
  assign n16808 = ~n16806 & ~n16807;
  assign n16809 = pi45  & pi63 ;
  assign n16810 = n5277 & n9567;
  assign n16811 = pi47  & pi61 ;
  assign n16812 = ~n14794 & ~n16811;
  assign n16813 = n16809 & ~n16810;
  assign n16814 = ~n16812 & n16813;
  assign n16815 = n16809 & ~n16814;
  assign n16816 = ~n16810 & ~n16814;
  assign n16817 = ~n16812 & n16816;
  assign n16818 = ~n16815 & ~n16817;
  assign n16819 = ~n16731 & ~n16737;
  assign n16820 = ~n16818 & n16819;
  assign n16821 = n16818 & ~n16819;
  assign n16822 = ~n16820 & ~n16821;
  assign n16823 = pi48  & pi60 ;
  assign n16824 = n5889 & n9402;
  assign n16825 = pi49  & pi59 ;
  assign n16826 = pi50  & pi58 ;
  assign n16827 = ~n16825 & ~n16826;
  assign n16828 = n16823 & ~n16824;
  assign n16829 = ~n16827 & n16828;
  assign n16830 = n16823 & ~n16829;
  assign n16831 = ~n16824 & ~n16829;
  assign n16832 = ~n16827 & n16831;
  assign n16833 = ~n16830 & ~n16832;
  assign n16834 = ~n16822 & ~n16833;
  assign n16835 = n16822 & n16833;
  assign n16836 = ~n16834 & ~n16835;
  assign n16837 = n16808 & n16836;
  assign n16838 = ~n16808 & ~n16836;
  assign n16839 = ~n16837 & ~n16838;
  assign n16840 = n16798 & n16839;
  assign n16841 = n16798 & ~n16840;
  assign n16842 = n16839 & ~n16840;
  assign n16843 = ~n16841 & ~n16842;
  assign n16844 = n16774 & n16843;
  assign n16845 = ~n16774 & ~n16843;
  assign n16846 = ~n16844 & ~n16845;
  assign n16847 = n16773 & ~n16846;
  assign n16848 = ~n16773 & ~n16844;
  assign n16849 = ~n16845 & n16848;
  assign po109  = ~n16847 & ~n16849;
  assign n16851 = ~n16845 & ~n16848;
  assign n16852 = ~n16800 & ~n16803;
  assign n16853 = pi55  & n15174;
  assign n16854 = n9891 & ~n16853;
  assign n16855 = n9891 & ~n16854;
  assign n16856 = ~n16853 & ~n16854;
  assign n16857 = ~pi55  & ~n15174;
  assign n16858 = n16856 & ~n16857;
  assign n16859 = ~n16855 & ~n16858;
  assign n16860 = ~n16852 & ~n16859;
  assign n16861 = ~n16852 & ~n16860;
  assign n16862 = ~n16859 & ~n16860;
  assign n16863 = ~n16861 & ~n16862;
  assign n16864 = ~n16818 & ~n16819;
  assign n16865 = ~n16834 & ~n16864;
  assign n16866 = n16863 & n16865;
  assign n16867 = ~n16863 & ~n16865;
  assign n16868 = ~n16866 & ~n16867;
  assign n16869 = ~n16807 & ~n16837;
  assign n16870 = n16868 & ~n16869;
  assign n16871 = ~n16868 & n16869;
  assign n16872 = ~n16870 & ~n16871;
  assign n16873 = pi46  & pi63 ;
  assign n16874 = ~n16782 & n16873;
  assign n16875 = n16782 & ~n16873;
  assign n16876 = ~n16874 & ~n16875;
  assign n16877 = n16831 & ~n16876;
  assign n16878 = ~n16831 & n16876;
  assign n16879 = ~n16877 & ~n16878;
  assign n16880 = ~n16785 & ~n16791;
  assign n16881 = ~n16879 & n16880;
  assign n16882 = n16879 & ~n16880;
  assign n16883 = ~n16881 & ~n16882;
  assign n16884 = pi48  & pi61 ;
  assign n16885 = n5889 & n8854;
  assign n16886 = pi49  & pi60 ;
  assign n16887 = pi50  & pi59 ;
  assign n16888 = ~n16886 & ~n16887;
  assign n16889 = n16884 & ~n16885;
  assign n16890 = ~n16888 & n16889;
  assign n16891 = n16884 & ~n16890;
  assign n16892 = ~n16885 & ~n16890;
  assign n16893 = ~n16888 & n16892;
  assign n16894 = ~n16891 & ~n16893;
  assign n16895 = n16816 & ~n16894;
  assign n16896 = ~n16816 & n16894;
  assign n16897 = ~n16895 & ~n16896;
  assign n16898 = pi51  & pi58 ;
  assign n16899 = n7643 & n9144;
  assign n16900 = pi53  & pi56 ;
  assign n16901 = pi52  & pi57 ;
  assign n16902 = ~n16900 & ~n16901;
  assign n16903 = n16898 & ~n16899;
  assign n16904 = ~n16902 & n16903;
  assign n16905 = n16898 & ~n16904;
  assign n16906 = ~n16899 & ~n16904;
  assign n16907 = ~n16902 & n16906;
  assign n16908 = ~n16905 & ~n16907;
  assign n16909 = ~n16897 & ~n16908;
  assign n16910 = n16897 & n16908;
  assign n16911 = ~n16909 & ~n16910;
  assign n16912 = n16883 & n16911;
  assign n16913 = ~n16883 & ~n16911;
  assign n16914 = ~n16912 & ~n16913;
  assign n16915 = n16872 & n16914;
  assign n16916 = n16872 & ~n16915;
  assign n16917 = n16914 & ~n16915;
  assign n16918 = ~n16916 & ~n16917;
  assign n16919 = ~n16797 & ~n16840;
  assign n16920 = ~n16918 & ~n16919;
  assign n16921 = n16918 & n16919;
  assign n16922 = ~n16920 & ~n16921;
  assign n16923 = ~n16851 & ~n16922;
  assign n16924 = n16851 & n16922;
  assign po110  = n16923 | n16924;
  assign n16926 = ~n16851 & ~n16921;
  assign n16927 = ~n16920 & ~n16926;
  assign n16928 = ~n16870 & ~n16915;
  assign n16929 = n16892 & n16906;
  assign n16930 = ~n16892 & ~n16906;
  assign n16931 = ~n16929 & ~n16930;
  assign n16932 = pi49  & pi61 ;
  assign n16933 = n6114 & n8854;
  assign n16934 = pi50  & pi60 ;
  assign n16935 = pi51  & pi59 ;
  assign n16936 = ~n16934 & ~n16935;
  assign n16937 = n16932 & ~n16933;
  assign n16938 = ~n16936 & n16937;
  assign n16939 = n16932 & ~n16938;
  assign n16940 = ~n16933 & ~n16938;
  assign n16941 = ~n16936 & n16940;
  assign n16942 = ~n16939 & ~n16941;
  assign n16943 = n16931 & ~n16942;
  assign n16944 = n16931 & ~n16943;
  assign n16945 = ~n16942 & ~n16943;
  assign n16946 = ~n16944 & ~n16945;
  assign n16947 = ~n16816 & ~n16894;
  assign n16948 = ~n16909 & ~n16947;
  assign n16949 = n16946 & n16948;
  assign n16950 = ~n16946 & ~n16948;
  assign n16951 = ~n16949 & ~n16950;
  assign n16952 = ~n16860 & ~n16867;
  assign n16953 = ~n16951 & n16952;
  assign n16954 = n16951 & ~n16952;
  assign n16955 = ~n16953 & ~n16954;
  assign n16956 = n5823 & n9123;
  assign n16957 = pi47  & pi63 ;
  assign n16958 = ~n15374 & ~n16957;
  assign n16959 = ~n16956 & ~n16958;
  assign n16960 = ~n16856 & n16959;
  assign n16961 = n16856 & ~n16959;
  assign n16962 = ~n16960 & ~n16961;
  assign n16963 = pi52  & pi58 ;
  assign n16964 = n7643 & n8092;
  assign n16965 = pi53  & pi57 ;
  assign n16966 = ~n6911 & ~n16965;
  assign n16967 = n16963 & ~n16964;
  assign n16968 = ~n16966 & n16967;
  assign n16969 = n16963 & ~n16968;
  assign n16970 = ~n16964 & ~n16968;
  assign n16971 = ~n16966 & n16970;
  assign n16972 = ~n16969 & ~n16971;
  assign n16973 = n16962 & ~n16972;
  assign n16974 = n16962 & ~n16973;
  assign n16975 = ~n16972 & ~n16973;
  assign n16976 = ~n16974 & ~n16975;
  assign n16977 = ~n16874 & ~n16878;
  assign n16978 = n16976 & n16977;
  assign n16979 = ~n16976 & ~n16977;
  assign n16980 = ~n16978 & ~n16979;
  assign n16981 = ~n16882 & ~n16912;
  assign n16982 = n16980 & ~n16981;
  assign n16983 = n16980 & ~n16982;
  assign n16984 = ~n16981 & ~n16982;
  assign n16985 = ~n16983 & ~n16984;
  assign n16986 = n16955 & ~n16985;
  assign n16987 = ~n16955 & n16985;
  assign n16988 = ~n16986 & ~n16987;
  assign n16989 = n16928 & ~n16988;
  assign n16990 = ~n16928 & n16988;
  assign n16991 = ~n16989 & ~n16990;
  assign n16992 = n16927 & ~n16991;
  assign n16993 = ~n16927 & ~n16989;
  assign n16994 = ~n16990 & n16993;
  assign po111  = ~n16992 & ~n16994;
  assign n16996 = ~n16990 & ~n16993;
  assign n16997 = ~n16982 & ~n16986;
  assign n16998 = n16940 & n16970;
  assign n16999 = ~n16940 & ~n16970;
  assign n17000 = ~n16998 & ~n16999;
  assign n17001 = ~n16956 & ~n16960;
  assign n17002 = ~n17000 & n17001;
  assign n17003 = n17000 & ~n17001;
  assign n17004 = ~n17002 & ~n17003;
  assign n17005 = ~n16930 & ~n16943;
  assign n17006 = ~n17004 & n17005;
  assign n17007 = n17004 & ~n17005;
  assign n17008 = ~n17006 & ~n17007;
  assign n17009 = ~n16973 & ~n16979;
  assign n17010 = ~n17008 & n17009;
  assign n17011 = n17008 & ~n17009;
  assign n17012 = ~n17010 & ~n17011;
  assign n17013 = pi50  & pi61 ;
  assign n17014 = pi51  & pi60 ;
  assign n17015 = ~n17013 & ~n17014;
  assign n17016 = n6114 & n9054;
  assign n17017 = pi48  & pi63 ;
  assign n17018 = ~n17015 & n17017;
  assign n17019 = ~n17016 & n17018;
  assign n17020 = ~n17016 & ~n17019;
  assign n17021 = ~n17015 & n17020;
  assign n17022 = n17017 & ~n17019;
  assign n17023 = ~n17021 & ~n17022;
  assign n17024 = pi56  & pi62 ;
  assign n17025 = pi49  & n17024;
  assign n17026 = n8521 & ~n17025;
  assign n17027 = n8521 & ~n17026;
  assign n17028 = ~n17025 & ~n17026;
  assign n17029 = ~pi56  & ~n15634;
  assign n17030 = n17028 & ~n17029;
  assign n17031 = ~n17027 & ~n17030;
  assign n17032 = ~n17023 & ~n17031;
  assign n17033 = ~n17023 & ~n17032;
  assign n17034 = ~n17031 & ~n17032;
  assign n17035 = ~n17033 & ~n17034;
  assign n17036 = pi52  & pi59 ;
  assign n17037 = n8092 & n8144;
  assign n17038 = pi53  & pi58 ;
  assign n17039 = ~n15118 & ~n17038;
  assign n17040 = n17036 & ~n17037;
  assign n17041 = ~n17039 & n17040;
  assign n17042 = n17036 & ~n17041;
  assign n17043 = ~n17037 & ~n17041;
  assign n17044 = ~n17039 & n17043;
  assign n17045 = ~n17042 & ~n17044;
  assign n17046 = ~n17035 & ~n17045;
  assign n17047 = ~n17035 & ~n17046;
  assign n17048 = ~n17045 & ~n17046;
  assign n17049 = ~n17047 & ~n17048;
  assign n17050 = ~n16950 & ~n16954;
  assign n17051 = n17049 & n17050;
  assign n17052 = ~n17049 & ~n17050;
  assign n17053 = ~n17051 & ~n17052;
  assign n17054 = n17012 & n17053;
  assign n17055 = ~n17012 & ~n17053;
  assign n17056 = ~n17054 & ~n17055;
  assign n17057 = ~n16997 & n17056;
  assign n17058 = n16997 & ~n17056;
  assign n17059 = ~n17057 & ~n17058;
  assign n17060 = ~n16996 & ~n17059;
  assign n17061 = n16996 & n17059;
  assign po112  = n17060 | n17061;
  assign n17063 = ~n16996 & ~n17058;
  assign n17064 = ~n17057 & ~n17063;
  assign n17065 = ~n17052 & ~n17054;
  assign n17066 = ~n17007 & ~n17011;
  assign n17067 = pi49  & pi63 ;
  assign n17068 = n9054 & n10319;
  assign n17069 = pi51  & pi61 ;
  assign n17070 = pi52  & pi60 ;
  assign n17071 = ~n17069 & ~n17070;
  assign n17072 = n17067 & ~n17068;
  assign n17073 = ~n17071 & n17072;
  assign n17074 = n17067 & ~n17073;
  assign n17075 = ~n17068 & ~n17073;
  assign n17076 = ~n17071 & n17075;
  assign n17077 = ~n17074 & ~n17076;
  assign n17078 = n17020 & ~n17077;
  assign n17079 = ~n17020 & n17077;
  assign n17080 = ~n17078 & ~n17079;
  assign n17081 = pi53  & pi59 ;
  assign n17082 = n8144 & n9891;
  assign n17083 = pi54  & pi58 ;
  assign n17084 = ~n13270 & ~n17083;
  assign n17085 = n17081 & ~n17082;
  assign n17086 = ~n17084 & n17085;
  assign n17087 = n17081 & ~n17086;
  assign n17088 = ~n17082 & ~n17086;
  assign n17089 = ~n17084 & n17088;
  assign n17090 = ~n17087 & ~n17089;
  assign n17091 = ~n17080 & ~n17090;
  assign n17092 = n17080 & n17090;
  assign n17093 = ~n17091 & ~n17092;
  assign n17094 = n17066 & ~n17093;
  assign n17095 = ~n17066 & n17093;
  assign n17096 = ~n17094 & ~n17095;
  assign n17097 = n15865 & ~n17028;
  assign n17098 = ~n15865 & n17028;
  assign n17099 = ~n17097 & ~n17098;
  assign n17100 = n17043 & ~n17099;
  assign n17101 = ~n17043 & n17099;
  assign n17102 = ~n17100 & ~n17101;
  assign n17103 = ~n16999 & ~n17003;
  assign n17104 = ~n17032 & ~n17046;
  assign n17105 = n17103 & n17104;
  assign n17106 = ~n17103 & ~n17104;
  assign n17107 = ~n17105 & ~n17106;
  assign n17108 = n17102 & n17107;
  assign n17109 = ~n17102 & ~n17107;
  assign n17110 = ~n17108 & ~n17109;
  assign n17111 = n17096 & n17110;
  assign n17112 = ~n17096 & ~n17110;
  assign n17113 = ~n17111 & ~n17112;
  assign n17114 = n17065 & ~n17113;
  assign n17115 = ~n17065 & n17113;
  assign n17116 = ~n17114 & ~n17115;
  assign n17117 = n17064 & ~n17116;
  assign n17118 = ~n17064 & ~n17114;
  assign n17119 = ~n17115 & n17118;
  assign po113  = ~n17117 & ~n17119;
  assign n17121 = ~n17115 & ~n17118;
  assign n17122 = ~n17095 & ~n17111;
  assign n17123 = n9054 & n9144;
  assign n17124 = pi53  & pi60 ;
  assign n17125 = ~n17123 & n17124;
  assign n17126 = pi52  & pi61 ;
  assign n17127 = ~n17123 & n17126;
  assign n17128 = ~n17125 & ~n17127;
  assign n17129 = ~n17088 & ~n17128;
  assign n17130 = ~n17088 & ~n17129;
  assign n17131 = ~n17128 & ~n17129;
  assign n17132 = ~n17130 & ~n17131;
  assign n17133 = ~n17097 & ~n17101;
  assign n17134 = n17132 & n17133;
  assign n17135 = ~n17132 & ~n17133;
  assign n17136 = ~n17134 & ~n17135;
  assign n17137 = ~n17020 & ~n17077;
  assign n17138 = ~n17091 & ~n17137;
  assign n17139 = ~n17136 & n17138;
  assign n17140 = n17136 & ~n17138;
  assign n17141 = ~n17139 & ~n17140;
  assign n17142 = ~n17106 & ~n17108;
  assign n17143 = pi50  & pi63 ;
  assign n17144 = n9402 & n9891;
  assign n17145 = pi55  & pi58 ;
  assign n17146 = pi54  & pi59 ;
  assign n17147 = ~n17145 & ~n17146;
  assign n17148 = n17143 & ~n17144;
  assign n17149 = ~n17147 & n17148;
  assign n17150 = n17143 & ~n17149;
  assign n17151 = ~n17144 & ~n17149;
  assign n17152 = ~n17147 & n17151;
  assign n17153 = ~n17150 & ~n17152;
  assign n17154 = n17075 & ~n17153;
  assign n17155 = ~n17075 & n17153;
  assign n17156 = ~n17154 & ~n17155;
  assign n17157 = pi62  & n13406;
  assign n17158 = n7643 & ~n17157;
  assign n17159 = n7643 & ~n17158;
  assign n17160 = ~n17157 & ~n17158;
  assign n17161 = pi51  & pi62 ;
  assign n17162 = ~pi57  & ~n17161;
  assign n17163 = n17160 & ~n17162;
  assign n17164 = ~n17159 & ~n17163;
  assign n17165 = ~n17156 & ~n17164;
  assign n17166 = n17156 & n17164;
  assign n17167 = ~n17165 & ~n17166;
  assign n17168 = ~n17142 & n17167;
  assign n17169 = n17142 & ~n17167;
  assign n17170 = ~n17168 & ~n17169;
  assign n17171 = ~n17141 & ~n17170;
  assign n17172 = n17141 & n17170;
  assign n17173 = ~n17171 & ~n17172;
  assign n17174 = n17122 & ~n17173;
  assign n17175 = ~n17122 & n17173;
  assign n17176 = ~n17174 & ~n17175;
  assign n17177 = ~n17121 & ~n17176;
  assign n17178 = n17121 & n17176;
  assign po114  = n17177 | n17178;
  assign n17180 = ~n17121 & ~n17174;
  assign n17181 = ~n17175 & ~n17180;
  assign n17182 = ~n17168 & ~n17172;
  assign n17183 = n17151 & n17160;
  assign n17184 = ~n17151 & ~n17160;
  assign n17185 = ~n17183 & ~n17184;
  assign n17186 = ~n17123 & ~n17129;
  assign n17187 = ~n17185 & n17186;
  assign n17188 = n17185 & ~n17186;
  assign n17189 = ~n17187 & ~n17188;
  assign n17190 = ~n17135 & ~n17140;
  assign n17191 = ~n17189 & n17190;
  assign n17192 = n17189 & ~n17190;
  assign n17193 = ~n17191 & ~n17192;
  assign n17194 = pi52  & pi62 ;
  assign n17195 = pi53  & pi61 ;
  assign n17196 = ~n17194 & ~n17195;
  assign n17197 = n9144 & n9567;
  assign n17198 = pi51  & pi63 ;
  assign n17199 = ~n17196 & n17198;
  assign n17200 = ~n17197 & n17199;
  assign n17201 = ~n17197 & ~n17200;
  assign n17202 = ~n17196 & n17201;
  assign n17203 = n17198 & ~n17200;
  assign n17204 = ~n17202 & ~n17203;
  assign n17205 = pi54  & pi60 ;
  assign n17206 = n8521 & n9402;
  assign n17207 = pi55  & pi59 ;
  assign n17208 = ~n12970 & ~n17207;
  assign n17209 = n17205 & ~n17206;
  assign n17210 = ~n17208 & n17209;
  assign n17211 = n17205 & ~n17210;
  assign n17212 = ~n17206 & ~n17210;
  assign n17213 = ~n17208 & n17212;
  assign n17214 = ~n17211 & ~n17213;
  assign n17215 = ~n17204 & ~n17214;
  assign n17216 = ~n17204 & ~n17215;
  assign n17217 = ~n17214 & ~n17215;
  assign n17218 = ~n17216 & ~n17217;
  assign n17219 = ~n17075 & ~n17153;
  assign n17220 = ~n17165 & ~n17219;
  assign n17221 = n17218 & n17220;
  assign n17222 = ~n17218 & ~n17220;
  assign n17223 = ~n17221 & ~n17222;
  assign n17224 = n17193 & n17223;
  assign n17225 = ~n17193 & ~n17223;
  assign n17226 = ~n17224 & ~n17225;
  assign n17227 = n17182 & ~n17226;
  assign n17228 = ~n17182 & n17226;
  assign n17229 = ~n17227 & ~n17228;
  assign n17230 = n17181 & ~n17229;
  assign n17231 = ~n17181 & ~n17227;
  assign n17232 = ~n17228 & n17231;
  assign po115  = ~n17230 & ~n17232;
  assign n17234 = ~n17228 & ~n17231;
  assign n17235 = ~n17192 & ~n17224;
  assign n17236 = pi53  & pi62 ;
  assign n17237 = pi58  & n17236;
  assign n17238 = n8144 & ~n17237;
  assign n17239 = ~n17237 & ~n17238;
  assign n17240 = ~pi58  & ~n17236;
  assign n17241 = n17239 & ~n17240;
  assign n17242 = n8144 & ~n17238;
  assign n17243 = ~n17241 & ~n17242;
  assign n17244 = pi54  & pi61 ;
  assign n17245 = n8521 & n8854;
  assign n17246 = pi55  & pi60 ;
  assign n17247 = ~n15489 & ~n17246;
  assign n17248 = n17244 & ~n17245;
  assign n17249 = ~n17247 & n17248;
  assign n17250 = n17244 & ~n17249;
  assign n17251 = ~n17245 & ~n17249;
  assign n17252 = ~n17247 & n17251;
  assign n17253 = ~n17250 & ~n17252;
  assign n17254 = ~n17243 & ~n17253;
  assign n17255 = ~n17243 & ~n17254;
  assign n17256 = ~n17253 & ~n17254;
  assign n17257 = ~n17255 & ~n17256;
  assign n17258 = ~n17184 & ~n17188;
  assign n17259 = n17257 & n17258;
  assign n17260 = ~n17257 & ~n17258;
  assign n17261 = ~n17259 & ~n17260;
  assign n17262 = pi52  & pi63 ;
  assign n17263 = ~n17212 & n17262;
  assign n17264 = n17212 & ~n17262;
  assign n17265 = ~n17263 & ~n17264;
  assign n17266 = n17201 & ~n17265;
  assign n17267 = ~n17201 & n17265;
  assign n17268 = ~n17266 & ~n17267;
  assign n17269 = ~n17215 & ~n17222;
  assign n17270 = ~n17268 & n17269;
  assign n17271 = n17268 & ~n17269;
  assign n17272 = ~n17270 & ~n17271;
  assign n17273 = n17261 & n17272;
  assign n17274 = ~n17261 & ~n17272;
  assign n17275 = ~n17273 & ~n17274;
  assign n17276 = ~n17235 & n17275;
  assign n17277 = n17235 & ~n17275;
  assign n17278 = ~n17276 & ~n17277;
  assign n17279 = ~n17234 & ~n17278;
  assign n17280 = n17234 & n17278;
  assign po116  = n17279 | n17280;
  assign n17282 = ~n17234 & ~n17277;
  assign n17283 = ~n17276 & ~n17282;
  assign n17284 = ~n17254 & ~n17260;
  assign n17285 = ~n17263 & ~n17267;
  assign n17286 = n17284 & n17285;
  assign n17287 = ~n17284 & ~n17285;
  assign n17288 = ~n17286 & ~n17287;
  assign n17289 = n8092 & n9123;
  assign n17290 = pi54  & pi62 ;
  assign n17291 = ~n17289 & n17290;
  assign n17292 = pi53  & pi63 ;
  assign n17293 = ~n17289 & n17292;
  assign n17294 = ~n17291 & ~n17293;
  assign n17295 = ~n17239 & ~n17294;
  assign n17296 = ~n17239 & ~n17295;
  assign n17297 = ~n17294 & ~n17295;
  assign n17298 = ~n17296 & ~n17297;
  assign n17299 = pi55  & pi61 ;
  assign n17300 = n7643 & n8854;
  assign n17301 = pi56  & pi60 ;
  assign n17302 = ~n12351 & ~n17301;
  assign n17303 = n17299 & ~n17300;
  assign n17304 = ~n17302 & n17303;
  assign n17305 = n17299 & ~n17304;
  assign n17306 = ~n17300 & ~n17304;
  assign n17307 = ~n17302 & n17306;
  assign n17308 = ~n17305 & ~n17307;
  assign n17309 = ~n17251 & ~n17308;
  assign n17310 = ~n17251 & ~n17309;
  assign n17311 = ~n17308 & ~n17309;
  assign n17312 = ~n17310 & ~n17311;
  assign n17313 = ~n17298 & ~n17312;
  assign n17314 = n17298 & n17312;
  assign n17315 = ~n17313 & ~n17314;
  assign n17316 = n17288 & n17315;
  assign n17317 = ~n17288 & ~n17315;
  assign n17318 = ~n17316 & ~n17317;
  assign n17319 = ~n17271 & ~n17273;
  assign n17320 = ~n17318 & n17319;
  assign n17321 = n17318 & ~n17319;
  assign n17322 = ~n17320 & ~n17321;
  assign n17323 = n17283 & ~n17322;
  assign n17324 = ~n17283 & ~n17320;
  assign n17325 = ~n17321 & n17324;
  assign po117  = ~n17323 & ~n17325;
  assign n17327 = ~n17321 & ~n17324;
  assign n17328 = ~n17287 & ~n17316;
  assign n17329 = ~n17289 & ~n17295;
  assign n17330 = n17306 & n17329;
  assign n17331 = ~n17306 & ~n17329;
  assign n17332 = ~n17330 & ~n17331;
  assign n17333 = pi54  & pi63 ;
  assign n17334 = n7643 & n9054;
  assign n17335 = pi57  & pi60 ;
  assign n17336 = pi56  & pi61 ;
  assign n17337 = ~n17335 & ~n17336;
  assign n17338 = n17333 & ~n17334;
  assign n17339 = ~n17337 & n17338;
  assign n17340 = n17333 & ~n17339;
  assign n17341 = ~n17334 & ~n17339;
  assign n17342 = ~n17337 & n17341;
  assign n17343 = ~n17340 & ~n17342;
  assign n17344 = n17332 & ~n17343;
  assign n17345 = n17332 & ~n17344;
  assign n17346 = ~n17343 & ~n17344;
  assign n17347 = ~n17345 & ~n17346;
  assign n17348 = ~n17309 & ~n17313;
  assign n17349 = pi59  & pi62 ;
  assign n17350 = pi55  & n17349;
  assign n17351 = n9402 & ~n17350;
  assign n17352 = n9402 & ~n17351;
  assign n17353 = ~n17350 & ~n17351;
  assign n17354 = pi55  & pi62 ;
  assign n17355 = ~pi59  & ~n17354;
  assign n17356 = n17353 & ~n17355;
  assign n17357 = ~n17352 & ~n17356;
  assign n17358 = ~n17348 & ~n17357;
  assign n17359 = ~n17348 & ~n17358;
  assign n17360 = ~n17357 & ~n17358;
  assign n17361 = ~n17359 & ~n17360;
  assign n17362 = ~n17347 & n17361;
  assign n17363 = n17347 & ~n17361;
  assign n17364 = ~n17362 & ~n17363;
  assign n17365 = ~n17328 & ~n17364;
  assign n17366 = n17328 & n17364;
  assign n17367 = ~n17365 & ~n17366;
  assign n17368 = ~n17327 & ~n17367;
  assign n17369 = n17327 & n17367;
  assign po118  = n17368 | n17369;
  assign n17371 = pi55  & pi63 ;
  assign n17372 = ~n17353 & n17371;
  assign n17373 = n17353 & ~n17371;
  assign n17374 = ~n17372 & ~n17373;
  assign n17375 = n17341 & ~n17374;
  assign n17376 = ~n17341 & n17374;
  assign n17377 = ~n17375 & ~n17376;
  assign n17378 = ~n17331 & ~n17344;
  assign n17379 = n8144 & n9054;
  assign n17380 = pi58  & pi60 ;
  assign n17381 = pi57  & pi61 ;
  assign n17382 = ~n17380 & ~n17381;
  assign n17383 = n17024 & ~n17379;
  assign n17384 = ~n17382 & n17383;
  assign n17385 = n17024 & ~n17384;
  assign n17386 = ~n17379 & ~n17384;
  assign n17387 = ~n17382 & n17386;
  assign n17388 = ~n17385 & ~n17387;
  assign n17389 = ~n17378 & ~n17388;
  assign n17390 = ~n17378 & ~n17389;
  assign n17391 = ~n17388 & ~n17389;
  assign n17392 = ~n17390 & ~n17391;
  assign n17393 = ~n17377 & n17392;
  assign n17394 = n17377 & ~n17392;
  assign n17395 = ~n17393 & ~n17394;
  assign n17396 = ~n17347 & ~n17361;
  assign n17397 = ~n17358 & ~n17396;
  assign n17398 = ~n17395 & n17397;
  assign n17399 = n17395 & ~n17397;
  assign n17400 = ~n17398 & ~n17399;
  assign n17401 = ~n17327 & ~n17366;
  assign n17402 = ~n17365 & ~n17401;
  assign n17403 = ~n17400 & n17402;
  assign n17404 = n17400 & ~n17402;
  assign po119  = ~n17403 & ~n17404;
  assign n17406 = n9236 & n12970;
  assign n17407 = pi58  & pi61 ;
  assign n17408 = ~n17406 & n17407;
  assign n17409 = pi56  & pi63 ;
  assign n17410 = ~n17406 & n17409;
  assign n17411 = ~n17408 & ~n17410;
  assign n17412 = ~n17386 & ~n17411;
  assign n17413 = ~n17386 & ~n17412;
  assign n17414 = ~n17411 & ~n17412;
  assign n17415 = ~n17413 & ~n17414;
  assign n17416 = pi57  & n8453;
  assign n17417 = n8854 & ~n17416;
  assign n17418 = n8854 & ~n17417;
  assign n17419 = ~n17416 & ~n17417;
  assign n17420 = pi57  & pi62 ;
  assign n17421 = ~pi60  & ~n17420;
  assign n17422 = n17419 & ~n17421;
  assign n17423 = ~n17418 & ~n17422;
  assign n17424 = ~n17415 & ~n17423;
  assign n17425 = ~n17415 & ~n17424;
  assign n17426 = ~n17423 & ~n17424;
  assign n17427 = ~n17425 & ~n17426;
  assign n17428 = ~n17372 & ~n17376;
  assign n17429 = n17427 & n17428;
  assign n17430 = ~n17427 & ~n17428;
  assign n17431 = ~n17429 & ~n17430;
  assign n17432 = ~n17389 & ~n17394;
  assign n17433 = n17431 & ~n17432;
  assign n17434 = ~n17431 & n17432;
  assign n17435 = ~n17433 & ~n17434;
  assign n17436 = ~n17399 & ~n17404;
  assign n17437 = ~n17435 & n17436;
  assign n17438 = n17435 & ~n17436;
  assign po120  = ~n17437 & ~n17438;
  assign n17440 = ~n17424 & ~n17430;
  assign n17441 = ~n17406 & ~n17412;
  assign n17442 = n17419 & n17441;
  assign n17443 = ~n17419 & ~n17441;
  assign n17444 = ~n17442 & ~n17443;
  assign n17445 = pi57  & pi63 ;
  assign n17446 = n9402 & n9567;
  assign n17447 = pi58  & pi62 ;
  assign n17448 = ~n15297 & ~n17447;
  assign n17449 = n17445 & ~n17446;
  assign n17450 = ~n17448 & n17449;
  assign n17451 = n17445 & ~n17450;
  assign n17452 = ~n17446 & ~n17450;
  assign n17453 = ~n17448 & n17452;
  assign n17454 = ~n17451 & ~n17453;
  assign n17455 = n17444 & ~n17454;
  assign n17456 = ~n17444 & n17454;
  assign n17457 = ~n17455 & ~n17456;
  assign n17458 = n17440 & ~n17457;
  assign n17459 = ~n17440 & n17457;
  assign n17460 = ~n17458 & ~n17459;
  assign n17461 = ~n17433 & ~n17438;
  assign n17462 = ~n17460 & n17461;
  assign n17463 = ~n17458 & ~n17461;
  assign n17464 = ~n17459 & n17463;
  assign po121  = ~n17462 & ~n17464;
  assign n17466 = ~pi60  & pi61 ;
  assign n17467 = ~n17349 & ~n17466;
  assign n17468 = n17349 & n17466;
  assign n17469 = ~n17467 & ~n17468;
  assign n17470 = n16694 & ~n17452;
  assign n17471 = ~n16694 & n17452;
  assign n17472 = ~n17470 & ~n17471;
  assign n17473 = ~n17469 & ~n17472;
  assign n17474 = n17469 & n17472;
  assign n17475 = ~n17473 & ~n17474;
  assign n17476 = ~n17443 & ~n17455;
  assign n17477 = ~n17475 & n17476;
  assign n17478 = n17475 & ~n17476;
  assign n17479 = ~n17477 & ~n17478;
  assign n17480 = ~n17459 & ~n17463;
  assign n17481 = ~n17479 & n17480;
  assign n17482 = n17479 & ~n17480;
  assign po122  = ~n17481 & ~n17482;
  assign n17484 = pi59  & pi63 ;
  assign n17485 = ~n8453 & ~n17484;
  assign n17486 = n8854 & n9123;
  assign n17487 = ~n9054 & ~n17468;
  assign n17488 = ~n17485 & ~n17486;
  assign n17489 = ~n17487 & n17488;
  assign n17490 = ~n17486 & ~n17489;
  assign n17491 = ~n17485 & n17490;
  assign n17492 = ~n17487 & ~n17489;
  assign n17493 = ~n17491 & ~n17492;
  assign n17494 = ~n17470 & ~n17474;
  assign n17495 = n17493 & n17494;
  assign n17496 = ~n17493 & ~n17494;
  assign n17497 = ~n17495 & ~n17496;
  assign n17498 = ~n17478 & ~n17482;
  assign n17499 = ~n17497 & n17498;
  assign n17500 = ~n17495 & ~n17498;
  assign n17501 = ~n17496 & n17500;
  assign po123  = ~n17499 & ~n17501;
  assign n17503 = pi60  & pi63 ;
  assign n17504 = ~pi61  & pi62 ;
  assign n17505 = ~n17503 & ~n17504;
  assign n17506 = n17503 & n17504;
  assign n17507 = ~n17505 & ~n17506;
  assign n17508 = n17490 & ~n17507;
  assign n17509 = ~n17490 & n17507;
  assign n17510 = ~n17508 & ~n17509;
  assign n17511 = ~n17496 & ~n17500;
  assign n17512 = ~n17510 & n17511;
  assign n17513 = n17510 & ~n17511;
  assign po124  = ~n17512 & ~n17513;
  assign n17515 = pi62  & n9236;
  assign n17516 = ~n9236 & ~n9567;
  assign n17517 = ~n17506 & n17516;
  assign n17518 = ~n17515 & ~n17517;
  assign n17519 = ~n17509 & ~n17513;
  assign n17520 = n17518 & ~n17519;
  assign n17521 = ~n17518 & n17519;
  assign po125  = ~n17520 & ~n17521;
  assign n17523 = ~pi62  & pi63 ;
  assign n17524 = ~n17515 & ~n17520;
  assign n17525 = ~n17523 & n17524;
  assign n17526 = n17523 & ~n17524;
  assign po126  = ~n17525 & ~n17526;
  assign po127  = n9123 | n17526;
  assign po1  = 1'b0;
  assign po0  = pi0 ;
endmodule
