module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 , pi132 ,
    pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 , pi140 ,
    pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 , pi148 ,
    pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 , pi156 ,
    pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 , pi164 ,
    pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 , pi172 ,
    pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 , pi180 ,
    pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 , pi188 ,
    pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 , pi196 ,
    pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 , pi204 ,
    pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 , pi212 ,
    pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 , pi220 ,
    pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 ,
    po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 ,
    po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 , po30 , po31 , po32 ,
    po33 , po34 , po35 , po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 , po46 , po47 , po48 ,
    po49 , po50 , po51 , po52 , po53 , po54 , po55 , po56 ,
    po57 , po58 , po59 , po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 , po70 , po71 , po72 ,
    po73 , po74 , po75 , po76 , po77 , po78 , po79 , po80 ,
    po81 , po82 , po83 , po84 , po85 , po86 , po87 , po88 ,
    po89 , po90 , po91 , po92 , po93 , po94 , po95 , po96 ,
    po97 , po98 , po99 , po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 , po108 , po109 , po110 ,
    po111 , po112 , po113 , po114 , po115 , po116 , po117 ,
    po118 , po119 , po120 , po121 , po122 , po123 , po124 ,
    po125 , po126 , po127 , po128  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 ,
    pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 ,
    pi140 , pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 ,
    pi148 , pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 ,
    pi156 , pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 ,
    pi164 , pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 ,
    pi172 , pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 ,
    pi180 , pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 ,
    pi188 , pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 ,
    pi196 , pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 ,
    pi204 , pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 ,
    pi212 , pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 ,
    pi220 , pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 , po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 , po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 , po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 , po100 , po101 , po102 ,
    po103 , po104 , po105 , po106 , po107 , po108 , po109 ,
    po110 , po111 , po112 , po113 , po114 , po115 , po116 ,
    po117 , po118 , po119 , po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 , po128;
  wire n386, n387, n389, n390, n391, n392, n393,
    n394, n396, n397, n398, n399, n400, n401,
    n402, n404, n405, n406, n407, n408, n409,
    n411, n412, n413, n414, n415, n416, n418,
    n419, n420, n421, n422, n423, n425, n426,
    n427, n428, n429, n430, n432, n433, n434,
    n435, n436, n437, n439, n440, n441, n442,
    n443, n444, n446, n447, n448, n449, n450,
    n451, n453, n454, n455, n456, n457, n458,
    n460, n461, n462, n463, n464, n465, n467,
    n468, n469, n470, n471, n472, n474, n475,
    n476, n477, n478, n479, n481, n482, n483,
    n484, n485, n486, n488, n489, n490, n491,
    n492, n493, n495, n496, n497, n498, n499,
    n500, n502, n503, n504, n505, n506, n507,
    n509, n510, n511, n512, n513, n514, n516,
    n517, n518, n519, n520, n521, n523, n524,
    n525, n526, n527, n528, n530, n531, n532,
    n533, n534, n535, n537, n538, n539, n540,
    n541, n542, n544, n545, n546, n547, n548,
    n549, n551, n552, n553, n554, n555, n556,
    n558, n559, n560, n561, n562, n563, n565,
    n566, n567, n568, n569, n570, n572, n573,
    n574, n575, n576, n577, n579, n580, n581,
    n582, n583, n584, n586, n587, n588, n589,
    n590, n591, n593, n594, n595, n596, n597,
    n598, n600, n601, n602, n603, n604, n605,
    n607, n608, n609, n610, n611, n612, n614,
    n615, n616, n617, n618, n619, n621, n622,
    n623, n624, n625, n626, n628, n629, n630,
    n631, n632, n633, n635, n636, n637, n638,
    n639, n640, n642, n643, n644, n645, n646,
    n647, n649, n650, n651, n652, n653, n654,
    n656, n657, n658, n659, n660, n661, n663,
    n664, n665, n666, n667, n668, n670, n671,
    n672, n673, n674, n675, n677, n678, n679,
    n680, n681, n682, n684, n685, n686, n687,
    n688, n689, n691, n692, n693, n694, n695,
    n696, n698, n699, n700, n701, n702, n703,
    n705, n706, n707, n708, n709, n710, n712,
    n713, n714, n715, n716, n717, n719, n720,
    n721, n722, n723, n724, n726, n727, n728,
    n729, n730, n731, n733, n734, n735, n736,
    n737, n738, n740, n741, n742, n743, n744,
    n745, n747, n748, n749, n750, n751, n752,
    n754, n755, n756, n757, n758, n759, n761,
    n762, n763, n764, n765, n766, n768, n769,
    n770, n771, n772, n773, n775, n776, n777,
    n778, n779, n780, n782, n783, n784, n785,
    n786, n787, n789, n790, n791, n792, n793,
    n794, n796, n797, n798, n799, n800, n801,
    n803, n804, n805, n806, n807, n808, n810,
    n811, n812, n813, n814, n815, n817, n818,
    n819, n820, n821, n822, n824, n825, n826,
    n827, n828, n829, n831, n832, n833, n834,
    n835, n836, n838, n839, n840, n841, n842,
    n843, n845, n846, n847, n848, n849, n850,
    n852, n853, n854, n855, n856, n857, n859,
    n860, n861, n862, n863, n864, n866, n867,
    n868, n869, n870, n871, n873, n874, n875,
    n876, n877, n878, n880, n881, n882, n883,
    n884, n885, n887, n888, n889, n890, n891,
    n892, n894, n895, n896, n897, n898, n899,
    n901, n902, n903, n904, n905, n906, n908,
    n909, n910, n911, n912, n913, n915, n916,
    n917, n918, n919, n920, n922, n923, n924,
    n925, n926, n927, n929, n930, n931, n932,
    n933, n934, n936, n937, n938, n939, n940,
    n941, n943, n944, n945, n946, n947, n948,
    n950, n951, n952, n953, n954, n955, n957,
    n958, n959, n960, n961, n962, n964, n965,
    n966, n967, n968, n969, n971, n972, n973,
    n974, n975, n976, n978, n979, n980, n981,
    n982, n983, n985, n986, n987, n988, n989,
    n990, n992, n993, n994, n995, n996, n997,
    n999, n1000, n1001, n1002, n1003, n1004,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1013, n1014, n1015, n1016, n1017, n1018,
    n1020, n1021, n1022, n1023, n1024, n1025,
    n1027, n1028, n1029, n1030, n1031, n1032,
    n1034, n1035, n1036, n1037, n1038, n1039,
    n1041, n1042, n1043, n1044, n1045, n1046,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1055, n1056, n1057, n1058, n1059, n1060,
    n1062, n1063, n1064, n1065, n1066, n1067,
    n1069, n1070, n1071, n1072, n1073, n1074,
    n1076, n1077, n1078, n1079, n1080, n1081,
    n1083, n1084, n1085, n1086, n1087, n1088,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1097, n1098, n1099, n1100, n1101, n1102,
    n1104, n1105, n1106, n1107, n1108, n1109,
    n1111, n1112, n1113, n1114, n1115, n1116,
    n1118, n1119, n1120, n1121, n1122, n1123,
    n1125, n1126, n1127, n1128, n1129, n1130,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1139, n1140, n1141, n1142, n1143, n1144,
    n1146, n1147, n1148, n1149, n1150, n1151,
    n1153, n1154, n1155, n1156, n1157, n1158,
    n1160, n1161, n1162, n1163, n1164, n1165,
    n1167, n1168, n1169, n1170, n1171, n1172,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1181, n1182, n1183, n1184, n1185, n1186,
    n1188, n1189, n1190, n1191, n1192, n1193,
    n1195, n1196, n1197, n1198, n1199, n1200,
    n1202, n1203, n1204, n1205, n1206, n1207,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1216, n1217, n1218, n1219, n1220, n1221,
    n1223, n1224, n1225, n1226, n1227, n1228,
    n1230, n1231, n1232, n1233, n1234, n1235,
    n1237, n1238, n1239, n1240, n1241, n1242,
    n1244, n1245, n1246, n1247, n1248, n1249,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1258, n1259, n1260, n1261, n1262, n1263,
    n1265, n1266, n1267, n1268, n1269, n1270,
    n1272, n1273, n1274, n1275, n1276, n1277;
  assign n386 = pi0  & ~pi128 ;
  assign n387 = ~pi0  & pi128 ;
  assign po0  = n386 | n387;
  assign n389 = pi0  & pi128 ;
  assign n390 = ~pi1  & ~pi129 ;
  assign n391 = pi1  & pi129 ;
  assign n392 = ~n390 & ~n391;
  assign n393 = n389 & ~n392;
  assign n394 = ~n389 & n392;
  assign po1  = n393 | n394;
  assign n396 = n389 & ~n390;
  assign n397 = ~n391 & ~n396;
  assign n398 = ~pi2  & ~pi130 ;
  assign n399 = pi2  & pi130 ;
  assign n400 = ~n398 & ~n399;
  assign n401 = n397 & ~n400;
  assign n402 = ~n397 & n400;
  assign po2  = ~n401 & ~n402;
  assign n404 = ~pi3  & ~pi131 ;
  assign n405 = pi3  & pi131 ;
  assign n406 = ~n404 & ~n405;
  assign n407 = ~n399 & ~n402;
  assign n408 = ~n406 & n407;
  assign n409 = n406 & ~n407;
  assign po3  = ~n408 & ~n409;
  assign n411 = ~pi4  & ~pi132 ;
  assign n412 = pi4  & pi132 ;
  assign n413 = ~n411 & ~n412;
  assign n414 = ~n405 & ~n409;
  assign n415 = ~n413 & n414;
  assign n416 = n413 & ~n414;
  assign po4  = ~n415 & ~n416;
  assign n418 = ~pi5  & ~pi133 ;
  assign n419 = pi5  & pi133 ;
  assign n420 = ~n418 & ~n419;
  assign n421 = ~n412 & ~n416;
  assign n422 = ~n420 & n421;
  assign n423 = n420 & ~n421;
  assign po5  = ~n422 & ~n423;
  assign n425 = ~pi6  & ~pi134 ;
  assign n426 = pi6  & pi134 ;
  assign n427 = ~n425 & ~n426;
  assign n428 = ~n419 & ~n423;
  assign n429 = ~n427 & n428;
  assign n430 = n427 & ~n428;
  assign po6  = ~n429 & ~n430;
  assign n432 = ~pi7  & ~pi135 ;
  assign n433 = pi7  & pi135 ;
  assign n434 = ~n432 & ~n433;
  assign n435 = ~n426 & ~n430;
  assign n436 = ~n434 & n435;
  assign n437 = n434 & ~n435;
  assign po7  = ~n436 & ~n437;
  assign n439 = ~pi8  & ~pi136 ;
  assign n440 = pi8  & pi136 ;
  assign n441 = ~n439 & ~n440;
  assign n442 = ~n433 & ~n437;
  assign n443 = ~n441 & n442;
  assign n444 = n441 & ~n442;
  assign po8  = ~n443 & ~n444;
  assign n446 = ~pi9  & ~pi137 ;
  assign n447 = pi9  & pi137 ;
  assign n448 = ~n446 & ~n447;
  assign n449 = ~n440 & ~n444;
  assign n450 = ~n448 & n449;
  assign n451 = n448 & ~n449;
  assign po9  = ~n450 & ~n451;
  assign n453 = ~pi10  & ~pi138 ;
  assign n454 = pi10  & pi138 ;
  assign n455 = ~n453 & ~n454;
  assign n456 = ~n447 & ~n451;
  assign n457 = ~n455 & n456;
  assign n458 = n455 & ~n456;
  assign po10  = ~n457 & ~n458;
  assign n460 = ~pi11  & ~pi139 ;
  assign n461 = pi11  & pi139 ;
  assign n462 = ~n460 & ~n461;
  assign n463 = ~n454 & ~n458;
  assign n464 = ~n462 & n463;
  assign n465 = n462 & ~n463;
  assign po11  = ~n464 & ~n465;
  assign n467 = ~pi12  & ~pi140 ;
  assign n468 = pi12  & pi140 ;
  assign n469 = ~n467 & ~n468;
  assign n470 = ~n461 & ~n465;
  assign n471 = ~n469 & n470;
  assign n472 = n469 & ~n470;
  assign po12  = ~n471 & ~n472;
  assign n474 = ~pi13  & ~pi141 ;
  assign n475 = pi13  & pi141 ;
  assign n476 = ~n474 & ~n475;
  assign n477 = ~n468 & ~n472;
  assign n478 = ~n476 & n477;
  assign n479 = n476 & ~n477;
  assign po13  = ~n478 & ~n479;
  assign n481 = ~pi14  & ~pi142 ;
  assign n482 = pi14  & pi142 ;
  assign n483 = ~n481 & ~n482;
  assign n484 = ~n475 & ~n479;
  assign n485 = ~n483 & n484;
  assign n486 = n483 & ~n484;
  assign po14  = ~n485 & ~n486;
  assign n488 = ~pi15  & ~pi143 ;
  assign n489 = pi15  & pi143 ;
  assign n490 = ~n488 & ~n489;
  assign n491 = ~n482 & ~n486;
  assign n492 = ~n490 & n491;
  assign n493 = n490 & ~n491;
  assign po15  = ~n492 & ~n493;
  assign n495 = ~pi16  & ~pi144 ;
  assign n496 = pi16  & pi144 ;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~n489 & ~n493;
  assign n499 = ~n497 & n498;
  assign n500 = n497 & ~n498;
  assign po16  = ~n499 & ~n500;
  assign n502 = ~pi17  & ~pi145 ;
  assign n503 = pi17  & pi145 ;
  assign n504 = ~n502 & ~n503;
  assign n505 = ~n496 & ~n500;
  assign n506 = ~n504 & n505;
  assign n507 = n504 & ~n505;
  assign po17  = ~n506 & ~n507;
  assign n509 = ~pi18  & ~pi146 ;
  assign n510 = pi18  & pi146 ;
  assign n511 = ~n509 & ~n510;
  assign n512 = ~n503 & ~n507;
  assign n513 = ~n511 & n512;
  assign n514 = n511 & ~n512;
  assign po18  = ~n513 & ~n514;
  assign n516 = ~pi19  & ~pi147 ;
  assign n517 = pi19  & pi147 ;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~n510 & ~n514;
  assign n520 = ~n518 & n519;
  assign n521 = n518 & ~n519;
  assign po19  = ~n520 & ~n521;
  assign n523 = ~pi20  & ~pi148 ;
  assign n524 = pi20  & pi148 ;
  assign n525 = ~n523 & ~n524;
  assign n526 = ~n517 & ~n521;
  assign n527 = ~n525 & n526;
  assign n528 = n525 & ~n526;
  assign po20  = ~n527 & ~n528;
  assign n530 = ~pi21  & ~pi149 ;
  assign n531 = pi21  & pi149 ;
  assign n532 = ~n530 & ~n531;
  assign n533 = ~n524 & ~n528;
  assign n534 = ~n532 & n533;
  assign n535 = n532 & ~n533;
  assign po21  = ~n534 & ~n535;
  assign n537 = ~pi22  & ~pi150 ;
  assign n538 = pi22  & pi150 ;
  assign n539 = ~n537 & ~n538;
  assign n540 = ~n531 & ~n535;
  assign n541 = ~n539 & n540;
  assign n542 = n539 & ~n540;
  assign po22  = ~n541 & ~n542;
  assign n544 = ~pi23  & ~pi151 ;
  assign n545 = pi23  & pi151 ;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~n538 & ~n542;
  assign n548 = ~n546 & n547;
  assign n549 = n546 & ~n547;
  assign po23  = ~n548 & ~n549;
  assign n551 = ~pi24  & ~pi152 ;
  assign n552 = pi24  & pi152 ;
  assign n553 = ~n551 & ~n552;
  assign n554 = ~n545 & ~n549;
  assign n555 = ~n553 & n554;
  assign n556 = n553 & ~n554;
  assign po24  = ~n555 & ~n556;
  assign n558 = ~pi25  & ~pi153 ;
  assign n559 = pi25  & pi153 ;
  assign n560 = ~n558 & ~n559;
  assign n561 = ~n552 & ~n556;
  assign n562 = ~n560 & n561;
  assign n563 = n560 & ~n561;
  assign po25  = ~n562 & ~n563;
  assign n565 = ~pi26  & ~pi154 ;
  assign n566 = pi26  & pi154 ;
  assign n567 = ~n565 & ~n566;
  assign n568 = ~n559 & ~n563;
  assign n569 = ~n567 & n568;
  assign n570 = n567 & ~n568;
  assign po26  = ~n569 & ~n570;
  assign n572 = ~pi27  & ~pi155 ;
  assign n573 = pi27  & pi155 ;
  assign n574 = ~n572 & ~n573;
  assign n575 = ~n566 & ~n570;
  assign n576 = ~n574 & n575;
  assign n577 = n574 & ~n575;
  assign po27  = ~n576 & ~n577;
  assign n579 = ~pi28  & ~pi156 ;
  assign n580 = pi28  & pi156 ;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~n573 & ~n577;
  assign n583 = ~n581 & n582;
  assign n584 = n581 & ~n582;
  assign po28  = ~n583 & ~n584;
  assign n586 = ~pi29  & ~pi157 ;
  assign n587 = pi29  & pi157 ;
  assign n588 = ~n586 & ~n587;
  assign n589 = ~n580 & ~n584;
  assign n590 = ~n588 & n589;
  assign n591 = n588 & ~n589;
  assign po29  = ~n590 & ~n591;
  assign n593 = ~pi30  & ~pi158 ;
  assign n594 = pi30  & pi158 ;
  assign n595 = ~n593 & ~n594;
  assign n596 = ~n587 & ~n591;
  assign n597 = ~n595 & n596;
  assign n598 = n595 & ~n596;
  assign po30  = ~n597 & ~n598;
  assign n600 = ~pi31  & ~pi159 ;
  assign n601 = pi31  & pi159 ;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~n594 & ~n598;
  assign n604 = ~n602 & n603;
  assign n605 = n602 & ~n603;
  assign po31  = ~n604 & ~n605;
  assign n607 = ~pi32  & ~pi160 ;
  assign n608 = pi32  & pi160 ;
  assign n609 = ~n607 & ~n608;
  assign n610 = ~n601 & ~n605;
  assign n611 = ~n609 & n610;
  assign n612 = n609 & ~n610;
  assign po32  = ~n611 & ~n612;
  assign n614 = ~pi33  & ~pi161 ;
  assign n615 = pi33  & pi161 ;
  assign n616 = ~n614 & ~n615;
  assign n617 = ~n608 & ~n612;
  assign n618 = ~n616 & n617;
  assign n619 = n616 & ~n617;
  assign po33  = ~n618 & ~n619;
  assign n621 = ~pi34  & ~pi162 ;
  assign n622 = pi34  & pi162 ;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~n615 & ~n619;
  assign n625 = ~n623 & n624;
  assign n626 = n623 & ~n624;
  assign po34  = ~n625 & ~n626;
  assign n628 = ~pi35  & ~pi163 ;
  assign n629 = pi35  & pi163 ;
  assign n630 = ~n628 & ~n629;
  assign n631 = ~n622 & ~n626;
  assign n632 = ~n630 & n631;
  assign n633 = n630 & ~n631;
  assign po35  = ~n632 & ~n633;
  assign n635 = ~pi36  & ~pi164 ;
  assign n636 = pi36  & pi164 ;
  assign n637 = ~n635 & ~n636;
  assign n638 = ~n629 & ~n633;
  assign n639 = ~n637 & n638;
  assign n640 = n637 & ~n638;
  assign po36  = ~n639 & ~n640;
  assign n642 = ~pi37  & ~pi165 ;
  assign n643 = pi37  & pi165 ;
  assign n644 = ~n642 & ~n643;
  assign n645 = ~n636 & ~n640;
  assign n646 = ~n644 & n645;
  assign n647 = n644 & ~n645;
  assign po37  = ~n646 & ~n647;
  assign n649 = ~pi38  & ~pi166 ;
  assign n650 = pi38  & pi166 ;
  assign n651 = ~n649 & ~n650;
  assign n652 = ~n643 & ~n647;
  assign n653 = ~n651 & n652;
  assign n654 = n651 & ~n652;
  assign po38  = ~n653 & ~n654;
  assign n656 = ~pi39  & ~pi167 ;
  assign n657 = pi39  & pi167 ;
  assign n658 = ~n656 & ~n657;
  assign n659 = ~n650 & ~n654;
  assign n660 = ~n658 & n659;
  assign n661 = n658 & ~n659;
  assign po39  = ~n660 & ~n661;
  assign n663 = ~pi40  & ~pi168 ;
  assign n664 = pi40  & pi168 ;
  assign n665 = ~n663 & ~n664;
  assign n666 = ~n657 & ~n661;
  assign n667 = ~n665 & n666;
  assign n668 = n665 & ~n666;
  assign po40  = ~n667 & ~n668;
  assign n670 = ~pi41  & ~pi169 ;
  assign n671 = pi41  & pi169 ;
  assign n672 = ~n670 & ~n671;
  assign n673 = ~n664 & ~n668;
  assign n674 = ~n672 & n673;
  assign n675 = n672 & ~n673;
  assign po41  = ~n674 & ~n675;
  assign n677 = ~pi42  & ~pi170 ;
  assign n678 = pi42  & pi170 ;
  assign n679 = ~n677 & ~n678;
  assign n680 = ~n671 & ~n675;
  assign n681 = ~n679 & n680;
  assign n682 = n679 & ~n680;
  assign po42  = ~n681 & ~n682;
  assign n684 = ~pi43  & ~pi171 ;
  assign n685 = pi43  & pi171 ;
  assign n686 = ~n684 & ~n685;
  assign n687 = ~n678 & ~n682;
  assign n688 = ~n686 & n687;
  assign n689 = n686 & ~n687;
  assign po43  = ~n688 & ~n689;
  assign n691 = ~pi44  & ~pi172 ;
  assign n692 = pi44  & pi172 ;
  assign n693 = ~n691 & ~n692;
  assign n694 = ~n685 & ~n689;
  assign n695 = ~n693 & n694;
  assign n696 = n693 & ~n694;
  assign po44  = ~n695 & ~n696;
  assign n698 = ~pi45  & ~pi173 ;
  assign n699 = pi45  & pi173 ;
  assign n700 = ~n698 & ~n699;
  assign n701 = ~n692 & ~n696;
  assign n702 = ~n700 & n701;
  assign n703 = n700 & ~n701;
  assign po45  = ~n702 & ~n703;
  assign n705 = ~pi46  & ~pi174 ;
  assign n706 = pi46  & pi174 ;
  assign n707 = ~n705 & ~n706;
  assign n708 = ~n699 & ~n703;
  assign n709 = ~n707 & n708;
  assign n710 = n707 & ~n708;
  assign po46  = ~n709 & ~n710;
  assign n712 = ~pi47  & ~pi175 ;
  assign n713 = pi47  & pi175 ;
  assign n714 = ~n712 & ~n713;
  assign n715 = ~n706 & ~n710;
  assign n716 = ~n714 & n715;
  assign n717 = n714 & ~n715;
  assign po47  = ~n716 & ~n717;
  assign n719 = ~pi48  & ~pi176 ;
  assign n720 = pi48  & pi176 ;
  assign n721 = ~n719 & ~n720;
  assign n722 = ~n713 & ~n717;
  assign n723 = ~n721 & n722;
  assign n724 = n721 & ~n722;
  assign po48  = ~n723 & ~n724;
  assign n726 = ~pi49  & ~pi177 ;
  assign n727 = pi49  & pi177 ;
  assign n728 = ~n726 & ~n727;
  assign n729 = ~n720 & ~n724;
  assign n730 = ~n728 & n729;
  assign n731 = n728 & ~n729;
  assign po49  = ~n730 & ~n731;
  assign n733 = ~pi50  & ~pi178 ;
  assign n734 = pi50  & pi178 ;
  assign n735 = ~n733 & ~n734;
  assign n736 = ~n727 & ~n731;
  assign n737 = ~n735 & n736;
  assign n738 = n735 & ~n736;
  assign po50  = ~n737 & ~n738;
  assign n740 = ~pi51  & ~pi179 ;
  assign n741 = pi51  & pi179 ;
  assign n742 = ~n740 & ~n741;
  assign n743 = ~n734 & ~n738;
  assign n744 = ~n742 & n743;
  assign n745 = n742 & ~n743;
  assign po51  = ~n744 & ~n745;
  assign n747 = ~pi52  & ~pi180 ;
  assign n748 = pi52  & pi180 ;
  assign n749 = ~n747 & ~n748;
  assign n750 = ~n741 & ~n745;
  assign n751 = ~n749 & n750;
  assign n752 = n749 & ~n750;
  assign po52  = ~n751 & ~n752;
  assign n754 = ~pi53  & ~pi181 ;
  assign n755 = pi53  & pi181 ;
  assign n756 = ~n754 & ~n755;
  assign n757 = ~n748 & ~n752;
  assign n758 = ~n756 & n757;
  assign n759 = n756 & ~n757;
  assign po53  = ~n758 & ~n759;
  assign n761 = ~pi54  & ~pi182 ;
  assign n762 = pi54  & pi182 ;
  assign n763 = ~n761 & ~n762;
  assign n764 = ~n755 & ~n759;
  assign n765 = ~n763 & n764;
  assign n766 = n763 & ~n764;
  assign po54  = ~n765 & ~n766;
  assign n768 = ~pi55  & ~pi183 ;
  assign n769 = pi55  & pi183 ;
  assign n770 = ~n768 & ~n769;
  assign n771 = ~n762 & ~n766;
  assign n772 = ~n770 & n771;
  assign n773 = n770 & ~n771;
  assign po55  = ~n772 & ~n773;
  assign n775 = ~pi56  & ~pi184 ;
  assign n776 = pi56  & pi184 ;
  assign n777 = ~n775 & ~n776;
  assign n778 = ~n769 & ~n773;
  assign n779 = ~n777 & n778;
  assign n780 = n777 & ~n778;
  assign po56  = ~n779 & ~n780;
  assign n782 = ~pi57  & ~pi185 ;
  assign n783 = pi57  & pi185 ;
  assign n784 = ~n782 & ~n783;
  assign n785 = ~n776 & ~n780;
  assign n786 = ~n784 & n785;
  assign n787 = n784 & ~n785;
  assign po57  = ~n786 & ~n787;
  assign n789 = ~pi58  & ~pi186 ;
  assign n790 = pi58  & pi186 ;
  assign n791 = ~n789 & ~n790;
  assign n792 = ~n783 & ~n787;
  assign n793 = ~n791 & n792;
  assign n794 = n791 & ~n792;
  assign po58  = ~n793 & ~n794;
  assign n796 = ~pi59  & ~pi187 ;
  assign n797 = pi59  & pi187 ;
  assign n798 = ~n796 & ~n797;
  assign n799 = ~n790 & ~n794;
  assign n800 = ~n798 & n799;
  assign n801 = n798 & ~n799;
  assign po59  = ~n800 & ~n801;
  assign n803 = ~pi60  & ~pi188 ;
  assign n804 = pi60  & pi188 ;
  assign n805 = ~n803 & ~n804;
  assign n806 = ~n797 & ~n801;
  assign n807 = ~n805 & n806;
  assign n808 = n805 & ~n806;
  assign po60  = ~n807 & ~n808;
  assign n810 = ~pi61  & ~pi189 ;
  assign n811 = pi61  & pi189 ;
  assign n812 = ~n810 & ~n811;
  assign n813 = ~n804 & ~n808;
  assign n814 = ~n812 & n813;
  assign n815 = n812 & ~n813;
  assign po61  = ~n814 & ~n815;
  assign n817 = ~pi62  & ~pi190 ;
  assign n818 = pi62  & pi190 ;
  assign n819 = ~n817 & ~n818;
  assign n820 = ~n811 & ~n815;
  assign n821 = ~n819 & n820;
  assign n822 = n819 & ~n820;
  assign po62  = ~n821 & ~n822;
  assign n824 = ~pi63  & ~pi191 ;
  assign n825 = pi63  & pi191 ;
  assign n826 = ~n824 & ~n825;
  assign n827 = ~n818 & ~n822;
  assign n828 = ~n826 & n827;
  assign n829 = n826 & ~n827;
  assign po63  = ~n828 & ~n829;
  assign n831 = ~pi64  & ~pi192 ;
  assign n832 = pi64  & pi192 ;
  assign n833 = ~n831 & ~n832;
  assign n834 = ~n825 & ~n829;
  assign n835 = ~n833 & n834;
  assign n836 = n833 & ~n834;
  assign po64  = ~n835 & ~n836;
  assign n838 = ~pi65  & ~pi193 ;
  assign n839 = pi65  & pi193 ;
  assign n840 = ~n838 & ~n839;
  assign n841 = ~n832 & ~n836;
  assign n842 = ~n840 & n841;
  assign n843 = n840 & ~n841;
  assign po65  = ~n842 & ~n843;
  assign n845 = ~pi66  & ~pi194 ;
  assign n846 = pi66  & pi194 ;
  assign n847 = ~n845 & ~n846;
  assign n848 = ~n839 & ~n843;
  assign n849 = ~n847 & n848;
  assign n850 = n847 & ~n848;
  assign po66  = ~n849 & ~n850;
  assign n852 = ~pi67  & ~pi195 ;
  assign n853 = pi67  & pi195 ;
  assign n854 = ~n852 & ~n853;
  assign n855 = ~n846 & ~n850;
  assign n856 = ~n854 & n855;
  assign n857 = n854 & ~n855;
  assign po67  = ~n856 & ~n857;
  assign n859 = ~pi68  & ~pi196 ;
  assign n860 = pi68  & pi196 ;
  assign n861 = ~n859 & ~n860;
  assign n862 = ~n853 & ~n857;
  assign n863 = ~n861 & n862;
  assign n864 = n861 & ~n862;
  assign po68  = ~n863 & ~n864;
  assign n866 = ~pi69  & ~pi197 ;
  assign n867 = pi69  & pi197 ;
  assign n868 = ~n866 & ~n867;
  assign n869 = ~n860 & ~n864;
  assign n870 = ~n868 & n869;
  assign n871 = n868 & ~n869;
  assign po69  = ~n870 & ~n871;
  assign n873 = ~pi70  & ~pi198 ;
  assign n874 = pi70  & pi198 ;
  assign n875 = ~n873 & ~n874;
  assign n876 = ~n867 & ~n871;
  assign n877 = ~n875 & n876;
  assign n878 = n875 & ~n876;
  assign po70  = ~n877 & ~n878;
  assign n880 = ~pi71  & ~pi199 ;
  assign n881 = pi71  & pi199 ;
  assign n882 = ~n880 & ~n881;
  assign n883 = ~n874 & ~n878;
  assign n884 = ~n882 & n883;
  assign n885 = n882 & ~n883;
  assign po71  = ~n884 & ~n885;
  assign n887 = ~pi72  & ~pi200 ;
  assign n888 = pi72  & pi200 ;
  assign n889 = ~n887 & ~n888;
  assign n890 = ~n881 & ~n885;
  assign n891 = ~n889 & n890;
  assign n892 = n889 & ~n890;
  assign po72  = ~n891 & ~n892;
  assign n894 = ~pi73  & ~pi201 ;
  assign n895 = pi73  & pi201 ;
  assign n896 = ~n894 & ~n895;
  assign n897 = ~n888 & ~n892;
  assign n898 = ~n896 & n897;
  assign n899 = n896 & ~n897;
  assign po73  = ~n898 & ~n899;
  assign n901 = ~pi74  & ~pi202 ;
  assign n902 = pi74  & pi202 ;
  assign n903 = ~n901 & ~n902;
  assign n904 = ~n895 & ~n899;
  assign n905 = ~n903 & n904;
  assign n906 = n903 & ~n904;
  assign po74  = ~n905 & ~n906;
  assign n908 = ~pi75  & ~pi203 ;
  assign n909 = pi75  & pi203 ;
  assign n910 = ~n908 & ~n909;
  assign n911 = ~n902 & ~n906;
  assign n912 = ~n910 & n911;
  assign n913 = n910 & ~n911;
  assign po75  = ~n912 & ~n913;
  assign n915 = ~pi76  & ~pi204 ;
  assign n916 = pi76  & pi204 ;
  assign n917 = ~n915 & ~n916;
  assign n918 = ~n909 & ~n913;
  assign n919 = ~n917 & n918;
  assign n920 = n917 & ~n918;
  assign po76  = ~n919 & ~n920;
  assign n922 = ~pi77  & ~pi205 ;
  assign n923 = pi77  & pi205 ;
  assign n924 = ~n922 & ~n923;
  assign n925 = ~n916 & ~n920;
  assign n926 = ~n924 & n925;
  assign n927 = n924 & ~n925;
  assign po77  = ~n926 & ~n927;
  assign n929 = ~pi78  & ~pi206 ;
  assign n930 = pi78  & pi206 ;
  assign n931 = ~n929 & ~n930;
  assign n932 = ~n923 & ~n927;
  assign n933 = ~n931 & n932;
  assign n934 = n931 & ~n932;
  assign po78  = ~n933 & ~n934;
  assign n936 = ~pi79  & ~pi207 ;
  assign n937 = pi79  & pi207 ;
  assign n938 = ~n936 & ~n937;
  assign n939 = ~n930 & ~n934;
  assign n940 = ~n938 & n939;
  assign n941 = n938 & ~n939;
  assign po79  = ~n940 & ~n941;
  assign n943 = ~pi80  & ~pi208 ;
  assign n944 = pi80  & pi208 ;
  assign n945 = ~n943 & ~n944;
  assign n946 = ~n937 & ~n941;
  assign n947 = ~n945 & n946;
  assign n948 = n945 & ~n946;
  assign po80  = ~n947 & ~n948;
  assign n950 = ~pi81  & ~pi209 ;
  assign n951 = pi81  & pi209 ;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~n944 & ~n948;
  assign n954 = ~n952 & n953;
  assign n955 = n952 & ~n953;
  assign po81  = ~n954 & ~n955;
  assign n957 = ~pi82  & ~pi210 ;
  assign n958 = pi82  & pi210 ;
  assign n959 = ~n957 & ~n958;
  assign n960 = ~n951 & ~n955;
  assign n961 = ~n959 & n960;
  assign n962 = n959 & ~n960;
  assign po82  = ~n961 & ~n962;
  assign n964 = ~pi83  & ~pi211 ;
  assign n965 = pi83  & pi211 ;
  assign n966 = ~n964 & ~n965;
  assign n967 = ~n958 & ~n962;
  assign n968 = ~n966 & n967;
  assign n969 = n966 & ~n967;
  assign po83  = ~n968 & ~n969;
  assign n971 = ~pi84  & ~pi212 ;
  assign n972 = pi84  & pi212 ;
  assign n973 = ~n971 & ~n972;
  assign n974 = ~n965 & ~n969;
  assign n975 = ~n973 & n974;
  assign n976 = n973 & ~n974;
  assign po84  = ~n975 & ~n976;
  assign n978 = ~pi85  & ~pi213 ;
  assign n979 = pi85  & pi213 ;
  assign n980 = ~n978 & ~n979;
  assign n981 = ~n972 & ~n976;
  assign n982 = ~n980 & n981;
  assign n983 = n980 & ~n981;
  assign po85  = ~n982 & ~n983;
  assign n985 = ~pi86  & ~pi214 ;
  assign n986 = pi86  & pi214 ;
  assign n987 = ~n985 & ~n986;
  assign n988 = ~n979 & ~n983;
  assign n989 = ~n987 & n988;
  assign n990 = n987 & ~n988;
  assign po86  = ~n989 & ~n990;
  assign n992 = ~pi87  & ~pi215 ;
  assign n993 = pi87  & pi215 ;
  assign n994 = ~n992 & ~n993;
  assign n995 = ~n986 & ~n990;
  assign n996 = ~n994 & n995;
  assign n997 = n994 & ~n995;
  assign po87  = ~n996 & ~n997;
  assign n999 = ~pi88  & ~pi216 ;
  assign n1000 = pi88  & pi216 ;
  assign n1001 = ~n999 & ~n1000;
  assign n1002 = ~n993 & ~n997;
  assign n1003 = ~n1001 & n1002;
  assign n1004 = n1001 & ~n1002;
  assign po88  = ~n1003 & ~n1004;
  assign n1006 = ~pi89  & ~pi217 ;
  assign n1007 = pi89  & pi217 ;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = ~n1000 & ~n1004;
  assign n1010 = ~n1008 & n1009;
  assign n1011 = n1008 & ~n1009;
  assign po89  = ~n1010 & ~n1011;
  assign n1013 = ~pi90  & ~pi218 ;
  assign n1014 = pi90  & pi218 ;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = ~n1007 & ~n1011;
  assign n1017 = ~n1015 & n1016;
  assign n1018 = n1015 & ~n1016;
  assign po90  = ~n1017 & ~n1018;
  assign n1020 = ~pi91  & ~pi219 ;
  assign n1021 = pi91  & pi219 ;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n1014 & ~n1018;
  assign n1024 = ~n1022 & n1023;
  assign n1025 = n1022 & ~n1023;
  assign po91  = ~n1024 & ~n1025;
  assign n1027 = ~pi92  & ~pi220 ;
  assign n1028 = pi92  & pi220 ;
  assign n1029 = ~n1027 & ~n1028;
  assign n1030 = ~n1021 & ~n1025;
  assign n1031 = ~n1029 & n1030;
  assign n1032 = n1029 & ~n1030;
  assign po92  = ~n1031 & ~n1032;
  assign n1034 = ~pi93  & ~pi221 ;
  assign n1035 = pi93  & pi221 ;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = ~n1028 & ~n1032;
  assign n1038 = ~n1036 & n1037;
  assign n1039 = n1036 & ~n1037;
  assign po93  = ~n1038 & ~n1039;
  assign n1041 = ~pi94  & ~pi222 ;
  assign n1042 = pi94  & pi222 ;
  assign n1043 = ~n1041 & ~n1042;
  assign n1044 = ~n1035 & ~n1039;
  assign n1045 = ~n1043 & n1044;
  assign n1046 = n1043 & ~n1044;
  assign po94  = ~n1045 & ~n1046;
  assign n1048 = ~pi95  & ~pi223 ;
  assign n1049 = pi95  & pi223 ;
  assign n1050 = ~n1048 & ~n1049;
  assign n1051 = ~n1042 & ~n1046;
  assign n1052 = ~n1050 & n1051;
  assign n1053 = n1050 & ~n1051;
  assign po95  = ~n1052 & ~n1053;
  assign n1055 = ~pi96  & ~pi224 ;
  assign n1056 = pi96  & pi224 ;
  assign n1057 = ~n1055 & ~n1056;
  assign n1058 = ~n1049 & ~n1053;
  assign n1059 = ~n1057 & n1058;
  assign n1060 = n1057 & ~n1058;
  assign po96  = ~n1059 & ~n1060;
  assign n1062 = ~pi97  & ~pi225 ;
  assign n1063 = pi97  & pi225 ;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = ~n1056 & ~n1060;
  assign n1066 = ~n1064 & n1065;
  assign n1067 = n1064 & ~n1065;
  assign po97  = ~n1066 & ~n1067;
  assign n1069 = ~pi98  & ~pi226 ;
  assign n1070 = pi98  & pi226 ;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = ~n1063 & ~n1067;
  assign n1073 = ~n1071 & n1072;
  assign n1074 = n1071 & ~n1072;
  assign po98  = ~n1073 & ~n1074;
  assign n1076 = ~pi99  & ~pi227 ;
  assign n1077 = pi99  & pi227 ;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = ~n1070 & ~n1074;
  assign n1080 = ~n1078 & n1079;
  assign n1081 = n1078 & ~n1079;
  assign po99  = ~n1080 & ~n1081;
  assign n1083 = ~pi100  & ~pi228 ;
  assign n1084 = pi100  & pi228 ;
  assign n1085 = ~n1083 & ~n1084;
  assign n1086 = ~n1077 & ~n1081;
  assign n1087 = ~n1085 & n1086;
  assign n1088 = n1085 & ~n1086;
  assign po100  = ~n1087 & ~n1088;
  assign n1090 = ~pi101  & ~pi229 ;
  assign n1091 = pi101  & pi229 ;
  assign n1092 = ~n1090 & ~n1091;
  assign n1093 = ~n1084 & ~n1088;
  assign n1094 = ~n1092 & n1093;
  assign n1095 = n1092 & ~n1093;
  assign po101  = ~n1094 & ~n1095;
  assign n1097 = ~pi102  & ~pi230 ;
  assign n1098 = pi102  & pi230 ;
  assign n1099 = ~n1097 & ~n1098;
  assign n1100 = ~n1091 & ~n1095;
  assign n1101 = ~n1099 & n1100;
  assign n1102 = n1099 & ~n1100;
  assign po102  = ~n1101 & ~n1102;
  assign n1104 = ~pi103  & ~pi231 ;
  assign n1105 = pi103  & pi231 ;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = ~n1098 & ~n1102;
  assign n1108 = ~n1106 & n1107;
  assign n1109 = n1106 & ~n1107;
  assign po103  = ~n1108 & ~n1109;
  assign n1111 = ~pi104  & ~pi232 ;
  assign n1112 = pi104  & pi232 ;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = ~n1105 & ~n1109;
  assign n1115 = ~n1113 & n1114;
  assign n1116 = n1113 & ~n1114;
  assign po104  = ~n1115 & ~n1116;
  assign n1118 = ~pi105  & ~pi233 ;
  assign n1119 = pi105  & pi233 ;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = ~n1112 & ~n1116;
  assign n1122 = ~n1120 & n1121;
  assign n1123 = n1120 & ~n1121;
  assign po105  = ~n1122 & ~n1123;
  assign n1125 = ~pi106  & ~pi234 ;
  assign n1126 = pi106  & pi234 ;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = ~n1119 & ~n1123;
  assign n1129 = ~n1127 & n1128;
  assign n1130 = n1127 & ~n1128;
  assign po106  = ~n1129 & ~n1130;
  assign n1132 = ~pi107  & ~pi235 ;
  assign n1133 = pi107  & pi235 ;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = ~n1126 & ~n1130;
  assign n1136 = ~n1134 & n1135;
  assign n1137 = n1134 & ~n1135;
  assign po107  = ~n1136 & ~n1137;
  assign n1139 = ~pi108  & ~pi236 ;
  assign n1140 = pi108  & pi236 ;
  assign n1141 = ~n1139 & ~n1140;
  assign n1142 = ~n1133 & ~n1137;
  assign n1143 = ~n1141 & n1142;
  assign n1144 = n1141 & ~n1142;
  assign po108  = ~n1143 & ~n1144;
  assign n1146 = ~pi109  & ~pi237 ;
  assign n1147 = pi109  & pi237 ;
  assign n1148 = ~n1146 & ~n1147;
  assign n1149 = ~n1140 & ~n1144;
  assign n1150 = ~n1148 & n1149;
  assign n1151 = n1148 & ~n1149;
  assign po109  = ~n1150 & ~n1151;
  assign n1153 = ~pi110  & ~pi238 ;
  assign n1154 = pi110  & pi238 ;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156 = ~n1147 & ~n1151;
  assign n1157 = ~n1155 & n1156;
  assign n1158 = n1155 & ~n1156;
  assign po110  = ~n1157 & ~n1158;
  assign n1160 = ~pi111  & ~pi239 ;
  assign n1161 = pi111  & pi239 ;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = ~n1154 & ~n1158;
  assign n1164 = ~n1162 & n1163;
  assign n1165 = n1162 & ~n1163;
  assign po111  = ~n1164 & ~n1165;
  assign n1167 = ~pi112  & ~pi240 ;
  assign n1168 = pi112  & pi240 ;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = ~n1161 & ~n1165;
  assign n1171 = ~n1169 & n1170;
  assign n1172 = n1169 & ~n1170;
  assign po112  = ~n1171 & ~n1172;
  assign n1174 = ~pi113  & ~pi241 ;
  assign n1175 = pi113  & pi241 ;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = ~n1168 & ~n1172;
  assign n1178 = ~n1176 & n1177;
  assign n1179 = n1176 & ~n1177;
  assign po113  = ~n1178 & ~n1179;
  assign n1181 = ~pi114  & ~pi242 ;
  assign n1182 = pi114  & pi242 ;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = ~n1175 & ~n1179;
  assign n1185 = ~n1183 & n1184;
  assign n1186 = n1183 & ~n1184;
  assign po114  = ~n1185 & ~n1186;
  assign n1188 = ~pi115  & ~pi243 ;
  assign n1189 = pi115  & pi243 ;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = ~n1182 & ~n1186;
  assign n1192 = ~n1190 & n1191;
  assign n1193 = n1190 & ~n1191;
  assign po115  = ~n1192 & ~n1193;
  assign n1195 = ~pi116  & ~pi244 ;
  assign n1196 = pi116  & pi244 ;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = ~n1189 & ~n1193;
  assign n1199 = ~n1197 & n1198;
  assign n1200 = n1197 & ~n1198;
  assign po116  = ~n1199 & ~n1200;
  assign n1202 = ~pi117  & ~pi245 ;
  assign n1203 = pi117  & pi245 ;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = ~n1196 & ~n1200;
  assign n1206 = ~n1204 & n1205;
  assign n1207 = n1204 & ~n1205;
  assign po117  = ~n1206 & ~n1207;
  assign n1209 = ~pi118  & ~pi246 ;
  assign n1210 = pi118  & pi246 ;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = ~n1203 & ~n1207;
  assign n1213 = ~n1211 & n1212;
  assign n1214 = n1211 & ~n1212;
  assign po118  = ~n1213 & ~n1214;
  assign n1216 = ~pi119  & ~pi247 ;
  assign n1217 = pi119  & pi247 ;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = ~n1210 & ~n1214;
  assign n1220 = ~n1218 & n1219;
  assign n1221 = n1218 & ~n1219;
  assign po119  = ~n1220 & ~n1221;
  assign n1223 = ~pi120  & ~pi248 ;
  assign n1224 = pi120  & pi248 ;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = ~n1217 & ~n1221;
  assign n1227 = ~n1225 & n1226;
  assign n1228 = n1225 & ~n1226;
  assign po120  = ~n1227 & ~n1228;
  assign n1230 = ~pi121  & ~pi249 ;
  assign n1231 = pi121  & pi249 ;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = ~n1224 & ~n1228;
  assign n1234 = ~n1232 & n1233;
  assign n1235 = n1232 & ~n1233;
  assign po121  = ~n1234 & ~n1235;
  assign n1237 = ~pi122  & ~pi250 ;
  assign n1238 = pi122  & pi250 ;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = ~n1231 & ~n1235;
  assign n1241 = ~n1239 & n1240;
  assign n1242 = n1239 & ~n1240;
  assign po122  = ~n1241 & ~n1242;
  assign n1244 = ~pi123  & ~pi251 ;
  assign n1245 = pi123  & pi251 ;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = ~n1238 & ~n1242;
  assign n1248 = ~n1246 & n1247;
  assign n1249 = n1246 & ~n1247;
  assign po123  = ~n1248 & ~n1249;
  assign n1251 = ~pi124  & ~pi252 ;
  assign n1252 = pi124  & pi252 ;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = ~n1245 & ~n1249;
  assign n1255 = ~n1253 & n1254;
  assign n1256 = n1253 & ~n1254;
  assign po124  = ~n1255 & ~n1256;
  assign n1258 = ~pi125  & ~pi253 ;
  assign n1259 = pi125  & pi253 ;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = ~n1252 & ~n1256;
  assign n1262 = ~n1260 & n1261;
  assign n1263 = n1260 & ~n1261;
  assign po125  = ~n1262 & ~n1263;
  assign n1265 = ~pi126  & ~pi254 ;
  assign n1266 = pi126  & pi254 ;
  assign n1267 = ~n1265 & ~n1266;
  assign n1268 = ~n1259 & ~n1263;
  assign n1269 = ~n1267 & n1268;
  assign n1270 = n1267 & ~n1268;
  assign po126  = ~n1269 & ~n1270;
  assign n1272 = ~pi127  & ~pi255 ;
  assign n1273 = pi127  & pi255 ;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = ~n1266 & ~n1270;
  assign n1276 = ~n1274 & n1275;
  assign n1277 = n1274 & ~n1275;
  assign po127  = ~n1276 & ~n1277;
  assign po128 = n1273 | n1277;
endmodule
