module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 ,
    pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 ,
    pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 ,
    pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 ,
    pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 ,
    pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 ,
    pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 ,
    pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 ,
    pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 ,
    pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 ,
    pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 ,
    pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 ,
    pi108 , pi109 , pi110 , pi111 ,
    pi112 , pi113 , pi114 , pi115 ,
    pi116 , pi117 , pi118 , pi119 ,
    pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ,
    pi128 , pi129 , pi130 , pi131 , pi132 , pi133 , pi134 ,
    pi135 , pi136 , pi137 , pi138 , pi139 , pi140 ,
    pi141 , pi142 , pi143 , pi144 , pi145 , pi146 ,
    pi147 , pi148 , pi149 , pi150 , pi151 , pi152 ,
    pi153 , pi154 , pi155 , pi156 , pi157 , pi158 ,
    pi159 , pi160 , pi161 , pi162 , pi163 , pi164 ,
    pi165 , pi166 , pi167 , pi168 , pi169 , pi170 ,
    pi171 , pi172 , pi173 , pi174 , pi175 , pi176 ,
    pi177 , pi178 , pi179 , pi180 , pi181 , pi182 ,
    pi183 , pi184 , pi185 , pi186 , pi187 , pi188 ,
    pi189 , pi190 , pi191 , pi192 , pi193 , pi194 ,
    pi195 , pi196 , pi197 , pi198 , pi199 , pi200 ,
    pi201 , pi202 , pi203 , pi204 , pi205 , pi206 ,
    pi207 , pi208 , pi209 , pi210 , pi211 , pi212 ,
    pi213 , pi214 , pi215 , pi216 , pi217 , pi218 ,
    pi219 , pi220 , pi221 , pi222 , pi223 , pi224 ,
    pi225 , pi226 , pi227 , pi228 , pi229 , pi230 ,
    pi231 , pi232 , pi233 , pi234 , pi235 , pi236 ,
    pi237 , pi238 , pi239 , pi240 , pi241 , pi242 ,
    pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 ,
    pi255 ,
    po0 , po1 , po2 , po3 , po4 , po5 ,
    po6 , po7 , po8 , po9 , po10 ,
    po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 ,
    po21 , po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 , po30 ,
    po31 , po32 , po33 , po34 , po35 ,
    po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 ,
    po46 , po47 , po48 , po49 , po50 ,
    po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 ,
    po61 , po62 , po63 , po64 , po65 ,
    po66 , po67 , po68 , po69 , po70 ,
    po71 , po72 , po73 , po74 , po75 ,
    po76 , po77 , po78 , po79 , po80 ,
    po81 , po82 , po83 , po84 , po85 ,
    po86 , po87 , po88 , po89 , po90 ,
    po91 , po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 , po100 ,
    po101 , po102 , po103 , po104 , po105 ,
    po106 , po107 , po108 , po109 , po110 ,
    po111 , po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 , po120 ,
    po121 , po122 , po123 , po124 , po125 ,
    po126 , po127 , po128  );
  input  pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 ,
    pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 ,
    pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 ,
    pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 ,
    pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 ,
    pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 ,
    pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 ,
    pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 ,
    pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 ,
    pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 ,
    pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 ,
    pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 ,
    pi108 , pi109 , pi110 , pi111 ,
    pi112 , pi113 , pi114 , pi115 ,
    pi116 , pi117 , pi118 , pi119 ,
    pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ,
    pi128 , pi129 , pi130 , pi131 , pi132 , pi133 , pi134 ,
    pi135 , pi136 , pi137 , pi138 , pi139 , pi140 ,
    pi141 , pi142 , pi143 , pi144 , pi145 , pi146 ,
    pi147 , pi148 , pi149 , pi150 , pi151 , pi152 ,
    pi153 , pi154 , pi155 , pi156 , pi157 , pi158 ,
    pi159 , pi160 , pi161 , pi162 , pi163 , pi164 ,
    pi165 , pi166 , pi167 , pi168 , pi169 , pi170 ,
    pi171 , pi172 , pi173 , pi174 , pi175 , pi176 ,
    pi177 , pi178 , pi179 , pi180 , pi181 , pi182 ,
    pi183 , pi184 , pi185 , pi186 , pi187 , pi188 ,
    pi189 , pi190 , pi191 , pi192 , pi193 , pi194 ,
    pi195 , pi196 , pi197 , pi198 , pi199 , pi200 ,
    pi201 , pi202 , pi203 , pi204 , pi205 , pi206 ,
    pi207 , pi208 , pi209 , pi210 , pi211 , pi212 ,
    pi213 , pi214 , pi215 , pi216 , pi217 , pi218 ,
    pi219 , pi220 , pi221 , pi222 , pi223 , pi224 ,
    pi225 , pi226 , pi227 , pi228 , pi229 , pi230 ,
    pi231 , pi232 , pi233 , pi234 , pi235 , pi236 ,
    pi237 , pi238 , pi239 , pi240 , pi241 , pi242 ,
    pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 ,
    pi255 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 , po104 ,
    po105 , po106 , po107 , po108 , po109 ,
    po110 , po111 , po112 , po113 , po114 ,
    po115 , po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 , po124 ,
    po125 , po126 , po127 , po128;
  wire n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511,
    n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925,
    n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988,
    n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061,
    n1062, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182,
    n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302,
    n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411,
    n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441,
    n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471,
    n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489,
    n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1668, n1669, n1670, n1671, n1672,
    n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702,
    n1703, n1704, n1705, n1706, n1707, n1708,
    n1709, n1710, n1711, n1712, n1713, n1714,
    n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726,
    n1727, n1728, n1729, n1730, n1731, n1732,
    n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1740, n1741, n1742, n1743, n1744,
    n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781,
    n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1811,
    n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823,
    n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926,
    n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951,
    n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981,
    n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2186, n2187, n2188,
    n2189, n2190, n2191, n2192, n2193, n2194,
    n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206,
    n2207, n2208, n2209, n2210, n2211, n2212,
    n2213, n2214, n2215, n2216, n2217, n2218,
    n2219, n2220, n2221, n2222, n2223, n2224,
    n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236,
    n2237, n2238, n2239, n2240, n2241, n2242,
    n2243, n2244, n2245, n2246, n2247, n2248,
    n2249, n2250, n2251, n2252, n2253, n2254,
    n2255, n2256, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266,
    n2267, n2268, n2269, n2270, n2272, n2273,
    n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291,
    n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303,
    n2304, n2305, n2306, n2307, n2308, n2309,
    n2310, n2311, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321,
    n2322, n2323, n2324, n2325, n2326, n2327,
    n2328, n2329, n2330, n2331, n2332, n2333,
    n2334, n2335, n2336, n2337, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351,
    n2352, n2353, n2354, n2355, n2356, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376,
    n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388,
    n2389, n2390, n2391, n2392, n2393, n2394,
    n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406,
    n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424,
    n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436,
    n2437, n2438, n2439, n2440, n2441, n2442,
    n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461,
    n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521,
    n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2702, n2703, n2704,
    n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716,
    n2717, n2718, n2719, n2720, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734,
    n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746,
    n2747, n2748, n2749, n2750, n2751, n2752,
    n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764,
    n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801,
    n2802, n2803, n2804, n2805, n2806, n2807,
    n2808, n2809, n2810, n2811, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831,
    n2832, n2833, n2834, n2835, n2836, n2837,
    n2838, n2839, n2840, n2841, n2842, n2843,
    n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861,
    n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904,
    n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2956, n2957, n2958,
    n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971,
    n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001,
    n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013,
    n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031,
    n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056,
    n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092,
    n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3218, n3219, n3220,
    n3221, n3222, n3223, n3224, n3225, n3226,
    n3227, n3228, n3229, n3230, n3231, n3232,
    n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244,
    n3245, n3246, n3247, n3248, n3249, n3250,
    n3251, n3252, n3253, n3254, n3255, n3256,
    n3257, n3258, n3259, n3260, n3261, n3262,
    n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274,
    n3275, n3276, n3277, n3278, n3279, n3280,
    n3281, n3282, n3283, n3284, n3285, n3286,
    n3287, n3288, n3289, n3290, n3291, n3292,
    n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3302, n3304, n3305,
    n3306, n3307, n3308, n3309, n3310, n3311,
    n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3321, n3322, n3323,
    n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335,
    n3336, n3337, n3338, n3339, n3340, n3341,
    n3342, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353,
    n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365,
    n3366, n3367, n3368, n3369, n3370, n3371,
    n3372, n3373, n3374, n3375, n3376, n3377,
    n3378, n3379, n3380, n3381, n3382, n3383,
    n3384, n3385, n3386, n3387, n3388, n3390,
    n3391, n3392, n3393, n3394, n3395, n3396,
    n3397, n3398, n3399, n3400, n3401, n3402,
    n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414,
    n3415, n3416, n3417, n3418, n3419, n3420,
    n3421, n3422, n3423, n3424, n3425, n3426,
    n3427, n3428, n3429, n3430, n3431, n3432,
    n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444,
    n3445, n3446, n3447, n3448, n3449, n3450,
    n3451, n3452, n3453, n3454, n3455, n3456,
    n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535,
    n3536, n3537, n3538, n3539, n3540, n3541,
    n3542, n3543, n3544, n3545, n3546, n3547,
    n3548, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3648, n3649, n3650, n3651,
    n3652, n3653, n3654, n3655, n3656, n3657,
    n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681,
    n3682, n3683, n3684, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3734, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742,
    n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772,
    n3773, n3774, n3775, n3776, n3777, n3778,
    n3779, n3780, n3781, n3782, n3783, n3784,
    n3785, n3786, n3787, n3788, n3789, n3790,
    n3791, n3792, n3793, n3794, n3795, n3796,
    n3797, n3798, n3799, n3800, n3801, n3802,
    n3803, n3804, n3805, n3806, n3807, n3808,
    n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818, n3820, n3821,
    n3822, n3823, n3824, n3825, n3826, n3827,
    n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3842, n3843, n3844, n3845,
    n3846, n3847, n3848, n3849, n3850, n3851,
    n3852, n3853, n3854, n3855, n3856, n3857,
    n3858, n3859, n3860, n3861, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881,
    n3882, n3883, n3884, n3885, n3886, n3887,
    n3888, n3889, n3890, n3891, n3892, n3893,
    n3894, n3895, n3896, n3897, n3898, n3899,
    n3900, n3901, n3902, n3903, n3904, n3906,
    n3907, n3908, n3909, n3910, n3911, n3912,
    n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924,
    n3925, n3926, n3927, n3928, n3929, n3930,
    n3931, n3932, n3933, n3934, n3935, n3936,
    n3937, n3938, n3939, n3940, n3941, n3942,
    n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954,
    n3955, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966,
    n3967, n3968, n3969, n3970, n3971, n3972,
    n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990,
    n3992, n3993, n3994, n3995, n3996, n3997,
    n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027,
    n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057,
    n4058, n4059, n4060, n4061, n4062, n4063,
    n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4078, n4079, n4080, n4081, n4082,
    n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4164, n4165, n4166, n4167,
    n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191,
    n4192, n4193, n4194, n4195, n4196, n4197,
    n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227,
    n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4250, n4251, n4252,
    n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264,
    n4265, n4266, n4267, n4268, n4269, n4270,
    n4271, n4272, n4273, n4274, n4275, n4276,
    n4277, n4278, n4279, n4280, n4281, n4282,
    n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294,
    n4295, n4296, n4297, n4298, n4299, n4300,
    n4301, n4302, n4303, n4304, n4305, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312,
    n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324,
    n4325, n4326, n4327, n4328, n4329, n4330,
    n4331, n4332, n4333, n4334, n4336, n4337,
    n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367,
    n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385,
    n4386, n4387, n4388, n4389, n4390, n4391,
    n4392, n4393, n4394, n4395, n4396, n4397,
    n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415,
    n4416, n4417, n4418, n4419, n4420, n4422,
    n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476,
    n4477, n4478, n4479, n4480, n4481, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4508, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525,
    n4526, n4527, n4528, n4529, n4530, n4531,
    n4532, n4533, n4534, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622,
    n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4680, n4681, n4682, n4683,
    n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707,
    n4708, n4709, n4710, n4711, n4712, n4713,
    n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737,
    n4738, n4739, n4740, n4741, n4742, n4743,
    n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761,
    n4762, n4763, n4764, n4766, n4767, n4768,
    n4769, n4770, n4771, n4772, n4773, n4774,
    n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786,
    n4787, n4788, n4789, n4790, n4791, n4792,
    n4793, n4794, n4795, n4796, n4797, n4798,
    n4799, n4800, n4801, n4802, n4803, n4804,
    n4805, n4806, n4807, n4808, n4809, n4810,
    n4811, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822,
    n4823, n4824, n4825, n4826, n4827, n4828,
    n4829, n4830, n4831, n4832, n4833, n4834,
    n4835, n4836, n4837, n4838, n4839, n4840,
    n4841, n4842, n4843, n4844, n4845, n4846,
    n4847, n4848, n4849, n4850, n4852, n4853,
    n4854, n4855, n4856, n4857, n4858, n4859,
    n4860, n4861, n4862, n4863, n4864, n4865,
    n4866, n4867, n4868, n4869, n4870, n4871,
    n4872, n4873, n4874, n4875, n4876, n4877,
    n4878, n4879, n4880, n4881, n4882, n4883,
    n4884, n4885, n4886, n4887, n4888, n4889,
    n4890, n4891, n4892, n4893, n4894, n4895,
    n4896, n4897, n4898, n4899, n4900, n4901,
    n4902, n4903, n4904, n4905, n4906, n4907,
    n4908, n4909, n4910, n4911, n4912, n4913,
    n4914, n4915, n4916, n4917, n4918, n4919,
    n4920, n4921, n4922, n4923, n4924, n4925,
    n4926, n4927, n4928, n4929, n4930, n4931,
    n4932, n4933, n4934, n4935, n4936, n4938,
    n4939, n4940, n4941, n4942, n4943, n4944,
    n4945, n4946, n4947, n4948, n4949, n4950,
    n4951, n4952, n4953, n4954, n4955, n4956,
    n4957, n4958, n4959, n4960, n4961, n4962,
    n4963, n4964, n4965, n4966, n4967, n4968,
    n4969, n4970, n4971, n4972, n4973, n4974,
    n4975, n4976, n4977, n4978, n4979, n4980,
    n4981, n4982, n4983, n4984, n4985, n4986,
    n4987, n4988, n4989, n4990, n4991, n4992,
    n4993, n4994, n4995, n4996, n4997, n4998,
    n4999, n5000, n5001, n5002, n5003, n5004,
    n5005, n5006, n5007, n5008, n5009, n5010,
    n5011, n5012, n5013, n5014, n5015, n5016,
    n5017, n5018, n5019, n5020, n5021, n5022,
    n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101,
    n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211,
    n5212, n5213, n5214, n5215, n5216, n5217,
    n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241,
    n5242, n5243, n5244, n5245, n5246, n5247,
    n5248, n5249, n5250, n5251, n5252, n5253,
    n5254, n5255, n5256, n5257, n5258, n5259,
    n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271,
    n5272, n5273, n5274, n5275, n5276, n5277,
    n5278, n5279, n5280, n5282, n5283, n5284,
    n5285, n5286, n5287, n5288, n5289, n5290,
    n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302,
    n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314,
    n5315, n5316, n5317, n5318, n5319, n5320,
    n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332,
    n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5344,
    n5345, n5346, n5347, n5348, n5349, n5350,
    n5351, n5352, n5353, n5354, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362,
    n5363, n5364, n5365, n5366, n5368, n5369,
    n5370, n5371, n5372, n5373, n5374, n5375,
    n5376, n5377, n5378, n5379, n5380, n5381,
    n5382, n5383, n5384, n5385, n5386, n5387,
    n5388, n5389, n5390, n5391, n5392, n5393,
    n5394, n5395, n5396, n5397, n5398, n5399,
    n5400, n5401, n5402, n5403, n5404, n5405,
    n5406, n5407, n5408, n5409, n5410, n5411,
    n5412, n5413, n5414, n5415, n5416, n5417,
    n5418, n5419, n5420, n5421, n5422, n5423,
    n5424, n5425, n5426, n5427, n5428, n5429,
    n5430, n5431, n5432, n5433, n5434, n5435,
    n5436, n5437, n5438, n5439, n5440, n5441,
    n5442, n5443, n5444, n5445, n5446, n5447,
    n5448, n5449, n5450, n5451, n5452, n5454,
    n5455, n5456, n5457, n5458, n5459, n5460,
    n5461, n5462, n5463, n5464, n5465, n5466,
    n5467, n5468, n5469, n5470, n5471, n5472,
    n5473, n5474, n5475, n5476, n5477, n5478,
    n5479, n5480, n5481, n5482, n5483, n5484,
    n5485, n5486, n5487, n5488, n5489, n5490,
    n5491, n5492, n5493, n5494, n5495, n5496,
    n5497, n5498, n5499, n5500, n5501, n5502,
    n5503, n5504, n5505, n5506, n5507, n5508,
    n5509, n5510, n5511, n5512, n5513, n5514,
    n5515, n5516, n5517, n5518, n5519, n5520,
    n5521, n5522, n5523, n5524, n5525, n5526,
    n5527, n5528, n5529, n5530, n5531, n5532,
    n5533, n5534, n5535, n5536, n5537, n5538,
    n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551,
    n5552, n5553, n5554, n5555, n5556, n5557,
    n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581,
    n5582, n5583, n5584, n5585, n5586, n5587,
    n5588, n5589, n5590, n5591, n5592, n5593,
    n5594, n5595, n5596, n5597, n5598, n5599,
    n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611,
    n5612, n5613, n5614, n5615, n5616, n5617,
    n5618, n5619, n5620, n5621, n5622, n5623,
    n5624, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636,
    n5637, n5638, n5639, n5640, n5641, n5642,
    n5643, n5644, n5645, n5646, n5647, n5648,
    n5649, n5650, n5651, n5652, n5653, n5654,
    n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666,
    n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678,
    n5679, n5680, n5681, n5682, n5683, n5684,
    n5685, n5686, n5687, n5688, n5689, n5690,
    n5691, n5692, n5693, n5694, n5695, n5696,
    n5697, n5698, n5699, n5700, n5701, n5702,
    n5703, n5704, n5705, n5706, n5707, n5708,
    n5709, n5710, n5712, n5713, n5714, n5715,
    n5716, n5717, n5718, n5719, n5720, n5721,
    n5722, n5723, n5724, n5725, n5726, n5727,
    n5728, n5729, n5730, n5731, n5732, n5733,
    n5734, n5735, n5736, n5737, n5738, n5739,
    n5740, n5741, n5742, n5743, n5744, n5745,
    n5746, n5747, n5748, n5749, n5750, n5751,
    n5752, n5753, n5754, n5755, n5756, n5757,
    n5758, n5759, n5760, n5761, n5762, n5763,
    n5764, n5765, n5766, n5767, n5768, n5769,
    n5770, n5771, n5772, n5773, n5774, n5775,
    n5776, n5777, n5778, n5779, n5780, n5781,
    n5782, n5783, n5784, n5785, n5786, n5787,
    n5788, n5789, n5790, n5791, n5792, n5793,
    n5794, n5795, n5796, n5798, n5799, n5800,
    n5801, n5802, n5803, n5804, n5805, n5806,
    n5807, n5808, n5809, n5810, n5811, n5812,
    n5813, n5814, n5815, n5816, n5817, n5818,
    n5819, n5820, n5821, n5822, n5823, n5824,
    n5825, n5826, n5827, n5828, n5829, n5830,
    n5831, n5832, n5833, n5834, n5835, n5836,
    n5837, n5838, n5839, n5840, n5841, n5842,
    n5843, n5844, n5845, n5846, n5847, n5848,
    n5849, n5850, n5851, n5852, n5853, n5854,
    n5855, n5856, n5857, n5858, n5859, n5860,
    n5861, n5862, n5863, n5864, n5865, n5866,
    n5867, n5868, n5869, n5870, n5871, n5872,
    n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5884, n5885,
    n5886, n5887, n5888, n5889, n5890, n5891,
    n5892, n5893, n5894, n5895, n5896, n5897,
    n5898, n5899, n5900, n5901, n5902, n5903,
    n5904, n5905, n5906, n5907, n5908, n5909,
    n5910, n5911, n5912, n5913, n5914, n5915,
    n5916, n5917, n5918, n5919, n5920, n5921,
    n5922, n5923, n5924, n5925, n5926, n5927,
    n5928, n5929, n5930, n5931, n5932, n5933,
    n5934, n5935, n5936, n5937, n5938, n5939,
    n5940, n5941, n5942, n5943, n5944, n5945,
    n5946, n5947, n5948, n5949, n5950, n5951,
    n5952, n5953, n5954, n5955, n5956, n5957,
    n5958, n5959, n5960, n5961, n5962, n5963,
    n5964, n5965, n5966, n5967, n5968, n5970,
    n5971, n5972, n5973, n5974, n5975, n5976,
    n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994,
    n5995, n5996, n5997, n5998, n5999, n6000,
    n6001, n6002, n6003, n6004, n6005, n6006,
    n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6022, n6023, n6024,
    n6025, n6026, n6027, n6028, n6029, n6030,
    n6031, n6032, n6033, n6034, n6035, n6036,
    n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054,
    n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067,
    n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079,
    n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097,
    n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6126, n6127,
    n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170,
    n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6228, n6229, n6230, n6231,
    n6232, n6233, n6234, n6235, n6236, n6237,
    n6238, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255,
    n6256, n6257, n6258, n6259, n6260, n6261,
    n6262, n6263, n6264, n6265, n6266, n6267,
    n6268, n6269, n6270, n6271, n6272, n6273,
    n6274, n6275, n6276, n6277, n6278, n6279,
    n6280, n6281, n6282, n6283, n6284, n6285,
    n6286, n6287, n6288, n6289, n6290, n6291,
    n6292, n6293, n6294, n6295, n6296, n6297,
    n6298, n6299, n6300, n6301, n6302, n6303,
    n6304, n6305, n6306, n6307, n6308, n6309,
    n6310, n6311, n6312, n6314, n6315, n6316,
    n6317, n6318, n6319, n6320, n6321, n6322,
    n6323, n6324, n6325, n6326, n6327, n6328,
    n6329, n6330, n6331, n6332, n6333, n6334,
    n6335, n6336, n6337, n6338, n6339, n6340,
    n6341, n6342, n6343, n6344, n6345, n6346,
    n6347, n6348, n6349, n6350, n6351, n6352,
    n6353, n6354, n6355, n6356, n6357, n6358,
    n6359, n6360, n6361, n6362, n6363, n6364,
    n6365, n6366, n6367, n6368, n6369, n6370,
    n6371, n6372, n6373, n6374, n6375, n6376,
    n6377, n6378, n6379, n6380, n6381, n6382,
    n6383, n6384, n6385, n6386, n6387, n6388,
    n6389, n6390, n6391, n6392, n6393, n6394,
    n6395, n6396, n6397, n6398, n6400, n6401,
    n6402, n6403, n6404, n6405, n6406, n6407,
    n6408, n6409, n6410, n6411, n6412, n6413,
    n6414, n6415, n6416, n6417, n6418, n6419,
    n6420, n6421, n6422, n6423, n6424, n6425,
    n6426, n6427, n6428, n6429, n6430, n6431,
    n6432, n6433, n6434, n6435, n6436, n6437,
    n6438, n6439, n6440, n6441, n6442, n6443,
    n6444, n6445, n6446, n6447, n6448, n6449,
    n6450, n6451, n6452, n6453, n6454, n6455,
    n6456, n6457, n6458, n6459, n6460, n6461,
    n6462, n6463, n6464, n6465, n6466, n6467,
    n6468, n6469, n6470, n6471, n6472, n6473,
    n6474, n6475, n6476, n6477, n6478, n6479,
    n6480, n6481, n6482, n6483, n6484, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546,
    n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558,
    n6559, n6560, n6561, n6562, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570,
    n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601,
    n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631,
    n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649,
    n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6744, n6745, n6746, n6747,
    n6748, n6749, n6750, n6751, n6752, n6753,
    n6754, n6755, n6756, n6757, n6758, n6759,
    n6760, n6761, n6762, n6763, n6764, n6765,
    n6766, n6767, n6768, n6769, n6770, n6771,
    n6772, n6773, n6774, n6775, n6776, n6777,
    n6778, n6779, n6780, n6781, n6782, n6783,
    n6784, n6785, n6786, n6787, n6788, n6789,
    n6790, n6791, n6792, n6793, n6794, n6795,
    n6796, n6797, n6798, n6799, n6800, n6801,
    n6802, n6803, n6804, n6805, n6806, n6807,
    n6808, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6830, n6831, n6832,
    n6833, n6834, n6835, n6836, n6837, n6838,
    n6839, n6840, n6841, n6842, n6843, n6844,
    n6845, n6846, n6847, n6848, n6849, n6850,
    n6851, n6852, n6853, n6854, n6855, n6856,
    n6857, n6858, n6859, n6860, n6861, n6862,
    n6863, n6864, n6865, n6866, n6867, n6868,
    n6869, n6870, n6871, n6872, n6873, n6874,
    n6875, n6876, n6877, n6878, n6879, n6880,
    n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n6891, n6892,
    n6893, n6894, n6895, n6896, n6897, n6898,
    n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6916, n6917,
    n6918, n6919, n6920, n6921, n6922, n6923,
    n6924, n6925, n6926, n6927, n6928, n6929,
    n6930, n6931, n6932, n6933, n6934, n6935,
    n6936, n6937, n6938, n6939, n6940, n6941,
    n6942, n6943, n6944, n6945, n6946, n6947,
    n6948, n6949, n6950, n6951, n6952, n6953,
    n6954, n6955, n6956, n6957, n6958, n6959,
    n6960, n6961, n6962, n6963, n6964, n6965,
    n6966, n6967, n6968, n6969, n6970, n6971,
    n6972, n6973, n6974, n6975, n6976, n6977,
    n6978, n6979, n6980, n6981, n6982, n6983,
    n6984, n6985, n6986, n6987, n6988, n6989,
    n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7002,
    n7003, n7004, n7005, n7006, n7007, n7008,
    n7009, n7010, n7011, n7012, n7013, n7014,
    n7015, n7016, n7017, n7018, n7019, n7020,
    n7021, n7022, n7023, n7024, n7025, n7026,
    n7027, n7028, n7029, n7030, n7031, n7032,
    n7033, n7034, n7035, n7036, n7037, n7038,
    n7039, n7040, n7041, n7042, n7043, n7044,
    n7045, n7046, n7047, n7048, n7049, n7050,
    n7051, n7052, n7053, n7054, n7055, n7056,
    n7057, n7058, n7059, n7060, n7061, n7062,
    n7063, n7064, n7065, n7066, n7067, n7068,
    n7069, n7070, n7071, n7072, n7073, n7074,
    n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086,
    n7088, n7089, n7090, n7091, n7092, n7093,
    n7094, n7095, n7096, n7097, n7098, n7099,
    n7100, n7101, n7102, n7103, n7104, n7105,
    n7106, n7107, n7108, n7109, n7110, n7111,
    n7112, n7113, n7114, n7115, n7116, n7117,
    n7118, n7119, n7120, n7121, n7122, n7123,
    n7124, n7125, n7126, n7127, n7128, n7129,
    n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7137, n7138, n7139, n7140, n7141,
    n7142, n7143, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153,
    n7154, n7155, n7156, n7157, n7158, n7159,
    n7160, n7161, n7162, n7163, n7164, n7165,
    n7166, n7167, n7168, n7169, n7170, n7171,
    n7172, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202,
    n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214,
    n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7260, n7261, n7262, n7263,
    n7264, n7265, n7266, n7267, n7268, n7269,
    n7270, n7271, n7272, n7273, n7274, n7275,
    n7276, n7277, n7278, n7279, n7280, n7281,
    n7282, n7283, n7284, n7285, n7286, n7287,
    n7288, n7289, n7290, n7291, n7292, n7293,
    n7294, n7295, n7296, n7297, n7298, n7299,
    n7300, n7301, n7302, n7303, n7304, n7305,
    n7306, n7307, n7308, n7309, n7310, n7311,
    n7312, n7313, n7314, n7315, n7316, n7317,
    n7318, n7319, n7320, n7321, n7322, n7323,
    n7324, n7325, n7326, n7327, n7328, n7329,
    n7330, n7331, n7332, n7333, n7334, n7335,
    n7336, n7337, n7338, n7339, n7340, n7341,
    n7342, n7343, n7344, n7346, n7347, n7348,
    n7349, n7350, n7351, n7352, n7353, n7354,
    n7355, n7356, n7357, n7358, n7359, n7360,
    n7361, n7362, n7363, n7364, n7365, n7366,
    n7367, n7368, n7369, n7370, n7371, n7372,
    n7373, n7374, n7375, n7376, n7377, n7378,
    n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390,
    n7391, n7392, n7393, n7394, n7395, n7396,
    n7397, n7398, n7399, n7400, n7401, n7402,
    n7403, n7404, n7405, n7406, n7407, n7408,
    n7409, n7410, n7411, n7412, n7413, n7414,
    n7415, n7416, n7417, n7418, n7419, n7420,
    n7421, n7422, n7423, n7424, n7425, n7426,
    n7427, n7428, n7429, n7430, n7432, n7433,
    n7434, n7435, n7436, n7437, n7438, n7439,
    n7440, n7441, n7442, n7443, n7444, n7445,
    n7446, n7447, n7448, n7449, n7450, n7451,
    n7452, n7453, n7454, n7455, n7456, n7457,
    n7458, n7459, n7460, n7461, n7462, n7463,
    n7464, n7465, n7466, n7467, n7468, n7469,
    n7470, n7471, n7472, n7473, n7474, n7475,
    n7476, n7477, n7478, n7479, n7480, n7481,
    n7482, n7483, n7484, n7485, n7486, n7487,
    n7488, n7489, n7490, n7491, n7492, n7493,
    n7494, n7495, n7496, n7497, n7498, n7499,
    n7500, n7501, n7502, n7503, n7504, n7505,
    n7506, n7507, n7508, n7509, n7510, n7511,
    n7512, n7513, n7514, n7515, n7516, n7518,
    n7519, n7520, n7521, n7522, n7523, n7524,
    n7525, n7526, n7527, n7528, n7529, n7530,
    n7531, n7532, n7533, n7534, n7535, n7536,
    n7537, n7538, n7539, n7540, n7541, n7542,
    n7543, n7544, n7545, n7546, n7547, n7548,
    n7549, n7550, n7551, n7552, n7553, n7554,
    n7555, n7556, n7557, n7558, n7559, n7560,
    n7561, n7562, n7563, n7564, n7565, n7566,
    n7567, n7568, n7569, n7570, n7571, n7572,
    n7573, n7574, n7575, n7576, n7577, n7578,
    n7579, n7580, n7581, n7582, n7583, n7584,
    n7585, n7586, n7587, n7588, n7589, n7590,
    n7591, n7592, n7593, n7594, n7595, n7596,
    n7597, n7598, n7599, n7600, n7601, n7602,
    n7604, n7605, n7606, n7607, n7608, n7609,
    n7610, n7611, n7612, n7613, n7614, n7615,
    n7616, n7617, n7618, n7619, n7620, n7621,
    n7622, n7623, n7624, n7625, n7626, n7627,
    n7628, n7629, n7630, n7631, n7632, n7633,
    n7634, n7635, n7636, n7637, n7638, n7639,
    n7640, n7641, n7642, n7643, n7644, n7645,
    n7646, n7647, n7648, n7649, n7650, n7651,
    n7652, n7653, n7654, n7655, n7656, n7657,
    n7658, n7659, n7660, n7661, n7662, n7663,
    n7664, n7665, n7666, n7667, n7668, n7669,
    n7670, n7671, n7672, n7673, n7674, n7675,
    n7676, n7677, n7678, n7679, n7680, n7681,
    n7682, n7683, n7684, n7685, n7686, n7687,
    n7688, n7690, n7691, n7692, n7693, n7694,
    n7695, n7696, n7697, n7698, n7699, n7700,
    n7701, n7702, n7703, n7704, n7705, n7706,
    n7707, n7708, n7709, n7710, n7711, n7712,
    n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7722, n7723, n7724,
    n7725, n7726, n7727, n7728, n7729, n7730,
    n7731, n7732, n7733, n7734, n7735, n7736,
    n7737, n7738, n7739, n7740, n7741, n7742,
    n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754,
    n7755, n7756, n7757, n7758, n7759, n7760,
    n7761, n7762, n7763, n7764, n7765, n7766,
    n7767, n7768, n7769, n7770, n7771, n7772,
    n7773, n7774, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785,
    n7786, n7787, n7788, n7789, n7790, n7791,
    n7792, n7793, n7794, n7795, n7796, n7797,
    n7798, n7799, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821,
    n7822, n7823, n7824, n7825, n7826, n7827,
    n7828, n7829, n7830, n7831, n7832, n7833,
    n7834, n7835, n7836, n7837, n7838, n7839,
    n7840, n7841, n7842, n7843, n7844, n7845,
    n7846, n7847, n7848, n7849, n7850, n7851,
    n7852, n7853, n7854, n7855, n7856, n7857,
    n7858, n7859, n7860, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912,
    n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7948, n7949,
    n7950, n7951, n7952, n7953, n7954, n7955,
    n7956, n7957, n7958, n7959, n7960, n7961,
    n7962, n7963, n7964, n7965, n7966, n7967,
    n7968, n7969, n7970, n7971, n7972, n7973,
    n7974, n7975, n7976, n7977, n7978, n7979,
    n7980, n7981, n7982, n7983, n7984, n7985,
    n7986, n7987, n7988, n7989, n7990, n7991,
    n7992, n7993, n7994, n7995, n7996, n7997,
    n7998, n7999, n8000, n8001, n8002, n8003,
    n8004, n8005, n8006, n8007, n8008, n8009,
    n8010, n8011, n8012, n8013, n8014, n8015,
    n8016, n8017, n8018, n8019, n8020, n8021,
    n8022, n8023, n8024, n8025, n8026, n8027,
    n8028, n8029, n8030, n8031, n8032, n8034,
    n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046,
    n8047, n8048, n8049, n8050, n8051, n8052,
    n8053, n8054, n8055, n8056, n8057, n8058,
    n8059, n8060, n8061, n8062, n8063, n8064,
    n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076,
    n8077, n8078, n8079, n8080, n8081, n8082,
    n8083, n8084, n8085, n8086, n8087, n8088,
    n8089, n8090, n8091, n8092, n8093, n8094,
    n8095, n8096, n8097, n8098, n8099, n8100,
    n8101, n8102, n8103, n8104, n8105, n8106,
    n8107, n8108, n8109, n8110, n8111, n8112,
    n8113, n8114, n8115, n8116, n8117, n8118,
    n8120, n8121, n8122, n8123, n8124, n8125,
    n8126, n8127, n8128, n8129, n8130, n8131,
    n8132, n8133, n8134, n8135, n8136, n8137,
    n8138, n8139, n8140, n8141, n8142, n8143,
    n8144, n8145, n8146, n8147, n8148, n8149,
    n8150, n8151, n8152, n8153, n8154, n8155,
    n8156, n8157, n8158, n8159, n8160, n8161,
    n8162, n8163, n8164, n8165, n8166, n8167,
    n8168, n8169, n8170, n8171, n8172, n8173,
    n8174, n8175, n8176, n8177, n8178, n8179,
    n8180, n8181, n8182, n8183, n8184, n8185,
    n8186, n8187, n8188, n8189, n8190, n8191,
    n8192, n8193, n8194, n8195, n8196, n8197,
    n8198, n8199, n8200, n8201, n8202, n8203,
    n8204, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216,
    n8217, n8218, n8219, n8220, n8221, n8222,
    n8223, n8224, n8225, n8226, n8227, n8228,
    n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246,
    n8247, n8248, n8249, n8250, n8251, n8252,
    n8253, n8254, n8255, n8256, n8257, n8258,
    n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276,
    n8277, n8278, n8279, n8280, n8281, n8282,
    n8283, n8284, n8285, n8286, n8287, n8288,
    n8289, n8290, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301,
    n8302, n8303, n8304, n8305, n8306, n8307,
    n8308, n8309, n8310, n8311, n8312, n8313,
    n8314, n8315, n8316, n8317, n8318, n8319,
    n8320, n8321, n8322, n8323, n8324, n8325,
    n8326, n8327, n8328, n8329, n8330, n8331,
    n8332, n8333, n8334, n8335, n8336, n8337,
    n8338, n8339, n8340, n8341, n8342, n8343,
    n8344, n8345, n8346, n8347, n8348, n8349,
    n8350, n8351, n8352, n8353, n8354, n8355,
    n8356, n8357, n8358, n8359, n8360, n8361,
    n8362, n8363, n8364, n8365, n8366, n8367,
    n8368, n8369, n8370, n8371, n8372, n8373,
    n8374, n8375, n8376, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386,
    n8387, n8388, n8389, n8390, n8391, n8392,
    n8393, n8394, n8395, n8396, n8397, n8398,
    n8399, n8400, n8401, n8402, n8403, n8404,
    n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8414, n8415, n8416,
    n8417, n8418, n8419, n8420, n8421, n8422,
    n8423, n8424, n8425, n8426, n8427, n8428,
    n8429, n8430, n8431, n8432, n8433, n8434,
    n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446,
    n8447, n8448, n8449, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8464, n8465,
    n8466, n8467, n8468, n8469, n8470, n8471,
    n8472, n8473, n8474, n8475, n8476, n8477,
    n8478, n8479, n8480, n8481, n8482, n8483,
    n8484, n8485, n8486, n8487, n8488, n8489,
    n8490, n8491, n8492, n8493, n8494, n8495,
    n8496, n8497, n8498, n8499, n8500, n8501,
    n8502, n8503, n8504, n8505, n8506, n8507,
    n8508, n8509, n8510, n8511, n8512, n8513,
    n8514, n8515, n8516, n8517, n8518, n8519,
    n8520, n8521, n8522, n8523, n8524, n8525,
    n8526, n8527, n8528, n8529, n8530, n8531,
    n8532, n8533, n8534, n8535, n8536, n8537,
    n8538, n8539, n8540, n8541, n8542, n8543,
    n8544, n8545, n8546, n8547, n8548, n8550,
    n8551, n8552, n8553, n8554, n8555, n8556,
    n8557, n8558, n8559, n8560, n8561, n8562,
    n8563, n8564, n8565, n8566, n8567, n8568,
    n8569, n8570, n8571, n8572, n8573, n8574,
    n8575, n8576, n8577, n8578, n8579, n8580,
    n8581, n8582, n8583, n8584, n8585, n8586,
    n8587, n8588, n8589, n8590, n8591, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598,
    n8599, n8600, n8601, n8602, n8603, n8604,
    n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8613, n8614, n8615, n8616,
    n8617, n8618, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8631, n8632, n8633, n8634,
    n8636, n8637, n8638, n8639, n8640, n8641,
    n8642, n8643, n8644, n8645, n8646, n8647,
    n8648, n8649, n8650, n8651, n8652, n8653,
    n8654, n8655, n8656, n8657, n8658, n8659,
    n8660, n8661, n8662, n8663, n8664, n8665,
    n8666, n8667, n8668, n8669, n8670, n8671,
    n8672, n8673, n8674, n8675, n8676, n8677,
    n8678, n8679, n8680, n8681, n8682, n8683,
    n8684, n8685, n8686, n8687, n8688, n8689,
    n8690, n8691, n8692, n8693, n8694, n8695,
    n8696, n8697, n8698, n8699, n8700, n8701,
    n8702, n8703, n8704, n8705, n8706, n8707,
    n8708, n8709, n8710, n8711, n8712, n8713,
    n8714, n8715, n8716, n8717, n8718, n8719,
    n8720, n8722, n8723, n8724, n8725, n8726,
    n8727, n8728, n8729, n8730, n8731, n8732,
    n8733, n8734, n8735, n8736, n8737, n8738,
    n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756,
    n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768,
    n8769, n8770, n8771, n8772, n8773, n8774,
    n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786,
    n8787, n8788, n8789, n8790, n8791, n8792,
    n8793, n8794, n8795, n8796, n8797, n8798,
    n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8808, n8809, n8810, n8811,
    n8812, n8813, n8814, n8815, n8816, n8817,
    n8818, n8819, n8820, n8821, n8822, n8823,
    n8824, n8825, n8826, n8827, n8828, n8829,
    n8830, n8831, n8832, n8833, n8834, n8835,
    n8836, n8837, n8838, n8839, n8840, n8841,
    n8842, n8843, n8844, n8845, n8846, n8847,
    n8848, n8849, n8850, n8851, n8852, n8853,
    n8854, n8855, n8856, n8857, n8858, n8859,
    n8860, n8861, n8862, n8863, n8864, n8865,
    n8866, n8867, n8868, n8869, n8870, n8871,
    n8872, n8873, n8874, n8875, n8876, n8877,
    n8878, n8879, n8880, n8881, n8882, n8883,
    n8884, n8885, n8886, n8887, n8888, n8889,
    n8890, n8891, n8892, n8894, n8895, n8896,
    n8897, n8898, n8899, n8900, n8901, n8902,
    n8903, n8904, n8905, n8906, n8907, n8908,
    n8909, n8910, n8911, n8912, n8913, n8914,
    n8915, n8916, n8917, n8918, n8919, n8920,
    n8921, n8922, n8923, n8924, n8925, n8926,
    n8927, n8928, n8929, n8930, n8931, n8932,
    n8933, n8934, n8935, n8936, n8937, n8938,
    n8939, n8940, n8941, n8942, n8943, n8944,
    n8945, n8946, n8947, n8948, n8949, n8950,
    n8951, n8952, n8953, n8954, n8955, n8956,
    n8957, n8958, n8959, n8960, n8961, n8962,
    n8963, n8964, n8965, n8966, n8967, n8968,
    n8969, n8970, n8971, n8972, n8973, n8974,
    n8975, n8976, n8977, n8978, n8980, n8981,
    n8982, n8983, n8984, n8985, n8986, n8987,
    n8988, n8989, n8990, n8991, n8992, n8993,
    n8994, n8995, n8996, n8997, n8998, n8999,
    n9000, n9001, n9002, n9003, n9004, n9005,
    n9006, n9007, n9008, n9009, n9010, n9011,
    n9012, n9013, n9014, n9015, n9016, n9017,
    n9018, n9019, n9020, n9021, n9022, n9023,
    n9024, n9025, n9026, n9027, n9028, n9029,
    n9030, n9031, n9032, n9033, n9034, n9035,
    n9036, n9037, n9038, n9039, n9040, n9041,
    n9042, n9043, n9044, n9045, n9046, n9047,
    n9048, n9049, n9050, n9051, n9052, n9053,
    n9054, n9055, n9056, n9057, n9058, n9059,
    n9060, n9061, n9062, n9063, n9064, n9066,
    n9067, n9068, n9069, n9070, n9071, n9072,
    n9073, n9074, n9075, n9076, n9077, n9078,
    n9079, n9080, n9081, n9082, n9083, n9084,
    n9085, n9086, n9087, n9088, n9089, n9090,
    n9091, n9092, n9093, n9094, n9095, n9096,
    n9097, n9098, n9099, n9100, n9101, n9102,
    n9103, n9104, n9105, n9106, n9107, n9108,
    n9109, n9110, n9111, n9112, n9113, n9114,
    n9115, n9116, n9117, n9118, n9119, n9120,
    n9121, n9122, n9123, n9124, n9125, n9126,
    n9127, n9128, n9129, n9130, n9131, n9132,
    n9133, n9134, n9135, n9136, n9137, n9138,
    n9139, n9140, n9141, n9142, n9143, n9144,
    n9145, n9146, n9147, n9148, n9149, n9150,
    n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9238, n9239, n9240, n9241, n9242,
    n9243, n9244, n9245, n9246, n9247, n9248,
    n9249, n9250, n9251, n9252, n9253, n9254,
    n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9265, n9266,
    n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278,
    n9279, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296,
    n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9307, n9308,
    n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9324, n9325, n9326, n9327,
    n9328, n9329, n9330, n9331, n9332, n9333,
    n9334, n9335, n9336, n9337, n9338, n9339,
    n9340, n9341, n9342, n9343, n9344, n9345,
    n9346, n9347, n9348, n9349, n9350, n9351,
    n9352, n9353, n9354, n9355, n9356, n9357,
    n9358, n9359, n9360, n9361, n9362, n9363,
    n9364, n9365, n9366, n9367, n9368, n9369,
    n9370, n9371, n9372, n9373, n9374, n9375,
    n9376, n9377, n9378, n9379, n9380, n9381,
    n9382, n9383, n9384, n9385, n9386, n9387,
    n9388, n9389, n9390, n9391, n9392, n9393,
    n9394, n9395, n9396, n9397, n9398, n9399,
    n9400, n9401, n9402, n9403, n9404, n9405,
    n9406, n9407, n9408, n9410, n9411, n9412,
    n9413, n9414, n9415, n9416, n9417, n9418,
    n9419, n9420, n9421, n9422, n9423, n9424,
    n9425, n9426, n9427, n9428, n9429, n9430,
    n9431, n9432, n9433, n9434, n9435, n9436,
    n9437, n9438, n9439, n9440, n9441, n9442,
    n9443, n9444, n9445, n9446, n9447, n9448,
    n9449, n9450, n9451, n9452, n9453, n9454,
    n9455, n9456, n9457, n9458, n9459, n9460,
    n9461, n9462, n9463, n9464, n9465, n9466,
    n9467, n9468, n9469, n9470, n9471, n9472,
    n9473, n9474, n9475, n9476, n9477, n9478,
    n9479, n9480, n9481, n9482, n9483, n9484,
    n9485, n9486, n9487, n9488, n9489, n9490,
    n9491, n9492, n9493, n9494, n9496, n9497,
    n9498, n9499, n9500, n9501, n9502, n9503,
    n9504, n9505, n9506, n9507, n9508, n9509,
    n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521,
    n9522, n9523, n9524, n9525, n9526, n9527,
    n9528, n9529, n9530, n9531, n9532, n9533,
    n9534, n9535, n9536, n9537, n9538, n9539,
    n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9547, n9548, n9549, n9550, n9551,
    n9552, n9553, n9554, n9555, n9556, n9557,
    n9558, n9559, n9560, n9561, n9562, n9563,
    n9564, n9565, n9566, n9567, n9568, n9569,
    n9570, n9571, n9572, n9573, n9574, n9575,
    n9576, n9577, n9578, n9579, n9580, n9582,
    n9583, n9584, n9585, n9586, n9587, n9588,
    n9589, n9590, n9591, n9592, n9593, n9594,
    n9595, n9596, n9597, n9598, n9599, n9600,
    n9601, n9602, n9603, n9604, n9605, n9606,
    n9607, n9608, n9609, n9610, n9611, n9612,
    n9613, n9614, n9615, n9616, n9617, n9618,
    n9619, n9620, n9621, n9622, n9623, n9624,
    n9625, n9626, n9627, n9628, n9629, n9630,
    n9631, n9632, n9633, n9634, n9635, n9636,
    n9637, n9638, n9639, n9640, n9641, n9642,
    n9643, n9644, n9645, n9646, n9647, n9648,
    n9649, n9650, n9651, n9652, n9653, n9654,
    n9655, n9656, n9657, n9658, n9659, n9660,
    n9661, n9662, n9663, n9664, n9665, n9666,
    n9668, n9669, n9670, n9671, n9672, n9673,
    n9674, n9675, n9676, n9677, n9678, n9679,
    n9680, n9681, n9682, n9683, n9684, n9685,
    n9686, n9687, n9688, n9689, n9690, n9691,
    n9692, n9693, n9694, n9695, n9696, n9697,
    n9698, n9699, n9700, n9701, n9702, n9703,
    n9704, n9705, n9706, n9707, n9708, n9709,
    n9710, n9711, n9712, n9713, n9714, n9715,
    n9716, n9717, n9718, n9719, n9720, n9721,
    n9722, n9723, n9724, n9725, n9726, n9727,
    n9728, n9729, n9730, n9731, n9732, n9733,
    n9734, n9735, n9736, n9737, n9738, n9739,
    n9740, n9741, n9742, n9743, n9744, n9745,
    n9746, n9747, n9748, n9749, n9750, n9751,
    n9752, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9840, n9841, n9842, n9843,
    n9844, n9845, n9846, n9847, n9848, n9849,
    n9850, n9851, n9852, n9853, n9854, n9855,
    n9856, n9857, n9858, n9859, n9860, n9861,
    n9862, n9863, n9864, n9865, n9866, n9867,
    n9868, n9869, n9870, n9871, n9872, n9873,
    n9874, n9875, n9876, n9877, n9878, n9879,
    n9880, n9881, n9882, n9883, n9884, n9885,
    n9886, n9887, n9888, n9889, n9890, n9891,
    n9892, n9893, n9894, n9895, n9896, n9897,
    n9898, n9899, n9900, n9901, n9902, n9903,
    n9904, n9905, n9906, n9907, n9908, n9909,
    n9910, n9911, n9912, n9913, n9914, n9915,
    n9916, n9917, n9918, n9919, n9920, n9921,
    n9922, n9923, n9924, n9926, n9927, n9928,
    n9929, n9930, n9931, n9932, n9933, n9934,
    n9935, n9936, n9937, n9938, n9939, n9940,
    n9941, n9942, n9943, n9944, n9945, n9946,
    n9947, n9948, n9949, n9950, n9951, n9952,
    n9953, n9954, n9955, n9956, n9957, n9958,
    n9959, n9960, n9961, n9962, n9963, n9964,
    n9965, n9966, n9967, n9968, n9969, n9970,
    n9971, n9972, n9973, n9974, n9975, n9976,
    n9977, n9978, n9979, n9980, n9981, n9982,
    n9983, n9984, n9985, n9986, n9987, n9988,
    n9989, n9990, n9991, n9992, n9993, n9994,
    n9995, n9996, n9997, n9998, n9999, n10000,
    n10001, n10002, n10003, n10004, n10005, n10006,
    n10007, n10008, n10009, n10010, n10012, n10013,
    n10014, n10015, n10016, n10017, n10018, n10019,
    n10020, n10021, n10022, n10023, n10024, n10025,
    n10026, n10027, n10028, n10029, n10030, n10031,
    n10032, n10033, n10034, n10035, n10036, n10037,
    n10038, n10039, n10040, n10041, n10042, n10043,
    n10044, n10045, n10046, n10047, n10048, n10049,
    n10050, n10051, n10052, n10053, n10054, n10055,
    n10056, n10057, n10058, n10059, n10060, n10061,
    n10062, n10063, n10064, n10065, n10066, n10067,
    n10068, n10069, n10070, n10071, n10072, n10073,
    n10074, n10075, n10076, n10077, n10078, n10079,
    n10080, n10081, n10082, n10083, n10084, n10085,
    n10086, n10087, n10088, n10089, n10090, n10091,
    n10092, n10093, n10094, n10095, n10096, n10098,
    n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116,
    n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134,
    n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146,
    n10147, n10148, n10149, n10150, n10151, n10152,
    n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170,
    n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182,
    n10184, n10185, n10186, n10187, n10188, n10189,
    n10190, n10191, n10192, n10193, n10194, n10195,
    n10196, n10197, n10198, n10199, n10200, n10201,
    n10202, n10203, n10204, n10205, n10206, n10207,
    n10208, n10209, n10210, n10211, n10212, n10213,
    n10214, n10215, n10216, n10217, n10218, n10219,
    n10220, n10221, n10222, n10223, n10224, n10225,
    n10226, n10227, n10228, n10229, n10230, n10231,
    n10232, n10233, n10234, n10235, n10236, n10237,
    n10238, n10239, n10240, n10241, n10242, n10243,
    n10244, n10245, n10246, n10247, n10248, n10249,
    n10250, n10251, n10252, n10253, n10254, n10255,
    n10256, n10257, n10258, n10259, n10260, n10261,
    n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10270, n10271, n10272, n10273, n10274,
    n10275, n10276, n10277, n10278, n10279, n10280,
    n10281, n10282, n10283, n10284, n10285, n10286,
    n10287, n10288, n10289, n10290, n10291, n10292,
    n10293, n10294, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10303, n10304,
    n10305, n10306, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10315, n10316,
    n10317, n10318, n10319, n10320, n10321, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328,
    n10329, n10330, n10331, n10332, n10333, n10334,
    n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346,
    n10347, n10348, n10349, n10350, n10351, n10352,
    n10353, n10354, n10356, n10357, n10358, n10359,
    n10360, n10361, n10362, n10363, n10364, n10365,
    n10366, n10367, n10368, n10369, n10370, n10371,
    n10372, n10373, n10374, n10375, n10376, n10377,
    n10378, n10379, n10380, n10381, n10382, n10383,
    n10384, n10385, n10386, n10387, n10388, n10389,
    n10390, n10391, n10392, n10393, n10394, n10395,
    n10396, n10397, n10398, n10399, n10400, n10401,
    n10402, n10403, n10404, n10405, n10406, n10407,
    n10408, n10409, n10410, n10411, n10412, n10413,
    n10414, n10415, n10416, n10417, n10418, n10419,
    n10420, n10421, n10422, n10423, n10424, n10425,
    n10426, n10427, n10428, n10429, n10430, n10431,
    n10432, n10433, n10434, n10435, n10436, n10437,
    n10438, n10439, n10440, n10442, n10443, n10444,
    n10445, n10446, n10447, n10448, n10449, n10450,
    n10451, n10452, n10453, n10454, n10455, n10456,
    n10457, n10458, n10459, n10460, n10461, n10462,
    n10463, n10464, n10465, n10466, n10467, n10468,
    n10469, n10470, n10471, n10472, n10473, n10474,
    n10475, n10476, n10477, n10478, n10479, n10480,
    n10481, n10482, n10483, n10484, n10485, n10486,
    n10487, n10488, n10489, n10490, n10491, n10492,
    n10493, n10494, n10495, n10496, n10497, n10498,
    n10499, n10500, n10501, n10502, n10503, n10504,
    n10505, n10506, n10507, n10508, n10509, n10510,
    n10511, n10512, n10513, n10514, n10515, n10516,
    n10517, n10518, n10519, n10520, n10521, n10522,
    n10523, n10524, n10525, n10526, n10528, n10529,
    n10530, n10531, n10532, n10533, n10534, n10535,
    n10536, n10537, n10538, n10539, n10540, n10541,
    n10542, n10543, n10544, n10545, n10546, n10547,
    n10548, n10549, n10550, n10551, n10552, n10553,
    n10554, n10555, n10556, n10557, n10558, n10559,
    n10560, n10561, n10562, n10563, n10564, n10565,
    n10566, n10567, n10568, n10569, n10570, n10571,
    n10572, n10573, n10574, n10575, n10576, n10577,
    n10578, n10579, n10580, n10581, n10582, n10583,
    n10584, n10585, n10586, n10587, n10588, n10589,
    n10590, n10591, n10592, n10593, n10594, n10595,
    n10596, n10597, n10598, n10599, n10600, n10601,
    n10602, n10603, n10604, n10605, n10606, n10607,
    n10608, n10609, n10610, n10611, n10612, n10614,
    n10615, n10616, n10617, n10618, n10619, n10620,
    n10621, n10622, n10623, n10624, n10625, n10626,
    n10627, n10628, n10629, n10630, n10631, n10632,
    n10633, n10634, n10635, n10636, n10637, n10638,
    n10639, n10640, n10641, n10642, n10643, n10644,
    n10645, n10646, n10647, n10648, n10649, n10650,
    n10651, n10652, n10653, n10654, n10655, n10656,
    n10657, n10658, n10659, n10660, n10661, n10662,
    n10663, n10664, n10665, n10666, n10667, n10668,
    n10669, n10670, n10671, n10672, n10673, n10674,
    n10675, n10676, n10677, n10678, n10679, n10680,
    n10681, n10682, n10683, n10684, n10685, n10686,
    n10687, n10688, n10689, n10690, n10691, n10692,
    n10693, n10694, n10695, n10696, n10697, n10698,
    n10700, n10701, n10702, n10703, n10704, n10705,
    n10706, n10707, n10708, n10709, n10710, n10711,
    n10712, n10713, n10714, n10715, n10716, n10717,
    n10718, n10719, n10720, n10721, n10722, n10723,
    n10724, n10725, n10726, n10727, n10728, n10729,
    n10730, n10731, n10732, n10733, n10734, n10735,
    n10736, n10737, n10738, n10739, n10740, n10741,
    n10742, n10743, n10744, n10745, n10746, n10747,
    n10748, n10749, n10750, n10751, n10752, n10753,
    n10754, n10755, n10756, n10757, n10758, n10759,
    n10760, n10761, n10762, n10763, n10764, n10765,
    n10766, n10767, n10768, n10769, n10770, n10771,
    n10772, n10773, n10774, n10775, n10776, n10777,
    n10778, n10779, n10780, n10781, n10782, n10783,
    n10784, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838,
    n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850,
    n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868,
    n10869, n10870, n10872, n10873, n10874, n10875,
    n10876, n10877, n10878, n10879, n10880, n10881,
    n10882, n10883, n10884, n10885, n10886, n10887,
    n10888, n10889, n10890, n10891, n10892, n10893,
    n10894, n10895, n10896, n10897, n10898, n10899,
    n10900, n10901, n10902, n10903, n10904, n10905,
    n10906, n10907, n10908, n10909, n10910, n10911,
    n10912, n10913, n10914, n10915, n10916, n10917,
    n10918, n10919, n10920, n10921, n10922, n10923,
    n10924, n10925, n10926, n10927, n10928, n10929,
    n10930, n10931, n10932, n10933, n10934, n10935,
    n10936, n10937, n10938, n10939, n10940, n10941,
    n10942, n10943, n10944, n10945, n10946, n10947,
    n10948, n10949, n10950, n10951, n10952, n10953,
    n10954, n10955, n10956, n10958, n10959, n10960,
    n10961, n10962, n10963, n10964, n10965, n10966,
    n10967, n10968, n10969, n10970, n10971, n10972,
    n10973, n10974, n10975, n10976, n10977, n10978,
    n10979, n10980, n10981, n10982, n10983, n10984,
    n10985, n10986, n10987, n10988, n10989, n10990,
    n10991, n10992, n10993, n10994, n10995, n10996,
    n10997, n10998, n10999, n11000, n11001, n11002,
    n11003, n11004, n11005, n11006, n11007, n11008,
    n11009, n11010, n11011, n11012, n11013, n11014,
    n11015, n11016, n11017, n11018, n11019, n11020,
    n11021, n11022, n11023, n11024, n11025, n11026,
    n11027, n11028, n11029, n11030, n11031, n11032,
    n11033, n11034, n11035, n11036, n11037, n11038,
    n11039, n11040, n11041, n11042, n11044, n11045,
    n11046, n11047, n11048, n11049, n11050, n11051,
    n11052, n11053, n11054, n11055, n11056, n11057,
    n11058, n11059, n11060, n11061, n11062, n11063,
    n11064, n11065, n11066, n11067, n11068, n11069,
    n11070, n11071, n11072, n11073, n11074, n11075,
    n11076, n11077, n11078, n11079, n11080, n11081,
    n11082, n11083, n11084, n11085, n11086, n11087,
    n11088, n11089, n11090, n11091, n11092, n11093,
    n11094, n11095, n11096, n11097, n11098, n11099,
    n11100, n11101, n11102, n11103, n11104, n11105,
    n11106, n11107, n11108, n11109, n11110, n11111,
    n11112, n11113, n11114, n11115, n11116, n11117,
    n11118, n11119, n11120, n11121, n11122, n11123,
    n11124, n11125, n11126, n11127, n11128, n11130,
    n11131, n11132, n11133, n11134, n11135, n11136,
    n11137, n11138, n11139, n11140, n11141, n11142,
    n11143, n11144, n11145, n11146, n11147, n11148,
    n11149, n11150, n11151, n11152, n11153, n11154,
    n11155, n11156, n11157, n11158, n11159, n11160,
    n11161, n11162, n11163, n11164, n11165, n11166,
    n11167, n11168, n11169, n11170, n11171, n11172,
    n11173, n11174, n11175, n11176, n11177, n11178,
    n11179, n11180, n11181, n11182, n11183, n11184,
    n11185, n11186, n11187, n11188, n11189, n11190,
    n11191, n11192, n11193, n11194, n11195, n11196,
    n11197, n11198, n11199, n11200, n11201, n11202,
    n11203, n11204, n11205, n11206, n11207, n11208,
    n11209, n11210, n11211, n11212, n11213, n11214,
    n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227,
    n11228, n11229, n11230, n11231, n11232, n11233,
    n11234, n11235, n11236, n11237, n11238, n11239,
    n11240, n11241, n11242, n11243, n11244, n11245,
    n11246, n11247, n11248, n11249, n11250, n11251,
    n11252, n11253, n11254, n11255, n11256, n11257,
    n11258, n11259, n11260, n11261, n11262, n11263,
    n11264, n11265, n11266, n11267, n11268, n11269,
    n11270, n11271, n11272, n11273, n11274, n11275,
    n11276, n11277, n11278, n11279, n11280, n11281,
    n11282, n11283, n11284, n11285, n11286, n11287,
    n11288, n11289, n11290, n11291, n11292, n11293,
    n11294, n11295, n11296, n11297, n11298, n11299,
    n11300, n11302, n11303, n11304, n11305, n11306,
    n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318,
    n11319, n11320, n11321, n11322, n11323, n11324,
    n11325, n11326, n11327, n11328, n11329, n11330,
    n11331, n11332, n11333, n11334, n11335, n11336,
    n11337, n11338, n11339, n11340, n11341, n11342,
    n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11350, n11351, n11352, n11353, n11354,
    n11355, n11356, n11357, n11358, n11359, n11360,
    n11361, n11362, n11363, n11364, n11365, n11366,
    n11367, n11368, n11369, n11370, n11371, n11372,
    n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11386, n11388, n11389, n11390, n11391,
    n11392, n11393, n11394, n11395, n11396, n11397,
    n11398, n11399, n11400, n11401, n11402, n11403,
    n11404, n11405, n11406, n11407, n11408, n11409,
    n11410, n11411, n11412, n11413, n11414, n11415,
    n11416, n11417, n11418, n11419, n11420, n11421,
    n11422, n11423, n11424, n11425, n11426, n11427,
    n11428, n11429, n11430, n11431, n11432, n11433,
    n11434, n11435, n11436, n11437, n11438, n11439,
    n11440, n11441, n11442, n11443, n11444, n11445,
    n11446, n11447, n11448, n11449, n11450, n11451,
    n11452, n11453, n11454, n11455, n11456, n11457,
    n11458, n11459, n11460, n11461, n11462, n11463,
    n11464, n11465, n11466, n11467, n11468, n11469,
    n11470, n11471, n11472, n11474, n11475, n11476,
    n11477, n11478, n11479, n11480, n11481, n11482,
    n11483, n11484, n11485, n11486, n11487, n11488,
    n11489, n11490, n11491, n11492, n11493, n11494,
    n11495, n11496, n11497, n11498, n11499, n11500,
    n11501, n11502, n11503, n11504, n11505, n11506,
    n11507, n11508, n11509, n11510, n11511, n11512,
    n11513, n11514, n11515, n11516, n11517, n11518,
    n11519, n11520, n11521, n11522, n11523, n11524,
    n11525, n11526, n11527, n11528, n11529, n11530,
    n11531, n11532, n11533, n11534, n11535, n11536,
    n11537, n11538, n11539, n11540, n11541, n11542,
    n11543, n11544, n11545, n11546, n11547, n11548,
    n11549, n11550, n11551, n11552, n11553, n11554,
    n11555, n11556, n11557, n11558, n11560, n11561,
    n11562, n11563, n11564, n11565, n11566, n11567,
    n11568, n11569, n11570, n11571, n11572, n11573,
    n11574, n11575, n11576, n11577, n11578, n11579,
    n11580, n11581, n11582, n11583, n11584, n11585,
    n11586, n11587, n11588, n11589, n11590, n11591,
    n11592, n11593, n11594, n11595, n11596, n11597,
    n11598, n11599, n11600, n11601, n11602, n11603,
    n11604, n11605, n11606, n11607, n11608, n11609,
    n11610, n11611, n11612, n11613, n11614, n11615,
    n11616, n11617, n11618, n11619, n11620, n11621,
    n11622, n11623, n11624, n11625, n11626, n11627,
    n11628, n11629, n11630, n11631, n11632, n11633,
    n11634, n11635, n11636, n11637, n11638, n11639,
    n11640, n11641, n11642, n11643, n11644, n11646,
    n11647, n11648, n11649, n11650, n11651, n11652,
    n11653, n11654, n11655, n11656, n11657, n11658,
    n11659, n11660, n11661, n11662, n11663, n11664,
    n11665, n11666, n11667, n11668, n11669, n11670,
    n11671, n11672, n11673, n11674, n11675, n11676,
    n11677, n11678, n11679, n11680, n11681, n11682,
    n11683, n11684, n11685, n11686, n11687, n11688,
    n11689, n11690, n11691, n11692, n11693, n11694,
    n11695, n11696, n11697, n11698, n11699, n11700,
    n11701, n11702, n11703, n11704, n11705, n11706,
    n11707, n11708, n11709, n11710, n11711, n11712,
    n11713, n11714, n11715, n11716, n11717, n11718,
    n11719, n11720, n11721, n11722, n11723, n11724,
    n11725, n11726, n11727, n11728, n11729, n11730,
    n11732, n11733, n11734, n11735, n11736, n11737,
    n11738, n11739, n11740, n11741, n11742, n11743,
    n11744, n11745, n11746, n11747, n11748, n11749,
    n11750, n11751, n11752, n11753, n11754, n11755,
    n11756, n11757, n11758, n11759, n11760, n11761,
    n11762, n11763, n11764, n11765, n11766, n11767,
    n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779,
    n11780, n11781, n11782, n11783, n11784, n11785,
    n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797,
    n11798, n11799, n11800, n11801, n11802, n11803,
    n11804, n11805, n11806, n11807, n11808, n11809,
    n11810, n11811, n11812, n11813, n11814, n11815,
    n11816, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834,
    n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846,
    n11847, n11848, n11849, n11850, n11851, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11904, n11905, n11906, n11907,
    n11908, n11909, n11910, n11911, n11912, n11913,
    n11914, n11915, n11916, n11917, n11918, n11919,
    n11920, n11921, n11922, n11923, n11924, n11925,
    n11926, n11927, n11928, n11929, n11930, n11931,
    n11932, n11933, n11934, n11935, n11936, n11937,
    n11938, n11939, n11940, n11941, n11942, n11943,
    n11944, n11945, n11946, n11947, n11948, n11949,
    n11950, n11951, n11952, n11953, n11954, n11955,
    n11956, n11957, n11958, n11959, n11960, n11961,
    n11962, n11963, n11964, n11965, n11966, n11967,
    n11968, n11969, n11970, n11971, n11972, n11973,
    n11974, n11975, n11976, n11977, n11978, n11979,
    n11980, n11981, n11982, n11983, n11984, n11985,
    n11986, n11987, n11988, n11990, n11991, n11992,
    n11993, n11994, n11995, n11996, n11997, n11998,
    n11999, n12000, n12001, n12002, n12003, n12004,
    n12005, n12006, n12007, n12008, n12009, n12010,
    n12011, n12012, n12013, n12014, n12015, n12016,
    n12017, n12018, n12019, n12020, n12021, n12022,
    n12023, n12024, n12025, n12026, n12027, n12028,
    n12029, n12030, n12031, n12032, n12033, n12034,
    n12035, n12036, n12037, n12038, n12039, n12040,
    n12041, n12042, n12043, n12044, n12045, n12046,
    n12047, n12048, n12049, n12050, n12051, n12052,
    n12053, n12054, n12055, n12056, n12057, n12058,
    n12059, n12060, n12061, n12062, n12063, n12064,
    n12065, n12066, n12067, n12068, n12069, n12070,
    n12071, n12072, n12073, n12074, n12076, n12077,
    n12078, n12079, n12080, n12081, n12082, n12083,
    n12084, n12085, n12086, n12087, n12088, n12089,
    n12090, n12091, n12092, n12093, n12094, n12095,
    n12096, n12097, n12098, n12099, n12100, n12101,
    n12102, n12103, n12104, n12105, n12106, n12107,
    n12108, n12109, n12110, n12111, n12112, n12113,
    n12114, n12115, n12116, n12117, n12118, n12119,
    n12120, n12121, n12122, n12123, n12124, n12125,
    n12126, n12127, n12128, n12129, n12130, n12131,
    n12132, n12133, n12134, n12135, n12136, n12137,
    n12138, n12139, n12140, n12141, n12142, n12143,
    n12144, n12145, n12146, n12147, n12148, n12149,
    n12150, n12151, n12152, n12153, n12154, n12155,
    n12156, n12157, n12158, n12159, n12160, n12162,
    n12163, n12164, n12165, n12166, n12167, n12168,
    n12169, n12170, n12171, n12172, n12173, n12174,
    n12175, n12176, n12177, n12178, n12179, n12180,
    n12181, n12182, n12183, n12184, n12185, n12186,
    n12187, n12188, n12189, n12190, n12191, n12192,
    n12193, n12194, n12195, n12196, n12197, n12198,
    n12199, n12200, n12201, n12202, n12203, n12204,
    n12205, n12206, n12207, n12208, n12209, n12210,
    n12211, n12212, n12213, n12214, n12215, n12216,
    n12217, n12218, n12219, n12220, n12221, n12222,
    n12223;
  assign n386 = pi1  & ~pi129 ;
  assign n387 = ~pi2  & ~n386;
  assign n388 = ~pi130  & ~pi131 ;
  assign n389 = ~n387 & n388;
  assign n390 = pi3  & ~pi131 ;
  assign n391 = ~pi4  & ~n390;
  assign n392 = ~pi5  & n391;
  assign n393 = ~n389 & n392;
  assign n394 = ~pi5  & pi132 ;
  assign n395 = ~pi133  & ~pi134 ;
  assign n396 = ~n394 & n395;
  assign n397 = ~n393 & n396;
  assign n398 = pi6  & ~pi134 ;
  assign n399 = ~pi7  & ~n398;
  assign n400 = ~pi8  & n399;
  assign n401 = ~n397 & n400;
  assign n402 = ~pi8  & pi135 ;
  assign n403 = ~pi136  & ~pi137 ;
  assign n404 = ~n402 & n403;
  assign n405 = ~n401 & n404;
  assign n406 = pi9  & ~pi137 ;
  assign n407 = ~pi10  & ~n406;
  assign n408 = ~pi11  & n407;
  assign n409 = ~n405 & n408;
  assign n410 = ~pi11  & pi138 ;
  assign n411 = ~pi139  & ~pi140 ;
  assign n412 = ~n410 & n411;
  assign n413 = ~n409 & n412;
  assign n414 = pi12  & ~pi140 ;
  assign n415 = ~pi13  & ~n414;
  assign n416 = ~pi14  & n415;
  assign n417 = ~n413 & n416;
  assign n418 = ~pi14  & pi141 ;
  assign n419 = ~pi142  & ~pi143 ;
  assign n420 = ~n418 & n419;
  assign n421 = ~n417 & n420;
  assign n422 = pi15  & ~pi143 ;
  assign n423 = ~pi16  & ~n422;
  assign n424 = ~pi17  & n423;
  assign n425 = ~n421 & n424;
  assign n426 = ~pi17  & pi144 ;
  assign n427 = ~pi145  & ~pi146 ;
  assign n428 = ~n426 & n427;
  assign n429 = ~n425 & n428;
  assign n430 = pi18  & ~pi146 ;
  assign n431 = ~pi19  & ~n430;
  assign n432 = ~pi20  & n431;
  assign n433 = ~n429 & n432;
  assign n434 = ~pi20  & pi147 ;
  assign n435 = ~pi148  & ~pi149 ;
  assign n436 = ~n434 & n435;
  assign n437 = ~n433 & n436;
  assign n438 = pi21  & ~pi149 ;
  assign n439 = ~pi22  & ~n438;
  assign n440 = ~pi23  & n439;
  assign n441 = ~n437 & n440;
  assign n442 = ~pi23  & pi150 ;
  assign n443 = ~pi151  & ~pi152 ;
  assign n444 = ~n442 & n443;
  assign n445 = ~n441 & n444;
  assign n446 = pi24  & ~pi152 ;
  assign n447 = ~pi25  & ~n446;
  assign n448 = ~pi26  & n447;
  assign n449 = ~n445 & n448;
  assign n450 = ~pi26  & pi153 ;
  assign n451 = ~pi154  & ~pi155 ;
  assign n452 = ~n450 & n451;
  assign n453 = ~n449 & n452;
  assign n454 = pi27  & ~pi155 ;
  assign n455 = ~pi28  & ~n454;
  assign n456 = ~pi29  & n455;
  assign n457 = ~n453 & n456;
  assign n458 = ~pi29  & pi156 ;
  assign n459 = ~pi157  & ~pi158 ;
  assign n460 = ~n458 & n459;
  assign n461 = ~n457 & n460;
  assign n462 = pi30  & ~pi158 ;
  assign n463 = ~pi31  & ~n462;
  assign n464 = ~pi32  & n463;
  assign n465 = ~n461 & n464;
  assign n466 = ~pi32  & pi159 ;
  assign n467 = ~pi160  & ~pi161 ;
  assign n468 = ~n466 & n467;
  assign n469 = ~n465 & n468;
  assign n470 = pi33  & ~pi161 ;
  assign n471 = ~pi34  & ~n470;
  assign n472 = ~pi35  & n471;
  assign n473 = ~n469 & n472;
  assign n474 = ~pi35  & pi162 ;
  assign n475 = ~pi163  & ~pi164 ;
  assign n476 = ~n474 & n475;
  assign n477 = ~n473 & n476;
  assign n478 = pi36  & ~pi164 ;
  assign n479 = ~pi37  & ~n478;
  assign n480 = ~pi38  & n479;
  assign n481 = ~n477 & n480;
  assign n482 = ~pi38  & pi165 ;
  assign n483 = ~pi166  & ~pi167 ;
  assign n484 = ~n482 & n483;
  assign n485 = ~n481 & n484;
  assign n486 = pi39  & ~pi167 ;
  assign n487 = ~pi40  & ~n486;
  assign n488 = ~pi41  & n487;
  assign n489 = ~n485 & n488;
  assign n490 = ~pi41  & pi168 ;
  assign n491 = ~pi169  & ~pi170 ;
  assign n492 = ~n490 & n491;
  assign n493 = ~n489 & n492;
  assign n494 = pi42  & ~pi170 ;
  assign n495 = ~pi43  & ~n494;
  assign n496 = ~pi44  & n495;
  assign n497 = ~n493 & n496;
  assign n498 = ~pi44  & pi171 ;
  assign n499 = ~pi172  & ~pi173 ;
  assign n500 = ~n498 & n499;
  assign n501 = ~n497 & n500;
  assign n502 = pi45  & ~pi173 ;
  assign n503 = ~pi46  & ~n502;
  assign n504 = ~pi47  & n503;
  assign n505 = ~n501 & n504;
  assign n506 = ~pi47  & pi174 ;
  assign n507 = ~pi175  & ~pi176 ;
  assign n508 = ~n506 & n507;
  assign n509 = ~n505 & n508;
  assign n510 = pi48  & ~pi176 ;
  assign n511 = ~pi49  & ~n510;
  assign n512 = ~pi50  & n511;
  assign n513 = ~n509 & n512;
  assign n514 = ~pi50  & pi177 ;
  assign n515 = ~pi178  & ~pi179 ;
  assign n516 = ~n514 & n515;
  assign n517 = ~n513 & n516;
  assign n518 = pi51  & ~pi179 ;
  assign n519 = ~pi52  & ~n518;
  assign n520 = ~pi53  & n519;
  assign n521 = ~n517 & n520;
  assign n522 = ~pi53  & pi180 ;
  assign n523 = ~pi181  & ~pi182 ;
  assign n524 = ~n522 & n523;
  assign n525 = ~n521 & n524;
  assign n526 = pi54  & ~pi182 ;
  assign n527 = ~pi55  & ~n526;
  assign n528 = ~pi56  & n527;
  assign n529 = ~n525 & n528;
  assign n530 = ~pi56  & pi183 ;
  assign n531 = ~pi184  & ~pi185 ;
  assign n532 = ~n530 & n531;
  assign n533 = ~n529 & n532;
  assign n534 = pi57  & ~pi185 ;
  assign n535 = ~pi58  & ~n534;
  assign n536 = ~pi59  & n535;
  assign n537 = ~n533 & n536;
  assign n538 = ~pi59  & pi186 ;
  assign n539 = ~pi187  & ~pi188 ;
  assign n540 = ~n538 & n539;
  assign n541 = ~n537 & n540;
  assign n542 = pi60  & ~pi188 ;
  assign n543 = ~pi61  & ~n542;
  assign n544 = ~pi62  & n543;
  assign n545 = ~n541 & n544;
  assign n546 = ~pi62  & pi189 ;
  assign n547 = ~pi190  & ~pi191 ;
  assign n548 = ~n546 & n547;
  assign n549 = ~n545 & n548;
  assign n550 = pi63  & ~pi191 ;
  assign n551 = ~pi64  & ~n550;
  assign n552 = ~pi65  & n551;
  assign n553 = ~n549 & n552;
  assign n554 = ~pi65  & pi192 ;
  assign n555 = ~pi193  & ~pi194 ;
  assign n556 = ~n554 & n555;
  assign n557 = ~n553 & n556;
  assign n558 = pi66  & ~pi194 ;
  assign n559 = ~pi67  & ~n558;
  assign n560 = ~pi68  & n559;
  assign n561 = ~n557 & n560;
  assign n562 = ~pi68  & pi195 ;
  assign n563 = ~pi196  & ~pi197 ;
  assign n564 = ~n562 & n563;
  assign n565 = ~n561 & n564;
  assign n566 = pi69  & ~pi197 ;
  assign n567 = ~pi70  & ~n566;
  assign n568 = ~pi71  & n567;
  assign n569 = ~n565 & n568;
  assign n570 = ~pi71  & pi198 ;
  assign n571 = ~pi199  & ~pi200 ;
  assign n572 = ~n570 & n571;
  assign n573 = ~n569 & n572;
  assign n574 = pi72  & ~pi200 ;
  assign n575 = ~pi73  & ~n574;
  assign n576 = ~pi74  & n575;
  assign n577 = ~n573 & n576;
  assign n578 = ~pi74  & pi201 ;
  assign n579 = ~pi202  & ~pi203 ;
  assign n580 = ~n578 & n579;
  assign n581 = ~n577 & n580;
  assign n582 = pi75  & ~pi203 ;
  assign n583 = ~pi76  & ~n582;
  assign n584 = ~pi77  & n583;
  assign n585 = ~n581 & n584;
  assign n586 = ~pi77  & pi204 ;
  assign n587 = ~pi205  & ~pi206 ;
  assign n588 = ~n586 & n587;
  assign n589 = ~n585 & n588;
  assign n590 = pi78  & ~pi206 ;
  assign n591 = ~pi79  & ~n590;
  assign n592 = ~pi80  & n591;
  assign n593 = ~n589 & n592;
  assign n594 = ~pi80  & pi207 ;
  assign n595 = ~pi208  & ~pi209 ;
  assign n596 = ~n594 & n595;
  assign n597 = ~n593 & n596;
  assign n598 = pi81  & ~pi209 ;
  assign n599 = ~pi82  & ~n598;
  assign n600 = ~pi83  & n599;
  assign n601 = ~n597 & n600;
  assign n602 = ~pi83  & pi210 ;
  assign n603 = ~pi211  & ~pi212 ;
  assign n604 = ~n602 & n603;
  assign n605 = ~n601 & n604;
  assign n606 = pi84  & ~pi212 ;
  assign n607 = ~pi85  & ~n606;
  assign n608 = ~pi86  & n607;
  assign n609 = ~n605 & n608;
  assign n610 = ~pi86  & pi213 ;
  assign n611 = ~pi214  & ~pi215 ;
  assign n612 = ~n610 & n611;
  assign n613 = ~n609 & n612;
  assign n614 = pi87  & ~pi215 ;
  assign n615 = ~pi88  & ~n614;
  assign n616 = ~pi89  & n615;
  assign n617 = ~n613 & n616;
  assign n618 = ~pi89  & pi216 ;
  assign n619 = ~pi217  & ~pi218 ;
  assign n620 = ~n618 & n619;
  assign n621 = ~n617 & n620;
  assign n622 = pi90  & ~pi218 ;
  assign n623 = ~pi91  & ~n622;
  assign n624 = ~pi92  & n623;
  assign n625 = ~n621 & n624;
  assign n626 = ~pi92  & pi219 ;
  assign n627 = ~pi220  & ~pi221 ;
  assign n628 = ~n626 & n627;
  assign n629 = ~n625 & n628;
  assign n630 = pi93  & ~pi221 ;
  assign n631 = ~pi94  & ~n630;
  assign n632 = ~pi95  & n631;
  assign n633 = ~n629 & n632;
  assign n634 = ~pi95  & pi222 ;
  assign n635 = ~pi223  & ~pi224 ;
  assign n636 = ~n634 & n635;
  assign n637 = ~n633 & n636;
  assign n638 = pi96  & ~pi224 ;
  assign n639 = ~pi97  & ~n638;
  assign n640 = ~pi98  & n639;
  assign n641 = ~n637 & n640;
  assign n642 = ~pi98  & pi225 ;
  assign n643 = ~pi226  & ~pi227 ;
  assign n644 = ~n642 & n643;
  assign n645 = ~n641 & n644;
  assign n646 = pi99  & ~pi227 ;
  assign n647 = ~pi100  & ~n646;
  assign n648 = ~pi101  & n647;
  assign n649 = ~n645 & n648;
  assign n650 = ~pi101  & pi228 ;
  assign n651 = ~pi229  & ~pi230 ;
  assign n652 = ~n650 & n651;
  assign n653 = ~n649 & n652;
  assign n654 = pi102  & ~pi230 ;
  assign n655 = ~pi103  & ~n654;
  assign n656 = ~pi104  & n655;
  assign n657 = ~n653 & n656;
  assign n658 = ~pi104  & pi231 ;
  assign n659 = ~pi232  & ~pi233 ;
  assign n660 = ~n658 & n659;
  assign n661 = ~n657 & n660;
  assign n662 = pi105  & ~pi233 ;
  assign n663 = ~pi106  & ~n662;
  assign n664 = ~pi107  & n663;
  assign n665 = ~n661 & n664;
  assign n666 = ~pi107  & pi234 ;
  assign n667 = ~pi235  & ~pi236 ;
  assign n668 = ~n666 & n667;
  assign n669 = ~n665 & n668;
  assign n670 = pi108  & ~pi236 ;
  assign n671 = ~pi109  & ~n670;
  assign n672 = ~pi110  & n671;
  assign n673 = ~n669 & n672;
  assign n674 = ~pi110  & pi237 ;
  assign n675 = ~pi238  & ~pi239 ;
  assign n676 = ~n674 & n675;
  assign n677 = ~n673 & n676;
  assign n678 = pi111  & ~pi239 ;
  assign n679 = ~pi112  & ~n678;
  assign n680 = ~pi113  & n679;
  assign n681 = ~n677 & n680;
  assign n682 = ~pi113  & pi240 ;
  assign n683 = ~pi241  & ~pi242 ;
  assign n684 = ~n682 & n683;
  assign n685 = ~n681 & n684;
  assign n686 = pi114  & ~pi242 ;
  assign n687 = ~pi115  & ~n686;
  assign n688 = ~pi116  & n687;
  assign n689 = ~n685 & n688;
  assign n690 = ~pi116  & pi243 ;
  assign n691 = ~pi244  & ~pi245 ;
  assign n692 = ~n690 & n691;
  assign n693 = ~n689 & n692;
  assign n694 = pi117  & ~pi245 ;
  assign n695 = ~pi118  & ~n694;
  assign n696 = ~pi119  & n695;
  assign n697 = ~n693 & n696;
  assign n698 = ~pi119  & pi246 ;
  assign n699 = ~pi247  & ~pi248 ;
  assign n700 = ~n698 & n699;
  assign n701 = ~n697 & n700;
  assign n702 = pi120  & ~pi248 ;
  assign n703 = ~pi121  & ~n702;
  assign n704 = ~pi122  & n703;
  assign n705 = ~n701 & n704;
  assign n706 = ~pi122  & pi249 ;
  assign n707 = ~pi250  & ~pi251 ;
  assign n708 = ~n706 & n707;
  assign n709 = ~n705 & n708;
  assign n710 = pi123  & ~pi251 ;
  assign n711 = ~pi124  & ~n710;
  assign n712 = ~pi125  & n711;
  assign n713 = ~n709 & n712;
  assign n714 = ~pi125  & pi252 ;
  assign n715 = ~pi253  & ~pi254 ;
  assign n716 = ~n714 & n715;
  assign n717 = ~n713 & n716;
  assign n718 = pi126  & ~pi254 ;
  assign n719 = ~pi127  & ~n718;
  assign n720 = ~pi0  & n719;
  assign n721 = ~n717 & n720;
  assign n722 = ~pi0  & pi255 ;
  assign n723 = pi128  & ~n722;
  assign po0  = ~n721 & n723;
  assign n725 = pi2  & ~pi130 ;
  assign n726 = ~pi3  & ~n725;
  assign n727 = ~pi131  & ~pi132 ;
  assign n728 = ~n726 & n727;
  assign n729 = pi4  & ~pi132 ;
  assign n730 = ~pi5  & ~n729;
  assign n731 = ~pi6  & n730;
  assign n732 = ~n728 & n731;
  assign n733 = ~pi6  & pi133 ;
  assign n734 = ~pi134  & ~pi135 ;
  assign n735 = ~n733 & n734;
  assign n736 = ~n732 & n735;
  assign n737 = pi7  & ~pi135 ;
  assign n738 = ~pi8  & ~n737;
  assign n739 = ~pi9  & n738;
  assign n740 = ~n736 & n739;
  assign n741 = ~pi9  & pi136 ;
  assign n742 = ~pi137  & ~pi138 ;
  assign n743 = ~n741 & n742;
  assign n744 = ~n740 & n743;
  assign n745 = pi10  & ~pi138 ;
  assign n746 = ~pi11  & ~n745;
  assign n747 = ~pi12  & n746;
  assign n748 = ~n744 & n747;
  assign n749 = ~pi12  & pi139 ;
  assign n750 = ~pi140  & ~pi141 ;
  assign n751 = ~n749 & n750;
  assign n752 = ~n748 & n751;
  assign n753 = pi13  & ~pi141 ;
  assign n754 = ~pi14  & ~n753;
  assign n755 = ~pi15  & n754;
  assign n756 = ~n752 & n755;
  assign n757 = ~pi15  & pi142 ;
  assign n758 = ~pi143  & ~pi144 ;
  assign n759 = ~n757 & n758;
  assign n760 = ~n756 & n759;
  assign n761 = pi16  & ~pi144 ;
  assign n762 = ~pi17  & ~n761;
  assign n763 = ~pi18  & n762;
  assign n764 = ~n760 & n763;
  assign n765 = ~pi18  & pi145 ;
  assign n766 = ~pi146  & ~pi147 ;
  assign n767 = ~n765 & n766;
  assign n768 = ~n764 & n767;
  assign n769 = pi19  & ~pi147 ;
  assign n770 = ~pi20  & ~n769;
  assign n771 = ~pi21  & n770;
  assign n772 = ~n768 & n771;
  assign n773 = ~pi21  & pi148 ;
  assign n774 = ~pi149  & ~pi150 ;
  assign n775 = ~n773 & n774;
  assign n776 = ~n772 & n775;
  assign n777 = pi22  & ~pi150 ;
  assign n778 = ~pi23  & ~n777;
  assign n779 = ~pi24  & n778;
  assign n780 = ~n776 & n779;
  assign n781 = ~pi24  & pi151 ;
  assign n782 = ~pi152  & ~pi153 ;
  assign n783 = ~n781 & n782;
  assign n784 = ~n780 & n783;
  assign n785 = pi25  & ~pi153 ;
  assign n786 = ~pi26  & ~n785;
  assign n787 = ~pi27  & n786;
  assign n788 = ~n784 & n787;
  assign n789 = ~pi27  & pi154 ;
  assign n790 = ~pi155  & ~pi156 ;
  assign n791 = ~n789 & n790;
  assign n792 = ~n788 & n791;
  assign n793 = pi28  & ~pi156 ;
  assign n794 = ~pi29  & ~n793;
  assign n795 = ~pi30  & n794;
  assign n796 = ~n792 & n795;
  assign n797 = ~pi30  & pi157 ;
  assign n798 = ~pi158  & ~pi159 ;
  assign n799 = ~n797 & n798;
  assign n800 = ~n796 & n799;
  assign n801 = pi31  & ~pi159 ;
  assign n802 = ~pi32  & ~n801;
  assign n803 = ~pi33  & n802;
  assign n804 = ~n800 & n803;
  assign n805 = ~pi33  & pi160 ;
  assign n806 = ~pi161  & ~pi162 ;
  assign n807 = ~n805 & n806;
  assign n808 = ~n804 & n807;
  assign n809 = pi34  & ~pi162 ;
  assign n810 = ~pi35  & ~n809;
  assign n811 = ~pi36  & n810;
  assign n812 = ~n808 & n811;
  assign n813 = ~pi36  & pi163 ;
  assign n814 = ~pi164  & ~pi165 ;
  assign n815 = ~n813 & n814;
  assign n816 = ~n812 & n815;
  assign n817 = pi37  & ~pi165 ;
  assign n818 = ~pi38  & ~n817;
  assign n819 = ~pi39  & n818;
  assign n820 = ~n816 & n819;
  assign n821 = ~pi39  & pi166 ;
  assign n822 = ~pi167  & ~pi168 ;
  assign n823 = ~n821 & n822;
  assign n824 = ~n820 & n823;
  assign n825 = pi40  & ~pi168 ;
  assign n826 = ~pi41  & ~n825;
  assign n827 = ~pi42  & n826;
  assign n828 = ~n824 & n827;
  assign n829 = ~pi42  & pi169 ;
  assign n830 = ~pi170  & ~pi171 ;
  assign n831 = ~n829 & n830;
  assign n832 = ~n828 & n831;
  assign n833 = pi43  & ~pi171 ;
  assign n834 = ~pi44  & ~n833;
  assign n835 = ~pi45  & n834;
  assign n836 = ~n832 & n835;
  assign n837 = ~pi45  & pi172 ;
  assign n838 = ~pi173  & ~pi174 ;
  assign n839 = ~n837 & n838;
  assign n840 = ~n836 & n839;
  assign n841 = pi46  & ~pi174 ;
  assign n842 = ~pi47  & ~n841;
  assign n843 = ~pi48  & n842;
  assign n844 = ~n840 & n843;
  assign n845 = ~pi48  & pi175 ;
  assign n846 = ~pi176  & ~pi177 ;
  assign n847 = ~n845 & n846;
  assign n848 = ~n844 & n847;
  assign n849 = pi49  & ~pi177 ;
  assign n850 = ~pi50  & ~n849;
  assign n851 = ~pi51  & n850;
  assign n852 = ~n848 & n851;
  assign n853 = ~pi51  & pi178 ;
  assign n854 = ~pi179  & ~pi180 ;
  assign n855 = ~n853 & n854;
  assign n856 = ~n852 & n855;
  assign n857 = pi52  & ~pi180 ;
  assign n858 = ~pi53  & ~n857;
  assign n859 = ~pi54  & n858;
  assign n860 = ~n856 & n859;
  assign n861 = ~pi54  & pi181 ;
  assign n862 = ~pi182  & ~pi183 ;
  assign n863 = ~n861 & n862;
  assign n864 = ~n860 & n863;
  assign n865 = pi55  & ~pi183 ;
  assign n866 = ~pi56  & ~n865;
  assign n867 = ~pi57  & n866;
  assign n868 = ~n864 & n867;
  assign n869 = ~pi57  & pi184 ;
  assign n870 = ~pi185  & ~pi186 ;
  assign n871 = ~n869 & n870;
  assign n872 = ~n868 & n871;
  assign n873 = pi58  & ~pi186 ;
  assign n874 = ~pi59  & ~n873;
  assign n875 = ~pi60  & n874;
  assign n876 = ~n872 & n875;
  assign n877 = ~pi60  & pi187 ;
  assign n878 = ~pi188  & ~pi189 ;
  assign n879 = ~n877 & n878;
  assign n880 = ~n876 & n879;
  assign n881 = pi61  & ~pi189 ;
  assign n882 = ~pi62  & ~n881;
  assign n883 = ~pi63  & n882;
  assign n884 = ~n880 & n883;
  assign n885 = ~pi63  & pi190 ;
  assign n886 = ~pi191  & ~pi192 ;
  assign n887 = ~n885 & n886;
  assign n888 = ~n884 & n887;
  assign n889 = pi64  & ~pi192 ;
  assign n890 = ~pi65  & ~n889;
  assign n891 = ~pi66  & n890;
  assign n892 = ~n888 & n891;
  assign n893 = ~pi66  & pi193 ;
  assign n894 = ~pi194  & ~pi195 ;
  assign n895 = ~n893 & n894;
  assign n896 = ~n892 & n895;
  assign n897 = pi67  & ~pi195 ;
  assign n898 = ~pi68  & ~n897;
  assign n899 = ~pi69  & n898;
  assign n900 = ~n896 & n899;
  assign n901 = ~pi69  & pi196 ;
  assign n902 = ~pi197  & ~pi198 ;
  assign n903 = ~n901 & n902;
  assign n904 = ~n900 & n903;
  assign n905 = pi70  & ~pi198 ;
  assign n906 = ~pi71  & ~n905;
  assign n907 = ~pi72  & n906;
  assign n908 = ~n904 & n907;
  assign n909 = ~pi72  & pi199 ;
  assign n910 = ~pi200  & ~pi201 ;
  assign n911 = ~n909 & n910;
  assign n912 = ~n908 & n911;
  assign n913 = pi73  & ~pi201 ;
  assign n914 = ~pi74  & ~n913;
  assign n915 = ~pi75  & n914;
  assign n916 = ~n912 & n915;
  assign n917 = ~pi75  & pi202 ;
  assign n918 = ~pi203  & ~pi204 ;
  assign n919 = ~n917 & n918;
  assign n920 = ~n916 & n919;
  assign n921 = pi76  & ~pi204 ;
  assign n922 = ~pi77  & ~n921;
  assign n923 = ~pi78  & n922;
  assign n924 = ~n920 & n923;
  assign n925 = ~pi78  & pi205 ;
  assign n926 = ~pi206  & ~pi207 ;
  assign n927 = ~n925 & n926;
  assign n928 = ~n924 & n927;
  assign n929 = pi79  & ~pi207 ;
  assign n930 = ~pi80  & ~n929;
  assign n931 = ~pi81  & n930;
  assign n932 = ~n928 & n931;
  assign n933 = ~pi81  & pi208 ;
  assign n934 = ~pi209  & ~pi210 ;
  assign n935 = ~n933 & n934;
  assign n936 = ~n932 & n935;
  assign n937 = pi82  & ~pi210 ;
  assign n938 = ~pi83  & ~n937;
  assign n939 = ~pi84  & n938;
  assign n940 = ~n936 & n939;
  assign n941 = ~pi84  & pi211 ;
  assign n942 = ~pi212  & ~pi213 ;
  assign n943 = ~n941 & n942;
  assign n944 = ~n940 & n943;
  assign n945 = pi85  & ~pi213 ;
  assign n946 = ~pi86  & ~n945;
  assign n947 = ~pi87  & n946;
  assign n948 = ~n944 & n947;
  assign n949 = ~pi87  & pi214 ;
  assign n950 = ~pi215  & ~pi216 ;
  assign n951 = ~n949 & n950;
  assign n952 = ~n948 & n951;
  assign n953 = pi88  & ~pi216 ;
  assign n954 = ~pi89  & ~n953;
  assign n955 = ~pi90  & n954;
  assign n956 = ~n952 & n955;
  assign n957 = ~pi90  & pi217 ;
  assign n958 = ~pi218  & ~pi219 ;
  assign n959 = ~n957 & n958;
  assign n960 = ~n956 & n959;
  assign n961 = pi91  & ~pi219 ;
  assign n962 = ~pi92  & ~n961;
  assign n963 = ~pi93  & n962;
  assign n964 = ~n960 & n963;
  assign n965 = ~pi93  & pi220 ;
  assign n966 = ~pi221  & ~pi222 ;
  assign n967 = ~n965 & n966;
  assign n968 = ~n964 & n967;
  assign n969 = pi94  & ~pi222 ;
  assign n970 = ~pi95  & ~n969;
  assign n971 = ~pi96  & n970;
  assign n972 = ~n968 & n971;
  assign n973 = ~pi96  & pi223 ;
  assign n974 = ~pi224  & ~pi225 ;
  assign n975 = ~n973 & n974;
  assign n976 = ~n972 & n975;
  assign n977 = pi97  & ~pi225 ;
  assign n978 = ~pi98  & ~n977;
  assign n979 = ~pi99  & n978;
  assign n980 = ~n976 & n979;
  assign n981 = ~pi99  & pi226 ;
  assign n982 = ~pi227  & ~pi228 ;
  assign n983 = ~n981 & n982;
  assign n984 = ~n980 & n983;
  assign n985 = pi100  & ~pi228 ;
  assign n986 = ~pi101  & ~n985;
  assign n987 = ~pi102  & n986;
  assign n988 = ~n984 & n987;
  assign n989 = ~pi102  & pi229 ;
  assign n990 = ~pi230  & ~pi231 ;
  assign n991 = ~n989 & n990;
  assign n992 = ~n988 & n991;
  assign n993 = pi103  & ~pi231 ;
  assign n994 = ~pi104  & ~n993;
  assign n995 = ~pi105  & n994;
  assign n996 = ~n992 & n995;
  assign n997 = ~pi105  & pi232 ;
  assign n998 = ~pi233  & ~pi234 ;
  assign n999 = ~n997 & n998;
  assign n1000 = ~n996 & n999;
  assign n1001 = pi106  & ~pi234 ;
  assign n1002 = ~pi107  & ~n1001;
  assign n1003 = ~pi108  & n1002;
  assign n1004 = ~n1000 & n1003;
  assign n1005 = ~pi108  & pi235 ;
  assign n1006 = ~pi236  & ~pi237 ;
  assign n1007 = ~n1005 & n1006;
  assign n1008 = ~n1004 & n1007;
  assign n1009 = pi109  & ~pi237 ;
  assign n1010 = ~pi110  & ~n1009;
  assign n1011 = ~pi111  & n1010;
  assign n1012 = ~n1008 & n1011;
  assign n1013 = ~pi111  & pi238 ;
  assign n1014 = ~pi239  & ~pi240 ;
  assign n1015 = ~n1013 & n1014;
  assign n1016 = ~n1012 & n1015;
  assign n1017 = pi112  & ~pi240 ;
  assign n1018 = ~pi113  & ~n1017;
  assign n1019 = ~pi114  & n1018;
  assign n1020 = ~n1016 & n1019;
  assign n1021 = ~pi114  & pi241 ;
  assign n1022 = ~pi242  & ~pi243 ;
  assign n1023 = ~n1021 & n1022;
  assign n1024 = ~n1020 & n1023;
  assign n1025 = pi115  & ~pi243 ;
  assign n1026 = ~pi116  & ~n1025;
  assign n1027 = ~pi117  & n1026;
  assign n1028 = ~n1024 & n1027;
  assign n1029 = ~pi117  & pi244 ;
  assign n1030 = ~pi245  & ~pi246 ;
  assign n1031 = ~n1029 & n1030;
  assign n1032 = ~n1028 & n1031;
  assign n1033 = pi118  & ~pi246 ;
  assign n1034 = ~pi119  & ~n1033;
  assign n1035 = ~pi120  & n1034;
  assign n1036 = ~n1032 & n1035;
  assign n1037 = ~pi120  & pi247 ;
  assign n1038 = ~pi248  & ~pi249 ;
  assign n1039 = ~n1037 & n1038;
  assign n1040 = ~n1036 & n1039;
  assign n1041 = pi121  & ~pi249 ;
  assign n1042 = ~pi122  & ~n1041;
  assign n1043 = ~pi123  & n1042;
  assign n1044 = ~n1040 & n1043;
  assign n1045 = ~pi123  & pi250 ;
  assign n1046 = ~pi251  & ~pi252 ;
  assign n1047 = ~n1045 & n1046;
  assign n1048 = ~n1044 & n1047;
  assign n1049 = pi124  & ~pi252 ;
  assign n1050 = ~pi125  & ~n1049;
  assign n1051 = ~pi126  & n1050;
  assign n1052 = ~n1048 & n1051;
  assign n1053 = ~pi126  & pi253 ;
  assign n1054 = ~pi254  & ~pi255 ;
  assign n1055 = ~n1053 & n1054;
  assign n1056 = ~n1052 & n1055;
  assign n1057 = pi127  & ~pi255 ;
  assign n1058 = ~pi0  & ~n1057;
  assign n1059 = ~pi1  & n1058;
  assign n1060 = ~n1056 & n1059;
  assign n1061 = ~pi1  & pi128 ;
  assign n1062 = pi129  & ~n1061;
  assign po1  = ~n1060 & n1062;
  assign n1064 = ~pi132  & ~pi133 ;
  assign n1065 = ~n391 & n1064;
  assign n1066 = pi5  & ~pi133 ;
  assign n1067 = ~pi6  & ~n1066;
  assign n1068 = ~pi7  & n1067;
  assign n1069 = ~n1065 & n1068;
  assign n1070 = ~pi7  & pi134 ;
  assign n1071 = ~pi135  & ~pi136 ;
  assign n1072 = ~n1070 & n1071;
  assign n1073 = ~n1069 & n1072;
  assign n1074 = pi8  & ~pi136 ;
  assign n1075 = ~pi9  & ~n1074;
  assign n1076 = ~pi10  & n1075;
  assign n1077 = ~n1073 & n1076;
  assign n1078 = ~pi10  & pi137 ;
  assign n1079 = ~pi138  & ~pi139 ;
  assign n1080 = ~n1078 & n1079;
  assign n1081 = ~n1077 & n1080;
  assign n1082 = pi11  & ~pi139 ;
  assign n1083 = ~pi12  & ~n1082;
  assign n1084 = ~pi13  & n1083;
  assign n1085 = ~n1081 & n1084;
  assign n1086 = ~pi13  & pi140 ;
  assign n1087 = ~pi141  & ~pi142 ;
  assign n1088 = ~n1086 & n1087;
  assign n1089 = ~n1085 & n1088;
  assign n1090 = pi14  & ~pi142 ;
  assign n1091 = ~pi15  & ~n1090;
  assign n1092 = ~pi16  & n1091;
  assign n1093 = ~n1089 & n1092;
  assign n1094 = ~pi16  & pi143 ;
  assign n1095 = ~pi144  & ~pi145 ;
  assign n1096 = ~n1094 & n1095;
  assign n1097 = ~n1093 & n1096;
  assign n1098 = pi17  & ~pi145 ;
  assign n1099 = ~pi18  & ~n1098;
  assign n1100 = ~pi19  & n1099;
  assign n1101 = ~n1097 & n1100;
  assign n1102 = ~pi19  & pi146 ;
  assign n1103 = ~pi147  & ~pi148 ;
  assign n1104 = ~n1102 & n1103;
  assign n1105 = ~n1101 & n1104;
  assign n1106 = pi20  & ~pi148 ;
  assign n1107 = ~pi21  & ~n1106;
  assign n1108 = ~pi22  & n1107;
  assign n1109 = ~n1105 & n1108;
  assign n1110 = ~pi22  & pi149 ;
  assign n1111 = ~pi150  & ~pi151 ;
  assign n1112 = ~n1110 & n1111;
  assign n1113 = ~n1109 & n1112;
  assign n1114 = pi23  & ~pi151 ;
  assign n1115 = ~pi24  & ~n1114;
  assign n1116 = ~pi25  & n1115;
  assign n1117 = ~n1113 & n1116;
  assign n1118 = ~pi25  & pi152 ;
  assign n1119 = ~pi153  & ~pi154 ;
  assign n1120 = ~n1118 & n1119;
  assign n1121 = ~n1117 & n1120;
  assign n1122 = pi26  & ~pi154 ;
  assign n1123 = ~pi27  & ~n1122;
  assign n1124 = ~pi28  & n1123;
  assign n1125 = ~n1121 & n1124;
  assign n1126 = ~pi28  & pi155 ;
  assign n1127 = ~pi156  & ~pi157 ;
  assign n1128 = ~n1126 & n1127;
  assign n1129 = ~n1125 & n1128;
  assign n1130 = pi29  & ~pi157 ;
  assign n1131 = ~pi30  & ~n1130;
  assign n1132 = ~pi31  & n1131;
  assign n1133 = ~n1129 & n1132;
  assign n1134 = ~pi31  & pi158 ;
  assign n1135 = ~pi159  & ~pi160 ;
  assign n1136 = ~n1134 & n1135;
  assign n1137 = ~n1133 & n1136;
  assign n1138 = pi32  & ~pi160 ;
  assign n1139 = ~pi33  & ~n1138;
  assign n1140 = ~pi34  & n1139;
  assign n1141 = ~n1137 & n1140;
  assign n1142 = ~pi34  & pi161 ;
  assign n1143 = ~pi162  & ~pi163 ;
  assign n1144 = ~n1142 & n1143;
  assign n1145 = ~n1141 & n1144;
  assign n1146 = pi35  & ~pi163 ;
  assign n1147 = ~pi36  & ~n1146;
  assign n1148 = ~pi37  & n1147;
  assign n1149 = ~n1145 & n1148;
  assign n1150 = ~pi37  & pi164 ;
  assign n1151 = ~pi165  & ~pi166 ;
  assign n1152 = ~n1150 & n1151;
  assign n1153 = ~n1149 & n1152;
  assign n1154 = pi38  & ~pi166 ;
  assign n1155 = ~pi39  & ~n1154;
  assign n1156 = ~pi40  & n1155;
  assign n1157 = ~n1153 & n1156;
  assign n1158 = ~pi40  & pi167 ;
  assign n1159 = ~pi168  & ~pi169 ;
  assign n1160 = ~n1158 & n1159;
  assign n1161 = ~n1157 & n1160;
  assign n1162 = pi41  & ~pi169 ;
  assign n1163 = ~pi42  & ~n1162;
  assign n1164 = ~pi43  & n1163;
  assign n1165 = ~n1161 & n1164;
  assign n1166 = ~pi43  & pi170 ;
  assign n1167 = ~pi171  & ~pi172 ;
  assign n1168 = ~n1166 & n1167;
  assign n1169 = ~n1165 & n1168;
  assign n1170 = pi44  & ~pi172 ;
  assign n1171 = ~pi45  & ~n1170;
  assign n1172 = ~pi46  & n1171;
  assign n1173 = ~n1169 & n1172;
  assign n1174 = ~pi46  & pi173 ;
  assign n1175 = ~pi174  & ~pi175 ;
  assign n1176 = ~n1174 & n1175;
  assign n1177 = ~n1173 & n1176;
  assign n1178 = pi47  & ~pi175 ;
  assign n1179 = ~pi48  & ~n1178;
  assign n1180 = ~pi49  & n1179;
  assign n1181 = ~n1177 & n1180;
  assign n1182 = ~pi49  & pi176 ;
  assign n1183 = ~pi177  & ~pi178 ;
  assign n1184 = ~n1182 & n1183;
  assign n1185 = ~n1181 & n1184;
  assign n1186 = pi50  & ~pi178 ;
  assign n1187 = ~pi51  & ~n1186;
  assign n1188 = ~pi52  & n1187;
  assign n1189 = ~n1185 & n1188;
  assign n1190 = ~pi52  & pi179 ;
  assign n1191 = ~pi180  & ~pi181 ;
  assign n1192 = ~n1190 & n1191;
  assign n1193 = ~n1189 & n1192;
  assign n1194 = pi53  & ~pi181 ;
  assign n1195 = ~pi54  & ~n1194;
  assign n1196 = ~pi55  & n1195;
  assign n1197 = ~n1193 & n1196;
  assign n1198 = ~pi55  & pi182 ;
  assign n1199 = ~pi183  & ~pi184 ;
  assign n1200 = ~n1198 & n1199;
  assign n1201 = ~n1197 & n1200;
  assign n1202 = pi56  & ~pi184 ;
  assign n1203 = ~pi57  & ~n1202;
  assign n1204 = ~pi58  & n1203;
  assign n1205 = ~n1201 & n1204;
  assign n1206 = ~pi58  & pi185 ;
  assign n1207 = ~pi186  & ~pi187 ;
  assign n1208 = ~n1206 & n1207;
  assign n1209 = ~n1205 & n1208;
  assign n1210 = pi59  & ~pi187 ;
  assign n1211 = ~pi60  & ~n1210;
  assign n1212 = ~pi61  & n1211;
  assign n1213 = ~n1209 & n1212;
  assign n1214 = ~pi61  & pi188 ;
  assign n1215 = ~pi189  & ~pi190 ;
  assign n1216 = ~n1214 & n1215;
  assign n1217 = ~n1213 & n1216;
  assign n1218 = pi62  & ~pi190 ;
  assign n1219 = ~pi63  & ~n1218;
  assign n1220 = ~pi64  & n1219;
  assign n1221 = ~n1217 & n1220;
  assign n1222 = ~pi64  & pi191 ;
  assign n1223 = ~pi192  & ~pi193 ;
  assign n1224 = ~n1222 & n1223;
  assign n1225 = ~n1221 & n1224;
  assign n1226 = pi65  & ~pi193 ;
  assign n1227 = ~pi66  & ~n1226;
  assign n1228 = ~pi67  & n1227;
  assign n1229 = ~n1225 & n1228;
  assign n1230 = ~pi67  & pi194 ;
  assign n1231 = ~pi195  & ~pi196 ;
  assign n1232 = ~n1230 & n1231;
  assign n1233 = ~n1229 & n1232;
  assign n1234 = pi68  & ~pi196 ;
  assign n1235 = ~pi69  & ~n1234;
  assign n1236 = ~pi70  & n1235;
  assign n1237 = ~n1233 & n1236;
  assign n1238 = ~pi70  & pi197 ;
  assign n1239 = ~pi198  & ~pi199 ;
  assign n1240 = ~n1238 & n1239;
  assign n1241 = ~n1237 & n1240;
  assign n1242 = pi71  & ~pi199 ;
  assign n1243 = ~pi72  & ~n1242;
  assign n1244 = ~pi73  & n1243;
  assign n1245 = ~n1241 & n1244;
  assign n1246 = ~pi73  & pi200 ;
  assign n1247 = ~pi201  & ~pi202 ;
  assign n1248 = ~n1246 & n1247;
  assign n1249 = ~n1245 & n1248;
  assign n1250 = pi74  & ~pi202 ;
  assign n1251 = ~pi75  & ~n1250;
  assign n1252 = ~pi76  & n1251;
  assign n1253 = ~n1249 & n1252;
  assign n1254 = ~pi76  & pi203 ;
  assign n1255 = ~pi204  & ~pi205 ;
  assign n1256 = ~n1254 & n1255;
  assign n1257 = ~n1253 & n1256;
  assign n1258 = pi77  & ~pi205 ;
  assign n1259 = ~pi78  & ~n1258;
  assign n1260 = ~pi79  & n1259;
  assign n1261 = ~n1257 & n1260;
  assign n1262 = ~pi79  & pi206 ;
  assign n1263 = ~pi207  & ~pi208 ;
  assign n1264 = ~n1262 & n1263;
  assign n1265 = ~n1261 & n1264;
  assign n1266 = pi80  & ~pi208 ;
  assign n1267 = ~pi81  & ~n1266;
  assign n1268 = ~pi82  & n1267;
  assign n1269 = ~n1265 & n1268;
  assign n1270 = ~pi82  & pi209 ;
  assign n1271 = ~pi210  & ~pi211 ;
  assign n1272 = ~n1270 & n1271;
  assign n1273 = ~n1269 & n1272;
  assign n1274 = pi83  & ~pi211 ;
  assign n1275 = ~pi84  & ~n1274;
  assign n1276 = ~pi85  & n1275;
  assign n1277 = ~n1273 & n1276;
  assign n1278 = ~pi85  & pi212 ;
  assign n1279 = ~pi213  & ~pi214 ;
  assign n1280 = ~n1278 & n1279;
  assign n1281 = ~n1277 & n1280;
  assign n1282 = pi86  & ~pi214 ;
  assign n1283 = ~pi87  & ~n1282;
  assign n1284 = ~pi88  & n1283;
  assign n1285 = ~n1281 & n1284;
  assign n1286 = ~pi88  & pi215 ;
  assign n1287 = ~pi216  & ~pi217 ;
  assign n1288 = ~n1286 & n1287;
  assign n1289 = ~n1285 & n1288;
  assign n1290 = pi89  & ~pi217 ;
  assign n1291 = ~pi90  & ~n1290;
  assign n1292 = ~pi91  & n1291;
  assign n1293 = ~n1289 & n1292;
  assign n1294 = ~pi91  & pi218 ;
  assign n1295 = ~pi219  & ~pi220 ;
  assign n1296 = ~n1294 & n1295;
  assign n1297 = ~n1293 & n1296;
  assign n1298 = pi92  & ~pi220 ;
  assign n1299 = ~pi93  & ~n1298;
  assign n1300 = ~pi94  & n1299;
  assign n1301 = ~n1297 & n1300;
  assign n1302 = ~pi94  & pi221 ;
  assign n1303 = ~pi222  & ~pi223 ;
  assign n1304 = ~n1302 & n1303;
  assign n1305 = ~n1301 & n1304;
  assign n1306 = pi95  & ~pi223 ;
  assign n1307 = ~pi96  & ~n1306;
  assign n1308 = ~pi97  & n1307;
  assign n1309 = ~n1305 & n1308;
  assign n1310 = ~pi97  & pi224 ;
  assign n1311 = ~pi225  & ~pi226 ;
  assign n1312 = ~n1310 & n1311;
  assign n1313 = ~n1309 & n1312;
  assign n1314 = pi98  & ~pi226 ;
  assign n1315 = ~pi99  & ~n1314;
  assign n1316 = ~pi100  & n1315;
  assign n1317 = ~n1313 & n1316;
  assign n1318 = ~pi100  & pi227 ;
  assign n1319 = ~pi228  & ~pi229 ;
  assign n1320 = ~n1318 & n1319;
  assign n1321 = ~n1317 & n1320;
  assign n1322 = pi101  & ~pi229 ;
  assign n1323 = ~pi102  & ~n1322;
  assign n1324 = ~pi103  & n1323;
  assign n1325 = ~n1321 & n1324;
  assign n1326 = ~pi103  & pi230 ;
  assign n1327 = ~pi231  & ~pi232 ;
  assign n1328 = ~n1326 & n1327;
  assign n1329 = ~n1325 & n1328;
  assign n1330 = pi104  & ~pi232 ;
  assign n1331 = ~pi105  & ~n1330;
  assign n1332 = ~pi106  & n1331;
  assign n1333 = ~n1329 & n1332;
  assign n1334 = ~pi106  & pi233 ;
  assign n1335 = ~pi234  & ~pi235 ;
  assign n1336 = ~n1334 & n1335;
  assign n1337 = ~n1333 & n1336;
  assign n1338 = pi107  & ~pi235 ;
  assign n1339 = ~pi108  & ~n1338;
  assign n1340 = ~pi109  & n1339;
  assign n1341 = ~n1337 & n1340;
  assign n1342 = ~pi109  & pi236 ;
  assign n1343 = ~pi237  & ~pi238 ;
  assign n1344 = ~n1342 & n1343;
  assign n1345 = ~n1341 & n1344;
  assign n1346 = pi110  & ~pi238 ;
  assign n1347 = ~pi111  & ~n1346;
  assign n1348 = ~pi112  & n1347;
  assign n1349 = ~n1345 & n1348;
  assign n1350 = ~pi112  & pi239 ;
  assign n1351 = ~pi240  & ~pi241 ;
  assign n1352 = ~n1350 & n1351;
  assign n1353 = ~n1349 & n1352;
  assign n1354 = pi113  & ~pi241 ;
  assign n1355 = ~pi114  & ~n1354;
  assign n1356 = ~pi115  & n1355;
  assign n1357 = ~n1353 & n1356;
  assign n1358 = ~pi115  & pi242 ;
  assign n1359 = ~pi243  & ~pi244 ;
  assign n1360 = ~n1358 & n1359;
  assign n1361 = ~n1357 & n1360;
  assign n1362 = pi116  & ~pi244 ;
  assign n1363 = ~pi117  & ~n1362;
  assign n1364 = ~pi118  & n1363;
  assign n1365 = ~n1361 & n1364;
  assign n1366 = ~pi118  & pi245 ;
  assign n1367 = ~pi246  & ~pi247 ;
  assign n1368 = ~n1366 & n1367;
  assign n1369 = ~n1365 & n1368;
  assign n1370 = pi119  & ~pi247 ;
  assign n1371 = ~pi120  & ~n1370;
  assign n1372 = ~pi121  & n1371;
  assign n1373 = ~n1369 & n1372;
  assign n1374 = ~pi121  & pi248 ;
  assign n1375 = ~pi249  & ~pi250 ;
  assign n1376 = ~n1374 & n1375;
  assign n1377 = ~n1373 & n1376;
  assign n1378 = pi122  & ~pi250 ;
  assign n1379 = ~pi123  & ~n1378;
  assign n1380 = ~pi124  & n1379;
  assign n1381 = ~n1377 & n1380;
  assign n1382 = ~pi124  & pi251 ;
  assign n1383 = ~pi252  & ~pi253 ;
  assign n1384 = ~n1382 & n1383;
  assign n1385 = ~n1381 & n1384;
  assign n1386 = pi125  & ~pi253 ;
  assign n1387 = ~pi126  & ~n1386;
  assign n1388 = ~pi127  & n1387;
  assign n1389 = ~n1385 & n1388;
  assign n1390 = ~pi127  & pi254 ;
  assign n1391 = ~pi128  & ~pi255 ;
  assign n1392 = ~n1390 & n1391;
  assign n1393 = ~n1389 & n1392;
  assign n1394 = pi0  & ~pi128 ;
  assign n1395 = ~pi1  & ~n1394;
  assign n1396 = ~pi2  & n1395;
  assign n1397 = ~n1393 & n1396;
  assign n1398 = ~pi2  & pi129 ;
  assign n1399 = pi130  & ~n1398;
  assign po2  = ~n1397 & n1399;
  assign n1401 = n395 & ~n730;
  assign n1402 = n400 & ~n1401;
  assign n1403 = n404 & ~n1402;
  assign n1404 = n408 & ~n1403;
  assign n1405 = n412 & ~n1404;
  assign n1406 = n416 & ~n1405;
  assign n1407 = n420 & ~n1406;
  assign n1408 = n424 & ~n1407;
  assign n1409 = n428 & ~n1408;
  assign n1410 = n432 & ~n1409;
  assign n1411 = n436 & ~n1410;
  assign n1412 = n440 & ~n1411;
  assign n1413 = n444 & ~n1412;
  assign n1414 = n448 & ~n1413;
  assign n1415 = n452 & ~n1414;
  assign n1416 = n456 & ~n1415;
  assign n1417 = n460 & ~n1416;
  assign n1418 = n464 & ~n1417;
  assign n1419 = n468 & ~n1418;
  assign n1420 = n472 & ~n1419;
  assign n1421 = n476 & ~n1420;
  assign n1422 = n480 & ~n1421;
  assign n1423 = n484 & ~n1422;
  assign n1424 = n488 & ~n1423;
  assign n1425 = n492 & ~n1424;
  assign n1426 = n496 & ~n1425;
  assign n1427 = n500 & ~n1426;
  assign n1428 = n504 & ~n1427;
  assign n1429 = n508 & ~n1428;
  assign n1430 = n512 & ~n1429;
  assign n1431 = n516 & ~n1430;
  assign n1432 = n520 & ~n1431;
  assign n1433 = n524 & ~n1432;
  assign n1434 = n528 & ~n1433;
  assign n1435 = n532 & ~n1434;
  assign n1436 = n536 & ~n1435;
  assign n1437 = n540 & ~n1436;
  assign n1438 = n544 & ~n1437;
  assign n1439 = n548 & ~n1438;
  assign n1440 = n552 & ~n1439;
  assign n1441 = n556 & ~n1440;
  assign n1442 = n560 & ~n1441;
  assign n1443 = n564 & ~n1442;
  assign n1444 = n568 & ~n1443;
  assign n1445 = n572 & ~n1444;
  assign n1446 = n576 & ~n1445;
  assign n1447 = n580 & ~n1446;
  assign n1448 = n584 & ~n1447;
  assign n1449 = n588 & ~n1448;
  assign n1450 = n592 & ~n1449;
  assign n1451 = n596 & ~n1450;
  assign n1452 = n600 & ~n1451;
  assign n1453 = n604 & ~n1452;
  assign n1454 = n608 & ~n1453;
  assign n1455 = n612 & ~n1454;
  assign n1456 = n616 & ~n1455;
  assign n1457 = n620 & ~n1456;
  assign n1458 = n624 & ~n1457;
  assign n1459 = n628 & ~n1458;
  assign n1460 = n632 & ~n1459;
  assign n1461 = n636 & ~n1460;
  assign n1462 = n640 & ~n1461;
  assign n1463 = n644 & ~n1462;
  assign n1464 = n648 & ~n1463;
  assign n1465 = n652 & ~n1464;
  assign n1466 = n656 & ~n1465;
  assign n1467 = n660 & ~n1466;
  assign n1468 = n664 & ~n1467;
  assign n1469 = n668 & ~n1468;
  assign n1470 = n672 & ~n1469;
  assign n1471 = n676 & ~n1470;
  assign n1472 = n680 & ~n1471;
  assign n1473 = n684 & ~n1472;
  assign n1474 = n688 & ~n1473;
  assign n1475 = n692 & ~n1474;
  assign n1476 = n696 & ~n1475;
  assign n1477 = n700 & ~n1476;
  assign n1478 = n704 & ~n1477;
  assign n1479 = n708 & ~n1478;
  assign n1480 = n712 & ~n1479;
  assign n1481 = n716 & ~n1480;
  assign n1482 = n720 & ~n1481;
  assign n1483 = ~pi128  & ~pi129 ;
  assign n1484 = ~n722 & n1483;
  assign n1485 = ~n1482 & n1484;
  assign n1486 = ~pi3  & n387;
  assign n1487 = ~n1485 & n1486;
  assign n1488 = ~pi3  & pi130 ;
  assign n1489 = pi131  & ~n1488;
  assign po3  = ~n1487 & n1489;
  assign n1491 = n734 & ~n1067;
  assign n1492 = n739 & ~n1491;
  assign n1493 = n743 & ~n1492;
  assign n1494 = n747 & ~n1493;
  assign n1495 = n751 & ~n1494;
  assign n1496 = n755 & ~n1495;
  assign n1497 = n759 & ~n1496;
  assign n1498 = n763 & ~n1497;
  assign n1499 = n767 & ~n1498;
  assign n1500 = n771 & ~n1499;
  assign n1501 = n775 & ~n1500;
  assign n1502 = n779 & ~n1501;
  assign n1503 = n783 & ~n1502;
  assign n1504 = n787 & ~n1503;
  assign n1505 = n791 & ~n1504;
  assign n1506 = n795 & ~n1505;
  assign n1507 = n799 & ~n1506;
  assign n1508 = n803 & ~n1507;
  assign n1509 = n807 & ~n1508;
  assign n1510 = n811 & ~n1509;
  assign n1511 = n815 & ~n1510;
  assign n1512 = n819 & ~n1511;
  assign n1513 = n823 & ~n1512;
  assign n1514 = n827 & ~n1513;
  assign n1515 = n831 & ~n1514;
  assign n1516 = n835 & ~n1515;
  assign n1517 = n839 & ~n1516;
  assign n1518 = n843 & ~n1517;
  assign n1519 = n847 & ~n1518;
  assign n1520 = n851 & ~n1519;
  assign n1521 = n855 & ~n1520;
  assign n1522 = n859 & ~n1521;
  assign n1523 = n863 & ~n1522;
  assign n1524 = n867 & ~n1523;
  assign n1525 = n871 & ~n1524;
  assign n1526 = n875 & ~n1525;
  assign n1527 = n879 & ~n1526;
  assign n1528 = n883 & ~n1527;
  assign n1529 = n887 & ~n1528;
  assign n1530 = n891 & ~n1529;
  assign n1531 = n895 & ~n1530;
  assign n1532 = n899 & ~n1531;
  assign n1533 = n903 & ~n1532;
  assign n1534 = n907 & ~n1533;
  assign n1535 = n911 & ~n1534;
  assign n1536 = n915 & ~n1535;
  assign n1537 = n919 & ~n1536;
  assign n1538 = n923 & ~n1537;
  assign n1539 = n927 & ~n1538;
  assign n1540 = n931 & ~n1539;
  assign n1541 = n935 & ~n1540;
  assign n1542 = n939 & ~n1541;
  assign n1543 = n943 & ~n1542;
  assign n1544 = n947 & ~n1543;
  assign n1545 = n951 & ~n1544;
  assign n1546 = n955 & ~n1545;
  assign n1547 = n959 & ~n1546;
  assign n1548 = n963 & ~n1547;
  assign n1549 = n967 & ~n1548;
  assign n1550 = n971 & ~n1549;
  assign n1551 = n975 & ~n1550;
  assign n1552 = n979 & ~n1551;
  assign n1553 = n983 & ~n1552;
  assign n1554 = n987 & ~n1553;
  assign n1555 = n991 & ~n1554;
  assign n1556 = n995 & ~n1555;
  assign n1557 = n999 & ~n1556;
  assign n1558 = n1003 & ~n1557;
  assign n1559 = n1007 & ~n1558;
  assign n1560 = n1011 & ~n1559;
  assign n1561 = n1015 & ~n1560;
  assign n1562 = n1019 & ~n1561;
  assign n1563 = n1023 & ~n1562;
  assign n1564 = n1027 & ~n1563;
  assign n1565 = n1031 & ~n1564;
  assign n1566 = n1035 & ~n1565;
  assign n1567 = n1039 & ~n1566;
  assign n1568 = n1043 & ~n1567;
  assign n1569 = n1047 & ~n1568;
  assign n1570 = n1051 & ~n1569;
  assign n1571 = n1055 & ~n1570;
  assign n1572 = n1059 & ~n1571;
  assign n1573 = ~pi129  & ~pi130 ;
  assign n1574 = ~n1061 & n1573;
  assign n1575 = ~n1572 & n1574;
  assign n1576 = ~pi4  & n726;
  assign n1577 = ~n1575 & n1576;
  assign n1578 = ~pi4  & pi131 ;
  assign n1579 = pi132  & ~n1578;
  assign po4  = ~n1577 & n1579;
  assign n1581 = ~n399 & n1071;
  assign n1582 = n1076 & ~n1581;
  assign n1583 = n1080 & ~n1582;
  assign n1584 = n1084 & ~n1583;
  assign n1585 = n1088 & ~n1584;
  assign n1586 = n1092 & ~n1585;
  assign n1587 = n1096 & ~n1586;
  assign n1588 = n1100 & ~n1587;
  assign n1589 = n1104 & ~n1588;
  assign n1590 = n1108 & ~n1589;
  assign n1591 = n1112 & ~n1590;
  assign n1592 = n1116 & ~n1591;
  assign n1593 = n1120 & ~n1592;
  assign n1594 = n1124 & ~n1593;
  assign n1595 = n1128 & ~n1594;
  assign n1596 = n1132 & ~n1595;
  assign n1597 = n1136 & ~n1596;
  assign n1598 = n1140 & ~n1597;
  assign n1599 = n1144 & ~n1598;
  assign n1600 = n1148 & ~n1599;
  assign n1601 = n1152 & ~n1600;
  assign n1602 = n1156 & ~n1601;
  assign n1603 = n1160 & ~n1602;
  assign n1604 = n1164 & ~n1603;
  assign n1605 = n1168 & ~n1604;
  assign n1606 = n1172 & ~n1605;
  assign n1607 = n1176 & ~n1606;
  assign n1608 = n1180 & ~n1607;
  assign n1609 = n1184 & ~n1608;
  assign n1610 = n1188 & ~n1609;
  assign n1611 = n1192 & ~n1610;
  assign n1612 = n1196 & ~n1611;
  assign n1613 = n1200 & ~n1612;
  assign n1614 = n1204 & ~n1613;
  assign n1615 = n1208 & ~n1614;
  assign n1616 = n1212 & ~n1615;
  assign n1617 = n1216 & ~n1616;
  assign n1618 = n1220 & ~n1617;
  assign n1619 = n1224 & ~n1618;
  assign n1620 = n1228 & ~n1619;
  assign n1621 = n1232 & ~n1620;
  assign n1622 = n1236 & ~n1621;
  assign n1623 = n1240 & ~n1622;
  assign n1624 = n1244 & ~n1623;
  assign n1625 = n1248 & ~n1624;
  assign n1626 = n1252 & ~n1625;
  assign n1627 = n1256 & ~n1626;
  assign n1628 = n1260 & ~n1627;
  assign n1629 = n1264 & ~n1628;
  assign n1630 = n1268 & ~n1629;
  assign n1631 = n1272 & ~n1630;
  assign n1632 = n1276 & ~n1631;
  assign n1633 = n1280 & ~n1632;
  assign n1634 = n1284 & ~n1633;
  assign n1635 = n1288 & ~n1634;
  assign n1636 = n1292 & ~n1635;
  assign n1637 = n1296 & ~n1636;
  assign n1638 = n1300 & ~n1637;
  assign n1639 = n1304 & ~n1638;
  assign n1640 = n1308 & ~n1639;
  assign n1641 = n1312 & ~n1640;
  assign n1642 = n1316 & ~n1641;
  assign n1643 = n1320 & ~n1642;
  assign n1644 = n1324 & ~n1643;
  assign n1645 = n1328 & ~n1644;
  assign n1646 = n1332 & ~n1645;
  assign n1647 = n1336 & ~n1646;
  assign n1648 = n1340 & ~n1647;
  assign n1649 = n1344 & ~n1648;
  assign n1650 = n1348 & ~n1649;
  assign n1651 = n1352 & ~n1650;
  assign n1652 = n1356 & ~n1651;
  assign n1653 = n1360 & ~n1652;
  assign n1654 = n1364 & ~n1653;
  assign n1655 = n1368 & ~n1654;
  assign n1656 = n1372 & ~n1655;
  assign n1657 = n1376 & ~n1656;
  assign n1658 = n1380 & ~n1657;
  assign n1659 = n1384 & ~n1658;
  assign n1660 = n1388 & ~n1659;
  assign n1661 = n1392 & ~n1660;
  assign n1662 = n1396 & ~n1661;
  assign n1663 = n388 & ~n1398;
  assign n1664 = ~n1662 & n1663;
  assign n1665 = n392 & ~n1664;
  assign n1666 = pi133  & ~n394;
  assign po5  = ~n1665 & n1666;
  assign n1668 = n403 & ~n738;
  assign n1669 = n408 & ~n1668;
  assign n1670 = n412 & ~n1669;
  assign n1671 = n416 & ~n1670;
  assign n1672 = n420 & ~n1671;
  assign n1673 = n424 & ~n1672;
  assign n1674 = n428 & ~n1673;
  assign n1675 = n432 & ~n1674;
  assign n1676 = n436 & ~n1675;
  assign n1677 = n440 & ~n1676;
  assign n1678 = n444 & ~n1677;
  assign n1679 = n448 & ~n1678;
  assign n1680 = n452 & ~n1679;
  assign n1681 = n456 & ~n1680;
  assign n1682 = n460 & ~n1681;
  assign n1683 = n464 & ~n1682;
  assign n1684 = n468 & ~n1683;
  assign n1685 = n472 & ~n1684;
  assign n1686 = n476 & ~n1685;
  assign n1687 = n480 & ~n1686;
  assign n1688 = n484 & ~n1687;
  assign n1689 = n488 & ~n1688;
  assign n1690 = n492 & ~n1689;
  assign n1691 = n496 & ~n1690;
  assign n1692 = n500 & ~n1691;
  assign n1693 = n504 & ~n1692;
  assign n1694 = n508 & ~n1693;
  assign n1695 = n512 & ~n1694;
  assign n1696 = n516 & ~n1695;
  assign n1697 = n520 & ~n1696;
  assign n1698 = n524 & ~n1697;
  assign n1699 = n528 & ~n1698;
  assign n1700 = n532 & ~n1699;
  assign n1701 = n536 & ~n1700;
  assign n1702 = n540 & ~n1701;
  assign n1703 = n544 & ~n1702;
  assign n1704 = n548 & ~n1703;
  assign n1705 = n552 & ~n1704;
  assign n1706 = n556 & ~n1705;
  assign n1707 = n560 & ~n1706;
  assign n1708 = n564 & ~n1707;
  assign n1709 = n568 & ~n1708;
  assign n1710 = n572 & ~n1709;
  assign n1711 = n576 & ~n1710;
  assign n1712 = n580 & ~n1711;
  assign n1713 = n584 & ~n1712;
  assign n1714 = n588 & ~n1713;
  assign n1715 = n592 & ~n1714;
  assign n1716 = n596 & ~n1715;
  assign n1717 = n600 & ~n1716;
  assign n1718 = n604 & ~n1717;
  assign n1719 = n608 & ~n1718;
  assign n1720 = n612 & ~n1719;
  assign n1721 = n616 & ~n1720;
  assign n1722 = n620 & ~n1721;
  assign n1723 = n624 & ~n1722;
  assign n1724 = n628 & ~n1723;
  assign n1725 = n632 & ~n1724;
  assign n1726 = n636 & ~n1725;
  assign n1727 = n640 & ~n1726;
  assign n1728 = n644 & ~n1727;
  assign n1729 = n648 & ~n1728;
  assign n1730 = n652 & ~n1729;
  assign n1731 = n656 & ~n1730;
  assign n1732 = n660 & ~n1731;
  assign n1733 = n664 & ~n1732;
  assign n1734 = n668 & ~n1733;
  assign n1735 = n672 & ~n1734;
  assign n1736 = n676 & ~n1735;
  assign n1737 = n680 & ~n1736;
  assign n1738 = n684 & ~n1737;
  assign n1739 = n688 & ~n1738;
  assign n1740 = n692 & ~n1739;
  assign n1741 = n696 & ~n1740;
  assign n1742 = n700 & ~n1741;
  assign n1743 = n704 & ~n1742;
  assign n1744 = n708 & ~n1743;
  assign n1745 = n712 & ~n1744;
  assign n1746 = n716 & ~n1745;
  assign n1747 = n720 & ~n1746;
  assign n1748 = n1484 & ~n1747;
  assign n1749 = n1486 & ~n1748;
  assign n1750 = n727 & ~n1488;
  assign n1751 = ~n1749 & n1750;
  assign n1752 = n731 & ~n1751;
  assign n1753 = pi134  & ~n733;
  assign po6  = ~n1752 & n1753;
  assign n1755 = n742 & ~n1075;
  assign n1756 = n747 & ~n1755;
  assign n1757 = n751 & ~n1756;
  assign n1758 = n755 & ~n1757;
  assign n1759 = n759 & ~n1758;
  assign n1760 = n763 & ~n1759;
  assign n1761 = n767 & ~n1760;
  assign n1762 = n771 & ~n1761;
  assign n1763 = n775 & ~n1762;
  assign n1764 = n779 & ~n1763;
  assign n1765 = n783 & ~n1764;
  assign n1766 = n787 & ~n1765;
  assign n1767 = n791 & ~n1766;
  assign n1768 = n795 & ~n1767;
  assign n1769 = n799 & ~n1768;
  assign n1770 = n803 & ~n1769;
  assign n1771 = n807 & ~n1770;
  assign n1772 = n811 & ~n1771;
  assign n1773 = n815 & ~n1772;
  assign n1774 = n819 & ~n1773;
  assign n1775 = n823 & ~n1774;
  assign n1776 = n827 & ~n1775;
  assign n1777 = n831 & ~n1776;
  assign n1778 = n835 & ~n1777;
  assign n1779 = n839 & ~n1778;
  assign n1780 = n843 & ~n1779;
  assign n1781 = n847 & ~n1780;
  assign n1782 = n851 & ~n1781;
  assign n1783 = n855 & ~n1782;
  assign n1784 = n859 & ~n1783;
  assign n1785 = n863 & ~n1784;
  assign n1786 = n867 & ~n1785;
  assign n1787 = n871 & ~n1786;
  assign n1788 = n875 & ~n1787;
  assign n1789 = n879 & ~n1788;
  assign n1790 = n883 & ~n1789;
  assign n1791 = n887 & ~n1790;
  assign n1792 = n891 & ~n1791;
  assign n1793 = n895 & ~n1792;
  assign n1794 = n899 & ~n1793;
  assign n1795 = n903 & ~n1794;
  assign n1796 = n907 & ~n1795;
  assign n1797 = n911 & ~n1796;
  assign n1798 = n915 & ~n1797;
  assign n1799 = n919 & ~n1798;
  assign n1800 = n923 & ~n1799;
  assign n1801 = n927 & ~n1800;
  assign n1802 = n931 & ~n1801;
  assign n1803 = n935 & ~n1802;
  assign n1804 = n939 & ~n1803;
  assign n1805 = n943 & ~n1804;
  assign n1806 = n947 & ~n1805;
  assign n1807 = n951 & ~n1806;
  assign n1808 = n955 & ~n1807;
  assign n1809 = n959 & ~n1808;
  assign n1810 = n963 & ~n1809;
  assign n1811 = n967 & ~n1810;
  assign n1812 = n971 & ~n1811;
  assign n1813 = n975 & ~n1812;
  assign n1814 = n979 & ~n1813;
  assign n1815 = n983 & ~n1814;
  assign n1816 = n987 & ~n1815;
  assign n1817 = n991 & ~n1816;
  assign n1818 = n995 & ~n1817;
  assign n1819 = n999 & ~n1818;
  assign n1820 = n1003 & ~n1819;
  assign n1821 = n1007 & ~n1820;
  assign n1822 = n1011 & ~n1821;
  assign n1823 = n1015 & ~n1822;
  assign n1824 = n1019 & ~n1823;
  assign n1825 = n1023 & ~n1824;
  assign n1826 = n1027 & ~n1825;
  assign n1827 = n1031 & ~n1826;
  assign n1828 = n1035 & ~n1827;
  assign n1829 = n1039 & ~n1828;
  assign n1830 = n1043 & ~n1829;
  assign n1831 = n1047 & ~n1830;
  assign n1832 = n1051 & ~n1831;
  assign n1833 = n1055 & ~n1832;
  assign n1834 = n1059 & ~n1833;
  assign n1835 = n1574 & ~n1834;
  assign n1836 = n1576 & ~n1835;
  assign n1837 = n1064 & ~n1578;
  assign n1838 = ~n1836 & n1837;
  assign n1839 = n1068 & ~n1838;
  assign n1840 = pi135  & ~n1070;
  assign po7  = ~n1839 & n1840;
  assign n1842 = ~n407 & n1079;
  assign n1843 = n1084 & ~n1842;
  assign n1844 = n1088 & ~n1843;
  assign n1845 = n1092 & ~n1844;
  assign n1846 = n1096 & ~n1845;
  assign n1847 = n1100 & ~n1846;
  assign n1848 = n1104 & ~n1847;
  assign n1849 = n1108 & ~n1848;
  assign n1850 = n1112 & ~n1849;
  assign n1851 = n1116 & ~n1850;
  assign n1852 = n1120 & ~n1851;
  assign n1853 = n1124 & ~n1852;
  assign n1854 = n1128 & ~n1853;
  assign n1855 = n1132 & ~n1854;
  assign n1856 = n1136 & ~n1855;
  assign n1857 = n1140 & ~n1856;
  assign n1858 = n1144 & ~n1857;
  assign n1859 = n1148 & ~n1858;
  assign n1860 = n1152 & ~n1859;
  assign n1861 = n1156 & ~n1860;
  assign n1862 = n1160 & ~n1861;
  assign n1863 = n1164 & ~n1862;
  assign n1864 = n1168 & ~n1863;
  assign n1865 = n1172 & ~n1864;
  assign n1866 = n1176 & ~n1865;
  assign n1867 = n1180 & ~n1866;
  assign n1868 = n1184 & ~n1867;
  assign n1869 = n1188 & ~n1868;
  assign n1870 = n1192 & ~n1869;
  assign n1871 = n1196 & ~n1870;
  assign n1872 = n1200 & ~n1871;
  assign n1873 = n1204 & ~n1872;
  assign n1874 = n1208 & ~n1873;
  assign n1875 = n1212 & ~n1874;
  assign n1876 = n1216 & ~n1875;
  assign n1877 = n1220 & ~n1876;
  assign n1878 = n1224 & ~n1877;
  assign n1879 = n1228 & ~n1878;
  assign n1880 = n1232 & ~n1879;
  assign n1881 = n1236 & ~n1880;
  assign n1882 = n1240 & ~n1881;
  assign n1883 = n1244 & ~n1882;
  assign n1884 = n1248 & ~n1883;
  assign n1885 = n1252 & ~n1884;
  assign n1886 = n1256 & ~n1885;
  assign n1887 = n1260 & ~n1886;
  assign n1888 = n1264 & ~n1887;
  assign n1889 = n1268 & ~n1888;
  assign n1890 = n1272 & ~n1889;
  assign n1891 = n1276 & ~n1890;
  assign n1892 = n1280 & ~n1891;
  assign n1893 = n1284 & ~n1892;
  assign n1894 = n1288 & ~n1893;
  assign n1895 = n1292 & ~n1894;
  assign n1896 = n1296 & ~n1895;
  assign n1897 = n1300 & ~n1896;
  assign n1898 = n1304 & ~n1897;
  assign n1899 = n1308 & ~n1898;
  assign n1900 = n1312 & ~n1899;
  assign n1901 = n1316 & ~n1900;
  assign n1902 = n1320 & ~n1901;
  assign n1903 = n1324 & ~n1902;
  assign n1904 = n1328 & ~n1903;
  assign n1905 = n1332 & ~n1904;
  assign n1906 = n1336 & ~n1905;
  assign n1907 = n1340 & ~n1906;
  assign n1908 = n1344 & ~n1907;
  assign n1909 = n1348 & ~n1908;
  assign n1910 = n1352 & ~n1909;
  assign n1911 = n1356 & ~n1910;
  assign n1912 = n1360 & ~n1911;
  assign n1913 = n1364 & ~n1912;
  assign n1914 = n1368 & ~n1913;
  assign n1915 = n1372 & ~n1914;
  assign n1916 = n1376 & ~n1915;
  assign n1917 = n1380 & ~n1916;
  assign n1918 = n1384 & ~n1917;
  assign n1919 = n1388 & ~n1918;
  assign n1920 = n1392 & ~n1919;
  assign n1921 = n1396 & ~n1920;
  assign n1922 = n1663 & ~n1921;
  assign n1923 = n392 & ~n1922;
  assign n1924 = n396 & ~n1923;
  assign n1925 = n400 & ~n1924;
  assign n1926 = pi136  & ~n402;
  assign po8  = ~n1925 & n1926;
  assign n1928 = n411 & ~n746;
  assign n1929 = n416 & ~n1928;
  assign n1930 = n420 & ~n1929;
  assign n1931 = n424 & ~n1930;
  assign n1932 = n428 & ~n1931;
  assign n1933 = n432 & ~n1932;
  assign n1934 = n436 & ~n1933;
  assign n1935 = n440 & ~n1934;
  assign n1936 = n444 & ~n1935;
  assign n1937 = n448 & ~n1936;
  assign n1938 = n452 & ~n1937;
  assign n1939 = n456 & ~n1938;
  assign n1940 = n460 & ~n1939;
  assign n1941 = n464 & ~n1940;
  assign n1942 = n468 & ~n1941;
  assign n1943 = n472 & ~n1942;
  assign n1944 = n476 & ~n1943;
  assign n1945 = n480 & ~n1944;
  assign n1946 = n484 & ~n1945;
  assign n1947 = n488 & ~n1946;
  assign n1948 = n492 & ~n1947;
  assign n1949 = n496 & ~n1948;
  assign n1950 = n500 & ~n1949;
  assign n1951 = n504 & ~n1950;
  assign n1952 = n508 & ~n1951;
  assign n1953 = n512 & ~n1952;
  assign n1954 = n516 & ~n1953;
  assign n1955 = n520 & ~n1954;
  assign n1956 = n524 & ~n1955;
  assign n1957 = n528 & ~n1956;
  assign n1958 = n532 & ~n1957;
  assign n1959 = n536 & ~n1958;
  assign n1960 = n540 & ~n1959;
  assign n1961 = n544 & ~n1960;
  assign n1962 = n548 & ~n1961;
  assign n1963 = n552 & ~n1962;
  assign n1964 = n556 & ~n1963;
  assign n1965 = n560 & ~n1964;
  assign n1966 = n564 & ~n1965;
  assign n1967 = n568 & ~n1966;
  assign n1968 = n572 & ~n1967;
  assign n1969 = n576 & ~n1968;
  assign n1970 = n580 & ~n1969;
  assign n1971 = n584 & ~n1970;
  assign n1972 = n588 & ~n1971;
  assign n1973 = n592 & ~n1972;
  assign n1974 = n596 & ~n1973;
  assign n1975 = n600 & ~n1974;
  assign n1976 = n604 & ~n1975;
  assign n1977 = n608 & ~n1976;
  assign n1978 = n612 & ~n1977;
  assign n1979 = n616 & ~n1978;
  assign n1980 = n620 & ~n1979;
  assign n1981 = n624 & ~n1980;
  assign n1982 = n628 & ~n1981;
  assign n1983 = n632 & ~n1982;
  assign n1984 = n636 & ~n1983;
  assign n1985 = n640 & ~n1984;
  assign n1986 = n644 & ~n1985;
  assign n1987 = n648 & ~n1986;
  assign n1988 = n652 & ~n1987;
  assign n1989 = n656 & ~n1988;
  assign n1990 = n660 & ~n1989;
  assign n1991 = n664 & ~n1990;
  assign n1992 = n668 & ~n1991;
  assign n1993 = n672 & ~n1992;
  assign n1994 = n676 & ~n1993;
  assign n1995 = n680 & ~n1994;
  assign n1996 = n684 & ~n1995;
  assign n1997 = n688 & ~n1996;
  assign n1998 = n692 & ~n1997;
  assign n1999 = n696 & ~n1998;
  assign n2000 = n700 & ~n1999;
  assign n2001 = n704 & ~n2000;
  assign n2002 = n708 & ~n2001;
  assign n2003 = n712 & ~n2002;
  assign n2004 = n716 & ~n2003;
  assign n2005 = n720 & ~n2004;
  assign n2006 = n1484 & ~n2005;
  assign n2007 = n1486 & ~n2006;
  assign n2008 = n1750 & ~n2007;
  assign n2009 = n731 & ~n2008;
  assign n2010 = n735 & ~n2009;
  assign n2011 = n739 & ~n2010;
  assign n2012 = pi137  & ~n741;
  assign po9  = ~n2011 & n2012;
  assign n2014 = n750 & ~n1083;
  assign n2015 = n755 & ~n2014;
  assign n2016 = n759 & ~n2015;
  assign n2017 = n763 & ~n2016;
  assign n2018 = n767 & ~n2017;
  assign n2019 = n771 & ~n2018;
  assign n2020 = n775 & ~n2019;
  assign n2021 = n779 & ~n2020;
  assign n2022 = n783 & ~n2021;
  assign n2023 = n787 & ~n2022;
  assign n2024 = n791 & ~n2023;
  assign n2025 = n795 & ~n2024;
  assign n2026 = n799 & ~n2025;
  assign n2027 = n803 & ~n2026;
  assign n2028 = n807 & ~n2027;
  assign n2029 = n811 & ~n2028;
  assign n2030 = n815 & ~n2029;
  assign n2031 = n819 & ~n2030;
  assign n2032 = n823 & ~n2031;
  assign n2033 = n827 & ~n2032;
  assign n2034 = n831 & ~n2033;
  assign n2035 = n835 & ~n2034;
  assign n2036 = n839 & ~n2035;
  assign n2037 = n843 & ~n2036;
  assign n2038 = n847 & ~n2037;
  assign n2039 = n851 & ~n2038;
  assign n2040 = n855 & ~n2039;
  assign n2041 = n859 & ~n2040;
  assign n2042 = n863 & ~n2041;
  assign n2043 = n867 & ~n2042;
  assign n2044 = n871 & ~n2043;
  assign n2045 = n875 & ~n2044;
  assign n2046 = n879 & ~n2045;
  assign n2047 = n883 & ~n2046;
  assign n2048 = n887 & ~n2047;
  assign n2049 = n891 & ~n2048;
  assign n2050 = n895 & ~n2049;
  assign n2051 = n899 & ~n2050;
  assign n2052 = n903 & ~n2051;
  assign n2053 = n907 & ~n2052;
  assign n2054 = n911 & ~n2053;
  assign n2055 = n915 & ~n2054;
  assign n2056 = n919 & ~n2055;
  assign n2057 = n923 & ~n2056;
  assign n2058 = n927 & ~n2057;
  assign n2059 = n931 & ~n2058;
  assign n2060 = n935 & ~n2059;
  assign n2061 = n939 & ~n2060;
  assign n2062 = n943 & ~n2061;
  assign n2063 = n947 & ~n2062;
  assign n2064 = n951 & ~n2063;
  assign n2065 = n955 & ~n2064;
  assign n2066 = n959 & ~n2065;
  assign n2067 = n963 & ~n2066;
  assign n2068 = n967 & ~n2067;
  assign n2069 = n971 & ~n2068;
  assign n2070 = n975 & ~n2069;
  assign n2071 = n979 & ~n2070;
  assign n2072 = n983 & ~n2071;
  assign n2073 = n987 & ~n2072;
  assign n2074 = n991 & ~n2073;
  assign n2075 = n995 & ~n2074;
  assign n2076 = n999 & ~n2075;
  assign n2077 = n1003 & ~n2076;
  assign n2078 = n1007 & ~n2077;
  assign n2079 = n1011 & ~n2078;
  assign n2080 = n1015 & ~n2079;
  assign n2081 = n1019 & ~n2080;
  assign n2082 = n1023 & ~n2081;
  assign n2083 = n1027 & ~n2082;
  assign n2084 = n1031 & ~n2083;
  assign n2085 = n1035 & ~n2084;
  assign n2086 = n1039 & ~n2085;
  assign n2087 = n1043 & ~n2086;
  assign n2088 = n1047 & ~n2087;
  assign n2089 = n1051 & ~n2088;
  assign n2090 = n1055 & ~n2089;
  assign n2091 = n1059 & ~n2090;
  assign n2092 = n1574 & ~n2091;
  assign n2093 = n1576 & ~n2092;
  assign n2094 = n1837 & ~n2093;
  assign n2095 = n1068 & ~n2094;
  assign n2096 = n1072 & ~n2095;
  assign n2097 = n1076 & ~n2096;
  assign n2098 = pi138  & ~n1078;
  assign po10  = ~n2097 & n2098;
  assign n2100 = ~n415 & n1087;
  assign n2101 = n1092 & ~n2100;
  assign n2102 = n1096 & ~n2101;
  assign n2103 = n1100 & ~n2102;
  assign n2104 = n1104 & ~n2103;
  assign n2105 = n1108 & ~n2104;
  assign n2106 = n1112 & ~n2105;
  assign n2107 = n1116 & ~n2106;
  assign n2108 = n1120 & ~n2107;
  assign n2109 = n1124 & ~n2108;
  assign n2110 = n1128 & ~n2109;
  assign n2111 = n1132 & ~n2110;
  assign n2112 = n1136 & ~n2111;
  assign n2113 = n1140 & ~n2112;
  assign n2114 = n1144 & ~n2113;
  assign n2115 = n1148 & ~n2114;
  assign n2116 = n1152 & ~n2115;
  assign n2117 = n1156 & ~n2116;
  assign n2118 = n1160 & ~n2117;
  assign n2119 = n1164 & ~n2118;
  assign n2120 = n1168 & ~n2119;
  assign n2121 = n1172 & ~n2120;
  assign n2122 = n1176 & ~n2121;
  assign n2123 = n1180 & ~n2122;
  assign n2124 = n1184 & ~n2123;
  assign n2125 = n1188 & ~n2124;
  assign n2126 = n1192 & ~n2125;
  assign n2127 = n1196 & ~n2126;
  assign n2128 = n1200 & ~n2127;
  assign n2129 = n1204 & ~n2128;
  assign n2130 = n1208 & ~n2129;
  assign n2131 = n1212 & ~n2130;
  assign n2132 = n1216 & ~n2131;
  assign n2133 = n1220 & ~n2132;
  assign n2134 = n1224 & ~n2133;
  assign n2135 = n1228 & ~n2134;
  assign n2136 = n1232 & ~n2135;
  assign n2137 = n1236 & ~n2136;
  assign n2138 = n1240 & ~n2137;
  assign n2139 = n1244 & ~n2138;
  assign n2140 = n1248 & ~n2139;
  assign n2141 = n1252 & ~n2140;
  assign n2142 = n1256 & ~n2141;
  assign n2143 = n1260 & ~n2142;
  assign n2144 = n1264 & ~n2143;
  assign n2145 = n1268 & ~n2144;
  assign n2146 = n1272 & ~n2145;
  assign n2147 = n1276 & ~n2146;
  assign n2148 = n1280 & ~n2147;
  assign n2149 = n1284 & ~n2148;
  assign n2150 = n1288 & ~n2149;
  assign n2151 = n1292 & ~n2150;
  assign n2152 = n1296 & ~n2151;
  assign n2153 = n1300 & ~n2152;
  assign n2154 = n1304 & ~n2153;
  assign n2155 = n1308 & ~n2154;
  assign n2156 = n1312 & ~n2155;
  assign n2157 = n1316 & ~n2156;
  assign n2158 = n1320 & ~n2157;
  assign n2159 = n1324 & ~n2158;
  assign n2160 = n1328 & ~n2159;
  assign n2161 = n1332 & ~n2160;
  assign n2162 = n1336 & ~n2161;
  assign n2163 = n1340 & ~n2162;
  assign n2164 = n1344 & ~n2163;
  assign n2165 = n1348 & ~n2164;
  assign n2166 = n1352 & ~n2165;
  assign n2167 = n1356 & ~n2166;
  assign n2168 = n1360 & ~n2167;
  assign n2169 = n1364 & ~n2168;
  assign n2170 = n1368 & ~n2169;
  assign n2171 = n1372 & ~n2170;
  assign n2172 = n1376 & ~n2171;
  assign n2173 = n1380 & ~n2172;
  assign n2174 = n1384 & ~n2173;
  assign n2175 = n1388 & ~n2174;
  assign n2176 = n1392 & ~n2175;
  assign n2177 = n1396 & ~n2176;
  assign n2178 = n1663 & ~n2177;
  assign n2179 = n392 & ~n2178;
  assign n2180 = n396 & ~n2179;
  assign n2181 = n400 & ~n2180;
  assign n2182 = n404 & ~n2181;
  assign n2183 = n408 & ~n2182;
  assign n2184 = pi139  & ~n410;
  assign po11  = ~n2183 & n2184;
  assign n2186 = n419 & ~n754;
  assign n2187 = n424 & ~n2186;
  assign n2188 = n428 & ~n2187;
  assign n2189 = n432 & ~n2188;
  assign n2190 = n436 & ~n2189;
  assign n2191 = n440 & ~n2190;
  assign n2192 = n444 & ~n2191;
  assign n2193 = n448 & ~n2192;
  assign n2194 = n452 & ~n2193;
  assign n2195 = n456 & ~n2194;
  assign n2196 = n460 & ~n2195;
  assign n2197 = n464 & ~n2196;
  assign n2198 = n468 & ~n2197;
  assign n2199 = n472 & ~n2198;
  assign n2200 = n476 & ~n2199;
  assign n2201 = n480 & ~n2200;
  assign n2202 = n484 & ~n2201;
  assign n2203 = n488 & ~n2202;
  assign n2204 = n492 & ~n2203;
  assign n2205 = n496 & ~n2204;
  assign n2206 = n500 & ~n2205;
  assign n2207 = n504 & ~n2206;
  assign n2208 = n508 & ~n2207;
  assign n2209 = n512 & ~n2208;
  assign n2210 = n516 & ~n2209;
  assign n2211 = n520 & ~n2210;
  assign n2212 = n524 & ~n2211;
  assign n2213 = n528 & ~n2212;
  assign n2214 = n532 & ~n2213;
  assign n2215 = n536 & ~n2214;
  assign n2216 = n540 & ~n2215;
  assign n2217 = n544 & ~n2216;
  assign n2218 = n548 & ~n2217;
  assign n2219 = n552 & ~n2218;
  assign n2220 = n556 & ~n2219;
  assign n2221 = n560 & ~n2220;
  assign n2222 = n564 & ~n2221;
  assign n2223 = n568 & ~n2222;
  assign n2224 = n572 & ~n2223;
  assign n2225 = n576 & ~n2224;
  assign n2226 = n580 & ~n2225;
  assign n2227 = n584 & ~n2226;
  assign n2228 = n588 & ~n2227;
  assign n2229 = n592 & ~n2228;
  assign n2230 = n596 & ~n2229;
  assign n2231 = n600 & ~n2230;
  assign n2232 = n604 & ~n2231;
  assign n2233 = n608 & ~n2232;
  assign n2234 = n612 & ~n2233;
  assign n2235 = n616 & ~n2234;
  assign n2236 = n620 & ~n2235;
  assign n2237 = n624 & ~n2236;
  assign n2238 = n628 & ~n2237;
  assign n2239 = n632 & ~n2238;
  assign n2240 = n636 & ~n2239;
  assign n2241 = n640 & ~n2240;
  assign n2242 = n644 & ~n2241;
  assign n2243 = n648 & ~n2242;
  assign n2244 = n652 & ~n2243;
  assign n2245 = n656 & ~n2244;
  assign n2246 = n660 & ~n2245;
  assign n2247 = n664 & ~n2246;
  assign n2248 = n668 & ~n2247;
  assign n2249 = n672 & ~n2248;
  assign n2250 = n676 & ~n2249;
  assign n2251 = n680 & ~n2250;
  assign n2252 = n684 & ~n2251;
  assign n2253 = n688 & ~n2252;
  assign n2254 = n692 & ~n2253;
  assign n2255 = n696 & ~n2254;
  assign n2256 = n700 & ~n2255;
  assign n2257 = n704 & ~n2256;
  assign n2258 = n708 & ~n2257;
  assign n2259 = n712 & ~n2258;
  assign n2260 = n716 & ~n2259;
  assign n2261 = n720 & ~n2260;
  assign n2262 = n1484 & ~n2261;
  assign n2263 = n1486 & ~n2262;
  assign n2264 = n1750 & ~n2263;
  assign n2265 = n731 & ~n2264;
  assign n2266 = n735 & ~n2265;
  assign n2267 = n739 & ~n2266;
  assign n2268 = n743 & ~n2267;
  assign n2269 = n747 & ~n2268;
  assign n2270 = pi140  & ~n749;
  assign po12  = ~n2269 & n2270;
  assign n2272 = n758 & ~n1091;
  assign n2273 = n763 & ~n2272;
  assign n2274 = n767 & ~n2273;
  assign n2275 = n771 & ~n2274;
  assign n2276 = n775 & ~n2275;
  assign n2277 = n779 & ~n2276;
  assign n2278 = n783 & ~n2277;
  assign n2279 = n787 & ~n2278;
  assign n2280 = n791 & ~n2279;
  assign n2281 = n795 & ~n2280;
  assign n2282 = n799 & ~n2281;
  assign n2283 = n803 & ~n2282;
  assign n2284 = n807 & ~n2283;
  assign n2285 = n811 & ~n2284;
  assign n2286 = n815 & ~n2285;
  assign n2287 = n819 & ~n2286;
  assign n2288 = n823 & ~n2287;
  assign n2289 = n827 & ~n2288;
  assign n2290 = n831 & ~n2289;
  assign n2291 = n835 & ~n2290;
  assign n2292 = n839 & ~n2291;
  assign n2293 = n843 & ~n2292;
  assign n2294 = n847 & ~n2293;
  assign n2295 = n851 & ~n2294;
  assign n2296 = n855 & ~n2295;
  assign n2297 = n859 & ~n2296;
  assign n2298 = n863 & ~n2297;
  assign n2299 = n867 & ~n2298;
  assign n2300 = n871 & ~n2299;
  assign n2301 = n875 & ~n2300;
  assign n2302 = n879 & ~n2301;
  assign n2303 = n883 & ~n2302;
  assign n2304 = n887 & ~n2303;
  assign n2305 = n891 & ~n2304;
  assign n2306 = n895 & ~n2305;
  assign n2307 = n899 & ~n2306;
  assign n2308 = n903 & ~n2307;
  assign n2309 = n907 & ~n2308;
  assign n2310 = n911 & ~n2309;
  assign n2311 = n915 & ~n2310;
  assign n2312 = n919 & ~n2311;
  assign n2313 = n923 & ~n2312;
  assign n2314 = n927 & ~n2313;
  assign n2315 = n931 & ~n2314;
  assign n2316 = n935 & ~n2315;
  assign n2317 = n939 & ~n2316;
  assign n2318 = n943 & ~n2317;
  assign n2319 = n947 & ~n2318;
  assign n2320 = n951 & ~n2319;
  assign n2321 = n955 & ~n2320;
  assign n2322 = n959 & ~n2321;
  assign n2323 = n963 & ~n2322;
  assign n2324 = n967 & ~n2323;
  assign n2325 = n971 & ~n2324;
  assign n2326 = n975 & ~n2325;
  assign n2327 = n979 & ~n2326;
  assign n2328 = n983 & ~n2327;
  assign n2329 = n987 & ~n2328;
  assign n2330 = n991 & ~n2329;
  assign n2331 = n995 & ~n2330;
  assign n2332 = n999 & ~n2331;
  assign n2333 = n1003 & ~n2332;
  assign n2334 = n1007 & ~n2333;
  assign n2335 = n1011 & ~n2334;
  assign n2336 = n1015 & ~n2335;
  assign n2337 = n1019 & ~n2336;
  assign n2338 = n1023 & ~n2337;
  assign n2339 = n1027 & ~n2338;
  assign n2340 = n1031 & ~n2339;
  assign n2341 = n1035 & ~n2340;
  assign n2342 = n1039 & ~n2341;
  assign n2343 = n1043 & ~n2342;
  assign n2344 = n1047 & ~n2343;
  assign n2345 = n1051 & ~n2344;
  assign n2346 = n1055 & ~n2345;
  assign n2347 = n1059 & ~n2346;
  assign n2348 = n1574 & ~n2347;
  assign n2349 = n1576 & ~n2348;
  assign n2350 = n1837 & ~n2349;
  assign n2351 = n1068 & ~n2350;
  assign n2352 = n1072 & ~n2351;
  assign n2353 = n1076 & ~n2352;
  assign n2354 = n1080 & ~n2353;
  assign n2355 = n1084 & ~n2354;
  assign n2356 = pi141  & ~n1086;
  assign po13  = ~n2355 & n2356;
  assign n2358 = ~n423 & n1095;
  assign n2359 = n1100 & ~n2358;
  assign n2360 = n1104 & ~n2359;
  assign n2361 = n1108 & ~n2360;
  assign n2362 = n1112 & ~n2361;
  assign n2363 = n1116 & ~n2362;
  assign n2364 = n1120 & ~n2363;
  assign n2365 = n1124 & ~n2364;
  assign n2366 = n1128 & ~n2365;
  assign n2367 = n1132 & ~n2366;
  assign n2368 = n1136 & ~n2367;
  assign n2369 = n1140 & ~n2368;
  assign n2370 = n1144 & ~n2369;
  assign n2371 = n1148 & ~n2370;
  assign n2372 = n1152 & ~n2371;
  assign n2373 = n1156 & ~n2372;
  assign n2374 = n1160 & ~n2373;
  assign n2375 = n1164 & ~n2374;
  assign n2376 = n1168 & ~n2375;
  assign n2377 = n1172 & ~n2376;
  assign n2378 = n1176 & ~n2377;
  assign n2379 = n1180 & ~n2378;
  assign n2380 = n1184 & ~n2379;
  assign n2381 = n1188 & ~n2380;
  assign n2382 = n1192 & ~n2381;
  assign n2383 = n1196 & ~n2382;
  assign n2384 = n1200 & ~n2383;
  assign n2385 = n1204 & ~n2384;
  assign n2386 = n1208 & ~n2385;
  assign n2387 = n1212 & ~n2386;
  assign n2388 = n1216 & ~n2387;
  assign n2389 = n1220 & ~n2388;
  assign n2390 = n1224 & ~n2389;
  assign n2391 = n1228 & ~n2390;
  assign n2392 = n1232 & ~n2391;
  assign n2393 = n1236 & ~n2392;
  assign n2394 = n1240 & ~n2393;
  assign n2395 = n1244 & ~n2394;
  assign n2396 = n1248 & ~n2395;
  assign n2397 = n1252 & ~n2396;
  assign n2398 = n1256 & ~n2397;
  assign n2399 = n1260 & ~n2398;
  assign n2400 = n1264 & ~n2399;
  assign n2401 = n1268 & ~n2400;
  assign n2402 = n1272 & ~n2401;
  assign n2403 = n1276 & ~n2402;
  assign n2404 = n1280 & ~n2403;
  assign n2405 = n1284 & ~n2404;
  assign n2406 = n1288 & ~n2405;
  assign n2407 = n1292 & ~n2406;
  assign n2408 = n1296 & ~n2407;
  assign n2409 = n1300 & ~n2408;
  assign n2410 = n1304 & ~n2409;
  assign n2411 = n1308 & ~n2410;
  assign n2412 = n1312 & ~n2411;
  assign n2413 = n1316 & ~n2412;
  assign n2414 = n1320 & ~n2413;
  assign n2415 = n1324 & ~n2414;
  assign n2416 = n1328 & ~n2415;
  assign n2417 = n1332 & ~n2416;
  assign n2418 = n1336 & ~n2417;
  assign n2419 = n1340 & ~n2418;
  assign n2420 = n1344 & ~n2419;
  assign n2421 = n1348 & ~n2420;
  assign n2422 = n1352 & ~n2421;
  assign n2423 = n1356 & ~n2422;
  assign n2424 = n1360 & ~n2423;
  assign n2425 = n1364 & ~n2424;
  assign n2426 = n1368 & ~n2425;
  assign n2427 = n1372 & ~n2426;
  assign n2428 = n1376 & ~n2427;
  assign n2429 = n1380 & ~n2428;
  assign n2430 = n1384 & ~n2429;
  assign n2431 = n1388 & ~n2430;
  assign n2432 = n1392 & ~n2431;
  assign n2433 = n1396 & ~n2432;
  assign n2434 = n1663 & ~n2433;
  assign n2435 = n392 & ~n2434;
  assign n2436 = n396 & ~n2435;
  assign n2437 = n400 & ~n2436;
  assign n2438 = n404 & ~n2437;
  assign n2439 = n408 & ~n2438;
  assign n2440 = n412 & ~n2439;
  assign n2441 = n416 & ~n2440;
  assign n2442 = pi142  & ~n418;
  assign po14  = ~n2441 & n2442;
  assign n2444 = n427 & ~n762;
  assign n2445 = n432 & ~n2444;
  assign n2446 = n436 & ~n2445;
  assign n2447 = n440 & ~n2446;
  assign n2448 = n444 & ~n2447;
  assign n2449 = n448 & ~n2448;
  assign n2450 = n452 & ~n2449;
  assign n2451 = n456 & ~n2450;
  assign n2452 = n460 & ~n2451;
  assign n2453 = n464 & ~n2452;
  assign n2454 = n468 & ~n2453;
  assign n2455 = n472 & ~n2454;
  assign n2456 = n476 & ~n2455;
  assign n2457 = n480 & ~n2456;
  assign n2458 = n484 & ~n2457;
  assign n2459 = n488 & ~n2458;
  assign n2460 = n492 & ~n2459;
  assign n2461 = n496 & ~n2460;
  assign n2462 = n500 & ~n2461;
  assign n2463 = n504 & ~n2462;
  assign n2464 = n508 & ~n2463;
  assign n2465 = n512 & ~n2464;
  assign n2466 = n516 & ~n2465;
  assign n2467 = n520 & ~n2466;
  assign n2468 = n524 & ~n2467;
  assign n2469 = n528 & ~n2468;
  assign n2470 = n532 & ~n2469;
  assign n2471 = n536 & ~n2470;
  assign n2472 = n540 & ~n2471;
  assign n2473 = n544 & ~n2472;
  assign n2474 = n548 & ~n2473;
  assign n2475 = n552 & ~n2474;
  assign n2476 = n556 & ~n2475;
  assign n2477 = n560 & ~n2476;
  assign n2478 = n564 & ~n2477;
  assign n2479 = n568 & ~n2478;
  assign n2480 = n572 & ~n2479;
  assign n2481 = n576 & ~n2480;
  assign n2482 = n580 & ~n2481;
  assign n2483 = n584 & ~n2482;
  assign n2484 = n588 & ~n2483;
  assign n2485 = n592 & ~n2484;
  assign n2486 = n596 & ~n2485;
  assign n2487 = n600 & ~n2486;
  assign n2488 = n604 & ~n2487;
  assign n2489 = n608 & ~n2488;
  assign n2490 = n612 & ~n2489;
  assign n2491 = n616 & ~n2490;
  assign n2492 = n620 & ~n2491;
  assign n2493 = n624 & ~n2492;
  assign n2494 = n628 & ~n2493;
  assign n2495 = n632 & ~n2494;
  assign n2496 = n636 & ~n2495;
  assign n2497 = n640 & ~n2496;
  assign n2498 = n644 & ~n2497;
  assign n2499 = n648 & ~n2498;
  assign n2500 = n652 & ~n2499;
  assign n2501 = n656 & ~n2500;
  assign n2502 = n660 & ~n2501;
  assign n2503 = n664 & ~n2502;
  assign n2504 = n668 & ~n2503;
  assign n2505 = n672 & ~n2504;
  assign n2506 = n676 & ~n2505;
  assign n2507 = n680 & ~n2506;
  assign n2508 = n684 & ~n2507;
  assign n2509 = n688 & ~n2508;
  assign n2510 = n692 & ~n2509;
  assign n2511 = n696 & ~n2510;
  assign n2512 = n700 & ~n2511;
  assign n2513 = n704 & ~n2512;
  assign n2514 = n708 & ~n2513;
  assign n2515 = n712 & ~n2514;
  assign n2516 = n716 & ~n2515;
  assign n2517 = n720 & ~n2516;
  assign n2518 = n1484 & ~n2517;
  assign n2519 = n1486 & ~n2518;
  assign n2520 = n1750 & ~n2519;
  assign n2521 = n731 & ~n2520;
  assign n2522 = n735 & ~n2521;
  assign n2523 = n739 & ~n2522;
  assign n2524 = n743 & ~n2523;
  assign n2525 = n747 & ~n2524;
  assign n2526 = n751 & ~n2525;
  assign n2527 = n755 & ~n2526;
  assign n2528 = pi143  & ~n757;
  assign po15  = ~n2527 & n2528;
  assign n2530 = n766 & ~n1099;
  assign n2531 = n771 & ~n2530;
  assign n2532 = n775 & ~n2531;
  assign n2533 = n779 & ~n2532;
  assign n2534 = n783 & ~n2533;
  assign n2535 = n787 & ~n2534;
  assign n2536 = n791 & ~n2535;
  assign n2537 = n795 & ~n2536;
  assign n2538 = n799 & ~n2537;
  assign n2539 = n803 & ~n2538;
  assign n2540 = n807 & ~n2539;
  assign n2541 = n811 & ~n2540;
  assign n2542 = n815 & ~n2541;
  assign n2543 = n819 & ~n2542;
  assign n2544 = n823 & ~n2543;
  assign n2545 = n827 & ~n2544;
  assign n2546 = n831 & ~n2545;
  assign n2547 = n835 & ~n2546;
  assign n2548 = n839 & ~n2547;
  assign n2549 = n843 & ~n2548;
  assign n2550 = n847 & ~n2549;
  assign n2551 = n851 & ~n2550;
  assign n2552 = n855 & ~n2551;
  assign n2553 = n859 & ~n2552;
  assign n2554 = n863 & ~n2553;
  assign n2555 = n867 & ~n2554;
  assign n2556 = n871 & ~n2555;
  assign n2557 = n875 & ~n2556;
  assign n2558 = n879 & ~n2557;
  assign n2559 = n883 & ~n2558;
  assign n2560 = n887 & ~n2559;
  assign n2561 = n891 & ~n2560;
  assign n2562 = n895 & ~n2561;
  assign n2563 = n899 & ~n2562;
  assign n2564 = n903 & ~n2563;
  assign n2565 = n907 & ~n2564;
  assign n2566 = n911 & ~n2565;
  assign n2567 = n915 & ~n2566;
  assign n2568 = n919 & ~n2567;
  assign n2569 = n923 & ~n2568;
  assign n2570 = n927 & ~n2569;
  assign n2571 = n931 & ~n2570;
  assign n2572 = n935 & ~n2571;
  assign n2573 = n939 & ~n2572;
  assign n2574 = n943 & ~n2573;
  assign n2575 = n947 & ~n2574;
  assign n2576 = n951 & ~n2575;
  assign n2577 = n955 & ~n2576;
  assign n2578 = n959 & ~n2577;
  assign n2579 = n963 & ~n2578;
  assign n2580 = n967 & ~n2579;
  assign n2581 = n971 & ~n2580;
  assign n2582 = n975 & ~n2581;
  assign n2583 = n979 & ~n2582;
  assign n2584 = n983 & ~n2583;
  assign n2585 = n987 & ~n2584;
  assign n2586 = n991 & ~n2585;
  assign n2587 = n995 & ~n2586;
  assign n2588 = n999 & ~n2587;
  assign n2589 = n1003 & ~n2588;
  assign n2590 = n1007 & ~n2589;
  assign n2591 = n1011 & ~n2590;
  assign n2592 = n1015 & ~n2591;
  assign n2593 = n1019 & ~n2592;
  assign n2594 = n1023 & ~n2593;
  assign n2595 = n1027 & ~n2594;
  assign n2596 = n1031 & ~n2595;
  assign n2597 = n1035 & ~n2596;
  assign n2598 = n1039 & ~n2597;
  assign n2599 = n1043 & ~n2598;
  assign n2600 = n1047 & ~n2599;
  assign n2601 = n1051 & ~n2600;
  assign n2602 = n1055 & ~n2601;
  assign n2603 = n1059 & ~n2602;
  assign n2604 = n1574 & ~n2603;
  assign n2605 = n1576 & ~n2604;
  assign n2606 = n1837 & ~n2605;
  assign n2607 = n1068 & ~n2606;
  assign n2608 = n1072 & ~n2607;
  assign n2609 = n1076 & ~n2608;
  assign n2610 = n1080 & ~n2609;
  assign n2611 = n1084 & ~n2610;
  assign n2612 = n1088 & ~n2611;
  assign n2613 = n1092 & ~n2612;
  assign n2614 = pi144  & ~n1094;
  assign po16  = ~n2613 & n2614;
  assign n2616 = ~n431 & n1103;
  assign n2617 = n1108 & ~n2616;
  assign n2618 = n1112 & ~n2617;
  assign n2619 = n1116 & ~n2618;
  assign n2620 = n1120 & ~n2619;
  assign n2621 = n1124 & ~n2620;
  assign n2622 = n1128 & ~n2621;
  assign n2623 = n1132 & ~n2622;
  assign n2624 = n1136 & ~n2623;
  assign n2625 = n1140 & ~n2624;
  assign n2626 = n1144 & ~n2625;
  assign n2627 = n1148 & ~n2626;
  assign n2628 = n1152 & ~n2627;
  assign n2629 = n1156 & ~n2628;
  assign n2630 = n1160 & ~n2629;
  assign n2631 = n1164 & ~n2630;
  assign n2632 = n1168 & ~n2631;
  assign n2633 = n1172 & ~n2632;
  assign n2634 = n1176 & ~n2633;
  assign n2635 = n1180 & ~n2634;
  assign n2636 = n1184 & ~n2635;
  assign n2637 = n1188 & ~n2636;
  assign n2638 = n1192 & ~n2637;
  assign n2639 = n1196 & ~n2638;
  assign n2640 = n1200 & ~n2639;
  assign n2641 = n1204 & ~n2640;
  assign n2642 = n1208 & ~n2641;
  assign n2643 = n1212 & ~n2642;
  assign n2644 = n1216 & ~n2643;
  assign n2645 = n1220 & ~n2644;
  assign n2646 = n1224 & ~n2645;
  assign n2647 = n1228 & ~n2646;
  assign n2648 = n1232 & ~n2647;
  assign n2649 = n1236 & ~n2648;
  assign n2650 = n1240 & ~n2649;
  assign n2651 = n1244 & ~n2650;
  assign n2652 = n1248 & ~n2651;
  assign n2653 = n1252 & ~n2652;
  assign n2654 = n1256 & ~n2653;
  assign n2655 = n1260 & ~n2654;
  assign n2656 = n1264 & ~n2655;
  assign n2657 = n1268 & ~n2656;
  assign n2658 = n1272 & ~n2657;
  assign n2659 = n1276 & ~n2658;
  assign n2660 = n1280 & ~n2659;
  assign n2661 = n1284 & ~n2660;
  assign n2662 = n1288 & ~n2661;
  assign n2663 = n1292 & ~n2662;
  assign n2664 = n1296 & ~n2663;
  assign n2665 = n1300 & ~n2664;
  assign n2666 = n1304 & ~n2665;
  assign n2667 = n1308 & ~n2666;
  assign n2668 = n1312 & ~n2667;
  assign n2669 = n1316 & ~n2668;
  assign n2670 = n1320 & ~n2669;
  assign n2671 = n1324 & ~n2670;
  assign n2672 = n1328 & ~n2671;
  assign n2673 = n1332 & ~n2672;
  assign n2674 = n1336 & ~n2673;
  assign n2675 = n1340 & ~n2674;
  assign n2676 = n1344 & ~n2675;
  assign n2677 = n1348 & ~n2676;
  assign n2678 = n1352 & ~n2677;
  assign n2679 = n1356 & ~n2678;
  assign n2680 = n1360 & ~n2679;
  assign n2681 = n1364 & ~n2680;
  assign n2682 = n1368 & ~n2681;
  assign n2683 = n1372 & ~n2682;
  assign n2684 = n1376 & ~n2683;
  assign n2685 = n1380 & ~n2684;
  assign n2686 = n1384 & ~n2685;
  assign n2687 = n1388 & ~n2686;
  assign n2688 = n1392 & ~n2687;
  assign n2689 = n1396 & ~n2688;
  assign n2690 = n1663 & ~n2689;
  assign n2691 = n392 & ~n2690;
  assign n2692 = n396 & ~n2691;
  assign n2693 = n400 & ~n2692;
  assign n2694 = n404 & ~n2693;
  assign n2695 = n408 & ~n2694;
  assign n2696 = n412 & ~n2695;
  assign n2697 = n416 & ~n2696;
  assign n2698 = n420 & ~n2697;
  assign n2699 = n424 & ~n2698;
  assign n2700 = pi145  & ~n426;
  assign po17  = ~n2699 & n2700;
  assign n2702 = n435 & ~n770;
  assign n2703 = n440 & ~n2702;
  assign n2704 = n444 & ~n2703;
  assign n2705 = n448 & ~n2704;
  assign n2706 = n452 & ~n2705;
  assign n2707 = n456 & ~n2706;
  assign n2708 = n460 & ~n2707;
  assign n2709 = n464 & ~n2708;
  assign n2710 = n468 & ~n2709;
  assign n2711 = n472 & ~n2710;
  assign n2712 = n476 & ~n2711;
  assign n2713 = n480 & ~n2712;
  assign n2714 = n484 & ~n2713;
  assign n2715 = n488 & ~n2714;
  assign n2716 = n492 & ~n2715;
  assign n2717 = n496 & ~n2716;
  assign n2718 = n500 & ~n2717;
  assign n2719 = n504 & ~n2718;
  assign n2720 = n508 & ~n2719;
  assign n2721 = n512 & ~n2720;
  assign n2722 = n516 & ~n2721;
  assign n2723 = n520 & ~n2722;
  assign n2724 = n524 & ~n2723;
  assign n2725 = n528 & ~n2724;
  assign n2726 = n532 & ~n2725;
  assign n2727 = n536 & ~n2726;
  assign n2728 = n540 & ~n2727;
  assign n2729 = n544 & ~n2728;
  assign n2730 = n548 & ~n2729;
  assign n2731 = n552 & ~n2730;
  assign n2732 = n556 & ~n2731;
  assign n2733 = n560 & ~n2732;
  assign n2734 = n564 & ~n2733;
  assign n2735 = n568 & ~n2734;
  assign n2736 = n572 & ~n2735;
  assign n2737 = n576 & ~n2736;
  assign n2738 = n580 & ~n2737;
  assign n2739 = n584 & ~n2738;
  assign n2740 = n588 & ~n2739;
  assign n2741 = n592 & ~n2740;
  assign n2742 = n596 & ~n2741;
  assign n2743 = n600 & ~n2742;
  assign n2744 = n604 & ~n2743;
  assign n2745 = n608 & ~n2744;
  assign n2746 = n612 & ~n2745;
  assign n2747 = n616 & ~n2746;
  assign n2748 = n620 & ~n2747;
  assign n2749 = n624 & ~n2748;
  assign n2750 = n628 & ~n2749;
  assign n2751 = n632 & ~n2750;
  assign n2752 = n636 & ~n2751;
  assign n2753 = n640 & ~n2752;
  assign n2754 = n644 & ~n2753;
  assign n2755 = n648 & ~n2754;
  assign n2756 = n652 & ~n2755;
  assign n2757 = n656 & ~n2756;
  assign n2758 = n660 & ~n2757;
  assign n2759 = n664 & ~n2758;
  assign n2760 = n668 & ~n2759;
  assign n2761 = n672 & ~n2760;
  assign n2762 = n676 & ~n2761;
  assign n2763 = n680 & ~n2762;
  assign n2764 = n684 & ~n2763;
  assign n2765 = n688 & ~n2764;
  assign n2766 = n692 & ~n2765;
  assign n2767 = n696 & ~n2766;
  assign n2768 = n700 & ~n2767;
  assign n2769 = n704 & ~n2768;
  assign n2770 = n708 & ~n2769;
  assign n2771 = n712 & ~n2770;
  assign n2772 = n716 & ~n2771;
  assign n2773 = n720 & ~n2772;
  assign n2774 = n1484 & ~n2773;
  assign n2775 = n1486 & ~n2774;
  assign n2776 = n1750 & ~n2775;
  assign n2777 = n731 & ~n2776;
  assign n2778 = n735 & ~n2777;
  assign n2779 = n739 & ~n2778;
  assign n2780 = n743 & ~n2779;
  assign n2781 = n747 & ~n2780;
  assign n2782 = n751 & ~n2781;
  assign n2783 = n755 & ~n2782;
  assign n2784 = n759 & ~n2783;
  assign n2785 = n763 & ~n2784;
  assign n2786 = pi146  & ~n765;
  assign po18  = ~n2785 & n2786;
  assign n2788 = n774 & ~n1107;
  assign n2789 = n779 & ~n2788;
  assign n2790 = n783 & ~n2789;
  assign n2791 = n787 & ~n2790;
  assign n2792 = n791 & ~n2791;
  assign n2793 = n795 & ~n2792;
  assign n2794 = n799 & ~n2793;
  assign n2795 = n803 & ~n2794;
  assign n2796 = n807 & ~n2795;
  assign n2797 = n811 & ~n2796;
  assign n2798 = n815 & ~n2797;
  assign n2799 = n819 & ~n2798;
  assign n2800 = n823 & ~n2799;
  assign n2801 = n827 & ~n2800;
  assign n2802 = n831 & ~n2801;
  assign n2803 = n835 & ~n2802;
  assign n2804 = n839 & ~n2803;
  assign n2805 = n843 & ~n2804;
  assign n2806 = n847 & ~n2805;
  assign n2807 = n851 & ~n2806;
  assign n2808 = n855 & ~n2807;
  assign n2809 = n859 & ~n2808;
  assign n2810 = n863 & ~n2809;
  assign n2811 = n867 & ~n2810;
  assign n2812 = n871 & ~n2811;
  assign n2813 = n875 & ~n2812;
  assign n2814 = n879 & ~n2813;
  assign n2815 = n883 & ~n2814;
  assign n2816 = n887 & ~n2815;
  assign n2817 = n891 & ~n2816;
  assign n2818 = n895 & ~n2817;
  assign n2819 = n899 & ~n2818;
  assign n2820 = n903 & ~n2819;
  assign n2821 = n907 & ~n2820;
  assign n2822 = n911 & ~n2821;
  assign n2823 = n915 & ~n2822;
  assign n2824 = n919 & ~n2823;
  assign n2825 = n923 & ~n2824;
  assign n2826 = n927 & ~n2825;
  assign n2827 = n931 & ~n2826;
  assign n2828 = n935 & ~n2827;
  assign n2829 = n939 & ~n2828;
  assign n2830 = n943 & ~n2829;
  assign n2831 = n947 & ~n2830;
  assign n2832 = n951 & ~n2831;
  assign n2833 = n955 & ~n2832;
  assign n2834 = n959 & ~n2833;
  assign n2835 = n963 & ~n2834;
  assign n2836 = n967 & ~n2835;
  assign n2837 = n971 & ~n2836;
  assign n2838 = n975 & ~n2837;
  assign n2839 = n979 & ~n2838;
  assign n2840 = n983 & ~n2839;
  assign n2841 = n987 & ~n2840;
  assign n2842 = n991 & ~n2841;
  assign n2843 = n995 & ~n2842;
  assign n2844 = n999 & ~n2843;
  assign n2845 = n1003 & ~n2844;
  assign n2846 = n1007 & ~n2845;
  assign n2847 = n1011 & ~n2846;
  assign n2848 = n1015 & ~n2847;
  assign n2849 = n1019 & ~n2848;
  assign n2850 = n1023 & ~n2849;
  assign n2851 = n1027 & ~n2850;
  assign n2852 = n1031 & ~n2851;
  assign n2853 = n1035 & ~n2852;
  assign n2854 = n1039 & ~n2853;
  assign n2855 = n1043 & ~n2854;
  assign n2856 = n1047 & ~n2855;
  assign n2857 = n1051 & ~n2856;
  assign n2858 = n1055 & ~n2857;
  assign n2859 = n1059 & ~n2858;
  assign n2860 = n1574 & ~n2859;
  assign n2861 = n1576 & ~n2860;
  assign n2862 = n1837 & ~n2861;
  assign n2863 = n1068 & ~n2862;
  assign n2864 = n1072 & ~n2863;
  assign n2865 = n1076 & ~n2864;
  assign n2866 = n1080 & ~n2865;
  assign n2867 = n1084 & ~n2866;
  assign n2868 = n1088 & ~n2867;
  assign n2869 = n1092 & ~n2868;
  assign n2870 = n1096 & ~n2869;
  assign n2871 = n1100 & ~n2870;
  assign n2872 = pi147  & ~n1102;
  assign po19  = ~n2871 & n2872;
  assign n2874 = ~n439 & n1111;
  assign n2875 = n1116 & ~n2874;
  assign n2876 = n1120 & ~n2875;
  assign n2877 = n1124 & ~n2876;
  assign n2878 = n1128 & ~n2877;
  assign n2879 = n1132 & ~n2878;
  assign n2880 = n1136 & ~n2879;
  assign n2881 = n1140 & ~n2880;
  assign n2882 = n1144 & ~n2881;
  assign n2883 = n1148 & ~n2882;
  assign n2884 = n1152 & ~n2883;
  assign n2885 = n1156 & ~n2884;
  assign n2886 = n1160 & ~n2885;
  assign n2887 = n1164 & ~n2886;
  assign n2888 = n1168 & ~n2887;
  assign n2889 = n1172 & ~n2888;
  assign n2890 = n1176 & ~n2889;
  assign n2891 = n1180 & ~n2890;
  assign n2892 = n1184 & ~n2891;
  assign n2893 = n1188 & ~n2892;
  assign n2894 = n1192 & ~n2893;
  assign n2895 = n1196 & ~n2894;
  assign n2896 = n1200 & ~n2895;
  assign n2897 = n1204 & ~n2896;
  assign n2898 = n1208 & ~n2897;
  assign n2899 = n1212 & ~n2898;
  assign n2900 = n1216 & ~n2899;
  assign n2901 = n1220 & ~n2900;
  assign n2902 = n1224 & ~n2901;
  assign n2903 = n1228 & ~n2902;
  assign n2904 = n1232 & ~n2903;
  assign n2905 = n1236 & ~n2904;
  assign n2906 = n1240 & ~n2905;
  assign n2907 = n1244 & ~n2906;
  assign n2908 = n1248 & ~n2907;
  assign n2909 = n1252 & ~n2908;
  assign n2910 = n1256 & ~n2909;
  assign n2911 = n1260 & ~n2910;
  assign n2912 = n1264 & ~n2911;
  assign n2913 = n1268 & ~n2912;
  assign n2914 = n1272 & ~n2913;
  assign n2915 = n1276 & ~n2914;
  assign n2916 = n1280 & ~n2915;
  assign n2917 = n1284 & ~n2916;
  assign n2918 = n1288 & ~n2917;
  assign n2919 = n1292 & ~n2918;
  assign n2920 = n1296 & ~n2919;
  assign n2921 = n1300 & ~n2920;
  assign n2922 = n1304 & ~n2921;
  assign n2923 = n1308 & ~n2922;
  assign n2924 = n1312 & ~n2923;
  assign n2925 = n1316 & ~n2924;
  assign n2926 = n1320 & ~n2925;
  assign n2927 = n1324 & ~n2926;
  assign n2928 = n1328 & ~n2927;
  assign n2929 = n1332 & ~n2928;
  assign n2930 = n1336 & ~n2929;
  assign n2931 = n1340 & ~n2930;
  assign n2932 = n1344 & ~n2931;
  assign n2933 = n1348 & ~n2932;
  assign n2934 = n1352 & ~n2933;
  assign n2935 = n1356 & ~n2934;
  assign n2936 = n1360 & ~n2935;
  assign n2937 = n1364 & ~n2936;
  assign n2938 = n1368 & ~n2937;
  assign n2939 = n1372 & ~n2938;
  assign n2940 = n1376 & ~n2939;
  assign n2941 = n1380 & ~n2940;
  assign n2942 = n1384 & ~n2941;
  assign n2943 = n1388 & ~n2942;
  assign n2944 = n1392 & ~n2943;
  assign n2945 = n1396 & ~n2944;
  assign n2946 = n1663 & ~n2945;
  assign n2947 = n392 & ~n2946;
  assign n2948 = n396 & ~n2947;
  assign n2949 = n400 & ~n2948;
  assign n2950 = n404 & ~n2949;
  assign n2951 = n408 & ~n2950;
  assign n2952 = n412 & ~n2951;
  assign n2953 = n416 & ~n2952;
  assign n2954 = n420 & ~n2953;
  assign n2955 = n424 & ~n2954;
  assign n2956 = n428 & ~n2955;
  assign n2957 = n432 & ~n2956;
  assign n2958 = pi148  & ~n434;
  assign po20  = ~n2957 & n2958;
  assign n2960 = n443 & ~n778;
  assign n2961 = n448 & ~n2960;
  assign n2962 = n452 & ~n2961;
  assign n2963 = n456 & ~n2962;
  assign n2964 = n460 & ~n2963;
  assign n2965 = n464 & ~n2964;
  assign n2966 = n468 & ~n2965;
  assign n2967 = n472 & ~n2966;
  assign n2968 = n476 & ~n2967;
  assign n2969 = n480 & ~n2968;
  assign n2970 = n484 & ~n2969;
  assign n2971 = n488 & ~n2970;
  assign n2972 = n492 & ~n2971;
  assign n2973 = n496 & ~n2972;
  assign n2974 = n500 & ~n2973;
  assign n2975 = n504 & ~n2974;
  assign n2976 = n508 & ~n2975;
  assign n2977 = n512 & ~n2976;
  assign n2978 = n516 & ~n2977;
  assign n2979 = n520 & ~n2978;
  assign n2980 = n524 & ~n2979;
  assign n2981 = n528 & ~n2980;
  assign n2982 = n532 & ~n2981;
  assign n2983 = n536 & ~n2982;
  assign n2984 = n540 & ~n2983;
  assign n2985 = n544 & ~n2984;
  assign n2986 = n548 & ~n2985;
  assign n2987 = n552 & ~n2986;
  assign n2988 = n556 & ~n2987;
  assign n2989 = n560 & ~n2988;
  assign n2990 = n564 & ~n2989;
  assign n2991 = n568 & ~n2990;
  assign n2992 = n572 & ~n2991;
  assign n2993 = n576 & ~n2992;
  assign n2994 = n580 & ~n2993;
  assign n2995 = n584 & ~n2994;
  assign n2996 = n588 & ~n2995;
  assign n2997 = n592 & ~n2996;
  assign n2998 = n596 & ~n2997;
  assign n2999 = n600 & ~n2998;
  assign n3000 = n604 & ~n2999;
  assign n3001 = n608 & ~n3000;
  assign n3002 = n612 & ~n3001;
  assign n3003 = n616 & ~n3002;
  assign n3004 = n620 & ~n3003;
  assign n3005 = n624 & ~n3004;
  assign n3006 = n628 & ~n3005;
  assign n3007 = n632 & ~n3006;
  assign n3008 = n636 & ~n3007;
  assign n3009 = n640 & ~n3008;
  assign n3010 = n644 & ~n3009;
  assign n3011 = n648 & ~n3010;
  assign n3012 = n652 & ~n3011;
  assign n3013 = n656 & ~n3012;
  assign n3014 = n660 & ~n3013;
  assign n3015 = n664 & ~n3014;
  assign n3016 = n668 & ~n3015;
  assign n3017 = n672 & ~n3016;
  assign n3018 = n676 & ~n3017;
  assign n3019 = n680 & ~n3018;
  assign n3020 = n684 & ~n3019;
  assign n3021 = n688 & ~n3020;
  assign n3022 = n692 & ~n3021;
  assign n3023 = n696 & ~n3022;
  assign n3024 = n700 & ~n3023;
  assign n3025 = n704 & ~n3024;
  assign n3026 = n708 & ~n3025;
  assign n3027 = n712 & ~n3026;
  assign n3028 = n716 & ~n3027;
  assign n3029 = n720 & ~n3028;
  assign n3030 = n1484 & ~n3029;
  assign n3031 = n1486 & ~n3030;
  assign n3032 = n1750 & ~n3031;
  assign n3033 = n731 & ~n3032;
  assign n3034 = n735 & ~n3033;
  assign n3035 = n739 & ~n3034;
  assign n3036 = n743 & ~n3035;
  assign n3037 = n747 & ~n3036;
  assign n3038 = n751 & ~n3037;
  assign n3039 = n755 & ~n3038;
  assign n3040 = n759 & ~n3039;
  assign n3041 = n763 & ~n3040;
  assign n3042 = n767 & ~n3041;
  assign n3043 = n771 & ~n3042;
  assign n3044 = pi149  & ~n773;
  assign po21  = ~n3043 & n3044;
  assign n3046 = n782 & ~n1115;
  assign n3047 = n787 & ~n3046;
  assign n3048 = n791 & ~n3047;
  assign n3049 = n795 & ~n3048;
  assign n3050 = n799 & ~n3049;
  assign n3051 = n803 & ~n3050;
  assign n3052 = n807 & ~n3051;
  assign n3053 = n811 & ~n3052;
  assign n3054 = n815 & ~n3053;
  assign n3055 = n819 & ~n3054;
  assign n3056 = n823 & ~n3055;
  assign n3057 = n827 & ~n3056;
  assign n3058 = n831 & ~n3057;
  assign n3059 = n835 & ~n3058;
  assign n3060 = n839 & ~n3059;
  assign n3061 = n843 & ~n3060;
  assign n3062 = n847 & ~n3061;
  assign n3063 = n851 & ~n3062;
  assign n3064 = n855 & ~n3063;
  assign n3065 = n859 & ~n3064;
  assign n3066 = n863 & ~n3065;
  assign n3067 = n867 & ~n3066;
  assign n3068 = n871 & ~n3067;
  assign n3069 = n875 & ~n3068;
  assign n3070 = n879 & ~n3069;
  assign n3071 = n883 & ~n3070;
  assign n3072 = n887 & ~n3071;
  assign n3073 = n891 & ~n3072;
  assign n3074 = n895 & ~n3073;
  assign n3075 = n899 & ~n3074;
  assign n3076 = n903 & ~n3075;
  assign n3077 = n907 & ~n3076;
  assign n3078 = n911 & ~n3077;
  assign n3079 = n915 & ~n3078;
  assign n3080 = n919 & ~n3079;
  assign n3081 = n923 & ~n3080;
  assign n3082 = n927 & ~n3081;
  assign n3083 = n931 & ~n3082;
  assign n3084 = n935 & ~n3083;
  assign n3085 = n939 & ~n3084;
  assign n3086 = n943 & ~n3085;
  assign n3087 = n947 & ~n3086;
  assign n3088 = n951 & ~n3087;
  assign n3089 = n955 & ~n3088;
  assign n3090 = n959 & ~n3089;
  assign n3091 = n963 & ~n3090;
  assign n3092 = n967 & ~n3091;
  assign n3093 = n971 & ~n3092;
  assign n3094 = n975 & ~n3093;
  assign n3095 = n979 & ~n3094;
  assign n3096 = n983 & ~n3095;
  assign n3097 = n987 & ~n3096;
  assign n3098 = n991 & ~n3097;
  assign n3099 = n995 & ~n3098;
  assign n3100 = n999 & ~n3099;
  assign n3101 = n1003 & ~n3100;
  assign n3102 = n1007 & ~n3101;
  assign n3103 = n1011 & ~n3102;
  assign n3104 = n1015 & ~n3103;
  assign n3105 = n1019 & ~n3104;
  assign n3106 = n1023 & ~n3105;
  assign n3107 = n1027 & ~n3106;
  assign n3108 = n1031 & ~n3107;
  assign n3109 = n1035 & ~n3108;
  assign n3110 = n1039 & ~n3109;
  assign n3111 = n1043 & ~n3110;
  assign n3112 = n1047 & ~n3111;
  assign n3113 = n1051 & ~n3112;
  assign n3114 = n1055 & ~n3113;
  assign n3115 = n1059 & ~n3114;
  assign n3116 = n1574 & ~n3115;
  assign n3117 = n1576 & ~n3116;
  assign n3118 = n1837 & ~n3117;
  assign n3119 = n1068 & ~n3118;
  assign n3120 = n1072 & ~n3119;
  assign n3121 = n1076 & ~n3120;
  assign n3122 = n1080 & ~n3121;
  assign n3123 = n1084 & ~n3122;
  assign n3124 = n1088 & ~n3123;
  assign n3125 = n1092 & ~n3124;
  assign n3126 = n1096 & ~n3125;
  assign n3127 = n1100 & ~n3126;
  assign n3128 = n1104 & ~n3127;
  assign n3129 = n1108 & ~n3128;
  assign n3130 = pi150  & ~n1110;
  assign po22  = ~n3129 & n3130;
  assign n3132 = ~n447 & n1119;
  assign n3133 = n1124 & ~n3132;
  assign n3134 = n1128 & ~n3133;
  assign n3135 = n1132 & ~n3134;
  assign n3136 = n1136 & ~n3135;
  assign n3137 = n1140 & ~n3136;
  assign n3138 = n1144 & ~n3137;
  assign n3139 = n1148 & ~n3138;
  assign n3140 = n1152 & ~n3139;
  assign n3141 = n1156 & ~n3140;
  assign n3142 = n1160 & ~n3141;
  assign n3143 = n1164 & ~n3142;
  assign n3144 = n1168 & ~n3143;
  assign n3145 = n1172 & ~n3144;
  assign n3146 = n1176 & ~n3145;
  assign n3147 = n1180 & ~n3146;
  assign n3148 = n1184 & ~n3147;
  assign n3149 = n1188 & ~n3148;
  assign n3150 = n1192 & ~n3149;
  assign n3151 = n1196 & ~n3150;
  assign n3152 = n1200 & ~n3151;
  assign n3153 = n1204 & ~n3152;
  assign n3154 = n1208 & ~n3153;
  assign n3155 = n1212 & ~n3154;
  assign n3156 = n1216 & ~n3155;
  assign n3157 = n1220 & ~n3156;
  assign n3158 = n1224 & ~n3157;
  assign n3159 = n1228 & ~n3158;
  assign n3160 = n1232 & ~n3159;
  assign n3161 = n1236 & ~n3160;
  assign n3162 = n1240 & ~n3161;
  assign n3163 = n1244 & ~n3162;
  assign n3164 = n1248 & ~n3163;
  assign n3165 = n1252 & ~n3164;
  assign n3166 = n1256 & ~n3165;
  assign n3167 = n1260 & ~n3166;
  assign n3168 = n1264 & ~n3167;
  assign n3169 = n1268 & ~n3168;
  assign n3170 = n1272 & ~n3169;
  assign n3171 = n1276 & ~n3170;
  assign n3172 = n1280 & ~n3171;
  assign n3173 = n1284 & ~n3172;
  assign n3174 = n1288 & ~n3173;
  assign n3175 = n1292 & ~n3174;
  assign n3176 = n1296 & ~n3175;
  assign n3177 = n1300 & ~n3176;
  assign n3178 = n1304 & ~n3177;
  assign n3179 = n1308 & ~n3178;
  assign n3180 = n1312 & ~n3179;
  assign n3181 = n1316 & ~n3180;
  assign n3182 = n1320 & ~n3181;
  assign n3183 = n1324 & ~n3182;
  assign n3184 = n1328 & ~n3183;
  assign n3185 = n1332 & ~n3184;
  assign n3186 = n1336 & ~n3185;
  assign n3187 = n1340 & ~n3186;
  assign n3188 = n1344 & ~n3187;
  assign n3189 = n1348 & ~n3188;
  assign n3190 = n1352 & ~n3189;
  assign n3191 = n1356 & ~n3190;
  assign n3192 = n1360 & ~n3191;
  assign n3193 = n1364 & ~n3192;
  assign n3194 = n1368 & ~n3193;
  assign n3195 = n1372 & ~n3194;
  assign n3196 = n1376 & ~n3195;
  assign n3197 = n1380 & ~n3196;
  assign n3198 = n1384 & ~n3197;
  assign n3199 = n1388 & ~n3198;
  assign n3200 = n1392 & ~n3199;
  assign n3201 = n1396 & ~n3200;
  assign n3202 = n1663 & ~n3201;
  assign n3203 = n392 & ~n3202;
  assign n3204 = n396 & ~n3203;
  assign n3205 = n400 & ~n3204;
  assign n3206 = n404 & ~n3205;
  assign n3207 = n408 & ~n3206;
  assign n3208 = n412 & ~n3207;
  assign n3209 = n416 & ~n3208;
  assign n3210 = n420 & ~n3209;
  assign n3211 = n424 & ~n3210;
  assign n3212 = n428 & ~n3211;
  assign n3213 = n432 & ~n3212;
  assign n3214 = n436 & ~n3213;
  assign n3215 = n440 & ~n3214;
  assign n3216 = pi151  & ~n442;
  assign po23  = ~n3215 & n3216;
  assign n3218 = n451 & ~n786;
  assign n3219 = n456 & ~n3218;
  assign n3220 = n460 & ~n3219;
  assign n3221 = n464 & ~n3220;
  assign n3222 = n468 & ~n3221;
  assign n3223 = n472 & ~n3222;
  assign n3224 = n476 & ~n3223;
  assign n3225 = n480 & ~n3224;
  assign n3226 = n484 & ~n3225;
  assign n3227 = n488 & ~n3226;
  assign n3228 = n492 & ~n3227;
  assign n3229 = n496 & ~n3228;
  assign n3230 = n500 & ~n3229;
  assign n3231 = n504 & ~n3230;
  assign n3232 = n508 & ~n3231;
  assign n3233 = n512 & ~n3232;
  assign n3234 = n516 & ~n3233;
  assign n3235 = n520 & ~n3234;
  assign n3236 = n524 & ~n3235;
  assign n3237 = n528 & ~n3236;
  assign n3238 = n532 & ~n3237;
  assign n3239 = n536 & ~n3238;
  assign n3240 = n540 & ~n3239;
  assign n3241 = n544 & ~n3240;
  assign n3242 = n548 & ~n3241;
  assign n3243 = n552 & ~n3242;
  assign n3244 = n556 & ~n3243;
  assign n3245 = n560 & ~n3244;
  assign n3246 = n564 & ~n3245;
  assign n3247 = n568 & ~n3246;
  assign n3248 = n572 & ~n3247;
  assign n3249 = n576 & ~n3248;
  assign n3250 = n580 & ~n3249;
  assign n3251 = n584 & ~n3250;
  assign n3252 = n588 & ~n3251;
  assign n3253 = n592 & ~n3252;
  assign n3254 = n596 & ~n3253;
  assign n3255 = n600 & ~n3254;
  assign n3256 = n604 & ~n3255;
  assign n3257 = n608 & ~n3256;
  assign n3258 = n612 & ~n3257;
  assign n3259 = n616 & ~n3258;
  assign n3260 = n620 & ~n3259;
  assign n3261 = n624 & ~n3260;
  assign n3262 = n628 & ~n3261;
  assign n3263 = n632 & ~n3262;
  assign n3264 = n636 & ~n3263;
  assign n3265 = n640 & ~n3264;
  assign n3266 = n644 & ~n3265;
  assign n3267 = n648 & ~n3266;
  assign n3268 = n652 & ~n3267;
  assign n3269 = n656 & ~n3268;
  assign n3270 = n660 & ~n3269;
  assign n3271 = n664 & ~n3270;
  assign n3272 = n668 & ~n3271;
  assign n3273 = n672 & ~n3272;
  assign n3274 = n676 & ~n3273;
  assign n3275 = n680 & ~n3274;
  assign n3276 = n684 & ~n3275;
  assign n3277 = n688 & ~n3276;
  assign n3278 = n692 & ~n3277;
  assign n3279 = n696 & ~n3278;
  assign n3280 = n700 & ~n3279;
  assign n3281 = n704 & ~n3280;
  assign n3282 = n708 & ~n3281;
  assign n3283 = n712 & ~n3282;
  assign n3284 = n716 & ~n3283;
  assign n3285 = n720 & ~n3284;
  assign n3286 = n1484 & ~n3285;
  assign n3287 = n1486 & ~n3286;
  assign n3288 = n1750 & ~n3287;
  assign n3289 = n731 & ~n3288;
  assign n3290 = n735 & ~n3289;
  assign n3291 = n739 & ~n3290;
  assign n3292 = n743 & ~n3291;
  assign n3293 = n747 & ~n3292;
  assign n3294 = n751 & ~n3293;
  assign n3295 = n755 & ~n3294;
  assign n3296 = n759 & ~n3295;
  assign n3297 = n763 & ~n3296;
  assign n3298 = n767 & ~n3297;
  assign n3299 = n771 & ~n3298;
  assign n3300 = n775 & ~n3299;
  assign n3301 = n779 & ~n3300;
  assign n3302 = pi152  & ~n781;
  assign po24  = ~n3301 & n3302;
  assign n3304 = n790 & ~n1123;
  assign n3305 = n795 & ~n3304;
  assign n3306 = n799 & ~n3305;
  assign n3307 = n803 & ~n3306;
  assign n3308 = n807 & ~n3307;
  assign n3309 = n811 & ~n3308;
  assign n3310 = n815 & ~n3309;
  assign n3311 = n819 & ~n3310;
  assign n3312 = n823 & ~n3311;
  assign n3313 = n827 & ~n3312;
  assign n3314 = n831 & ~n3313;
  assign n3315 = n835 & ~n3314;
  assign n3316 = n839 & ~n3315;
  assign n3317 = n843 & ~n3316;
  assign n3318 = n847 & ~n3317;
  assign n3319 = n851 & ~n3318;
  assign n3320 = n855 & ~n3319;
  assign n3321 = n859 & ~n3320;
  assign n3322 = n863 & ~n3321;
  assign n3323 = n867 & ~n3322;
  assign n3324 = n871 & ~n3323;
  assign n3325 = n875 & ~n3324;
  assign n3326 = n879 & ~n3325;
  assign n3327 = n883 & ~n3326;
  assign n3328 = n887 & ~n3327;
  assign n3329 = n891 & ~n3328;
  assign n3330 = n895 & ~n3329;
  assign n3331 = n899 & ~n3330;
  assign n3332 = n903 & ~n3331;
  assign n3333 = n907 & ~n3332;
  assign n3334 = n911 & ~n3333;
  assign n3335 = n915 & ~n3334;
  assign n3336 = n919 & ~n3335;
  assign n3337 = n923 & ~n3336;
  assign n3338 = n927 & ~n3337;
  assign n3339 = n931 & ~n3338;
  assign n3340 = n935 & ~n3339;
  assign n3341 = n939 & ~n3340;
  assign n3342 = n943 & ~n3341;
  assign n3343 = n947 & ~n3342;
  assign n3344 = n951 & ~n3343;
  assign n3345 = n955 & ~n3344;
  assign n3346 = n959 & ~n3345;
  assign n3347 = n963 & ~n3346;
  assign n3348 = n967 & ~n3347;
  assign n3349 = n971 & ~n3348;
  assign n3350 = n975 & ~n3349;
  assign n3351 = n979 & ~n3350;
  assign n3352 = n983 & ~n3351;
  assign n3353 = n987 & ~n3352;
  assign n3354 = n991 & ~n3353;
  assign n3355 = n995 & ~n3354;
  assign n3356 = n999 & ~n3355;
  assign n3357 = n1003 & ~n3356;
  assign n3358 = n1007 & ~n3357;
  assign n3359 = n1011 & ~n3358;
  assign n3360 = n1015 & ~n3359;
  assign n3361 = n1019 & ~n3360;
  assign n3362 = n1023 & ~n3361;
  assign n3363 = n1027 & ~n3362;
  assign n3364 = n1031 & ~n3363;
  assign n3365 = n1035 & ~n3364;
  assign n3366 = n1039 & ~n3365;
  assign n3367 = n1043 & ~n3366;
  assign n3368 = n1047 & ~n3367;
  assign n3369 = n1051 & ~n3368;
  assign n3370 = n1055 & ~n3369;
  assign n3371 = n1059 & ~n3370;
  assign n3372 = n1574 & ~n3371;
  assign n3373 = n1576 & ~n3372;
  assign n3374 = n1837 & ~n3373;
  assign n3375 = n1068 & ~n3374;
  assign n3376 = n1072 & ~n3375;
  assign n3377 = n1076 & ~n3376;
  assign n3378 = n1080 & ~n3377;
  assign n3379 = n1084 & ~n3378;
  assign n3380 = n1088 & ~n3379;
  assign n3381 = n1092 & ~n3380;
  assign n3382 = n1096 & ~n3381;
  assign n3383 = n1100 & ~n3382;
  assign n3384 = n1104 & ~n3383;
  assign n3385 = n1108 & ~n3384;
  assign n3386 = n1112 & ~n3385;
  assign n3387 = n1116 & ~n3386;
  assign n3388 = pi153  & ~n1118;
  assign po25  = ~n3387 & n3388;
  assign n3390 = ~n455 & n1127;
  assign n3391 = n1132 & ~n3390;
  assign n3392 = n1136 & ~n3391;
  assign n3393 = n1140 & ~n3392;
  assign n3394 = n1144 & ~n3393;
  assign n3395 = n1148 & ~n3394;
  assign n3396 = n1152 & ~n3395;
  assign n3397 = n1156 & ~n3396;
  assign n3398 = n1160 & ~n3397;
  assign n3399 = n1164 & ~n3398;
  assign n3400 = n1168 & ~n3399;
  assign n3401 = n1172 & ~n3400;
  assign n3402 = n1176 & ~n3401;
  assign n3403 = n1180 & ~n3402;
  assign n3404 = n1184 & ~n3403;
  assign n3405 = n1188 & ~n3404;
  assign n3406 = n1192 & ~n3405;
  assign n3407 = n1196 & ~n3406;
  assign n3408 = n1200 & ~n3407;
  assign n3409 = n1204 & ~n3408;
  assign n3410 = n1208 & ~n3409;
  assign n3411 = n1212 & ~n3410;
  assign n3412 = n1216 & ~n3411;
  assign n3413 = n1220 & ~n3412;
  assign n3414 = n1224 & ~n3413;
  assign n3415 = n1228 & ~n3414;
  assign n3416 = n1232 & ~n3415;
  assign n3417 = n1236 & ~n3416;
  assign n3418 = n1240 & ~n3417;
  assign n3419 = n1244 & ~n3418;
  assign n3420 = n1248 & ~n3419;
  assign n3421 = n1252 & ~n3420;
  assign n3422 = n1256 & ~n3421;
  assign n3423 = n1260 & ~n3422;
  assign n3424 = n1264 & ~n3423;
  assign n3425 = n1268 & ~n3424;
  assign n3426 = n1272 & ~n3425;
  assign n3427 = n1276 & ~n3426;
  assign n3428 = n1280 & ~n3427;
  assign n3429 = n1284 & ~n3428;
  assign n3430 = n1288 & ~n3429;
  assign n3431 = n1292 & ~n3430;
  assign n3432 = n1296 & ~n3431;
  assign n3433 = n1300 & ~n3432;
  assign n3434 = n1304 & ~n3433;
  assign n3435 = n1308 & ~n3434;
  assign n3436 = n1312 & ~n3435;
  assign n3437 = n1316 & ~n3436;
  assign n3438 = n1320 & ~n3437;
  assign n3439 = n1324 & ~n3438;
  assign n3440 = n1328 & ~n3439;
  assign n3441 = n1332 & ~n3440;
  assign n3442 = n1336 & ~n3441;
  assign n3443 = n1340 & ~n3442;
  assign n3444 = n1344 & ~n3443;
  assign n3445 = n1348 & ~n3444;
  assign n3446 = n1352 & ~n3445;
  assign n3447 = n1356 & ~n3446;
  assign n3448 = n1360 & ~n3447;
  assign n3449 = n1364 & ~n3448;
  assign n3450 = n1368 & ~n3449;
  assign n3451 = n1372 & ~n3450;
  assign n3452 = n1376 & ~n3451;
  assign n3453 = n1380 & ~n3452;
  assign n3454 = n1384 & ~n3453;
  assign n3455 = n1388 & ~n3454;
  assign n3456 = n1392 & ~n3455;
  assign n3457 = n1396 & ~n3456;
  assign n3458 = n1663 & ~n3457;
  assign n3459 = n392 & ~n3458;
  assign n3460 = n396 & ~n3459;
  assign n3461 = n400 & ~n3460;
  assign n3462 = n404 & ~n3461;
  assign n3463 = n408 & ~n3462;
  assign n3464 = n412 & ~n3463;
  assign n3465 = n416 & ~n3464;
  assign n3466 = n420 & ~n3465;
  assign n3467 = n424 & ~n3466;
  assign n3468 = n428 & ~n3467;
  assign n3469 = n432 & ~n3468;
  assign n3470 = n436 & ~n3469;
  assign n3471 = n440 & ~n3470;
  assign n3472 = n444 & ~n3471;
  assign n3473 = n448 & ~n3472;
  assign n3474 = pi154  & ~n450;
  assign po26  = ~n3473 & n3474;
  assign n3476 = n459 & ~n794;
  assign n3477 = n464 & ~n3476;
  assign n3478 = n468 & ~n3477;
  assign n3479 = n472 & ~n3478;
  assign n3480 = n476 & ~n3479;
  assign n3481 = n480 & ~n3480;
  assign n3482 = n484 & ~n3481;
  assign n3483 = n488 & ~n3482;
  assign n3484 = n492 & ~n3483;
  assign n3485 = n496 & ~n3484;
  assign n3486 = n500 & ~n3485;
  assign n3487 = n504 & ~n3486;
  assign n3488 = n508 & ~n3487;
  assign n3489 = n512 & ~n3488;
  assign n3490 = n516 & ~n3489;
  assign n3491 = n520 & ~n3490;
  assign n3492 = n524 & ~n3491;
  assign n3493 = n528 & ~n3492;
  assign n3494 = n532 & ~n3493;
  assign n3495 = n536 & ~n3494;
  assign n3496 = n540 & ~n3495;
  assign n3497 = n544 & ~n3496;
  assign n3498 = n548 & ~n3497;
  assign n3499 = n552 & ~n3498;
  assign n3500 = n556 & ~n3499;
  assign n3501 = n560 & ~n3500;
  assign n3502 = n564 & ~n3501;
  assign n3503 = n568 & ~n3502;
  assign n3504 = n572 & ~n3503;
  assign n3505 = n576 & ~n3504;
  assign n3506 = n580 & ~n3505;
  assign n3507 = n584 & ~n3506;
  assign n3508 = n588 & ~n3507;
  assign n3509 = n592 & ~n3508;
  assign n3510 = n596 & ~n3509;
  assign n3511 = n600 & ~n3510;
  assign n3512 = n604 & ~n3511;
  assign n3513 = n608 & ~n3512;
  assign n3514 = n612 & ~n3513;
  assign n3515 = n616 & ~n3514;
  assign n3516 = n620 & ~n3515;
  assign n3517 = n624 & ~n3516;
  assign n3518 = n628 & ~n3517;
  assign n3519 = n632 & ~n3518;
  assign n3520 = n636 & ~n3519;
  assign n3521 = n640 & ~n3520;
  assign n3522 = n644 & ~n3521;
  assign n3523 = n648 & ~n3522;
  assign n3524 = n652 & ~n3523;
  assign n3525 = n656 & ~n3524;
  assign n3526 = n660 & ~n3525;
  assign n3527 = n664 & ~n3526;
  assign n3528 = n668 & ~n3527;
  assign n3529 = n672 & ~n3528;
  assign n3530 = n676 & ~n3529;
  assign n3531 = n680 & ~n3530;
  assign n3532 = n684 & ~n3531;
  assign n3533 = n688 & ~n3532;
  assign n3534 = n692 & ~n3533;
  assign n3535 = n696 & ~n3534;
  assign n3536 = n700 & ~n3535;
  assign n3537 = n704 & ~n3536;
  assign n3538 = n708 & ~n3537;
  assign n3539 = n712 & ~n3538;
  assign n3540 = n716 & ~n3539;
  assign n3541 = n720 & ~n3540;
  assign n3542 = n1484 & ~n3541;
  assign n3543 = n1486 & ~n3542;
  assign n3544 = n1750 & ~n3543;
  assign n3545 = n731 & ~n3544;
  assign n3546 = n735 & ~n3545;
  assign n3547 = n739 & ~n3546;
  assign n3548 = n743 & ~n3547;
  assign n3549 = n747 & ~n3548;
  assign n3550 = n751 & ~n3549;
  assign n3551 = n755 & ~n3550;
  assign n3552 = n759 & ~n3551;
  assign n3553 = n763 & ~n3552;
  assign n3554 = n767 & ~n3553;
  assign n3555 = n771 & ~n3554;
  assign n3556 = n775 & ~n3555;
  assign n3557 = n779 & ~n3556;
  assign n3558 = n783 & ~n3557;
  assign n3559 = n787 & ~n3558;
  assign n3560 = pi155  & ~n789;
  assign po27  = ~n3559 & n3560;
  assign n3562 = n798 & ~n1131;
  assign n3563 = n803 & ~n3562;
  assign n3564 = n807 & ~n3563;
  assign n3565 = n811 & ~n3564;
  assign n3566 = n815 & ~n3565;
  assign n3567 = n819 & ~n3566;
  assign n3568 = n823 & ~n3567;
  assign n3569 = n827 & ~n3568;
  assign n3570 = n831 & ~n3569;
  assign n3571 = n835 & ~n3570;
  assign n3572 = n839 & ~n3571;
  assign n3573 = n843 & ~n3572;
  assign n3574 = n847 & ~n3573;
  assign n3575 = n851 & ~n3574;
  assign n3576 = n855 & ~n3575;
  assign n3577 = n859 & ~n3576;
  assign n3578 = n863 & ~n3577;
  assign n3579 = n867 & ~n3578;
  assign n3580 = n871 & ~n3579;
  assign n3581 = n875 & ~n3580;
  assign n3582 = n879 & ~n3581;
  assign n3583 = n883 & ~n3582;
  assign n3584 = n887 & ~n3583;
  assign n3585 = n891 & ~n3584;
  assign n3586 = n895 & ~n3585;
  assign n3587 = n899 & ~n3586;
  assign n3588 = n903 & ~n3587;
  assign n3589 = n907 & ~n3588;
  assign n3590 = n911 & ~n3589;
  assign n3591 = n915 & ~n3590;
  assign n3592 = n919 & ~n3591;
  assign n3593 = n923 & ~n3592;
  assign n3594 = n927 & ~n3593;
  assign n3595 = n931 & ~n3594;
  assign n3596 = n935 & ~n3595;
  assign n3597 = n939 & ~n3596;
  assign n3598 = n943 & ~n3597;
  assign n3599 = n947 & ~n3598;
  assign n3600 = n951 & ~n3599;
  assign n3601 = n955 & ~n3600;
  assign n3602 = n959 & ~n3601;
  assign n3603 = n963 & ~n3602;
  assign n3604 = n967 & ~n3603;
  assign n3605 = n971 & ~n3604;
  assign n3606 = n975 & ~n3605;
  assign n3607 = n979 & ~n3606;
  assign n3608 = n983 & ~n3607;
  assign n3609 = n987 & ~n3608;
  assign n3610 = n991 & ~n3609;
  assign n3611 = n995 & ~n3610;
  assign n3612 = n999 & ~n3611;
  assign n3613 = n1003 & ~n3612;
  assign n3614 = n1007 & ~n3613;
  assign n3615 = n1011 & ~n3614;
  assign n3616 = n1015 & ~n3615;
  assign n3617 = n1019 & ~n3616;
  assign n3618 = n1023 & ~n3617;
  assign n3619 = n1027 & ~n3618;
  assign n3620 = n1031 & ~n3619;
  assign n3621 = n1035 & ~n3620;
  assign n3622 = n1039 & ~n3621;
  assign n3623 = n1043 & ~n3622;
  assign n3624 = n1047 & ~n3623;
  assign n3625 = n1051 & ~n3624;
  assign n3626 = n1055 & ~n3625;
  assign n3627 = n1059 & ~n3626;
  assign n3628 = n1574 & ~n3627;
  assign n3629 = n1576 & ~n3628;
  assign n3630 = n1837 & ~n3629;
  assign n3631 = n1068 & ~n3630;
  assign n3632 = n1072 & ~n3631;
  assign n3633 = n1076 & ~n3632;
  assign n3634 = n1080 & ~n3633;
  assign n3635 = n1084 & ~n3634;
  assign n3636 = n1088 & ~n3635;
  assign n3637 = n1092 & ~n3636;
  assign n3638 = n1096 & ~n3637;
  assign n3639 = n1100 & ~n3638;
  assign n3640 = n1104 & ~n3639;
  assign n3641 = n1108 & ~n3640;
  assign n3642 = n1112 & ~n3641;
  assign n3643 = n1116 & ~n3642;
  assign n3644 = n1120 & ~n3643;
  assign n3645 = n1124 & ~n3644;
  assign n3646 = pi156  & ~n1126;
  assign po28  = ~n3645 & n3646;
  assign n3648 = ~n463 & n1135;
  assign n3649 = n1140 & ~n3648;
  assign n3650 = n1144 & ~n3649;
  assign n3651 = n1148 & ~n3650;
  assign n3652 = n1152 & ~n3651;
  assign n3653 = n1156 & ~n3652;
  assign n3654 = n1160 & ~n3653;
  assign n3655 = n1164 & ~n3654;
  assign n3656 = n1168 & ~n3655;
  assign n3657 = n1172 & ~n3656;
  assign n3658 = n1176 & ~n3657;
  assign n3659 = n1180 & ~n3658;
  assign n3660 = n1184 & ~n3659;
  assign n3661 = n1188 & ~n3660;
  assign n3662 = n1192 & ~n3661;
  assign n3663 = n1196 & ~n3662;
  assign n3664 = n1200 & ~n3663;
  assign n3665 = n1204 & ~n3664;
  assign n3666 = n1208 & ~n3665;
  assign n3667 = n1212 & ~n3666;
  assign n3668 = n1216 & ~n3667;
  assign n3669 = n1220 & ~n3668;
  assign n3670 = n1224 & ~n3669;
  assign n3671 = n1228 & ~n3670;
  assign n3672 = n1232 & ~n3671;
  assign n3673 = n1236 & ~n3672;
  assign n3674 = n1240 & ~n3673;
  assign n3675 = n1244 & ~n3674;
  assign n3676 = n1248 & ~n3675;
  assign n3677 = n1252 & ~n3676;
  assign n3678 = n1256 & ~n3677;
  assign n3679 = n1260 & ~n3678;
  assign n3680 = n1264 & ~n3679;
  assign n3681 = n1268 & ~n3680;
  assign n3682 = n1272 & ~n3681;
  assign n3683 = n1276 & ~n3682;
  assign n3684 = n1280 & ~n3683;
  assign n3685 = n1284 & ~n3684;
  assign n3686 = n1288 & ~n3685;
  assign n3687 = n1292 & ~n3686;
  assign n3688 = n1296 & ~n3687;
  assign n3689 = n1300 & ~n3688;
  assign n3690 = n1304 & ~n3689;
  assign n3691 = n1308 & ~n3690;
  assign n3692 = n1312 & ~n3691;
  assign n3693 = n1316 & ~n3692;
  assign n3694 = n1320 & ~n3693;
  assign n3695 = n1324 & ~n3694;
  assign n3696 = n1328 & ~n3695;
  assign n3697 = n1332 & ~n3696;
  assign n3698 = n1336 & ~n3697;
  assign n3699 = n1340 & ~n3698;
  assign n3700 = n1344 & ~n3699;
  assign n3701 = n1348 & ~n3700;
  assign n3702 = n1352 & ~n3701;
  assign n3703 = n1356 & ~n3702;
  assign n3704 = n1360 & ~n3703;
  assign n3705 = n1364 & ~n3704;
  assign n3706 = n1368 & ~n3705;
  assign n3707 = n1372 & ~n3706;
  assign n3708 = n1376 & ~n3707;
  assign n3709 = n1380 & ~n3708;
  assign n3710 = n1384 & ~n3709;
  assign n3711 = n1388 & ~n3710;
  assign n3712 = n1392 & ~n3711;
  assign n3713 = n1396 & ~n3712;
  assign n3714 = n1663 & ~n3713;
  assign n3715 = n392 & ~n3714;
  assign n3716 = n396 & ~n3715;
  assign n3717 = n400 & ~n3716;
  assign n3718 = n404 & ~n3717;
  assign n3719 = n408 & ~n3718;
  assign n3720 = n412 & ~n3719;
  assign n3721 = n416 & ~n3720;
  assign n3722 = n420 & ~n3721;
  assign n3723 = n424 & ~n3722;
  assign n3724 = n428 & ~n3723;
  assign n3725 = n432 & ~n3724;
  assign n3726 = n436 & ~n3725;
  assign n3727 = n440 & ~n3726;
  assign n3728 = n444 & ~n3727;
  assign n3729 = n448 & ~n3728;
  assign n3730 = n452 & ~n3729;
  assign n3731 = n456 & ~n3730;
  assign n3732 = pi157  & ~n458;
  assign po29  = ~n3731 & n3732;
  assign n3734 = n467 & ~n802;
  assign n3735 = n472 & ~n3734;
  assign n3736 = n476 & ~n3735;
  assign n3737 = n480 & ~n3736;
  assign n3738 = n484 & ~n3737;
  assign n3739 = n488 & ~n3738;
  assign n3740 = n492 & ~n3739;
  assign n3741 = n496 & ~n3740;
  assign n3742 = n500 & ~n3741;
  assign n3743 = n504 & ~n3742;
  assign n3744 = n508 & ~n3743;
  assign n3745 = n512 & ~n3744;
  assign n3746 = n516 & ~n3745;
  assign n3747 = n520 & ~n3746;
  assign n3748 = n524 & ~n3747;
  assign n3749 = n528 & ~n3748;
  assign n3750 = n532 & ~n3749;
  assign n3751 = n536 & ~n3750;
  assign n3752 = n540 & ~n3751;
  assign n3753 = n544 & ~n3752;
  assign n3754 = n548 & ~n3753;
  assign n3755 = n552 & ~n3754;
  assign n3756 = n556 & ~n3755;
  assign n3757 = n560 & ~n3756;
  assign n3758 = n564 & ~n3757;
  assign n3759 = n568 & ~n3758;
  assign n3760 = n572 & ~n3759;
  assign n3761 = n576 & ~n3760;
  assign n3762 = n580 & ~n3761;
  assign n3763 = n584 & ~n3762;
  assign n3764 = n588 & ~n3763;
  assign n3765 = n592 & ~n3764;
  assign n3766 = n596 & ~n3765;
  assign n3767 = n600 & ~n3766;
  assign n3768 = n604 & ~n3767;
  assign n3769 = n608 & ~n3768;
  assign n3770 = n612 & ~n3769;
  assign n3771 = n616 & ~n3770;
  assign n3772 = n620 & ~n3771;
  assign n3773 = n624 & ~n3772;
  assign n3774 = n628 & ~n3773;
  assign n3775 = n632 & ~n3774;
  assign n3776 = n636 & ~n3775;
  assign n3777 = n640 & ~n3776;
  assign n3778 = n644 & ~n3777;
  assign n3779 = n648 & ~n3778;
  assign n3780 = n652 & ~n3779;
  assign n3781 = n656 & ~n3780;
  assign n3782 = n660 & ~n3781;
  assign n3783 = n664 & ~n3782;
  assign n3784 = n668 & ~n3783;
  assign n3785 = n672 & ~n3784;
  assign n3786 = n676 & ~n3785;
  assign n3787 = n680 & ~n3786;
  assign n3788 = n684 & ~n3787;
  assign n3789 = n688 & ~n3788;
  assign n3790 = n692 & ~n3789;
  assign n3791 = n696 & ~n3790;
  assign n3792 = n700 & ~n3791;
  assign n3793 = n704 & ~n3792;
  assign n3794 = n708 & ~n3793;
  assign n3795 = n712 & ~n3794;
  assign n3796 = n716 & ~n3795;
  assign n3797 = n720 & ~n3796;
  assign n3798 = n1484 & ~n3797;
  assign n3799 = n1486 & ~n3798;
  assign n3800 = n1750 & ~n3799;
  assign n3801 = n731 & ~n3800;
  assign n3802 = n735 & ~n3801;
  assign n3803 = n739 & ~n3802;
  assign n3804 = n743 & ~n3803;
  assign n3805 = n747 & ~n3804;
  assign n3806 = n751 & ~n3805;
  assign n3807 = n755 & ~n3806;
  assign n3808 = n759 & ~n3807;
  assign n3809 = n763 & ~n3808;
  assign n3810 = n767 & ~n3809;
  assign n3811 = n771 & ~n3810;
  assign n3812 = n775 & ~n3811;
  assign n3813 = n779 & ~n3812;
  assign n3814 = n783 & ~n3813;
  assign n3815 = n787 & ~n3814;
  assign n3816 = n791 & ~n3815;
  assign n3817 = n795 & ~n3816;
  assign n3818 = pi158  & ~n797;
  assign po30  = ~n3817 & n3818;
  assign n3820 = n806 & ~n1139;
  assign n3821 = n811 & ~n3820;
  assign n3822 = n815 & ~n3821;
  assign n3823 = n819 & ~n3822;
  assign n3824 = n823 & ~n3823;
  assign n3825 = n827 & ~n3824;
  assign n3826 = n831 & ~n3825;
  assign n3827 = n835 & ~n3826;
  assign n3828 = n839 & ~n3827;
  assign n3829 = n843 & ~n3828;
  assign n3830 = n847 & ~n3829;
  assign n3831 = n851 & ~n3830;
  assign n3832 = n855 & ~n3831;
  assign n3833 = n859 & ~n3832;
  assign n3834 = n863 & ~n3833;
  assign n3835 = n867 & ~n3834;
  assign n3836 = n871 & ~n3835;
  assign n3837 = n875 & ~n3836;
  assign n3838 = n879 & ~n3837;
  assign n3839 = n883 & ~n3838;
  assign n3840 = n887 & ~n3839;
  assign n3841 = n891 & ~n3840;
  assign n3842 = n895 & ~n3841;
  assign n3843 = n899 & ~n3842;
  assign n3844 = n903 & ~n3843;
  assign n3845 = n907 & ~n3844;
  assign n3846 = n911 & ~n3845;
  assign n3847 = n915 & ~n3846;
  assign n3848 = n919 & ~n3847;
  assign n3849 = n923 & ~n3848;
  assign n3850 = n927 & ~n3849;
  assign n3851 = n931 & ~n3850;
  assign n3852 = n935 & ~n3851;
  assign n3853 = n939 & ~n3852;
  assign n3854 = n943 & ~n3853;
  assign n3855 = n947 & ~n3854;
  assign n3856 = n951 & ~n3855;
  assign n3857 = n955 & ~n3856;
  assign n3858 = n959 & ~n3857;
  assign n3859 = n963 & ~n3858;
  assign n3860 = n967 & ~n3859;
  assign n3861 = n971 & ~n3860;
  assign n3862 = n975 & ~n3861;
  assign n3863 = n979 & ~n3862;
  assign n3864 = n983 & ~n3863;
  assign n3865 = n987 & ~n3864;
  assign n3866 = n991 & ~n3865;
  assign n3867 = n995 & ~n3866;
  assign n3868 = n999 & ~n3867;
  assign n3869 = n1003 & ~n3868;
  assign n3870 = n1007 & ~n3869;
  assign n3871 = n1011 & ~n3870;
  assign n3872 = n1015 & ~n3871;
  assign n3873 = n1019 & ~n3872;
  assign n3874 = n1023 & ~n3873;
  assign n3875 = n1027 & ~n3874;
  assign n3876 = n1031 & ~n3875;
  assign n3877 = n1035 & ~n3876;
  assign n3878 = n1039 & ~n3877;
  assign n3879 = n1043 & ~n3878;
  assign n3880 = n1047 & ~n3879;
  assign n3881 = n1051 & ~n3880;
  assign n3882 = n1055 & ~n3881;
  assign n3883 = n1059 & ~n3882;
  assign n3884 = n1574 & ~n3883;
  assign n3885 = n1576 & ~n3884;
  assign n3886 = n1837 & ~n3885;
  assign n3887 = n1068 & ~n3886;
  assign n3888 = n1072 & ~n3887;
  assign n3889 = n1076 & ~n3888;
  assign n3890 = n1080 & ~n3889;
  assign n3891 = n1084 & ~n3890;
  assign n3892 = n1088 & ~n3891;
  assign n3893 = n1092 & ~n3892;
  assign n3894 = n1096 & ~n3893;
  assign n3895 = n1100 & ~n3894;
  assign n3896 = n1104 & ~n3895;
  assign n3897 = n1108 & ~n3896;
  assign n3898 = n1112 & ~n3897;
  assign n3899 = n1116 & ~n3898;
  assign n3900 = n1120 & ~n3899;
  assign n3901 = n1124 & ~n3900;
  assign n3902 = n1128 & ~n3901;
  assign n3903 = n1132 & ~n3902;
  assign n3904 = pi159  & ~n1134;
  assign po31  = ~n3903 & n3904;
  assign n3906 = ~n471 & n1143;
  assign n3907 = n1148 & ~n3906;
  assign n3908 = n1152 & ~n3907;
  assign n3909 = n1156 & ~n3908;
  assign n3910 = n1160 & ~n3909;
  assign n3911 = n1164 & ~n3910;
  assign n3912 = n1168 & ~n3911;
  assign n3913 = n1172 & ~n3912;
  assign n3914 = n1176 & ~n3913;
  assign n3915 = n1180 & ~n3914;
  assign n3916 = n1184 & ~n3915;
  assign n3917 = n1188 & ~n3916;
  assign n3918 = n1192 & ~n3917;
  assign n3919 = n1196 & ~n3918;
  assign n3920 = n1200 & ~n3919;
  assign n3921 = n1204 & ~n3920;
  assign n3922 = n1208 & ~n3921;
  assign n3923 = n1212 & ~n3922;
  assign n3924 = n1216 & ~n3923;
  assign n3925 = n1220 & ~n3924;
  assign n3926 = n1224 & ~n3925;
  assign n3927 = n1228 & ~n3926;
  assign n3928 = n1232 & ~n3927;
  assign n3929 = n1236 & ~n3928;
  assign n3930 = n1240 & ~n3929;
  assign n3931 = n1244 & ~n3930;
  assign n3932 = n1248 & ~n3931;
  assign n3933 = n1252 & ~n3932;
  assign n3934 = n1256 & ~n3933;
  assign n3935 = n1260 & ~n3934;
  assign n3936 = n1264 & ~n3935;
  assign n3937 = n1268 & ~n3936;
  assign n3938 = n1272 & ~n3937;
  assign n3939 = n1276 & ~n3938;
  assign n3940 = n1280 & ~n3939;
  assign n3941 = n1284 & ~n3940;
  assign n3942 = n1288 & ~n3941;
  assign n3943 = n1292 & ~n3942;
  assign n3944 = n1296 & ~n3943;
  assign n3945 = n1300 & ~n3944;
  assign n3946 = n1304 & ~n3945;
  assign n3947 = n1308 & ~n3946;
  assign n3948 = n1312 & ~n3947;
  assign n3949 = n1316 & ~n3948;
  assign n3950 = n1320 & ~n3949;
  assign n3951 = n1324 & ~n3950;
  assign n3952 = n1328 & ~n3951;
  assign n3953 = n1332 & ~n3952;
  assign n3954 = n1336 & ~n3953;
  assign n3955 = n1340 & ~n3954;
  assign n3956 = n1344 & ~n3955;
  assign n3957 = n1348 & ~n3956;
  assign n3958 = n1352 & ~n3957;
  assign n3959 = n1356 & ~n3958;
  assign n3960 = n1360 & ~n3959;
  assign n3961 = n1364 & ~n3960;
  assign n3962 = n1368 & ~n3961;
  assign n3963 = n1372 & ~n3962;
  assign n3964 = n1376 & ~n3963;
  assign n3965 = n1380 & ~n3964;
  assign n3966 = n1384 & ~n3965;
  assign n3967 = n1388 & ~n3966;
  assign n3968 = n1392 & ~n3967;
  assign n3969 = n1396 & ~n3968;
  assign n3970 = n1663 & ~n3969;
  assign n3971 = n392 & ~n3970;
  assign n3972 = n396 & ~n3971;
  assign n3973 = n400 & ~n3972;
  assign n3974 = n404 & ~n3973;
  assign n3975 = n408 & ~n3974;
  assign n3976 = n412 & ~n3975;
  assign n3977 = n416 & ~n3976;
  assign n3978 = n420 & ~n3977;
  assign n3979 = n424 & ~n3978;
  assign n3980 = n428 & ~n3979;
  assign n3981 = n432 & ~n3980;
  assign n3982 = n436 & ~n3981;
  assign n3983 = n440 & ~n3982;
  assign n3984 = n444 & ~n3983;
  assign n3985 = n448 & ~n3984;
  assign n3986 = n452 & ~n3985;
  assign n3987 = n456 & ~n3986;
  assign n3988 = n460 & ~n3987;
  assign n3989 = n464 & ~n3988;
  assign n3990 = pi160  & ~n466;
  assign po32  = ~n3989 & n3990;
  assign n3992 = n475 & ~n810;
  assign n3993 = n480 & ~n3992;
  assign n3994 = n484 & ~n3993;
  assign n3995 = n488 & ~n3994;
  assign n3996 = n492 & ~n3995;
  assign n3997 = n496 & ~n3996;
  assign n3998 = n500 & ~n3997;
  assign n3999 = n504 & ~n3998;
  assign n4000 = n508 & ~n3999;
  assign n4001 = n512 & ~n4000;
  assign n4002 = n516 & ~n4001;
  assign n4003 = n520 & ~n4002;
  assign n4004 = n524 & ~n4003;
  assign n4005 = n528 & ~n4004;
  assign n4006 = n532 & ~n4005;
  assign n4007 = n536 & ~n4006;
  assign n4008 = n540 & ~n4007;
  assign n4009 = n544 & ~n4008;
  assign n4010 = n548 & ~n4009;
  assign n4011 = n552 & ~n4010;
  assign n4012 = n556 & ~n4011;
  assign n4013 = n560 & ~n4012;
  assign n4014 = n564 & ~n4013;
  assign n4015 = n568 & ~n4014;
  assign n4016 = n572 & ~n4015;
  assign n4017 = n576 & ~n4016;
  assign n4018 = n580 & ~n4017;
  assign n4019 = n584 & ~n4018;
  assign n4020 = n588 & ~n4019;
  assign n4021 = n592 & ~n4020;
  assign n4022 = n596 & ~n4021;
  assign n4023 = n600 & ~n4022;
  assign n4024 = n604 & ~n4023;
  assign n4025 = n608 & ~n4024;
  assign n4026 = n612 & ~n4025;
  assign n4027 = n616 & ~n4026;
  assign n4028 = n620 & ~n4027;
  assign n4029 = n624 & ~n4028;
  assign n4030 = n628 & ~n4029;
  assign n4031 = n632 & ~n4030;
  assign n4032 = n636 & ~n4031;
  assign n4033 = n640 & ~n4032;
  assign n4034 = n644 & ~n4033;
  assign n4035 = n648 & ~n4034;
  assign n4036 = n652 & ~n4035;
  assign n4037 = n656 & ~n4036;
  assign n4038 = n660 & ~n4037;
  assign n4039 = n664 & ~n4038;
  assign n4040 = n668 & ~n4039;
  assign n4041 = n672 & ~n4040;
  assign n4042 = n676 & ~n4041;
  assign n4043 = n680 & ~n4042;
  assign n4044 = n684 & ~n4043;
  assign n4045 = n688 & ~n4044;
  assign n4046 = n692 & ~n4045;
  assign n4047 = n696 & ~n4046;
  assign n4048 = n700 & ~n4047;
  assign n4049 = n704 & ~n4048;
  assign n4050 = n708 & ~n4049;
  assign n4051 = n712 & ~n4050;
  assign n4052 = n716 & ~n4051;
  assign n4053 = n720 & ~n4052;
  assign n4054 = n1484 & ~n4053;
  assign n4055 = n1486 & ~n4054;
  assign n4056 = n1750 & ~n4055;
  assign n4057 = n731 & ~n4056;
  assign n4058 = n735 & ~n4057;
  assign n4059 = n739 & ~n4058;
  assign n4060 = n743 & ~n4059;
  assign n4061 = n747 & ~n4060;
  assign n4062 = n751 & ~n4061;
  assign n4063 = n755 & ~n4062;
  assign n4064 = n759 & ~n4063;
  assign n4065 = n763 & ~n4064;
  assign n4066 = n767 & ~n4065;
  assign n4067 = n771 & ~n4066;
  assign n4068 = n775 & ~n4067;
  assign n4069 = n779 & ~n4068;
  assign n4070 = n783 & ~n4069;
  assign n4071 = n787 & ~n4070;
  assign n4072 = n791 & ~n4071;
  assign n4073 = n795 & ~n4072;
  assign n4074 = n799 & ~n4073;
  assign n4075 = n803 & ~n4074;
  assign n4076 = pi161  & ~n805;
  assign po33  = ~n4075 & n4076;
  assign n4078 = n814 & ~n1147;
  assign n4079 = n819 & ~n4078;
  assign n4080 = n823 & ~n4079;
  assign n4081 = n827 & ~n4080;
  assign n4082 = n831 & ~n4081;
  assign n4083 = n835 & ~n4082;
  assign n4084 = n839 & ~n4083;
  assign n4085 = n843 & ~n4084;
  assign n4086 = n847 & ~n4085;
  assign n4087 = n851 & ~n4086;
  assign n4088 = n855 & ~n4087;
  assign n4089 = n859 & ~n4088;
  assign n4090 = n863 & ~n4089;
  assign n4091 = n867 & ~n4090;
  assign n4092 = n871 & ~n4091;
  assign n4093 = n875 & ~n4092;
  assign n4094 = n879 & ~n4093;
  assign n4095 = n883 & ~n4094;
  assign n4096 = n887 & ~n4095;
  assign n4097 = n891 & ~n4096;
  assign n4098 = n895 & ~n4097;
  assign n4099 = n899 & ~n4098;
  assign n4100 = n903 & ~n4099;
  assign n4101 = n907 & ~n4100;
  assign n4102 = n911 & ~n4101;
  assign n4103 = n915 & ~n4102;
  assign n4104 = n919 & ~n4103;
  assign n4105 = n923 & ~n4104;
  assign n4106 = n927 & ~n4105;
  assign n4107 = n931 & ~n4106;
  assign n4108 = n935 & ~n4107;
  assign n4109 = n939 & ~n4108;
  assign n4110 = n943 & ~n4109;
  assign n4111 = n947 & ~n4110;
  assign n4112 = n951 & ~n4111;
  assign n4113 = n955 & ~n4112;
  assign n4114 = n959 & ~n4113;
  assign n4115 = n963 & ~n4114;
  assign n4116 = n967 & ~n4115;
  assign n4117 = n971 & ~n4116;
  assign n4118 = n975 & ~n4117;
  assign n4119 = n979 & ~n4118;
  assign n4120 = n983 & ~n4119;
  assign n4121 = n987 & ~n4120;
  assign n4122 = n991 & ~n4121;
  assign n4123 = n995 & ~n4122;
  assign n4124 = n999 & ~n4123;
  assign n4125 = n1003 & ~n4124;
  assign n4126 = n1007 & ~n4125;
  assign n4127 = n1011 & ~n4126;
  assign n4128 = n1015 & ~n4127;
  assign n4129 = n1019 & ~n4128;
  assign n4130 = n1023 & ~n4129;
  assign n4131 = n1027 & ~n4130;
  assign n4132 = n1031 & ~n4131;
  assign n4133 = n1035 & ~n4132;
  assign n4134 = n1039 & ~n4133;
  assign n4135 = n1043 & ~n4134;
  assign n4136 = n1047 & ~n4135;
  assign n4137 = n1051 & ~n4136;
  assign n4138 = n1055 & ~n4137;
  assign n4139 = n1059 & ~n4138;
  assign n4140 = n1574 & ~n4139;
  assign n4141 = n1576 & ~n4140;
  assign n4142 = n1837 & ~n4141;
  assign n4143 = n1068 & ~n4142;
  assign n4144 = n1072 & ~n4143;
  assign n4145 = n1076 & ~n4144;
  assign n4146 = n1080 & ~n4145;
  assign n4147 = n1084 & ~n4146;
  assign n4148 = n1088 & ~n4147;
  assign n4149 = n1092 & ~n4148;
  assign n4150 = n1096 & ~n4149;
  assign n4151 = n1100 & ~n4150;
  assign n4152 = n1104 & ~n4151;
  assign n4153 = n1108 & ~n4152;
  assign n4154 = n1112 & ~n4153;
  assign n4155 = n1116 & ~n4154;
  assign n4156 = n1120 & ~n4155;
  assign n4157 = n1124 & ~n4156;
  assign n4158 = n1128 & ~n4157;
  assign n4159 = n1132 & ~n4158;
  assign n4160 = n1136 & ~n4159;
  assign n4161 = n1140 & ~n4160;
  assign n4162 = pi162  & ~n1142;
  assign po34  = ~n4161 & n4162;
  assign n4164 = ~n479 & n1151;
  assign n4165 = n1156 & ~n4164;
  assign n4166 = n1160 & ~n4165;
  assign n4167 = n1164 & ~n4166;
  assign n4168 = n1168 & ~n4167;
  assign n4169 = n1172 & ~n4168;
  assign n4170 = n1176 & ~n4169;
  assign n4171 = n1180 & ~n4170;
  assign n4172 = n1184 & ~n4171;
  assign n4173 = n1188 & ~n4172;
  assign n4174 = n1192 & ~n4173;
  assign n4175 = n1196 & ~n4174;
  assign n4176 = n1200 & ~n4175;
  assign n4177 = n1204 & ~n4176;
  assign n4178 = n1208 & ~n4177;
  assign n4179 = n1212 & ~n4178;
  assign n4180 = n1216 & ~n4179;
  assign n4181 = n1220 & ~n4180;
  assign n4182 = n1224 & ~n4181;
  assign n4183 = n1228 & ~n4182;
  assign n4184 = n1232 & ~n4183;
  assign n4185 = n1236 & ~n4184;
  assign n4186 = n1240 & ~n4185;
  assign n4187 = n1244 & ~n4186;
  assign n4188 = n1248 & ~n4187;
  assign n4189 = n1252 & ~n4188;
  assign n4190 = n1256 & ~n4189;
  assign n4191 = n1260 & ~n4190;
  assign n4192 = n1264 & ~n4191;
  assign n4193 = n1268 & ~n4192;
  assign n4194 = n1272 & ~n4193;
  assign n4195 = n1276 & ~n4194;
  assign n4196 = n1280 & ~n4195;
  assign n4197 = n1284 & ~n4196;
  assign n4198 = n1288 & ~n4197;
  assign n4199 = n1292 & ~n4198;
  assign n4200 = n1296 & ~n4199;
  assign n4201 = n1300 & ~n4200;
  assign n4202 = n1304 & ~n4201;
  assign n4203 = n1308 & ~n4202;
  assign n4204 = n1312 & ~n4203;
  assign n4205 = n1316 & ~n4204;
  assign n4206 = n1320 & ~n4205;
  assign n4207 = n1324 & ~n4206;
  assign n4208 = n1328 & ~n4207;
  assign n4209 = n1332 & ~n4208;
  assign n4210 = n1336 & ~n4209;
  assign n4211 = n1340 & ~n4210;
  assign n4212 = n1344 & ~n4211;
  assign n4213 = n1348 & ~n4212;
  assign n4214 = n1352 & ~n4213;
  assign n4215 = n1356 & ~n4214;
  assign n4216 = n1360 & ~n4215;
  assign n4217 = n1364 & ~n4216;
  assign n4218 = n1368 & ~n4217;
  assign n4219 = n1372 & ~n4218;
  assign n4220 = n1376 & ~n4219;
  assign n4221 = n1380 & ~n4220;
  assign n4222 = n1384 & ~n4221;
  assign n4223 = n1388 & ~n4222;
  assign n4224 = n1392 & ~n4223;
  assign n4225 = n1396 & ~n4224;
  assign n4226 = n1663 & ~n4225;
  assign n4227 = n392 & ~n4226;
  assign n4228 = n396 & ~n4227;
  assign n4229 = n400 & ~n4228;
  assign n4230 = n404 & ~n4229;
  assign n4231 = n408 & ~n4230;
  assign n4232 = n412 & ~n4231;
  assign n4233 = n416 & ~n4232;
  assign n4234 = n420 & ~n4233;
  assign n4235 = n424 & ~n4234;
  assign n4236 = n428 & ~n4235;
  assign n4237 = n432 & ~n4236;
  assign n4238 = n436 & ~n4237;
  assign n4239 = n440 & ~n4238;
  assign n4240 = n444 & ~n4239;
  assign n4241 = n448 & ~n4240;
  assign n4242 = n452 & ~n4241;
  assign n4243 = n456 & ~n4242;
  assign n4244 = n460 & ~n4243;
  assign n4245 = n464 & ~n4244;
  assign n4246 = n468 & ~n4245;
  assign n4247 = n472 & ~n4246;
  assign n4248 = pi163  & ~n474;
  assign po35  = ~n4247 & n4248;
  assign n4250 = n483 & ~n818;
  assign n4251 = n488 & ~n4250;
  assign n4252 = n492 & ~n4251;
  assign n4253 = n496 & ~n4252;
  assign n4254 = n500 & ~n4253;
  assign n4255 = n504 & ~n4254;
  assign n4256 = n508 & ~n4255;
  assign n4257 = n512 & ~n4256;
  assign n4258 = n516 & ~n4257;
  assign n4259 = n520 & ~n4258;
  assign n4260 = n524 & ~n4259;
  assign n4261 = n528 & ~n4260;
  assign n4262 = n532 & ~n4261;
  assign n4263 = n536 & ~n4262;
  assign n4264 = n540 & ~n4263;
  assign n4265 = n544 & ~n4264;
  assign n4266 = n548 & ~n4265;
  assign n4267 = n552 & ~n4266;
  assign n4268 = n556 & ~n4267;
  assign n4269 = n560 & ~n4268;
  assign n4270 = n564 & ~n4269;
  assign n4271 = n568 & ~n4270;
  assign n4272 = n572 & ~n4271;
  assign n4273 = n576 & ~n4272;
  assign n4274 = n580 & ~n4273;
  assign n4275 = n584 & ~n4274;
  assign n4276 = n588 & ~n4275;
  assign n4277 = n592 & ~n4276;
  assign n4278 = n596 & ~n4277;
  assign n4279 = n600 & ~n4278;
  assign n4280 = n604 & ~n4279;
  assign n4281 = n608 & ~n4280;
  assign n4282 = n612 & ~n4281;
  assign n4283 = n616 & ~n4282;
  assign n4284 = n620 & ~n4283;
  assign n4285 = n624 & ~n4284;
  assign n4286 = n628 & ~n4285;
  assign n4287 = n632 & ~n4286;
  assign n4288 = n636 & ~n4287;
  assign n4289 = n640 & ~n4288;
  assign n4290 = n644 & ~n4289;
  assign n4291 = n648 & ~n4290;
  assign n4292 = n652 & ~n4291;
  assign n4293 = n656 & ~n4292;
  assign n4294 = n660 & ~n4293;
  assign n4295 = n664 & ~n4294;
  assign n4296 = n668 & ~n4295;
  assign n4297 = n672 & ~n4296;
  assign n4298 = n676 & ~n4297;
  assign n4299 = n680 & ~n4298;
  assign n4300 = n684 & ~n4299;
  assign n4301 = n688 & ~n4300;
  assign n4302 = n692 & ~n4301;
  assign n4303 = n696 & ~n4302;
  assign n4304 = n700 & ~n4303;
  assign n4305 = n704 & ~n4304;
  assign n4306 = n708 & ~n4305;
  assign n4307 = n712 & ~n4306;
  assign n4308 = n716 & ~n4307;
  assign n4309 = n720 & ~n4308;
  assign n4310 = n1484 & ~n4309;
  assign n4311 = n1486 & ~n4310;
  assign n4312 = n1750 & ~n4311;
  assign n4313 = n731 & ~n4312;
  assign n4314 = n735 & ~n4313;
  assign n4315 = n739 & ~n4314;
  assign n4316 = n743 & ~n4315;
  assign n4317 = n747 & ~n4316;
  assign n4318 = n751 & ~n4317;
  assign n4319 = n755 & ~n4318;
  assign n4320 = n759 & ~n4319;
  assign n4321 = n763 & ~n4320;
  assign n4322 = n767 & ~n4321;
  assign n4323 = n771 & ~n4322;
  assign n4324 = n775 & ~n4323;
  assign n4325 = n779 & ~n4324;
  assign n4326 = n783 & ~n4325;
  assign n4327 = n787 & ~n4326;
  assign n4328 = n791 & ~n4327;
  assign n4329 = n795 & ~n4328;
  assign n4330 = n799 & ~n4329;
  assign n4331 = n803 & ~n4330;
  assign n4332 = n807 & ~n4331;
  assign n4333 = n811 & ~n4332;
  assign n4334 = pi164  & ~n813;
  assign po36  = ~n4333 & n4334;
  assign n4336 = n822 & ~n1155;
  assign n4337 = n827 & ~n4336;
  assign n4338 = n831 & ~n4337;
  assign n4339 = n835 & ~n4338;
  assign n4340 = n839 & ~n4339;
  assign n4341 = n843 & ~n4340;
  assign n4342 = n847 & ~n4341;
  assign n4343 = n851 & ~n4342;
  assign n4344 = n855 & ~n4343;
  assign n4345 = n859 & ~n4344;
  assign n4346 = n863 & ~n4345;
  assign n4347 = n867 & ~n4346;
  assign n4348 = n871 & ~n4347;
  assign n4349 = n875 & ~n4348;
  assign n4350 = n879 & ~n4349;
  assign n4351 = n883 & ~n4350;
  assign n4352 = n887 & ~n4351;
  assign n4353 = n891 & ~n4352;
  assign n4354 = n895 & ~n4353;
  assign n4355 = n899 & ~n4354;
  assign n4356 = n903 & ~n4355;
  assign n4357 = n907 & ~n4356;
  assign n4358 = n911 & ~n4357;
  assign n4359 = n915 & ~n4358;
  assign n4360 = n919 & ~n4359;
  assign n4361 = n923 & ~n4360;
  assign n4362 = n927 & ~n4361;
  assign n4363 = n931 & ~n4362;
  assign n4364 = n935 & ~n4363;
  assign n4365 = n939 & ~n4364;
  assign n4366 = n943 & ~n4365;
  assign n4367 = n947 & ~n4366;
  assign n4368 = n951 & ~n4367;
  assign n4369 = n955 & ~n4368;
  assign n4370 = n959 & ~n4369;
  assign n4371 = n963 & ~n4370;
  assign n4372 = n967 & ~n4371;
  assign n4373 = n971 & ~n4372;
  assign n4374 = n975 & ~n4373;
  assign n4375 = n979 & ~n4374;
  assign n4376 = n983 & ~n4375;
  assign n4377 = n987 & ~n4376;
  assign n4378 = n991 & ~n4377;
  assign n4379 = n995 & ~n4378;
  assign n4380 = n999 & ~n4379;
  assign n4381 = n1003 & ~n4380;
  assign n4382 = n1007 & ~n4381;
  assign n4383 = n1011 & ~n4382;
  assign n4384 = n1015 & ~n4383;
  assign n4385 = n1019 & ~n4384;
  assign n4386 = n1023 & ~n4385;
  assign n4387 = n1027 & ~n4386;
  assign n4388 = n1031 & ~n4387;
  assign n4389 = n1035 & ~n4388;
  assign n4390 = n1039 & ~n4389;
  assign n4391 = n1043 & ~n4390;
  assign n4392 = n1047 & ~n4391;
  assign n4393 = n1051 & ~n4392;
  assign n4394 = n1055 & ~n4393;
  assign n4395 = n1059 & ~n4394;
  assign n4396 = n1574 & ~n4395;
  assign n4397 = n1576 & ~n4396;
  assign n4398 = n1837 & ~n4397;
  assign n4399 = n1068 & ~n4398;
  assign n4400 = n1072 & ~n4399;
  assign n4401 = n1076 & ~n4400;
  assign n4402 = n1080 & ~n4401;
  assign n4403 = n1084 & ~n4402;
  assign n4404 = n1088 & ~n4403;
  assign n4405 = n1092 & ~n4404;
  assign n4406 = n1096 & ~n4405;
  assign n4407 = n1100 & ~n4406;
  assign n4408 = n1104 & ~n4407;
  assign n4409 = n1108 & ~n4408;
  assign n4410 = n1112 & ~n4409;
  assign n4411 = n1116 & ~n4410;
  assign n4412 = n1120 & ~n4411;
  assign n4413 = n1124 & ~n4412;
  assign n4414 = n1128 & ~n4413;
  assign n4415 = n1132 & ~n4414;
  assign n4416 = n1136 & ~n4415;
  assign n4417 = n1140 & ~n4416;
  assign n4418 = n1144 & ~n4417;
  assign n4419 = n1148 & ~n4418;
  assign n4420 = pi165  & ~n1150;
  assign po37  = ~n4419 & n4420;
  assign n4422 = ~n487 & n1159;
  assign n4423 = n1164 & ~n4422;
  assign n4424 = n1168 & ~n4423;
  assign n4425 = n1172 & ~n4424;
  assign n4426 = n1176 & ~n4425;
  assign n4427 = n1180 & ~n4426;
  assign n4428 = n1184 & ~n4427;
  assign n4429 = n1188 & ~n4428;
  assign n4430 = n1192 & ~n4429;
  assign n4431 = n1196 & ~n4430;
  assign n4432 = n1200 & ~n4431;
  assign n4433 = n1204 & ~n4432;
  assign n4434 = n1208 & ~n4433;
  assign n4435 = n1212 & ~n4434;
  assign n4436 = n1216 & ~n4435;
  assign n4437 = n1220 & ~n4436;
  assign n4438 = n1224 & ~n4437;
  assign n4439 = n1228 & ~n4438;
  assign n4440 = n1232 & ~n4439;
  assign n4441 = n1236 & ~n4440;
  assign n4442 = n1240 & ~n4441;
  assign n4443 = n1244 & ~n4442;
  assign n4444 = n1248 & ~n4443;
  assign n4445 = n1252 & ~n4444;
  assign n4446 = n1256 & ~n4445;
  assign n4447 = n1260 & ~n4446;
  assign n4448 = n1264 & ~n4447;
  assign n4449 = n1268 & ~n4448;
  assign n4450 = n1272 & ~n4449;
  assign n4451 = n1276 & ~n4450;
  assign n4452 = n1280 & ~n4451;
  assign n4453 = n1284 & ~n4452;
  assign n4454 = n1288 & ~n4453;
  assign n4455 = n1292 & ~n4454;
  assign n4456 = n1296 & ~n4455;
  assign n4457 = n1300 & ~n4456;
  assign n4458 = n1304 & ~n4457;
  assign n4459 = n1308 & ~n4458;
  assign n4460 = n1312 & ~n4459;
  assign n4461 = n1316 & ~n4460;
  assign n4462 = n1320 & ~n4461;
  assign n4463 = n1324 & ~n4462;
  assign n4464 = n1328 & ~n4463;
  assign n4465 = n1332 & ~n4464;
  assign n4466 = n1336 & ~n4465;
  assign n4467 = n1340 & ~n4466;
  assign n4468 = n1344 & ~n4467;
  assign n4469 = n1348 & ~n4468;
  assign n4470 = n1352 & ~n4469;
  assign n4471 = n1356 & ~n4470;
  assign n4472 = n1360 & ~n4471;
  assign n4473 = n1364 & ~n4472;
  assign n4474 = n1368 & ~n4473;
  assign n4475 = n1372 & ~n4474;
  assign n4476 = n1376 & ~n4475;
  assign n4477 = n1380 & ~n4476;
  assign n4478 = n1384 & ~n4477;
  assign n4479 = n1388 & ~n4478;
  assign n4480 = n1392 & ~n4479;
  assign n4481 = n1396 & ~n4480;
  assign n4482 = n1663 & ~n4481;
  assign n4483 = n392 & ~n4482;
  assign n4484 = n396 & ~n4483;
  assign n4485 = n400 & ~n4484;
  assign n4486 = n404 & ~n4485;
  assign n4487 = n408 & ~n4486;
  assign n4488 = n412 & ~n4487;
  assign n4489 = n416 & ~n4488;
  assign n4490 = n420 & ~n4489;
  assign n4491 = n424 & ~n4490;
  assign n4492 = n428 & ~n4491;
  assign n4493 = n432 & ~n4492;
  assign n4494 = n436 & ~n4493;
  assign n4495 = n440 & ~n4494;
  assign n4496 = n444 & ~n4495;
  assign n4497 = n448 & ~n4496;
  assign n4498 = n452 & ~n4497;
  assign n4499 = n456 & ~n4498;
  assign n4500 = n460 & ~n4499;
  assign n4501 = n464 & ~n4500;
  assign n4502 = n468 & ~n4501;
  assign n4503 = n472 & ~n4502;
  assign n4504 = n476 & ~n4503;
  assign n4505 = n480 & ~n4504;
  assign n4506 = pi166  & ~n482;
  assign po38  = ~n4505 & n4506;
  assign n4508 = n491 & ~n826;
  assign n4509 = n496 & ~n4508;
  assign n4510 = n500 & ~n4509;
  assign n4511 = n504 & ~n4510;
  assign n4512 = n508 & ~n4511;
  assign n4513 = n512 & ~n4512;
  assign n4514 = n516 & ~n4513;
  assign n4515 = n520 & ~n4514;
  assign n4516 = n524 & ~n4515;
  assign n4517 = n528 & ~n4516;
  assign n4518 = n532 & ~n4517;
  assign n4519 = n536 & ~n4518;
  assign n4520 = n540 & ~n4519;
  assign n4521 = n544 & ~n4520;
  assign n4522 = n548 & ~n4521;
  assign n4523 = n552 & ~n4522;
  assign n4524 = n556 & ~n4523;
  assign n4525 = n560 & ~n4524;
  assign n4526 = n564 & ~n4525;
  assign n4527 = n568 & ~n4526;
  assign n4528 = n572 & ~n4527;
  assign n4529 = n576 & ~n4528;
  assign n4530 = n580 & ~n4529;
  assign n4531 = n584 & ~n4530;
  assign n4532 = n588 & ~n4531;
  assign n4533 = n592 & ~n4532;
  assign n4534 = n596 & ~n4533;
  assign n4535 = n600 & ~n4534;
  assign n4536 = n604 & ~n4535;
  assign n4537 = n608 & ~n4536;
  assign n4538 = n612 & ~n4537;
  assign n4539 = n616 & ~n4538;
  assign n4540 = n620 & ~n4539;
  assign n4541 = n624 & ~n4540;
  assign n4542 = n628 & ~n4541;
  assign n4543 = n632 & ~n4542;
  assign n4544 = n636 & ~n4543;
  assign n4545 = n640 & ~n4544;
  assign n4546 = n644 & ~n4545;
  assign n4547 = n648 & ~n4546;
  assign n4548 = n652 & ~n4547;
  assign n4549 = n656 & ~n4548;
  assign n4550 = n660 & ~n4549;
  assign n4551 = n664 & ~n4550;
  assign n4552 = n668 & ~n4551;
  assign n4553 = n672 & ~n4552;
  assign n4554 = n676 & ~n4553;
  assign n4555 = n680 & ~n4554;
  assign n4556 = n684 & ~n4555;
  assign n4557 = n688 & ~n4556;
  assign n4558 = n692 & ~n4557;
  assign n4559 = n696 & ~n4558;
  assign n4560 = n700 & ~n4559;
  assign n4561 = n704 & ~n4560;
  assign n4562 = n708 & ~n4561;
  assign n4563 = n712 & ~n4562;
  assign n4564 = n716 & ~n4563;
  assign n4565 = n720 & ~n4564;
  assign n4566 = n1484 & ~n4565;
  assign n4567 = n1486 & ~n4566;
  assign n4568 = n1750 & ~n4567;
  assign n4569 = n731 & ~n4568;
  assign n4570 = n735 & ~n4569;
  assign n4571 = n739 & ~n4570;
  assign n4572 = n743 & ~n4571;
  assign n4573 = n747 & ~n4572;
  assign n4574 = n751 & ~n4573;
  assign n4575 = n755 & ~n4574;
  assign n4576 = n759 & ~n4575;
  assign n4577 = n763 & ~n4576;
  assign n4578 = n767 & ~n4577;
  assign n4579 = n771 & ~n4578;
  assign n4580 = n775 & ~n4579;
  assign n4581 = n779 & ~n4580;
  assign n4582 = n783 & ~n4581;
  assign n4583 = n787 & ~n4582;
  assign n4584 = n791 & ~n4583;
  assign n4585 = n795 & ~n4584;
  assign n4586 = n799 & ~n4585;
  assign n4587 = n803 & ~n4586;
  assign n4588 = n807 & ~n4587;
  assign n4589 = n811 & ~n4588;
  assign n4590 = n815 & ~n4589;
  assign n4591 = n819 & ~n4590;
  assign n4592 = pi167  & ~n821;
  assign po39  = ~n4591 & n4592;
  assign n4594 = n830 & ~n1163;
  assign n4595 = n835 & ~n4594;
  assign n4596 = n839 & ~n4595;
  assign n4597 = n843 & ~n4596;
  assign n4598 = n847 & ~n4597;
  assign n4599 = n851 & ~n4598;
  assign n4600 = n855 & ~n4599;
  assign n4601 = n859 & ~n4600;
  assign n4602 = n863 & ~n4601;
  assign n4603 = n867 & ~n4602;
  assign n4604 = n871 & ~n4603;
  assign n4605 = n875 & ~n4604;
  assign n4606 = n879 & ~n4605;
  assign n4607 = n883 & ~n4606;
  assign n4608 = n887 & ~n4607;
  assign n4609 = n891 & ~n4608;
  assign n4610 = n895 & ~n4609;
  assign n4611 = n899 & ~n4610;
  assign n4612 = n903 & ~n4611;
  assign n4613 = n907 & ~n4612;
  assign n4614 = n911 & ~n4613;
  assign n4615 = n915 & ~n4614;
  assign n4616 = n919 & ~n4615;
  assign n4617 = n923 & ~n4616;
  assign n4618 = n927 & ~n4617;
  assign n4619 = n931 & ~n4618;
  assign n4620 = n935 & ~n4619;
  assign n4621 = n939 & ~n4620;
  assign n4622 = n943 & ~n4621;
  assign n4623 = n947 & ~n4622;
  assign n4624 = n951 & ~n4623;
  assign n4625 = n955 & ~n4624;
  assign n4626 = n959 & ~n4625;
  assign n4627 = n963 & ~n4626;
  assign n4628 = n967 & ~n4627;
  assign n4629 = n971 & ~n4628;
  assign n4630 = n975 & ~n4629;
  assign n4631 = n979 & ~n4630;
  assign n4632 = n983 & ~n4631;
  assign n4633 = n987 & ~n4632;
  assign n4634 = n991 & ~n4633;
  assign n4635 = n995 & ~n4634;
  assign n4636 = n999 & ~n4635;
  assign n4637 = n1003 & ~n4636;
  assign n4638 = n1007 & ~n4637;
  assign n4639 = n1011 & ~n4638;
  assign n4640 = n1015 & ~n4639;
  assign n4641 = n1019 & ~n4640;
  assign n4642 = n1023 & ~n4641;
  assign n4643 = n1027 & ~n4642;
  assign n4644 = n1031 & ~n4643;
  assign n4645 = n1035 & ~n4644;
  assign n4646 = n1039 & ~n4645;
  assign n4647 = n1043 & ~n4646;
  assign n4648 = n1047 & ~n4647;
  assign n4649 = n1051 & ~n4648;
  assign n4650 = n1055 & ~n4649;
  assign n4651 = n1059 & ~n4650;
  assign n4652 = n1574 & ~n4651;
  assign n4653 = n1576 & ~n4652;
  assign n4654 = n1837 & ~n4653;
  assign n4655 = n1068 & ~n4654;
  assign n4656 = n1072 & ~n4655;
  assign n4657 = n1076 & ~n4656;
  assign n4658 = n1080 & ~n4657;
  assign n4659 = n1084 & ~n4658;
  assign n4660 = n1088 & ~n4659;
  assign n4661 = n1092 & ~n4660;
  assign n4662 = n1096 & ~n4661;
  assign n4663 = n1100 & ~n4662;
  assign n4664 = n1104 & ~n4663;
  assign n4665 = n1108 & ~n4664;
  assign n4666 = n1112 & ~n4665;
  assign n4667 = n1116 & ~n4666;
  assign n4668 = n1120 & ~n4667;
  assign n4669 = n1124 & ~n4668;
  assign n4670 = n1128 & ~n4669;
  assign n4671 = n1132 & ~n4670;
  assign n4672 = n1136 & ~n4671;
  assign n4673 = n1140 & ~n4672;
  assign n4674 = n1144 & ~n4673;
  assign n4675 = n1148 & ~n4674;
  assign n4676 = n1152 & ~n4675;
  assign n4677 = n1156 & ~n4676;
  assign n4678 = pi168  & ~n1158;
  assign po40  = ~n4677 & n4678;
  assign n4680 = ~n495 & n1167;
  assign n4681 = n1172 & ~n4680;
  assign n4682 = n1176 & ~n4681;
  assign n4683 = n1180 & ~n4682;
  assign n4684 = n1184 & ~n4683;
  assign n4685 = n1188 & ~n4684;
  assign n4686 = n1192 & ~n4685;
  assign n4687 = n1196 & ~n4686;
  assign n4688 = n1200 & ~n4687;
  assign n4689 = n1204 & ~n4688;
  assign n4690 = n1208 & ~n4689;
  assign n4691 = n1212 & ~n4690;
  assign n4692 = n1216 & ~n4691;
  assign n4693 = n1220 & ~n4692;
  assign n4694 = n1224 & ~n4693;
  assign n4695 = n1228 & ~n4694;
  assign n4696 = n1232 & ~n4695;
  assign n4697 = n1236 & ~n4696;
  assign n4698 = n1240 & ~n4697;
  assign n4699 = n1244 & ~n4698;
  assign n4700 = n1248 & ~n4699;
  assign n4701 = n1252 & ~n4700;
  assign n4702 = n1256 & ~n4701;
  assign n4703 = n1260 & ~n4702;
  assign n4704 = n1264 & ~n4703;
  assign n4705 = n1268 & ~n4704;
  assign n4706 = n1272 & ~n4705;
  assign n4707 = n1276 & ~n4706;
  assign n4708 = n1280 & ~n4707;
  assign n4709 = n1284 & ~n4708;
  assign n4710 = n1288 & ~n4709;
  assign n4711 = n1292 & ~n4710;
  assign n4712 = n1296 & ~n4711;
  assign n4713 = n1300 & ~n4712;
  assign n4714 = n1304 & ~n4713;
  assign n4715 = n1308 & ~n4714;
  assign n4716 = n1312 & ~n4715;
  assign n4717 = n1316 & ~n4716;
  assign n4718 = n1320 & ~n4717;
  assign n4719 = n1324 & ~n4718;
  assign n4720 = n1328 & ~n4719;
  assign n4721 = n1332 & ~n4720;
  assign n4722 = n1336 & ~n4721;
  assign n4723 = n1340 & ~n4722;
  assign n4724 = n1344 & ~n4723;
  assign n4725 = n1348 & ~n4724;
  assign n4726 = n1352 & ~n4725;
  assign n4727 = n1356 & ~n4726;
  assign n4728 = n1360 & ~n4727;
  assign n4729 = n1364 & ~n4728;
  assign n4730 = n1368 & ~n4729;
  assign n4731 = n1372 & ~n4730;
  assign n4732 = n1376 & ~n4731;
  assign n4733 = n1380 & ~n4732;
  assign n4734 = n1384 & ~n4733;
  assign n4735 = n1388 & ~n4734;
  assign n4736 = n1392 & ~n4735;
  assign n4737 = n1396 & ~n4736;
  assign n4738 = n1663 & ~n4737;
  assign n4739 = n392 & ~n4738;
  assign n4740 = n396 & ~n4739;
  assign n4741 = n400 & ~n4740;
  assign n4742 = n404 & ~n4741;
  assign n4743 = n408 & ~n4742;
  assign n4744 = n412 & ~n4743;
  assign n4745 = n416 & ~n4744;
  assign n4746 = n420 & ~n4745;
  assign n4747 = n424 & ~n4746;
  assign n4748 = n428 & ~n4747;
  assign n4749 = n432 & ~n4748;
  assign n4750 = n436 & ~n4749;
  assign n4751 = n440 & ~n4750;
  assign n4752 = n444 & ~n4751;
  assign n4753 = n448 & ~n4752;
  assign n4754 = n452 & ~n4753;
  assign n4755 = n456 & ~n4754;
  assign n4756 = n460 & ~n4755;
  assign n4757 = n464 & ~n4756;
  assign n4758 = n468 & ~n4757;
  assign n4759 = n472 & ~n4758;
  assign n4760 = n476 & ~n4759;
  assign n4761 = n480 & ~n4760;
  assign n4762 = n484 & ~n4761;
  assign n4763 = n488 & ~n4762;
  assign n4764 = pi169  & ~n490;
  assign po41  = ~n4763 & n4764;
  assign n4766 = n499 & ~n834;
  assign n4767 = n504 & ~n4766;
  assign n4768 = n508 & ~n4767;
  assign n4769 = n512 & ~n4768;
  assign n4770 = n516 & ~n4769;
  assign n4771 = n520 & ~n4770;
  assign n4772 = n524 & ~n4771;
  assign n4773 = n528 & ~n4772;
  assign n4774 = n532 & ~n4773;
  assign n4775 = n536 & ~n4774;
  assign n4776 = n540 & ~n4775;
  assign n4777 = n544 & ~n4776;
  assign n4778 = n548 & ~n4777;
  assign n4779 = n552 & ~n4778;
  assign n4780 = n556 & ~n4779;
  assign n4781 = n560 & ~n4780;
  assign n4782 = n564 & ~n4781;
  assign n4783 = n568 & ~n4782;
  assign n4784 = n572 & ~n4783;
  assign n4785 = n576 & ~n4784;
  assign n4786 = n580 & ~n4785;
  assign n4787 = n584 & ~n4786;
  assign n4788 = n588 & ~n4787;
  assign n4789 = n592 & ~n4788;
  assign n4790 = n596 & ~n4789;
  assign n4791 = n600 & ~n4790;
  assign n4792 = n604 & ~n4791;
  assign n4793 = n608 & ~n4792;
  assign n4794 = n612 & ~n4793;
  assign n4795 = n616 & ~n4794;
  assign n4796 = n620 & ~n4795;
  assign n4797 = n624 & ~n4796;
  assign n4798 = n628 & ~n4797;
  assign n4799 = n632 & ~n4798;
  assign n4800 = n636 & ~n4799;
  assign n4801 = n640 & ~n4800;
  assign n4802 = n644 & ~n4801;
  assign n4803 = n648 & ~n4802;
  assign n4804 = n652 & ~n4803;
  assign n4805 = n656 & ~n4804;
  assign n4806 = n660 & ~n4805;
  assign n4807 = n664 & ~n4806;
  assign n4808 = n668 & ~n4807;
  assign n4809 = n672 & ~n4808;
  assign n4810 = n676 & ~n4809;
  assign n4811 = n680 & ~n4810;
  assign n4812 = n684 & ~n4811;
  assign n4813 = n688 & ~n4812;
  assign n4814 = n692 & ~n4813;
  assign n4815 = n696 & ~n4814;
  assign n4816 = n700 & ~n4815;
  assign n4817 = n704 & ~n4816;
  assign n4818 = n708 & ~n4817;
  assign n4819 = n712 & ~n4818;
  assign n4820 = n716 & ~n4819;
  assign n4821 = n720 & ~n4820;
  assign n4822 = n1484 & ~n4821;
  assign n4823 = n1486 & ~n4822;
  assign n4824 = n1750 & ~n4823;
  assign n4825 = n731 & ~n4824;
  assign n4826 = n735 & ~n4825;
  assign n4827 = n739 & ~n4826;
  assign n4828 = n743 & ~n4827;
  assign n4829 = n747 & ~n4828;
  assign n4830 = n751 & ~n4829;
  assign n4831 = n755 & ~n4830;
  assign n4832 = n759 & ~n4831;
  assign n4833 = n763 & ~n4832;
  assign n4834 = n767 & ~n4833;
  assign n4835 = n771 & ~n4834;
  assign n4836 = n775 & ~n4835;
  assign n4837 = n779 & ~n4836;
  assign n4838 = n783 & ~n4837;
  assign n4839 = n787 & ~n4838;
  assign n4840 = n791 & ~n4839;
  assign n4841 = n795 & ~n4840;
  assign n4842 = n799 & ~n4841;
  assign n4843 = n803 & ~n4842;
  assign n4844 = n807 & ~n4843;
  assign n4845 = n811 & ~n4844;
  assign n4846 = n815 & ~n4845;
  assign n4847 = n819 & ~n4846;
  assign n4848 = n823 & ~n4847;
  assign n4849 = n827 & ~n4848;
  assign n4850 = pi170  & ~n829;
  assign po42  = ~n4849 & n4850;
  assign n4852 = n838 & ~n1171;
  assign n4853 = n843 & ~n4852;
  assign n4854 = n847 & ~n4853;
  assign n4855 = n851 & ~n4854;
  assign n4856 = n855 & ~n4855;
  assign n4857 = n859 & ~n4856;
  assign n4858 = n863 & ~n4857;
  assign n4859 = n867 & ~n4858;
  assign n4860 = n871 & ~n4859;
  assign n4861 = n875 & ~n4860;
  assign n4862 = n879 & ~n4861;
  assign n4863 = n883 & ~n4862;
  assign n4864 = n887 & ~n4863;
  assign n4865 = n891 & ~n4864;
  assign n4866 = n895 & ~n4865;
  assign n4867 = n899 & ~n4866;
  assign n4868 = n903 & ~n4867;
  assign n4869 = n907 & ~n4868;
  assign n4870 = n911 & ~n4869;
  assign n4871 = n915 & ~n4870;
  assign n4872 = n919 & ~n4871;
  assign n4873 = n923 & ~n4872;
  assign n4874 = n927 & ~n4873;
  assign n4875 = n931 & ~n4874;
  assign n4876 = n935 & ~n4875;
  assign n4877 = n939 & ~n4876;
  assign n4878 = n943 & ~n4877;
  assign n4879 = n947 & ~n4878;
  assign n4880 = n951 & ~n4879;
  assign n4881 = n955 & ~n4880;
  assign n4882 = n959 & ~n4881;
  assign n4883 = n963 & ~n4882;
  assign n4884 = n967 & ~n4883;
  assign n4885 = n971 & ~n4884;
  assign n4886 = n975 & ~n4885;
  assign n4887 = n979 & ~n4886;
  assign n4888 = n983 & ~n4887;
  assign n4889 = n987 & ~n4888;
  assign n4890 = n991 & ~n4889;
  assign n4891 = n995 & ~n4890;
  assign n4892 = n999 & ~n4891;
  assign n4893 = n1003 & ~n4892;
  assign n4894 = n1007 & ~n4893;
  assign n4895 = n1011 & ~n4894;
  assign n4896 = n1015 & ~n4895;
  assign n4897 = n1019 & ~n4896;
  assign n4898 = n1023 & ~n4897;
  assign n4899 = n1027 & ~n4898;
  assign n4900 = n1031 & ~n4899;
  assign n4901 = n1035 & ~n4900;
  assign n4902 = n1039 & ~n4901;
  assign n4903 = n1043 & ~n4902;
  assign n4904 = n1047 & ~n4903;
  assign n4905 = n1051 & ~n4904;
  assign n4906 = n1055 & ~n4905;
  assign n4907 = n1059 & ~n4906;
  assign n4908 = n1574 & ~n4907;
  assign n4909 = n1576 & ~n4908;
  assign n4910 = n1837 & ~n4909;
  assign n4911 = n1068 & ~n4910;
  assign n4912 = n1072 & ~n4911;
  assign n4913 = n1076 & ~n4912;
  assign n4914 = n1080 & ~n4913;
  assign n4915 = n1084 & ~n4914;
  assign n4916 = n1088 & ~n4915;
  assign n4917 = n1092 & ~n4916;
  assign n4918 = n1096 & ~n4917;
  assign n4919 = n1100 & ~n4918;
  assign n4920 = n1104 & ~n4919;
  assign n4921 = n1108 & ~n4920;
  assign n4922 = n1112 & ~n4921;
  assign n4923 = n1116 & ~n4922;
  assign n4924 = n1120 & ~n4923;
  assign n4925 = n1124 & ~n4924;
  assign n4926 = n1128 & ~n4925;
  assign n4927 = n1132 & ~n4926;
  assign n4928 = n1136 & ~n4927;
  assign n4929 = n1140 & ~n4928;
  assign n4930 = n1144 & ~n4929;
  assign n4931 = n1148 & ~n4930;
  assign n4932 = n1152 & ~n4931;
  assign n4933 = n1156 & ~n4932;
  assign n4934 = n1160 & ~n4933;
  assign n4935 = n1164 & ~n4934;
  assign n4936 = pi171  & ~n1166;
  assign po43  = ~n4935 & n4936;
  assign n4938 = ~n503 & n1175;
  assign n4939 = n1180 & ~n4938;
  assign n4940 = n1184 & ~n4939;
  assign n4941 = n1188 & ~n4940;
  assign n4942 = n1192 & ~n4941;
  assign n4943 = n1196 & ~n4942;
  assign n4944 = n1200 & ~n4943;
  assign n4945 = n1204 & ~n4944;
  assign n4946 = n1208 & ~n4945;
  assign n4947 = n1212 & ~n4946;
  assign n4948 = n1216 & ~n4947;
  assign n4949 = n1220 & ~n4948;
  assign n4950 = n1224 & ~n4949;
  assign n4951 = n1228 & ~n4950;
  assign n4952 = n1232 & ~n4951;
  assign n4953 = n1236 & ~n4952;
  assign n4954 = n1240 & ~n4953;
  assign n4955 = n1244 & ~n4954;
  assign n4956 = n1248 & ~n4955;
  assign n4957 = n1252 & ~n4956;
  assign n4958 = n1256 & ~n4957;
  assign n4959 = n1260 & ~n4958;
  assign n4960 = n1264 & ~n4959;
  assign n4961 = n1268 & ~n4960;
  assign n4962 = n1272 & ~n4961;
  assign n4963 = n1276 & ~n4962;
  assign n4964 = n1280 & ~n4963;
  assign n4965 = n1284 & ~n4964;
  assign n4966 = n1288 & ~n4965;
  assign n4967 = n1292 & ~n4966;
  assign n4968 = n1296 & ~n4967;
  assign n4969 = n1300 & ~n4968;
  assign n4970 = n1304 & ~n4969;
  assign n4971 = n1308 & ~n4970;
  assign n4972 = n1312 & ~n4971;
  assign n4973 = n1316 & ~n4972;
  assign n4974 = n1320 & ~n4973;
  assign n4975 = n1324 & ~n4974;
  assign n4976 = n1328 & ~n4975;
  assign n4977 = n1332 & ~n4976;
  assign n4978 = n1336 & ~n4977;
  assign n4979 = n1340 & ~n4978;
  assign n4980 = n1344 & ~n4979;
  assign n4981 = n1348 & ~n4980;
  assign n4982 = n1352 & ~n4981;
  assign n4983 = n1356 & ~n4982;
  assign n4984 = n1360 & ~n4983;
  assign n4985 = n1364 & ~n4984;
  assign n4986 = n1368 & ~n4985;
  assign n4987 = n1372 & ~n4986;
  assign n4988 = n1376 & ~n4987;
  assign n4989 = n1380 & ~n4988;
  assign n4990 = n1384 & ~n4989;
  assign n4991 = n1388 & ~n4990;
  assign n4992 = n1392 & ~n4991;
  assign n4993 = n1396 & ~n4992;
  assign n4994 = n1663 & ~n4993;
  assign n4995 = n392 & ~n4994;
  assign n4996 = n396 & ~n4995;
  assign n4997 = n400 & ~n4996;
  assign n4998 = n404 & ~n4997;
  assign n4999 = n408 & ~n4998;
  assign n5000 = n412 & ~n4999;
  assign n5001 = n416 & ~n5000;
  assign n5002 = n420 & ~n5001;
  assign n5003 = n424 & ~n5002;
  assign n5004 = n428 & ~n5003;
  assign n5005 = n432 & ~n5004;
  assign n5006 = n436 & ~n5005;
  assign n5007 = n440 & ~n5006;
  assign n5008 = n444 & ~n5007;
  assign n5009 = n448 & ~n5008;
  assign n5010 = n452 & ~n5009;
  assign n5011 = n456 & ~n5010;
  assign n5012 = n460 & ~n5011;
  assign n5013 = n464 & ~n5012;
  assign n5014 = n468 & ~n5013;
  assign n5015 = n472 & ~n5014;
  assign n5016 = n476 & ~n5015;
  assign n5017 = n480 & ~n5016;
  assign n5018 = n484 & ~n5017;
  assign n5019 = n488 & ~n5018;
  assign n5020 = n492 & ~n5019;
  assign n5021 = n496 & ~n5020;
  assign n5022 = pi172  & ~n498;
  assign po44  = ~n5021 & n5022;
  assign n5024 = n507 & ~n842;
  assign n5025 = n512 & ~n5024;
  assign n5026 = n516 & ~n5025;
  assign n5027 = n520 & ~n5026;
  assign n5028 = n524 & ~n5027;
  assign n5029 = n528 & ~n5028;
  assign n5030 = n532 & ~n5029;
  assign n5031 = n536 & ~n5030;
  assign n5032 = n540 & ~n5031;
  assign n5033 = n544 & ~n5032;
  assign n5034 = n548 & ~n5033;
  assign n5035 = n552 & ~n5034;
  assign n5036 = n556 & ~n5035;
  assign n5037 = n560 & ~n5036;
  assign n5038 = n564 & ~n5037;
  assign n5039 = n568 & ~n5038;
  assign n5040 = n572 & ~n5039;
  assign n5041 = n576 & ~n5040;
  assign n5042 = n580 & ~n5041;
  assign n5043 = n584 & ~n5042;
  assign n5044 = n588 & ~n5043;
  assign n5045 = n592 & ~n5044;
  assign n5046 = n596 & ~n5045;
  assign n5047 = n600 & ~n5046;
  assign n5048 = n604 & ~n5047;
  assign n5049 = n608 & ~n5048;
  assign n5050 = n612 & ~n5049;
  assign n5051 = n616 & ~n5050;
  assign n5052 = n620 & ~n5051;
  assign n5053 = n624 & ~n5052;
  assign n5054 = n628 & ~n5053;
  assign n5055 = n632 & ~n5054;
  assign n5056 = n636 & ~n5055;
  assign n5057 = n640 & ~n5056;
  assign n5058 = n644 & ~n5057;
  assign n5059 = n648 & ~n5058;
  assign n5060 = n652 & ~n5059;
  assign n5061 = n656 & ~n5060;
  assign n5062 = n660 & ~n5061;
  assign n5063 = n664 & ~n5062;
  assign n5064 = n668 & ~n5063;
  assign n5065 = n672 & ~n5064;
  assign n5066 = n676 & ~n5065;
  assign n5067 = n680 & ~n5066;
  assign n5068 = n684 & ~n5067;
  assign n5069 = n688 & ~n5068;
  assign n5070 = n692 & ~n5069;
  assign n5071 = n696 & ~n5070;
  assign n5072 = n700 & ~n5071;
  assign n5073 = n704 & ~n5072;
  assign n5074 = n708 & ~n5073;
  assign n5075 = n712 & ~n5074;
  assign n5076 = n716 & ~n5075;
  assign n5077 = n720 & ~n5076;
  assign n5078 = n1484 & ~n5077;
  assign n5079 = n1486 & ~n5078;
  assign n5080 = n1750 & ~n5079;
  assign n5081 = n731 & ~n5080;
  assign n5082 = n735 & ~n5081;
  assign n5083 = n739 & ~n5082;
  assign n5084 = n743 & ~n5083;
  assign n5085 = n747 & ~n5084;
  assign n5086 = n751 & ~n5085;
  assign n5087 = n755 & ~n5086;
  assign n5088 = n759 & ~n5087;
  assign n5089 = n763 & ~n5088;
  assign n5090 = n767 & ~n5089;
  assign n5091 = n771 & ~n5090;
  assign n5092 = n775 & ~n5091;
  assign n5093 = n779 & ~n5092;
  assign n5094 = n783 & ~n5093;
  assign n5095 = n787 & ~n5094;
  assign n5096 = n791 & ~n5095;
  assign n5097 = n795 & ~n5096;
  assign n5098 = n799 & ~n5097;
  assign n5099 = n803 & ~n5098;
  assign n5100 = n807 & ~n5099;
  assign n5101 = n811 & ~n5100;
  assign n5102 = n815 & ~n5101;
  assign n5103 = n819 & ~n5102;
  assign n5104 = n823 & ~n5103;
  assign n5105 = n827 & ~n5104;
  assign n5106 = n831 & ~n5105;
  assign n5107 = n835 & ~n5106;
  assign n5108 = pi173  & ~n837;
  assign po45  = ~n5107 & n5108;
  assign n5110 = n846 & ~n1179;
  assign n5111 = n851 & ~n5110;
  assign n5112 = n855 & ~n5111;
  assign n5113 = n859 & ~n5112;
  assign n5114 = n863 & ~n5113;
  assign n5115 = n867 & ~n5114;
  assign n5116 = n871 & ~n5115;
  assign n5117 = n875 & ~n5116;
  assign n5118 = n879 & ~n5117;
  assign n5119 = n883 & ~n5118;
  assign n5120 = n887 & ~n5119;
  assign n5121 = n891 & ~n5120;
  assign n5122 = n895 & ~n5121;
  assign n5123 = n899 & ~n5122;
  assign n5124 = n903 & ~n5123;
  assign n5125 = n907 & ~n5124;
  assign n5126 = n911 & ~n5125;
  assign n5127 = n915 & ~n5126;
  assign n5128 = n919 & ~n5127;
  assign n5129 = n923 & ~n5128;
  assign n5130 = n927 & ~n5129;
  assign n5131 = n931 & ~n5130;
  assign n5132 = n935 & ~n5131;
  assign n5133 = n939 & ~n5132;
  assign n5134 = n943 & ~n5133;
  assign n5135 = n947 & ~n5134;
  assign n5136 = n951 & ~n5135;
  assign n5137 = n955 & ~n5136;
  assign n5138 = n959 & ~n5137;
  assign n5139 = n963 & ~n5138;
  assign n5140 = n967 & ~n5139;
  assign n5141 = n971 & ~n5140;
  assign n5142 = n975 & ~n5141;
  assign n5143 = n979 & ~n5142;
  assign n5144 = n983 & ~n5143;
  assign n5145 = n987 & ~n5144;
  assign n5146 = n991 & ~n5145;
  assign n5147 = n995 & ~n5146;
  assign n5148 = n999 & ~n5147;
  assign n5149 = n1003 & ~n5148;
  assign n5150 = n1007 & ~n5149;
  assign n5151 = n1011 & ~n5150;
  assign n5152 = n1015 & ~n5151;
  assign n5153 = n1019 & ~n5152;
  assign n5154 = n1023 & ~n5153;
  assign n5155 = n1027 & ~n5154;
  assign n5156 = n1031 & ~n5155;
  assign n5157 = n1035 & ~n5156;
  assign n5158 = n1039 & ~n5157;
  assign n5159 = n1043 & ~n5158;
  assign n5160 = n1047 & ~n5159;
  assign n5161 = n1051 & ~n5160;
  assign n5162 = n1055 & ~n5161;
  assign n5163 = n1059 & ~n5162;
  assign n5164 = n1574 & ~n5163;
  assign n5165 = n1576 & ~n5164;
  assign n5166 = n1837 & ~n5165;
  assign n5167 = n1068 & ~n5166;
  assign n5168 = n1072 & ~n5167;
  assign n5169 = n1076 & ~n5168;
  assign n5170 = n1080 & ~n5169;
  assign n5171 = n1084 & ~n5170;
  assign n5172 = n1088 & ~n5171;
  assign n5173 = n1092 & ~n5172;
  assign n5174 = n1096 & ~n5173;
  assign n5175 = n1100 & ~n5174;
  assign n5176 = n1104 & ~n5175;
  assign n5177 = n1108 & ~n5176;
  assign n5178 = n1112 & ~n5177;
  assign n5179 = n1116 & ~n5178;
  assign n5180 = n1120 & ~n5179;
  assign n5181 = n1124 & ~n5180;
  assign n5182 = n1128 & ~n5181;
  assign n5183 = n1132 & ~n5182;
  assign n5184 = n1136 & ~n5183;
  assign n5185 = n1140 & ~n5184;
  assign n5186 = n1144 & ~n5185;
  assign n5187 = n1148 & ~n5186;
  assign n5188 = n1152 & ~n5187;
  assign n5189 = n1156 & ~n5188;
  assign n5190 = n1160 & ~n5189;
  assign n5191 = n1164 & ~n5190;
  assign n5192 = n1168 & ~n5191;
  assign n5193 = n1172 & ~n5192;
  assign n5194 = pi174  & ~n1174;
  assign po46  = ~n5193 & n5194;
  assign n5196 = ~n511 & n1183;
  assign n5197 = n1188 & ~n5196;
  assign n5198 = n1192 & ~n5197;
  assign n5199 = n1196 & ~n5198;
  assign n5200 = n1200 & ~n5199;
  assign n5201 = n1204 & ~n5200;
  assign n5202 = n1208 & ~n5201;
  assign n5203 = n1212 & ~n5202;
  assign n5204 = n1216 & ~n5203;
  assign n5205 = n1220 & ~n5204;
  assign n5206 = n1224 & ~n5205;
  assign n5207 = n1228 & ~n5206;
  assign n5208 = n1232 & ~n5207;
  assign n5209 = n1236 & ~n5208;
  assign n5210 = n1240 & ~n5209;
  assign n5211 = n1244 & ~n5210;
  assign n5212 = n1248 & ~n5211;
  assign n5213 = n1252 & ~n5212;
  assign n5214 = n1256 & ~n5213;
  assign n5215 = n1260 & ~n5214;
  assign n5216 = n1264 & ~n5215;
  assign n5217 = n1268 & ~n5216;
  assign n5218 = n1272 & ~n5217;
  assign n5219 = n1276 & ~n5218;
  assign n5220 = n1280 & ~n5219;
  assign n5221 = n1284 & ~n5220;
  assign n5222 = n1288 & ~n5221;
  assign n5223 = n1292 & ~n5222;
  assign n5224 = n1296 & ~n5223;
  assign n5225 = n1300 & ~n5224;
  assign n5226 = n1304 & ~n5225;
  assign n5227 = n1308 & ~n5226;
  assign n5228 = n1312 & ~n5227;
  assign n5229 = n1316 & ~n5228;
  assign n5230 = n1320 & ~n5229;
  assign n5231 = n1324 & ~n5230;
  assign n5232 = n1328 & ~n5231;
  assign n5233 = n1332 & ~n5232;
  assign n5234 = n1336 & ~n5233;
  assign n5235 = n1340 & ~n5234;
  assign n5236 = n1344 & ~n5235;
  assign n5237 = n1348 & ~n5236;
  assign n5238 = n1352 & ~n5237;
  assign n5239 = n1356 & ~n5238;
  assign n5240 = n1360 & ~n5239;
  assign n5241 = n1364 & ~n5240;
  assign n5242 = n1368 & ~n5241;
  assign n5243 = n1372 & ~n5242;
  assign n5244 = n1376 & ~n5243;
  assign n5245 = n1380 & ~n5244;
  assign n5246 = n1384 & ~n5245;
  assign n5247 = n1388 & ~n5246;
  assign n5248 = n1392 & ~n5247;
  assign n5249 = n1396 & ~n5248;
  assign n5250 = n1663 & ~n5249;
  assign n5251 = n392 & ~n5250;
  assign n5252 = n396 & ~n5251;
  assign n5253 = n400 & ~n5252;
  assign n5254 = n404 & ~n5253;
  assign n5255 = n408 & ~n5254;
  assign n5256 = n412 & ~n5255;
  assign n5257 = n416 & ~n5256;
  assign n5258 = n420 & ~n5257;
  assign n5259 = n424 & ~n5258;
  assign n5260 = n428 & ~n5259;
  assign n5261 = n432 & ~n5260;
  assign n5262 = n436 & ~n5261;
  assign n5263 = n440 & ~n5262;
  assign n5264 = n444 & ~n5263;
  assign n5265 = n448 & ~n5264;
  assign n5266 = n452 & ~n5265;
  assign n5267 = n456 & ~n5266;
  assign n5268 = n460 & ~n5267;
  assign n5269 = n464 & ~n5268;
  assign n5270 = n468 & ~n5269;
  assign n5271 = n472 & ~n5270;
  assign n5272 = n476 & ~n5271;
  assign n5273 = n480 & ~n5272;
  assign n5274 = n484 & ~n5273;
  assign n5275 = n488 & ~n5274;
  assign n5276 = n492 & ~n5275;
  assign n5277 = n496 & ~n5276;
  assign n5278 = n500 & ~n5277;
  assign n5279 = n504 & ~n5278;
  assign n5280 = pi175  & ~n506;
  assign po47  = ~n5279 & n5280;
  assign n5282 = n515 & ~n850;
  assign n5283 = n520 & ~n5282;
  assign n5284 = n524 & ~n5283;
  assign n5285 = n528 & ~n5284;
  assign n5286 = n532 & ~n5285;
  assign n5287 = n536 & ~n5286;
  assign n5288 = n540 & ~n5287;
  assign n5289 = n544 & ~n5288;
  assign n5290 = n548 & ~n5289;
  assign n5291 = n552 & ~n5290;
  assign n5292 = n556 & ~n5291;
  assign n5293 = n560 & ~n5292;
  assign n5294 = n564 & ~n5293;
  assign n5295 = n568 & ~n5294;
  assign n5296 = n572 & ~n5295;
  assign n5297 = n576 & ~n5296;
  assign n5298 = n580 & ~n5297;
  assign n5299 = n584 & ~n5298;
  assign n5300 = n588 & ~n5299;
  assign n5301 = n592 & ~n5300;
  assign n5302 = n596 & ~n5301;
  assign n5303 = n600 & ~n5302;
  assign n5304 = n604 & ~n5303;
  assign n5305 = n608 & ~n5304;
  assign n5306 = n612 & ~n5305;
  assign n5307 = n616 & ~n5306;
  assign n5308 = n620 & ~n5307;
  assign n5309 = n624 & ~n5308;
  assign n5310 = n628 & ~n5309;
  assign n5311 = n632 & ~n5310;
  assign n5312 = n636 & ~n5311;
  assign n5313 = n640 & ~n5312;
  assign n5314 = n644 & ~n5313;
  assign n5315 = n648 & ~n5314;
  assign n5316 = n652 & ~n5315;
  assign n5317 = n656 & ~n5316;
  assign n5318 = n660 & ~n5317;
  assign n5319 = n664 & ~n5318;
  assign n5320 = n668 & ~n5319;
  assign n5321 = n672 & ~n5320;
  assign n5322 = n676 & ~n5321;
  assign n5323 = n680 & ~n5322;
  assign n5324 = n684 & ~n5323;
  assign n5325 = n688 & ~n5324;
  assign n5326 = n692 & ~n5325;
  assign n5327 = n696 & ~n5326;
  assign n5328 = n700 & ~n5327;
  assign n5329 = n704 & ~n5328;
  assign n5330 = n708 & ~n5329;
  assign n5331 = n712 & ~n5330;
  assign n5332 = n716 & ~n5331;
  assign n5333 = n720 & ~n5332;
  assign n5334 = n1484 & ~n5333;
  assign n5335 = n1486 & ~n5334;
  assign n5336 = n1750 & ~n5335;
  assign n5337 = n731 & ~n5336;
  assign n5338 = n735 & ~n5337;
  assign n5339 = n739 & ~n5338;
  assign n5340 = n743 & ~n5339;
  assign n5341 = n747 & ~n5340;
  assign n5342 = n751 & ~n5341;
  assign n5343 = n755 & ~n5342;
  assign n5344 = n759 & ~n5343;
  assign n5345 = n763 & ~n5344;
  assign n5346 = n767 & ~n5345;
  assign n5347 = n771 & ~n5346;
  assign n5348 = n775 & ~n5347;
  assign n5349 = n779 & ~n5348;
  assign n5350 = n783 & ~n5349;
  assign n5351 = n787 & ~n5350;
  assign n5352 = n791 & ~n5351;
  assign n5353 = n795 & ~n5352;
  assign n5354 = n799 & ~n5353;
  assign n5355 = n803 & ~n5354;
  assign n5356 = n807 & ~n5355;
  assign n5357 = n811 & ~n5356;
  assign n5358 = n815 & ~n5357;
  assign n5359 = n819 & ~n5358;
  assign n5360 = n823 & ~n5359;
  assign n5361 = n827 & ~n5360;
  assign n5362 = n831 & ~n5361;
  assign n5363 = n835 & ~n5362;
  assign n5364 = n839 & ~n5363;
  assign n5365 = n843 & ~n5364;
  assign n5366 = pi176  & ~n845;
  assign po48  = ~n5365 & n5366;
  assign n5368 = n854 & ~n1187;
  assign n5369 = n859 & ~n5368;
  assign n5370 = n863 & ~n5369;
  assign n5371 = n867 & ~n5370;
  assign n5372 = n871 & ~n5371;
  assign n5373 = n875 & ~n5372;
  assign n5374 = n879 & ~n5373;
  assign n5375 = n883 & ~n5374;
  assign n5376 = n887 & ~n5375;
  assign n5377 = n891 & ~n5376;
  assign n5378 = n895 & ~n5377;
  assign n5379 = n899 & ~n5378;
  assign n5380 = n903 & ~n5379;
  assign n5381 = n907 & ~n5380;
  assign n5382 = n911 & ~n5381;
  assign n5383 = n915 & ~n5382;
  assign n5384 = n919 & ~n5383;
  assign n5385 = n923 & ~n5384;
  assign n5386 = n927 & ~n5385;
  assign n5387 = n931 & ~n5386;
  assign n5388 = n935 & ~n5387;
  assign n5389 = n939 & ~n5388;
  assign n5390 = n943 & ~n5389;
  assign n5391 = n947 & ~n5390;
  assign n5392 = n951 & ~n5391;
  assign n5393 = n955 & ~n5392;
  assign n5394 = n959 & ~n5393;
  assign n5395 = n963 & ~n5394;
  assign n5396 = n967 & ~n5395;
  assign n5397 = n971 & ~n5396;
  assign n5398 = n975 & ~n5397;
  assign n5399 = n979 & ~n5398;
  assign n5400 = n983 & ~n5399;
  assign n5401 = n987 & ~n5400;
  assign n5402 = n991 & ~n5401;
  assign n5403 = n995 & ~n5402;
  assign n5404 = n999 & ~n5403;
  assign n5405 = n1003 & ~n5404;
  assign n5406 = n1007 & ~n5405;
  assign n5407 = n1011 & ~n5406;
  assign n5408 = n1015 & ~n5407;
  assign n5409 = n1019 & ~n5408;
  assign n5410 = n1023 & ~n5409;
  assign n5411 = n1027 & ~n5410;
  assign n5412 = n1031 & ~n5411;
  assign n5413 = n1035 & ~n5412;
  assign n5414 = n1039 & ~n5413;
  assign n5415 = n1043 & ~n5414;
  assign n5416 = n1047 & ~n5415;
  assign n5417 = n1051 & ~n5416;
  assign n5418 = n1055 & ~n5417;
  assign n5419 = n1059 & ~n5418;
  assign n5420 = n1574 & ~n5419;
  assign n5421 = n1576 & ~n5420;
  assign n5422 = n1837 & ~n5421;
  assign n5423 = n1068 & ~n5422;
  assign n5424 = n1072 & ~n5423;
  assign n5425 = n1076 & ~n5424;
  assign n5426 = n1080 & ~n5425;
  assign n5427 = n1084 & ~n5426;
  assign n5428 = n1088 & ~n5427;
  assign n5429 = n1092 & ~n5428;
  assign n5430 = n1096 & ~n5429;
  assign n5431 = n1100 & ~n5430;
  assign n5432 = n1104 & ~n5431;
  assign n5433 = n1108 & ~n5432;
  assign n5434 = n1112 & ~n5433;
  assign n5435 = n1116 & ~n5434;
  assign n5436 = n1120 & ~n5435;
  assign n5437 = n1124 & ~n5436;
  assign n5438 = n1128 & ~n5437;
  assign n5439 = n1132 & ~n5438;
  assign n5440 = n1136 & ~n5439;
  assign n5441 = n1140 & ~n5440;
  assign n5442 = n1144 & ~n5441;
  assign n5443 = n1148 & ~n5442;
  assign n5444 = n1152 & ~n5443;
  assign n5445 = n1156 & ~n5444;
  assign n5446 = n1160 & ~n5445;
  assign n5447 = n1164 & ~n5446;
  assign n5448 = n1168 & ~n5447;
  assign n5449 = n1172 & ~n5448;
  assign n5450 = n1176 & ~n5449;
  assign n5451 = n1180 & ~n5450;
  assign n5452 = pi177  & ~n1182;
  assign po49  = ~n5451 & n5452;
  assign n5454 = ~n519 & n1191;
  assign n5455 = n1196 & ~n5454;
  assign n5456 = n1200 & ~n5455;
  assign n5457 = n1204 & ~n5456;
  assign n5458 = n1208 & ~n5457;
  assign n5459 = n1212 & ~n5458;
  assign n5460 = n1216 & ~n5459;
  assign n5461 = n1220 & ~n5460;
  assign n5462 = n1224 & ~n5461;
  assign n5463 = n1228 & ~n5462;
  assign n5464 = n1232 & ~n5463;
  assign n5465 = n1236 & ~n5464;
  assign n5466 = n1240 & ~n5465;
  assign n5467 = n1244 & ~n5466;
  assign n5468 = n1248 & ~n5467;
  assign n5469 = n1252 & ~n5468;
  assign n5470 = n1256 & ~n5469;
  assign n5471 = n1260 & ~n5470;
  assign n5472 = n1264 & ~n5471;
  assign n5473 = n1268 & ~n5472;
  assign n5474 = n1272 & ~n5473;
  assign n5475 = n1276 & ~n5474;
  assign n5476 = n1280 & ~n5475;
  assign n5477 = n1284 & ~n5476;
  assign n5478 = n1288 & ~n5477;
  assign n5479 = n1292 & ~n5478;
  assign n5480 = n1296 & ~n5479;
  assign n5481 = n1300 & ~n5480;
  assign n5482 = n1304 & ~n5481;
  assign n5483 = n1308 & ~n5482;
  assign n5484 = n1312 & ~n5483;
  assign n5485 = n1316 & ~n5484;
  assign n5486 = n1320 & ~n5485;
  assign n5487 = n1324 & ~n5486;
  assign n5488 = n1328 & ~n5487;
  assign n5489 = n1332 & ~n5488;
  assign n5490 = n1336 & ~n5489;
  assign n5491 = n1340 & ~n5490;
  assign n5492 = n1344 & ~n5491;
  assign n5493 = n1348 & ~n5492;
  assign n5494 = n1352 & ~n5493;
  assign n5495 = n1356 & ~n5494;
  assign n5496 = n1360 & ~n5495;
  assign n5497 = n1364 & ~n5496;
  assign n5498 = n1368 & ~n5497;
  assign n5499 = n1372 & ~n5498;
  assign n5500 = n1376 & ~n5499;
  assign n5501 = n1380 & ~n5500;
  assign n5502 = n1384 & ~n5501;
  assign n5503 = n1388 & ~n5502;
  assign n5504 = n1392 & ~n5503;
  assign n5505 = n1396 & ~n5504;
  assign n5506 = n1663 & ~n5505;
  assign n5507 = n392 & ~n5506;
  assign n5508 = n396 & ~n5507;
  assign n5509 = n400 & ~n5508;
  assign n5510 = n404 & ~n5509;
  assign n5511 = n408 & ~n5510;
  assign n5512 = n412 & ~n5511;
  assign n5513 = n416 & ~n5512;
  assign n5514 = n420 & ~n5513;
  assign n5515 = n424 & ~n5514;
  assign n5516 = n428 & ~n5515;
  assign n5517 = n432 & ~n5516;
  assign n5518 = n436 & ~n5517;
  assign n5519 = n440 & ~n5518;
  assign n5520 = n444 & ~n5519;
  assign n5521 = n448 & ~n5520;
  assign n5522 = n452 & ~n5521;
  assign n5523 = n456 & ~n5522;
  assign n5524 = n460 & ~n5523;
  assign n5525 = n464 & ~n5524;
  assign n5526 = n468 & ~n5525;
  assign n5527 = n472 & ~n5526;
  assign n5528 = n476 & ~n5527;
  assign n5529 = n480 & ~n5528;
  assign n5530 = n484 & ~n5529;
  assign n5531 = n488 & ~n5530;
  assign n5532 = n492 & ~n5531;
  assign n5533 = n496 & ~n5532;
  assign n5534 = n500 & ~n5533;
  assign n5535 = n504 & ~n5534;
  assign n5536 = n508 & ~n5535;
  assign n5537 = n512 & ~n5536;
  assign n5538 = pi178  & ~n514;
  assign po50  = ~n5537 & n5538;
  assign n5540 = n523 & ~n858;
  assign n5541 = n528 & ~n5540;
  assign n5542 = n532 & ~n5541;
  assign n5543 = n536 & ~n5542;
  assign n5544 = n540 & ~n5543;
  assign n5545 = n544 & ~n5544;
  assign n5546 = n548 & ~n5545;
  assign n5547 = n552 & ~n5546;
  assign n5548 = n556 & ~n5547;
  assign n5549 = n560 & ~n5548;
  assign n5550 = n564 & ~n5549;
  assign n5551 = n568 & ~n5550;
  assign n5552 = n572 & ~n5551;
  assign n5553 = n576 & ~n5552;
  assign n5554 = n580 & ~n5553;
  assign n5555 = n584 & ~n5554;
  assign n5556 = n588 & ~n5555;
  assign n5557 = n592 & ~n5556;
  assign n5558 = n596 & ~n5557;
  assign n5559 = n600 & ~n5558;
  assign n5560 = n604 & ~n5559;
  assign n5561 = n608 & ~n5560;
  assign n5562 = n612 & ~n5561;
  assign n5563 = n616 & ~n5562;
  assign n5564 = n620 & ~n5563;
  assign n5565 = n624 & ~n5564;
  assign n5566 = n628 & ~n5565;
  assign n5567 = n632 & ~n5566;
  assign n5568 = n636 & ~n5567;
  assign n5569 = n640 & ~n5568;
  assign n5570 = n644 & ~n5569;
  assign n5571 = n648 & ~n5570;
  assign n5572 = n652 & ~n5571;
  assign n5573 = n656 & ~n5572;
  assign n5574 = n660 & ~n5573;
  assign n5575 = n664 & ~n5574;
  assign n5576 = n668 & ~n5575;
  assign n5577 = n672 & ~n5576;
  assign n5578 = n676 & ~n5577;
  assign n5579 = n680 & ~n5578;
  assign n5580 = n684 & ~n5579;
  assign n5581 = n688 & ~n5580;
  assign n5582 = n692 & ~n5581;
  assign n5583 = n696 & ~n5582;
  assign n5584 = n700 & ~n5583;
  assign n5585 = n704 & ~n5584;
  assign n5586 = n708 & ~n5585;
  assign n5587 = n712 & ~n5586;
  assign n5588 = n716 & ~n5587;
  assign n5589 = n720 & ~n5588;
  assign n5590 = n1484 & ~n5589;
  assign n5591 = n1486 & ~n5590;
  assign n5592 = n1750 & ~n5591;
  assign n5593 = n731 & ~n5592;
  assign n5594 = n735 & ~n5593;
  assign n5595 = n739 & ~n5594;
  assign n5596 = n743 & ~n5595;
  assign n5597 = n747 & ~n5596;
  assign n5598 = n751 & ~n5597;
  assign n5599 = n755 & ~n5598;
  assign n5600 = n759 & ~n5599;
  assign n5601 = n763 & ~n5600;
  assign n5602 = n767 & ~n5601;
  assign n5603 = n771 & ~n5602;
  assign n5604 = n775 & ~n5603;
  assign n5605 = n779 & ~n5604;
  assign n5606 = n783 & ~n5605;
  assign n5607 = n787 & ~n5606;
  assign n5608 = n791 & ~n5607;
  assign n5609 = n795 & ~n5608;
  assign n5610 = n799 & ~n5609;
  assign n5611 = n803 & ~n5610;
  assign n5612 = n807 & ~n5611;
  assign n5613 = n811 & ~n5612;
  assign n5614 = n815 & ~n5613;
  assign n5615 = n819 & ~n5614;
  assign n5616 = n823 & ~n5615;
  assign n5617 = n827 & ~n5616;
  assign n5618 = n831 & ~n5617;
  assign n5619 = n835 & ~n5618;
  assign n5620 = n839 & ~n5619;
  assign n5621 = n843 & ~n5620;
  assign n5622 = n847 & ~n5621;
  assign n5623 = n851 & ~n5622;
  assign n5624 = pi179  & ~n853;
  assign po51  = ~n5623 & n5624;
  assign n5626 = n862 & ~n1195;
  assign n5627 = n867 & ~n5626;
  assign n5628 = n871 & ~n5627;
  assign n5629 = n875 & ~n5628;
  assign n5630 = n879 & ~n5629;
  assign n5631 = n883 & ~n5630;
  assign n5632 = n887 & ~n5631;
  assign n5633 = n891 & ~n5632;
  assign n5634 = n895 & ~n5633;
  assign n5635 = n899 & ~n5634;
  assign n5636 = n903 & ~n5635;
  assign n5637 = n907 & ~n5636;
  assign n5638 = n911 & ~n5637;
  assign n5639 = n915 & ~n5638;
  assign n5640 = n919 & ~n5639;
  assign n5641 = n923 & ~n5640;
  assign n5642 = n927 & ~n5641;
  assign n5643 = n931 & ~n5642;
  assign n5644 = n935 & ~n5643;
  assign n5645 = n939 & ~n5644;
  assign n5646 = n943 & ~n5645;
  assign n5647 = n947 & ~n5646;
  assign n5648 = n951 & ~n5647;
  assign n5649 = n955 & ~n5648;
  assign n5650 = n959 & ~n5649;
  assign n5651 = n963 & ~n5650;
  assign n5652 = n967 & ~n5651;
  assign n5653 = n971 & ~n5652;
  assign n5654 = n975 & ~n5653;
  assign n5655 = n979 & ~n5654;
  assign n5656 = n983 & ~n5655;
  assign n5657 = n987 & ~n5656;
  assign n5658 = n991 & ~n5657;
  assign n5659 = n995 & ~n5658;
  assign n5660 = n999 & ~n5659;
  assign n5661 = n1003 & ~n5660;
  assign n5662 = n1007 & ~n5661;
  assign n5663 = n1011 & ~n5662;
  assign n5664 = n1015 & ~n5663;
  assign n5665 = n1019 & ~n5664;
  assign n5666 = n1023 & ~n5665;
  assign n5667 = n1027 & ~n5666;
  assign n5668 = n1031 & ~n5667;
  assign n5669 = n1035 & ~n5668;
  assign n5670 = n1039 & ~n5669;
  assign n5671 = n1043 & ~n5670;
  assign n5672 = n1047 & ~n5671;
  assign n5673 = n1051 & ~n5672;
  assign n5674 = n1055 & ~n5673;
  assign n5675 = n1059 & ~n5674;
  assign n5676 = n1574 & ~n5675;
  assign n5677 = n1576 & ~n5676;
  assign n5678 = n1837 & ~n5677;
  assign n5679 = n1068 & ~n5678;
  assign n5680 = n1072 & ~n5679;
  assign n5681 = n1076 & ~n5680;
  assign n5682 = n1080 & ~n5681;
  assign n5683 = n1084 & ~n5682;
  assign n5684 = n1088 & ~n5683;
  assign n5685 = n1092 & ~n5684;
  assign n5686 = n1096 & ~n5685;
  assign n5687 = n1100 & ~n5686;
  assign n5688 = n1104 & ~n5687;
  assign n5689 = n1108 & ~n5688;
  assign n5690 = n1112 & ~n5689;
  assign n5691 = n1116 & ~n5690;
  assign n5692 = n1120 & ~n5691;
  assign n5693 = n1124 & ~n5692;
  assign n5694 = n1128 & ~n5693;
  assign n5695 = n1132 & ~n5694;
  assign n5696 = n1136 & ~n5695;
  assign n5697 = n1140 & ~n5696;
  assign n5698 = n1144 & ~n5697;
  assign n5699 = n1148 & ~n5698;
  assign n5700 = n1152 & ~n5699;
  assign n5701 = n1156 & ~n5700;
  assign n5702 = n1160 & ~n5701;
  assign n5703 = n1164 & ~n5702;
  assign n5704 = n1168 & ~n5703;
  assign n5705 = n1172 & ~n5704;
  assign n5706 = n1176 & ~n5705;
  assign n5707 = n1180 & ~n5706;
  assign n5708 = n1184 & ~n5707;
  assign n5709 = n1188 & ~n5708;
  assign n5710 = pi180  & ~n1190;
  assign po52  = ~n5709 & n5710;
  assign n5712 = ~n527 & n1199;
  assign n5713 = n1204 & ~n5712;
  assign n5714 = n1208 & ~n5713;
  assign n5715 = n1212 & ~n5714;
  assign n5716 = n1216 & ~n5715;
  assign n5717 = n1220 & ~n5716;
  assign n5718 = n1224 & ~n5717;
  assign n5719 = n1228 & ~n5718;
  assign n5720 = n1232 & ~n5719;
  assign n5721 = n1236 & ~n5720;
  assign n5722 = n1240 & ~n5721;
  assign n5723 = n1244 & ~n5722;
  assign n5724 = n1248 & ~n5723;
  assign n5725 = n1252 & ~n5724;
  assign n5726 = n1256 & ~n5725;
  assign n5727 = n1260 & ~n5726;
  assign n5728 = n1264 & ~n5727;
  assign n5729 = n1268 & ~n5728;
  assign n5730 = n1272 & ~n5729;
  assign n5731 = n1276 & ~n5730;
  assign n5732 = n1280 & ~n5731;
  assign n5733 = n1284 & ~n5732;
  assign n5734 = n1288 & ~n5733;
  assign n5735 = n1292 & ~n5734;
  assign n5736 = n1296 & ~n5735;
  assign n5737 = n1300 & ~n5736;
  assign n5738 = n1304 & ~n5737;
  assign n5739 = n1308 & ~n5738;
  assign n5740 = n1312 & ~n5739;
  assign n5741 = n1316 & ~n5740;
  assign n5742 = n1320 & ~n5741;
  assign n5743 = n1324 & ~n5742;
  assign n5744 = n1328 & ~n5743;
  assign n5745 = n1332 & ~n5744;
  assign n5746 = n1336 & ~n5745;
  assign n5747 = n1340 & ~n5746;
  assign n5748 = n1344 & ~n5747;
  assign n5749 = n1348 & ~n5748;
  assign n5750 = n1352 & ~n5749;
  assign n5751 = n1356 & ~n5750;
  assign n5752 = n1360 & ~n5751;
  assign n5753 = n1364 & ~n5752;
  assign n5754 = n1368 & ~n5753;
  assign n5755 = n1372 & ~n5754;
  assign n5756 = n1376 & ~n5755;
  assign n5757 = n1380 & ~n5756;
  assign n5758 = n1384 & ~n5757;
  assign n5759 = n1388 & ~n5758;
  assign n5760 = n1392 & ~n5759;
  assign n5761 = n1396 & ~n5760;
  assign n5762 = n1663 & ~n5761;
  assign n5763 = n392 & ~n5762;
  assign n5764 = n396 & ~n5763;
  assign n5765 = n400 & ~n5764;
  assign n5766 = n404 & ~n5765;
  assign n5767 = n408 & ~n5766;
  assign n5768 = n412 & ~n5767;
  assign n5769 = n416 & ~n5768;
  assign n5770 = n420 & ~n5769;
  assign n5771 = n424 & ~n5770;
  assign n5772 = n428 & ~n5771;
  assign n5773 = n432 & ~n5772;
  assign n5774 = n436 & ~n5773;
  assign n5775 = n440 & ~n5774;
  assign n5776 = n444 & ~n5775;
  assign n5777 = n448 & ~n5776;
  assign n5778 = n452 & ~n5777;
  assign n5779 = n456 & ~n5778;
  assign n5780 = n460 & ~n5779;
  assign n5781 = n464 & ~n5780;
  assign n5782 = n468 & ~n5781;
  assign n5783 = n472 & ~n5782;
  assign n5784 = n476 & ~n5783;
  assign n5785 = n480 & ~n5784;
  assign n5786 = n484 & ~n5785;
  assign n5787 = n488 & ~n5786;
  assign n5788 = n492 & ~n5787;
  assign n5789 = n496 & ~n5788;
  assign n5790 = n500 & ~n5789;
  assign n5791 = n504 & ~n5790;
  assign n5792 = n508 & ~n5791;
  assign n5793 = n512 & ~n5792;
  assign n5794 = n516 & ~n5793;
  assign n5795 = n520 & ~n5794;
  assign n5796 = pi181  & ~n522;
  assign po53  = ~n5795 & n5796;
  assign n5798 = n531 & ~n866;
  assign n5799 = n536 & ~n5798;
  assign n5800 = n540 & ~n5799;
  assign n5801 = n544 & ~n5800;
  assign n5802 = n548 & ~n5801;
  assign n5803 = n552 & ~n5802;
  assign n5804 = n556 & ~n5803;
  assign n5805 = n560 & ~n5804;
  assign n5806 = n564 & ~n5805;
  assign n5807 = n568 & ~n5806;
  assign n5808 = n572 & ~n5807;
  assign n5809 = n576 & ~n5808;
  assign n5810 = n580 & ~n5809;
  assign n5811 = n584 & ~n5810;
  assign n5812 = n588 & ~n5811;
  assign n5813 = n592 & ~n5812;
  assign n5814 = n596 & ~n5813;
  assign n5815 = n600 & ~n5814;
  assign n5816 = n604 & ~n5815;
  assign n5817 = n608 & ~n5816;
  assign n5818 = n612 & ~n5817;
  assign n5819 = n616 & ~n5818;
  assign n5820 = n620 & ~n5819;
  assign n5821 = n624 & ~n5820;
  assign n5822 = n628 & ~n5821;
  assign n5823 = n632 & ~n5822;
  assign n5824 = n636 & ~n5823;
  assign n5825 = n640 & ~n5824;
  assign n5826 = n644 & ~n5825;
  assign n5827 = n648 & ~n5826;
  assign n5828 = n652 & ~n5827;
  assign n5829 = n656 & ~n5828;
  assign n5830 = n660 & ~n5829;
  assign n5831 = n664 & ~n5830;
  assign n5832 = n668 & ~n5831;
  assign n5833 = n672 & ~n5832;
  assign n5834 = n676 & ~n5833;
  assign n5835 = n680 & ~n5834;
  assign n5836 = n684 & ~n5835;
  assign n5837 = n688 & ~n5836;
  assign n5838 = n692 & ~n5837;
  assign n5839 = n696 & ~n5838;
  assign n5840 = n700 & ~n5839;
  assign n5841 = n704 & ~n5840;
  assign n5842 = n708 & ~n5841;
  assign n5843 = n712 & ~n5842;
  assign n5844 = n716 & ~n5843;
  assign n5845 = n720 & ~n5844;
  assign n5846 = n1484 & ~n5845;
  assign n5847 = n1486 & ~n5846;
  assign n5848 = n1750 & ~n5847;
  assign n5849 = n731 & ~n5848;
  assign n5850 = n735 & ~n5849;
  assign n5851 = n739 & ~n5850;
  assign n5852 = n743 & ~n5851;
  assign n5853 = n747 & ~n5852;
  assign n5854 = n751 & ~n5853;
  assign n5855 = n755 & ~n5854;
  assign n5856 = n759 & ~n5855;
  assign n5857 = n763 & ~n5856;
  assign n5858 = n767 & ~n5857;
  assign n5859 = n771 & ~n5858;
  assign n5860 = n775 & ~n5859;
  assign n5861 = n779 & ~n5860;
  assign n5862 = n783 & ~n5861;
  assign n5863 = n787 & ~n5862;
  assign n5864 = n791 & ~n5863;
  assign n5865 = n795 & ~n5864;
  assign n5866 = n799 & ~n5865;
  assign n5867 = n803 & ~n5866;
  assign n5868 = n807 & ~n5867;
  assign n5869 = n811 & ~n5868;
  assign n5870 = n815 & ~n5869;
  assign n5871 = n819 & ~n5870;
  assign n5872 = n823 & ~n5871;
  assign n5873 = n827 & ~n5872;
  assign n5874 = n831 & ~n5873;
  assign n5875 = n835 & ~n5874;
  assign n5876 = n839 & ~n5875;
  assign n5877 = n843 & ~n5876;
  assign n5878 = n847 & ~n5877;
  assign n5879 = n851 & ~n5878;
  assign n5880 = n855 & ~n5879;
  assign n5881 = n859 & ~n5880;
  assign n5882 = pi182  & ~n861;
  assign po54  = ~n5881 & n5882;
  assign n5884 = n870 & ~n1203;
  assign n5885 = n875 & ~n5884;
  assign n5886 = n879 & ~n5885;
  assign n5887 = n883 & ~n5886;
  assign n5888 = n887 & ~n5887;
  assign n5889 = n891 & ~n5888;
  assign n5890 = n895 & ~n5889;
  assign n5891 = n899 & ~n5890;
  assign n5892 = n903 & ~n5891;
  assign n5893 = n907 & ~n5892;
  assign n5894 = n911 & ~n5893;
  assign n5895 = n915 & ~n5894;
  assign n5896 = n919 & ~n5895;
  assign n5897 = n923 & ~n5896;
  assign n5898 = n927 & ~n5897;
  assign n5899 = n931 & ~n5898;
  assign n5900 = n935 & ~n5899;
  assign n5901 = n939 & ~n5900;
  assign n5902 = n943 & ~n5901;
  assign n5903 = n947 & ~n5902;
  assign n5904 = n951 & ~n5903;
  assign n5905 = n955 & ~n5904;
  assign n5906 = n959 & ~n5905;
  assign n5907 = n963 & ~n5906;
  assign n5908 = n967 & ~n5907;
  assign n5909 = n971 & ~n5908;
  assign n5910 = n975 & ~n5909;
  assign n5911 = n979 & ~n5910;
  assign n5912 = n983 & ~n5911;
  assign n5913 = n987 & ~n5912;
  assign n5914 = n991 & ~n5913;
  assign n5915 = n995 & ~n5914;
  assign n5916 = n999 & ~n5915;
  assign n5917 = n1003 & ~n5916;
  assign n5918 = n1007 & ~n5917;
  assign n5919 = n1011 & ~n5918;
  assign n5920 = n1015 & ~n5919;
  assign n5921 = n1019 & ~n5920;
  assign n5922 = n1023 & ~n5921;
  assign n5923 = n1027 & ~n5922;
  assign n5924 = n1031 & ~n5923;
  assign n5925 = n1035 & ~n5924;
  assign n5926 = n1039 & ~n5925;
  assign n5927 = n1043 & ~n5926;
  assign n5928 = n1047 & ~n5927;
  assign n5929 = n1051 & ~n5928;
  assign n5930 = n1055 & ~n5929;
  assign n5931 = n1059 & ~n5930;
  assign n5932 = n1574 & ~n5931;
  assign n5933 = n1576 & ~n5932;
  assign n5934 = n1837 & ~n5933;
  assign n5935 = n1068 & ~n5934;
  assign n5936 = n1072 & ~n5935;
  assign n5937 = n1076 & ~n5936;
  assign n5938 = n1080 & ~n5937;
  assign n5939 = n1084 & ~n5938;
  assign n5940 = n1088 & ~n5939;
  assign n5941 = n1092 & ~n5940;
  assign n5942 = n1096 & ~n5941;
  assign n5943 = n1100 & ~n5942;
  assign n5944 = n1104 & ~n5943;
  assign n5945 = n1108 & ~n5944;
  assign n5946 = n1112 & ~n5945;
  assign n5947 = n1116 & ~n5946;
  assign n5948 = n1120 & ~n5947;
  assign n5949 = n1124 & ~n5948;
  assign n5950 = n1128 & ~n5949;
  assign n5951 = n1132 & ~n5950;
  assign n5952 = n1136 & ~n5951;
  assign n5953 = n1140 & ~n5952;
  assign n5954 = n1144 & ~n5953;
  assign n5955 = n1148 & ~n5954;
  assign n5956 = n1152 & ~n5955;
  assign n5957 = n1156 & ~n5956;
  assign n5958 = n1160 & ~n5957;
  assign n5959 = n1164 & ~n5958;
  assign n5960 = n1168 & ~n5959;
  assign n5961 = n1172 & ~n5960;
  assign n5962 = n1176 & ~n5961;
  assign n5963 = n1180 & ~n5962;
  assign n5964 = n1184 & ~n5963;
  assign n5965 = n1188 & ~n5964;
  assign n5966 = n1192 & ~n5965;
  assign n5967 = n1196 & ~n5966;
  assign n5968 = pi183  & ~n1198;
  assign po55  = ~n5967 & n5968;
  assign n5970 = ~n535 & n1207;
  assign n5971 = n1212 & ~n5970;
  assign n5972 = n1216 & ~n5971;
  assign n5973 = n1220 & ~n5972;
  assign n5974 = n1224 & ~n5973;
  assign n5975 = n1228 & ~n5974;
  assign n5976 = n1232 & ~n5975;
  assign n5977 = n1236 & ~n5976;
  assign n5978 = n1240 & ~n5977;
  assign n5979 = n1244 & ~n5978;
  assign n5980 = n1248 & ~n5979;
  assign n5981 = n1252 & ~n5980;
  assign n5982 = n1256 & ~n5981;
  assign n5983 = n1260 & ~n5982;
  assign n5984 = n1264 & ~n5983;
  assign n5985 = n1268 & ~n5984;
  assign n5986 = n1272 & ~n5985;
  assign n5987 = n1276 & ~n5986;
  assign n5988 = n1280 & ~n5987;
  assign n5989 = n1284 & ~n5988;
  assign n5990 = n1288 & ~n5989;
  assign n5991 = n1292 & ~n5990;
  assign n5992 = n1296 & ~n5991;
  assign n5993 = n1300 & ~n5992;
  assign n5994 = n1304 & ~n5993;
  assign n5995 = n1308 & ~n5994;
  assign n5996 = n1312 & ~n5995;
  assign n5997 = n1316 & ~n5996;
  assign n5998 = n1320 & ~n5997;
  assign n5999 = n1324 & ~n5998;
  assign n6000 = n1328 & ~n5999;
  assign n6001 = n1332 & ~n6000;
  assign n6002 = n1336 & ~n6001;
  assign n6003 = n1340 & ~n6002;
  assign n6004 = n1344 & ~n6003;
  assign n6005 = n1348 & ~n6004;
  assign n6006 = n1352 & ~n6005;
  assign n6007 = n1356 & ~n6006;
  assign n6008 = n1360 & ~n6007;
  assign n6009 = n1364 & ~n6008;
  assign n6010 = n1368 & ~n6009;
  assign n6011 = n1372 & ~n6010;
  assign n6012 = n1376 & ~n6011;
  assign n6013 = n1380 & ~n6012;
  assign n6014 = n1384 & ~n6013;
  assign n6015 = n1388 & ~n6014;
  assign n6016 = n1392 & ~n6015;
  assign n6017 = n1396 & ~n6016;
  assign n6018 = n1663 & ~n6017;
  assign n6019 = n392 & ~n6018;
  assign n6020 = n396 & ~n6019;
  assign n6021 = n400 & ~n6020;
  assign n6022 = n404 & ~n6021;
  assign n6023 = n408 & ~n6022;
  assign n6024 = n412 & ~n6023;
  assign n6025 = n416 & ~n6024;
  assign n6026 = n420 & ~n6025;
  assign n6027 = n424 & ~n6026;
  assign n6028 = n428 & ~n6027;
  assign n6029 = n432 & ~n6028;
  assign n6030 = n436 & ~n6029;
  assign n6031 = n440 & ~n6030;
  assign n6032 = n444 & ~n6031;
  assign n6033 = n448 & ~n6032;
  assign n6034 = n452 & ~n6033;
  assign n6035 = n456 & ~n6034;
  assign n6036 = n460 & ~n6035;
  assign n6037 = n464 & ~n6036;
  assign n6038 = n468 & ~n6037;
  assign n6039 = n472 & ~n6038;
  assign n6040 = n476 & ~n6039;
  assign n6041 = n480 & ~n6040;
  assign n6042 = n484 & ~n6041;
  assign n6043 = n488 & ~n6042;
  assign n6044 = n492 & ~n6043;
  assign n6045 = n496 & ~n6044;
  assign n6046 = n500 & ~n6045;
  assign n6047 = n504 & ~n6046;
  assign n6048 = n508 & ~n6047;
  assign n6049 = n512 & ~n6048;
  assign n6050 = n516 & ~n6049;
  assign n6051 = n520 & ~n6050;
  assign n6052 = n524 & ~n6051;
  assign n6053 = n528 & ~n6052;
  assign n6054 = pi184  & ~n530;
  assign po56  = ~n6053 & n6054;
  assign n6056 = n539 & ~n874;
  assign n6057 = n544 & ~n6056;
  assign n6058 = n548 & ~n6057;
  assign n6059 = n552 & ~n6058;
  assign n6060 = n556 & ~n6059;
  assign n6061 = n560 & ~n6060;
  assign n6062 = n564 & ~n6061;
  assign n6063 = n568 & ~n6062;
  assign n6064 = n572 & ~n6063;
  assign n6065 = n576 & ~n6064;
  assign n6066 = n580 & ~n6065;
  assign n6067 = n584 & ~n6066;
  assign n6068 = n588 & ~n6067;
  assign n6069 = n592 & ~n6068;
  assign n6070 = n596 & ~n6069;
  assign n6071 = n600 & ~n6070;
  assign n6072 = n604 & ~n6071;
  assign n6073 = n608 & ~n6072;
  assign n6074 = n612 & ~n6073;
  assign n6075 = n616 & ~n6074;
  assign n6076 = n620 & ~n6075;
  assign n6077 = n624 & ~n6076;
  assign n6078 = n628 & ~n6077;
  assign n6079 = n632 & ~n6078;
  assign n6080 = n636 & ~n6079;
  assign n6081 = n640 & ~n6080;
  assign n6082 = n644 & ~n6081;
  assign n6083 = n648 & ~n6082;
  assign n6084 = n652 & ~n6083;
  assign n6085 = n656 & ~n6084;
  assign n6086 = n660 & ~n6085;
  assign n6087 = n664 & ~n6086;
  assign n6088 = n668 & ~n6087;
  assign n6089 = n672 & ~n6088;
  assign n6090 = n676 & ~n6089;
  assign n6091 = n680 & ~n6090;
  assign n6092 = n684 & ~n6091;
  assign n6093 = n688 & ~n6092;
  assign n6094 = n692 & ~n6093;
  assign n6095 = n696 & ~n6094;
  assign n6096 = n700 & ~n6095;
  assign n6097 = n704 & ~n6096;
  assign n6098 = n708 & ~n6097;
  assign n6099 = n712 & ~n6098;
  assign n6100 = n716 & ~n6099;
  assign n6101 = n720 & ~n6100;
  assign n6102 = n1484 & ~n6101;
  assign n6103 = n1486 & ~n6102;
  assign n6104 = n1750 & ~n6103;
  assign n6105 = n731 & ~n6104;
  assign n6106 = n735 & ~n6105;
  assign n6107 = n739 & ~n6106;
  assign n6108 = n743 & ~n6107;
  assign n6109 = n747 & ~n6108;
  assign n6110 = n751 & ~n6109;
  assign n6111 = n755 & ~n6110;
  assign n6112 = n759 & ~n6111;
  assign n6113 = n763 & ~n6112;
  assign n6114 = n767 & ~n6113;
  assign n6115 = n771 & ~n6114;
  assign n6116 = n775 & ~n6115;
  assign n6117 = n779 & ~n6116;
  assign n6118 = n783 & ~n6117;
  assign n6119 = n787 & ~n6118;
  assign n6120 = n791 & ~n6119;
  assign n6121 = n795 & ~n6120;
  assign n6122 = n799 & ~n6121;
  assign n6123 = n803 & ~n6122;
  assign n6124 = n807 & ~n6123;
  assign n6125 = n811 & ~n6124;
  assign n6126 = n815 & ~n6125;
  assign n6127 = n819 & ~n6126;
  assign n6128 = n823 & ~n6127;
  assign n6129 = n827 & ~n6128;
  assign n6130 = n831 & ~n6129;
  assign n6131 = n835 & ~n6130;
  assign n6132 = n839 & ~n6131;
  assign n6133 = n843 & ~n6132;
  assign n6134 = n847 & ~n6133;
  assign n6135 = n851 & ~n6134;
  assign n6136 = n855 & ~n6135;
  assign n6137 = n859 & ~n6136;
  assign n6138 = n863 & ~n6137;
  assign n6139 = n867 & ~n6138;
  assign n6140 = pi185  & ~n869;
  assign po57  = ~n6139 & n6140;
  assign n6142 = n878 & ~n1211;
  assign n6143 = n883 & ~n6142;
  assign n6144 = n887 & ~n6143;
  assign n6145 = n891 & ~n6144;
  assign n6146 = n895 & ~n6145;
  assign n6147 = n899 & ~n6146;
  assign n6148 = n903 & ~n6147;
  assign n6149 = n907 & ~n6148;
  assign n6150 = n911 & ~n6149;
  assign n6151 = n915 & ~n6150;
  assign n6152 = n919 & ~n6151;
  assign n6153 = n923 & ~n6152;
  assign n6154 = n927 & ~n6153;
  assign n6155 = n931 & ~n6154;
  assign n6156 = n935 & ~n6155;
  assign n6157 = n939 & ~n6156;
  assign n6158 = n943 & ~n6157;
  assign n6159 = n947 & ~n6158;
  assign n6160 = n951 & ~n6159;
  assign n6161 = n955 & ~n6160;
  assign n6162 = n959 & ~n6161;
  assign n6163 = n963 & ~n6162;
  assign n6164 = n967 & ~n6163;
  assign n6165 = n971 & ~n6164;
  assign n6166 = n975 & ~n6165;
  assign n6167 = n979 & ~n6166;
  assign n6168 = n983 & ~n6167;
  assign n6169 = n987 & ~n6168;
  assign n6170 = n991 & ~n6169;
  assign n6171 = n995 & ~n6170;
  assign n6172 = n999 & ~n6171;
  assign n6173 = n1003 & ~n6172;
  assign n6174 = n1007 & ~n6173;
  assign n6175 = n1011 & ~n6174;
  assign n6176 = n1015 & ~n6175;
  assign n6177 = n1019 & ~n6176;
  assign n6178 = n1023 & ~n6177;
  assign n6179 = n1027 & ~n6178;
  assign n6180 = n1031 & ~n6179;
  assign n6181 = n1035 & ~n6180;
  assign n6182 = n1039 & ~n6181;
  assign n6183 = n1043 & ~n6182;
  assign n6184 = n1047 & ~n6183;
  assign n6185 = n1051 & ~n6184;
  assign n6186 = n1055 & ~n6185;
  assign n6187 = n1059 & ~n6186;
  assign n6188 = n1574 & ~n6187;
  assign n6189 = n1576 & ~n6188;
  assign n6190 = n1837 & ~n6189;
  assign n6191 = n1068 & ~n6190;
  assign n6192 = n1072 & ~n6191;
  assign n6193 = n1076 & ~n6192;
  assign n6194 = n1080 & ~n6193;
  assign n6195 = n1084 & ~n6194;
  assign n6196 = n1088 & ~n6195;
  assign n6197 = n1092 & ~n6196;
  assign n6198 = n1096 & ~n6197;
  assign n6199 = n1100 & ~n6198;
  assign n6200 = n1104 & ~n6199;
  assign n6201 = n1108 & ~n6200;
  assign n6202 = n1112 & ~n6201;
  assign n6203 = n1116 & ~n6202;
  assign n6204 = n1120 & ~n6203;
  assign n6205 = n1124 & ~n6204;
  assign n6206 = n1128 & ~n6205;
  assign n6207 = n1132 & ~n6206;
  assign n6208 = n1136 & ~n6207;
  assign n6209 = n1140 & ~n6208;
  assign n6210 = n1144 & ~n6209;
  assign n6211 = n1148 & ~n6210;
  assign n6212 = n1152 & ~n6211;
  assign n6213 = n1156 & ~n6212;
  assign n6214 = n1160 & ~n6213;
  assign n6215 = n1164 & ~n6214;
  assign n6216 = n1168 & ~n6215;
  assign n6217 = n1172 & ~n6216;
  assign n6218 = n1176 & ~n6217;
  assign n6219 = n1180 & ~n6218;
  assign n6220 = n1184 & ~n6219;
  assign n6221 = n1188 & ~n6220;
  assign n6222 = n1192 & ~n6221;
  assign n6223 = n1196 & ~n6222;
  assign n6224 = n1200 & ~n6223;
  assign n6225 = n1204 & ~n6224;
  assign n6226 = pi186  & ~n1206;
  assign po58  = ~n6225 & n6226;
  assign n6228 = ~n543 & n1215;
  assign n6229 = n1220 & ~n6228;
  assign n6230 = n1224 & ~n6229;
  assign n6231 = n1228 & ~n6230;
  assign n6232 = n1232 & ~n6231;
  assign n6233 = n1236 & ~n6232;
  assign n6234 = n1240 & ~n6233;
  assign n6235 = n1244 & ~n6234;
  assign n6236 = n1248 & ~n6235;
  assign n6237 = n1252 & ~n6236;
  assign n6238 = n1256 & ~n6237;
  assign n6239 = n1260 & ~n6238;
  assign n6240 = n1264 & ~n6239;
  assign n6241 = n1268 & ~n6240;
  assign n6242 = n1272 & ~n6241;
  assign n6243 = n1276 & ~n6242;
  assign n6244 = n1280 & ~n6243;
  assign n6245 = n1284 & ~n6244;
  assign n6246 = n1288 & ~n6245;
  assign n6247 = n1292 & ~n6246;
  assign n6248 = n1296 & ~n6247;
  assign n6249 = n1300 & ~n6248;
  assign n6250 = n1304 & ~n6249;
  assign n6251 = n1308 & ~n6250;
  assign n6252 = n1312 & ~n6251;
  assign n6253 = n1316 & ~n6252;
  assign n6254 = n1320 & ~n6253;
  assign n6255 = n1324 & ~n6254;
  assign n6256 = n1328 & ~n6255;
  assign n6257 = n1332 & ~n6256;
  assign n6258 = n1336 & ~n6257;
  assign n6259 = n1340 & ~n6258;
  assign n6260 = n1344 & ~n6259;
  assign n6261 = n1348 & ~n6260;
  assign n6262 = n1352 & ~n6261;
  assign n6263 = n1356 & ~n6262;
  assign n6264 = n1360 & ~n6263;
  assign n6265 = n1364 & ~n6264;
  assign n6266 = n1368 & ~n6265;
  assign n6267 = n1372 & ~n6266;
  assign n6268 = n1376 & ~n6267;
  assign n6269 = n1380 & ~n6268;
  assign n6270 = n1384 & ~n6269;
  assign n6271 = n1388 & ~n6270;
  assign n6272 = n1392 & ~n6271;
  assign n6273 = n1396 & ~n6272;
  assign n6274 = n1663 & ~n6273;
  assign n6275 = n392 & ~n6274;
  assign n6276 = n396 & ~n6275;
  assign n6277 = n400 & ~n6276;
  assign n6278 = n404 & ~n6277;
  assign n6279 = n408 & ~n6278;
  assign n6280 = n412 & ~n6279;
  assign n6281 = n416 & ~n6280;
  assign n6282 = n420 & ~n6281;
  assign n6283 = n424 & ~n6282;
  assign n6284 = n428 & ~n6283;
  assign n6285 = n432 & ~n6284;
  assign n6286 = n436 & ~n6285;
  assign n6287 = n440 & ~n6286;
  assign n6288 = n444 & ~n6287;
  assign n6289 = n448 & ~n6288;
  assign n6290 = n452 & ~n6289;
  assign n6291 = n456 & ~n6290;
  assign n6292 = n460 & ~n6291;
  assign n6293 = n464 & ~n6292;
  assign n6294 = n468 & ~n6293;
  assign n6295 = n472 & ~n6294;
  assign n6296 = n476 & ~n6295;
  assign n6297 = n480 & ~n6296;
  assign n6298 = n484 & ~n6297;
  assign n6299 = n488 & ~n6298;
  assign n6300 = n492 & ~n6299;
  assign n6301 = n496 & ~n6300;
  assign n6302 = n500 & ~n6301;
  assign n6303 = n504 & ~n6302;
  assign n6304 = n508 & ~n6303;
  assign n6305 = n512 & ~n6304;
  assign n6306 = n516 & ~n6305;
  assign n6307 = n520 & ~n6306;
  assign n6308 = n524 & ~n6307;
  assign n6309 = n528 & ~n6308;
  assign n6310 = n532 & ~n6309;
  assign n6311 = n536 & ~n6310;
  assign n6312 = pi187  & ~n538;
  assign po59  = ~n6311 & n6312;
  assign n6314 = n547 & ~n882;
  assign n6315 = n552 & ~n6314;
  assign n6316 = n556 & ~n6315;
  assign n6317 = n560 & ~n6316;
  assign n6318 = n564 & ~n6317;
  assign n6319 = n568 & ~n6318;
  assign n6320 = n572 & ~n6319;
  assign n6321 = n576 & ~n6320;
  assign n6322 = n580 & ~n6321;
  assign n6323 = n584 & ~n6322;
  assign n6324 = n588 & ~n6323;
  assign n6325 = n592 & ~n6324;
  assign n6326 = n596 & ~n6325;
  assign n6327 = n600 & ~n6326;
  assign n6328 = n604 & ~n6327;
  assign n6329 = n608 & ~n6328;
  assign n6330 = n612 & ~n6329;
  assign n6331 = n616 & ~n6330;
  assign n6332 = n620 & ~n6331;
  assign n6333 = n624 & ~n6332;
  assign n6334 = n628 & ~n6333;
  assign n6335 = n632 & ~n6334;
  assign n6336 = n636 & ~n6335;
  assign n6337 = n640 & ~n6336;
  assign n6338 = n644 & ~n6337;
  assign n6339 = n648 & ~n6338;
  assign n6340 = n652 & ~n6339;
  assign n6341 = n656 & ~n6340;
  assign n6342 = n660 & ~n6341;
  assign n6343 = n664 & ~n6342;
  assign n6344 = n668 & ~n6343;
  assign n6345 = n672 & ~n6344;
  assign n6346 = n676 & ~n6345;
  assign n6347 = n680 & ~n6346;
  assign n6348 = n684 & ~n6347;
  assign n6349 = n688 & ~n6348;
  assign n6350 = n692 & ~n6349;
  assign n6351 = n696 & ~n6350;
  assign n6352 = n700 & ~n6351;
  assign n6353 = n704 & ~n6352;
  assign n6354 = n708 & ~n6353;
  assign n6355 = n712 & ~n6354;
  assign n6356 = n716 & ~n6355;
  assign n6357 = n720 & ~n6356;
  assign n6358 = n1484 & ~n6357;
  assign n6359 = n1486 & ~n6358;
  assign n6360 = n1750 & ~n6359;
  assign n6361 = n731 & ~n6360;
  assign n6362 = n735 & ~n6361;
  assign n6363 = n739 & ~n6362;
  assign n6364 = n743 & ~n6363;
  assign n6365 = n747 & ~n6364;
  assign n6366 = n751 & ~n6365;
  assign n6367 = n755 & ~n6366;
  assign n6368 = n759 & ~n6367;
  assign n6369 = n763 & ~n6368;
  assign n6370 = n767 & ~n6369;
  assign n6371 = n771 & ~n6370;
  assign n6372 = n775 & ~n6371;
  assign n6373 = n779 & ~n6372;
  assign n6374 = n783 & ~n6373;
  assign n6375 = n787 & ~n6374;
  assign n6376 = n791 & ~n6375;
  assign n6377 = n795 & ~n6376;
  assign n6378 = n799 & ~n6377;
  assign n6379 = n803 & ~n6378;
  assign n6380 = n807 & ~n6379;
  assign n6381 = n811 & ~n6380;
  assign n6382 = n815 & ~n6381;
  assign n6383 = n819 & ~n6382;
  assign n6384 = n823 & ~n6383;
  assign n6385 = n827 & ~n6384;
  assign n6386 = n831 & ~n6385;
  assign n6387 = n835 & ~n6386;
  assign n6388 = n839 & ~n6387;
  assign n6389 = n843 & ~n6388;
  assign n6390 = n847 & ~n6389;
  assign n6391 = n851 & ~n6390;
  assign n6392 = n855 & ~n6391;
  assign n6393 = n859 & ~n6392;
  assign n6394 = n863 & ~n6393;
  assign n6395 = n867 & ~n6394;
  assign n6396 = n871 & ~n6395;
  assign n6397 = n875 & ~n6396;
  assign n6398 = pi188  & ~n877;
  assign po60  = ~n6397 & n6398;
  assign n6400 = n886 & ~n1219;
  assign n6401 = n891 & ~n6400;
  assign n6402 = n895 & ~n6401;
  assign n6403 = n899 & ~n6402;
  assign n6404 = n903 & ~n6403;
  assign n6405 = n907 & ~n6404;
  assign n6406 = n911 & ~n6405;
  assign n6407 = n915 & ~n6406;
  assign n6408 = n919 & ~n6407;
  assign n6409 = n923 & ~n6408;
  assign n6410 = n927 & ~n6409;
  assign n6411 = n931 & ~n6410;
  assign n6412 = n935 & ~n6411;
  assign n6413 = n939 & ~n6412;
  assign n6414 = n943 & ~n6413;
  assign n6415 = n947 & ~n6414;
  assign n6416 = n951 & ~n6415;
  assign n6417 = n955 & ~n6416;
  assign n6418 = n959 & ~n6417;
  assign n6419 = n963 & ~n6418;
  assign n6420 = n967 & ~n6419;
  assign n6421 = n971 & ~n6420;
  assign n6422 = n975 & ~n6421;
  assign n6423 = n979 & ~n6422;
  assign n6424 = n983 & ~n6423;
  assign n6425 = n987 & ~n6424;
  assign n6426 = n991 & ~n6425;
  assign n6427 = n995 & ~n6426;
  assign n6428 = n999 & ~n6427;
  assign n6429 = n1003 & ~n6428;
  assign n6430 = n1007 & ~n6429;
  assign n6431 = n1011 & ~n6430;
  assign n6432 = n1015 & ~n6431;
  assign n6433 = n1019 & ~n6432;
  assign n6434 = n1023 & ~n6433;
  assign n6435 = n1027 & ~n6434;
  assign n6436 = n1031 & ~n6435;
  assign n6437 = n1035 & ~n6436;
  assign n6438 = n1039 & ~n6437;
  assign n6439 = n1043 & ~n6438;
  assign n6440 = n1047 & ~n6439;
  assign n6441 = n1051 & ~n6440;
  assign n6442 = n1055 & ~n6441;
  assign n6443 = n1059 & ~n6442;
  assign n6444 = n1574 & ~n6443;
  assign n6445 = n1576 & ~n6444;
  assign n6446 = n1837 & ~n6445;
  assign n6447 = n1068 & ~n6446;
  assign n6448 = n1072 & ~n6447;
  assign n6449 = n1076 & ~n6448;
  assign n6450 = n1080 & ~n6449;
  assign n6451 = n1084 & ~n6450;
  assign n6452 = n1088 & ~n6451;
  assign n6453 = n1092 & ~n6452;
  assign n6454 = n1096 & ~n6453;
  assign n6455 = n1100 & ~n6454;
  assign n6456 = n1104 & ~n6455;
  assign n6457 = n1108 & ~n6456;
  assign n6458 = n1112 & ~n6457;
  assign n6459 = n1116 & ~n6458;
  assign n6460 = n1120 & ~n6459;
  assign n6461 = n1124 & ~n6460;
  assign n6462 = n1128 & ~n6461;
  assign n6463 = n1132 & ~n6462;
  assign n6464 = n1136 & ~n6463;
  assign n6465 = n1140 & ~n6464;
  assign n6466 = n1144 & ~n6465;
  assign n6467 = n1148 & ~n6466;
  assign n6468 = n1152 & ~n6467;
  assign n6469 = n1156 & ~n6468;
  assign n6470 = n1160 & ~n6469;
  assign n6471 = n1164 & ~n6470;
  assign n6472 = n1168 & ~n6471;
  assign n6473 = n1172 & ~n6472;
  assign n6474 = n1176 & ~n6473;
  assign n6475 = n1180 & ~n6474;
  assign n6476 = n1184 & ~n6475;
  assign n6477 = n1188 & ~n6476;
  assign n6478 = n1192 & ~n6477;
  assign n6479 = n1196 & ~n6478;
  assign n6480 = n1200 & ~n6479;
  assign n6481 = n1204 & ~n6480;
  assign n6482 = n1208 & ~n6481;
  assign n6483 = n1212 & ~n6482;
  assign n6484 = pi189  & ~n1214;
  assign po61  = ~n6483 & n6484;
  assign n6486 = ~n551 & n1223;
  assign n6487 = n1228 & ~n6486;
  assign n6488 = n1232 & ~n6487;
  assign n6489 = n1236 & ~n6488;
  assign n6490 = n1240 & ~n6489;
  assign n6491 = n1244 & ~n6490;
  assign n6492 = n1248 & ~n6491;
  assign n6493 = n1252 & ~n6492;
  assign n6494 = n1256 & ~n6493;
  assign n6495 = n1260 & ~n6494;
  assign n6496 = n1264 & ~n6495;
  assign n6497 = n1268 & ~n6496;
  assign n6498 = n1272 & ~n6497;
  assign n6499 = n1276 & ~n6498;
  assign n6500 = n1280 & ~n6499;
  assign n6501 = n1284 & ~n6500;
  assign n6502 = n1288 & ~n6501;
  assign n6503 = n1292 & ~n6502;
  assign n6504 = n1296 & ~n6503;
  assign n6505 = n1300 & ~n6504;
  assign n6506 = n1304 & ~n6505;
  assign n6507 = n1308 & ~n6506;
  assign n6508 = n1312 & ~n6507;
  assign n6509 = n1316 & ~n6508;
  assign n6510 = n1320 & ~n6509;
  assign n6511 = n1324 & ~n6510;
  assign n6512 = n1328 & ~n6511;
  assign n6513 = n1332 & ~n6512;
  assign n6514 = n1336 & ~n6513;
  assign n6515 = n1340 & ~n6514;
  assign n6516 = n1344 & ~n6515;
  assign n6517 = n1348 & ~n6516;
  assign n6518 = n1352 & ~n6517;
  assign n6519 = n1356 & ~n6518;
  assign n6520 = n1360 & ~n6519;
  assign n6521 = n1364 & ~n6520;
  assign n6522 = n1368 & ~n6521;
  assign n6523 = n1372 & ~n6522;
  assign n6524 = n1376 & ~n6523;
  assign n6525 = n1380 & ~n6524;
  assign n6526 = n1384 & ~n6525;
  assign n6527 = n1388 & ~n6526;
  assign n6528 = n1392 & ~n6527;
  assign n6529 = n1396 & ~n6528;
  assign n6530 = n1663 & ~n6529;
  assign n6531 = n392 & ~n6530;
  assign n6532 = n396 & ~n6531;
  assign n6533 = n400 & ~n6532;
  assign n6534 = n404 & ~n6533;
  assign n6535 = n408 & ~n6534;
  assign n6536 = n412 & ~n6535;
  assign n6537 = n416 & ~n6536;
  assign n6538 = n420 & ~n6537;
  assign n6539 = n424 & ~n6538;
  assign n6540 = n428 & ~n6539;
  assign n6541 = n432 & ~n6540;
  assign n6542 = n436 & ~n6541;
  assign n6543 = n440 & ~n6542;
  assign n6544 = n444 & ~n6543;
  assign n6545 = n448 & ~n6544;
  assign n6546 = n452 & ~n6545;
  assign n6547 = n456 & ~n6546;
  assign n6548 = n460 & ~n6547;
  assign n6549 = n464 & ~n6548;
  assign n6550 = n468 & ~n6549;
  assign n6551 = n472 & ~n6550;
  assign n6552 = n476 & ~n6551;
  assign n6553 = n480 & ~n6552;
  assign n6554 = n484 & ~n6553;
  assign n6555 = n488 & ~n6554;
  assign n6556 = n492 & ~n6555;
  assign n6557 = n496 & ~n6556;
  assign n6558 = n500 & ~n6557;
  assign n6559 = n504 & ~n6558;
  assign n6560 = n508 & ~n6559;
  assign n6561 = n512 & ~n6560;
  assign n6562 = n516 & ~n6561;
  assign n6563 = n520 & ~n6562;
  assign n6564 = n524 & ~n6563;
  assign n6565 = n528 & ~n6564;
  assign n6566 = n532 & ~n6565;
  assign n6567 = n536 & ~n6566;
  assign n6568 = n540 & ~n6567;
  assign n6569 = n544 & ~n6568;
  assign n6570 = pi190  & ~n546;
  assign po62  = ~n6569 & n6570;
  assign n6572 = n555 & ~n890;
  assign n6573 = n560 & ~n6572;
  assign n6574 = n564 & ~n6573;
  assign n6575 = n568 & ~n6574;
  assign n6576 = n572 & ~n6575;
  assign n6577 = n576 & ~n6576;
  assign n6578 = n580 & ~n6577;
  assign n6579 = n584 & ~n6578;
  assign n6580 = n588 & ~n6579;
  assign n6581 = n592 & ~n6580;
  assign n6582 = n596 & ~n6581;
  assign n6583 = n600 & ~n6582;
  assign n6584 = n604 & ~n6583;
  assign n6585 = n608 & ~n6584;
  assign n6586 = n612 & ~n6585;
  assign n6587 = n616 & ~n6586;
  assign n6588 = n620 & ~n6587;
  assign n6589 = n624 & ~n6588;
  assign n6590 = n628 & ~n6589;
  assign n6591 = n632 & ~n6590;
  assign n6592 = n636 & ~n6591;
  assign n6593 = n640 & ~n6592;
  assign n6594 = n644 & ~n6593;
  assign n6595 = n648 & ~n6594;
  assign n6596 = n652 & ~n6595;
  assign n6597 = n656 & ~n6596;
  assign n6598 = n660 & ~n6597;
  assign n6599 = n664 & ~n6598;
  assign n6600 = n668 & ~n6599;
  assign n6601 = n672 & ~n6600;
  assign n6602 = n676 & ~n6601;
  assign n6603 = n680 & ~n6602;
  assign n6604 = n684 & ~n6603;
  assign n6605 = n688 & ~n6604;
  assign n6606 = n692 & ~n6605;
  assign n6607 = n696 & ~n6606;
  assign n6608 = n700 & ~n6607;
  assign n6609 = n704 & ~n6608;
  assign n6610 = n708 & ~n6609;
  assign n6611 = n712 & ~n6610;
  assign n6612 = n716 & ~n6611;
  assign n6613 = n720 & ~n6612;
  assign n6614 = n1484 & ~n6613;
  assign n6615 = n1486 & ~n6614;
  assign n6616 = n1750 & ~n6615;
  assign n6617 = n731 & ~n6616;
  assign n6618 = n735 & ~n6617;
  assign n6619 = n739 & ~n6618;
  assign n6620 = n743 & ~n6619;
  assign n6621 = n747 & ~n6620;
  assign n6622 = n751 & ~n6621;
  assign n6623 = n755 & ~n6622;
  assign n6624 = n759 & ~n6623;
  assign n6625 = n763 & ~n6624;
  assign n6626 = n767 & ~n6625;
  assign n6627 = n771 & ~n6626;
  assign n6628 = n775 & ~n6627;
  assign n6629 = n779 & ~n6628;
  assign n6630 = n783 & ~n6629;
  assign n6631 = n787 & ~n6630;
  assign n6632 = n791 & ~n6631;
  assign n6633 = n795 & ~n6632;
  assign n6634 = n799 & ~n6633;
  assign n6635 = n803 & ~n6634;
  assign n6636 = n807 & ~n6635;
  assign n6637 = n811 & ~n6636;
  assign n6638 = n815 & ~n6637;
  assign n6639 = n819 & ~n6638;
  assign n6640 = n823 & ~n6639;
  assign n6641 = n827 & ~n6640;
  assign n6642 = n831 & ~n6641;
  assign n6643 = n835 & ~n6642;
  assign n6644 = n839 & ~n6643;
  assign n6645 = n843 & ~n6644;
  assign n6646 = n847 & ~n6645;
  assign n6647 = n851 & ~n6646;
  assign n6648 = n855 & ~n6647;
  assign n6649 = n859 & ~n6648;
  assign n6650 = n863 & ~n6649;
  assign n6651 = n867 & ~n6650;
  assign n6652 = n871 & ~n6651;
  assign n6653 = n875 & ~n6652;
  assign n6654 = n879 & ~n6653;
  assign n6655 = n883 & ~n6654;
  assign n6656 = pi191  & ~n885;
  assign po63  = ~n6655 & n6656;
  assign n6658 = n894 & ~n1227;
  assign n6659 = n899 & ~n6658;
  assign n6660 = n903 & ~n6659;
  assign n6661 = n907 & ~n6660;
  assign n6662 = n911 & ~n6661;
  assign n6663 = n915 & ~n6662;
  assign n6664 = n919 & ~n6663;
  assign n6665 = n923 & ~n6664;
  assign n6666 = n927 & ~n6665;
  assign n6667 = n931 & ~n6666;
  assign n6668 = n935 & ~n6667;
  assign n6669 = n939 & ~n6668;
  assign n6670 = n943 & ~n6669;
  assign n6671 = n947 & ~n6670;
  assign n6672 = n951 & ~n6671;
  assign n6673 = n955 & ~n6672;
  assign n6674 = n959 & ~n6673;
  assign n6675 = n963 & ~n6674;
  assign n6676 = n967 & ~n6675;
  assign n6677 = n971 & ~n6676;
  assign n6678 = n975 & ~n6677;
  assign n6679 = n979 & ~n6678;
  assign n6680 = n983 & ~n6679;
  assign n6681 = n987 & ~n6680;
  assign n6682 = n991 & ~n6681;
  assign n6683 = n995 & ~n6682;
  assign n6684 = n999 & ~n6683;
  assign n6685 = n1003 & ~n6684;
  assign n6686 = n1007 & ~n6685;
  assign n6687 = n1011 & ~n6686;
  assign n6688 = n1015 & ~n6687;
  assign n6689 = n1019 & ~n6688;
  assign n6690 = n1023 & ~n6689;
  assign n6691 = n1027 & ~n6690;
  assign n6692 = n1031 & ~n6691;
  assign n6693 = n1035 & ~n6692;
  assign n6694 = n1039 & ~n6693;
  assign n6695 = n1043 & ~n6694;
  assign n6696 = n1047 & ~n6695;
  assign n6697 = n1051 & ~n6696;
  assign n6698 = n1055 & ~n6697;
  assign n6699 = n1059 & ~n6698;
  assign n6700 = n1574 & ~n6699;
  assign n6701 = n1576 & ~n6700;
  assign n6702 = n1837 & ~n6701;
  assign n6703 = n1068 & ~n6702;
  assign n6704 = n1072 & ~n6703;
  assign n6705 = n1076 & ~n6704;
  assign n6706 = n1080 & ~n6705;
  assign n6707 = n1084 & ~n6706;
  assign n6708 = n1088 & ~n6707;
  assign n6709 = n1092 & ~n6708;
  assign n6710 = n1096 & ~n6709;
  assign n6711 = n1100 & ~n6710;
  assign n6712 = n1104 & ~n6711;
  assign n6713 = n1108 & ~n6712;
  assign n6714 = n1112 & ~n6713;
  assign n6715 = n1116 & ~n6714;
  assign n6716 = n1120 & ~n6715;
  assign n6717 = n1124 & ~n6716;
  assign n6718 = n1128 & ~n6717;
  assign n6719 = n1132 & ~n6718;
  assign n6720 = n1136 & ~n6719;
  assign n6721 = n1140 & ~n6720;
  assign n6722 = n1144 & ~n6721;
  assign n6723 = n1148 & ~n6722;
  assign n6724 = n1152 & ~n6723;
  assign n6725 = n1156 & ~n6724;
  assign n6726 = n1160 & ~n6725;
  assign n6727 = n1164 & ~n6726;
  assign n6728 = n1168 & ~n6727;
  assign n6729 = n1172 & ~n6728;
  assign n6730 = n1176 & ~n6729;
  assign n6731 = n1180 & ~n6730;
  assign n6732 = n1184 & ~n6731;
  assign n6733 = n1188 & ~n6732;
  assign n6734 = n1192 & ~n6733;
  assign n6735 = n1196 & ~n6734;
  assign n6736 = n1200 & ~n6735;
  assign n6737 = n1204 & ~n6736;
  assign n6738 = n1208 & ~n6737;
  assign n6739 = n1212 & ~n6738;
  assign n6740 = n1216 & ~n6739;
  assign n6741 = n1220 & ~n6740;
  assign n6742 = pi192  & ~n1222;
  assign po64  = ~n6741 & n6742;
  assign n6744 = ~n559 & n1231;
  assign n6745 = n1236 & ~n6744;
  assign n6746 = n1240 & ~n6745;
  assign n6747 = n1244 & ~n6746;
  assign n6748 = n1248 & ~n6747;
  assign n6749 = n1252 & ~n6748;
  assign n6750 = n1256 & ~n6749;
  assign n6751 = n1260 & ~n6750;
  assign n6752 = n1264 & ~n6751;
  assign n6753 = n1268 & ~n6752;
  assign n6754 = n1272 & ~n6753;
  assign n6755 = n1276 & ~n6754;
  assign n6756 = n1280 & ~n6755;
  assign n6757 = n1284 & ~n6756;
  assign n6758 = n1288 & ~n6757;
  assign n6759 = n1292 & ~n6758;
  assign n6760 = n1296 & ~n6759;
  assign n6761 = n1300 & ~n6760;
  assign n6762 = n1304 & ~n6761;
  assign n6763 = n1308 & ~n6762;
  assign n6764 = n1312 & ~n6763;
  assign n6765 = n1316 & ~n6764;
  assign n6766 = n1320 & ~n6765;
  assign n6767 = n1324 & ~n6766;
  assign n6768 = n1328 & ~n6767;
  assign n6769 = n1332 & ~n6768;
  assign n6770 = n1336 & ~n6769;
  assign n6771 = n1340 & ~n6770;
  assign n6772 = n1344 & ~n6771;
  assign n6773 = n1348 & ~n6772;
  assign n6774 = n1352 & ~n6773;
  assign n6775 = n1356 & ~n6774;
  assign n6776 = n1360 & ~n6775;
  assign n6777 = n1364 & ~n6776;
  assign n6778 = n1368 & ~n6777;
  assign n6779 = n1372 & ~n6778;
  assign n6780 = n1376 & ~n6779;
  assign n6781 = n1380 & ~n6780;
  assign n6782 = n1384 & ~n6781;
  assign n6783 = n1388 & ~n6782;
  assign n6784 = n1392 & ~n6783;
  assign n6785 = n1396 & ~n6784;
  assign n6786 = n1663 & ~n6785;
  assign n6787 = n392 & ~n6786;
  assign n6788 = n396 & ~n6787;
  assign n6789 = n400 & ~n6788;
  assign n6790 = n404 & ~n6789;
  assign n6791 = n408 & ~n6790;
  assign n6792 = n412 & ~n6791;
  assign n6793 = n416 & ~n6792;
  assign n6794 = n420 & ~n6793;
  assign n6795 = n424 & ~n6794;
  assign n6796 = n428 & ~n6795;
  assign n6797 = n432 & ~n6796;
  assign n6798 = n436 & ~n6797;
  assign n6799 = n440 & ~n6798;
  assign n6800 = n444 & ~n6799;
  assign n6801 = n448 & ~n6800;
  assign n6802 = n452 & ~n6801;
  assign n6803 = n456 & ~n6802;
  assign n6804 = n460 & ~n6803;
  assign n6805 = n464 & ~n6804;
  assign n6806 = n468 & ~n6805;
  assign n6807 = n472 & ~n6806;
  assign n6808 = n476 & ~n6807;
  assign n6809 = n480 & ~n6808;
  assign n6810 = n484 & ~n6809;
  assign n6811 = n488 & ~n6810;
  assign n6812 = n492 & ~n6811;
  assign n6813 = n496 & ~n6812;
  assign n6814 = n500 & ~n6813;
  assign n6815 = n504 & ~n6814;
  assign n6816 = n508 & ~n6815;
  assign n6817 = n512 & ~n6816;
  assign n6818 = n516 & ~n6817;
  assign n6819 = n520 & ~n6818;
  assign n6820 = n524 & ~n6819;
  assign n6821 = n528 & ~n6820;
  assign n6822 = n532 & ~n6821;
  assign n6823 = n536 & ~n6822;
  assign n6824 = n540 & ~n6823;
  assign n6825 = n544 & ~n6824;
  assign n6826 = n548 & ~n6825;
  assign n6827 = n552 & ~n6826;
  assign n6828 = pi193  & ~n554;
  assign po65  = ~n6827 & n6828;
  assign n6830 = n563 & ~n898;
  assign n6831 = n568 & ~n6830;
  assign n6832 = n572 & ~n6831;
  assign n6833 = n576 & ~n6832;
  assign n6834 = n580 & ~n6833;
  assign n6835 = n584 & ~n6834;
  assign n6836 = n588 & ~n6835;
  assign n6837 = n592 & ~n6836;
  assign n6838 = n596 & ~n6837;
  assign n6839 = n600 & ~n6838;
  assign n6840 = n604 & ~n6839;
  assign n6841 = n608 & ~n6840;
  assign n6842 = n612 & ~n6841;
  assign n6843 = n616 & ~n6842;
  assign n6844 = n620 & ~n6843;
  assign n6845 = n624 & ~n6844;
  assign n6846 = n628 & ~n6845;
  assign n6847 = n632 & ~n6846;
  assign n6848 = n636 & ~n6847;
  assign n6849 = n640 & ~n6848;
  assign n6850 = n644 & ~n6849;
  assign n6851 = n648 & ~n6850;
  assign n6852 = n652 & ~n6851;
  assign n6853 = n656 & ~n6852;
  assign n6854 = n660 & ~n6853;
  assign n6855 = n664 & ~n6854;
  assign n6856 = n668 & ~n6855;
  assign n6857 = n672 & ~n6856;
  assign n6858 = n676 & ~n6857;
  assign n6859 = n680 & ~n6858;
  assign n6860 = n684 & ~n6859;
  assign n6861 = n688 & ~n6860;
  assign n6862 = n692 & ~n6861;
  assign n6863 = n696 & ~n6862;
  assign n6864 = n700 & ~n6863;
  assign n6865 = n704 & ~n6864;
  assign n6866 = n708 & ~n6865;
  assign n6867 = n712 & ~n6866;
  assign n6868 = n716 & ~n6867;
  assign n6869 = n720 & ~n6868;
  assign n6870 = n1484 & ~n6869;
  assign n6871 = n1486 & ~n6870;
  assign n6872 = n1750 & ~n6871;
  assign n6873 = n731 & ~n6872;
  assign n6874 = n735 & ~n6873;
  assign n6875 = n739 & ~n6874;
  assign n6876 = n743 & ~n6875;
  assign n6877 = n747 & ~n6876;
  assign n6878 = n751 & ~n6877;
  assign n6879 = n755 & ~n6878;
  assign n6880 = n759 & ~n6879;
  assign n6881 = n763 & ~n6880;
  assign n6882 = n767 & ~n6881;
  assign n6883 = n771 & ~n6882;
  assign n6884 = n775 & ~n6883;
  assign n6885 = n779 & ~n6884;
  assign n6886 = n783 & ~n6885;
  assign n6887 = n787 & ~n6886;
  assign n6888 = n791 & ~n6887;
  assign n6889 = n795 & ~n6888;
  assign n6890 = n799 & ~n6889;
  assign n6891 = n803 & ~n6890;
  assign n6892 = n807 & ~n6891;
  assign n6893 = n811 & ~n6892;
  assign n6894 = n815 & ~n6893;
  assign n6895 = n819 & ~n6894;
  assign n6896 = n823 & ~n6895;
  assign n6897 = n827 & ~n6896;
  assign n6898 = n831 & ~n6897;
  assign n6899 = n835 & ~n6898;
  assign n6900 = n839 & ~n6899;
  assign n6901 = n843 & ~n6900;
  assign n6902 = n847 & ~n6901;
  assign n6903 = n851 & ~n6902;
  assign n6904 = n855 & ~n6903;
  assign n6905 = n859 & ~n6904;
  assign n6906 = n863 & ~n6905;
  assign n6907 = n867 & ~n6906;
  assign n6908 = n871 & ~n6907;
  assign n6909 = n875 & ~n6908;
  assign n6910 = n879 & ~n6909;
  assign n6911 = n883 & ~n6910;
  assign n6912 = n887 & ~n6911;
  assign n6913 = n891 & ~n6912;
  assign n6914 = pi194  & ~n893;
  assign po66  = ~n6913 & n6914;
  assign n6916 = n902 & ~n1235;
  assign n6917 = n907 & ~n6916;
  assign n6918 = n911 & ~n6917;
  assign n6919 = n915 & ~n6918;
  assign n6920 = n919 & ~n6919;
  assign n6921 = n923 & ~n6920;
  assign n6922 = n927 & ~n6921;
  assign n6923 = n931 & ~n6922;
  assign n6924 = n935 & ~n6923;
  assign n6925 = n939 & ~n6924;
  assign n6926 = n943 & ~n6925;
  assign n6927 = n947 & ~n6926;
  assign n6928 = n951 & ~n6927;
  assign n6929 = n955 & ~n6928;
  assign n6930 = n959 & ~n6929;
  assign n6931 = n963 & ~n6930;
  assign n6932 = n967 & ~n6931;
  assign n6933 = n971 & ~n6932;
  assign n6934 = n975 & ~n6933;
  assign n6935 = n979 & ~n6934;
  assign n6936 = n983 & ~n6935;
  assign n6937 = n987 & ~n6936;
  assign n6938 = n991 & ~n6937;
  assign n6939 = n995 & ~n6938;
  assign n6940 = n999 & ~n6939;
  assign n6941 = n1003 & ~n6940;
  assign n6942 = n1007 & ~n6941;
  assign n6943 = n1011 & ~n6942;
  assign n6944 = n1015 & ~n6943;
  assign n6945 = n1019 & ~n6944;
  assign n6946 = n1023 & ~n6945;
  assign n6947 = n1027 & ~n6946;
  assign n6948 = n1031 & ~n6947;
  assign n6949 = n1035 & ~n6948;
  assign n6950 = n1039 & ~n6949;
  assign n6951 = n1043 & ~n6950;
  assign n6952 = n1047 & ~n6951;
  assign n6953 = n1051 & ~n6952;
  assign n6954 = n1055 & ~n6953;
  assign n6955 = n1059 & ~n6954;
  assign n6956 = n1574 & ~n6955;
  assign n6957 = n1576 & ~n6956;
  assign n6958 = n1837 & ~n6957;
  assign n6959 = n1068 & ~n6958;
  assign n6960 = n1072 & ~n6959;
  assign n6961 = n1076 & ~n6960;
  assign n6962 = n1080 & ~n6961;
  assign n6963 = n1084 & ~n6962;
  assign n6964 = n1088 & ~n6963;
  assign n6965 = n1092 & ~n6964;
  assign n6966 = n1096 & ~n6965;
  assign n6967 = n1100 & ~n6966;
  assign n6968 = n1104 & ~n6967;
  assign n6969 = n1108 & ~n6968;
  assign n6970 = n1112 & ~n6969;
  assign n6971 = n1116 & ~n6970;
  assign n6972 = n1120 & ~n6971;
  assign n6973 = n1124 & ~n6972;
  assign n6974 = n1128 & ~n6973;
  assign n6975 = n1132 & ~n6974;
  assign n6976 = n1136 & ~n6975;
  assign n6977 = n1140 & ~n6976;
  assign n6978 = n1144 & ~n6977;
  assign n6979 = n1148 & ~n6978;
  assign n6980 = n1152 & ~n6979;
  assign n6981 = n1156 & ~n6980;
  assign n6982 = n1160 & ~n6981;
  assign n6983 = n1164 & ~n6982;
  assign n6984 = n1168 & ~n6983;
  assign n6985 = n1172 & ~n6984;
  assign n6986 = n1176 & ~n6985;
  assign n6987 = n1180 & ~n6986;
  assign n6988 = n1184 & ~n6987;
  assign n6989 = n1188 & ~n6988;
  assign n6990 = n1192 & ~n6989;
  assign n6991 = n1196 & ~n6990;
  assign n6992 = n1200 & ~n6991;
  assign n6993 = n1204 & ~n6992;
  assign n6994 = n1208 & ~n6993;
  assign n6995 = n1212 & ~n6994;
  assign n6996 = n1216 & ~n6995;
  assign n6997 = n1220 & ~n6996;
  assign n6998 = n1224 & ~n6997;
  assign n6999 = n1228 & ~n6998;
  assign n7000 = pi195  & ~n1230;
  assign po67  = ~n6999 & n7000;
  assign n7002 = ~n567 & n1239;
  assign n7003 = n1244 & ~n7002;
  assign n7004 = n1248 & ~n7003;
  assign n7005 = n1252 & ~n7004;
  assign n7006 = n1256 & ~n7005;
  assign n7007 = n1260 & ~n7006;
  assign n7008 = n1264 & ~n7007;
  assign n7009 = n1268 & ~n7008;
  assign n7010 = n1272 & ~n7009;
  assign n7011 = n1276 & ~n7010;
  assign n7012 = n1280 & ~n7011;
  assign n7013 = n1284 & ~n7012;
  assign n7014 = n1288 & ~n7013;
  assign n7015 = n1292 & ~n7014;
  assign n7016 = n1296 & ~n7015;
  assign n7017 = n1300 & ~n7016;
  assign n7018 = n1304 & ~n7017;
  assign n7019 = n1308 & ~n7018;
  assign n7020 = n1312 & ~n7019;
  assign n7021 = n1316 & ~n7020;
  assign n7022 = n1320 & ~n7021;
  assign n7023 = n1324 & ~n7022;
  assign n7024 = n1328 & ~n7023;
  assign n7025 = n1332 & ~n7024;
  assign n7026 = n1336 & ~n7025;
  assign n7027 = n1340 & ~n7026;
  assign n7028 = n1344 & ~n7027;
  assign n7029 = n1348 & ~n7028;
  assign n7030 = n1352 & ~n7029;
  assign n7031 = n1356 & ~n7030;
  assign n7032 = n1360 & ~n7031;
  assign n7033 = n1364 & ~n7032;
  assign n7034 = n1368 & ~n7033;
  assign n7035 = n1372 & ~n7034;
  assign n7036 = n1376 & ~n7035;
  assign n7037 = n1380 & ~n7036;
  assign n7038 = n1384 & ~n7037;
  assign n7039 = n1388 & ~n7038;
  assign n7040 = n1392 & ~n7039;
  assign n7041 = n1396 & ~n7040;
  assign n7042 = n1663 & ~n7041;
  assign n7043 = n392 & ~n7042;
  assign n7044 = n396 & ~n7043;
  assign n7045 = n400 & ~n7044;
  assign n7046 = n404 & ~n7045;
  assign n7047 = n408 & ~n7046;
  assign n7048 = n412 & ~n7047;
  assign n7049 = n416 & ~n7048;
  assign n7050 = n420 & ~n7049;
  assign n7051 = n424 & ~n7050;
  assign n7052 = n428 & ~n7051;
  assign n7053 = n432 & ~n7052;
  assign n7054 = n436 & ~n7053;
  assign n7055 = n440 & ~n7054;
  assign n7056 = n444 & ~n7055;
  assign n7057 = n448 & ~n7056;
  assign n7058 = n452 & ~n7057;
  assign n7059 = n456 & ~n7058;
  assign n7060 = n460 & ~n7059;
  assign n7061 = n464 & ~n7060;
  assign n7062 = n468 & ~n7061;
  assign n7063 = n472 & ~n7062;
  assign n7064 = n476 & ~n7063;
  assign n7065 = n480 & ~n7064;
  assign n7066 = n484 & ~n7065;
  assign n7067 = n488 & ~n7066;
  assign n7068 = n492 & ~n7067;
  assign n7069 = n496 & ~n7068;
  assign n7070 = n500 & ~n7069;
  assign n7071 = n504 & ~n7070;
  assign n7072 = n508 & ~n7071;
  assign n7073 = n512 & ~n7072;
  assign n7074 = n516 & ~n7073;
  assign n7075 = n520 & ~n7074;
  assign n7076 = n524 & ~n7075;
  assign n7077 = n528 & ~n7076;
  assign n7078 = n532 & ~n7077;
  assign n7079 = n536 & ~n7078;
  assign n7080 = n540 & ~n7079;
  assign n7081 = n544 & ~n7080;
  assign n7082 = n548 & ~n7081;
  assign n7083 = n552 & ~n7082;
  assign n7084 = n556 & ~n7083;
  assign n7085 = n560 & ~n7084;
  assign n7086 = pi196  & ~n562;
  assign po68  = ~n7085 & n7086;
  assign n7088 = n571 & ~n906;
  assign n7089 = n576 & ~n7088;
  assign n7090 = n580 & ~n7089;
  assign n7091 = n584 & ~n7090;
  assign n7092 = n588 & ~n7091;
  assign n7093 = n592 & ~n7092;
  assign n7094 = n596 & ~n7093;
  assign n7095 = n600 & ~n7094;
  assign n7096 = n604 & ~n7095;
  assign n7097 = n608 & ~n7096;
  assign n7098 = n612 & ~n7097;
  assign n7099 = n616 & ~n7098;
  assign n7100 = n620 & ~n7099;
  assign n7101 = n624 & ~n7100;
  assign n7102 = n628 & ~n7101;
  assign n7103 = n632 & ~n7102;
  assign n7104 = n636 & ~n7103;
  assign n7105 = n640 & ~n7104;
  assign n7106 = n644 & ~n7105;
  assign n7107 = n648 & ~n7106;
  assign n7108 = n652 & ~n7107;
  assign n7109 = n656 & ~n7108;
  assign n7110 = n660 & ~n7109;
  assign n7111 = n664 & ~n7110;
  assign n7112 = n668 & ~n7111;
  assign n7113 = n672 & ~n7112;
  assign n7114 = n676 & ~n7113;
  assign n7115 = n680 & ~n7114;
  assign n7116 = n684 & ~n7115;
  assign n7117 = n688 & ~n7116;
  assign n7118 = n692 & ~n7117;
  assign n7119 = n696 & ~n7118;
  assign n7120 = n700 & ~n7119;
  assign n7121 = n704 & ~n7120;
  assign n7122 = n708 & ~n7121;
  assign n7123 = n712 & ~n7122;
  assign n7124 = n716 & ~n7123;
  assign n7125 = n720 & ~n7124;
  assign n7126 = n1484 & ~n7125;
  assign n7127 = n1486 & ~n7126;
  assign n7128 = n1750 & ~n7127;
  assign n7129 = n731 & ~n7128;
  assign n7130 = n735 & ~n7129;
  assign n7131 = n739 & ~n7130;
  assign n7132 = n743 & ~n7131;
  assign n7133 = n747 & ~n7132;
  assign n7134 = n751 & ~n7133;
  assign n7135 = n755 & ~n7134;
  assign n7136 = n759 & ~n7135;
  assign n7137 = n763 & ~n7136;
  assign n7138 = n767 & ~n7137;
  assign n7139 = n771 & ~n7138;
  assign n7140 = n775 & ~n7139;
  assign n7141 = n779 & ~n7140;
  assign n7142 = n783 & ~n7141;
  assign n7143 = n787 & ~n7142;
  assign n7144 = n791 & ~n7143;
  assign n7145 = n795 & ~n7144;
  assign n7146 = n799 & ~n7145;
  assign n7147 = n803 & ~n7146;
  assign n7148 = n807 & ~n7147;
  assign n7149 = n811 & ~n7148;
  assign n7150 = n815 & ~n7149;
  assign n7151 = n819 & ~n7150;
  assign n7152 = n823 & ~n7151;
  assign n7153 = n827 & ~n7152;
  assign n7154 = n831 & ~n7153;
  assign n7155 = n835 & ~n7154;
  assign n7156 = n839 & ~n7155;
  assign n7157 = n843 & ~n7156;
  assign n7158 = n847 & ~n7157;
  assign n7159 = n851 & ~n7158;
  assign n7160 = n855 & ~n7159;
  assign n7161 = n859 & ~n7160;
  assign n7162 = n863 & ~n7161;
  assign n7163 = n867 & ~n7162;
  assign n7164 = n871 & ~n7163;
  assign n7165 = n875 & ~n7164;
  assign n7166 = n879 & ~n7165;
  assign n7167 = n883 & ~n7166;
  assign n7168 = n887 & ~n7167;
  assign n7169 = n891 & ~n7168;
  assign n7170 = n895 & ~n7169;
  assign n7171 = n899 & ~n7170;
  assign n7172 = pi197  & ~n901;
  assign po69  = ~n7171 & n7172;
  assign n7174 = n910 & ~n1243;
  assign n7175 = n915 & ~n7174;
  assign n7176 = n919 & ~n7175;
  assign n7177 = n923 & ~n7176;
  assign n7178 = n927 & ~n7177;
  assign n7179 = n931 & ~n7178;
  assign n7180 = n935 & ~n7179;
  assign n7181 = n939 & ~n7180;
  assign n7182 = n943 & ~n7181;
  assign n7183 = n947 & ~n7182;
  assign n7184 = n951 & ~n7183;
  assign n7185 = n955 & ~n7184;
  assign n7186 = n959 & ~n7185;
  assign n7187 = n963 & ~n7186;
  assign n7188 = n967 & ~n7187;
  assign n7189 = n971 & ~n7188;
  assign n7190 = n975 & ~n7189;
  assign n7191 = n979 & ~n7190;
  assign n7192 = n983 & ~n7191;
  assign n7193 = n987 & ~n7192;
  assign n7194 = n991 & ~n7193;
  assign n7195 = n995 & ~n7194;
  assign n7196 = n999 & ~n7195;
  assign n7197 = n1003 & ~n7196;
  assign n7198 = n1007 & ~n7197;
  assign n7199 = n1011 & ~n7198;
  assign n7200 = n1015 & ~n7199;
  assign n7201 = n1019 & ~n7200;
  assign n7202 = n1023 & ~n7201;
  assign n7203 = n1027 & ~n7202;
  assign n7204 = n1031 & ~n7203;
  assign n7205 = n1035 & ~n7204;
  assign n7206 = n1039 & ~n7205;
  assign n7207 = n1043 & ~n7206;
  assign n7208 = n1047 & ~n7207;
  assign n7209 = n1051 & ~n7208;
  assign n7210 = n1055 & ~n7209;
  assign n7211 = n1059 & ~n7210;
  assign n7212 = n1574 & ~n7211;
  assign n7213 = n1576 & ~n7212;
  assign n7214 = n1837 & ~n7213;
  assign n7215 = n1068 & ~n7214;
  assign n7216 = n1072 & ~n7215;
  assign n7217 = n1076 & ~n7216;
  assign n7218 = n1080 & ~n7217;
  assign n7219 = n1084 & ~n7218;
  assign n7220 = n1088 & ~n7219;
  assign n7221 = n1092 & ~n7220;
  assign n7222 = n1096 & ~n7221;
  assign n7223 = n1100 & ~n7222;
  assign n7224 = n1104 & ~n7223;
  assign n7225 = n1108 & ~n7224;
  assign n7226 = n1112 & ~n7225;
  assign n7227 = n1116 & ~n7226;
  assign n7228 = n1120 & ~n7227;
  assign n7229 = n1124 & ~n7228;
  assign n7230 = n1128 & ~n7229;
  assign n7231 = n1132 & ~n7230;
  assign n7232 = n1136 & ~n7231;
  assign n7233 = n1140 & ~n7232;
  assign n7234 = n1144 & ~n7233;
  assign n7235 = n1148 & ~n7234;
  assign n7236 = n1152 & ~n7235;
  assign n7237 = n1156 & ~n7236;
  assign n7238 = n1160 & ~n7237;
  assign n7239 = n1164 & ~n7238;
  assign n7240 = n1168 & ~n7239;
  assign n7241 = n1172 & ~n7240;
  assign n7242 = n1176 & ~n7241;
  assign n7243 = n1180 & ~n7242;
  assign n7244 = n1184 & ~n7243;
  assign n7245 = n1188 & ~n7244;
  assign n7246 = n1192 & ~n7245;
  assign n7247 = n1196 & ~n7246;
  assign n7248 = n1200 & ~n7247;
  assign n7249 = n1204 & ~n7248;
  assign n7250 = n1208 & ~n7249;
  assign n7251 = n1212 & ~n7250;
  assign n7252 = n1216 & ~n7251;
  assign n7253 = n1220 & ~n7252;
  assign n7254 = n1224 & ~n7253;
  assign n7255 = n1228 & ~n7254;
  assign n7256 = n1232 & ~n7255;
  assign n7257 = n1236 & ~n7256;
  assign n7258 = pi198  & ~n1238;
  assign po70  = ~n7257 & n7258;
  assign n7260 = ~n575 & n1247;
  assign n7261 = n1252 & ~n7260;
  assign n7262 = n1256 & ~n7261;
  assign n7263 = n1260 & ~n7262;
  assign n7264 = n1264 & ~n7263;
  assign n7265 = n1268 & ~n7264;
  assign n7266 = n1272 & ~n7265;
  assign n7267 = n1276 & ~n7266;
  assign n7268 = n1280 & ~n7267;
  assign n7269 = n1284 & ~n7268;
  assign n7270 = n1288 & ~n7269;
  assign n7271 = n1292 & ~n7270;
  assign n7272 = n1296 & ~n7271;
  assign n7273 = n1300 & ~n7272;
  assign n7274 = n1304 & ~n7273;
  assign n7275 = n1308 & ~n7274;
  assign n7276 = n1312 & ~n7275;
  assign n7277 = n1316 & ~n7276;
  assign n7278 = n1320 & ~n7277;
  assign n7279 = n1324 & ~n7278;
  assign n7280 = n1328 & ~n7279;
  assign n7281 = n1332 & ~n7280;
  assign n7282 = n1336 & ~n7281;
  assign n7283 = n1340 & ~n7282;
  assign n7284 = n1344 & ~n7283;
  assign n7285 = n1348 & ~n7284;
  assign n7286 = n1352 & ~n7285;
  assign n7287 = n1356 & ~n7286;
  assign n7288 = n1360 & ~n7287;
  assign n7289 = n1364 & ~n7288;
  assign n7290 = n1368 & ~n7289;
  assign n7291 = n1372 & ~n7290;
  assign n7292 = n1376 & ~n7291;
  assign n7293 = n1380 & ~n7292;
  assign n7294 = n1384 & ~n7293;
  assign n7295 = n1388 & ~n7294;
  assign n7296 = n1392 & ~n7295;
  assign n7297 = n1396 & ~n7296;
  assign n7298 = n1663 & ~n7297;
  assign n7299 = n392 & ~n7298;
  assign n7300 = n396 & ~n7299;
  assign n7301 = n400 & ~n7300;
  assign n7302 = n404 & ~n7301;
  assign n7303 = n408 & ~n7302;
  assign n7304 = n412 & ~n7303;
  assign n7305 = n416 & ~n7304;
  assign n7306 = n420 & ~n7305;
  assign n7307 = n424 & ~n7306;
  assign n7308 = n428 & ~n7307;
  assign n7309 = n432 & ~n7308;
  assign n7310 = n436 & ~n7309;
  assign n7311 = n440 & ~n7310;
  assign n7312 = n444 & ~n7311;
  assign n7313 = n448 & ~n7312;
  assign n7314 = n452 & ~n7313;
  assign n7315 = n456 & ~n7314;
  assign n7316 = n460 & ~n7315;
  assign n7317 = n464 & ~n7316;
  assign n7318 = n468 & ~n7317;
  assign n7319 = n472 & ~n7318;
  assign n7320 = n476 & ~n7319;
  assign n7321 = n480 & ~n7320;
  assign n7322 = n484 & ~n7321;
  assign n7323 = n488 & ~n7322;
  assign n7324 = n492 & ~n7323;
  assign n7325 = n496 & ~n7324;
  assign n7326 = n500 & ~n7325;
  assign n7327 = n504 & ~n7326;
  assign n7328 = n508 & ~n7327;
  assign n7329 = n512 & ~n7328;
  assign n7330 = n516 & ~n7329;
  assign n7331 = n520 & ~n7330;
  assign n7332 = n524 & ~n7331;
  assign n7333 = n528 & ~n7332;
  assign n7334 = n532 & ~n7333;
  assign n7335 = n536 & ~n7334;
  assign n7336 = n540 & ~n7335;
  assign n7337 = n544 & ~n7336;
  assign n7338 = n548 & ~n7337;
  assign n7339 = n552 & ~n7338;
  assign n7340 = n556 & ~n7339;
  assign n7341 = n560 & ~n7340;
  assign n7342 = n564 & ~n7341;
  assign n7343 = n568 & ~n7342;
  assign n7344 = pi199  & ~n570;
  assign po71  = ~n7343 & n7344;
  assign n7346 = n579 & ~n914;
  assign n7347 = n584 & ~n7346;
  assign n7348 = n588 & ~n7347;
  assign n7349 = n592 & ~n7348;
  assign n7350 = n596 & ~n7349;
  assign n7351 = n600 & ~n7350;
  assign n7352 = n604 & ~n7351;
  assign n7353 = n608 & ~n7352;
  assign n7354 = n612 & ~n7353;
  assign n7355 = n616 & ~n7354;
  assign n7356 = n620 & ~n7355;
  assign n7357 = n624 & ~n7356;
  assign n7358 = n628 & ~n7357;
  assign n7359 = n632 & ~n7358;
  assign n7360 = n636 & ~n7359;
  assign n7361 = n640 & ~n7360;
  assign n7362 = n644 & ~n7361;
  assign n7363 = n648 & ~n7362;
  assign n7364 = n652 & ~n7363;
  assign n7365 = n656 & ~n7364;
  assign n7366 = n660 & ~n7365;
  assign n7367 = n664 & ~n7366;
  assign n7368 = n668 & ~n7367;
  assign n7369 = n672 & ~n7368;
  assign n7370 = n676 & ~n7369;
  assign n7371 = n680 & ~n7370;
  assign n7372 = n684 & ~n7371;
  assign n7373 = n688 & ~n7372;
  assign n7374 = n692 & ~n7373;
  assign n7375 = n696 & ~n7374;
  assign n7376 = n700 & ~n7375;
  assign n7377 = n704 & ~n7376;
  assign n7378 = n708 & ~n7377;
  assign n7379 = n712 & ~n7378;
  assign n7380 = n716 & ~n7379;
  assign n7381 = n720 & ~n7380;
  assign n7382 = n1484 & ~n7381;
  assign n7383 = n1486 & ~n7382;
  assign n7384 = n1750 & ~n7383;
  assign n7385 = n731 & ~n7384;
  assign n7386 = n735 & ~n7385;
  assign n7387 = n739 & ~n7386;
  assign n7388 = n743 & ~n7387;
  assign n7389 = n747 & ~n7388;
  assign n7390 = n751 & ~n7389;
  assign n7391 = n755 & ~n7390;
  assign n7392 = n759 & ~n7391;
  assign n7393 = n763 & ~n7392;
  assign n7394 = n767 & ~n7393;
  assign n7395 = n771 & ~n7394;
  assign n7396 = n775 & ~n7395;
  assign n7397 = n779 & ~n7396;
  assign n7398 = n783 & ~n7397;
  assign n7399 = n787 & ~n7398;
  assign n7400 = n791 & ~n7399;
  assign n7401 = n795 & ~n7400;
  assign n7402 = n799 & ~n7401;
  assign n7403 = n803 & ~n7402;
  assign n7404 = n807 & ~n7403;
  assign n7405 = n811 & ~n7404;
  assign n7406 = n815 & ~n7405;
  assign n7407 = n819 & ~n7406;
  assign n7408 = n823 & ~n7407;
  assign n7409 = n827 & ~n7408;
  assign n7410 = n831 & ~n7409;
  assign n7411 = n835 & ~n7410;
  assign n7412 = n839 & ~n7411;
  assign n7413 = n843 & ~n7412;
  assign n7414 = n847 & ~n7413;
  assign n7415 = n851 & ~n7414;
  assign n7416 = n855 & ~n7415;
  assign n7417 = n859 & ~n7416;
  assign n7418 = n863 & ~n7417;
  assign n7419 = n867 & ~n7418;
  assign n7420 = n871 & ~n7419;
  assign n7421 = n875 & ~n7420;
  assign n7422 = n879 & ~n7421;
  assign n7423 = n883 & ~n7422;
  assign n7424 = n887 & ~n7423;
  assign n7425 = n891 & ~n7424;
  assign n7426 = n895 & ~n7425;
  assign n7427 = n899 & ~n7426;
  assign n7428 = n903 & ~n7427;
  assign n7429 = n907 & ~n7428;
  assign n7430 = pi200  & ~n909;
  assign po72  = ~n7429 & n7430;
  assign n7432 = n918 & ~n1251;
  assign n7433 = n923 & ~n7432;
  assign n7434 = n927 & ~n7433;
  assign n7435 = n931 & ~n7434;
  assign n7436 = n935 & ~n7435;
  assign n7437 = n939 & ~n7436;
  assign n7438 = n943 & ~n7437;
  assign n7439 = n947 & ~n7438;
  assign n7440 = n951 & ~n7439;
  assign n7441 = n955 & ~n7440;
  assign n7442 = n959 & ~n7441;
  assign n7443 = n963 & ~n7442;
  assign n7444 = n967 & ~n7443;
  assign n7445 = n971 & ~n7444;
  assign n7446 = n975 & ~n7445;
  assign n7447 = n979 & ~n7446;
  assign n7448 = n983 & ~n7447;
  assign n7449 = n987 & ~n7448;
  assign n7450 = n991 & ~n7449;
  assign n7451 = n995 & ~n7450;
  assign n7452 = n999 & ~n7451;
  assign n7453 = n1003 & ~n7452;
  assign n7454 = n1007 & ~n7453;
  assign n7455 = n1011 & ~n7454;
  assign n7456 = n1015 & ~n7455;
  assign n7457 = n1019 & ~n7456;
  assign n7458 = n1023 & ~n7457;
  assign n7459 = n1027 & ~n7458;
  assign n7460 = n1031 & ~n7459;
  assign n7461 = n1035 & ~n7460;
  assign n7462 = n1039 & ~n7461;
  assign n7463 = n1043 & ~n7462;
  assign n7464 = n1047 & ~n7463;
  assign n7465 = n1051 & ~n7464;
  assign n7466 = n1055 & ~n7465;
  assign n7467 = n1059 & ~n7466;
  assign n7468 = n1574 & ~n7467;
  assign n7469 = n1576 & ~n7468;
  assign n7470 = n1837 & ~n7469;
  assign n7471 = n1068 & ~n7470;
  assign n7472 = n1072 & ~n7471;
  assign n7473 = n1076 & ~n7472;
  assign n7474 = n1080 & ~n7473;
  assign n7475 = n1084 & ~n7474;
  assign n7476 = n1088 & ~n7475;
  assign n7477 = n1092 & ~n7476;
  assign n7478 = n1096 & ~n7477;
  assign n7479 = n1100 & ~n7478;
  assign n7480 = n1104 & ~n7479;
  assign n7481 = n1108 & ~n7480;
  assign n7482 = n1112 & ~n7481;
  assign n7483 = n1116 & ~n7482;
  assign n7484 = n1120 & ~n7483;
  assign n7485 = n1124 & ~n7484;
  assign n7486 = n1128 & ~n7485;
  assign n7487 = n1132 & ~n7486;
  assign n7488 = n1136 & ~n7487;
  assign n7489 = n1140 & ~n7488;
  assign n7490 = n1144 & ~n7489;
  assign n7491 = n1148 & ~n7490;
  assign n7492 = n1152 & ~n7491;
  assign n7493 = n1156 & ~n7492;
  assign n7494 = n1160 & ~n7493;
  assign n7495 = n1164 & ~n7494;
  assign n7496 = n1168 & ~n7495;
  assign n7497 = n1172 & ~n7496;
  assign n7498 = n1176 & ~n7497;
  assign n7499 = n1180 & ~n7498;
  assign n7500 = n1184 & ~n7499;
  assign n7501 = n1188 & ~n7500;
  assign n7502 = n1192 & ~n7501;
  assign n7503 = n1196 & ~n7502;
  assign n7504 = n1200 & ~n7503;
  assign n7505 = n1204 & ~n7504;
  assign n7506 = n1208 & ~n7505;
  assign n7507 = n1212 & ~n7506;
  assign n7508 = n1216 & ~n7507;
  assign n7509 = n1220 & ~n7508;
  assign n7510 = n1224 & ~n7509;
  assign n7511 = n1228 & ~n7510;
  assign n7512 = n1232 & ~n7511;
  assign n7513 = n1236 & ~n7512;
  assign n7514 = n1240 & ~n7513;
  assign n7515 = n1244 & ~n7514;
  assign n7516 = pi201  & ~n1246;
  assign po73  = ~n7515 & n7516;
  assign n7518 = ~n583 & n1255;
  assign n7519 = n1260 & ~n7518;
  assign n7520 = n1264 & ~n7519;
  assign n7521 = n1268 & ~n7520;
  assign n7522 = n1272 & ~n7521;
  assign n7523 = n1276 & ~n7522;
  assign n7524 = n1280 & ~n7523;
  assign n7525 = n1284 & ~n7524;
  assign n7526 = n1288 & ~n7525;
  assign n7527 = n1292 & ~n7526;
  assign n7528 = n1296 & ~n7527;
  assign n7529 = n1300 & ~n7528;
  assign n7530 = n1304 & ~n7529;
  assign n7531 = n1308 & ~n7530;
  assign n7532 = n1312 & ~n7531;
  assign n7533 = n1316 & ~n7532;
  assign n7534 = n1320 & ~n7533;
  assign n7535 = n1324 & ~n7534;
  assign n7536 = n1328 & ~n7535;
  assign n7537 = n1332 & ~n7536;
  assign n7538 = n1336 & ~n7537;
  assign n7539 = n1340 & ~n7538;
  assign n7540 = n1344 & ~n7539;
  assign n7541 = n1348 & ~n7540;
  assign n7542 = n1352 & ~n7541;
  assign n7543 = n1356 & ~n7542;
  assign n7544 = n1360 & ~n7543;
  assign n7545 = n1364 & ~n7544;
  assign n7546 = n1368 & ~n7545;
  assign n7547 = n1372 & ~n7546;
  assign n7548 = n1376 & ~n7547;
  assign n7549 = n1380 & ~n7548;
  assign n7550 = n1384 & ~n7549;
  assign n7551 = n1388 & ~n7550;
  assign n7552 = n1392 & ~n7551;
  assign n7553 = n1396 & ~n7552;
  assign n7554 = n1663 & ~n7553;
  assign n7555 = n392 & ~n7554;
  assign n7556 = n396 & ~n7555;
  assign n7557 = n400 & ~n7556;
  assign n7558 = n404 & ~n7557;
  assign n7559 = n408 & ~n7558;
  assign n7560 = n412 & ~n7559;
  assign n7561 = n416 & ~n7560;
  assign n7562 = n420 & ~n7561;
  assign n7563 = n424 & ~n7562;
  assign n7564 = n428 & ~n7563;
  assign n7565 = n432 & ~n7564;
  assign n7566 = n436 & ~n7565;
  assign n7567 = n440 & ~n7566;
  assign n7568 = n444 & ~n7567;
  assign n7569 = n448 & ~n7568;
  assign n7570 = n452 & ~n7569;
  assign n7571 = n456 & ~n7570;
  assign n7572 = n460 & ~n7571;
  assign n7573 = n464 & ~n7572;
  assign n7574 = n468 & ~n7573;
  assign n7575 = n472 & ~n7574;
  assign n7576 = n476 & ~n7575;
  assign n7577 = n480 & ~n7576;
  assign n7578 = n484 & ~n7577;
  assign n7579 = n488 & ~n7578;
  assign n7580 = n492 & ~n7579;
  assign n7581 = n496 & ~n7580;
  assign n7582 = n500 & ~n7581;
  assign n7583 = n504 & ~n7582;
  assign n7584 = n508 & ~n7583;
  assign n7585 = n512 & ~n7584;
  assign n7586 = n516 & ~n7585;
  assign n7587 = n520 & ~n7586;
  assign n7588 = n524 & ~n7587;
  assign n7589 = n528 & ~n7588;
  assign n7590 = n532 & ~n7589;
  assign n7591 = n536 & ~n7590;
  assign n7592 = n540 & ~n7591;
  assign n7593 = n544 & ~n7592;
  assign n7594 = n548 & ~n7593;
  assign n7595 = n552 & ~n7594;
  assign n7596 = n556 & ~n7595;
  assign n7597 = n560 & ~n7596;
  assign n7598 = n564 & ~n7597;
  assign n7599 = n568 & ~n7598;
  assign n7600 = n572 & ~n7599;
  assign n7601 = n576 & ~n7600;
  assign n7602 = pi202  & ~n578;
  assign po74  = ~n7601 & n7602;
  assign n7604 = n587 & ~n922;
  assign n7605 = n592 & ~n7604;
  assign n7606 = n596 & ~n7605;
  assign n7607 = n600 & ~n7606;
  assign n7608 = n604 & ~n7607;
  assign n7609 = n608 & ~n7608;
  assign n7610 = n612 & ~n7609;
  assign n7611 = n616 & ~n7610;
  assign n7612 = n620 & ~n7611;
  assign n7613 = n624 & ~n7612;
  assign n7614 = n628 & ~n7613;
  assign n7615 = n632 & ~n7614;
  assign n7616 = n636 & ~n7615;
  assign n7617 = n640 & ~n7616;
  assign n7618 = n644 & ~n7617;
  assign n7619 = n648 & ~n7618;
  assign n7620 = n652 & ~n7619;
  assign n7621 = n656 & ~n7620;
  assign n7622 = n660 & ~n7621;
  assign n7623 = n664 & ~n7622;
  assign n7624 = n668 & ~n7623;
  assign n7625 = n672 & ~n7624;
  assign n7626 = n676 & ~n7625;
  assign n7627 = n680 & ~n7626;
  assign n7628 = n684 & ~n7627;
  assign n7629 = n688 & ~n7628;
  assign n7630 = n692 & ~n7629;
  assign n7631 = n696 & ~n7630;
  assign n7632 = n700 & ~n7631;
  assign n7633 = n704 & ~n7632;
  assign n7634 = n708 & ~n7633;
  assign n7635 = n712 & ~n7634;
  assign n7636 = n716 & ~n7635;
  assign n7637 = n720 & ~n7636;
  assign n7638 = n1484 & ~n7637;
  assign n7639 = n1486 & ~n7638;
  assign n7640 = n1750 & ~n7639;
  assign n7641 = n731 & ~n7640;
  assign n7642 = n735 & ~n7641;
  assign n7643 = n739 & ~n7642;
  assign n7644 = n743 & ~n7643;
  assign n7645 = n747 & ~n7644;
  assign n7646 = n751 & ~n7645;
  assign n7647 = n755 & ~n7646;
  assign n7648 = n759 & ~n7647;
  assign n7649 = n763 & ~n7648;
  assign n7650 = n767 & ~n7649;
  assign n7651 = n771 & ~n7650;
  assign n7652 = n775 & ~n7651;
  assign n7653 = n779 & ~n7652;
  assign n7654 = n783 & ~n7653;
  assign n7655 = n787 & ~n7654;
  assign n7656 = n791 & ~n7655;
  assign n7657 = n795 & ~n7656;
  assign n7658 = n799 & ~n7657;
  assign n7659 = n803 & ~n7658;
  assign n7660 = n807 & ~n7659;
  assign n7661 = n811 & ~n7660;
  assign n7662 = n815 & ~n7661;
  assign n7663 = n819 & ~n7662;
  assign n7664 = n823 & ~n7663;
  assign n7665 = n827 & ~n7664;
  assign n7666 = n831 & ~n7665;
  assign n7667 = n835 & ~n7666;
  assign n7668 = n839 & ~n7667;
  assign n7669 = n843 & ~n7668;
  assign n7670 = n847 & ~n7669;
  assign n7671 = n851 & ~n7670;
  assign n7672 = n855 & ~n7671;
  assign n7673 = n859 & ~n7672;
  assign n7674 = n863 & ~n7673;
  assign n7675 = n867 & ~n7674;
  assign n7676 = n871 & ~n7675;
  assign n7677 = n875 & ~n7676;
  assign n7678 = n879 & ~n7677;
  assign n7679 = n883 & ~n7678;
  assign n7680 = n887 & ~n7679;
  assign n7681 = n891 & ~n7680;
  assign n7682 = n895 & ~n7681;
  assign n7683 = n899 & ~n7682;
  assign n7684 = n903 & ~n7683;
  assign n7685 = n907 & ~n7684;
  assign n7686 = n911 & ~n7685;
  assign n7687 = n915 & ~n7686;
  assign n7688 = pi203  & ~n917;
  assign po75  = ~n7687 & n7688;
  assign n7690 = n926 & ~n1259;
  assign n7691 = n931 & ~n7690;
  assign n7692 = n935 & ~n7691;
  assign n7693 = n939 & ~n7692;
  assign n7694 = n943 & ~n7693;
  assign n7695 = n947 & ~n7694;
  assign n7696 = n951 & ~n7695;
  assign n7697 = n955 & ~n7696;
  assign n7698 = n959 & ~n7697;
  assign n7699 = n963 & ~n7698;
  assign n7700 = n967 & ~n7699;
  assign n7701 = n971 & ~n7700;
  assign n7702 = n975 & ~n7701;
  assign n7703 = n979 & ~n7702;
  assign n7704 = n983 & ~n7703;
  assign n7705 = n987 & ~n7704;
  assign n7706 = n991 & ~n7705;
  assign n7707 = n995 & ~n7706;
  assign n7708 = n999 & ~n7707;
  assign n7709 = n1003 & ~n7708;
  assign n7710 = n1007 & ~n7709;
  assign n7711 = n1011 & ~n7710;
  assign n7712 = n1015 & ~n7711;
  assign n7713 = n1019 & ~n7712;
  assign n7714 = n1023 & ~n7713;
  assign n7715 = n1027 & ~n7714;
  assign n7716 = n1031 & ~n7715;
  assign n7717 = n1035 & ~n7716;
  assign n7718 = n1039 & ~n7717;
  assign n7719 = n1043 & ~n7718;
  assign n7720 = n1047 & ~n7719;
  assign n7721 = n1051 & ~n7720;
  assign n7722 = n1055 & ~n7721;
  assign n7723 = n1059 & ~n7722;
  assign n7724 = n1574 & ~n7723;
  assign n7725 = n1576 & ~n7724;
  assign n7726 = n1837 & ~n7725;
  assign n7727 = n1068 & ~n7726;
  assign n7728 = n1072 & ~n7727;
  assign n7729 = n1076 & ~n7728;
  assign n7730 = n1080 & ~n7729;
  assign n7731 = n1084 & ~n7730;
  assign n7732 = n1088 & ~n7731;
  assign n7733 = n1092 & ~n7732;
  assign n7734 = n1096 & ~n7733;
  assign n7735 = n1100 & ~n7734;
  assign n7736 = n1104 & ~n7735;
  assign n7737 = n1108 & ~n7736;
  assign n7738 = n1112 & ~n7737;
  assign n7739 = n1116 & ~n7738;
  assign n7740 = n1120 & ~n7739;
  assign n7741 = n1124 & ~n7740;
  assign n7742 = n1128 & ~n7741;
  assign n7743 = n1132 & ~n7742;
  assign n7744 = n1136 & ~n7743;
  assign n7745 = n1140 & ~n7744;
  assign n7746 = n1144 & ~n7745;
  assign n7747 = n1148 & ~n7746;
  assign n7748 = n1152 & ~n7747;
  assign n7749 = n1156 & ~n7748;
  assign n7750 = n1160 & ~n7749;
  assign n7751 = n1164 & ~n7750;
  assign n7752 = n1168 & ~n7751;
  assign n7753 = n1172 & ~n7752;
  assign n7754 = n1176 & ~n7753;
  assign n7755 = n1180 & ~n7754;
  assign n7756 = n1184 & ~n7755;
  assign n7757 = n1188 & ~n7756;
  assign n7758 = n1192 & ~n7757;
  assign n7759 = n1196 & ~n7758;
  assign n7760 = n1200 & ~n7759;
  assign n7761 = n1204 & ~n7760;
  assign n7762 = n1208 & ~n7761;
  assign n7763 = n1212 & ~n7762;
  assign n7764 = n1216 & ~n7763;
  assign n7765 = n1220 & ~n7764;
  assign n7766 = n1224 & ~n7765;
  assign n7767 = n1228 & ~n7766;
  assign n7768 = n1232 & ~n7767;
  assign n7769 = n1236 & ~n7768;
  assign n7770 = n1240 & ~n7769;
  assign n7771 = n1244 & ~n7770;
  assign n7772 = n1248 & ~n7771;
  assign n7773 = n1252 & ~n7772;
  assign n7774 = pi204  & ~n1254;
  assign po76  = ~n7773 & n7774;
  assign n7776 = ~n591 & n1263;
  assign n7777 = n1268 & ~n7776;
  assign n7778 = n1272 & ~n7777;
  assign n7779 = n1276 & ~n7778;
  assign n7780 = n1280 & ~n7779;
  assign n7781 = n1284 & ~n7780;
  assign n7782 = n1288 & ~n7781;
  assign n7783 = n1292 & ~n7782;
  assign n7784 = n1296 & ~n7783;
  assign n7785 = n1300 & ~n7784;
  assign n7786 = n1304 & ~n7785;
  assign n7787 = n1308 & ~n7786;
  assign n7788 = n1312 & ~n7787;
  assign n7789 = n1316 & ~n7788;
  assign n7790 = n1320 & ~n7789;
  assign n7791 = n1324 & ~n7790;
  assign n7792 = n1328 & ~n7791;
  assign n7793 = n1332 & ~n7792;
  assign n7794 = n1336 & ~n7793;
  assign n7795 = n1340 & ~n7794;
  assign n7796 = n1344 & ~n7795;
  assign n7797 = n1348 & ~n7796;
  assign n7798 = n1352 & ~n7797;
  assign n7799 = n1356 & ~n7798;
  assign n7800 = n1360 & ~n7799;
  assign n7801 = n1364 & ~n7800;
  assign n7802 = n1368 & ~n7801;
  assign n7803 = n1372 & ~n7802;
  assign n7804 = n1376 & ~n7803;
  assign n7805 = n1380 & ~n7804;
  assign n7806 = n1384 & ~n7805;
  assign n7807 = n1388 & ~n7806;
  assign n7808 = n1392 & ~n7807;
  assign n7809 = n1396 & ~n7808;
  assign n7810 = n1663 & ~n7809;
  assign n7811 = n392 & ~n7810;
  assign n7812 = n396 & ~n7811;
  assign n7813 = n400 & ~n7812;
  assign n7814 = n404 & ~n7813;
  assign n7815 = n408 & ~n7814;
  assign n7816 = n412 & ~n7815;
  assign n7817 = n416 & ~n7816;
  assign n7818 = n420 & ~n7817;
  assign n7819 = n424 & ~n7818;
  assign n7820 = n428 & ~n7819;
  assign n7821 = n432 & ~n7820;
  assign n7822 = n436 & ~n7821;
  assign n7823 = n440 & ~n7822;
  assign n7824 = n444 & ~n7823;
  assign n7825 = n448 & ~n7824;
  assign n7826 = n452 & ~n7825;
  assign n7827 = n456 & ~n7826;
  assign n7828 = n460 & ~n7827;
  assign n7829 = n464 & ~n7828;
  assign n7830 = n468 & ~n7829;
  assign n7831 = n472 & ~n7830;
  assign n7832 = n476 & ~n7831;
  assign n7833 = n480 & ~n7832;
  assign n7834 = n484 & ~n7833;
  assign n7835 = n488 & ~n7834;
  assign n7836 = n492 & ~n7835;
  assign n7837 = n496 & ~n7836;
  assign n7838 = n500 & ~n7837;
  assign n7839 = n504 & ~n7838;
  assign n7840 = n508 & ~n7839;
  assign n7841 = n512 & ~n7840;
  assign n7842 = n516 & ~n7841;
  assign n7843 = n520 & ~n7842;
  assign n7844 = n524 & ~n7843;
  assign n7845 = n528 & ~n7844;
  assign n7846 = n532 & ~n7845;
  assign n7847 = n536 & ~n7846;
  assign n7848 = n540 & ~n7847;
  assign n7849 = n544 & ~n7848;
  assign n7850 = n548 & ~n7849;
  assign n7851 = n552 & ~n7850;
  assign n7852 = n556 & ~n7851;
  assign n7853 = n560 & ~n7852;
  assign n7854 = n564 & ~n7853;
  assign n7855 = n568 & ~n7854;
  assign n7856 = n572 & ~n7855;
  assign n7857 = n576 & ~n7856;
  assign n7858 = n580 & ~n7857;
  assign n7859 = n584 & ~n7858;
  assign n7860 = pi205  & ~n586;
  assign po77  = ~n7859 & n7860;
  assign n7862 = n595 & ~n930;
  assign n7863 = n600 & ~n7862;
  assign n7864 = n604 & ~n7863;
  assign n7865 = n608 & ~n7864;
  assign n7866 = n612 & ~n7865;
  assign n7867 = n616 & ~n7866;
  assign n7868 = n620 & ~n7867;
  assign n7869 = n624 & ~n7868;
  assign n7870 = n628 & ~n7869;
  assign n7871 = n632 & ~n7870;
  assign n7872 = n636 & ~n7871;
  assign n7873 = n640 & ~n7872;
  assign n7874 = n644 & ~n7873;
  assign n7875 = n648 & ~n7874;
  assign n7876 = n652 & ~n7875;
  assign n7877 = n656 & ~n7876;
  assign n7878 = n660 & ~n7877;
  assign n7879 = n664 & ~n7878;
  assign n7880 = n668 & ~n7879;
  assign n7881 = n672 & ~n7880;
  assign n7882 = n676 & ~n7881;
  assign n7883 = n680 & ~n7882;
  assign n7884 = n684 & ~n7883;
  assign n7885 = n688 & ~n7884;
  assign n7886 = n692 & ~n7885;
  assign n7887 = n696 & ~n7886;
  assign n7888 = n700 & ~n7887;
  assign n7889 = n704 & ~n7888;
  assign n7890 = n708 & ~n7889;
  assign n7891 = n712 & ~n7890;
  assign n7892 = n716 & ~n7891;
  assign n7893 = n720 & ~n7892;
  assign n7894 = n1484 & ~n7893;
  assign n7895 = n1486 & ~n7894;
  assign n7896 = n1750 & ~n7895;
  assign n7897 = n731 & ~n7896;
  assign n7898 = n735 & ~n7897;
  assign n7899 = n739 & ~n7898;
  assign n7900 = n743 & ~n7899;
  assign n7901 = n747 & ~n7900;
  assign n7902 = n751 & ~n7901;
  assign n7903 = n755 & ~n7902;
  assign n7904 = n759 & ~n7903;
  assign n7905 = n763 & ~n7904;
  assign n7906 = n767 & ~n7905;
  assign n7907 = n771 & ~n7906;
  assign n7908 = n775 & ~n7907;
  assign n7909 = n779 & ~n7908;
  assign n7910 = n783 & ~n7909;
  assign n7911 = n787 & ~n7910;
  assign n7912 = n791 & ~n7911;
  assign n7913 = n795 & ~n7912;
  assign n7914 = n799 & ~n7913;
  assign n7915 = n803 & ~n7914;
  assign n7916 = n807 & ~n7915;
  assign n7917 = n811 & ~n7916;
  assign n7918 = n815 & ~n7917;
  assign n7919 = n819 & ~n7918;
  assign n7920 = n823 & ~n7919;
  assign n7921 = n827 & ~n7920;
  assign n7922 = n831 & ~n7921;
  assign n7923 = n835 & ~n7922;
  assign n7924 = n839 & ~n7923;
  assign n7925 = n843 & ~n7924;
  assign n7926 = n847 & ~n7925;
  assign n7927 = n851 & ~n7926;
  assign n7928 = n855 & ~n7927;
  assign n7929 = n859 & ~n7928;
  assign n7930 = n863 & ~n7929;
  assign n7931 = n867 & ~n7930;
  assign n7932 = n871 & ~n7931;
  assign n7933 = n875 & ~n7932;
  assign n7934 = n879 & ~n7933;
  assign n7935 = n883 & ~n7934;
  assign n7936 = n887 & ~n7935;
  assign n7937 = n891 & ~n7936;
  assign n7938 = n895 & ~n7937;
  assign n7939 = n899 & ~n7938;
  assign n7940 = n903 & ~n7939;
  assign n7941 = n907 & ~n7940;
  assign n7942 = n911 & ~n7941;
  assign n7943 = n915 & ~n7942;
  assign n7944 = n919 & ~n7943;
  assign n7945 = n923 & ~n7944;
  assign n7946 = pi206  & ~n925;
  assign po78  = ~n7945 & n7946;
  assign n7948 = n934 & ~n1267;
  assign n7949 = n939 & ~n7948;
  assign n7950 = n943 & ~n7949;
  assign n7951 = n947 & ~n7950;
  assign n7952 = n951 & ~n7951;
  assign n7953 = n955 & ~n7952;
  assign n7954 = n959 & ~n7953;
  assign n7955 = n963 & ~n7954;
  assign n7956 = n967 & ~n7955;
  assign n7957 = n971 & ~n7956;
  assign n7958 = n975 & ~n7957;
  assign n7959 = n979 & ~n7958;
  assign n7960 = n983 & ~n7959;
  assign n7961 = n987 & ~n7960;
  assign n7962 = n991 & ~n7961;
  assign n7963 = n995 & ~n7962;
  assign n7964 = n999 & ~n7963;
  assign n7965 = n1003 & ~n7964;
  assign n7966 = n1007 & ~n7965;
  assign n7967 = n1011 & ~n7966;
  assign n7968 = n1015 & ~n7967;
  assign n7969 = n1019 & ~n7968;
  assign n7970 = n1023 & ~n7969;
  assign n7971 = n1027 & ~n7970;
  assign n7972 = n1031 & ~n7971;
  assign n7973 = n1035 & ~n7972;
  assign n7974 = n1039 & ~n7973;
  assign n7975 = n1043 & ~n7974;
  assign n7976 = n1047 & ~n7975;
  assign n7977 = n1051 & ~n7976;
  assign n7978 = n1055 & ~n7977;
  assign n7979 = n1059 & ~n7978;
  assign n7980 = n1574 & ~n7979;
  assign n7981 = n1576 & ~n7980;
  assign n7982 = n1837 & ~n7981;
  assign n7983 = n1068 & ~n7982;
  assign n7984 = n1072 & ~n7983;
  assign n7985 = n1076 & ~n7984;
  assign n7986 = n1080 & ~n7985;
  assign n7987 = n1084 & ~n7986;
  assign n7988 = n1088 & ~n7987;
  assign n7989 = n1092 & ~n7988;
  assign n7990 = n1096 & ~n7989;
  assign n7991 = n1100 & ~n7990;
  assign n7992 = n1104 & ~n7991;
  assign n7993 = n1108 & ~n7992;
  assign n7994 = n1112 & ~n7993;
  assign n7995 = n1116 & ~n7994;
  assign n7996 = n1120 & ~n7995;
  assign n7997 = n1124 & ~n7996;
  assign n7998 = n1128 & ~n7997;
  assign n7999 = n1132 & ~n7998;
  assign n8000 = n1136 & ~n7999;
  assign n8001 = n1140 & ~n8000;
  assign n8002 = n1144 & ~n8001;
  assign n8003 = n1148 & ~n8002;
  assign n8004 = n1152 & ~n8003;
  assign n8005 = n1156 & ~n8004;
  assign n8006 = n1160 & ~n8005;
  assign n8007 = n1164 & ~n8006;
  assign n8008 = n1168 & ~n8007;
  assign n8009 = n1172 & ~n8008;
  assign n8010 = n1176 & ~n8009;
  assign n8011 = n1180 & ~n8010;
  assign n8012 = n1184 & ~n8011;
  assign n8013 = n1188 & ~n8012;
  assign n8014 = n1192 & ~n8013;
  assign n8015 = n1196 & ~n8014;
  assign n8016 = n1200 & ~n8015;
  assign n8017 = n1204 & ~n8016;
  assign n8018 = n1208 & ~n8017;
  assign n8019 = n1212 & ~n8018;
  assign n8020 = n1216 & ~n8019;
  assign n8021 = n1220 & ~n8020;
  assign n8022 = n1224 & ~n8021;
  assign n8023 = n1228 & ~n8022;
  assign n8024 = n1232 & ~n8023;
  assign n8025 = n1236 & ~n8024;
  assign n8026 = n1240 & ~n8025;
  assign n8027 = n1244 & ~n8026;
  assign n8028 = n1248 & ~n8027;
  assign n8029 = n1252 & ~n8028;
  assign n8030 = n1256 & ~n8029;
  assign n8031 = n1260 & ~n8030;
  assign n8032 = pi207  & ~n1262;
  assign po79  = ~n8031 & n8032;
  assign n8034 = ~n599 & n1271;
  assign n8035 = n1276 & ~n8034;
  assign n8036 = n1280 & ~n8035;
  assign n8037 = n1284 & ~n8036;
  assign n8038 = n1288 & ~n8037;
  assign n8039 = n1292 & ~n8038;
  assign n8040 = n1296 & ~n8039;
  assign n8041 = n1300 & ~n8040;
  assign n8042 = n1304 & ~n8041;
  assign n8043 = n1308 & ~n8042;
  assign n8044 = n1312 & ~n8043;
  assign n8045 = n1316 & ~n8044;
  assign n8046 = n1320 & ~n8045;
  assign n8047 = n1324 & ~n8046;
  assign n8048 = n1328 & ~n8047;
  assign n8049 = n1332 & ~n8048;
  assign n8050 = n1336 & ~n8049;
  assign n8051 = n1340 & ~n8050;
  assign n8052 = n1344 & ~n8051;
  assign n8053 = n1348 & ~n8052;
  assign n8054 = n1352 & ~n8053;
  assign n8055 = n1356 & ~n8054;
  assign n8056 = n1360 & ~n8055;
  assign n8057 = n1364 & ~n8056;
  assign n8058 = n1368 & ~n8057;
  assign n8059 = n1372 & ~n8058;
  assign n8060 = n1376 & ~n8059;
  assign n8061 = n1380 & ~n8060;
  assign n8062 = n1384 & ~n8061;
  assign n8063 = n1388 & ~n8062;
  assign n8064 = n1392 & ~n8063;
  assign n8065 = n1396 & ~n8064;
  assign n8066 = n1663 & ~n8065;
  assign n8067 = n392 & ~n8066;
  assign n8068 = n396 & ~n8067;
  assign n8069 = n400 & ~n8068;
  assign n8070 = n404 & ~n8069;
  assign n8071 = n408 & ~n8070;
  assign n8072 = n412 & ~n8071;
  assign n8073 = n416 & ~n8072;
  assign n8074 = n420 & ~n8073;
  assign n8075 = n424 & ~n8074;
  assign n8076 = n428 & ~n8075;
  assign n8077 = n432 & ~n8076;
  assign n8078 = n436 & ~n8077;
  assign n8079 = n440 & ~n8078;
  assign n8080 = n444 & ~n8079;
  assign n8081 = n448 & ~n8080;
  assign n8082 = n452 & ~n8081;
  assign n8083 = n456 & ~n8082;
  assign n8084 = n460 & ~n8083;
  assign n8085 = n464 & ~n8084;
  assign n8086 = n468 & ~n8085;
  assign n8087 = n472 & ~n8086;
  assign n8088 = n476 & ~n8087;
  assign n8089 = n480 & ~n8088;
  assign n8090 = n484 & ~n8089;
  assign n8091 = n488 & ~n8090;
  assign n8092 = n492 & ~n8091;
  assign n8093 = n496 & ~n8092;
  assign n8094 = n500 & ~n8093;
  assign n8095 = n504 & ~n8094;
  assign n8096 = n508 & ~n8095;
  assign n8097 = n512 & ~n8096;
  assign n8098 = n516 & ~n8097;
  assign n8099 = n520 & ~n8098;
  assign n8100 = n524 & ~n8099;
  assign n8101 = n528 & ~n8100;
  assign n8102 = n532 & ~n8101;
  assign n8103 = n536 & ~n8102;
  assign n8104 = n540 & ~n8103;
  assign n8105 = n544 & ~n8104;
  assign n8106 = n548 & ~n8105;
  assign n8107 = n552 & ~n8106;
  assign n8108 = n556 & ~n8107;
  assign n8109 = n560 & ~n8108;
  assign n8110 = n564 & ~n8109;
  assign n8111 = n568 & ~n8110;
  assign n8112 = n572 & ~n8111;
  assign n8113 = n576 & ~n8112;
  assign n8114 = n580 & ~n8113;
  assign n8115 = n584 & ~n8114;
  assign n8116 = n588 & ~n8115;
  assign n8117 = n592 & ~n8116;
  assign n8118 = pi208  & ~n594;
  assign po80  = ~n8117 & n8118;
  assign n8120 = n603 & ~n938;
  assign n8121 = n608 & ~n8120;
  assign n8122 = n612 & ~n8121;
  assign n8123 = n616 & ~n8122;
  assign n8124 = n620 & ~n8123;
  assign n8125 = n624 & ~n8124;
  assign n8126 = n628 & ~n8125;
  assign n8127 = n632 & ~n8126;
  assign n8128 = n636 & ~n8127;
  assign n8129 = n640 & ~n8128;
  assign n8130 = n644 & ~n8129;
  assign n8131 = n648 & ~n8130;
  assign n8132 = n652 & ~n8131;
  assign n8133 = n656 & ~n8132;
  assign n8134 = n660 & ~n8133;
  assign n8135 = n664 & ~n8134;
  assign n8136 = n668 & ~n8135;
  assign n8137 = n672 & ~n8136;
  assign n8138 = n676 & ~n8137;
  assign n8139 = n680 & ~n8138;
  assign n8140 = n684 & ~n8139;
  assign n8141 = n688 & ~n8140;
  assign n8142 = n692 & ~n8141;
  assign n8143 = n696 & ~n8142;
  assign n8144 = n700 & ~n8143;
  assign n8145 = n704 & ~n8144;
  assign n8146 = n708 & ~n8145;
  assign n8147 = n712 & ~n8146;
  assign n8148 = n716 & ~n8147;
  assign n8149 = n720 & ~n8148;
  assign n8150 = n1484 & ~n8149;
  assign n8151 = n1486 & ~n8150;
  assign n8152 = n1750 & ~n8151;
  assign n8153 = n731 & ~n8152;
  assign n8154 = n735 & ~n8153;
  assign n8155 = n739 & ~n8154;
  assign n8156 = n743 & ~n8155;
  assign n8157 = n747 & ~n8156;
  assign n8158 = n751 & ~n8157;
  assign n8159 = n755 & ~n8158;
  assign n8160 = n759 & ~n8159;
  assign n8161 = n763 & ~n8160;
  assign n8162 = n767 & ~n8161;
  assign n8163 = n771 & ~n8162;
  assign n8164 = n775 & ~n8163;
  assign n8165 = n779 & ~n8164;
  assign n8166 = n783 & ~n8165;
  assign n8167 = n787 & ~n8166;
  assign n8168 = n791 & ~n8167;
  assign n8169 = n795 & ~n8168;
  assign n8170 = n799 & ~n8169;
  assign n8171 = n803 & ~n8170;
  assign n8172 = n807 & ~n8171;
  assign n8173 = n811 & ~n8172;
  assign n8174 = n815 & ~n8173;
  assign n8175 = n819 & ~n8174;
  assign n8176 = n823 & ~n8175;
  assign n8177 = n827 & ~n8176;
  assign n8178 = n831 & ~n8177;
  assign n8179 = n835 & ~n8178;
  assign n8180 = n839 & ~n8179;
  assign n8181 = n843 & ~n8180;
  assign n8182 = n847 & ~n8181;
  assign n8183 = n851 & ~n8182;
  assign n8184 = n855 & ~n8183;
  assign n8185 = n859 & ~n8184;
  assign n8186 = n863 & ~n8185;
  assign n8187 = n867 & ~n8186;
  assign n8188 = n871 & ~n8187;
  assign n8189 = n875 & ~n8188;
  assign n8190 = n879 & ~n8189;
  assign n8191 = n883 & ~n8190;
  assign n8192 = n887 & ~n8191;
  assign n8193 = n891 & ~n8192;
  assign n8194 = n895 & ~n8193;
  assign n8195 = n899 & ~n8194;
  assign n8196 = n903 & ~n8195;
  assign n8197 = n907 & ~n8196;
  assign n8198 = n911 & ~n8197;
  assign n8199 = n915 & ~n8198;
  assign n8200 = n919 & ~n8199;
  assign n8201 = n923 & ~n8200;
  assign n8202 = n927 & ~n8201;
  assign n8203 = n931 & ~n8202;
  assign n8204 = pi209  & ~n933;
  assign po81  = ~n8203 & n8204;
  assign n8206 = n942 & ~n1275;
  assign n8207 = n947 & ~n8206;
  assign n8208 = n951 & ~n8207;
  assign n8209 = n955 & ~n8208;
  assign n8210 = n959 & ~n8209;
  assign n8211 = n963 & ~n8210;
  assign n8212 = n967 & ~n8211;
  assign n8213 = n971 & ~n8212;
  assign n8214 = n975 & ~n8213;
  assign n8215 = n979 & ~n8214;
  assign n8216 = n983 & ~n8215;
  assign n8217 = n987 & ~n8216;
  assign n8218 = n991 & ~n8217;
  assign n8219 = n995 & ~n8218;
  assign n8220 = n999 & ~n8219;
  assign n8221 = n1003 & ~n8220;
  assign n8222 = n1007 & ~n8221;
  assign n8223 = n1011 & ~n8222;
  assign n8224 = n1015 & ~n8223;
  assign n8225 = n1019 & ~n8224;
  assign n8226 = n1023 & ~n8225;
  assign n8227 = n1027 & ~n8226;
  assign n8228 = n1031 & ~n8227;
  assign n8229 = n1035 & ~n8228;
  assign n8230 = n1039 & ~n8229;
  assign n8231 = n1043 & ~n8230;
  assign n8232 = n1047 & ~n8231;
  assign n8233 = n1051 & ~n8232;
  assign n8234 = n1055 & ~n8233;
  assign n8235 = n1059 & ~n8234;
  assign n8236 = n1574 & ~n8235;
  assign n8237 = n1576 & ~n8236;
  assign n8238 = n1837 & ~n8237;
  assign n8239 = n1068 & ~n8238;
  assign n8240 = n1072 & ~n8239;
  assign n8241 = n1076 & ~n8240;
  assign n8242 = n1080 & ~n8241;
  assign n8243 = n1084 & ~n8242;
  assign n8244 = n1088 & ~n8243;
  assign n8245 = n1092 & ~n8244;
  assign n8246 = n1096 & ~n8245;
  assign n8247 = n1100 & ~n8246;
  assign n8248 = n1104 & ~n8247;
  assign n8249 = n1108 & ~n8248;
  assign n8250 = n1112 & ~n8249;
  assign n8251 = n1116 & ~n8250;
  assign n8252 = n1120 & ~n8251;
  assign n8253 = n1124 & ~n8252;
  assign n8254 = n1128 & ~n8253;
  assign n8255 = n1132 & ~n8254;
  assign n8256 = n1136 & ~n8255;
  assign n8257 = n1140 & ~n8256;
  assign n8258 = n1144 & ~n8257;
  assign n8259 = n1148 & ~n8258;
  assign n8260 = n1152 & ~n8259;
  assign n8261 = n1156 & ~n8260;
  assign n8262 = n1160 & ~n8261;
  assign n8263 = n1164 & ~n8262;
  assign n8264 = n1168 & ~n8263;
  assign n8265 = n1172 & ~n8264;
  assign n8266 = n1176 & ~n8265;
  assign n8267 = n1180 & ~n8266;
  assign n8268 = n1184 & ~n8267;
  assign n8269 = n1188 & ~n8268;
  assign n8270 = n1192 & ~n8269;
  assign n8271 = n1196 & ~n8270;
  assign n8272 = n1200 & ~n8271;
  assign n8273 = n1204 & ~n8272;
  assign n8274 = n1208 & ~n8273;
  assign n8275 = n1212 & ~n8274;
  assign n8276 = n1216 & ~n8275;
  assign n8277 = n1220 & ~n8276;
  assign n8278 = n1224 & ~n8277;
  assign n8279 = n1228 & ~n8278;
  assign n8280 = n1232 & ~n8279;
  assign n8281 = n1236 & ~n8280;
  assign n8282 = n1240 & ~n8281;
  assign n8283 = n1244 & ~n8282;
  assign n8284 = n1248 & ~n8283;
  assign n8285 = n1252 & ~n8284;
  assign n8286 = n1256 & ~n8285;
  assign n8287 = n1260 & ~n8286;
  assign n8288 = n1264 & ~n8287;
  assign n8289 = n1268 & ~n8288;
  assign n8290 = pi210  & ~n1270;
  assign po82  = ~n8289 & n8290;
  assign n8292 = ~n607 & n1279;
  assign n8293 = n1284 & ~n8292;
  assign n8294 = n1288 & ~n8293;
  assign n8295 = n1292 & ~n8294;
  assign n8296 = n1296 & ~n8295;
  assign n8297 = n1300 & ~n8296;
  assign n8298 = n1304 & ~n8297;
  assign n8299 = n1308 & ~n8298;
  assign n8300 = n1312 & ~n8299;
  assign n8301 = n1316 & ~n8300;
  assign n8302 = n1320 & ~n8301;
  assign n8303 = n1324 & ~n8302;
  assign n8304 = n1328 & ~n8303;
  assign n8305 = n1332 & ~n8304;
  assign n8306 = n1336 & ~n8305;
  assign n8307 = n1340 & ~n8306;
  assign n8308 = n1344 & ~n8307;
  assign n8309 = n1348 & ~n8308;
  assign n8310 = n1352 & ~n8309;
  assign n8311 = n1356 & ~n8310;
  assign n8312 = n1360 & ~n8311;
  assign n8313 = n1364 & ~n8312;
  assign n8314 = n1368 & ~n8313;
  assign n8315 = n1372 & ~n8314;
  assign n8316 = n1376 & ~n8315;
  assign n8317 = n1380 & ~n8316;
  assign n8318 = n1384 & ~n8317;
  assign n8319 = n1388 & ~n8318;
  assign n8320 = n1392 & ~n8319;
  assign n8321 = n1396 & ~n8320;
  assign n8322 = n1663 & ~n8321;
  assign n8323 = n392 & ~n8322;
  assign n8324 = n396 & ~n8323;
  assign n8325 = n400 & ~n8324;
  assign n8326 = n404 & ~n8325;
  assign n8327 = n408 & ~n8326;
  assign n8328 = n412 & ~n8327;
  assign n8329 = n416 & ~n8328;
  assign n8330 = n420 & ~n8329;
  assign n8331 = n424 & ~n8330;
  assign n8332 = n428 & ~n8331;
  assign n8333 = n432 & ~n8332;
  assign n8334 = n436 & ~n8333;
  assign n8335 = n440 & ~n8334;
  assign n8336 = n444 & ~n8335;
  assign n8337 = n448 & ~n8336;
  assign n8338 = n452 & ~n8337;
  assign n8339 = n456 & ~n8338;
  assign n8340 = n460 & ~n8339;
  assign n8341 = n464 & ~n8340;
  assign n8342 = n468 & ~n8341;
  assign n8343 = n472 & ~n8342;
  assign n8344 = n476 & ~n8343;
  assign n8345 = n480 & ~n8344;
  assign n8346 = n484 & ~n8345;
  assign n8347 = n488 & ~n8346;
  assign n8348 = n492 & ~n8347;
  assign n8349 = n496 & ~n8348;
  assign n8350 = n500 & ~n8349;
  assign n8351 = n504 & ~n8350;
  assign n8352 = n508 & ~n8351;
  assign n8353 = n512 & ~n8352;
  assign n8354 = n516 & ~n8353;
  assign n8355 = n520 & ~n8354;
  assign n8356 = n524 & ~n8355;
  assign n8357 = n528 & ~n8356;
  assign n8358 = n532 & ~n8357;
  assign n8359 = n536 & ~n8358;
  assign n8360 = n540 & ~n8359;
  assign n8361 = n544 & ~n8360;
  assign n8362 = n548 & ~n8361;
  assign n8363 = n552 & ~n8362;
  assign n8364 = n556 & ~n8363;
  assign n8365 = n560 & ~n8364;
  assign n8366 = n564 & ~n8365;
  assign n8367 = n568 & ~n8366;
  assign n8368 = n572 & ~n8367;
  assign n8369 = n576 & ~n8368;
  assign n8370 = n580 & ~n8369;
  assign n8371 = n584 & ~n8370;
  assign n8372 = n588 & ~n8371;
  assign n8373 = n592 & ~n8372;
  assign n8374 = n596 & ~n8373;
  assign n8375 = n600 & ~n8374;
  assign n8376 = pi211  & ~n602;
  assign po83  = ~n8375 & n8376;
  assign n8378 = n611 & ~n946;
  assign n8379 = n616 & ~n8378;
  assign n8380 = n620 & ~n8379;
  assign n8381 = n624 & ~n8380;
  assign n8382 = n628 & ~n8381;
  assign n8383 = n632 & ~n8382;
  assign n8384 = n636 & ~n8383;
  assign n8385 = n640 & ~n8384;
  assign n8386 = n644 & ~n8385;
  assign n8387 = n648 & ~n8386;
  assign n8388 = n652 & ~n8387;
  assign n8389 = n656 & ~n8388;
  assign n8390 = n660 & ~n8389;
  assign n8391 = n664 & ~n8390;
  assign n8392 = n668 & ~n8391;
  assign n8393 = n672 & ~n8392;
  assign n8394 = n676 & ~n8393;
  assign n8395 = n680 & ~n8394;
  assign n8396 = n684 & ~n8395;
  assign n8397 = n688 & ~n8396;
  assign n8398 = n692 & ~n8397;
  assign n8399 = n696 & ~n8398;
  assign n8400 = n700 & ~n8399;
  assign n8401 = n704 & ~n8400;
  assign n8402 = n708 & ~n8401;
  assign n8403 = n712 & ~n8402;
  assign n8404 = n716 & ~n8403;
  assign n8405 = n720 & ~n8404;
  assign n8406 = n1484 & ~n8405;
  assign n8407 = n1486 & ~n8406;
  assign n8408 = n1750 & ~n8407;
  assign n8409 = n731 & ~n8408;
  assign n8410 = n735 & ~n8409;
  assign n8411 = n739 & ~n8410;
  assign n8412 = n743 & ~n8411;
  assign n8413 = n747 & ~n8412;
  assign n8414 = n751 & ~n8413;
  assign n8415 = n755 & ~n8414;
  assign n8416 = n759 & ~n8415;
  assign n8417 = n763 & ~n8416;
  assign n8418 = n767 & ~n8417;
  assign n8419 = n771 & ~n8418;
  assign n8420 = n775 & ~n8419;
  assign n8421 = n779 & ~n8420;
  assign n8422 = n783 & ~n8421;
  assign n8423 = n787 & ~n8422;
  assign n8424 = n791 & ~n8423;
  assign n8425 = n795 & ~n8424;
  assign n8426 = n799 & ~n8425;
  assign n8427 = n803 & ~n8426;
  assign n8428 = n807 & ~n8427;
  assign n8429 = n811 & ~n8428;
  assign n8430 = n815 & ~n8429;
  assign n8431 = n819 & ~n8430;
  assign n8432 = n823 & ~n8431;
  assign n8433 = n827 & ~n8432;
  assign n8434 = n831 & ~n8433;
  assign n8435 = n835 & ~n8434;
  assign n8436 = n839 & ~n8435;
  assign n8437 = n843 & ~n8436;
  assign n8438 = n847 & ~n8437;
  assign n8439 = n851 & ~n8438;
  assign n8440 = n855 & ~n8439;
  assign n8441 = n859 & ~n8440;
  assign n8442 = n863 & ~n8441;
  assign n8443 = n867 & ~n8442;
  assign n8444 = n871 & ~n8443;
  assign n8445 = n875 & ~n8444;
  assign n8446 = n879 & ~n8445;
  assign n8447 = n883 & ~n8446;
  assign n8448 = n887 & ~n8447;
  assign n8449 = n891 & ~n8448;
  assign n8450 = n895 & ~n8449;
  assign n8451 = n899 & ~n8450;
  assign n8452 = n903 & ~n8451;
  assign n8453 = n907 & ~n8452;
  assign n8454 = n911 & ~n8453;
  assign n8455 = n915 & ~n8454;
  assign n8456 = n919 & ~n8455;
  assign n8457 = n923 & ~n8456;
  assign n8458 = n927 & ~n8457;
  assign n8459 = n931 & ~n8458;
  assign n8460 = n935 & ~n8459;
  assign n8461 = n939 & ~n8460;
  assign n8462 = pi212  & ~n941;
  assign po84  = ~n8461 & n8462;
  assign n8464 = n950 & ~n1283;
  assign n8465 = n955 & ~n8464;
  assign n8466 = n959 & ~n8465;
  assign n8467 = n963 & ~n8466;
  assign n8468 = n967 & ~n8467;
  assign n8469 = n971 & ~n8468;
  assign n8470 = n975 & ~n8469;
  assign n8471 = n979 & ~n8470;
  assign n8472 = n983 & ~n8471;
  assign n8473 = n987 & ~n8472;
  assign n8474 = n991 & ~n8473;
  assign n8475 = n995 & ~n8474;
  assign n8476 = n999 & ~n8475;
  assign n8477 = n1003 & ~n8476;
  assign n8478 = n1007 & ~n8477;
  assign n8479 = n1011 & ~n8478;
  assign n8480 = n1015 & ~n8479;
  assign n8481 = n1019 & ~n8480;
  assign n8482 = n1023 & ~n8481;
  assign n8483 = n1027 & ~n8482;
  assign n8484 = n1031 & ~n8483;
  assign n8485 = n1035 & ~n8484;
  assign n8486 = n1039 & ~n8485;
  assign n8487 = n1043 & ~n8486;
  assign n8488 = n1047 & ~n8487;
  assign n8489 = n1051 & ~n8488;
  assign n8490 = n1055 & ~n8489;
  assign n8491 = n1059 & ~n8490;
  assign n8492 = n1574 & ~n8491;
  assign n8493 = n1576 & ~n8492;
  assign n8494 = n1837 & ~n8493;
  assign n8495 = n1068 & ~n8494;
  assign n8496 = n1072 & ~n8495;
  assign n8497 = n1076 & ~n8496;
  assign n8498 = n1080 & ~n8497;
  assign n8499 = n1084 & ~n8498;
  assign n8500 = n1088 & ~n8499;
  assign n8501 = n1092 & ~n8500;
  assign n8502 = n1096 & ~n8501;
  assign n8503 = n1100 & ~n8502;
  assign n8504 = n1104 & ~n8503;
  assign n8505 = n1108 & ~n8504;
  assign n8506 = n1112 & ~n8505;
  assign n8507 = n1116 & ~n8506;
  assign n8508 = n1120 & ~n8507;
  assign n8509 = n1124 & ~n8508;
  assign n8510 = n1128 & ~n8509;
  assign n8511 = n1132 & ~n8510;
  assign n8512 = n1136 & ~n8511;
  assign n8513 = n1140 & ~n8512;
  assign n8514 = n1144 & ~n8513;
  assign n8515 = n1148 & ~n8514;
  assign n8516 = n1152 & ~n8515;
  assign n8517 = n1156 & ~n8516;
  assign n8518 = n1160 & ~n8517;
  assign n8519 = n1164 & ~n8518;
  assign n8520 = n1168 & ~n8519;
  assign n8521 = n1172 & ~n8520;
  assign n8522 = n1176 & ~n8521;
  assign n8523 = n1180 & ~n8522;
  assign n8524 = n1184 & ~n8523;
  assign n8525 = n1188 & ~n8524;
  assign n8526 = n1192 & ~n8525;
  assign n8527 = n1196 & ~n8526;
  assign n8528 = n1200 & ~n8527;
  assign n8529 = n1204 & ~n8528;
  assign n8530 = n1208 & ~n8529;
  assign n8531 = n1212 & ~n8530;
  assign n8532 = n1216 & ~n8531;
  assign n8533 = n1220 & ~n8532;
  assign n8534 = n1224 & ~n8533;
  assign n8535 = n1228 & ~n8534;
  assign n8536 = n1232 & ~n8535;
  assign n8537 = n1236 & ~n8536;
  assign n8538 = n1240 & ~n8537;
  assign n8539 = n1244 & ~n8538;
  assign n8540 = n1248 & ~n8539;
  assign n8541 = n1252 & ~n8540;
  assign n8542 = n1256 & ~n8541;
  assign n8543 = n1260 & ~n8542;
  assign n8544 = n1264 & ~n8543;
  assign n8545 = n1268 & ~n8544;
  assign n8546 = n1272 & ~n8545;
  assign n8547 = n1276 & ~n8546;
  assign n8548 = pi213  & ~n1278;
  assign po85  = ~n8547 & n8548;
  assign n8550 = ~n615 & n1287;
  assign n8551 = n1292 & ~n8550;
  assign n8552 = n1296 & ~n8551;
  assign n8553 = n1300 & ~n8552;
  assign n8554 = n1304 & ~n8553;
  assign n8555 = n1308 & ~n8554;
  assign n8556 = n1312 & ~n8555;
  assign n8557 = n1316 & ~n8556;
  assign n8558 = n1320 & ~n8557;
  assign n8559 = n1324 & ~n8558;
  assign n8560 = n1328 & ~n8559;
  assign n8561 = n1332 & ~n8560;
  assign n8562 = n1336 & ~n8561;
  assign n8563 = n1340 & ~n8562;
  assign n8564 = n1344 & ~n8563;
  assign n8565 = n1348 & ~n8564;
  assign n8566 = n1352 & ~n8565;
  assign n8567 = n1356 & ~n8566;
  assign n8568 = n1360 & ~n8567;
  assign n8569 = n1364 & ~n8568;
  assign n8570 = n1368 & ~n8569;
  assign n8571 = n1372 & ~n8570;
  assign n8572 = n1376 & ~n8571;
  assign n8573 = n1380 & ~n8572;
  assign n8574 = n1384 & ~n8573;
  assign n8575 = n1388 & ~n8574;
  assign n8576 = n1392 & ~n8575;
  assign n8577 = n1396 & ~n8576;
  assign n8578 = n1663 & ~n8577;
  assign n8579 = n392 & ~n8578;
  assign n8580 = n396 & ~n8579;
  assign n8581 = n400 & ~n8580;
  assign n8582 = n404 & ~n8581;
  assign n8583 = n408 & ~n8582;
  assign n8584 = n412 & ~n8583;
  assign n8585 = n416 & ~n8584;
  assign n8586 = n420 & ~n8585;
  assign n8587 = n424 & ~n8586;
  assign n8588 = n428 & ~n8587;
  assign n8589 = n432 & ~n8588;
  assign n8590 = n436 & ~n8589;
  assign n8591 = n440 & ~n8590;
  assign n8592 = n444 & ~n8591;
  assign n8593 = n448 & ~n8592;
  assign n8594 = n452 & ~n8593;
  assign n8595 = n456 & ~n8594;
  assign n8596 = n460 & ~n8595;
  assign n8597 = n464 & ~n8596;
  assign n8598 = n468 & ~n8597;
  assign n8599 = n472 & ~n8598;
  assign n8600 = n476 & ~n8599;
  assign n8601 = n480 & ~n8600;
  assign n8602 = n484 & ~n8601;
  assign n8603 = n488 & ~n8602;
  assign n8604 = n492 & ~n8603;
  assign n8605 = n496 & ~n8604;
  assign n8606 = n500 & ~n8605;
  assign n8607 = n504 & ~n8606;
  assign n8608 = n508 & ~n8607;
  assign n8609 = n512 & ~n8608;
  assign n8610 = n516 & ~n8609;
  assign n8611 = n520 & ~n8610;
  assign n8612 = n524 & ~n8611;
  assign n8613 = n528 & ~n8612;
  assign n8614 = n532 & ~n8613;
  assign n8615 = n536 & ~n8614;
  assign n8616 = n540 & ~n8615;
  assign n8617 = n544 & ~n8616;
  assign n8618 = n548 & ~n8617;
  assign n8619 = n552 & ~n8618;
  assign n8620 = n556 & ~n8619;
  assign n8621 = n560 & ~n8620;
  assign n8622 = n564 & ~n8621;
  assign n8623 = n568 & ~n8622;
  assign n8624 = n572 & ~n8623;
  assign n8625 = n576 & ~n8624;
  assign n8626 = n580 & ~n8625;
  assign n8627 = n584 & ~n8626;
  assign n8628 = n588 & ~n8627;
  assign n8629 = n592 & ~n8628;
  assign n8630 = n596 & ~n8629;
  assign n8631 = n600 & ~n8630;
  assign n8632 = n604 & ~n8631;
  assign n8633 = n608 & ~n8632;
  assign n8634 = pi214  & ~n610;
  assign po86  = ~n8633 & n8634;
  assign n8636 = n619 & ~n954;
  assign n8637 = n624 & ~n8636;
  assign n8638 = n628 & ~n8637;
  assign n8639 = n632 & ~n8638;
  assign n8640 = n636 & ~n8639;
  assign n8641 = n640 & ~n8640;
  assign n8642 = n644 & ~n8641;
  assign n8643 = n648 & ~n8642;
  assign n8644 = n652 & ~n8643;
  assign n8645 = n656 & ~n8644;
  assign n8646 = n660 & ~n8645;
  assign n8647 = n664 & ~n8646;
  assign n8648 = n668 & ~n8647;
  assign n8649 = n672 & ~n8648;
  assign n8650 = n676 & ~n8649;
  assign n8651 = n680 & ~n8650;
  assign n8652 = n684 & ~n8651;
  assign n8653 = n688 & ~n8652;
  assign n8654 = n692 & ~n8653;
  assign n8655 = n696 & ~n8654;
  assign n8656 = n700 & ~n8655;
  assign n8657 = n704 & ~n8656;
  assign n8658 = n708 & ~n8657;
  assign n8659 = n712 & ~n8658;
  assign n8660 = n716 & ~n8659;
  assign n8661 = n720 & ~n8660;
  assign n8662 = n1484 & ~n8661;
  assign n8663 = n1486 & ~n8662;
  assign n8664 = n1750 & ~n8663;
  assign n8665 = n731 & ~n8664;
  assign n8666 = n735 & ~n8665;
  assign n8667 = n739 & ~n8666;
  assign n8668 = n743 & ~n8667;
  assign n8669 = n747 & ~n8668;
  assign n8670 = n751 & ~n8669;
  assign n8671 = n755 & ~n8670;
  assign n8672 = n759 & ~n8671;
  assign n8673 = n763 & ~n8672;
  assign n8674 = n767 & ~n8673;
  assign n8675 = n771 & ~n8674;
  assign n8676 = n775 & ~n8675;
  assign n8677 = n779 & ~n8676;
  assign n8678 = n783 & ~n8677;
  assign n8679 = n787 & ~n8678;
  assign n8680 = n791 & ~n8679;
  assign n8681 = n795 & ~n8680;
  assign n8682 = n799 & ~n8681;
  assign n8683 = n803 & ~n8682;
  assign n8684 = n807 & ~n8683;
  assign n8685 = n811 & ~n8684;
  assign n8686 = n815 & ~n8685;
  assign n8687 = n819 & ~n8686;
  assign n8688 = n823 & ~n8687;
  assign n8689 = n827 & ~n8688;
  assign n8690 = n831 & ~n8689;
  assign n8691 = n835 & ~n8690;
  assign n8692 = n839 & ~n8691;
  assign n8693 = n843 & ~n8692;
  assign n8694 = n847 & ~n8693;
  assign n8695 = n851 & ~n8694;
  assign n8696 = n855 & ~n8695;
  assign n8697 = n859 & ~n8696;
  assign n8698 = n863 & ~n8697;
  assign n8699 = n867 & ~n8698;
  assign n8700 = n871 & ~n8699;
  assign n8701 = n875 & ~n8700;
  assign n8702 = n879 & ~n8701;
  assign n8703 = n883 & ~n8702;
  assign n8704 = n887 & ~n8703;
  assign n8705 = n891 & ~n8704;
  assign n8706 = n895 & ~n8705;
  assign n8707 = n899 & ~n8706;
  assign n8708 = n903 & ~n8707;
  assign n8709 = n907 & ~n8708;
  assign n8710 = n911 & ~n8709;
  assign n8711 = n915 & ~n8710;
  assign n8712 = n919 & ~n8711;
  assign n8713 = n923 & ~n8712;
  assign n8714 = n927 & ~n8713;
  assign n8715 = n931 & ~n8714;
  assign n8716 = n935 & ~n8715;
  assign n8717 = n939 & ~n8716;
  assign n8718 = n943 & ~n8717;
  assign n8719 = n947 & ~n8718;
  assign n8720 = pi215  & ~n949;
  assign po87  = ~n8719 & n8720;
  assign n8722 = n958 & ~n1291;
  assign n8723 = n963 & ~n8722;
  assign n8724 = n967 & ~n8723;
  assign n8725 = n971 & ~n8724;
  assign n8726 = n975 & ~n8725;
  assign n8727 = n979 & ~n8726;
  assign n8728 = n983 & ~n8727;
  assign n8729 = n987 & ~n8728;
  assign n8730 = n991 & ~n8729;
  assign n8731 = n995 & ~n8730;
  assign n8732 = n999 & ~n8731;
  assign n8733 = n1003 & ~n8732;
  assign n8734 = n1007 & ~n8733;
  assign n8735 = n1011 & ~n8734;
  assign n8736 = n1015 & ~n8735;
  assign n8737 = n1019 & ~n8736;
  assign n8738 = n1023 & ~n8737;
  assign n8739 = n1027 & ~n8738;
  assign n8740 = n1031 & ~n8739;
  assign n8741 = n1035 & ~n8740;
  assign n8742 = n1039 & ~n8741;
  assign n8743 = n1043 & ~n8742;
  assign n8744 = n1047 & ~n8743;
  assign n8745 = n1051 & ~n8744;
  assign n8746 = n1055 & ~n8745;
  assign n8747 = n1059 & ~n8746;
  assign n8748 = n1574 & ~n8747;
  assign n8749 = n1576 & ~n8748;
  assign n8750 = n1837 & ~n8749;
  assign n8751 = n1068 & ~n8750;
  assign n8752 = n1072 & ~n8751;
  assign n8753 = n1076 & ~n8752;
  assign n8754 = n1080 & ~n8753;
  assign n8755 = n1084 & ~n8754;
  assign n8756 = n1088 & ~n8755;
  assign n8757 = n1092 & ~n8756;
  assign n8758 = n1096 & ~n8757;
  assign n8759 = n1100 & ~n8758;
  assign n8760 = n1104 & ~n8759;
  assign n8761 = n1108 & ~n8760;
  assign n8762 = n1112 & ~n8761;
  assign n8763 = n1116 & ~n8762;
  assign n8764 = n1120 & ~n8763;
  assign n8765 = n1124 & ~n8764;
  assign n8766 = n1128 & ~n8765;
  assign n8767 = n1132 & ~n8766;
  assign n8768 = n1136 & ~n8767;
  assign n8769 = n1140 & ~n8768;
  assign n8770 = n1144 & ~n8769;
  assign n8771 = n1148 & ~n8770;
  assign n8772 = n1152 & ~n8771;
  assign n8773 = n1156 & ~n8772;
  assign n8774 = n1160 & ~n8773;
  assign n8775 = n1164 & ~n8774;
  assign n8776 = n1168 & ~n8775;
  assign n8777 = n1172 & ~n8776;
  assign n8778 = n1176 & ~n8777;
  assign n8779 = n1180 & ~n8778;
  assign n8780 = n1184 & ~n8779;
  assign n8781 = n1188 & ~n8780;
  assign n8782 = n1192 & ~n8781;
  assign n8783 = n1196 & ~n8782;
  assign n8784 = n1200 & ~n8783;
  assign n8785 = n1204 & ~n8784;
  assign n8786 = n1208 & ~n8785;
  assign n8787 = n1212 & ~n8786;
  assign n8788 = n1216 & ~n8787;
  assign n8789 = n1220 & ~n8788;
  assign n8790 = n1224 & ~n8789;
  assign n8791 = n1228 & ~n8790;
  assign n8792 = n1232 & ~n8791;
  assign n8793 = n1236 & ~n8792;
  assign n8794 = n1240 & ~n8793;
  assign n8795 = n1244 & ~n8794;
  assign n8796 = n1248 & ~n8795;
  assign n8797 = n1252 & ~n8796;
  assign n8798 = n1256 & ~n8797;
  assign n8799 = n1260 & ~n8798;
  assign n8800 = n1264 & ~n8799;
  assign n8801 = n1268 & ~n8800;
  assign n8802 = n1272 & ~n8801;
  assign n8803 = n1276 & ~n8802;
  assign n8804 = n1280 & ~n8803;
  assign n8805 = n1284 & ~n8804;
  assign n8806 = pi216  & ~n1286;
  assign po88  = ~n8805 & n8806;
  assign n8808 = ~n623 & n1295;
  assign n8809 = n1300 & ~n8808;
  assign n8810 = n1304 & ~n8809;
  assign n8811 = n1308 & ~n8810;
  assign n8812 = n1312 & ~n8811;
  assign n8813 = n1316 & ~n8812;
  assign n8814 = n1320 & ~n8813;
  assign n8815 = n1324 & ~n8814;
  assign n8816 = n1328 & ~n8815;
  assign n8817 = n1332 & ~n8816;
  assign n8818 = n1336 & ~n8817;
  assign n8819 = n1340 & ~n8818;
  assign n8820 = n1344 & ~n8819;
  assign n8821 = n1348 & ~n8820;
  assign n8822 = n1352 & ~n8821;
  assign n8823 = n1356 & ~n8822;
  assign n8824 = n1360 & ~n8823;
  assign n8825 = n1364 & ~n8824;
  assign n8826 = n1368 & ~n8825;
  assign n8827 = n1372 & ~n8826;
  assign n8828 = n1376 & ~n8827;
  assign n8829 = n1380 & ~n8828;
  assign n8830 = n1384 & ~n8829;
  assign n8831 = n1388 & ~n8830;
  assign n8832 = n1392 & ~n8831;
  assign n8833 = n1396 & ~n8832;
  assign n8834 = n1663 & ~n8833;
  assign n8835 = n392 & ~n8834;
  assign n8836 = n396 & ~n8835;
  assign n8837 = n400 & ~n8836;
  assign n8838 = n404 & ~n8837;
  assign n8839 = n408 & ~n8838;
  assign n8840 = n412 & ~n8839;
  assign n8841 = n416 & ~n8840;
  assign n8842 = n420 & ~n8841;
  assign n8843 = n424 & ~n8842;
  assign n8844 = n428 & ~n8843;
  assign n8845 = n432 & ~n8844;
  assign n8846 = n436 & ~n8845;
  assign n8847 = n440 & ~n8846;
  assign n8848 = n444 & ~n8847;
  assign n8849 = n448 & ~n8848;
  assign n8850 = n452 & ~n8849;
  assign n8851 = n456 & ~n8850;
  assign n8852 = n460 & ~n8851;
  assign n8853 = n464 & ~n8852;
  assign n8854 = n468 & ~n8853;
  assign n8855 = n472 & ~n8854;
  assign n8856 = n476 & ~n8855;
  assign n8857 = n480 & ~n8856;
  assign n8858 = n484 & ~n8857;
  assign n8859 = n488 & ~n8858;
  assign n8860 = n492 & ~n8859;
  assign n8861 = n496 & ~n8860;
  assign n8862 = n500 & ~n8861;
  assign n8863 = n504 & ~n8862;
  assign n8864 = n508 & ~n8863;
  assign n8865 = n512 & ~n8864;
  assign n8866 = n516 & ~n8865;
  assign n8867 = n520 & ~n8866;
  assign n8868 = n524 & ~n8867;
  assign n8869 = n528 & ~n8868;
  assign n8870 = n532 & ~n8869;
  assign n8871 = n536 & ~n8870;
  assign n8872 = n540 & ~n8871;
  assign n8873 = n544 & ~n8872;
  assign n8874 = n548 & ~n8873;
  assign n8875 = n552 & ~n8874;
  assign n8876 = n556 & ~n8875;
  assign n8877 = n560 & ~n8876;
  assign n8878 = n564 & ~n8877;
  assign n8879 = n568 & ~n8878;
  assign n8880 = n572 & ~n8879;
  assign n8881 = n576 & ~n8880;
  assign n8882 = n580 & ~n8881;
  assign n8883 = n584 & ~n8882;
  assign n8884 = n588 & ~n8883;
  assign n8885 = n592 & ~n8884;
  assign n8886 = n596 & ~n8885;
  assign n8887 = n600 & ~n8886;
  assign n8888 = n604 & ~n8887;
  assign n8889 = n608 & ~n8888;
  assign n8890 = n612 & ~n8889;
  assign n8891 = n616 & ~n8890;
  assign n8892 = pi217  & ~n618;
  assign po89  = ~n8891 & n8892;
  assign n8894 = n627 & ~n962;
  assign n8895 = n632 & ~n8894;
  assign n8896 = n636 & ~n8895;
  assign n8897 = n640 & ~n8896;
  assign n8898 = n644 & ~n8897;
  assign n8899 = n648 & ~n8898;
  assign n8900 = n652 & ~n8899;
  assign n8901 = n656 & ~n8900;
  assign n8902 = n660 & ~n8901;
  assign n8903 = n664 & ~n8902;
  assign n8904 = n668 & ~n8903;
  assign n8905 = n672 & ~n8904;
  assign n8906 = n676 & ~n8905;
  assign n8907 = n680 & ~n8906;
  assign n8908 = n684 & ~n8907;
  assign n8909 = n688 & ~n8908;
  assign n8910 = n692 & ~n8909;
  assign n8911 = n696 & ~n8910;
  assign n8912 = n700 & ~n8911;
  assign n8913 = n704 & ~n8912;
  assign n8914 = n708 & ~n8913;
  assign n8915 = n712 & ~n8914;
  assign n8916 = n716 & ~n8915;
  assign n8917 = n720 & ~n8916;
  assign n8918 = n1484 & ~n8917;
  assign n8919 = n1486 & ~n8918;
  assign n8920 = n1750 & ~n8919;
  assign n8921 = n731 & ~n8920;
  assign n8922 = n735 & ~n8921;
  assign n8923 = n739 & ~n8922;
  assign n8924 = n743 & ~n8923;
  assign n8925 = n747 & ~n8924;
  assign n8926 = n751 & ~n8925;
  assign n8927 = n755 & ~n8926;
  assign n8928 = n759 & ~n8927;
  assign n8929 = n763 & ~n8928;
  assign n8930 = n767 & ~n8929;
  assign n8931 = n771 & ~n8930;
  assign n8932 = n775 & ~n8931;
  assign n8933 = n779 & ~n8932;
  assign n8934 = n783 & ~n8933;
  assign n8935 = n787 & ~n8934;
  assign n8936 = n791 & ~n8935;
  assign n8937 = n795 & ~n8936;
  assign n8938 = n799 & ~n8937;
  assign n8939 = n803 & ~n8938;
  assign n8940 = n807 & ~n8939;
  assign n8941 = n811 & ~n8940;
  assign n8942 = n815 & ~n8941;
  assign n8943 = n819 & ~n8942;
  assign n8944 = n823 & ~n8943;
  assign n8945 = n827 & ~n8944;
  assign n8946 = n831 & ~n8945;
  assign n8947 = n835 & ~n8946;
  assign n8948 = n839 & ~n8947;
  assign n8949 = n843 & ~n8948;
  assign n8950 = n847 & ~n8949;
  assign n8951 = n851 & ~n8950;
  assign n8952 = n855 & ~n8951;
  assign n8953 = n859 & ~n8952;
  assign n8954 = n863 & ~n8953;
  assign n8955 = n867 & ~n8954;
  assign n8956 = n871 & ~n8955;
  assign n8957 = n875 & ~n8956;
  assign n8958 = n879 & ~n8957;
  assign n8959 = n883 & ~n8958;
  assign n8960 = n887 & ~n8959;
  assign n8961 = n891 & ~n8960;
  assign n8962 = n895 & ~n8961;
  assign n8963 = n899 & ~n8962;
  assign n8964 = n903 & ~n8963;
  assign n8965 = n907 & ~n8964;
  assign n8966 = n911 & ~n8965;
  assign n8967 = n915 & ~n8966;
  assign n8968 = n919 & ~n8967;
  assign n8969 = n923 & ~n8968;
  assign n8970 = n927 & ~n8969;
  assign n8971 = n931 & ~n8970;
  assign n8972 = n935 & ~n8971;
  assign n8973 = n939 & ~n8972;
  assign n8974 = n943 & ~n8973;
  assign n8975 = n947 & ~n8974;
  assign n8976 = n951 & ~n8975;
  assign n8977 = n955 & ~n8976;
  assign n8978 = pi218  & ~n957;
  assign po90  = ~n8977 & n8978;
  assign n8980 = n966 & ~n1299;
  assign n8981 = n971 & ~n8980;
  assign n8982 = n975 & ~n8981;
  assign n8983 = n979 & ~n8982;
  assign n8984 = n983 & ~n8983;
  assign n8985 = n987 & ~n8984;
  assign n8986 = n991 & ~n8985;
  assign n8987 = n995 & ~n8986;
  assign n8988 = n999 & ~n8987;
  assign n8989 = n1003 & ~n8988;
  assign n8990 = n1007 & ~n8989;
  assign n8991 = n1011 & ~n8990;
  assign n8992 = n1015 & ~n8991;
  assign n8993 = n1019 & ~n8992;
  assign n8994 = n1023 & ~n8993;
  assign n8995 = n1027 & ~n8994;
  assign n8996 = n1031 & ~n8995;
  assign n8997 = n1035 & ~n8996;
  assign n8998 = n1039 & ~n8997;
  assign n8999 = n1043 & ~n8998;
  assign n9000 = n1047 & ~n8999;
  assign n9001 = n1051 & ~n9000;
  assign n9002 = n1055 & ~n9001;
  assign n9003 = n1059 & ~n9002;
  assign n9004 = n1574 & ~n9003;
  assign n9005 = n1576 & ~n9004;
  assign n9006 = n1837 & ~n9005;
  assign n9007 = n1068 & ~n9006;
  assign n9008 = n1072 & ~n9007;
  assign n9009 = n1076 & ~n9008;
  assign n9010 = n1080 & ~n9009;
  assign n9011 = n1084 & ~n9010;
  assign n9012 = n1088 & ~n9011;
  assign n9013 = n1092 & ~n9012;
  assign n9014 = n1096 & ~n9013;
  assign n9015 = n1100 & ~n9014;
  assign n9016 = n1104 & ~n9015;
  assign n9017 = n1108 & ~n9016;
  assign n9018 = n1112 & ~n9017;
  assign n9019 = n1116 & ~n9018;
  assign n9020 = n1120 & ~n9019;
  assign n9021 = n1124 & ~n9020;
  assign n9022 = n1128 & ~n9021;
  assign n9023 = n1132 & ~n9022;
  assign n9024 = n1136 & ~n9023;
  assign n9025 = n1140 & ~n9024;
  assign n9026 = n1144 & ~n9025;
  assign n9027 = n1148 & ~n9026;
  assign n9028 = n1152 & ~n9027;
  assign n9029 = n1156 & ~n9028;
  assign n9030 = n1160 & ~n9029;
  assign n9031 = n1164 & ~n9030;
  assign n9032 = n1168 & ~n9031;
  assign n9033 = n1172 & ~n9032;
  assign n9034 = n1176 & ~n9033;
  assign n9035 = n1180 & ~n9034;
  assign n9036 = n1184 & ~n9035;
  assign n9037 = n1188 & ~n9036;
  assign n9038 = n1192 & ~n9037;
  assign n9039 = n1196 & ~n9038;
  assign n9040 = n1200 & ~n9039;
  assign n9041 = n1204 & ~n9040;
  assign n9042 = n1208 & ~n9041;
  assign n9043 = n1212 & ~n9042;
  assign n9044 = n1216 & ~n9043;
  assign n9045 = n1220 & ~n9044;
  assign n9046 = n1224 & ~n9045;
  assign n9047 = n1228 & ~n9046;
  assign n9048 = n1232 & ~n9047;
  assign n9049 = n1236 & ~n9048;
  assign n9050 = n1240 & ~n9049;
  assign n9051 = n1244 & ~n9050;
  assign n9052 = n1248 & ~n9051;
  assign n9053 = n1252 & ~n9052;
  assign n9054 = n1256 & ~n9053;
  assign n9055 = n1260 & ~n9054;
  assign n9056 = n1264 & ~n9055;
  assign n9057 = n1268 & ~n9056;
  assign n9058 = n1272 & ~n9057;
  assign n9059 = n1276 & ~n9058;
  assign n9060 = n1280 & ~n9059;
  assign n9061 = n1284 & ~n9060;
  assign n9062 = n1288 & ~n9061;
  assign n9063 = n1292 & ~n9062;
  assign n9064 = pi219  & ~n1294;
  assign po91  = ~n9063 & n9064;
  assign n9066 = ~n631 & n1303;
  assign n9067 = n1308 & ~n9066;
  assign n9068 = n1312 & ~n9067;
  assign n9069 = n1316 & ~n9068;
  assign n9070 = n1320 & ~n9069;
  assign n9071 = n1324 & ~n9070;
  assign n9072 = n1328 & ~n9071;
  assign n9073 = n1332 & ~n9072;
  assign n9074 = n1336 & ~n9073;
  assign n9075 = n1340 & ~n9074;
  assign n9076 = n1344 & ~n9075;
  assign n9077 = n1348 & ~n9076;
  assign n9078 = n1352 & ~n9077;
  assign n9079 = n1356 & ~n9078;
  assign n9080 = n1360 & ~n9079;
  assign n9081 = n1364 & ~n9080;
  assign n9082 = n1368 & ~n9081;
  assign n9083 = n1372 & ~n9082;
  assign n9084 = n1376 & ~n9083;
  assign n9085 = n1380 & ~n9084;
  assign n9086 = n1384 & ~n9085;
  assign n9087 = n1388 & ~n9086;
  assign n9088 = n1392 & ~n9087;
  assign n9089 = n1396 & ~n9088;
  assign n9090 = n1663 & ~n9089;
  assign n9091 = n392 & ~n9090;
  assign n9092 = n396 & ~n9091;
  assign n9093 = n400 & ~n9092;
  assign n9094 = n404 & ~n9093;
  assign n9095 = n408 & ~n9094;
  assign n9096 = n412 & ~n9095;
  assign n9097 = n416 & ~n9096;
  assign n9098 = n420 & ~n9097;
  assign n9099 = n424 & ~n9098;
  assign n9100 = n428 & ~n9099;
  assign n9101 = n432 & ~n9100;
  assign n9102 = n436 & ~n9101;
  assign n9103 = n440 & ~n9102;
  assign n9104 = n444 & ~n9103;
  assign n9105 = n448 & ~n9104;
  assign n9106 = n452 & ~n9105;
  assign n9107 = n456 & ~n9106;
  assign n9108 = n460 & ~n9107;
  assign n9109 = n464 & ~n9108;
  assign n9110 = n468 & ~n9109;
  assign n9111 = n472 & ~n9110;
  assign n9112 = n476 & ~n9111;
  assign n9113 = n480 & ~n9112;
  assign n9114 = n484 & ~n9113;
  assign n9115 = n488 & ~n9114;
  assign n9116 = n492 & ~n9115;
  assign n9117 = n496 & ~n9116;
  assign n9118 = n500 & ~n9117;
  assign n9119 = n504 & ~n9118;
  assign n9120 = n508 & ~n9119;
  assign n9121 = n512 & ~n9120;
  assign n9122 = n516 & ~n9121;
  assign n9123 = n520 & ~n9122;
  assign n9124 = n524 & ~n9123;
  assign n9125 = n528 & ~n9124;
  assign n9126 = n532 & ~n9125;
  assign n9127 = n536 & ~n9126;
  assign n9128 = n540 & ~n9127;
  assign n9129 = n544 & ~n9128;
  assign n9130 = n548 & ~n9129;
  assign n9131 = n552 & ~n9130;
  assign n9132 = n556 & ~n9131;
  assign n9133 = n560 & ~n9132;
  assign n9134 = n564 & ~n9133;
  assign n9135 = n568 & ~n9134;
  assign n9136 = n572 & ~n9135;
  assign n9137 = n576 & ~n9136;
  assign n9138 = n580 & ~n9137;
  assign n9139 = n584 & ~n9138;
  assign n9140 = n588 & ~n9139;
  assign n9141 = n592 & ~n9140;
  assign n9142 = n596 & ~n9141;
  assign n9143 = n600 & ~n9142;
  assign n9144 = n604 & ~n9143;
  assign n9145 = n608 & ~n9144;
  assign n9146 = n612 & ~n9145;
  assign n9147 = n616 & ~n9146;
  assign n9148 = n620 & ~n9147;
  assign n9149 = n624 & ~n9148;
  assign n9150 = pi220  & ~n626;
  assign po92  = ~n9149 & n9150;
  assign n9152 = n635 & ~n970;
  assign n9153 = n640 & ~n9152;
  assign n9154 = n644 & ~n9153;
  assign n9155 = n648 & ~n9154;
  assign n9156 = n652 & ~n9155;
  assign n9157 = n656 & ~n9156;
  assign n9158 = n660 & ~n9157;
  assign n9159 = n664 & ~n9158;
  assign n9160 = n668 & ~n9159;
  assign n9161 = n672 & ~n9160;
  assign n9162 = n676 & ~n9161;
  assign n9163 = n680 & ~n9162;
  assign n9164 = n684 & ~n9163;
  assign n9165 = n688 & ~n9164;
  assign n9166 = n692 & ~n9165;
  assign n9167 = n696 & ~n9166;
  assign n9168 = n700 & ~n9167;
  assign n9169 = n704 & ~n9168;
  assign n9170 = n708 & ~n9169;
  assign n9171 = n712 & ~n9170;
  assign n9172 = n716 & ~n9171;
  assign n9173 = n720 & ~n9172;
  assign n9174 = n1484 & ~n9173;
  assign n9175 = n1486 & ~n9174;
  assign n9176 = n1750 & ~n9175;
  assign n9177 = n731 & ~n9176;
  assign n9178 = n735 & ~n9177;
  assign n9179 = n739 & ~n9178;
  assign n9180 = n743 & ~n9179;
  assign n9181 = n747 & ~n9180;
  assign n9182 = n751 & ~n9181;
  assign n9183 = n755 & ~n9182;
  assign n9184 = n759 & ~n9183;
  assign n9185 = n763 & ~n9184;
  assign n9186 = n767 & ~n9185;
  assign n9187 = n771 & ~n9186;
  assign n9188 = n775 & ~n9187;
  assign n9189 = n779 & ~n9188;
  assign n9190 = n783 & ~n9189;
  assign n9191 = n787 & ~n9190;
  assign n9192 = n791 & ~n9191;
  assign n9193 = n795 & ~n9192;
  assign n9194 = n799 & ~n9193;
  assign n9195 = n803 & ~n9194;
  assign n9196 = n807 & ~n9195;
  assign n9197 = n811 & ~n9196;
  assign n9198 = n815 & ~n9197;
  assign n9199 = n819 & ~n9198;
  assign n9200 = n823 & ~n9199;
  assign n9201 = n827 & ~n9200;
  assign n9202 = n831 & ~n9201;
  assign n9203 = n835 & ~n9202;
  assign n9204 = n839 & ~n9203;
  assign n9205 = n843 & ~n9204;
  assign n9206 = n847 & ~n9205;
  assign n9207 = n851 & ~n9206;
  assign n9208 = n855 & ~n9207;
  assign n9209 = n859 & ~n9208;
  assign n9210 = n863 & ~n9209;
  assign n9211 = n867 & ~n9210;
  assign n9212 = n871 & ~n9211;
  assign n9213 = n875 & ~n9212;
  assign n9214 = n879 & ~n9213;
  assign n9215 = n883 & ~n9214;
  assign n9216 = n887 & ~n9215;
  assign n9217 = n891 & ~n9216;
  assign n9218 = n895 & ~n9217;
  assign n9219 = n899 & ~n9218;
  assign n9220 = n903 & ~n9219;
  assign n9221 = n907 & ~n9220;
  assign n9222 = n911 & ~n9221;
  assign n9223 = n915 & ~n9222;
  assign n9224 = n919 & ~n9223;
  assign n9225 = n923 & ~n9224;
  assign n9226 = n927 & ~n9225;
  assign n9227 = n931 & ~n9226;
  assign n9228 = n935 & ~n9227;
  assign n9229 = n939 & ~n9228;
  assign n9230 = n943 & ~n9229;
  assign n9231 = n947 & ~n9230;
  assign n9232 = n951 & ~n9231;
  assign n9233 = n955 & ~n9232;
  assign n9234 = n959 & ~n9233;
  assign n9235 = n963 & ~n9234;
  assign n9236 = pi221  & ~n965;
  assign po93  = ~n9235 & n9236;
  assign n9238 = n974 & ~n1307;
  assign n9239 = n979 & ~n9238;
  assign n9240 = n983 & ~n9239;
  assign n9241 = n987 & ~n9240;
  assign n9242 = n991 & ~n9241;
  assign n9243 = n995 & ~n9242;
  assign n9244 = n999 & ~n9243;
  assign n9245 = n1003 & ~n9244;
  assign n9246 = n1007 & ~n9245;
  assign n9247 = n1011 & ~n9246;
  assign n9248 = n1015 & ~n9247;
  assign n9249 = n1019 & ~n9248;
  assign n9250 = n1023 & ~n9249;
  assign n9251 = n1027 & ~n9250;
  assign n9252 = n1031 & ~n9251;
  assign n9253 = n1035 & ~n9252;
  assign n9254 = n1039 & ~n9253;
  assign n9255 = n1043 & ~n9254;
  assign n9256 = n1047 & ~n9255;
  assign n9257 = n1051 & ~n9256;
  assign n9258 = n1055 & ~n9257;
  assign n9259 = n1059 & ~n9258;
  assign n9260 = n1574 & ~n9259;
  assign n9261 = n1576 & ~n9260;
  assign n9262 = n1837 & ~n9261;
  assign n9263 = n1068 & ~n9262;
  assign n9264 = n1072 & ~n9263;
  assign n9265 = n1076 & ~n9264;
  assign n9266 = n1080 & ~n9265;
  assign n9267 = n1084 & ~n9266;
  assign n9268 = n1088 & ~n9267;
  assign n9269 = n1092 & ~n9268;
  assign n9270 = n1096 & ~n9269;
  assign n9271 = n1100 & ~n9270;
  assign n9272 = n1104 & ~n9271;
  assign n9273 = n1108 & ~n9272;
  assign n9274 = n1112 & ~n9273;
  assign n9275 = n1116 & ~n9274;
  assign n9276 = n1120 & ~n9275;
  assign n9277 = n1124 & ~n9276;
  assign n9278 = n1128 & ~n9277;
  assign n9279 = n1132 & ~n9278;
  assign n9280 = n1136 & ~n9279;
  assign n9281 = n1140 & ~n9280;
  assign n9282 = n1144 & ~n9281;
  assign n9283 = n1148 & ~n9282;
  assign n9284 = n1152 & ~n9283;
  assign n9285 = n1156 & ~n9284;
  assign n9286 = n1160 & ~n9285;
  assign n9287 = n1164 & ~n9286;
  assign n9288 = n1168 & ~n9287;
  assign n9289 = n1172 & ~n9288;
  assign n9290 = n1176 & ~n9289;
  assign n9291 = n1180 & ~n9290;
  assign n9292 = n1184 & ~n9291;
  assign n9293 = n1188 & ~n9292;
  assign n9294 = n1192 & ~n9293;
  assign n9295 = n1196 & ~n9294;
  assign n9296 = n1200 & ~n9295;
  assign n9297 = n1204 & ~n9296;
  assign n9298 = n1208 & ~n9297;
  assign n9299 = n1212 & ~n9298;
  assign n9300 = n1216 & ~n9299;
  assign n9301 = n1220 & ~n9300;
  assign n9302 = n1224 & ~n9301;
  assign n9303 = n1228 & ~n9302;
  assign n9304 = n1232 & ~n9303;
  assign n9305 = n1236 & ~n9304;
  assign n9306 = n1240 & ~n9305;
  assign n9307 = n1244 & ~n9306;
  assign n9308 = n1248 & ~n9307;
  assign n9309 = n1252 & ~n9308;
  assign n9310 = n1256 & ~n9309;
  assign n9311 = n1260 & ~n9310;
  assign n9312 = n1264 & ~n9311;
  assign n9313 = n1268 & ~n9312;
  assign n9314 = n1272 & ~n9313;
  assign n9315 = n1276 & ~n9314;
  assign n9316 = n1280 & ~n9315;
  assign n9317 = n1284 & ~n9316;
  assign n9318 = n1288 & ~n9317;
  assign n9319 = n1292 & ~n9318;
  assign n9320 = n1296 & ~n9319;
  assign n9321 = n1300 & ~n9320;
  assign n9322 = pi222  & ~n1302;
  assign po94  = ~n9321 & n9322;
  assign n9324 = ~n639 & n1311;
  assign n9325 = n1316 & ~n9324;
  assign n9326 = n1320 & ~n9325;
  assign n9327 = n1324 & ~n9326;
  assign n9328 = n1328 & ~n9327;
  assign n9329 = n1332 & ~n9328;
  assign n9330 = n1336 & ~n9329;
  assign n9331 = n1340 & ~n9330;
  assign n9332 = n1344 & ~n9331;
  assign n9333 = n1348 & ~n9332;
  assign n9334 = n1352 & ~n9333;
  assign n9335 = n1356 & ~n9334;
  assign n9336 = n1360 & ~n9335;
  assign n9337 = n1364 & ~n9336;
  assign n9338 = n1368 & ~n9337;
  assign n9339 = n1372 & ~n9338;
  assign n9340 = n1376 & ~n9339;
  assign n9341 = n1380 & ~n9340;
  assign n9342 = n1384 & ~n9341;
  assign n9343 = n1388 & ~n9342;
  assign n9344 = n1392 & ~n9343;
  assign n9345 = n1396 & ~n9344;
  assign n9346 = n1663 & ~n9345;
  assign n9347 = n392 & ~n9346;
  assign n9348 = n396 & ~n9347;
  assign n9349 = n400 & ~n9348;
  assign n9350 = n404 & ~n9349;
  assign n9351 = n408 & ~n9350;
  assign n9352 = n412 & ~n9351;
  assign n9353 = n416 & ~n9352;
  assign n9354 = n420 & ~n9353;
  assign n9355 = n424 & ~n9354;
  assign n9356 = n428 & ~n9355;
  assign n9357 = n432 & ~n9356;
  assign n9358 = n436 & ~n9357;
  assign n9359 = n440 & ~n9358;
  assign n9360 = n444 & ~n9359;
  assign n9361 = n448 & ~n9360;
  assign n9362 = n452 & ~n9361;
  assign n9363 = n456 & ~n9362;
  assign n9364 = n460 & ~n9363;
  assign n9365 = n464 & ~n9364;
  assign n9366 = n468 & ~n9365;
  assign n9367 = n472 & ~n9366;
  assign n9368 = n476 & ~n9367;
  assign n9369 = n480 & ~n9368;
  assign n9370 = n484 & ~n9369;
  assign n9371 = n488 & ~n9370;
  assign n9372 = n492 & ~n9371;
  assign n9373 = n496 & ~n9372;
  assign n9374 = n500 & ~n9373;
  assign n9375 = n504 & ~n9374;
  assign n9376 = n508 & ~n9375;
  assign n9377 = n512 & ~n9376;
  assign n9378 = n516 & ~n9377;
  assign n9379 = n520 & ~n9378;
  assign n9380 = n524 & ~n9379;
  assign n9381 = n528 & ~n9380;
  assign n9382 = n532 & ~n9381;
  assign n9383 = n536 & ~n9382;
  assign n9384 = n540 & ~n9383;
  assign n9385 = n544 & ~n9384;
  assign n9386 = n548 & ~n9385;
  assign n9387 = n552 & ~n9386;
  assign n9388 = n556 & ~n9387;
  assign n9389 = n560 & ~n9388;
  assign n9390 = n564 & ~n9389;
  assign n9391 = n568 & ~n9390;
  assign n9392 = n572 & ~n9391;
  assign n9393 = n576 & ~n9392;
  assign n9394 = n580 & ~n9393;
  assign n9395 = n584 & ~n9394;
  assign n9396 = n588 & ~n9395;
  assign n9397 = n592 & ~n9396;
  assign n9398 = n596 & ~n9397;
  assign n9399 = n600 & ~n9398;
  assign n9400 = n604 & ~n9399;
  assign n9401 = n608 & ~n9400;
  assign n9402 = n612 & ~n9401;
  assign n9403 = n616 & ~n9402;
  assign n9404 = n620 & ~n9403;
  assign n9405 = n624 & ~n9404;
  assign n9406 = n628 & ~n9405;
  assign n9407 = n632 & ~n9406;
  assign n9408 = pi223  & ~n634;
  assign po95  = ~n9407 & n9408;
  assign n9410 = n643 & ~n978;
  assign n9411 = n648 & ~n9410;
  assign n9412 = n652 & ~n9411;
  assign n9413 = n656 & ~n9412;
  assign n9414 = n660 & ~n9413;
  assign n9415 = n664 & ~n9414;
  assign n9416 = n668 & ~n9415;
  assign n9417 = n672 & ~n9416;
  assign n9418 = n676 & ~n9417;
  assign n9419 = n680 & ~n9418;
  assign n9420 = n684 & ~n9419;
  assign n9421 = n688 & ~n9420;
  assign n9422 = n692 & ~n9421;
  assign n9423 = n696 & ~n9422;
  assign n9424 = n700 & ~n9423;
  assign n9425 = n704 & ~n9424;
  assign n9426 = n708 & ~n9425;
  assign n9427 = n712 & ~n9426;
  assign n9428 = n716 & ~n9427;
  assign n9429 = n720 & ~n9428;
  assign n9430 = n1484 & ~n9429;
  assign n9431 = n1486 & ~n9430;
  assign n9432 = n1750 & ~n9431;
  assign n9433 = n731 & ~n9432;
  assign n9434 = n735 & ~n9433;
  assign n9435 = n739 & ~n9434;
  assign n9436 = n743 & ~n9435;
  assign n9437 = n747 & ~n9436;
  assign n9438 = n751 & ~n9437;
  assign n9439 = n755 & ~n9438;
  assign n9440 = n759 & ~n9439;
  assign n9441 = n763 & ~n9440;
  assign n9442 = n767 & ~n9441;
  assign n9443 = n771 & ~n9442;
  assign n9444 = n775 & ~n9443;
  assign n9445 = n779 & ~n9444;
  assign n9446 = n783 & ~n9445;
  assign n9447 = n787 & ~n9446;
  assign n9448 = n791 & ~n9447;
  assign n9449 = n795 & ~n9448;
  assign n9450 = n799 & ~n9449;
  assign n9451 = n803 & ~n9450;
  assign n9452 = n807 & ~n9451;
  assign n9453 = n811 & ~n9452;
  assign n9454 = n815 & ~n9453;
  assign n9455 = n819 & ~n9454;
  assign n9456 = n823 & ~n9455;
  assign n9457 = n827 & ~n9456;
  assign n9458 = n831 & ~n9457;
  assign n9459 = n835 & ~n9458;
  assign n9460 = n839 & ~n9459;
  assign n9461 = n843 & ~n9460;
  assign n9462 = n847 & ~n9461;
  assign n9463 = n851 & ~n9462;
  assign n9464 = n855 & ~n9463;
  assign n9465 = n859 & ~n9464;
  assign n9466 = n863 & ~n9465;
  assign n9467 = n867 & ~n9466;
  assign n9468 = n871 & ~n9467;
  assign n9469 = n875 & ~n9468;
  assign n9470 = n879 & ~n9469;
  assign n9471 = n883 & ~n9470;
  assign n9472 = n887 & ~n9471;
  assign n9473 = n891 & ~n9472;
  assign n9474 = n895 & ~n9473;
  assign n9475 = n899 & ~n9474;
  assign n9476 = n903 & ~n9475;
  assign n9477 = n907 & ~n9476;
  assign n9478 = n911 & ~n9477;
  assign n9479 = n915 & ~n9478;
  assign n9480 = n919 & ~n9479;
  assign n9481 = n923 & ~n9480;
  assign n9482 = n927 & ~n9481;
  assign n9483 = n931 & ~n9482;
  assign n9484 = n935 & ~n9483;
  assign n9485 = n939 & ~n9484;
  assign n9486 = n943 & ~n9485;
  assign n9487 = n947 & ~n9486;
  assign n9488 = n951 & ~n9487;
  assign n9489 = n955 & ~n9488;
  assign n9490 = n959 & ~n9489;
  assign n9491 = n963 & ~n9490;
  assign n9492 = n967 & ~n9491;
  assign n9493 = n971 & ~n9492;
  assign n9494 = pi224  & ~n973;
  assign po96  = ~n9493 & n9494;
  assign n9496 = n982 & ~n1315;
  assign n9497 = n987 & ~n9496;
  assign n9498 = n991 & ~n9497;
  assign n9499 = n995 & ~n9498;
  assign n9500 = n999 & ~n9499;
  assign n9501 = n1003 & ~n9500;
  assign n9502 = n1007 & ~n9501;
  assign n9503 = n1011 & ~n9502;
  assign n9504 = n1015 & ~n9503;
  assign n9505 = n1019 & ~n9504;
  assign n9506 = n1023 & ~n9505;
  assign n9507 = n1027 & ~n9506;
  assign n9508 = n1031 & ~n9507;
  assign n9509 = n1035 & ~n9508;
  assign n9510 = n1039 & ~n9509;
  assign n9511 = n1043 & ~n9510;
  assign n9512 = n1047 & ~n9511;
  assign n9513 = n1051 & ~n9512;
  assign n9514 = n1055 & ~n9513;
  assign n9515 = n1059 & ~n9514;
  assign n9516 = n1574 & ~n9515;
  assign n9517 = n1576 & ~n9516;
  assign n9518 = n1837 & ~n9517;
  assign n9519 = n1068 & ~n9518;
  assign n9520 = n1072 & ~n9519;
  assign n9521 = n1076 & ~n9520;
  assign n9522 = n1080 & ~n9521;
  assign n9523 = n1084 & ~n9522;
  assign n9524 = n1088 & ~n9523;
  assign n9525 = n1092 & ~n9524;
  assign n9526 = n1096 & ~n9525;
  assign n9527 = n1100 & ~n9526;
  assign n9528 = n1104 & ~n9527;
  assign n9529 = n1108 & ~n9528;
  assign n9530 = n1112 & ~n9529;
  assign n9531 = n1116 & ~n9530;
  assign n9532 = n1120 & ~n9531;
  assign n9533 = n1124 & ~n9532;
  assign n9534 = n1128 & ~n9533;
  assign n9535 = n1132 & ~n9534;
  assign n9536 = n1136 & ~n9535;
  assign n9537 = n1140 & ~n9536;
  assign n9538 = n1144 & ~n9537;
  assign n9539 = n1148 & ~n9538;
  assign n9540 = n1152 & ~n9539;
  assign n9541 = n1156 & ~n9540;
  assign n9542 = n1160 & ~n9541;
  assign n9543 = n1164 & ~n9542;
  assign n9544 = n1168 & ~n9543;
  assign n9545 = n1172 & ~n9544;
  assign n9546 = n1176 & ~n9545;
  assign n9547 = n1180 & ~n9546;
  assign n9548 = n1184 & ~n9547;
  assign n9549 = n1188 & ~n9548;
  assign n9550 = n1192 & ~n9549;
  assign n9551 = n1196 & ~n9550;
  assign n9552 = n1200 & ~n9551;
  assign n9553 = n1204 & ~n9552;
  assign n9554 = n1208 & ~n9553;
  assign n9555 = n1212 & ~n9554;
  assign n9556 = n1216 & ~n9555;
  assign n9557 = n1220 & ~n9556;
  assign n9558 = n1224 & ~n9557;
  assign n9559 = n1228 & ~n9558;
  assign n9560 = n1232 & ~n9559;
  assign n9561 = n1236 & ~n9560;
  assign n9562 = n1240 & ~n9561;
  assign n9563 = n1244 & ~n9562;
  assign n9564 = n1248 & ~n9563;
  assign n9565 = n1252 & ~n9564;
  assign n9566 = n1256 & ~n9565;
  assign n9567 = n1260 & ~n9566;
  assign n9568 = n1264 & ~n9567;
  assign n9569 = n1268 & ~n9568;
  assign n9570 = n1272 & ~n9569;
  assign n9571 = n1276 & ~n9570;
  assign n9572 = n1280 & ~n9571;
  assign n9573 = n1284 & ~n9572;
  assign n9574 = n1288 & ~n9573;
  assign n9575 = n1292 & ~n9574;
  assign n9576 = n1296 & ~n9575;
  assign n9577 = n1300 & ~n9576;
  assign n9578 = n1304 & ~n9577;
  assign n9579 = n1308 & ~n9578;
  assign n9580 = pi225  & ~n1310;
  assign po97  = ~n9579 & n9580;
  assign n9582 = ~n647 & n1319;
  assign n9583 = n1324 & ~n9582;
  assign n9584 = n1328 & ~n9583;
  assign n9585 = n1332 & ~n9584;
  assign n9586 = n1336 & ~n9585;
  assign n9587 = n1340 & ~n9586;
  assign n9588 = n1344 & ~n9587;
  assign n9589 = n1348 & ~n9588;
  assign n9590 = n1352 & ~n9589;
  assign n9591 = n1356 & ~n9590;
  assign n9592 = n1360 & ~n9591;
  assign n9593 = n1364 & ~n9592;
  assign n9594 = n1368 & ~n9593;
  assign n9595 = n1372 & ~n9594;
  assign n9596 = n1376 & ~n9595;
  assign n9597 = n1380 & ~n9596;
  assign n9598 = n1384 & ~n9597;
  assign n9599 = n1388 & ~n9598;
  assign n9600 = n1392 & ~n9599;
  assign n9601 = n1396 & ~n9600;
  assign n9602 = n1663 & ~n9601;
  assign n9603 = n392 & ~n9602;
  assign n9604 = n396 & ~n9603;
  assign n9605 = n400 & ~n9604;
  assign n9606 = n404 & ~n9605;
  assign n9607 = n408 & ~n9606;
  assign n9608 = n412 & ~n9607;
  assign n9609 = n416 & ~n9608;
  assign n9610 = n420 & ~n9609;
  assign n9611 = n424 & ~n9610;
  assign n9612 = n428 & ~n9611;
  assign n9613 = n432 & ~n9612;
  assign n9614 = n436 & ~n9613;
  assign n9615 = n440 & ~n9614;
  assign n9616 = n444 & ~n9615;
  assign n9617 = n448 & ~n9616;
  assign n9618 = n452 & ~n9617;
  assign n9619 = n456 & ~n9618;
  assign n9620 = n460 & ~n9619;
  assign n9621 = n464 & ~n9620;
  assign n9622 = n468 & ~n9621;
  assign n9623 = n472 & ~n9622;
  assign n9624 = n476 & ~n9623;
  assign n9625 = n480 & ~n9624;
  assign n9626 = n484 & ~n9625;
  assign n9627 = n488 & ~n9626;
  assign n9628 = n492 & ~n9627;
  assign n9629 = n496 & ~n9628;
  assign n9630 = n500 & ~n9629;
  assign n9631 = n504 & ~n9630;
  assign n9632 = n508 & ~n9631;
  assign n9633 = n512 & ~n9632;
  assign n9634 = n516 & ~n9633;
  assign n9635 = n520 & ~n9634;
  assign n9636 = n524 & ~n9635;
  assign n9637 = n528 & ~n9636;
  assign n9638 = n532 & ~n9637;
  assign n9639 = n536 & ~n9638;
  assign n9640 = n540 & ~n9639;
  assign n9641 = n544 & ~n9640;
  assign n9642 = n548 & ~n9641;
  assign n9643 = n552 & ~n9642;
  assign n9644 = n556 & ~n9643;
  assign n9645 = n560 & ~n9644;
  assign n9646 = n564 & ~n9645;
  assign n9647 = n568 & ~n9646;
  assign n9648 = n572 & ~n9647;
  assign n9649 = n576 & ~n9648;
  assign n9650 = n580 & ~n9649;
  assign n9651 = n584 & ~n9650;
  assign n9652 = n588 & ~n9651;
  assign n9653 = n592 & ~n9652;
  assign n9654 = n596 & ~n9653;
  assign n9655 = n600 & ~n9654;
  assign n9656 = n604 & ~n9655;
  assign n9657 = n608 & ~n9656;
  assign n9658 = n612 & ~n9657;
  assign n9659 = n616 & ~n9658;
  assign n9660 = n620 & ~n9659;
  assign n9661 = n624 & ~n9660;
  assign n9662 = n628 & ~n9661;
  assign n9663 = n632 & ~n9662;
  assign n9664 = n636 & ~n9663;
  assign n9665 = n640 & ~n9664;
  assign n9666 = pi226  & ~n642;
  assign po98  = ~n9665 & n9666;
  assign n9668 = n651 & ~n986;
  assign n9669 = n656 & ~n9668;
  assign n9670 = n660 & ~n9669;
  assign n9671 = n664 & ~n9670;
  assign n9672 = n668 & ~n9671;
  assign n9673 = n672 & ~n9672;
  assign n9674 = n676 & ~n9673;
  assign n9675 = n680 & ~n9674;
  assign n9676 = n684 & ~n9675;
  assign n9677 = n688 & ~n9676;
  assign n9678 = n692 & ~n9677;
  assign n9679 = n696 & ~n9678;
  assign n9680 = n700 & ~n9679;
  assign n9681 = n704 & ~n9680;
  assign n9682 = n708 & ~n9681;
  assign n9683 = n712 & ~n9682;
  assign n9684 = n716 & ~n9683;
  assign n9685 = n720 & ~n9684;
  assign n9686 = n1484 & ~n9685;
  assign n9687 = n1486 & ~n9686;
  assign n9688 = n1750 & ~n9687;
  assign n9689 = n731 & ~n9688;
  assign n9690 = n735 & ~n9689;
  assign n9691 = n739 & ~n9690;
  assign n9692 = n743 & ~n9691;
  assign n9693 = n747 & ~n9692;
  assign n9694 = n751 & ~n9693;
  assign n9695 = n755 & ~n9694;
  assign n9696 = n759 & ~n9695;
  assign n9697 = n763 & ~n9696;
  assign n9698 = n767 & ~n9697;
  assign n9699 = n771 & ~n9698;
  assign n9700 = n775 & ~n9699;
  assign n9701 = n779 & ~n9700;
  assign n9702 = n783 & ~n9701;
  assign n9703 = n787 & ~n9702;
  assign n9704 = n791 & ~n9703;
  assign n9705 = n795 & ~n9704;
  assign n9706 = n799 & ~n9705;
  assign n9707 = n803 & ~n9706;
  assign n9708 = n807 & ~n9707;
  assign n9709 = n811 & ~n9708;
  assign n9710 = n815 & ~n9709;
  assign n9711 = n819 & ~n9710;
  assign n9712 = n823 & ~n9711;
  assign n9713 = n827 & ~n9712;
  assign n9714 = n831 & ~n9713;
  assign n9715 = n835 & ~n9714;
  assign n9716 = n839 & ~n9715;
  assign n9717 = n843 & ~n9716;
  assign n9718 = n847 & ~n9717;
  assign n9719 = n851 & ~n9718;
  assign n9720 = n855 & ~n9719;
  assign n9721 = n859 & ~n9720;
  assign n9722 = n863 & ~n9721;
  assign n9723 = n867 & ~n9722;
  assign n9724 = n871 & ~n9723;
  assign n9725 = n875 & ~n9724;
  assign n9726 = n879 & ~n9725;
  assign n9727 = n883 & ~n9726;
  assign n9728 = n887 & ~n9727;
  assign n9729 = n891 & ~n9728;
  assign n9730 = n895 & ~n9729;
  assign n9731 = n899 & ~n9730;
  assign n9732 = n903 & ~n9731;
  assign n9733 = n907 & ~n9732;
  assign n9734 = n911 & ~n9733;
  assign n9735 = n915 & ~n9734;
  assign n9736 = n919 & ~n9735;
  assign n9737 = n923 & ~n9736;
  assign n9738 = n927 & ~n9737;
  assign n9739 = n931 & ~n9738;
  assign n9740 = n935 & ~n9739;
  assign n9741 = n939 & ~n9740;
  assign n9742 = n943 & ~n9741;
  assign n9743 = n947 & ~n9742;
  assign n9744 = n951 & ~n9743;
  assign n9745 = n955 & ~n9744;
  assign n9746 = n959 & ~n9745;
  assign n9747 = n963 & ~n9746;
  assign n9748 = n967 & ~n9747;
  assign n9749 = n971 & ~n9748;
  assign n9750 = n975 & ~n9749;
  assign n9751 = n979 & ~n9750;
  assign n9752 = pi227  & ~n981;
  assign po99  = ~n9751 & n9752;
  assign n9754 = n990 & ~n1323;
  assign n9755 = n995 & ~n9754;
  assign n9756 = n999 & ~n9755;
  assign n9757 = n1003 & ~n9756;
  assign n9758 = n1007 & ~n9757;
  assign n9759 = n1011 & ~n9758;
  assign n9760 = n1015 & ~n9759;
  assign n9761 = n1019 & ~n9760;
  assign n9762 = n1023 & ~n9761;
  assign n9763 = n1027 & ~n9762;
  assign n9764 = n1031 & ~n9763;
  assign n9765 = n1035 & ~n9764;
  assign n9766 = n1039 & ~n9765;
  assign n9767 = n1043 & ~n9766;
  assign n9768 = n1047 & ~n9767;
  assign n9769 = n1051 & ~n9768;
  assign n9770 = n1055 & ~n9769;
  assign n9771 = n1059 & ~n9770;
  assign n9772 = n1574 & ~n9771;
  assign n9773 = n1576 & ~n9772;
  assign n9774 = n1837 & ~n9773;
  assign n9775 = n1068 & ~n9774;
  assign n9776 = n1072 & ~n9775;
  assign n9777 = n1076 & ~n9776;
  assign n9778 = n1080 & ~n9777;
  assign n9779 = n1084 & ~n9778;
  assign n9780 = n1088 & ~n9779;
  assign n9781 = n1092 & ~n9780;
  assign n9782 = n1096 & ~n9781;
  assign n9783 = n1100 & ~n9782;
  assign n9784 = n1104 & ~n9783;
  assign n9785 = n1108 & ~n9784;
  assign n9786 = n1112 & ~n9785;
  assign n9787 = n1116 & ~n9786;
  assign n9788 = n1120 & ~n9787;
  assign n9789 = n1124 & ~n9788;
  assign n9790 = n1128 & ~n9789;
  assign n9791 = n1132 & ~n9790;
  assign n9792 = n1136 & ~n9791;
  assign n9793 = n1140 & ~n9792;
  assign n9794 = n1144 & ~n9793;
  assign n9795 = n1148 & ~n9794;
  assign n9796 = n1152 & ~n9795;
  assign n9797 = n1156 & ~n9796;
  assign n9798 = n1160 & ~n9797;
  assign n9799 = n1164 & ~n9798;
  assign n9800 = n1168 & ~n9799;
  assign n9801 = n1172 & ~n9800;
  assign n9802 = n1176 & ~n9801;
  assign n9803 = n1180 & ~n9802;
  assign n9804 = n1184 & ~n9803;
  assign n9805 = n1188 & ~n9804;
  assign n9806 = n1192 & ~n9805;
  assign n9807 = n1196 & ~n9806;
  assign n9808 = n1200 & ~n9807;
  assign n9809 = n1204 & ~n9808;
  assign n9810 = n1208 & ~n9809;
  assign n9811 = n1212 & ~n9810;
  assign n9812 = n1216 & ~n9811;
  assign n9813 = n1220 & ~n9812;
  assign n9814 = n1224 & ~n9813;
  assign n9815 = n1228 & ~n9814;
  assign n9816 = n1232 & ~n9815;
  assign n9817 = n1236 & ~n9816;
  assign n9818 = n1240 & ~n9817;
  assign n9819 = n1244 & ~n9818;
  assign n9820 = n1248 & ~n9819;
  assign n9821 = n1252 & ~n9820;
  assign n9822 = n1256 & ~n9821;
  assign n9823 = n1260 & ~n9822;
  assign n9824 = n1264 & ~n9823;
  assign n9825 = n1268 & ~n9824;
  assign n9826 = n1272 & ~n9825;
  assign n9827 = n1276 & ~n9826;
  assign n9828 = n1280 & ~n9827;
  assign n9829 = n1284 & ~n9828;
  assign n9830 = n1288 & ~n9829;
  assign n9831 = n1292 & ~n9830;
  assign n9832 = n1296 & ~n9831;
  assign n9833 = n1300 & ~n9832;
  assign n9834 = n1304 & ~n9833;
  assign n9835 = n1308 & ~n9834;
  assign n9836 = n1312 & ~n9835;
  assign n9837 = n1316 & ~n9836;
  assign n9838 = pi228  & ~n1318;
  assign po100  = ~n9837 & n9838;
  assign n9840 = ~n655 & n1327;
  assign n9841 = n1332 & ~n9840;
  assign n9842 = n1336 & ~n9841;
  assign n9843 = n1340 & ~n9842;
  assign n9844 = n1344 & ~n9843;
  assign n9845 = n1348 & ~n9844;
  assign n9846 = n1352 & ~n9845;
  assign n9847 = n1356 & ~n9846;
  assign n9848 = n1360 & ~n9847;
  assign n9849 = n1364 & ~n9848;
  assign n9850 = n1368 & ~n9849;
  assign n9851 = n1372 & ~n9850;
  assign n9852 = n1376 & ~n9851;
  assign n9853 = n1380 & ~n9852;
  assign n9854 = n1384 & ~n9853;
  assign n9855 = n1388 & ~n9854;
  assign n9856 = n1392 & ~n9855;
  assign n9857 = n1396 & ~n9856;
  assign n9858 = n1663 & ~n9857;
  assign n9859 = n392 & ~n9858;
  assign n9860 = n396 & ~n9859;
  assign n9861 = n400 & ~n9860;
  assign n9862 = n404 & ~n9861;
  assign n9863 = n408 & ~n9862;
  assign n9864 = n412 & ~n9863;
  assign n9865 = n416 & ~n9864;
  assign n9866 = n420 & ~n9865;
  assign n9867 = n424 & ~n9866;
  assign n9868 = n428 & ~n9867;
  assign n9869 = n432 & ~n9868;
  assign n9870 = n436 & ~n9869;
  assign n9871 = n440 & ~n9870;
  assign n9872 = n444 & ~n9871;
  assign n9873 = n448 & ~n9872;
  assign n9874 = n452 & ~n9873;
  assign n9875 = n456 & ~n9874;
  assign n9876 = n460 & ~n9875;
  assign n9877 = n464 & ~n9876;
  assign n9878 = n468 & ~n9877;
  assign n9879 = n472 & ~n9878;
  assign n9880 = n476 & ~n9879;
  assign n9881 = n480 & ~n9880;
  assign n9882 = n484 & ~n9881;
  assign n9883 = n488 & ~n9882;
  assign n9884 = n492 & ~n9883;
  assign n9885 = n496 & ~n9884;
  assign n9886 = n500 & ~n9885;
  assign n9887 = n504 & ~n9886;
  assign n9888 = n508 & ~n9887;
  assign n9889 = n512 & ~n9888;
  assign n9890 = n516 & ~n9889;
  assign n9891 = n520 & ~n9890;
  assign n9892 = n524 & ~n9891;
  assign n9893 = n528 & ~n9892;
  assign n9894 = n532 & ~n9893;
  assign n9895 = n536 & ~n9894;
  assign n9896 = n540 & ~n9895;
  assign n9897 = n544 & ~n9896;
  assign n9898 = n548 & ~n9897;
  assign n9899 = n552 & ~n9898;
  assign n9900 = n556 & ~n9899;
  assign n9901 = n560 & ~n9900;
  assign n9902 = n564 & ~n9901;
  assign n9903 = n568 & ~n9902;
  assign n9904 = n572 & ~n9903;
  assign n9905 = n576 & ~n9904;
  assign n9906 = n580 & ~n9905;
  assign n9907 = n584 & ~n9906;
  assign n9908 = n588 & ~n9907;
  assign n9909 = n592 & ~n9908;
  assign n9910 = n596 & ~n9909;
  assign n9911 = n600 & ~n9910;
  assign n9912 = n604 & ~n9911;
  assign n9913 = n608 & ~n9912;
  assign n9914 = n612 & ~n9913;
  assign n9915 = n616 & ~n9914;
  assign n9916 = n620 & ~n9915;
  assign n9917 = n624 & ~n9916;
  assign n9918 = n628 & ~n9917;
  assign n9919 = n632 & ~n9918;
  assign n9920 = n636 & ~n9919;
  assign n9921 = n640 & ~n9920;
  assign n9922 = n644 & ~n9921;
  assign n9923 = n648 & ~n9922;
  assign n9924 = pi229  & ~n650;
  assign po101  = ~n9923 & n9924;
  assign n9926 = n659 & ~n994;
  assign n9927 = n664 & ~n9926;
  assign n9928 = n668 & ~n9927;
  assign n9929 = n672 & ~n9928;
  assign n9930 = n676 & ~n9929;
  assign n9931 = n680 & ~n9930;
  assign n9932 = n684 & ~n9931;
  assign n9933 = n688 & ~n9932;
  assign n9934 = n692 & ~n9933;
  assign n9935 = n696 & ~n9934;
  assign n9936 = n700 & ~n9935;
  assign n9937 = n704 & ~n9936;
  assign n9938 = n708 & ~n9937;
  assign n9939 = n712 & ~n9938;
  assign n9940 = n716 & ~n9939;
  assign n9941 = n720 & ~n9940;
  assign n9942 = n1484 & ~n9941;
  assign n9943 = n1486 & ~n9942;
  assign n9944 = n1750 & ~n9943;
  assign n9945 = n731 & ~n9944;
  assign n9946 = n735 & ~n9945;
  assign n9947 = n739 & ~n9946;
  assign n9948 = n743 & ~n9947;
  assign n9949 = n747 & ~n9948;
  assign n9950 = n751 & ~n9949;
  assign n9951 = n755 & ~n9950;
  assign n9952 = n759 & ~n9951;
  assign n9953 = n763 & ~n9952;
  assign n9954 = n767 & ~n9953;
  assign n9955 = n771 & ~n9954;
  assign n9956 = n775 & ~n9955;
  assign n9957 = n779 & ~n9956;
  assign n9958 = n783 & ~n9957;
  assign n9959 = n787 & ~n9958;
  assign n9960 = n791 & ~n9959;
  assign n9961 = n795 & ~n9960;
  assign n9962 = n799 & ~n9961;
  assign n9963 = n803 & ~n9962;
  assign n9964 = n807 & ~n9963;
  assign n9965 = n811 & ~n9964;
  assign n9966 = n815 & ~n9965;
  assign n9967 = n819 & ~n9966;
  assign n9968 = n823 & ~n9967;
  assign n9969 = n827 & ~n9968;
  assign n9970 = n831 & ~n9969;
  assign n9971 = n835 & ~n9970;
  assign n9972 = n839 & ~n9971;
  assign n9973 = n843 & ~n9972;
  assign n9974 = n847 & ~n9973;
  assign n9975 = n851 & ~n9974;
  assign n9976 = n855 & ~n9975;
  assign n9977 = n859 & ~n9976;
  assign n9978 = n863 & ~n9977;
  assign n9979 = n867 & ~n9978;
  assign n9980 = n871 & ~n9979;
  assign n9981 = n875 & ~n9980;
  assign n9982 = n879 & ~n9981;
  assign n9983 = n883 & ~n9982;
  assign n9984 = n887 & ~n9983;
  assign n9985 = n891 & ~n9984;
  assign n9986 = n895 & ~n9985;
  assign n9987 = n899 & ~n9986;
  assign n9988 = n903 & ~n9987;
  assign n9989 = n907 & ~n9988;
  assign n9990 = n911 & ~n9989;
  assign n9991 = n915 & ~n9990;
  assign n9992 = n919 & ~n9991;
  assign n9993 = n923 & ~n9992;
  assign n9994 = n927 & ~n9993;
  assign n9995 = n931 & ~n9994;
  assign n9996 = n935 & ~n9995;
  assign n9997 = n939 & ~n9996;
  assign n9998 = n943 & ~n9997;
  assign n9999 = n947 & ~n9998;
  assign n10000 = n951 & ~n9999;
  assign n10001 = n955 & ~n10000;
  assign n10002 = n959 & ~n10001;
  assign n10003 = n963 & ~n10002;
  assign n10004 = n967 & ~n10003;
  assign n10005 = n971 & ~n10004;
  assign n10006 = n975 & ~n10005;
  assign n10007 = n979 & ~n10006;
  assign n10008 = n983 & ~n10007;
  assign n10009 = n987 & ~n10008;
  assign n10010 = pi230  & ~n989;
  assign po102  = ~n10009 & n10010;
  assign n10012 = n998 & ~n1331;
  assign n10013 = n1003 & ~n10012;
  assign n10014 = n1007 & ~n10013;
  assign n10015 = n1011 & ~n10014;
  assign n10016 = n1015 & ~n10015;
  assign n10017 = n1019 & ~n10016;
  assign n10018 = n1023 & ~n10017;
  assign n10019 = n1027 & ~n10018;
  assign n10020 = n1031 & ~n10019;
  assign n10021 = n1035 & ~n10020;
  assign n10022 = n1039 & ~n10021;
  assign n10023 = n1043 & ~n10022;
  assign n10024 = n1047 & ~n10023;
  assign n10025 = n1051 & ~n10024;
  assign n10026 = n1055 & ~n10025;
  assign n10027 = n1059 & ~n10026;
  assign n10028 = n1574 & ~n10027;
  assign n10029 = n1576 & ~n10028;
  assign n10030 = n1837 & ~n10029;
  assign n10031 = n1068 & ~n10030;
  assign n10032 = n1072 & ~n10031;
  assign n10033 = n1076 & ~n10032;
  assign n10034 = n1080 & ~n10033;
  assign n10035 = n1084 & ~n10034;
  assign n10036 = n1088 & ~n10035;
  assign n10037 = n1092 & ~n10036;
  assign n10038 = n1096 & ~n10037;
  assign n10039 = n1100 & ~n10038;
  assign n10040 = n1104 & ~n10039;
  assign n10041 = n1108 & ~n10040;
  assign n10042 = n1112 & ~n10041;
  assign n10043 = n1116 & ~n10042;
  assign n10044 = n1120 & ~n10043;
  assign n10045 = n1124 & ~n10044;
  assign n10046 = n1128 & ~n10045;
  assign n10047 = n1132 & ~n10046;
  assign n10048 = n1136 & ~n10047;
  assign n10049 = n1140 & ~n10048;
  assign n10050 = n1144 & ~n10049;
  assign n10051 = n1148 & ~n10050;
  assign n10052 = n1152 & ~n10051;
  assign n10053 = n1156 & ~n10052;
  assign n10054 = n1160 & ~n10053;
  assign n10055 = n1164 & ~n10054;
  assign n10056 = n1168 & ~n10055;
  assign n10057 = n1172 & ~n10056;
  assign n10058 = n1176 & ~n10057;
  assign n10059 = n1180 & ~n10058;
  assign n10060 = n1184 & ~n10059;
  assign n10061 = n1188 & ~n10060;
  assign n10062 = n1192 & ~n10061;
  assign n10063 = n1196 & ~n10062;
  assign n10064 = n1200 & ~n10063;
  assign n10065 = n1204 & ~n10064;
  assign n10066 = n1208 & ~n10065;
  assign n10067 = n1212 & ~n10066;
  assign n10068 = n1216 & ~n10067;
  assign n10069 = n1220 & ~n10068;
  assign n10070 = n1224 & ~n10069;
  assign n10071 = n1228 & ~n10070;
  assign n10072 = n1232 & ~n10071;
  assign n10073 = n1236 & ~n10072;
  assign n10074 = n1240 & ~n10073;
  assign n10075 = n1244 & ~n10074;
  assign n10076 = n1248 & ~n10075;
  assign n10077 = n1252 & ~n10076;
  assign n10078 = n1256 & ~n10077;
  assign n10079 = n1260 & ~n10078;
  assign n10080 = n1264 & ~n10079;
  assign n10081 = n1268 & ~n10080;
  assign n10082 = n1272 & ~n10081;
  assign n10083 = n1276 & ~n10082;
  assign n10084 = n1280 & ~n10083;
  assign n10085 = n1284 & ~n10084;
  assign n10086 = n1288 & ~n10085;
  assign n10087 = n1292 & ~n10086;
  assign n10088 = n1296 & ~n10087;
  assign n10089 = n1300 & ~n10088;
  assign n10090 = n1304 & ~n10089;
  assign n10091 = n1308 & ~n10090;
  assign n10092 = n1312 & ~n10091;
  assign n10093 = n1316 & ~n10092;
  assign n10094 = n1320 & ~n10093;
  assign n10095 = n1324 & ~n10094;
  assign n10096 = pi231  & ~n1326;
  assign po103  = ~n10095 & n10096;
  assign n10098 = ~n663 & n1335;
  assign n10099 = n1340 & ~n10098;
  assign n10100 = n1344 & ~n10099;
  assign n10101 = n1348 & ~n10100;
  assign n10102 = n1352 & ~n10101;
  assign n10103 = n1356 & ~n10102;
  assign n10104 = n1360 & ~n10103;
  assign n10105 = n1364 & ~n10104;
  assign n10106 = n1368 & ~n10105;
  assign n10107 = n1372 & ~n10106;
  assign n10108 = n1376 & ~n10107;
  assign n10109 = n1380 & ~n10108;
  assign n10110 = n1384 & ~n10109;
  assign n10111 = n1388 & ~n10110;
  assign n10112 = n1392 & ~n10111;
  assign n10113 = n1396 & ~n10112;
  assign n10114 = n1663 & ~n10113;
  assign n10115 = n392 & ~n10114;
  assign n10116 = n396 & ~n10115;
  assign n10117 = n400 & ~n10116;
  assign n10118 = n404 & ~n10117;
  assign n10119 = n408 & ~n10118;
  assign n10120 = n412 & ~n10119;
  assign n10121 = n416 & ~n10120;
  assign n10122 = n420 & ~n10121;
  assign n10123 = n424 & ~n10122;
  assign n10124 = n428 & ~n10123;
  assign n10125 = n432 & ~n10124;
  assign n10126 = n436 & ~n10125;
  assign n10127 = n440 & ~n10126;
  assign n10128 = n444 & ~n10127;
  assign n10129 = n448 & ~n10128;
  assign n10130 = n452 & ~n10129;
  assign n10131 = n456 & ~n10130;
  assign n10132 = n460 & ~n10131;
  assign n10133 = n464 & ~n10132;
  assign n10134 = n468 & ~n10133;
  assign n10135 = n472 & ~n10134;
  assign n10136 = n476 & ~n10135;
  assign n10137 = n480 & ~n10136;
  assign n10138 = n484 & ~n10137;
  assign n10139 = n488 & ~n10138;
  assign n10140 = n492 & ~n10139;
  assign n10141 = n496 & ~n10140;
  assign n10142 = n500 & ~n10141;
  assign n10143 = n504 & ~n10142;
  assign n10144 = n508 & ~n10143;
  assign n10145 = n512 & ~n10144;
  assign n10146 = n516 & ~n10145;
  assign n10147 = n520 & ~n10146;
  assign n10148 = n524 & ~n10147;
  assign n10149 = n528 & ~n10148;
  assign n10150 = n532 & ~n10149;
  assign n10151 = n536 & ~n10150;
  assign n10152 = n540 & ~n10151;
  assign n10153 = n544 & ~n10152;
  assign n10154 = n548 & ~n10153;
  assign n10155 = n552 & ~n10154;
  assign n10156 = n556 & ~n10155;
  assign n10157 = n560 & ~n10156;
  assign n10158 = n564 & ~n10157;
  assign n10159 = n568 & ~n10158;
  assign n10160 = n572 & ~n10159;
  assign n10161 = n576 & ~n10160;
  assign n10162 = n580 & ~n10161;
  assign n10163 = n584 & ~n10162;
  assign n10164 = n588 & ~n10163;
  assign n10165 = n592 & ~n10164;
  assign n10166 = n596 & ~n10165;
  assign n10167 = n600 & ~n10166;
  assign n10168 = n604 & ~n10167;
  assign n10169 = n608 & ~n10168;
  assign n10170 = n612 & ~n10169;
  assign n10171 = n616 & ~n10170;
  assign n10172 = n620 & ~n10171;
  assign n10173 = n624 & ~n10172;
  assign n10174 = n628 & ~n10173;
  assign n10175 = n632 & ~n10174;
  assign n10176 = n636 & ~n10175;
  assign n10177 = n640 & ~n10176;
  assign n10178 = n644 & ~n10177;
  assign n10179 = n648 & ~n10178;
  assign n10180 = n652 & ~n10179;
  assign n10181 = n656 & ~n10180;
  assign n10182 = pi232  & ~n658;
  assign po104  = ~n10181 & n10182;
  assign n10184 = n667 & ~n1002;
  assign n10185 = n672 & ~n10184;
  assign n10186 = n676 & ~n10185;
  assign n10187 = n680 & ~n10186;
  assign n10188 = n684 & ~n10187;
  assign n10189 = n688 & ~n10188;
  assign n10190 = n692 & ~n10189;
  assign n10191 = n696 & ~n10190;
  assign n10192 = n700 & ~n10191;
  assign n10193 = n704 & ~n10192;
  assign n10194 = n708 & ~n10193;
  assign n10195 = n712 & ~n10194;
  assign n10196 = n716 & ~n10195;
  assign n10197 = n720 & ~n10196;
  assign n10198 = n1484 & ~n10197;
  assign n10199 = n1486 & ~n10198;
  assign n10200 = n1750 & ~n10199;
  assign n10201 = n731 & ~n10200;
  assign n10202 = n735 & ~n10201;
  assign n10203 = n739 & ~n10202;
  assign n10204 = n743 & ~n10203;
  assign n10205 = n747 & ~n10204;
  assign n10206 = n751 & ~n10205;
  assign n10207 = n755 & ~n10206;
  assign n10208 = n759 & ~n10207;
  assign n10209 = n763 & ~n10208;
  assign n10210 = n767 & ~n10209;
  assign n10211 = n771 & ~n10210;
  assign n10212 = n775 & ~n10211;
  assign n10213 = n779 & ~n10212;
  assign n10214 = n783 & ~n10213;
  assign n10215 = n787 & ~n10214;
  assign n10216 = n791 & ~n10215;
  assign n10217 = n795 & ~n10216;
  assign n10218 = n799 & ~n10217;
  assign n10219 = n803 & ~n10218;
  assign n10220 = n807 & ~n10219;
  assign n10221 = n811 & ~n10220;
  assign n10222 = n815 & ~n10221;
  assign n10223 = n819 & ~n10222;
  assign n10224 = n823 & ~n10223;
  assign n10225 = n827 & ~n10224;
  assign n10226 = n831 & ~n10225;
  assign n10227 = n835 & ~n10226;
  assign n10228 = n839 & ~n10227;
  assign n10229 = n843 & ~n10228;
  assign n10230 = n847 & ~n10229;
  assign n10231 = n851 & ~n10230;
  assign n10232 = n855 & ~n10231;
  assign n10233 = n859 & ~n10232;
  assign n10234 = n863 & ~n10233;
  assign n10235 = n867 & ~n10234;
  assign n10236 = n871 & ~n10235;
  assign n10237 = n875 & ~n10236;
  assign n10238 = n879 & ~n10237;
  assign n10239 = n883 & ~n10238;
  assign n10240 = n887 & ~n10239;
  assign n10241 = n891 & ~n10240;
  assign n10242 = n895 & ~n10241;
  assign n10243 = n899 & ~n10242;
  assign n10244 = n903 & ~n10243;
  assign n10245 = n907 & ~n10244;
  assign n10246 = n911 & ~n10245;
  assign n10247 = n915 & ~n10246;
  assign n10248 = n919 & ~n10247;
  assign n10249 = n923 & ~n10248;
  assign n10250 = n927 & ~n10249;
  assign n10251 = n931 & ~n10250;
  assign n10252 = n935 & ~n10251;
  assign n10253 = n939 & ~n10252;
  assign n10254 = n943 & ~n10253;
  assign n10255 = n947 & ~n10254;
  assign n10256 = n951 & ~n10255;
  assign n10257 = n955 & ~n10256;
  assign n10258 = n959 & ~n10257;
  assign n10259 = n963 & ~n10258;
  assign n10260 = n967 & ~n10259;
  assign n10261 = n971 & ~n10260;
  assign n10262 = n975 & ~n10261;
  assign n10263 = n979 & ~n10262;
  assign n10264 = n983 & ~n10263;
  assign n10265 = n987 & ~n10264;
  assign n10266 = n991 & ~n10265;
  assign n10267 = n995 & ~n10266;
  assign n10268 = pi233  & ~n997;
  assign po105  = ~n10267 & n10268;
  assign n10270 = n1006 & ~n1339;
  assign n10271 = n1011 & ~n10270;
  assign n10272 = n1015 & ~n10271;
  assign n10273 = n1019 & ~n10272;
  assign n10274 = n1023 & ~n10273;
  assign n10275 = n1027 & ~n10274;
  assign n10276 = n1031 & ~n10275;
  assign n10277 = n1035 & ~n10276;
  assign n10278 = n1039 & ~n10277;
  assign n10279 = n1043 & ~n10278;
  assign n10280 = n1047 & ~n10279;
  assign n10281 = n1051 & ~n10280;
  assign n10282 = n1055 & ~n10281;
  assign n10283 = n1059 & ~n10282;
  assign n10284 = n1574 & ~n10283;
  assign n10285 = n1576 & ~n10284;
  assign n10286 = n1837 & ~n10285;
  assign n10287 = n1068 & ~n10286;
  assign n10288 = n1072 & ~n10287;
  assign n10289 = n1076 & ~n10288;
  assign n10290 = n1080 & ~n10289;
  assign n10291 = n1084 & ~n10290;
  assign n10292 = n1088 & ~n10291;
  assign n10293 = n1092 & ~n10292;
  assign n10294 = n1096 & ~n10293;
  assign n10295 = n1100 & ~n10294;
  assign n10296 = n1104 & ~n10295;
  assign n10297 = n1108 & ~n10296;
  assign n10298 = n1112 & ~n10297;
  assign n10299 = n1116 & ~n10298;
  assign n10300 = n1120 & ~n10299;
  assign n10301 = n1124 & ~n10300;
  assign n10302 = n1128 & ~n10301;
  assign n10303 = n1132 & ~n10302;
  assign n10304 = n1136 & ~n10303;
  assign n10305 = n1140 & ~n10304;
  assign n10306 = n1144 & ~n10305;
  assign n10307 = n1148 & ~n10306;
  assign n10308 = n1152 & ~n10307;
  assign n10309 = n1156 & ~n10308;
  assign n10310 = n1160 & ~n10309;
  assign n10311 = n1164 & ~n10310;
  assign n10312 = n1168 & ~n10311;
  assign n10313 = n1172 & ~n10312;
  assign n10314 = n1176 & ~n10313;
  assign n10315 = n1180 & ~n10314;
  assign n10316 = n1184 & ~n10315;
  assign n10317 = n1188 & ~n10316;
  assign n10318 = n1192 & ~n10317;
  assign n10319 = n1196 & ~n10318;
  assign n10320 = n1200 & ~n10319;
  assign n10321 = n1204 & ~n10320;
  assign n10322 = n1208 & ~n10321;
  assign n10323 = n1212 & ~n10322;
  assign n10324 = n1216 & ~n10323;
  assign n10325 = n1220 & ~n10324;
  assign n10326 = n1224 & ~n10325;
  assign n10327 = n1228 & ~n10326;
  assign n10328 = n1232 & ~n10327;
  assign n10329 = n1236 & ~n10328;
  assign n10330 = n1240 & ~n10329;
  assign n10331 = n1244 & ~n10330;
  assign n10332 = n1248 & ~n10331;
  assign n10333 = n1252 & ~n10332;
  assign n10334 = n1256 & ~n10333;
  assign n10335 = n1260 & ~n10334;
  assign n10336 = n1264 & ~n10335;
  assign n10337 = n1268 & ~n10336;
  assign n10338 = n1272 & ~n10337;
  assign n10339 = n1276 & ~n10338;
  assign n10340 = n1280 & ~n10339;
  assign n10341 = n1284 & ~n10340;
  assign n10342 = n1288 & ~n10341;
  assign n10343 = n1292 & ~n10342;
  assign n10344 = n1296 & ~n10343;
  assign n10345 = n1300 & ~n10344;
  assign n10346 = n1304 & ~n10345;
  assign n10347 = n1308 & ~n10346;
  assign n10348 = n1312 & ~n10347;
  assign n10349 = n1316 & ~n10348;
  assign n10350 = n1320 & ~n10349;
  assign n10351 = n1324 & ~n10350;
  assign n10352 = n1328 & ~n10351;
  assign n10353 = n1332 & ~n10352;
  assign n10354 = pi234  & ~n1334;
  assign po106  = ~n10353 & n10354;
  assign n10356 = ~n671 & n1343;
  assign n10357 = n1348 & ~n10356;
  assign n10358 = n1352 & ~n10357;
  assign n10359 = n1356 & ~n10358;
  assign n10360 = n1360 & ~n10359;
  assign n10361 = n1364 & ~n10360;
  assign n10362 = n1368 & ~n10361;
  assign n10363 = n1372 & ~n10362;
  assign n10364 = n1376 & ~n10363;
  assign n10365 = n1380 & ~n10364;
  assign n10366 = n1384 & ~n10365;
  assign n10367 = n1388 & ~n10366;
  assign n10368 = n1392 & ~n10367;
  assign n10369 = n1396 & ~n10368;
  assign n10370 = n1663 & ~n10369;
  assign n10371 = n392 & ~n10370;
  assign n10372 = n396 & ~n10371;
  assign n10373 = n400 & ~n10372;
  assign n10374 = n404 & ~n10373;
  assign n10375 = n408 & ~n10374;
  assign n10376 = n412 & ~n10375;
  assign n10377 = n416 & ~n10376;
  assign n10378 = n420 & ~n10377;
  assign n10379 = n424 & ~n10378;
  assign n10380 = n428 & ~n10379;
  assign n10381 = n432 & ~n10380;
  assign n10382 = n436 & ~n10381;
  assign n10383 = n440 & ~n10382;
  assign n10384 = n444 & ~n10383;
  assign n10385 = n448 & ~n10384;
  assign n10386 = n452 & ~n10385;
  assign n10387 = n456 & ~n10386;
  assign n10388 = n460 & ~n10387;
  assign n10389 = n464 & ~n10388;
  assign n10390 = n468 & ~n10389;
  assign n10391 = n472 & ~n10390;
  assign n10392 = n476 & ~n10391;
  assign n10393 = n480 & ~n10392;
  assign n10394 = n484 & ~n10393;
  assign n10395 = n488 & ~n10394;
  assign n10396 = n492 & ~n10395;
  assign n10397 = n496 & ~n10396;
  assign n10398 = n500 & ~n10397;
  assign n10399 = n504 & ~n10398;
  assign n10400 = n508 & ~n10399;
  assign n10401 = n512 & ~n10400;
  assign n10402 = n516 & ~n10401;
  assign n10403 = n520 & ~n10402;
  assign n10404 = n524 & ~n10403;
  assign n10405 = n528 & ~n10404;
  assign n10406 = n532 & ~n10405;
  assign n10407 = n536 & ~n10406;
  assign n10408 = n540 & ~n10407;
  assign n10409 = n544 & ~n10408;
  assign n10410 = n548 & ~n10409;
  assign n10411 = n552 & ~n10410;
  assign n10412 = n556 & ~n10411;
  assign n10413 = n560 & ~n10412;
  assign n10414 = n564 & ~n10413;
  assign n10415 = n568 & ~n10414;
  assign n10416 = n572 & ~n10415;
  assign n10417 = n576 & ~n10416;
  assign n10418 = n580 & ~n10417;
  assign n10419 = n584 & ~n10418;
  assign n10420 = n588 & ~n10419;
  assign n10421 = n592 & ~n10420;
  assign n10422 = n596 & ~n10421;
  assign n10423 = n600 & ~n10422;
  assign n10424 = n604 & ~n10423;
  assign n10425 = n608 & ~n10424;
  assign n10426 = n612 & ~n10425;
  assign n10427 = n616 & ~n10426;
  assign n10428 = n620 & ~n10427;
  assign n10429 = n624 & ~n10428;
  assign n10430 = n628 & ~n10429;
  assign n10431 = n632 & ~n10430;
  assign n10432 = n636 & ~n10431;
  assign n10433 = n640 & ~n10432;
  assign n10434 = n644 & ~n10433;
  assign n10435 = n648 & ~n10434;
  assign n10436 = n652 & ~n10435;
  assign n10437 = n656 & ~n10436;
  assign n10438 = n660 & ~n10437;
  assign n10439 = n664 & ~n10438;
  assign n10440 = pi235  & ~n666;
  assign po107  = ~n10439 & n10440;
  assign n10442 = n675 & ~n1010;
  assign n10443 = n680 & ~n10442;
  assign n10444 = n684 & ~n10443;
  assign n10445 = n688 & ~n10444;
  assign n10446 = n692 & ~n10445;
  assign n10447 = n696 & ~n10446;
  assign n10448 = n700 & ~n10447;
  assign n10449 = n704 & ~n10448;
  assign n10450 = n708 & ~n10449;
  assign n10451 = n712 & ~n10450;
  assign n10452 = n716 & ~n10451;
  assign n10453 = n720 & ~n10452;
  assign n10454 = n1484 & ~n10453;
  assign n10455 = n1486 & ~n10454;
  assign n10456 = n1750 & ~n10455;
  assign n10457 = n731 & ~n10456;
  assign n10458 = n735 & ~n10457;
  assign n10459 = n739 & ~n10458;
  assign n10460 = n743 & ~n10459;
  assign n10461 = n747 & ~n10460;
  assign n10462 = n751 & ~n10461;
  assign n10463 = n755 & ~n10462;
  assign n10464 = n759 & ~n10463;
  assign n10465 = n763 & ~n10464;
  assign n10466 = n767 & ~n10465;
  assign n10467 = n771 & ~n10466;
  assign n10468 = n775 & ~n10467;
  assign n10469 = n779 & ~n10468;
  assign n10470 = n783 & ~n10469;
  assign n10471 = n787 & ~n10470;
  assign n10472 = n791 & ~n10471;
  assign n10473 = n795 & ~n10472;
  assign n10474 = n799 & ~n10473;
  assign n10475 = n803 & ~n10474;
  assign n10476 = n807 & ~n10475;
  assign n10477 = n811 & ~n10476;
  assign n10478 = n815 & ~n10477;
  assign n10479 = n819 & ~n10478;
  assign n10480 = n823 & ~n10479;
  assign n10481 = n827 & ~n10480;
  assign n10482 = n831 & ~n10481;
  assign n10483 = n835 & ~n10482;
  assign n10484 = n839 & ~n10483;
  assign n10485 = n843 & ~n10484;
  assign n10486 = n847 & ~n10485;
  assign n10487 = n851 & ~n10486;
  assign n10488 = n855 & ~n10487;
  assign n10489 = n859 & ~n10488;
  assign n10490 = n863 & ~n10489;
  assign n10491 = n867 & ~n10490;
  assign n10492 = n871 & ~n10491;
  assign n10493 = n875 & ~n10492;
  assign n10494 = n879 & ~n10493;
  assign n10495 = n883 & ~n10494;
  assign n10496 = n887 & ~n10495;
  assign n10497 = n891 & ~n10496;
  assign n10498 = n895 & ~n10497;
  assign n10499 = n899 & ~n10498;
  assign n10500 = n903 & ~n10499;
  assign n10501 = n907 & ~n10500;
  assign n10502 = n911 & ~n10501;
  assign n10503 = n915 & ~n10502;
  assign n10504 = n919 & ~n10503;
  assign n10505 = n923 & ~n10504;
  assign n10506 = n927 & ~n10505;
  assign n10507 = n931 & ~n10506;
  assign n10508 = n935 & ~n10507;
  assign n10509 = n939 & ~n10508;
  assign n10510 = n943 & ~n10509;
  assign n10511 = n947 & ~n10510;
  assign n10512 = n951 & ~n10511;
  assign n10513 = n955 & ~n10512;
  assign n10514 = n959 & ~n10513;
  assign n10515 = n963 & ~n10514;
  assign n10516 = n967 & ~n10515;
  assign n10517 = n971 & ~n10516;
  assign n10518 = n975 & ~n10517;
  assign n10519 = n979 & ~n10518;
  assign n10520 = n983 & ~n10519;
  assign n10521 = n987 & ~n10520;
  assign n10522 = n991 & ~n10521;
  assign n10523 = n995 & ~n10522;
  assign n10524 = n999 & ~n10523;
  assign n10525 = n1003 & ~n10524;
  assign n10526 = pi236  & ~n1005;
  assign po108  = ~n10525 & n10526;
  assign n10528 = n1014 & ~n1347;
  assign n10529 = n1019 & ~n10528;
  assign n10530 = n1023 & ~n10529;
  assign n10531 = n1027 & ~n10530;
  assign n10532 = n1031 & ~n10531;
  assign n10533 = n1035 & ~n10532;
  assign n10534 = n1039 & ~n10533;
  assign n10535 = n1043 & ~n10534;
  assign n10536 = n1047 & ~n10535;
  assign n10537 = n1051 & ~n10536;
  assign n10538 = n1055 & ~n10537;
  assign n10539 = n1059 & ~n10538;
  assign n10540 = n1574 & ~n10539;
  assign n10541 = n1576 & ~n10540;
  assign n10542 = n1837 & ~n10541;
  assign n10543 = n1068 & ~n10542;
  assign n10544 = n1072 & ~n10543;
  assign n10545 = n1076 & ~n10544;
  assign n10546 = n1080 & ~n10545;
  assign n10547 = n1084 & ~n10546;
  assign n10548 = n1088 & ~n10547;
  assign n10549 = n1092 & ~n10548;
  assign n10550 = n1096 & ~n10549;
  assign n10551 = n1100 & ~n10550;
  assign n10552 = n1104 & ~n10551;
  assign n10553 = n1108 & ~n10552;
  assign n10554 = n1112 & ~n10553;
  assign n10555 = n1116 & ~n10554;
  assign n10556 = n1120 & ~n10555;
  assign n10557 = n1124 & ~n10556;
  assign n10558 = n1128 & ~n10557;
  assign n10559 = n1132 & ~n10558;
  assign n10560 = n1136 & ~n10559;
  assign n10561 = n1140 & ~n10560;
  assign n10562 = n1144 & ~n10561;
  assign n10563 = n1148 & ~n10562;
  assign n10564 = n1152 & ~n10563;
  assign n10565 = n1156 & ~n10564;
  assign n10566 = n1160 & ~n10565;
  assign n10567 = n1164 & ~n10566;
  assign n10568 = n1168 & ~n10567;
  assign n10569 = n1172 & ~n10568;
  assign n10570 = n1176 & ~n10569;
  assign n10571 = n1180 & ~n10570;
  assign n10572 = n1184 & ~n10571;
  assign n10573 = n1188 & ~n10572;
  assign n10574 = n1192 & ~n10573;
  assign n10575 = n1196 & ~n10574;
  assign n10576 = n1200 & ~n10575;
  assign n10577 = n1204 & ~n10576;
  assign n10578 = n1208 & ~n10577;
  assign n10579 = n1212 & ~n10578;
  assign n10580 = n1216 & ~n10579;
  assign n10581 = n1220 & ~n10580;
  assign n10582 = n1224 & ~n10581;
  assign n10583 = n1228 & ~n10582;
  assign n10584 = n1232 & ~n10583;
  assign n10585 = n1236 & ~n10584;
  assign n10586 = n1240 & ~n10585;
  assign n10587 = n1244 & ~n10586;
  assign n10588 = n1248 & ~n10587;
  assign n10589 = n1252 & ~n10588;
  assign n10590 = n1256 & ~n10589;
  assign n10591 = n1260 & ~n10590;
  assign n10592 = n1264 & ~n10591;
  assign n10593 = n1268 & ~n10592;
  assign n10594 = n1272 & ~n10593;
  assign n10595 = n1276 & ~n10594;
  assign n10596 = n1280 & ~n10595;
  assign n10597 = n1284 & ~n10596;
  assign n10598 = n1288 & ~n10597;
  assign n10599 = n1292 & ~n10598;
  assign n10600 = n1296 & ~n10599;
  assign n10601 = n1300 & ~n10600;
  assign n10602 = n1304 & ~n10601;
  assign n10603 = n1308 & ~n10602;
  assign n10604 = n1312 & ~n10603;
  assign n10605 = n1316 & ~n10604;
  assign n10606 = n1320 & ~n10605;
  assign n10607 = n1324 & ~n10606;
  assign n10608 = n1328 & ~n10607;
  assign n10609 = n1332 & ~n10608;
  assign n10610 = n1336 & ~n10609;
  assign n10611 = n1340 & ~n10610;
  assign n10612 = pi237  & ~n1342;
  assign po109  = ~n10611 & n10612;
  assign n10614 = ~n679 & n1351;
  assign n10615 = n1356 & ~n10614;
  assign n10616 = n1360 & ~n10615;
  assign n10617 = n1364 & ~n10616;
  assign n10618 = n1368 & ~n10617;
  assign n10619 = n1372 & ~n10618;
  assign n10620 = n1376 & ~n10619;
  assign n10621 = n1380 & ~n10620;
  assign n10622 = n1384 & ~n10621;
  assign n10623 = n1388 & ~n10622;
  assign n10624 = n1392 & ~n10623;
  assign n10625 = n1396 & ~n10624;
  assign n10626 = n1663 & ~n10625;
  assign n10627 = n392 & ~n10626;
  assign n10628 = n396 & ~n10627;
  assign n10629 = n400 & ~n10628;
  assign n10630 = n404 & ~n10629;
  assign n10631 = n408 & ~n10630;
  assign n10632 = n412 & ~n10631;
  assign n10633 = n416 & ~n10632;
  assign n10634 = n420 & ~n10633;
  assign n10635 = n424 & ~n10634;
  assign n10636 = n428 & ~n10635;
  assign n10637 = n432 & ~n10636;
  assign n10638 = n436 & ~n10637;
  assign n10639 = n440 & ~n10638;
  assign n10640 = n444 & ~n10639;
  assign n10641 = n448 & ~n10640;
  assign n10642 = n452 & ~n10641;
  assign n10643 = n456 & ~n10642;
  assign n10644 = n460 & ~n10643;
  assign n10645 = n464 & ~n10644;
  assign n10646 = n468 & ~n10645;
  assign n10647 = n472 & ~n10646;
  assign n10648 = n476 & ~n10647;
  assign n10649 = n480 & ~n10648;
  assign n10650 = n484 & ~n10649;
  assign n10651 = n488 & ~n10650;
  assign n10652 = n492 & ~n10651;
  assign n10653 = n496 & ~n10652;
  assign n10654 = n500 & ~n10653;
  assign n10655 = n504 & ~n10654;
  assign n10656 = n508 & ~n10655;
  assign n10657 = n512 & ~n10656;
  assign n10658 = n516 & ~n10657;
  assign n10659 = n520 & ~n10658;
  assign n10660 = n524 & ~n10659;
  assign n10661 = n528 & ~n10660;
  assign n10662 = n532 & ~n10661;
  assign n10663 = n536 & ~n10662;
  assign n10664 = n540 & ~n10663;
  assign n10665 = n544 & ~n10664;
  assign n10666 = n548 & ~n10665;
  assign n10667 = n552 & ~n10666;
  assign n10668 = n556 & ~n10667;
  assign n10669 = n560 & ~n10668;
  assign n10670 = n564 & ~n10669;
  assign n10671 = n568 & ~n10670;
  assign n10672 = n572 & ~n10671;
  assign n10673 = n576 & ~n10672;
  assign n10674 = n580 & ~n10673;
  assign n10675 = n584 & ~n10674;
  assign n10676 = n588 & ~n10675;
  assign n10677 = n592 & ~n10676;
  assign n10678 = n596 & ~n10677;
  assign n10679 = n600 & ~n10678;
  assign n10680 = n604 & ~n10679;
  assign n10681 = n608 & ~n10680;
  assign n10682 = n612 & ~n10681;
  assign n10683 = n616 & ~n10682;
  assign n10684 = n620 & ~n10683;
  assign n10685 = n624 & ~n10684;
  assign n10686 = n628 & ~n10685;
  assign n10687 = n632 & ~n10686;
  assign n10688 = n636 & ~n10687;
  assign n10689 = n640 & ~n10688;
  assign n10690 = n644 & ~n10689;
  assign n10691 = n648 & ~n10690;
  assign n10692 = n652 & ~n10691;
  assign n10693 = n656 & ~n10692;
  assign n10694 = n660 & ~n10693;
  assign n10695 = n664 & ~n10694;
  assign n10696 = n668 & ~n10695;
  assign n10697 = n672 & ~n10696;
  assign n10698 = pi238  & ~n674;
  assign po110  = ~n10697 & n10698;
  assign n10700 = n683 & ~n1018;
  assign n10701 = n688 & ~n10700;
  assign n10702 = n692 & ~n10701;
  assign n10703 = n696 & ~n10702;
  assign n10704 = n700 & ~n10703;
  assign n10705 = n704 & ~n10704;
  assign n10706 = n708 & ~n10705;
  assign n10707 = n712 & ~n10706;
  assign n10708 = n716 & ~n10707;
  assign n10709 = n720 & ~n10708;
  assign n10710 = n1484 & ~n10709;
  assign n10711 = n1486 & ~n10710;
  assign n10712 = n1750 & ~n10711;
  assign n10713 = n731 & ~n10712;
  assign n10714 = n735 & ~n10713;
  assign n10715 = n739 & ~n10714;
  assign n10716 = n743 & ~n10715;
  assign n10717 = n747 & ~n10716;
  assign n10718 = n751 & ~n10717;
  assign n10719 = n755 & ~n10718;
  assign n10720 = n759 & ~n10719;
  assign n10721 = n763 & ~n10720;
  assign n10722 = n767 & ~n10721;
  assign n10723 = n771 & ~n10722;
  assign n10724 = n775 & ~n10723;
  assign n10725 = n779 & ~n10724;
  assign n10726 = n783 & ~n10725;
  assign n10727 = n787 & ~n10726;
  assign n10728 = n791 & ~n10727;
  assign n10729 = n795 & ~n10728;
  assign n10730 = n799 & ~n10729;
  assign n10731 = n803 & ~n10730;
  assign n10732 = n807 & ~n10731;
  assign n10733 = n811 & ~n10732;
  assign n10734 = n815 & ~n10733;
  assign n10735 = n819 & ~n10734;
  assign n10736 = n823 & ~n10735;
  assign n10737 = n827 & ~n10736;
  assign n10738 = n831 & ~n10737;
  assign n10739 = n835 & ~n10738;
  assign n10740 = n839 & ~n10739;
  assign n10741 = n843 & ~n10740;
  assign n10742 = n847 & ~n10741;
  assign n10743 = n851 & ~n10742;
  assign n10744 = n855 & ~n10743;
  assign n10745 = n859 & ~n10744;
  assign n10746 = n863 & ~n10745;
  assign n10747 = n867 & ~n10746;
  assign n10748 = n871 & ~n10747;
  assign n10749 = n875 & ~n10748;
  assign n10750 = n879 & ~n10749;
  assign n10751 = n883 & ~n10750;
  assign n10752 = n887 & ~n10751;
  assign n10753 = n891 & ~n10752;
  assign n10754 = n895 & ~n10753;
  assign n10755 = n899 & ~n10754;
  assign n10756 = n903 & ~n10755;
  assign n10757 = n907 & ~n10756;
  assign n10758 = n911 & ~n10757;
  assign n10759 = n915 & ~n10758;
  assign n10760 = n919 & ~n10759;
  assign n10761 = n923 & ~n10760;
  assign n10762 = n927 & ~n10761;
  assign n10763 = n931 & ~n10762;
  assign n10764 = n935 & ~n10763;
  assign n10765 = n939 & ~n10764;
  assign n10766 = n943 & ~n10765;
  assign n10767 = n947 & ~n10766;
  assign n10768 = n951 & ~n10767;
  assign n10769 = n955 & ~n10768;
  assign n10770 = n959 & ~n10769;
  assign n10771 = n963 & ~n10770;
  assign n10772 = n967 & ~n10771;
  assign n10773 = n971 & ~n10772;
  assign n10774 = n975 & ~n10773;
  assign n10775 = n979 & ~n10774;
  assign n10776 = n983 & ~n10775;
  assign n10777 = n987 & ~n10776;
  assign n10778 = n991 & ~n10777;
  assign n10779 = n995 & ~n10778;
  assign n10780 = n999 & ~n10779;
  assign n10781 = n1003 & ~n10780;
  assign n10782 = n1007 & ~n10781;
  assign n10783 = n1011 & ~n10782;
  assign n10784 = pi239  & ~n1013;
  assign po111  = ~n10783 & n10784;
  assign n10786 = n1022 & ~n1355;
  assign n10787 = n1027 & ~n10786;
  assign n10788 = n1031 & ~n10787;
  assign n10789 = n1035 & ~n10788;
  assign n10790 = n1039 & ~n10789;
  assign n10791 = n1043 & ~n10790;
  assign n10792 = n1047 & ~n10791;
  assign n10793 = n1051 & ~n10792;
  assign n10794 = n1055 & ~n10793;
  assign n10795 = n1059 & ~n10794;
  assign n10796 = n1574 & ~n10795;
  assign n10797 = n1576 & ~n10796;
  assign n10798 = n1837 & ~n10797;
  assign n10799 = n1068 & ~n10798;
  assign n10800 = n1072 & ~n10799;
  assign n10801 = n1076 & ~n10800;
  assign n10802 = n1080 & ~n10801;
  assign n10803 = n1084 & ~n10802;
  assign n10804 = n1088 & ~n10803;
  assign n10805 = n1092 & ~n10804;
  assign n10806 = n1096 & ~n10805;
  assign n10807 = n1100 & ~n10806;
  assign n10808 = n1104 & ~n10807;
  assign n10809 = n1108 & ~n10808;
  assign n10810 = n1112 & ~n10809;
  assign n10811 = n1116 & ~n10810;
  assign n10812 = n1120 & ~n10811;
  assign n10813 = n1124 & ~n10812;
  assign n10814 = n1128 & ~n10813;
  assign n10815 = n1132 & ~n10814;
  assign n10816 = n1136 & ~n10815;
  assign n10817 = n1140 & ~n10816;
  assign n10818 = n1144 & ~n10817;
  assign n10819 = n1148 & ~n10818;
  assign n10820 = n1152 & ~n10819;
  assign n10821 = n1156 & ~n10820;
  assign n10822 = n1160 & ~n10821;
  assign n10823 = n1164 & ~n10822;
  assign n10824 = n1168 & ~n10823;
  assign n10825 = n1172 & ~n10824;
  assign n10826 = n1176 & ~n10825;
  assign n10827 = n1180 & ~n10826;
  assign n10828 = n1184 & ~n10827;
  assign n10829 = n1188 & ~n10828;
  assign n10830 = n1192 & ~n10829;
  assign n10831 = n1196 & ~n10830;
  assign n10832 = n1200 & ~n10831;
  assign n10833 = n1204 & ~n10832;
  assign n10834 = n1208 & ~n10833;
  assign n10835 = n1212 & ~n10834;
  assign n10836 = n1216 & ~n10835;
  assign n10837 = n1220 & ~n10836;
  assign n10838 = n1224 & ~n10837;
  assign n10839 = n1228 & ~n10838;
  assign n10840 = n1232 & ~n10839;
  assign n10841 = n1236 & ~n10840;
  assign n10842 = n1240 & ~n10841;
  assign n10843 = n1244 & ~n10842;
  assign n10844 = n1248 & ~n10843;
  assign n10845 = n1252 & ~n10844;
  assign n10846 = n1256 & ~n10845;
  assign n10847 = n1260 & ~n10846;
  assign n10848 = n1264 & ~n10847;
  assign n10849 = n1268 & ~n10848;
  assign n10850 = n1272 & ~n10849;
  assign n10851 = n1276 & ~n10850;
  assign n10852 = n1280 & ~n10851;
  assign n10853 = n1284 & ~n10852;
  assign n10854 = n1288 & ~n10853;
  assign n10855 = n1292 & ~n10854;
  assign n10856 = n1296 & ~n10855;
  assign n10857 = n1300 & ~n10856;
  assign n10858 = n1304 & ~n10857;
  assign n10859 = n1308 & ~n10858;
  assign n10860 = n1312 & ~n10859;
  assign n10861 = n1316 & ~n10860;
  assign n10862 = n1320 & ~n10861;
  assign n10863 = n1324 & ~n10862;
  assign n10864 = n1328 & ~n10863;
  assign n10865 = n1332 & ~n10864;
  assign n10866 = n1336 & ~n10865;
  assign n10867 = n1340 & ~n10866;
  assign n10868 = n1344 & ~n10867;
  assign n10869 = n1348 & ~n10868;
  assign n10870 = pi240  & ~n1350;
  assign po112  = ~n10869 & n10870;
  assign n10872 = ~n687 & n1359;
  assign n10873 = n1364 & ~n10872;
  assign n10874 = n1368 & ~n10873;
  assign n10875 = n1372 & ~n10874;
  assign n10876 = n1376 & ~n10875;
  assign n10877 = n1380 & ~n10876;
  assign n10878 = n1384 & ~n10877;
  assign n10879 = n1388 & ~n10878;
  assign n10880 = n1392 & ~n10879;
  assign n10881 = n1396 & ~n10880;
  assign n10882 = n1663 & ~n10881;
  assign n10883 = n392 & ~n10882;
  assign n10884 = n396 & ~n10883;
  assign n10885 = n400 & ~n10884;
  assign n10886 = n404 & ~n10885;
  assign n10887 = n408 & ~n10886;
  assign n10888 = n412 & ~n10887;
  assign n10889 = n416 & ~n10888;
  assign n10890 = n420 & ~n10889;
  assign n10891 = n424 & ~n10890;
  assign n10892 = n428 & ~n10891;
  assign n10893 = n432 & ~n10892;
  assign n10894 = n436 & ~n10893;
  assign n10895 = n440 & ~n10894;
  assign n10896 = n444 & ~n10895;
  assign n10897 = n448 & ~n10896;
  assign n10898 = n452 & ~n10897;
  assign n10899 = n456 & ~n10898;
  assign n10900 = n460 & ~n10899;
  assign n10901 = n464 & ~n10900;
  assign n10902 = n468 & ~n10901;
  assign n10903 = n472 & ~n10902;
  assign n10904 = n476 & ~n10903;
  assign n10905 = n480 & ~n10904;
  assign n10906 = n484 & ~n10905;
  assign n10907 = n488 & ~n10906;
  assign n10908 = n492 & ~n10907;
  assign n10909 = n496 & ~n10908;
  assign n10910 = n500 & ~n10909;
  assign n10911 = n504 & ~n10910;
  assign n10912 = n508 & ~n10911;
  assign n10913 = n512 & ~n10912;
  assign n10914 = n516 & ~n10913;
  assign n10915 = n520 & ~n10914;
  assign n10916 = n524 & ~n10915;
  assign n10917 = n528 & ~n10916;
  assign n10918 = n532 & ~n10917;
  assign n10919 = n536 & ~n10918;
  assign n10920 = n540 & ~n10919;
  assign n10921 = n544 & ~n10920;
  assign n10922 = n548 & ~n10921;
  assign n10923 = n552 & ~n10922;
  assign n10924 = n556 & ~n10923;
  assign n10925 = n560 & ~n10924;
  assign n10926 = n564 & ~n10925;
  assign n10927 = n568 & ~n10926;
  assign n10928 = n572 & ~n10927;
  assign n10929 = n576 & ~n10928;
  assign n10930 = n580 & ~n10929;
  assign n10931 = n584 & ~n10930;
  assign n10932 = n588 & ~n10931;
  assign n10933 = n592 & ~n10932;
  assign n10934 = n596 & ~n10933;
  assign n10935 = n600 & ~n10934;
  assign n10936 = n604 & ~n10935;
  assign n10937 = n608 & ~n10936;
  assign n10938 = n612 & ~n10937;
  assign n10939 = n616 & ~n10938;
  assign n10940 = n620 & ~n10939;
  assign n10941 = n624 & ~n10940;
  assign n10942 = n628 & ~n10941;
  assign n10943 = n632 & ~n10942;
  assign n10944 = n636 & ~n10943;
  assign n10945 = n640 & ~n10944;
  assign n10946 = n644 & ~n10945;
  assign n10947 = n648 & ~n10946;
  assign n10948 = n652 & ~n10947;
  assign n10949 = n656 & ~n10948;
  assign n10950 = n660 & ~n10949;
  assign n10951 = n664 & ~n10950;
  assign n10952 = n668 & ~n10951;
  assign n10953 = n672 & ~n10952;
  assign n10954 = n676 & ~n10953;
  assign n10955 = n680 & ~n10954;
  assign n10956 = pi241  & ~n682;
  assign po113  = ~n10955 & n10956;
  assign n10958 = n691 & ~n1026;
  assign n10959 = n696 & ~n10958;
  assign n10960 = n700 & ~n10959;
  assign n10961 = n704 & ~n10960;
  assign n10962 = n708 & ~n10961;
  assign n10963 = n712 & ~n10962;
  assign n10964 = n716 & ~n10963;
  assign n10965 = n720 & ~n10964;
  assign n10966 = n1484 & ~n10965;
  assign n10967 = n1486 & ~n10966;
  assign n10968 = n1750 & ~n10967;
  assign n10969 = n731 & ~n10968;
  assign n10970 = n735 & ~n10969;
  assign n10971 = n739 & ~n10970;
  assign n10972 = n743 & ~n10971;
  assign n10973 = n747 & ~n10972;
  assign n10974 = n751 & ~n10973;
  assign n10975 = n755 & ~n10974;
  assign n10976 = n759 & ~n10975;
  assign n10977 = n763 & ~n10976;
  assign n10978 = n767 & ~n10977;
  assign n10979 = n771 & ~n10978;
  assign n10980 = n775 & ~n10979;
  assign n10981 = n779 & ~n10980;
  assign n10982 = n783 & ~n10981;
  assign n10983 = n787 & ~n10982;
  assign n10984 = n791 & ~n10983;
  assign n10985 = n795 & ~n10984;
  assign n10986 = n799 & ~n10985;
  assign n10987 = n803 & ~n10986;
  assign n10988 = n807 & ~n10987;
  assign n10989 = n811 & ~n10988;
  assign n10990 = n815 & ~n10989;
  assign n10991 = n819 & ~n10990;
  assign n10992 = n823 & ~n10991;
  assign n10993 = n827 & ~n10992;
  assign n10994 = n831 & ~n10993;
  assign n10995 = n835 & ~n10994;
  assign n10996 = n839 & ~n10995;
  assign n10997 = n843 & ~n10996;
  assign n10998 = n847 & ~n10997;
  assign n10999 = n851 & ~n10998;
  assign n11000 = n855 & ~n10999;
  assign n11001 = n859 & ~n11000;
  assign n11002 = n863 & ~n11001;
  assign n11003 = n867 & ~n11002;
  assign n11004 = n871 & ~n11003;
  assign n11005 = n875 & ~n11004;
  assign n11006 = n879 & ~n11005;
  assign n11007 = n883 & ~n11006;
  assign n11008 = n887 & ~n11007;
  assign n11009 = n891 & ~n11008;
  assign n11010 = n895 & ~n11009;
  assign n11011 = n899 & ~n11010;
  assign n11012 = n903 & ~n11011;
  assign n11013 = n907 & ~n11012;
  assign n11014 = n911 & ~n11013;
  assign n11015 = n915 & ~n11014;
  assign n11016 = n919 & ~n11015;
  assign n11017 = n923 & ~n11016;
  assign n11018 = n927 & ~n11017;
  assign n11019 = n931 & ~n11018;
  assign n11020 = n935 & ~n11019;
  assign n11021 = n939 & ~n11020;
  assign n11022 = n943 & ~n11021;
  assign n11023 = n947 & ~n11022;
  assign n11024 = n951 & ~n11023;
  assign n11025 = n955 & ~n11024;
  assign n11026 = n959 & ~n11025;
  assign n11027 = n963 & ~n11026;
  assign n11028 = n967 & ~n11027;
  assign n11029 = n971 & ~n11028;
  assign n11030 = n975 & ~n11029;
  assign n11031 = n979 & ~n11030;
  assign n11032 = n983 & ~n11031;
  assign n11033 = n987 & ~n11032;
  assign n11034 = n991 & ~n11033;
  assign n11035 = n995 & ~n11034;
  assign n11036 = n999 & ~n11035;
  assign n11037 = n1003 & ~n11036;
  assign n11038 = n1007 & ~n11037;
  assign n11039 = n1011 & ~n11038;
  assign n11040 = n1015 & ~n11039;
  assign n11041 = n1019 & ~n11040;
  assign n11042 = pi242  & ~n1021;
  assign po114  = ~n11041 & n11042;
  assign n11044 = n1030 & ~n1363;
  assign n11045 = n1035 & ~n11044;
  assign n11046 = n1039 & ~n11045;
  assign n11047 = n1043 & ~n11046;
  assign n11048 = n1047 & ~n11047;
  assign n11049 = n1051 & ~n11048;
  assign n11050 = n1055 & ~n11049;
  assign n11051 = n1059 & ~n11050;
  assign n11052 = n1574 & ~n11051;
  assign n11053 = n1576 & ~n11052;
  assign n11054 = n1837 & ~n11053;
  assign n11055 = n1068 & ~n11054;
  assign n11056 = n1072 & ~n11055;
  assign n11057 = n1076 & ~n11056;
  assign n11058 = n1080 & ~n11057;
  assign n11059 = n1084 & ~n11058;
  assign n11060 = n1088 & ~n11059;
  assign n11061 = n1092 & ~n11060;
  assign n11062 = n1096 & ~n11061;
  assign n11063 = n1100 & ~n11062;
  assign n11064 = n1104 & ~n11063;
  assign n11065 = n1108 & ~n11064;
  assign n11066 = n1112 & ~n11065;
  assign n11067 = n1116 & ~n11066;
  assign n11068 = n1120 & ~n11067;
  assign n11069 = n1124 & ~n11068;
  assign n11070 = n1128 & ~n11069;
  assign n11071 = n1132 & ~n11070;
  assign n11072 = n1136 & ~n11071;
  assign n11073 = n1140 & ~n11072;
  assign n11074 = n1144 & ~n11073;
  assign n11075 = n1148 & ~n11074;
  assign n11076 = n1152 & ~n11075;
  assign n11077 = n1156 & ~n11076;
  assign n11078 = n1160 & ~n11077;
  assign n11079 = n1164 & ~n11078;
  assign n11080 = n1168 & ~n11079;
  assign n11081 = n1172 & ~n11080;
  assign n11082 = n1176 & ~n11081;
  assign n11083 = n1180 & ~n11082;
  assign n11084 = n1184 & ~n11083;
  assign n11085 = n1188 & ~n11084;
  assign n11086 = n1192 & ~n11085;
  assign n11087 = n1196 & ~n11086;
  assign n11088 = n1200 & ~n11087;
  assign n11089 = n1204 & ~n11088;
  assign n11090 = n1208 & ~n11089;
  assign n11091 = n1212 & ~n11090;
  assign n11092 = n1216 & ~n11091;
  assign n11093 = n1220 & ~n11092;
  assign n11094 = n1224 & ~n11093;
  assign n11095 = n1228 & ~n11094;
  assign n11096 = n1232 & ~n11095;
  assign n11097 = n1236 & ~n11096;
  assign n11098 = n1240 & ~n11097;
  assign n11099 = n1244 & ~n11098;
  assign n11100 = n1248 & ~n11099;
  assign n11101 = n1252 & ~n11100;
  assign n11102 = n1256 & ~n11101;
  assign n11103 = n1260 & ~n11102;
  assign n11104 = n1264 & ~n11103;
  assign n11105 = n1268 & ~n11104;
  assign n11106 = n1272 & ~n11105;
  assign n11107 = n1276 & ~n11106;
  assign n11108 = n1280 & ~n11107;
  assign n11109 = n1284 & ~n11108;
  assign n11110 = n1288 & ~n11109;
  assign n11111 = n1292 & ~n11110;
  assign n11112 = n1296 & ~n11111;
  assign n11113 = n1300 & ~n11112;
  assign n11114 = n1304 & ~n11113;
  assign n11115 = n1308 & ~n11114;
  assign n11116 = n1312 & ~n11115;
  assign n11117 = n1316 & ~n11116;
  assign n11118 = n1320 & ~n11117;
  assign n11119 = n1324 & ~n11118;
  assign n11120 = n1328 & ~n11119;
  assign n11121 = n1332 & ~n11120;
  assign n11122 = n1336 & ~n11121;
  assign n11123 = n1340 & ~n11122;
  assign n11124 = n1344 & ~n11123;
  assign n11125 = n1348 & ~n11124;
  assign n11126 = n1352 & ~n11125;
  assign n11127 = n1356 & ~n11126;
  assign n11128 = pi243  & ~n1358;
  assign po115  = ~n11127 & n11128;
  assign n11130 = ~n695 & n1367;
  assign n11131 = n1372 & ~n11130;
  assign n11132 = n1376 & ~n11131;
  assign n11133 = n1380 & ~n11132;
  assign n11134 = n1384 & ~n11133;
  assign n11135 = n1388 & ~n11134;
  assign n11136 = n1392 & ~n11135;
  assign n11137 = n1396 & ~n11136;
  assign n11138 = n1663 & ~n11137;
  assign n11139 = n392 & ~n11138;
  assign n11140 = n396 & ~n11139;
  assign n11141 = n400 & ~n11140;
  assign n11142 = n404 & ~n11141;
  assign n11143 = n408 & ~n11142;
  assign n11144 = n412 & ~n11143;
  assign n11145 = n416 & ~n11144;
  assign n11146 = n420 & ~n11145;
  assign n11147 = n424 & ~n11146;
  assign n11148 = n428 & ~n11147;
  assign n11149 = n432 & ~n11148;
  assign n11150 = n436 & ~n11149;
  assign n11151 = n440 & ~n11150;
  assign n11152 = n444 & ~n11151;
  assign n11153 = n448 & ~n11152;
  assign n11154 = n452 & ~n11153;
  assign n11155 = n456 & ~n11154;
  assign n11156 = n460 & ~n11155;
  assign n11157 = n464 & ~n11156;
  assign n11158 = n468 & ~n11157;
  assign n11159 = n472 & ~n11158;
  assign n11160 = n476 & ~n11159;
  assign n11161 = n480 & ~n11160;
  assign n11162 = n484 & ~n11161;
  assign n11163 = n488 & ~n11162;
  assign n11164 = n492 & ~n11163;
  assign n11165 = n496 & ~n11164;
  assign n11166 = n500 & ~n11165;
  assign n11167 = n504 & ~n11166;
  assign n11168 = n508 & ~n11167;
  assign n11169 = n512 & ~n11168;
  assign n11170 = n516 & ~n11169;
  assign n11171 = n520 & ~n11170;
  assign n11172 = n524 & ~n11171;
  assign n11173 = n528 & ~n11172;
  assign n11174 = n532 & ~n11173;
  assign n11175 = n536 & ~n11174;
  assign n11176 = n540 & ~n11175;
  assign n11177 = n544 & ~n11176;
  assign n11178 = n548 & ~n11177;
  assign n11179 = n552 & ~n11178;
  assign n11180 = n556 & ~n11179;
  assign n11181 = n560 & ~n11180;
  assign n11182 = n564 & ~n11181;
  assign n11183 = n568 & ~n11182;
  assign n11184 = n572 & ~n11183;
  assign n11185 = n576 & ~n11184;
  assign n11186 = n580 & ~n11185;
  assign n11187 = n584 & ~n11186;
  assign n11188 = n588 & ~n11187;
  assign n11189 = n592 & ~n11188;
  assign n11190 = n596 & ~n11189;
  assign n11191 = n600 & ~n11190;
  assign n11192 = n604 & ~n11191;
  assign n11193 = n608 & ~n11192;
  assign n11194 = n612 & ~n11193;
  assign n11195 = n616 & ~n11194;
  assign n11196 = n620 & ~n11195;
  assign n11197 = n624 & ~n11196;
  assign n11198 = n628 & ~n11197;
  assign n11199 = n632 & ~n11198;
  assign n11200 = n636 & ~n11199;
  assign n11201 = n640 & ~n11200;
  assign n11202 = n644 & ~n11201;
  assign n11203 = n648 & ~n11202;
  assign n11204 = n652 & ~n11203;
  assign n11205 = n656 & ~n11204;
  assign n11206 = n660 & ~n11205;
  assign n11207 = n664 & ~n11206;
  assign n11208 = n668 & ~n11207;
  assign n11209 = n672 & ~n11208;
  assign n11210 = n676 & ~n11209;
  assign n11211 = n680 & ~n11210;
  assign n11212 = n684 & ~n11211;
  assign n11213 = n688 & ~n11212;
  assign n11214 = pi244  & ~n690;
  assign po116  = ~n11213 & n11214;
  assign n11216 = n699 & ~n1034;
  assign n11217 = n704 & ~n11216;
  assign n11218 = n708 & ~n11217;
  assign n11219 = n712 & ~n11218;
  assign n11220 = n716 & ~n11219;
  assign n11221 = n720 & ~n11220;
  assign n11222 = n1484 & ~n11221;
  assign n11223 = n1486 & ~n11222;
  assign n11224 = n1750 & ~n11223;
  assign n11225 = n731 & ~n11224;
  assign n11226 = n735 & ~n11225;
  assign n11227 = n739 & ~n11226;
  assign n11228 = n743 & ~n11227;
  assign n11229 = n747 & ~n11228;
  assign n11230 = n751 & ~n11229;
  assign n11231 = n755 & ~n11230;
  assign n11232 = n759 & ~n11231;
  assign n11233 = n763 & ~n11232;
  assign n11234 = n767 & ~n11233;
  assign n11235 = n771 & ~n11234;
  assign n11236 = n775 & ~n11235;
  assign n11237 = n779 & ~n11236;
  assign n11238 = n783 & ~n11237;
  assign n11239 = n787 & ~n11238;
  assign n11240 = n791 & ~n11239;
  assign n11241 = n795 & ~n11240;
  assign n11242 = n799 & ~n11241;
  assign n11243 = n803 & ~n11242;
  assign n11244 = n807 & ~n11243;
  assign n11245 = n811 & ~n11244;
  assign n11246 = n815 & ~n11245;
  assign n11247 = n819 & ~n11246;
  assign n11248 = n823 & ~n11247;
  assign n11249 = n827 & ~n11248;
  assign n11250 = n831 & ~n11249;
  assign n11251 = n835 & ~n11250;
  assign n11252 = n839 & ~n11251;
  assign n11253 = n843 & ~n11252;
  assign n11254 = n847 & ~n11253;
  assign n11255 = n851 & ~n11254;
  assign n11256 = n855 & ~n11255;
  assign n11257 = n859 & ~n11256;
  assign n11258 = n863 & ~n11257;
  assign n11259 = n867 & ~n11258;
  assign n11260 = n871 & ~n11259;
  assign n11261 = n875 & ~n11260;
  assign n11262 = n879 & ~n11261;
  assign n11263 = n883 & ~n11262;
  assign n11264 = n887 & ~n11263;
  assign n11265 = n891 & ~n11264;
  assign n11266 = n895 & ~n11265;
  assign n11267 = n899 & ~n11266;
  assign n11268 = n903 & ~n11267;
  assign n11269 = n907 & ~n11268;
  assign n11270 = n911 & ~n11269;
  assign n11271 = n915 & ~n11270;
  assign n11272 = n919 & ~n11271;
  assign n11273 = n923 & ~n11272;
  assign n11274 = n927 & ~n11273;
  assign n11275 = n931 & ~n11274;
  assign n11276 = n935 & ~n11275;
  assign n11277 = n939 & ~n11276;
  assign n11278 = n943 & ~n11277;
  assign n11279 = n947 & ~n11278;
  assign n11280 = n951 & ~n11279;
  assign n11281 = n955 & ~n11280;
  assign n11282 = n959 & ~n11281;
  assign n11283 = n963 & ~n11282;
  assign n11284 = n967 & ~n11283;
  assign n11285 = n971 & ~n11284;
  assign n11286 = n975 & ~n11285;
  assign n11287 = n979 & ~n11286;
  assign n11288 = n983 & ~n11287;
  assign n11289 = n987 & ~n11288;
  assign n11290 = n991 & ~n11289;
  assign n11291 = n995 & ~n11290;
  assign n11292 = n999 & ~n11291;
  assign n11293 = n1003 & ~n11292;
  assign n11294 = n1007 & ~n11293;
  assign n11295 = n1011 & ~n11294;
  assign n11296 = n1015 & ~n11295;
  assign n11297 = n1019 & ~n11296;
  assign n11298 = n1023 & ~n11297;
  assign n11299 = n1027 & ~n11298;
  assign n11300 = pi245  & ~n1029;
  assign po117  = ~n11299 & n11300;
  assign n11302 = n1038 & ~n1371;
  assign n11303 = n1043 & ~n11302;
  assign n11304 = n1047 & ~n11303;
  assign n11305 = n1051 & ~n11304;
  assign n11306 = n1055 & ~n11305;
  assign n11307 = n1059 & ~n11306;
  assign n11308 = n1574 & ~n11307;
  assign n11309 = n1576 & ~n11308;
  assign n11310 = n1837 & ~n11309;
  assign n11311 = n1068 & ~n11310;
  assign n11312 = n1072 & ~n11311;
  assign n11313 = n1076 & ~n11312;
  assign n11314 = n1080 & ~n11313;
  assign n11315 = n1084 & ~n11314;
  assign n11316 = n1088 & ~n11315;
  assign n11317 = n1092 & ~n11316;
  assign n11318 = n1096 & ~n11317;
  assign n11319 = n1100 & ~n11318;
  assign n11320 = n1104 & ~n11319;
  assign n11321 = n1108 & ~n11320;
  assign n11322 = n1112 & ~n11321;
  assign n11323 = n1116 & ~n11322;
  assign n11324 = n1120 & ~n11323;
  assign n11325 = n1124 & ~n11324;
  assign n11326 = n1128 & ~n11325;
  assign n11327 = n1132 & ~n11326;
  assign n11328 = n1136 & ~n11327;
  assign n11329 = n1140 & ~n11328;
  assign n11330 = n1144 & ~n11329;
  assign n11331 = n1148 & ~n11330;
  assign n11332 = n1152 & ~n11331;
  assign n11333 = n1156 & ~n11332;
  assign n11334 = n1160 & ~n11333;
  assign n11335 = n1164 & ~n11334;
  assign n11336 = n1168 & ~n11335;
  assign n11337 = n1172 & ~n11336;
  assign n11338 = n1176 & ~n11337;
  assign n11339 = n1180 & ~n11338;
  assign n11340 = n1184 & ~n11339;
  assign n11341 = n1188 & ~n11340;
  assign n11342 = n1192 & ~n11341;
  assign n11343 = n1196 & ~n11342;
  assign n11344 = n1200 & ~n11343;
  assign n11345 = n1204 & ~n11344;
  assign n11346 = n1208 & ~n11345;
  assign n11347 = n1212 & ~n11346;
  assign n11348 = n1216 & ~n11347;
  assign n11349 = n1220 & ~n11348;
  assign n11350 = n1224 & ~n11349;
  assign n11351 = n1228 & ~n11350;
  assign n11352 = n1232 & ~n11351;
  assign n11353 = n1236 & ~n11352;
  assign n11354 = n1240 & ~n11353;
  assign n11355 = n1244 & ~n11354;
  assign n11356 = n1248 & ~n11355;
  assign n11357 = n1252 & ~n11356;
  assign n11358 = n1256 & ~n11357;
  assign n11359 = n1260 & ~n11358;
  assign n11360 = n1264 & ~n11359;
  assign n11361 = n1268 & ~n11360;
  assign n11362 = n1272 & ~n11361;
  assign n11363 = n1276 & ~n11362;
  assign n11364 = n1280 & ~n11363;
  assign n11365 = n1284 & ~n11364;
  assign n11366 = n1288 & ~n11365;
  assign n11367 = n1292 & ~n11366;
  assign n11368 = n1296 & ~n11367;
  assign n11369 = n1300 & ~n11368;
  assign n11370 = n1304 & ~n11369;
  assign n11371 = n1308 & ~n11370;
  assign n11372 = n1312 & ~n11371;
  assign n11373 = n1316 & ~n11372;
  assign n11374 = n1320 & ~n11373;
  assign n11375 = n1324 & ~n11374;
  assign n11376 = n1328 & ~n11375;
  assign n11377 = n1332 & ~n11376;
  assign n11378 = n1336 & ~n11377;
  assign n11379 = n1340 & ~n11378;
  assign n11380 = n1344 & ~n11379;
  assign n11381 = n1348 & ~n11380;
  assign n11382 = n1352 & ~n11381;
  assign n11383 = n1356 & ~n11382;
  assign n11384 = n1360 & ~n11383;
  assign n11385 = n1364 & ~n11384;
  assign n11386 = pi246  & ~n1366;
  assign po118  = ~n11385 & n11386;
  assign n11388 = ~n703 & n1375;
  assign n11389 = n1380 & ~n11388;
  assign n11390 = n1384 & ~n11389;
  assign n11391 = n1388 & ~n11390;
  assign n11392 = n1392 & ~n11391;
  assign n11393 = n1396 & ~n11392;
  assign n11394 = n1663 & ~n11393;
  assign n11395 = n392 & ~n11394;
  assign n11396 = n396 & ~n11395;
  assign n11397 = n400 & ~n11396;
  assign n11398 = n404 & ~n11397;
  assign n11399 = n408 & ~n11398;
  assign n11400 = n412 & ~n11399;
  assign n11401 = n416 & ~n11400;
  assign n11402 = n420 & ~n11401;
  assign n11403 = n424 & ~n11402;
  assign n11404 = n428 & ~n11403;
  assign n11405 = n432 & ~n11404;
  assign n11406 = n436 & ~n11405;
  assign n11407 = n440 & ~n11406;
  assign n11408 = n444 & ~n11407;
  assign n11409 = n448 & ~n11408;
  assign n11410 = n452 & ~n11409;
  assign n11411 = n456 & ~n11410;
  assign n11412 = n460 & ~n11411;
  assign n11413 = n464 & ~n11412;
  assign n11414 = n468 & ~n11413;
  assign n11415 = n472 & ~n11414;
  assign n11416 = n476 & ~n11415;
  assign n11417 = n480 & ~n11416;
  assign n11418 = n484 & ~n11417;
  assign n11419 = n488 & ~n11418;
  assign n11420 = n492 & ~n11419;
  assign n11421 = n496 & ~n11420;
  assign n11422 = n500 & ~n11421;
  assign n11423 = n504 & ~n11422;
  assign n11424 = n508 & ~n11423;
  assign n11425 = n512 & ~n11424;
  assign n11426 = n516 & ~n11425;
  assign n11427 = n520 & ~n11426;
  assign n11428 = n524 & ~n11427;
  assign n11429 = n528 & ~n11428;
  assign n11430 = n532 & ~n11429;
  assign n11431 = n536 & ~n11430;
  assign n11432 = n540 & ~n11431;
  assign n11433 = n544 & ~n11432;
  assign n11434 = n548 & ~n11433;
  assign n11435 = n552 & ~n11434;
  assign n11436 = n556 & ~n11435;
  assign n11437 = n560 & ~n11436;
  assign n11438 = n564 & ~n11437;
  assign n11439 = n568 & ~n11438;
  assign n11440 = n572 & ~n11439;
  assign n11441 = n576 & ~n11440;
  assign n11442 = n580 & ~n11441;
  assign n11443 = n584 & ~n11442;
  assign n11444 = n588 & ~n11443;
  assign n11445 = n592 & ~n11444;
  assign n11446 = n596 & ~n11445;
  assign n11447 = n600 & ~n11446;
  assign n11448 = n604 & ~n11447;
  assign n11449 = n608 & ~n11448;
  assign n11450 = n612 & ~n11449;
  assign n11451 = n616 & ~n11450;
  assign n11452 = n620 & ~n11451;
  assign n11453 = n624 & ~n11452;
  assign n11454 = n628 & ~n11453;
  assign n11455 = n632 & ~n11454;
  assign n11456 = n636 & ~n11455;
  assign n11457 = n640 & ~n11456;
  assign n11458 = n644 & ~n11457;
  assign n11459 = n648 & ~n11458;
  assign n11460 = n652 & ~n11459;
  assign n11461 = n656 & ~n11460;
  assign n11462 = n660 & ~n11461;
  assign n11463 = n664 & ~n11462;
  assign n11464 = n668 & ~n11463;
  assign n11465 = n672 & ~n11464;
  assign n11466 = n676 & ~n11465;
  assign n11467 = n680 & ~n11466;
  assign n11468 = n684 & ~n11467;
  assign n11469 = n688 & ~n11468;
  assign n11470 = n692 & ~n11469;
  assign n11471 = n696 & ~n11470;
  assign n11472 = pi247  & ~n698;
  assign po119  = ~n11471 & n11472;
  assign n11474 = n707 & ~n1042;
  assign n11475 = n712 & ~n11474;
  assign n11476 = n716 & ~n11475;
  assign n11477 = n720 & ~n11476;
  assign n11478 = n1484 & ~n11477;
  assign n11479 = n1486 & ~n11478;
  assign n11480 = n1750 & ~n11479;
  assign n11481 = n731 & ~n11480;
  assign n11482 = n735 & ~n11481;
  assign n11483 = n739 & ~n11482;
  assign n11484 = n743 & ~n11483;
  assign n11485 = n747 & ~n11484;
  assign n11486 = n751 & ~n11485;
  assign n11487 = n755 & ~n11486;
  assign n11488 = n759 & ~n11487;
  assign n11489 = n763 & ~n11488;
  assign n11490 = n767 & ~n11489;
  assign n11491 = n771 & ~n11490;
  assign n11492 = n775 & ~n11491;
  assign n11493 = n779 & ~n11492;
  assign n11494 = n783 & ~n11493;
  assign n11495 = n787 & ~n11494;
  assign n11496 = n791 & ~n11495;
  assign n11497 = n795 & ~n11496;
  assign n11498 = n799 & ~n11497;
  assign n11499 = n803 & ~n11498;
  assign n11500 = n807 & ~n11499;
  assign n11501 = n811 & ~n11500;
  assign n11502 = n815 & ~n11501;
  assign n11503 = n819 & ~n11502;
  assign n11504 = n823 & ~n11503;
  assign n11505 = n827 & ~n11504;
  assign n11506 = n831 & ~n11505;
  assign n11507 = n835 & ~n11506;
  assign n11508 = n839 & ~n11507;
  assign n11509 = n843 & ~n11508;
  assign n11510 = n847 & ~n11509;
  assign n11511 = n851 & ~n11510;
  assign n11512 = n855 & ~n11511;
  assign n11513 = n859 & ~n11512;
  assign n11514 = n863 & ~n11513;
  assign n11515 = n867 & ~n11514;
  assign n11516 = n871 & ~n11515;
  assign n11517 = n875 & ~n11516;
  assign n11518 = n879 & ~n11517;
  assign n11519 = n883 & ~n11518;
  assign n11520 = n887 & ~n11519;
  assign n11521 = n891 & ~n11520;
  assign n11522 = n895 & ~n11521;
  assign n11523 = n899 & ~n11522;
  assign n11524 = n903 & ~n11523;
  assign n11525 = n907 & ~n11524;
  assign n11526 = n911 & ~n11525;
  assign n11527 = n915 & ~n11526;
  assign n11528 = n919 & ~n11527;
  assign n11529 = n923 & ~n11528;
  assign n11530 = n927 & ~n11529;
  assign n11531 = n931 & ~n11530;
  assign n11532 = n935 & ~n11531;
  assign n11533 = n939 & ~n11532;
  assign n11534 = n943 & ~n11533;
  assign n11535 = n947 & ~n11534;
  assign n11536 = n951 & ~n11535;
  assign n11537 = n955 & ~n11536;
  assign n11538 = n959 & ~n11537;
  assign n11539 = n963 & ~n11538;
  assign n11540 = n967 & ~n11539;
  assign n11541 = n971 & ~n11540;
  assign n11542 = n975 & ~n11541;
  assign n11543 = n979 & ~n11542;
  assign n11544 = n983 & ~n11543;
  assign n11545 = n987 & ~n11544;
  assign n11546 = n991 & ~n11545;
  assign n11547 = n995 & ~n11546;
  assign n11548 = n999 & ~n11547;
  assign n11549 = n1003 & ~n11548;
  assign n11550 = n1007 & ~n11549;
  assign n11551 = n1011 & ~n11550;
  assign n11552 = n1015 & ~n11551;
  assign n11553 = n1019 & ~n11552;
  assign n11554 = n1023 & ~n11553;
  assign n11555 = n1027 & ~n11554;
  assign n11556 = n1031 & ~n11555;
  assign n11557 = n1035 & ~n11556;
  assign n11558 = pi248  & ~n1037;
  assign po120  = ~n11557 & n11558;
  assign n11560 = n1046 & ~n1379;
  assign n11561 = n1051 & ~n11560;
  assign n11562 = n1055 & ~n11561;
  assign n11563 = n1059 & ~n11562;
  assign n11564 = n1574 & ~n11563;
  assign n11565 = n1576 & ~n11564;
  assign n11566 = n1837 & ~n11565;
  assign n11567 = n1068 & ~n11566;
  assign n11568 = n1072 & ~n11567;
  assign n11569 = n1076 & ~n11568;
  assign n11570 = n1080 & ~n11569;
  assign n11571 = n1084 & ~n11570;
  assign n11572 = n1088 & ~n11571;
  assign n11573 = n1092 & ~n11572;
  assign n11574 = n1096 & ~n11573;
  assign n11575 = n1100 & ~n11574;
  assign n11576 = n1104 & ~n11575;
  assign n11577 = n1108 & ~n11576;
  assign n11578 = n1112 & ~n11577;
  assign n11579 = n1116 & ~n11578;
  assign n11580 = n1120 & ~n11579;
  assign n11581 = n1124 & ~n11580;
  assign n11582 = n1128 & ~n11581;
  assign n11583 = n1132 & ~n11582;
  assign n11584 = n1136 & ~n11583;
  assign n11585 = n1140 & ~n11584;
  assign n11586 = n1144 & ~n11585;
  assign n11587 = n1148 & ~n11586;
  assign n11588 = n1152 & ~n11587;
  assign n11589 = n1156 & ~n11588;
  assign n11590 = n1160 & ~n11589;
  assign n11591 = n1164 & ~n11590;
  assign n11592 = n1168 & ~n11591;
  assign n11593 = n1172 & ~n11592;
  assign n11594 = n1176 & ~n11593;
  assign n11595 = n1180 & ~n11594;
  assign n11596 = n1184 & ~n11595;
  assign n11597 = n1188 & ~n11596;
  assign n11598 = n1192 & ~n11597;
  assign n11599 = n1196 & ~n11598;
  assign n11600 = n1200 & ~n11599;
  assign n11601 = n1204 & ~n11600;
  assign n11602 = n1208 & ~n11601;
  assign n11603 = n1212 & ~n11602;
  assign n11604 = n1216 & ~n11603;
  assign n11605 = n1220 & ~n11604;
  assign n11606 = n1224 & ~n11605;
  assign n11607 = n1228 & ~n11606;
  assign n11608 = n1232 & ~n11607;
  assign n11609 = n1236 & ~n11608;
  assign n11610 = n1240 & ~n11609;
  assign n11611 = n1244 & ~n11610;
  assign n11612 = n1248 & ~n11611;
  assign n11613 = n1252 & ~n11612;
  assign n11614 = n1256 & ~n11613;
  assign n11615 = n1260 & ~n11614;
  assign n11616 = n1264 & ~n11615;
  assign n11617 = n1268 & ~n11616;
  assign n11618 = n1272 & ~n11617;
  assign n11619 = n1276 & ~n11618;
  assign n11620 = n1280 & ~n11619;
  assign n11621 = n1284 & ~n11620;
  assign n11622 = n1288 & ~n11621;
  assign n11623 = n1292 & ~n11622;
  assign n11624 = n1296 & ~n11623;
  assign n11625 = n1300 & ~n11624;
  assign n11626 = n1304 & ~n11625;
  assign n11627 = n1308 & ~n11626;
  assign n11628 = n1312 & ~n11627;
  assign n11629 = n1316 & ~n11628;
  assign n11630 = n1320 & ~n11629;
  assign n11631 = n1324 & ~n11630;
  assign n11632 = n1328 & ~n11631;
  assign n11633 = n1332 & ~n11632;
  assign n11634 = n1336 & ~n11633;
  assign n11635 = n1340 & ~n11634;
  assign n11636 = n1344 & ~n11635;
  assign n11637 = n1348 & ~n11636;
  assign n11638 = n1352 & ~n11637;
  assign n11639 = n1356 & ~n11638;
  assign n11640 = n1360 & ~n11639;
  assign n11641 = n1364 & ~n11640;
  assign n11642 = n1368 & ~n11641;
  assign n11643 = n1372 & ~n11642;
  assign n11644 = pi249  & ~n1374;
  assign po121  = ~n11643 & n11644;
  assign n11646 = ~n711 & n1383;
  assign n11647 = n1388 & ~n11646;
  assign n11648 = n1392 & ~n11647;
  assign n11649 = n1396 & ~n11648;
  assign n11650 = n1663 & ~n11649;
  assign n11651 = n392 & ~n11650;
  assign n11652 = n396 & ~n11651;
  assign n11653 = n400 & ~n11652;
  assign n11654 = n404 & ~n11653;
  assign n11655 = n408 & ~n11654;
  assign n11656 = n412 & ~n11655;
  assign n11657 = n416 & ~n11656;
  assign n11658 = n420 & ~n11657;
  assign n11659 = n424 & ~n11658;
  assign n11660 = n428 & ~n11659;
  assign n11661 = n432 & ~n11660;
  assign n11662 = n436 & ~n11661;
  assign n11663 = n440 & ~n11662;
  assign n11664 = n444 & ~n11663;
  assign n11665 = n448 & ~n11664;
  assign n11666 = n452 & ~n11665;
  assign n11667 = n456 & ~n11666;
  assign n11668 = n460 & ~n11667;
  assign n11669 = n464 & ~n11668;
  assign n11670 = n468 & ~n11669;
  assign n11671 = n472 & ~n11670;
  assign n11672 = n476 & ~n11671;
  assign n11673 = n480 & ~n11672;
  assign n11674 = n484 & ~n11673;
  assign n11675 = n488 & ~n11674;
  assign n11676 = n492 & ~n11675;
  assign n11677 = n496 & ~n11676;
  assign n11678 = n500 & ~n11677;
  assign n11679 = n504 & ~n11678;
  assign n11680 = n508 & ~n11679;
  assign n11681 = n512 & ~n11680;
  assign n11682 = n516 & ~n11681;
  assign n11683 = n520 & ~n11682;
  assign n11684 = n524 & ~n11683;
  assign n11685 = n528 & ~n11684;
  assign n11686 = n532 & ~n11685;
  assign n11687 = n536 & ~n11686;
  assign n11688 = n540 & ~n11687;
  assign n11689 = n544 & ~n11688;
  assign n11690 = n548 & ~n11689;
  assign n11691 = n552 & ~n11690;
  assign n11692 = n556 & ~n11691;
  assign n11693 = n560 & ~n11692;
  assign n11694 = n564 & ~n11693;
  assign n11695 = n568 & ~n11694;
  assign n11696 = n572 & ~n11695;
  assign n11697 = n576 & ~n11696;
  assign n11698 = n580 & ~n11697;
  assign n11699 = n584 & ~n11698;
  assign n11700 = n588 & ~n11699;
  assign n11701 = n592 & ~n11700;
  assign n11702 = n596 & ~n11701;
  assign n11703 = n600 & ~n11702;
  assign n11704 = n604 & ~n11703;
  assign n11705 = n608 & ~n11704;
  assign n11706 = n612 & ~n11705;
  assign n11707 = n616 & ~n11706;
  assign n11708 = n620 & ~n11707;
  assign n11709 = n624 & ~n11708;
  assign n11710 = n628 & ~n11709;
  assign n11711 = n632 & ~n11710;
  assign n11712 = n636 & ~n11711;
  assign n11713 = n640 & ~n11712;
  assign n11714 = n644 & ~n11713;
  assign n11715 = n648 & ~n11714;
  assign n11716 = n652 & ~n11715;
  assign n11717 = n656 & ~n11716;
  assign n11718 = n660 & ~n11717;
  assign n11719 = n664 & ~n11718;
  assign n11720 = n668 & ~n11719;
  assign n11721 = n672 & ~n11720;
  assign n11722 = n676 & ~n11721;
  assign n11723 = n680 & ~n11722;
  assign n11724 = n684 & ~n11723;
  assign n11725 = n688 & ~n11724;
  assign n11726 = n692 & ~n11725;
  assign n11727 = n696 & ~n11726;
  assign n11728 = n700 & ~n11727;
  assign n11729 = n704 & ~n11728;
  assign n11730 = pi250  & ~n706;
  assign po122  = ~n11729 & n11730;
  assign n11732 = n715 & ~n1050;
  assign n11733 = n720 & ~n11732;
  assign n11734 = n1484 & ~n11733;
  assign n11735 = n1486 & ~n11734;
  assign n11736 = n1750 & ~n11735;
  assign n11737 = n731 & ~n11736;
  assign n11738 = n735 & ~n11737;
  assign n11739 = n739 & ~n11738;
  assign n11740 = n743 & ~n11739;
  assign n11741 = n747 & ~n11740;
  assign n11742 = n751 & ~n11741;
  assign n11743 = n755 & ~n11742;
  assign n11744 = n759 & ~n11743;
  assign n11745 = n763 & ~n11744;
  assign n11746 = n767 & ~n11745;
  assign n11747 = n771 & ~n11746;
  assign n11748 = n775 & ~n11747;
  assign n11749 = n779 & ~n11748;
  assign n11750 = n783 & ~n11749;
  assign n11751 = n787 & ~n11750;
  assign n11752 = n791 & ~n11751;
  assign n11753 = n795 & ~n11752;
  assign n11754 = n799 & ~n11753;
  assign n11755 = n803 & ~n11754;
  assign n11756 = n807 & ~n11755;
  assign n11757 = n811 & ~n11756;
  assign n11758 = n815 & ~n11757;
  assign n11759 = n819 & ~n11758;
  assign n11760 = n823 & ~n11759;
  assign n11761 = n827 & ~n11760;
  assign n11762 = n831 & ~n11761;
  assign n11763 = n835 & ~n11762;
  assign n11764 = n839 & ~n11763;
  assign n11765 = n843 & ~n11764;
  assign n11766 = n847 & ~n11765;
  assign n11767 = n851 & ~n11766;
  assign n11768 = n855 & ~n11767;
  assign n11769 = n859 & ~n11768;
  assign n11770 = n863 & ~n11769;
  assign n11771 = n867 & ~n11770;
  assign n11772 = n871 & ~n11771;
  assign n11773 = n875 & ~n11772;
  assign n11774 = n879 & ~n11773;
  assign n11775 = n883 & ~n11774;
  assign n11776 = n887 & ~n11775;
  assign n11777 = n891 & ~n11776;
  assign n11778 = n895 & ~n11777;
  assign n11779 = n899 & ~n11778;
  assign n11780 = n903 & ~n11779;
  assign n11781 = n907 & ~n11780;
  assign n11782 = n911 & ~n11781;
  assign n11783 = n915 & ~n11782;
  assign n11784 = n919 & ~n11783;
  assign n11785 = n923 & ~n11784;
  assign n11786 = n927 & ~n11785;
  assign n11787 = n931 & ~n11786;
  assign n11788 = n935 & ~n11787;
  assign n11789 = n939 & ~n11788;
  assign n11790 = n943 & ~n11789;
  assign n11791 = n947 & ~n11790;
  assign n11792 = n951 & ~n11791;
  assign n11793 = n955 & ~n11792;
  assign n11794 = n959 & ~n11793;
  assign n11795 = n963 & ~n11794;
  assign n11796 = n967 & ~n11795;
  assign n11797 = n971 & ~n11796;
  assign n11798 = n975 & ~n11797;
  assign n11799 = n979 & ~n11798;
  assign n11800 = n983 & ~n11799;
  assign n11801 = n987 & ~n11800;
  assign n11802 = n991 & ~n11801;
  assign n11803 = n995 & ~n11802;
  assign n11804 = n999 & ~n11803;
  assign n11805 = n1003 & ~n11804;
  assign n11806 = n1007 & ~n11805;
  assign n11807 = n1011 & ~n11806;
  assign n11808 = n1015 & ~n11807;
  assign n11809 = n1019 & ~n11808;
  assign n11810 = n1023 & ~n11809;
  assign n11811 = n1027 & ~n11810;
  assign n11812 = n1031 & ~n11811;
  assign n11813 = n1035 & ~n11812;
  assign n11814 = n1039 & ~n11813;
  assign n11815 = n1043 & ~n11814;
  assign n11816 = pi251  & ~n1045;
  assign po123  = ~n11815 & n11816;
  assign n11818 = n1054 & ~n1387;
  assign n11819 = n1059 & ~n11818;
  assign n11820 = n1574 & ~n11819;
  assign n11821 = n1576 & ~n11820;
  assign n11822 = n1837 & ~n11821;
  assign n11823 = n1068 & ~n11822;
  assign n11824 = n1072 & ~n11823;
  assign n11825 = n1076 & ~n11824;
  assign n11826 = n1080 & ~n11825;
  assign n11827 = n1084 & ~n11826;
  assign n11828 = n1088 & ~n11827;
  assign n11829 = n1092 & ~n11828;
  assign n11830 = n1096 & ~n11829;
  assign n11831 = n1100 & ~n11830;
  assign n11832 = n1104 & ~n11831;
  assign n11833 = n1108 & ~n11832;
  assign n11834 = n1112 & ~n11833;
  assign n11835 = n1116 & ~n11834;
  assign n11836 = n1120 & ~n11835;
  assign n11837 = n1124 & ~n11836;
  assign n11838 = n1128 & ~n11837;
  assign n11839 = n1132 & ~n11838;
  assign n11840 = n1136 & ~n11839;
  assign n11841 = n1140 & ~n11840;
  assign n11842 = n1144 & ~n11841;
  assign n11843 = n1148 & ~n11842;
  assign n11844 = n1152 & ~n11843;
  assign n11845 = n1156 & ~n11844;
  assign n11846 = n1160 & ~n11845;
  assign n11847 = n1164 & ~n11846;
  assign n11848 = n1168 & ~n11847;
  assign n11849 = n1172 & ~n11848;
  assign n11850 = n1176 & ~n11849;
  assign n11851 = n1180 & ~n11850;
  assign n11852 = n1184 & ~n11851;
  assign n11853 = n1188 & ~n11852;
  assign n11854 = n1192 & ~n11853;
  assign n11855 = n1196 & ~n11854;
  assign n11856 = n1200 & ~n11855;
  assign n11857 = n1204 & ~n11856;
  assign n11858 = n1208 & ~n11857;
  assign n11859 = n1212 & ~n11858;
  assign n11860 = n1216 & ~n11859;
  assign n11861 = n1220 & ~n11860;
  assign n11862 = n1224 & ~n11861;
  assign n11863 = n1228 & ~n11862;
  assign n11864 = n1232 & ~n11863;
  assign n11865 = n1236 & ~n11864;
  assign n11866 = n1240 & ~n11865;
  assign n11867 = n1244 & ~n11866;
  assign n11868 = n1248 & ~n11867;
  assign n11869 = n1252 & ~n11868;
  assign n11870 = n1256 & ~n11869;
  assign n11871 = n1260 & ~n11870;
  assign n11872 = n1264 & ~n11871;
  assign n11873 = n1268 & ~n11872;
  assign n11874 = n1272 & ~n11873;
  assign n11875 = n1276 & ~n11874;
  assign n11876 = n1280 & ~n11875;
  assign n11877 = n1284 & ~n11876;
  assign n11878 = n1288 & ~n11877;
  assign n11879 = n1292 & ~n11878;
  assign n11880 = n1296 & ~n11879;
  assign n11881 = n1300 & ~n11880;
  assign n11882 = n1304 & ~n11881;
  assign n11883 = n1308 & ~n11882;
  assign n11884 = n1312 & ~n11883;
  assign n11885 = n1316 & ~n11884;
  assign n11886 = n1320 & ~n11885;
  assign n11887 = n1324 & ~n11886;
  assign n11888 = n1328 & ~n11887;
  assign n11889 = n1332 & ~n11888;
  assign n11890 = n1336 & ~n11889;
  assign n11891 = n1340 & ~n11890;
  assign n11892 = n1344 & ~n11891;
  assign n11893 = n1348 & ~n11892;
  assign n11894 = n1352 & ~n11893;
  assign n11895 = n1356 & ~n11894;
  assign n11896 = n1360 & ~n11895;
  assign n11897 = n1364 & ~n11896;
  assign n11898 = n1368 & ~n11897;
  assign n11899 = n1372 & ~n11898;
  assign n11900 = n1376 & ~n11899;
  assign n11901 = n1380 & ~n11900;
  assign n11902 = pi252  & ~n1382;
  assign po124  = ~n11901 & n11902;
  assign n11904 = ~n719 & n1391;
  assign n11905 = n1396 & ~n11904;
  assign n11906 = n1663 & ~n11905;
  assign n11907 = n392 & ~n11906;
  assign n11908 = n396 & ~n11907;
  assign n11909 = n400 & ~n11908;
  assign n11910 = n404 & ~n11909;
  assign n11911 = n408 & ~n11910;
  assign n11912 = n412 & ~n11911;
  assign n11913 = n416 & ~n11912;
  assign n11914 = n420 & ~n11913;
  assign n11915 = n424 & ~n11914;
  assign n11916 = n428 & ~n11915;
  assign n11917 = n432 & ~n11916;
  assign n11918 = n436 & ~n11917;
  assign n11919 = n440 & ~n11918;
  assign n11920 = n444 & ~n11919;
  assign n11921 = n448 & ~n11920;
  assign n11922 = n452 & ~n11921;
  assign n11923 = n456 & ~n11922;
  assign n11924 = n460 & ~n11923;
  assign n11925 = n464 & ~n11924;
  assign n11926 = n468 & ~n11925;
  assign n11927 = n472 & ~n11926;
  assign n11928 = n476 & ~n11927;
  assign n11929 = n480 & ~n11928;
  assign n11930 = n484 & ~n11929;
  assign n11931 = n488 & ~n11930;
  assign n11932 = n492 & ~n11931;
  assign n11933 = n496 & ~n11932;
  assign n11934 = n500 & ~n11933;
  assign n11935 = n504 & ~n11934;
  assign n11936 = n508 & ~n11935;
  assign n11937 = n512 & ~n11936;
  assign n11938 = n516 & ~n11937;
  assign n11939 = n520 & ~n11938;
  assign n11940 = n524 & ~n11939;
  assign n11941 = n528 & ~n11940;
  assign n11942 = n532 & ~n11941;
  assign n11943 = n536 & ~n11942;
  assign n11944 = n540 & ~n11943;
  assign n11945 = n544 & ~n11944;
  assign n11946 = n548 & ~n11945;
  assign n11947 = n552 & ~n11946;
  assign n11948 = n556 & ~n11947;
  assign n11949 = n560 & ~n11948;
  assign n11950 = n564 & ~n11949;
  assign n11951 = n568 & ~n11950;
  assign n11952 = n572 & ~n11951;
  assign n11953 = n576 & ~n11952;
  assign n11954 = n580 & ~n11953;
  assign n11955 = n584 & ~n11954;
  assign n11956 = n588 & ~n11955;
  assign n11957 = n592 & ~n11956;
  assign n11958 = n596 & ~n11957;
  assign n11959 = n600 & ~n11958;
  assign n11960 = n604 & ~n11959;
  assign n11961 = n608 & ~n11960;
  assign n11962 = n612 & ~n11961;
  assign n11963 = n616 & ~n11962;
  assign n11964 = n620 & ~n11963;
  assign n11965 = n624 & ~n11964;
  assign n11966 = n628 & ~n11965;
  assign n11967 = n632 & ~n11966;
  assign n11968 = n636 & ~n11967;
  assign n11969 = n640 & ~n11968;
  assign n11970 = n644 & ~n11969;
  assign n11971 = n648 & ~n11970;
  assign n11972 = n652 & ~n11971;
  assign n11973 = n656 & ~n11972;
  assign n11974 = n660 & ~n11973;
  assign n11975 = n664 & ~n11974;
  assign n11976 = n668 & ~n11975;
  assign n11977 = n672 & ~n11976;
  assign n11978 = n676 & ~n11977;
  assign n11979 = n680 & ~n11978;
  assign n11980 = n684 & ~n11979;
  assign n11981 = n688 & ~n11980;
  assign n11982 = n692 & ~n11981;
  assign n11983 = n696 & ~n11982;
  assign n11984 = n700 & ~n11983;
  assign n11985 = n704 & ~n11984;
  assign n11986 = n708 & ~n11985;
  assign n11987 = n712 & ~n11986;
  assign n11988 = pi253  & ~n714;
  assign po125  = ~n11987 & n11988;
  assign n11990 = ~n1058 & n1483;
  assign n11991 = n1486 & ~n11990;
  assign n11992 = n1750 & ~n11991;
  assign n11993 = n731 & ~n11992;
  assign n11994 = n735 & ~n11993;
  assign n11995 = n739 & ~n11994;
  assign n11996 = n743 & ~n11995;
  assign n11997 = n747 & ~n11996;
  assign n11998 = n751 & ~n11997;
  assign n11999 = n755 & ~n11998;
  assign n12000 = n759 & ~n11999;
  assign n12001 = n763 & ~n12000;
  assign n12002 = n767 & ~n12001;
  assign n12003 = n771 & ~n12002;
  assign n12004 = n775 & ~n12003;
  assign n12005 = n779 & ~n12004;
  assign n12006 = n783 & ~n12005;
  assign n12007 = n787 & ~n12006;
  assign n12008 = n791 & ~n12007;
  assign n12009 = n795 & ~n12008;
  assign n12010 = n799 & ~n12009;
  assign n12011 = n803 & ~n12010;
  assign n12012 = n807 & ~n12011;
  assign n12013 = n811 & ~n12012;
  assign n12014 = n815 & ~n12013;
  assign n12015 = n819 & ~n12014;
  assign n12016 = n823 & ~n12015;
  assign n12017 = n827 & ~n12016;
  assign n12018 = n831 & ~n12017;
  assign n12019 = n835 & ~n12018;
  assign n12020 = n839 & ~n12019;
  assign n12021 = n843 & ~n12020;
  assign n12022 = n847 & ~n12021;
  assign n12023 = n851 & ~n12022;
  assign n12024 = n855 & ~n12023;
  assign n12025 = n859 & ~n12024;
  assign n12026 = n863 & ~n12025;
  assign n12027 = n867 & ~n12026;
  assign n12028 = n871 & ~n12027;
  assign n12029 = n875 & ~n12028;
  assign n12030 = n879 & ~n12029;
  assign n12031 = n883 & ~n12030;
  assign n12032 = n887 & ~n12031;
  assign n12033 = n891 & ~n12032;
  assign n12034 = n895 & ~n12033;
  assign n12035 = n899 & ~n12034;
  assign n12036 = n903 & ~n12035;
  assign n12037 = n907 & ~n12036;
  assign n12038 = n911 & ~n12037;
  assign n12039 = n915 & ~n12038;
  assign n12040 = n919 & ~n12039;
  assign n12041 = n923 & ~n12040;
  assign n12042 = n927 & ~n12041;
  assign n12043 = n931 & ~n12042;
  assign n12044 = n935 & ~n12043;
  assign n12045 = n939 & ~n12044;
  assign n12046 = n943 & ~n12045;
  assign n12047 = n947 & ~n12046;
  assign n12048 = n951 & ~n12047;
  assign n12049 = n955 & ~n12048;
  assign n12050 = n959 & ~n12049;
  assign n12051 = n963 & ~n12050;
  assign n12052 = n967 & ~n12051;
  assign n12053 = n971 & ~n12052;
  assign n12054 = n975 & ~n12053;
  assign n12055 = n979 & ~n12054;
  assign n12056 = n983 & ~n12055;
  assign n12057 = n987 & ~n12056;
  assign n12058 = n991 & ~n12057;
  assign n12059 = n995 & ~n12058;
  assign n12060 = n999 & ~n12059;
  assign n12061 = n1003 & ~n12060;
  assign n12062 = n1007 & ~n12061;
  assign n12063 = n1011 & ~n12062;
  assign n12064 = n1015 & ~n12063;
  assign n12065 = n1019 & ~n12064;
  assign n12066 = n1023 & ~n12065;
  assign n12067 = n1027 & ~n12066;
  assign n12068 = n1031 & ~n12067;
  assign n12069 = n1035 & ~n12068;
  assign n12070 = n1039 & ~n12069;
  assign n12071 = n1043 & ~n12070;
  assign n12072 = n1047 & ~n12071;
  assign n12073 = n1051 & ~n12072;
  assign n12074 = pi254  & ~n1053;
  assign po126  = ~n12073 & n12074;
  assign n12076 = ~n1395 & n1573;
  assign n12077 = n1576 & ~n12076;
  assign n12078 = n1837 & ~n12077;
  assign n12079 = n1068 & ~n12078;
  assign n12080 = n1072 & ~n12079;
  assign n12081 = n1076 & ~n12080;
  assign n12082 = n1080 & ~n12081;
  assign n12083 = n1084 & ~n12082;
  assign n12084 = n1088 & ~n12083;
  assign n12085 = n1092 & ~n12084;
  assign n12086 = n1096 & ~n12085;
  assign n12087 = n1100 & ~n12086;
  assign n12088 = n1104 & ~n12087;
  assign n12089 = n1108 & ~n12088;
  assign n12090 = n1112 & ~n12089;
  assign n12091 = n1116 & ~n12090;
  assign n12092 = n1120 & ~n12091;
  assign n12093 = n1124 & ~n12092;
  assign n12094 = n1128 & ~n12093;
  assign n12095 = n1132 & ~n12094;
  assign n12096 = n1136 & ~n12095;
  assign n12097 = n1140 & ~n12096;
  assign n12098 = n1144 & ~n12097;
  assign n12099 = n1148 & ~n12098;
  assign n12100 = n1152 & ~n12099;
  assign n12101 = n1156 & ~n12100;
  assign n12102 = n1160 & ~n12101;
  assign n12103 = n1164 & ~n12102;
  assign n12104 = n1168 & ~n12103;
  assign n12105 = n1172 & ~n12104;
  assign n12106 = n1176 & ~n12105;
  assign n12107 = n1180 & ~n12106;
  assign n12108 = n1184 & ~n12107;
  assign n12109 = n1188 & ~n12108;
  assign n12110 = n1192 & ~n12109;
  assign n12111 = n1196 & ~n12110;
  assign n12112 = n1200 & ~n12111;
  assign n12113 = n1204 & ~n12112;
  assign n12114 = n1208 & ~n12113;
  assign n12115 = n1212 & ~n12114;
  assign n12116 = n1216 & ~n12115;
  assign n12117 = n1220 & ~n12116;
  assign n12118 = n1224 & ~n12117;
  assign n12119 = n1228 & ~n12118;
  assign n12120 = n1232 & ~n12119;
  assign n12121 = n1236 & ~n12120;
  assign n12122 = n1240 & ~n12121;
  assign n12123 = n1244 & ~n12122;
  assign n12124 = n1248 & ~n12123;
  assign n12125 = n1252 & ~n12124;
  assign n12126 = n1256 & ~n12125;
  assign n12127 = n1260 & ~n12126;
  assign n12128 = n1264 & ~n12127;
  assign n12129 = n1268 & ~n12128;
  assign n12130 = n1272 & ~n12129;
  assign n12131 = n1276 & ~n12130;
  assign n12132 = n1280 & ~n12131;
  assign n12133 = n1284 & ~n12132;
  assign n12134 = n1288 & ~n12133;
  assign n12135 = n1292 & ~n12134;
  assign n12136 = n1296 & ~n12135;
  assign n12137 = n1300 & ~n12136;
  assign n12138 = n1304 & ~n12137;
  assign n12139 = n1308 & ~n12138;
  assign n12140 = n1312 & ~n12139;
  assign n12141 = n1316 & ~n12140;
  assign n12142 = n1320 & ~n12141;
  assign n12143 = n1324 & ~n12142;
  assign n12144 = n1328 & ~n12143;
  assign n12145 = n1332 & ~n12144;
  assign n12146 = n1336 & ~n12145;
  assign n12147 = n1340 & ~n12146;
  assign n12148 = n1344 & ~n12147;
  assign n12149 = n1348 & ~n12148;
  assign n12150 = n1352 & ~n12149;
  assign n12151 = n1356 & ~n12150;
  assign n12152 = n1360 & ~n12151;
  assign n12153 = n1364 & ~n12152;
  assign n12154 = n1368 & ~n12153;
  assign n12155 = n1372 & ~n12154;
  assign n12156 = n1376 & ~n12155;
  assign n12157 = n1380 & ~n12156;
  assign n12158 = n1384 & ~n12157;
  assign n12159 = n1388 & ~n12158;
  assign n12160 = pi255  & ~n1390;
  assign po127  = ~n12159 & n12160;
  assign n12162 = n862 & n878;
  assign n12163 = n846 & n894;
  assign n12164 = n814 & n12163;
  assign n12165 = n12162 & n12164;
  assign n12166 = n782 & n12165;
  assign n12167 = n798 & n12166;
  assign n12168 = n734 & n750;
  assign n12169 = n707 & n766;
  assign n12170 = n675 & n12169;
  assign n12171 = n12168 & n12170;
  assign n12172 = n643 & n12171;
  assign n12173 = n659 & n691;
  assign n12174 = n12172 & n12173;
  assign n12175 = n830 & n12174;
  assign n12176 = n12167 & n12175;
  assign n12177 = n595 & n611;
  assign n12178 = n579 & n627;
  assign n12179 = n547 & n12178;
  assign n12180 = n12177 & n12179;
  assign n12181 = n515 & n12180;
  assign n12182 = n531 & n12181;
  assign n12183 = n467 & n483;
  assign n12184 = n451 & n499;
  assign n12185 = n419 & n12184;
  assign n12186 = n12183 & n12185;
  assign n12187 = n388 & n12186;
  assign n12188 = n403 & n435;
  assign n12189 = n12187 & n12188;
  assign n12190 = n563 & n12189;
  assign n12191 = n12182 & n12190;
  assign n12192 = n12176 & n12191;
  assign n12193 = n1367 & n1383;
  assign n12194 = n1351 & n1483;
  assign n12195 = n1319 & n12194;
  assign n12196 = n12193 & n12195;
  assign n12197 = n1287 & n12196;
  assign n12198 = n1303 & n12197;
  assign n12199 = n1239 & n1255;
  assign n12200 = n1223 & n1271;
  assign n12201 = n1191 & n12200;
  assign n12202 = n12199 & n12201;
  assign n12203 = n1159 & n12202;
  assign n12204 = n1175 & n1207;
  assign n12205 = n12203 & n12204;
  assign n12206 = n1335 & n12205;
  assign n12207 = n12198 & n12206;
  assign n12208 = n1111 & n1127;
  assign n12209 = n1095 & n1143;
  assign n12210 = n1064 & n12209;
  assign n12211 = n12208 & n12210;
  assign n12212 = n1038 & n12211;
  assign n12213 = n1054 & n12212;
  assign n12214 = n990 & n1006;
  assign n12215 = n974 & n1022;
  assign n12216 = n942 & n12215;
  assign n12217 = n12214 & n12216;
  assign n12218 = n910 & n12217;
  assign n12219 = n926 & n958;
  assign n12220 = n12218 & n12219;
  assign n12221 = n1079 & n12220;
  assign n12222 = n12213 & n12221;
  assign n12223 = n12207 & n12222;
  assign po128 = ~n12192 | ~n12223;
endmodule
