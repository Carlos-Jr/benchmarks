module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 ,
    po6 , po7 , po8 , po9 , po10 ,
    po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 ,
    po21 , po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 , po30 ,
    po31 , po32 , po33 , po34 , po35 ,
    po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 ,
    po46 , po47 , po48 , po49 , po50 ,
    po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 ,
    po61 , po62 , po63   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 ;
  wire n194, n195, n196, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n245,
    n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366,
    n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408,
    n409, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486,
    n487, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n677, n678,
    n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847,
    n848, n849, n850, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n861,
    n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889,
    n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903,
    n904, n905, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925,
    n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988,
    n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201,
    n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231,
    n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291,
    n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321,
    n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672,
    n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702,
    n1703, n1704, n1705, n1706, n1707, n1708,
    n1709, n1710, n1711, n1712, n1713, n1714,
    n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726,
    n1727, n1728, n1729, n1730, n1731, n1732,
    n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1740, n1741, n1742, n1743, n1744,
    n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756,
    n1757, n1758, n1759, n1760, n1761, n1762,
    n1763, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774,
    n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786,
    n1787, n1788, n1789, n1790, n1791, n1792,
    n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816,
    n1817, n1818, n1819, n1820, n1821, n1822,
    n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834,
    n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1849, n1850, n1851, n1852, n1853,
    n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871,
    n1872, n1873, n1874, n1875, n1876, n1877,
    n1878, n1879, n1880, n1881, n1882, n1883,
    n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901,
    n1902, n1903, n1904, n1905, n1906, n1907,
    n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931,
    n1932, n1933, n1934, n1935, n1936, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1959, n1960, n1961,
    n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973,
    n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991,
    n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003,
    n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2017, n2018, n2019, n2020, n2021,
    n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2029, n2030, n2031, n2032, n2033,
    n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2043, n2044, n2045, n2046,
    n2047, n2048, n2049, n2050, n2051, n2052,
    n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076,
    n2077, n2078, n2079, n2080, n2081, n2082,
    n2083, n2084, n2085, n2086, n2087, n2088,
    n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106,
    n2107, n2108, n2109, n2110, n2111, n2112,
    n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142,
    n2143, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202,
    n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232,
    n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2244,
    n2245, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281,
    n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311,
    n2312, n2313, n2314, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2323,
    n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341,
    n2342, n2343, n2344, n2345, n2346, n2347,
    n2348, n2349, n2350, n2351, n2352, n2353,
    n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371,
    n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401,
    n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2923, n2924, n2925, n2926,
    n2927, n2928, n2929, n2930, n2931, n2932,
    n2933, n2934, n2935, n2936, n2937, n2938,
    n2939, n2940, n2941, n2942, n2943, n2944,
    n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956,
    n2957, n2958, n2959, n2960, n2961, n2962,
    n2963, n2964, n2965, n2966, n2967, n2968,
    n2969, n2970, n2971, n2972, n2973, n2974,
    n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986,
    n2987, n2988, n2989, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2997, n2998,
    n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016,
    n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3025, n3026, n3027, n3028,
    n3029, n3030, n3031, n3032, n3033, n3034,
    n3035, n3036, n3037, n3038, n3039, n3040,
    n3041, n3042, n3043, n3044, n3045, n3046,
    n3047, n3048, n3049, n3050, n3051, n3052,
    n3053, n3054, n3055, n3056, n3057, n3058,
    n3059, n3060, n3061, n3062, n3063, n3064,
    n3065, n3066, n3067, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076,
    n3077, n3078, n3079, n3080, n3081, n3082,
    n3083, n3084, n3085, n3086, n3087, n3088,
    n3089, n3090, n3091, n3092, n3093, n3094,
    n3095, n3096, n3097, n3098, n3099, n3100,
    n3101, n3102, n3103, n3104, n3105, n3106,
    n3107, n3108, n3109, n3110, n3111, n3112,
    n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3130,
    n3131, n3132, n3133, n3134, n3135, n3136,
    n3137, n3138, n3139, n3140, n3141, n3142,
    n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154,
    n3155, n3156, n3157, n3158, n3159, n3160,
    n3161, n3162, n3163, n3164, n3165, n3166,
    n3167, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179,
    n3180, n3181, n3182, n3183, n3184, n3185,
    n3186, n3187, n3188, n3189, n3190, n3191,
    n3192, n3193, n3194, n3195, n3196, n3197,
    n3198, n3199, n3200, n3201, n3202, n3203,
    n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215,
    n3216, n3217, n3218, n3219, n3220, n3221,
    n3222, n3223, n3224, n3225, n3226, n3227,
    n3228, n3229, n3230, n3231, n3232, n3233,
    n3234, n3235, n3236, n3237, n3238, n3239,
    n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251,
    n3252, n3253, n3254, n3255, n3256, n3257,
    n3258, n3259, n3260, n3261, n3262, n3263,
    n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3272, n3273, n3274, n3275,
    n3276, n3277, n3278, n3279, n3280, n3281,
    n3282, n3283, n3284, n3285, n3286, n3287,
    n3288, n3289, n3290, n3291, n3292, n3293,
    n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305,
    n3306, n3307, n3308, n3309, n3310, n3311,
    n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3321, n3322, n3323,
    n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335,
    n3336, n3337, n3338, n3339, n3340, n3341,
    n3342, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353,
    n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365,
    n3366, n3367, n3368, n3369, n3370, n3371,
    n3372, n3373, n3374, n3375, n3376, n3377,
    n3378, n3379, n3380, n3381, n3382, n3383,
    n3384, n3385, n3386, n3387, n3388, n3389,
    n3390, n3391, n3392, n3393, n3394, n3395,
    n3396, n3397, n3398, n3399, n3400, n3401,
    n3402, n3403, n3404, n3405, n3406, n3407,
    n3408, n3409, n3410, n3411, n3412, n3413,
    n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3426,
    n3427, n3428, n3429, n3430, n3431, n3432,
    n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444,
    n3445, n3446, n3447, n3448, n3449, n3450,
    n3451, n3452, n3453, n3454, n3455, n3456,
    n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474,
    n3475, n3476, n3477, n3478, n3479, n3480,
    n3481, n3482, n3483, n3484, n3485, n3486,
    n3487, n3488, n3489, n3490, n3491, n3492,
    n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504,
    n3505, n3506, n3507, n3508, n3509, n3510,
    n3511, n3512, n3513, n3514, n3515, n3516,
    n3517, n3518, n3519, n3520, n3521, n3522,
    n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534,
    n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546,
    n3547, n3548, n3549, n3550, n3551, n3552,
    n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564,
    n3565, n3566, n3567, n3568, n3569, n3570,
    n3571, n3572, n3573, n3574, n3575, n3576,
    n3577, n3578, n3579, n3580, n3581, n3582,
    n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594,
    n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3603, n3604, n3605, n3606,
    n3607, n3608, n3609, n3610, n3611, n3612,
    n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624,
    n3625, n3626, n3627, n3628, n3629, n3630,
    n3631, n3632, n3633, n3634, n3635, n3636,
    n3637, n3638, n3639, n3640, n3641, n3642,
    n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654,
    n3655, n3656, n3657, n3658, n3659, n3660,
    n3661, n3662, n3663, n3664, n3665, n3666,
    n3667, n3668, n3669, n3670, n3671, n3672,
    n3673, n3674, n3675, n3676, n3677, n3678,
    n3679, n3680, n3681, n3682, n3683, n3684,
    n3685, n3686, n3687, n3688, n3689, n3690,
    n3691, n3693, n3694, n3695, n3696, n3697,
    n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721,
    n3722, n3723, n3724, n3725, n3726, n3727,
    n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751,
    n3752, n3753, n3754, n3755, n3756, n3757,
    n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775,
    n3776, n3777, n3778, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787,
    n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805,
    n3806, n3807, n3808, n3809, n3810, n3811,
    n3812, n3813, n3814, n3815, n3816, n3817,
    n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835,
    n3836, n3837, n3838, n3839, n3840, n3841,
    n3842, n3843, n3844, n3845, n3846, n3847,
    n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865,
    n3866, n3867, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877,
    n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901,
    n3902, n3903, n3904, n3905, n3906, n3907,
    n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931,
    n3932, n3933, n3934, n3935, n3936, n3937,
    n3938, n3939, n3940, n3941, n3942, n3943,
    n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961,
    n3962, n3963, n3964, n3965, n3966, n3967,
    n3968, n3969, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016,
    n4017, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046,
    n4047, n4048, n4049, n4050, n4051, n4052,
    n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082,
    n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214,
    n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232,
    n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317,
    n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341,
    n4342, n4343, n4344, n4345, n4346, n4347,
    n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371,
    n4372, n4373, n4374, n4375, n4376, n4377,
    n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4394, n4395,
    n4396, n4397, n4398, n4399, n4400, n4401,
    n4402, n4403, n4404, n4405, n4406, n4407,
    n4408, n4409, n4410, n4411, n4412, n4413,
    n4414, n4415, n4416, n4417, n4418, n4419,
    n4420, n4421, n4422, n4423, n4424, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431,
    n4432, n4433, n4434, n4435, n4436, n4437,
    n4438, n4439, n4440, n4441, n4442, n4443,
    n4444, n4445, n4446, n4447, n4448, n4449,
    n4450, n4451, n4452, n4453, n4454, n4455,
    n4456, n4457, n4458, n4459, n4460, n4461,
    n4462, n4463, n4464, n4465, n4466, n4467,
    n4468, n4469, n4470, n4471, n4472, n4473,
    n4474, n4475, n4476, n4477, n4478, n4479,
    n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491,
    n4492, n4493, n4494, n4495, n4496, n4497,
    n4498, n4499, n4500, n4501, n4502, n4503,
    n4504, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515,
    n4516, n4517, n4518, n4519, n4520, n4521,
    n4522, n4523, n4524, n4525, n4526, n4527,
    n4528, n4529, n4530, n4531, n4532, n4533,
    n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551,
    n4552, n4553, n4554, n4555, n4556, n4558,
    n4559, n4560, n4561, n4562, n4563, n4564,
    n4565, n4566, n4567, n4568, n4569, n4570,
    n4571, n4572, n4573, n4574, n4575, n4576,
    n4577, n4578, n4579, n4580, n4581, n4582,
    n4583, n4584, n4585, n4586, n4587, n4588,
    n4589, n4590, n4591, n4592, n4593, n4594,
    n4595, n4596, n4597, n4598, n4599, n4600,
    n4601, n4602, n4603, n4604, n4605, n4606,
    n4607, n4608, n4609, n4610, n4611, n4612,
    n4613, n4614, n4615, n4616, n4617, n4618,
    n4619, n4620, n4621, n4622, n4623, n4624,
    n4625, n4626, n4627, n4628, n4629, n4630,
    n4631, n4632, n4633, n4634, n4635, n4636,
    n4637, n4638, n4639, n4640, n4641, n4642,
    n4643, n4644, n4645, n4646, n4647, n4648,
    n4649, n4650, n4651, n4652, n4653, n4654,
    n4655, n4656, n4657, n4658, n4659, n4660,
    n4661, n4662, n4663, n4664, n4665, n4666,
    n4667, n4668, n4669, n4670, n4671, n4672,
    n4673, n4674, n4675, n4676, n4677, n4678,
    n4679, n4680, n4681, n4682, n4683, n4684,
    n4685, n4686, n4687, n4688, n4689, n4690,
    n4691, n4692, n4693, n4694, n4695, n4696,
    n4697, n4698, n4699, n4700, n4701, n4702,
    n4703, n4704, n4705, n4706, n4707, n4708,
    n4709, n4710, n4711, n4712, n4713, n4714,
    n4715, n4716, n4717, n4718, n4719, n4720,
    n4721, n4722, n4723, n4724, n4725, n4726,
    n4727, n4728, n4729, n4730, n4731, n4732,
    n4733, n4734, n4735, n4736, n4737, n4738,
    n4739, n4740, n4741, n4742, n4743, n4744,
    n4745, n4746, n4747, n4748, n4749, n4750,
    n4751, n4752, n4753, n4754, n4755, n4756,
    n4757, n4758, n4759, n4760, n4761, n4762,
    n4763, n4764, n4765, n4766, n4767, n4768,
    n4769, n4770, n4771, n4772, n4773, n4774,
    n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786,
    n4787, n4788, n4789, n4790, n4791, n4792,
    n4793, n4794, n4795, n4796, n4797, n4798,
    n4799, n4800, n4801, n4802, n4803, n4804,
    n4805, n4806, n4807, n4808, n4809, n4810,
    n4811, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822,
    n4823, n4824, n4825, n4826, n4827, n4828,
    n4829, n4830, n4831, n4832, n4833, n4834,
    n4835, n4836, n4837, n4838, n4839, n4840,
    n4841, n4842, n4843, n4844, n4845, n4846,
    n4847, n4848, n4849, n4850, n4851, n4852,
    n4853, n4854, n4855, n4856, n4857, n4858,
    n4859, n4860, n4861, n4862, n4863, n4864,
    n4865, n4867, n4868, n4869, n4870, n4871,
    n4872, n4873, n4874, n4875, n4876, n4877,
    n4878, n4879, n4880, n4881, n4882, n4883,
    n4884, n4885, n4886, n4887, n4888, n4889,
    n4890, n4891, n4892, n4893, n4894, n4895,
    n4896, n4897, n4898, n4899, n4900, n4901,
    n4902, n4903, n4904, n4905, n4906, n4907,
    n4908, n4909, n4910, n4911, n4912, n4913,
    n4914, n4915, n4916, n4917, n4918, n4919,
    n4920, n4921, n4922, n4923, n4924, n4925,
    n4926, n4927, n4928, n4929, n4930, n4931,
    n4932, n4933, n4934, n4935, n4936, n4937,
    n4938, n4939, n4940, n4941, n4942, n4943,
    n4944, n4945, n4946, n4947, n4948, n4949,
    n4950, n4951, n4952, n4953, n4954, n4955,
    n4956, n4957, n4958, n4959, n4960, n4961,
    n4962, n4963, n4964, n4965, n4966, n4967,
    n4968, n4969, n4970, n4971, n4972, n4973,
    n4974, n4975, n4976, n4977, n4978, n4979,
    n4980, n4981, n4982, n4983, n4984, n4985,
    n4986, n4987, n4988, n4989, n4990, n4991,
    n4992, n4993, n4994, n4995, n4996, n4997,
    n4998, n4999, n5000, n5001, n5002, n5003,
    n5004, n5005, n5006, n5007, n5008, n5009,
    n5010, n5011, n5012, n5013, n5014, n5015,
    n5016, n5017, n5018, n5019, n5020, n5021,
    n5022, n5023, n5024, n5025, n5026, n5027,
    n5028, n5029, n5030, n5031, n5032, n5033,
    n5034, n5035, n5036, n5037, n5038, n5039,
    n5040, n5041, n5042, n5043, n5044, n5045,
    n5046, n5047, n5048, n5049, n5050, n5051,
    n5052, n5053, n5054, n5055, n5056, n5057,
    n5058, n5059, n5060, n5061, n5062, n5063,
    n5064, n5065, n5066, n5067, n5068, n5069,
    n5070, n5071, n5072, n5073, n5074, n5075,
    n5076, n5077, n5078, n5079, n5080, n5081,
    n5082, n5083, n5084, n5085, n5086, n5087,
    n5088, n5089, n5090, n5091, n5092, n5093,
    n5094, n5095, n5096, n5097, n5098, n5099,
    n5100, n5101, n5102, n5103, n5104, n5105,
    n5106, n5107, n5108, n5109, n5110, n5111,
    n5112, n5113, n5114, n5115, n5116, n5117,
    n5118, n5119, n5120, n5121, n5122, n5123,
    n5124, n5125, n5126, n5127, n5128, n5129,
    n5130, n5131, n5132, n5133, n5134, n5135,
    n5136, n5137, n5138, n5139, n5140, n5141,
    n5142, n5143, n5144, n5145, n5146, n5147,
    n5148, n5149, n5150, n5151, n5152, n5153,
    n5154, n5155, n5156, n5157, n5158, n5159,
    n5160, n5161, n5162, n5163, n5164, n5165,
    n5166, n5167, n5168, n5169, n5170, n5171,
    n5172, n5173, n5174, n5175, n5176, n5177,
    n5178, n5179, n5180, n5181, n5182, n5183,
    n5184, n5185, n5187, n5188, n5189, n5190,
    n5191, n5192, n5193, n5194, n5195, n5196,
    n5197, n5198, n5199, n5200, n5201, n5202,
    n5203, n5204, n5205, n5206, n5207, n5208,
    n5209, n5210, n5211, n5212, n5213, n5214,
    n5215, n5216, n5217, n5218, n5219, n5220,
    n5221, n5222, n5223, n5224, n5225, n5226,
    n5227, n5228, n5229, n5230, n5231, n5232,
    n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5244,
    n5245, n5246, n5247, n5248, n5249, n5250,
    n5251, n5252, n5253, n5254, n5255, n5256,
    n5257, n5258, n5259, n5260, n5261, n5262,
    n5263, n5264, n5265, n5266, n5267, n5268,
    n5269, n5270, n5271, n5272, n5273, n5274,
    n5275, n5276, n5277, n5278, n5279, n5280,
    n5281, n5282, n5283, n5284, n5285, n5286,
    n5287, n5288, n5289, n5290, n5291, n5292,
    n5293, n5294, n5295, n5296, n5297, n5298,
    n5299, n5300, n5301, n5302, n5303, n5304,
    n5305, n5306, n5307, n5308, n5309, n5310,
    n5311, n5312, n5313, n5314, n5315, n5316,
    n5317, n5318, n5319, n5320, n5321, n5322,
    n5323, n5324, n5325, n5326, n5327, n5328,
    n5329, n5330, n5331, n5332, n5333, n5334,
    n5335, n5336, n5337, n5338, n5339, n5340,
    n5341, n5342, n5343, n5344, n5345, n5346,
    n5347, n5348, n5349, n5350, n5351, n5352,
    n5353, n5354, n5355, n5356, n5357, n5358,
    n5359, n5360, n5361, n5362, n5363, n5364,
    n5365, n5366, n5367, n5368, n5369, n5370,
    n5371, n5372, n5373, n5374, n5375, n5376,
    n5377, n5378, n5379, n5380, n5381, n5382,
    n5383, n5384, n5385, n5386, n5387, n5388,
    n5389, n5390, n5391, n5392, n5393, n5394,
    n5395, n5396, n5397, n5398, n5399, n5400,
    n5401, n5402, n5403, n5404, n5405, n5406,
    n5407, n5408, n5409, n5410, n5411, n5412,
    n5413, n5414, n5415, n5416, n5417, n5418,
    n5419, n5420, n5421, n5422, n5423, n5424,
    n5425, n5426, n5427, n5428, n5429, n5430,
    n5431, n5432, n5433, n5434, n5435, n5436,
    n5437, n5438, n5439, n5440, n5441, n5442,
    n5443, n5444, n5445, n5446, n5447, n5448,
    n5449, n5450, n5451, n5452, n5453, n5454,
    n5455, n5456, n5457, n5458, n5459, n5460,
    n5461, n5462, n5463, n5464, n5465, n5466,
    n5467, n5468, n5469, n5470, n5471, n5472,
    n5473, n5474, n5475, n5476, n5477, n5478,
    n5479, n5480, n5481, n5482, n5483, n5484,
    n5485, n5486, n5487, n5488, n5489, n5490,
    n5491, n5492, n5493, n5494, n5495, n5496,
    n5497, n5498, n5499, n5500, n5501, n5502,
    n5503, n5504, n5505, n5506, n5507, n5508,
    n5509, n5510, n5511, n5512, n5513, n5514,
    n5515, n5517, n5518, n5519, n5520, n5521,
    n5522, n5523, n5524, n5525, n5526, n5527,
    n5528, n5529, n5530, n5531, n5532, n5533,
    n5534, n5535, n5536, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551,
    n5552, n5553, n5554, n5555, n5556, n5557,
    n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581,
    n5582, n5583, n5584, n5585, n5586, n5587,
    n5588, n5589, n5590, n5591, n5592, n5593,
    n5594, n5595, n5596, n5597, n5598, n5599,
    n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611,
    n5612, n5613, n5614, n5615, n5616, n5617,
    n5618, n5619, n5620, n5621, n5622, n5623,
    n5624, n5625, n5626, n5627, n5628, n5629,
    n5630, n5631, n5632, n5633, n5634, n5635,
    n5636, n5637, n5638, n5639, n5640, n5641,
    n5642, n5643, n5644, n5645, n5646, n5647,
    n5648, n5649, n5650, n5651, n5652, n5653,
    n5654, n5655, n5656, n5657, n5658, n5659,
    n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5667, n5668, n5669, n5670, n5671,
    n5672, n5673, n5674, n5675, n5676, n5677,
    n5678, n5679, n5680, n5681, n5682, n5683,
    n5684, n5685, n5686, n5687, n5688, n5689,
    n5690, n5691, n5692, n5693, n5694, n5695,
    n5696, n5697, n5698, n5699, n5700, n5701,
    n5702, n5703, n5704, n5705, n5706, n5707,
    n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5715, n5716, n5717, n5718, n5719,
    n5720, n5721, n5722, n5723, n5724, n5725,
    n5726, n5727, n5728, n5729, n5730, n5731,
    n5732, n5733, n5734, n5735, n5736, n5737,
    n5738, n5739, n5740, n5741, n5742, n5743,
    n5744, n5745, n5746, n5747, n5748, n5749,
    n5750, n5751, n5752, n5753, n5754, n5755,
    n5756, n5757, n5758, n5759, n5760, n5761,
    n5762, n5763, n5764, n5765, n5766, n5767,
    n5768, n5769, n5770, n5771, n5772, n5773,
    n5774, n5775, n5776, n5777, n5778, n5779,
    n5780, n5781, n5782, n5783, n5784, n5785,
    n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5794, n5795, n5796, n5797,
    n5798, n5799, n5800, n5801, n5802, n5803,
    n5804, n5805, n5806, n5807, n5808, n5809,
    n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5817, n5818, n5819, n5820, n5821,
    n5822, n5823, n5824, n5825, n5826, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833,
    n5834, n5835, n5836, n5837, n5838, n5839,
    n5840, n5841, n5842, n5843, n5844, n5845,
    n5846, n5847, n5848, n5849, n5850, n5851,
    n5852, n5853, n5854, n5855, n5856, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864,
    n5865, n5866, n5867, n5868, n5869, n5870,
    n5871, n5872, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5881, n5882,
    n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894,
    n5895, n5896, n5897, n5898, n5899, n5900,
    n5901, n5902, n5903, n5904, n5905, n5906,
    n5907, n5908, n5909, n5910, n5911, n5912,
    n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924,
    n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954,
    n5955, n5956, n5957, n5958, n5959, n5960,
    n5961, n5962, n5963, n5964, n5965, n5966,
    n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984,
    n5985, n5986, n5987, n5988, n5989, n5990,
    n5991, n5992, n5993, n5994, n5995, n5996,
    n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008,
    n6009, n6010, n6011, n6012, n6013, n6014,
    n6015, n6016, n6017, n6018, n6019, n6020,
    n6021, n6022, n6023, n6024, n6025, n6026,
    n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038,
    n6039, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050,
    n6051, n6052, n6053, n6054, n6055, n6056,
    n6057, n6058, n6059, n6060, n6061, n6062,
    n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074,
    n6075, n6076, n6077, n6078, n6079, n6080,
    n6081, n6082, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6090, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6107, n6108, n6109, n6110,
    n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6119, n6120, n6121, n6122,
    n6123, n6124, n6125, n6126, n6127, n6128,
    n6129, n6130, n6131, n6132, n6133, n6134,
    n6135, n6136, n6137, n6138, n6139, n6140,
    n6141, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170,
    n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6209, n6210, n6211, n6212, n6213,
    n6214, n6215, n6216, n6217, n6218, n6219,
    n6220, n6221, n6222, n6223, n6224, n6225,
    n6226, n6227, n6228, n6229, n6230, n6231,
    n6232, n6233, n6234, n6235, n6236, n6237,
    n6238, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255,
    n6256, n6257, n6258, n6259, n6260, n6261,
    n6262, n6263, n6264, n6265, n6266, n6267,
    n6268, n6269, n6270, n6271, n6272, n6273,
    n6274, n6275, n6276, n6277, n6278, n6279,
    n6280, n6281, n6282, n6283, n6284, n6285,
    n6286, n6287, n6288, n6289, n6290, n6291,
    n6292, n6293, n6294, n6295, n6296, n6297,
    n6298, n6299, n6300, n6301, n6302, n6303,
    n6304, n6305, n6306, n6307, n6308, n6309,
    n6310, n6311, n6312, n6313, n6314, n6315,
    n6316, n6317, n6318, n6319, n6320, n6321,
    n6322, n6323, n6324, n6325, n6326, n6327,
    n6328, n6329, n6330, n6331, n6332, n6333,
    n6334, n6335, n6336, n6337, n6338, n6339,
    n6340, n6341, n6342, n6343, n6344, n6345,
    n6346, n6347, n6348, n6349, n6350, n6351,
    n6352, n6353, n6354, n6355, n6356, n6357,
    n6358, n6359, n6360, n6361, n6362, n6363,
    n6364, n6365, n6366, n6367, n6368, n6369,
    n6370, n6371, n6372, n6373, n6374, n6375,
    n6376, n6377, n6378, n6379, n6380, n6381,
    n6382, n6383, n6384, n6385, n6386, n6387,
    n6388, n6389, n6390, n6391, n6392, n6393,
    n6394, n6395, n6396, n6397, n6398, n6399,
    n6400, n6401, n6402, n6403, n6404, n6405,
    n6406, n6407, n6408, n6409, n6410, n6411,
    n6412, n6413, n6414, n6415, n6416, n6417,
    n6418, n6419, n6420, n6421, n6422, n6423,
    n6424, n6425, n6426, n6427, n6428, n6429,
    n6430, n6431, n6432, n6433, n6434, n6435,
    n6436, n6437, n6438, n6439, n6440, n6441,
    n6442, n6443, n6444, n6445, n6446, n6447,
    n6448, n6449, n6450, n6451, n6452, n6453,
    n6454, n6455, n6456, n6457, n6458, n6459,
    n6460, n6461, n6462, n6463, n6464, n6465,
    n6466, n6467, n6468, n6469, n6470, n6471,
    n6472, n6473, n6474, n6475, n6476, n6477,
    n6478, n6479, n6480, n6481, n6482, n6483,
    n6484, n6485, n6486, n6487, n6488, n6489,
    n6490, n6491, n6492, n6493, n6494, n6495,
    n6496, n6497, n6498, n6499, n6500, n6501,
    n6502, n6503, n6504, n6505, n6506, n6507,
    n6508, n6509, n6510, n6511, n6512, n6513,
    n6514, n6515, n6516, n6517, n6518, n6519,
    n6520, n6521, n6522, n6523, n6524, n6525,
    n6526, n6527, n6528, n6529, n6530, n6531,
    n6532, n6533, n6534, n6535, n6536, n6537,
    n6538, n6539, n6540, n6541, n6542, n6543,
    n6544, n6545, n6546, n6547, n6548, n6549,
    n6550, n6551, n6552, n6553, n6554, n6555,
    n6556, n6557, n6558, n6559, n6560, n6561,
    n6562, n6563, n6564, n6565, n6566, n6567,
    n6568, n6569, n6571, n6572, n6573, n6574,
    n6575, n6576, n6577, n6578, n6579, n6580,
    n6581, n6582, n6583, n6584, n6585, n6586,
    n6587, n6588, n6589, n6590, n6591, n6592,
    n6593, n6594, n6595, n6596, n6597, n6598,
    n6599, n6600, n6601, n6602, n6603, n6604,
    n6605, n6606, n6607, n6608, n6609, n6610,
    n6611, n6612, n6613, n6614, n6615, n6616,
    n6617, n6618, n6619, n6620, n6621, n6622,
    n6623, n6624, n6625, n6626, n6627, n6628,
    n6629, n6630, n6631, n6632, n6633, n6634,
    n6635, n6636, n6637, n6638, n6639, n6640,
    n6641, n6642, n6643, n6644, n6645, n6646,
    n6647, n6648, n6649, n6650, n6651, n6652,
    n6653, n6654, n6655, n6656, n6657, n6658,
    n6659, n6660, n6661, n6662, n6663, n6664,
    n6665, n6666, n6667, n6668, n6669, n6670,
    n6671, n6672, n6673, n6674, n6675, n6676,
    n6677, n6678, n6679, n6680, n6681, n6682,
    n6683, n6684, n6685, n6686, n6687, n6688,
    n6689, n6690, n6691, n6692, n6693, n6694,
    n6695, n6696, n6697, n6698, n6699, n6700,
    n6701, n6702, n6703, n6704, n6705, n6706,
    n6707, n6708, n6709, n6710, n6711, n6712,
    n6713, n6714, n6715, n6716, n6717, n6718,
    n6719, n6720, n6721, n6722, n6723, n6724,
    n6725, n6726, n6727, n6728, n6729, n6730,
    n6731, n6732, n6733, n6734, n6735, n6736,
    n6737, n6738, n6739, n6740, n6741, n6742,
    n6743, n6744, n6745, n6746, n6747, n6748,
    n6749, n6750, n6751, n6752, n6753, n6754,
    n6755, n6756, n6757, n6758, n6759, n6760,
    n6761, n6762, n6763, n6764, n6765, n6766,
    n6767, n6768, n6769, n6770, n6771, n6772,
    n6773, n6774, n6775, n6776, n6777, n6778,
    n6779, n6780, n6781, n6782, n6783, n6784,
    n6785, n6786, n6787, n6788, n6789, n6790,
    n6791, n6792, n6793, n6794, n6795, n6796,
    n6797, n6798, n6799, n6800, n6801, n6802,
    n6803, n6804, n6805, n6806, n6807, n6808,
    n6809, n6810, n6811, n6812, n6813, n6814,
    n6815, n6816, n6817, n6818, n6819, n6820,
    n6821, n6822, n6823, n6824, n6825, n6826,
    n6827, n6828, n6829, n6830, n6831, n6832,
    n6833, n6834, n6835, n6836, n6837, n6838,
    n6839, n6840, n6841, n6842, n6843, n6844,
    n6845, n6846, n6847, n6848, n6849, n6850,
    n6851, n6852, n6853, n6854, n6855, n6856,
    n6857, n6858, n6859, n6860, n6861, n6862,
    n6863, n6864, n6865, n6866, n6867, n6868,
    n6869, n6870, n6871, n6872, n6873, n6874,
    n6875, n6876, n6877, n6878, n6879, n6880,
    n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n6891, n6892,
    n6893, n6894, n6895, n6896, n6897, n6898,
    n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6943, n6944, n6945, n6946, n6947,
    n6948, n6949, n6950, n6951, n6952, n6953,
    n6954, n6955, n6956, n6957, n6958, n6959,
    n6960, n6961, n6962, n6963, n6964, n6965,
    n6966, n6967, n6968, n6969, n6970, n6971,
    n6972, n6973, n6974, n6975, n6976, n6977,
    n6978, n6979, n6980, n6981, n6982, n6983,
    n6984, n6985, n6986, n6987, n6988, n6989,
    n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7001,
    n7002, n7003, n7004, n7005, n7006, n7007,
    n7008, n7009, n7010, n7011, n7012, n7013,
    n7014, n7015, n7016, n7017, n7018, n7019,
    n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031,
    n7032, n7033, n7034, n7035, n7036, n7037,
    n7038, n7039, n7040, n7041, n7042, n7043,
    n7044, n7045, n7046, n7047, n7048, n7049,
    n7050, n7051, n7052, n7053, n7054, n7055,
    n7056, n7057, n7058, n7059, n7060, n7061,
    n7062, n7063, n7064, n7065, n7066, n7067,
    n7068, n7069, n7070, n7071, n7072, n7073,
    n7074, n7075, n7076, n7077, n7078, n7079,
    n7080, n7081, n7082, n7083, n7084, n7085,
    n7086, n7087, n7088, n7089, n7090, n7091,
    n7092, n7093, n7094, n7095, n7096, n7097,
    n7098, n7099, n7100, n7101, n7102, n7103,
    n7104, n7105, n7106, n7107, n7108, n7109,
    n7110, n7111, n7112, n7113, n7114, n7115,
    n7116, n7117, n7118, n7119, n7120, n7121,
    n7122, n7123, n7124, n7125, n7126, n7127,
    n7128, n7129, n7130, n7131, n7132, n7133,
    n7134, n7135, n7136, n7137, n7138, n7139,
    n7140, n7141, n7142, n7143, n7144, n7145,
    n7146, n7147, n7148, n7149, n7150, n7151,
    n7152, n7153, n7154, n7155, n7156, n7157,
    n7158, n7159, n7160, n7161, n7162, n7163,
    n7164, n7165, n7166, n7167, n7168, n7169,
    n7170, n7171, n7172, n7173, n7174, n7175,
    n7176, n7177, n7178, n7179, n7180, n7181,
    n7182, n7183, n7184, n7185, n7186, n7187,
    n7188, n7189, n7190, n7191, n7192, n7193,
    n7194, n7195, n7196, n7197, n7198, n7199,
    n7200, n7201, n7202, n7203, n7204, n7205,
    n7206, n7207, n7208, n7209, n7210, n7211,
    n7212, n7213, n7214, n7215, n7216, n7217,
    n7218, n7219, n7220, n7221, n7222, n7223,
    n7224, n7225, n7226, n7227, n7228, n7229,
    n7230, n7231, n7232, n7233, n7234, n7235,
    n7236, n7237, n7238, n7239, n7240, n7241,
    n7242, n7243, n7244, n7245, n7246, n7247,
    n7248, n7249, n7250, n7251, n7252, n7253,
    n7254, n7255, n7256, n7257, n7258, n7259,
    n7260, n7261, n7262, n7263, n7264, n7265,
    n7266, n7267, n7268, n7269, n7270, n7271,
    n7272, n7273, n7274, n7275, n7276, n7277,
    n7278, n7279, n7280, n7281, n7282, n7283,
    n7284, n7285, n7286, n7287, n7288, n7289,
    n7290, n7291, n7292, n7293, n7294, n7295,
    n7296, n7297, n7298, n7299, n7300, n7301,
    n7302, n7303, n7304, n7305, n7306, n7307,
    n7308, n7309, n7310, n7311, n7312, n7313,
    n7314, n7315, n7316, n7317, n7318, n7319,
    n7320, n7321, n7322, n7323, n7324, n7326,
    n7327, n7328, n7329, n7330, n7331, n7332,
    n7333, n7334, n7335, n7336, n7337, n7338,
    n7339, n7340, n7341, n7342, n7343, n7344,
    n7345, n7346, n7347, n7348, n7349, n7350,
    n7351, n7352, n7353, n7354, n7355, n7356,
    n7357, n7358, n7359, n7360, n7361, n7362,
    n7363, n7364, n7365, n7366, n7367, n7368,
    n7369, n7370, n7371, n7372, n7373, n7374,
    n7375, n7376, n7377, n7378, n7379, n7380,
    n7381, n7382, n7383, n7384, n7385, n7386,
    n7387, n7388, n7389, n7390, n7391, n7392,
    n7393, n7394, n7395, n7396, n7397, n7398,
    n7399, n7400, n7401, n7402, n7403, n7404,
    n7405, n7406, n7407, n7408, n7409, n7410,
    n7411, n7412, n7413, n7414, n7415, n7416,
    n7417, n7418, n7419, n7420, n7421, n7422,
    n7423, n7424, n7425, n7426, n7427, n7428,
    n7429, n7430, n7431, n7432, n7433, n7434,
    n7435, n7436, n7437, n7438, n7439, n7440,
    n7441, n7442, n7443, n7444, n7445, n7446,
    n7447, n7448, n7449, n7450, n7451, n7452,
    n7453, n7454, n7455, n7456, n7457, n7458,
    n7459, n7460, n7461, n7462, n7463, n7464,
    n7465, n7466, n7467, n7468, n7469, n7470,
    n7471, n7472, n7473, n7474, n7475, n7476,
    n7477, n7478, n7479, n7480, n7481, n7482,
    n7483, n7484, n7485, n7486, n7487, n7488,
    n7489, n7490, n7491, n7492, n7493, n7494,
    n7495, n7496, n7497, n7498, n7499, n7500,
    n7501, n7502, n7503, n7504, n7505, n7506,
    n7507, n7508, n7509, n7510, n7511, n7512,
    n7513, n7514, n7515, n7516, n7517, n7518,
    n7519, n7520, n7521, n7522, n7523, n7524,
    n7525, n7526, n7527, n7528, n7529, n7530,
    n7531, n7532, n7533, n7534, n7535, n7536,
    n7537, n7538, n7539, n7540, n7541, n7542,
    n7543, n7544, n7545, n7546, n7547, n7548,
    n7549, n7550, n7551, n7552, n7553, n7554,
    n7555, n7556, n7557, n7558, n7559, n7560,
    n7561, n7562, n7563, n7564, n7565, n7566,
    n7567, n7568, n7569, n7570, n7571, n7572,
    n7573, n7574, n7575, n7576, n7577, n7578,
    n7579, n7580, n7581, n7582, n7583, n7584,
    n7585, n7586, n7587, n7588, n7589, n7590,
    n7591, n7592, n7593, n7594, n7595, n7596,
    n7597, n7598, n7599, n7600, n7601, n7602,
    n7603, n7604, n7605, n7606, n7607, n7608,
    n7609, n7610, n7611, n7612, n7613, n7614,
    n7615, n7616, n7617, n7618, n7619, n7620,
    n7621, n7622, n7623, n7624, n7625, n7626,
    n7627, n7628, n7629, n7630, n7631, n7632,
    n7633, n7634, n7635, n7636, n7637, n7638,
    n7639, n7640, n7641, n7642, n7643, n7644,
    n7645, n7646, n7647, n7648, n7649, n7650,
    n7651, n7652, n7653, n7654, n7655, n7656,
    n7657, n7658, n7659, n7660, n7661, n7662,
    n7663, n7664, n7665, n7666, n7667, n7668,
    n7669, n7670, n7671, n7672, n7673, n7674,
    n7675, n7676, n7677, n7678, n7679, n7680,
    n7681, n7682, n7683, n7684, n7685, n7686,
    n7687, n7688, n7689, n7690, n7691, n7692,
    n7693, n7694, n7695, n7696, n7697, n7698,
    n7699, n7700, n7701, n7702, n7703, n7704,
    n7705, n7706, n7707, n7708, n7709, n7710,
    n7711, n7712, n7713, n7714, n7715, n7716,
    n7717, n7719, n7720, n7721, n7722, n7723,
    n7724, n7725, n7726, n7727, n7728, n7729,
    n7730, n7731, n7732, n7733, n7734, n7735,
    n7736, n7737, n7738, n7739, n7740, n7741,
    n7742, n7743, n7744, n7745, n7746, n7747,
    n7748, n7749, n7750, n7751, n7752, n7753,
    n7754, n7755, n7756, n7757, n7758, n7759,
    n7760, n7761, n7762, n7763, n7764, n7765,
    n7766, n7767, n7768, n7769, n7770, n7771,
    n7772, n7773, n7774, n7775, n7776, n7777,
    n7778, n7779, n7780, n7781, n7782, n7783,
    n7784, n7785, n7786, n7787, n7788, n7789,
    n7790, n7791, n7792, n7793, n7794, n7795,
    n7796, n7797, n7798, n7799, n7800, n7801,
    n7802, n7803, n7804, n7805, n7806, n7807,
    n7808, n7809, n7810, n7811, n7812, n7813,
    n7814, n7815, n7816, n7817, n7818, n7819,
    n7820, n7821, n7822, n7823, n7824, n7825,
    n7826, n7827, n7828, n7829, n7830, n7831,
    n7832, n7833, n7834, n7835, n7836, n7837,
    n7838, n7839, n7840, n7841, n7842, n7843,
    n7844, n7845, n7846, n7847, n7848, n7849,
    n7850, n7851, n7852, n7853, n7854, n7855,
    n7856, n7857, n7858, n7859, n7860, n7861,
    n7862, n7863, n7864, n7865, n7866, n7867,
    n7868, n7869, n7870, n7871, n7872, n7873,
    n7874, n7875, n7876, n7877, n7878, n7879,
    n7880, n7881, n7882, n7883, n7884, n7885,
    n7886, n7887, n7888, n7889, n7890, n7891,
    n7892, n7893, n7894, n7895, n7896, n7897,
    n7898, n7899, n7900, n7901, n7902, n7903,
    n7904, n7905, n7906, n7907, n7908, n7909,
    n7910, n7911, n7912, n7913, n7914, n7915,
    n7916, n7917, n7918, n7919, n7920, n7921,
    n7922, n7923, n7924, n7925, n7926, n7927,
    n7928, n7929, n7930, n7931, n7932, n7933,
    n7934, n7935, n7936, n7937, n7938, n7939,
    n7940, n7941, n7942, n7943, n7944, n7945,
    n7946, n7947, n7948, n7949, n7950, n7951,
    n7952, n7953, n7954, n7955, n7956, n7957,
    n7958, n7959, n7960, n7961, n7962, n7963,
    n7964, n7965, n7966, n7967, n7968, n7969,
    n7970, n7971, n7972, n7973, n7974, n7975,
    n7976, n7977, n7978, n7979, n7980, n7981,
    n7982, n7983, n7984, n7985, n7986, n7987,
    n7988, n7989, n7990, n7991, n7992, n7993,
    n7994, n7995, n7996, n7997, n7998, n7999,
    n8000, n8001, n8002, n8003, n8004, n8005,
    n8006, n8007, n8008, n8009, n8010, n8011,
    n8012, n8013, n8014, n8015, n8016, n8017,
    n8018, n8019, n8020, n8021, n8022, n8023,
    n8024, n8025, n8026, n8027, n8028, n8029,
    n8030, n8031, n8032, n8033, n8034, n8035,
    n8036, n8037, n8038, n8039, n8040, n8041,
    n8042, n8043, n8044, n8045, n8046, n8047,
    n8048, n8049, n8050, n8051, n8052, n8053,
    n8054, n8055, n8056, n8057, n8058, n8059,
    n8060, n8061, n8062, n8063, n8064, n8065,
    n8066, n8067, n8068, n8069, n8070, n8071,
    n8072, n8073, n8074, n8075, n8076, n8077,
    n8078, n8079, n8080, n8081, n8082, n8083,
    n8084, n8085, n8086, n8087, n8088, n8089,
    n8090, n8091, n8092, n8093, n8094, n8095,
    n8096, n8097, n8098, n8099, n8100, n8101,
    n8102, n8103, n8104, n8105, n8106, n8107,
    n8108, n8109, n8110, n8111, n8112, n8113,
    n8114, n8115, n8116, n8117, n8118, n8119,
    n8120, n8121, n8123, n8124, n8125, n8126,
    n8127, n8128, n8129, n8130, n8131, n8132,
    n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144,
    n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156,
    n8157, n8158, n8159, n8160, n8161, n8162,
    n8163, n8164, n8165, n8166, n8167, n8168,
    n8169, n8170, n8171, n8172, n8173, n8174,
    n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186,
    n8187, n8188, n8189, n8190, n8191, n8192,
    n8193, n8194, n8195, n8196, n8197, n8198,
    n8199, n8200, n8201, n8202, n8203, n8204,
    n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216,
    n8217, n8218, n8219, n8220, n8221, n8222,
    n8223, n8224, n8225, n8226, n8227, n8228,
    n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246,
    n8247, n8248, n8249, n8250, n8251, n8252,
    n8253, n8254, n8255, n8256, n8257, n8258,
    n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276,
    n8277, n8278, n8279, n8280, n8281, n8282,
    n8283, n8284, n8285, n8286, n8287, n8288,
    n8289, n8290, n8291, n8292, n8293, n8294,
    n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306,
    n8307, n8308, n8309, n8310, n8311, n8312,
    n8313, n8314, n8315, n8316, n8317, n8318,
    n8319, n8320, n8321, n8322, n8323, n8324,
    n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336,
    n8337, n8338, n8339, n8340, n8341, n8342,
    n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360,
    n8361, n8362, n8363, n8364, n8365, n8366,
    n8367, n8368, n8369, n8370, n8371, n8372,
    n8373, n8374, n8375, n8376, n8377, n8378,
    n8379, n8380, n8381, n8382, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396,
    n8397, n8398, n8399, n8400, n8401, n8402,
    n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414,
    n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444,
    n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456,
    n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486,
    n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504,
    n8505, n8506, n8507, n8508, n8509, n8510,
    n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528,
    n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8537, n8538, n8539, n8540, n8541,
    n8542, n8543, n8544, n8545, n8546, n8547,
    n8548, n8549, n8550, n8551, n8552, n8553,
    n8554, n8555, n8556, n8557, n8558, n8559,
    n8560, n8561, n8562, n8563, n8564, n8565,
    n8566, n8567, n8568, n8569, n8570, n8571,
    n8572, n8573, n8574, n8575, n8576, n8577,
    n8578, n8579, n8580, n8581, n8582, n8583,
    n8584, n8585, n8586, n8587, n8588, n8589,
    n8590, n8591, n8592, n8593, n8594, n8595,
    n8596, n8597, n8598, n8599, n8600, n8601,
    n8602, n8603, n8604, n8605, n8606, n8607,
    n8608, n8609, n8610, n8611, n8612, n8613,
    n8614, n8615, n8616, n8617, n8618, n8619,
    n8620, n8621, n8622, n8623, n8624, n8625,
    n8626, n8627, n8628, n8629, n8630, n8631,
    n8632, n8633, n8634, n8635, n8636, n8637,
    n8638, n8639, n8640, n8641, n8642, n8643,
    n8644, n8645, n8646, n8647, n8648, n8649,
    n8650, n8651, n8652, n8653, n8654, n8655,
    n8656, n8657, n8658, n8659, n8660, n8661,
    n8662, n8663, n8664, n8665, n8666, n8667,
    n8668, n8669, n8670, n8671, n8672, n8673,
    n8674, n8675, n8676, n8677, n8678, n8679,
    n8680, n8681, n8682, n8683, n8684, n8685,
    n8686, n8687, n8688, n8689, n8690, n8691,
    n8692, n8693, n8694, n8695, n8696, n8697,
    n8698, n8699, n8700, n8701, n8702, n8703,
    n8704, n8705, n8706, n8707, n8708, n8709,
    n8710, n8711, n8712, n8713, n8714, n8715,
    n8716, n8717, n8718, n8719, n8720, n8721,
    n8722, n8723, n8724, n8725, n8726, n8727,
    n8728, n8729, n8730, n8731, n8732, n8733,
    n8734, n8735, n8736, n8737, n8738, n8739,
    n8740, n8741, n8742, n8743, n8744, n8745,
    n8746, n8747, n8748, n8749, n8750, n8751,
    n8752, n8753, n8754, n8755, n8756, n8757,
    n8758, n8759, n8760, n8761, n8762, n8763,
    n8764, n8765, n8766, n8767, n8768, n8769,
    n8770, n8771, n8772, n8773, n8774, n8775,
    n8776, n8777, n8778, n8779, n8780, n8781,
    n8782, n8783, n8784, n8785, n8786, n8787,
    n8788, n8789, n8790, n8791, n8792, n8793,
    n8794, n8795, n8796, n8797, n8798, n8799,
    n8800, n8801, n8802, n8803, n8804, n8805,
    n8806, n8807, n8808, n8809, n8810, n8811,
    n8812, n8813, n8814, n8815, n8816, n8817,
    n8818, n8819, n8820, n8821, n8822, n8823,
    n8824, n8825, n8826, n8827, n8828, n8829,
    n8830, n8831, n8832, n8833, n8834, n8835,
    n8836, n8837, n8838, n8839, n8840, n8841,
    n8842, n8843, n8844, n8845, n8846, n8847,
    n8848, n8849, n8850, n8851, n8852, n8853,
    n8854, n8855, n8856, n8857, n8858, n8859,
    n8860, n8861, n8862, n8863, n8864, n8865,
    n8866, n8867, n8868, n8869, n8870, n8871,
    n8872, n8873, n8874, n8875, n8876, n8877,
    n8878, n8879, n8880, n8881, n8882, n8883,
    n8884, n8885, n8886, n8887, n8888, n8889,
    n8890, n8891, n8892, n8893, n8894, n8895,
    n8896, n8897, n8898, n8899, n8900, n8901,
    n8902, n8903, n8904, n8905, n8906, n8907,
    n8908, n8909, n8910, n8911, n8912, n8913,
    n8914, n8915, n8916, n8917, n8918, n8919,
    n8920, n8921, n8922, n8923, n8924, n8925,
    n8926, n8927, n8928, n8929, n8930, n8931,
    n8932, n8933, n8934, n8935, n8936, n8937,
    n8938, n8939, n8940, n8941, n8942, n8943,
    n8944, n8945, n8946, n8947, n8948, n8949,
    n8950, n8951, n8952, n8953, n8954, n8955,
    n8956, n8957, n8958, n8959, n8960, n8962,
    n8963, n8964, n8965, n8966, n8967, n8968,
    n8969, n8970, n8971, n8972, n8973, n8974,
    n8975, n8976, n8977, n8978, n8979, n8980,
    n8981, n8982, n8983, n8984, n8985, n8986,
    n8987, n8988, n8989, n8990, n8991, n8992,
    n8993, n8994, n8995, n8996, n8997, n8998,
    n8999, n9000, n9001, n9002, n9003, n9004,
    n9005, n9006, n9007, n9008, n9009, n9010,
    n9011, n9012, n9013, n9014, n9015, n9016,
    n9017, n9018, n9019, n9020, n9021, n9022,
    n9023, n9024, n9025, n9026, n9027, n9028,
    n9029, n9030, n9031, n9032, n9033, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040,
    n9041, n9042, n9043, n9044, n9045, n9046,
    n9047, n9048, n9049, n9050, n9051, n9052,
    n9053, n9054, n9055, n9056, n9057, n9058,
    n9059, n9060, n9061, n9062, n9063, n9064,
    n9065, n9066, n9067, n9068, n9069, n9070,
    n9071, n9072, n9073, n9074, n9075, n9076,
    n9077, n9078, n9079, n9080, n9081, n9082,
    n9083, n9084, n9085, n9086, n9087, n9088,
    n9089, n9090, n9091, n9092, n9093, n9094,
    n9095, n9096, n9097, n9098, n9099, n9100,
    n9101, n9102, n9103, n9104, n9105, n9106,
    n9107, n9108, n9109, n9110, n9111, n9112,
    n9113, n9114, n9115, n9116, n9117, n9118,
    n9119, n9120, n9121, n9122, n9123, n9124,
    n9125, n9126, n9127, n9128, n9129, n9130,
    n9131, n9132, n9133, n9134, n9135, n9136,
    n9137, n9138, n9139, n9140, n9141, n9142,
    n9143, n9144, n9145, n9146, n9147, n9148,
    n9149, n9150, n9151, n9152, n9153, n9154,
    n9155, n9156, n9157, n9158, n9159, n9160,
    n9161, n9162, n9163, n9164, n9165, n9166,
    n9167, n9168, n9169, n9170, n9171, n9172,
    n9173, n9174, n9175, n9176, n9177, n9178,
    n9179, n9180, n9181, n9182, n9183, n9184,
    n9185, n9186, n9187, n9188, n9189, n9190,
    n9191, n9192, n9193, n9194, n9195, n9196,
    n9197, n9198, n9199, n9200, n9201, n9202,
    n9203, n9204, n9205, n9206, n9207, n9208,
    n9209, n9210, n9211, n9212, n9213, n9214,
    n9215, n9216, n9217, n9218, n9219, n9220,
    n9221, n9222, n9223, n9224, n9225, n9226,
    n9227, n9228, n9229, n9230, n9231, n9232,
    n9233, n9234, n9235, n9236, n9237, n9238,
    n9239, n9240, n9241, n9242, n9243, n9244,
    n9245, n9246, n9247, n9248, n9249, n9250,
    n9251, n9252, n9253, n9254, n9255, n9256,
    n9257, n9258, n9259, n9260, n9261, n9262,
    n9263, n9264, n9265, n9266, n9267, n9268,
    n9269, n9270, n9271, n9272, n9273, n9274,
    n9275, n9276, n9277, n9278, n9279, n9280,
    n9281, n9282, n9283, n9284, n9285, n9286,
    n9287, n9288, n9289, n9290, n9291, n9292,
    n9293, n9294, n9295, n9296, n9297, n9298,
    n9299, n9300, n9301, n9302, n9303, n9304,
    n9305, n9306, n9307, n9308, n9309, n9310,
    n9311, n9312, n9313, n9314, n9315, n9316,
    n9317, n9318, n9319, n9320, n9321, n9322,
    n9323, n9324, n9325, n9326, n9327, n9328,
    n9329, n9330, n9331, n9332, n9333, n9334,
    n9335, n9336, n9337, n9338, n9339, n9340,
    n9341, n9342, n9343, n9344, n9345, n9346,
    n9347, n9348, n9349, n9350, n9351, n9352,
    n9353, n9354, n9355, n9356, n9357, n9358,
    n9359, n9360, n9361, n9362, n9363, n9364,
    n9365, n9366, n9367, n9368, n9369, n9370,
    n9371, n9372, n9373, n9374, n9375, n9376,
    n9377, n9378, n9379, n9380, n9381, n9382,
    n9383, n9384, n9385, n9386, n9387, n9388,
    n9389, n9390, n9391, n9392, n9393, n9394,
    n9395, n9397, n9398, n9399, n9400, n9401,
    n9402, n9403, n9404, n9405, n9406, n9407,
    n9408, n9409, n9410, n9411, n9412, n9413,
    n9414, n9415, n9416, n9417, n9418, n9419,
    n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431,
    n9432, n9433, n9434, n9435, n9436, n9437,
    n9438, n9439, n9440, n9441, n9442, n9443,
    n9444, n9445, n9446, n9447, n9448, n9449,
    n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461,
    n9462, n9463, n9464, n9465, n9466, n9467,
    n9468, n9469, n9470, n9471, n9472, n9473,
    n9474, n9475, n9476, n9477, n9478, n9479,
    n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491,
    n9492, n9493, n9494, n9495, n9496, n9497,
    n9498, n9499, n9500, n9501, n9502, n9503,
    n9504, n9505, n9506, n9507, n9508, n9509,
    n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521,
    n9522, n9523, n9524, n9525, n9526, n9527,
    n9528, n9529, n9530, n9531, n9532, n9533,
    n9534, n9535, n9536, n9537, n9538, n9539,
    n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9547, n9548, n9549, n9550, n9551,
    n9552, n9553, n9554, n9555, n9556, n9557,
    n9558, n9559, n9560, n9561, n9562, n9563,
    n9564, n9565, n9566, n9567, n9568, n9569,
    n9570, n9571, n9572, n9573, n9574, n9575,
    n9576, n9577, n9578, n9579, n9580, n9581,
    n9582, n9583, n9584, n9585, n9586, n9587,
    n9588, n9589, n9590, n9591, n9592, n9593,
    n9594, n9595, n9596, n9597, n9598, n9599,
    n9600, n9601, n9602, n9603, n9604, n9605,
    n9606, n9607, n9608, n9609, n9610, n9611,
    n9612, n9613, n9614, n9615, n9616, n9617,
    n9618, n9619, n9620, n9621, n9622, n9623,
    n9624, n9625, n9626, n9627, n9628, n9629,
    n9630, n9631, n9632, n9633, n9634, n9635,
    n9636, n9637, n9638, n9639, n9640, n9641,
    n9642, n9643, n9644, n9645, n9646, n9647,
    n9648, n9649, n9650, n9651, n9652, n9653,
    n9654, n9655, n9656, n9657, n9658, n9659,
    n9660, n9661, n9662, n9663, n9664, n9665,
    n9666, n9667, n9668, n9669, n9670, n9671,
    n9672, n9673, n9674, n9675, n9676, n9677,
    n9678, n9679, n9680, n9681, n9682, n9683,
    n9684, n9685, n9686, n9687, n9688, n9689,
    n9690, n9691, n9692, n9693, n9694, n9695,
    n9696, n9697, n9698, n9699, n9700, n9701,
    n9702, n9703, n9704, n9705, n9706, n9707,
    n9708, n9709, n9710, n9711, n9712, n9713,
    n9714, n9715, n9716, n9717, n9718, n9719,
    n9720, n9721, n9722, n9723, n9724, n9725,
    n9726, n9727, n9728, n9729, n9730, n9731,
    n9732, n9733, n9734, n9735, n9736, n9737,
    n9738, n9739, n9740, n9741, n9742, n9743,
    n9744, n9745, n9746, n9747, n9748, n9749,
    n9750, n9751, n9752, n9753, n9754, n9755,
    n9756, n9757, n9758, n9759, n9760, n9761,
    n9762, n9763, n9764, n9765, n9766, n9767,
    n9768, n9769, n9770, n9771, n9772, n9773,
    n9774, n9775, n9776, n9777, n9778, n9779,
    n9780, n9781, n9782, n9783, n9784, n9785,
    n9786, n9787, n9788, n9789, n9790, n9791,
    n9792, n9793, n9794, n9795, n9796, n9797,
    n9798, n9799, n9800, n9801, n9802, n9803,
    n9804, n9805, n9806, n9807, n9808, n9809,
    n9810, n9811, n9812, n9813, n9814, n9815,
    n9816, n9817, n9818, n9819, n9820, n9821,
    n9822, n9823, n9824, n9825, n9826, n9827,
    n9828, n9829, n9830, n9831, n9832, n9833,
    n9834, n9835, n9836, n9837, n9838, n9839,
    n9840, n9841, n9843, n9844, n9845, n9846,
    n9847, n9848, n9849, n9850, n9851, n9852,
    n9853, n9854, n9855, n9856, n9857, n9858,
    n9859, n9860, n9861, n9862, n9863, n9864,
    n9865, n9866, n9867, n9868, n9869, n9870,
    n9871, n9872, n9873, n9874, n9875, n9876,
    n9877, n9878, n9879, n9880, n9881, n9882,
    n9883, n9884, n9885, n9886, n9887, n9888,
    n9889, n9890, n9891, n9892, n9893, n9894,
    n9895, n9896, n9897, n9898, n9899, n9900,
    n9901, n9902, n9903, n9904, n9905, n9906,
    n9907, n9908, n9909, n9910, n9911, n9912,
    n9913, n9914, n9915, n9916, n9917, n9918,
    n9919, n9920, n9921, n9922, n9923, n9924,
    n9925, n9926, n9927, n9928, n9929, n9930,
    n9931, n9932, n9933, n9934, n9935, n9936,
    n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948,
    n9949, n9950, n9951, n9952, n9953, n9954,
    n9955, n9956, n9957, n9958, n9959, n9960,
    n9961, n9962, n9963, n9964, n9965, n9966,
    n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9990,
    n9991, n9992, n9993, n9994, n9995, n9996,
    n9997, n9998, n9999, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026,
    n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044,
    n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062,
    n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074,
    n10075, n10076, n10077, n10078, n10079, n10080,
    n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092,
    n10093, n10094, n10095, n10096, n10097, n10098,
    n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116,
    n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134,
    n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146,
    n10147, n10148, n10149, n10150, n10151, n10152,
    n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170,
    n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188,
    n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200,
    n10201, n10202, n10203, n10204, n10205, n10206,
    n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218,
    n10219, n10220, n10221, n10222, n10223, n10224,
    n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236,
    n10237, n10238, n10239, n10240, n10241, n10242,
    n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254,
    n10255, n10256, n10257, n10258, n10259, n10260,
    n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272,
    n10273, n10274, n10275, n10276, n10277, n10278,
    n10279, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290,
    n10291, n10292, n10293, n10294, n10295, n10296,
    n10297, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309,
    n10310, n10311, n10312, n10313, n10314, n10315,
    n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327,
    n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345,
    n10346, n10347, n10348, n10349, n10350, n10351,
    n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363,
    n10364, n10365, n10366, n10367, n10368, n10369,
    n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381,
    n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10395, n10396, n10397, n10398, n10399,
    n10400, n10401, n10402, n10403, n10404, n10405,
    n10406, n10407, n10408, n10409, n10410, n10411,
    n10412, n10413, n10414, n10415, n10416, n10417,
    n10418, n10419, n10420, n10421, n10422, n10423,
    n10424, n10425, n10426, n10427, n10428, n10429,
    n10430, n10431, n10432, n10433, n10434, n10435,
    n10436, n10437, n10438, n10439, n10440, n10441,
    n10442, n10443, n10444, n10445, n10446, n10447,
    n10448, n10449, n10450, n10451, n10452, n10453,
    n10454, n10455, n10456, n10457, n10458, n10459,
    n10460, n10461, n10462, n10463, n10464, n10465,
    n10466, n10467, n10468, n10469, n10470, n10471,
    n10472, n10473, n10474, n10475, n10476, n10477,
    n10478, n10479, n10480, n10481, n10482, n10483,
    n10484, n10485, n10486, n10487, n10488, n10489,
    n10490, n10491, n10492, n10493, n10494, n10495,
    n10496, n10497, n10498, n10499, n10500, n10501,
    n10502, n10503, n10504, n10505, n10506, n10507,
    n10508, n10509, n10510, n10511, n10512, n10513,
    n10514, n10515, n10516, n10517, n10518, n10519,
    n10520, n10521, n10522, n10523, n10524, n10525,
    n10526, n10527, n10528, n10529, n10530, n10531,
    n10532, n10533, n10534, n10535, n10536, n10537,
    n10538, n10539, n10540, n10541, n10542, n10543,
    n10544, n10545, n10546, n10547, n10548, n10549,
    n10550, n10551, n10552, n10553, n10554, n10555,
    n10556, n10557, n10558, n10559, n10560, n10561,
    n10562, n10563, n10564, n10565, n10566, n10567,
    n10568, n10569, n10570, n10571, n10572, n10573,
    n10574, n10575, n10576, n10577, n10578, n10579,
    n10580, n10581, n10582, n10583, n10584, n10585,
    n10586, n10587, n10588, n10589, n10590, n10591,
    n10592, n10593, n10594, n10595, n10596, n10597,
    n10598, n10599, n10600, n10601, n10602, n10603,
    n10604, n10605, n10606, n10607, n10608, n10609,
    n10610, n10611, n10612, n10613, n10614, n10615,
    n10616, n10617, n10618, n10619, n10620, n10621,
    n10622, n10623, n10624, n10625, n10626, n10627,
    n10628, n10629, n10630, n10631, n10632, n10633,
    n10634, n10635, n10636, n10637, n10638, n10639,
    n10640, n10641, n10642, n10643, n10644, n10645,
    n10646, n10647, n10648, n10649, n10650, n10651,
    n10652, n10653, n10654, n10655, n10656, n10657,
    n10658, n10659, n10660, n10661, n10662, n10663,
    n10664, n10665, n10666, n10667, n10668, n10669,
    n10670, n10671, n10672, n10673, n10674, n10675,
    n10676, n10677, n10678, n10679, n10680, n10681,
    n10682, n10683, n10684, n10685, n10686, n10687,
    n10688, n10689, n10690, n10691, n10692, n10693,
    n10694, n10695, n10696, n10697, n10698, n10699,
    n10700, n10701, n10702, n10703, n10704, n10705,
    n10706, n10707, n10708, n10709, n10710, n10711,
    n10712, n10713, n10714, n10715, n10716, n10717,
    n10718, n10719, n10720, n10721, n10722, n10723,
    n10724, n10725, n10726, n10727, n10728, n10729,
    n10730, n10731, n10732, n10733, n10734, n10735,
    n10736, n10737, n10738, n10739, n10740, n10741,
    n10742, n10743, n10744, n10745, n10746, n10747,
    n10748, n10749, n10750, n10751, n10752, n10753,
    n10754, n10755, n10756, n10757, n10758, n10759,
    n10760, n10761, n10762, n10763, n10764, n10766,
    n10767, n10768, n10769, n10770, n10771, n10772,
    n10773, n10774, n10775, n10776, n10777, n10778,
    n10779, n10780, n10781, n10782, n10783, n10784,
    n10785, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838,
    n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850,
    n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868,
    n10869, n10870, n10871, n10872, n10873, n10874,
    n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886,
    n10887, n10888, n10889, n10890, n10891, n10892,
    n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904,
    n10905, n10906, n10907, n10908, n10909, n10910,
    n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922,
    n10923, n10924, n10925, n10926, n10927, n10928,
    n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940,
    n10941, n10942, n10943, n10944, n10945, n10946,
    n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958,
    n10959, n10960, n10961, n10962, n10963, n10964,
    n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10981, n10982,
    n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994,
    n10995, n10996, n10997, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012,
    n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030,
    n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048,
    n11049, n11050, n11051, n11052, n11053, n11054,
    n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066,
    n11067, n11068, n11069, n11070, n11071, n11072,
    n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084,
    n11085, n11086, n11087, n11088, n11089, n11090,
    n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102,
    n11103, n11104, n11105, n11106, n11107, n11108,
    n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120,
    n11121, n11122, n11123, n11124, n11125, n11126,
    n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138,
    n11139, n11140, n11141, n11142, n11143, n11144,
    n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11152, n11153, n11154, n11155, n11156,
    n11157, n11158, n11159, n11160, n11161, n11162,
    n11163, n11164, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174,
    n11175, n11176, n11177, n11178, n11179, n11180,
    n11181, n11182, n11183, n11184, n11185, n11186,
    n11187, n11188, n11189, n11190, n11191, n11192,
    n11193, n11194, n11195, n11196, n11197, n11198,
    n11199, n11200, n11201, n11202, n11203, n11204,
    n11205, n11206, n11207, n11208, n11209, n11210,
    n11211, n11212, n11213, n11214, n11215, n11216,
    n11217, n11218, n11219, n11220, n11221, n11222,
    n11223, n11224, n11225, n11226, n11227, n11228,
    n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240,
    n11241, n11243, n11244, n11245, n11246, n11247,
    n11248, n11249, n11250, n11251, n11252, n11253,
    n11254, n11255, n11256, n11257, n11258, n11259,
    n11260, n11261, n11262, n11263, n11264, n11265,
    n11266, n11267, n11268, n11269, n11270, n11271,
    n11272, n11273, n11274, n11275, n11276, n11277,
    n11278, n11279, n11280, n11281, n11282, n11283,
    n11284, n11285, n11286, n11287, n11288, n11289,
    n11290, n11291, n11292, n11293, n11294, n11295,
    n11296, n11297, n11298, n11299, n11300, n11301,
    n11302, n11303, n11304, n11305, n11306, n11307,
    n11308, n11309, n11310, n11311, n11312, n11313,
    n11314, n11315, n11316, n11317, n11318, n11319,
    n11320, n11321, n11322, n11323, n11324, n11325,
    n11326, n11327, n11328, n11329, n11330, n11331,
    n11332, n11333, n11334, n11335, n11336, n11337,
    n11338, n11339, n11340, n11341, n11342, n11343,
    n11344, n11345, n11346, n11347, n11348, n11349,
    n11350, n11351, n11352, n11353, n11354, n11355,
    n11356, n11357, n11358, n11359, n11360, n11361,
    n11362, n11363, n11364, n11365, n11366, n11367,
    n11368, n11369, n11370, n11371, n11372, n11373,
    n11374, n11375, n11376, n11377, n11378, n11379,
    n11380, n11381, n11382, n11383, n11384, n11385,
    n11386, n11387, n11388, n11389, n11390, n11391,
    n11392, n11393, n11394, n11395, n11396, n11397,
    n11398, n11399, n11400, n11401, n11402, n11403,
    n11404, n11405, n11406, n11407, n11408, n11409,
    n11410, n11411, n11412, n11413, n11414, n11415,
    n11416, n11417, n11418, n11419, n11420, n11421,
    n11422, n11423, n11424, n11425, n11426, n11427,
    n11428, n11429, n11430, n11431, n11432, n11433,
    n11434, n11435, n11436, n11437, n11438, n11439,
    n11440, n11441, n11442, n11443, n11444, n11445,
    n11446, n11447, n11448, n11449, n11450, n11451,
    n11452, n11453, n11454, n11455, n11456, n11457,
    n11458, n11459, n11460, n11461, n11462, n11463,
    n11464, n11465, n11466, n11467, n11468, n11469,
    n11470, n11471, n11472, n11473, n11474, n11475,
    n11476, n11477, n11478, n11479, n11480, n11481,
    n11482, n11483, n11484, n11485, n11486, n11487,
    n11488, n11489, n11490, n11491, n11492, n11493,
    n11494, n11495, n11496, n11497, n11498, n11499,
    n11500, n11501, n11502, n11503, n11504, n11505,
    n11506, n11507, n11508, n11509, n11510, n11511,
    n11512, n11513, n11514, n11515, n11516, n11517,
    n11518, n11519, n11520, n11521, n11522, n11523,
    n11524, n11525, n11526, n11527, n11528, n11529,
    n11530, n11531, n11532, n11533, n11534, n11535,
    n11536, n11537, n11538, n11539, n11540, n11541,
    n11542, n11543, n11544, n11545, n11546, n11547,
    n11548, n11549, n11550, n11551, n11552, n11553,
    n11554, n11555, n11556, n11557, n11558, n11559,
    n11560, n11561, n11562, n11563, n11564, n11565,
    n11566, n11567, n11568, n11569, n11570, n11571,
    n11572, n11573, n11574, n11575, n11576, n11577,
    n11578, n11579, n11580, n11581, n11582, n11583,
    n11584, n11585, n11586, n11587, n11588, n11589,
    n11590, n11591, n11592, n11593, n11594, n11595,
    n11596, n11597, n11598, n11599, n11600, n11601,
    n11602, n11603, n11604, n11605, n11606, n11607,
    n11608, n11609, n11610, n11611, n11612, n11613,
    n11614, n11615, n11616, n11617, n11618, n11619,
    n11620, n11621, n11622, n11623, n11624, n11625,
    n11626, n11627, n11628, n11629, n11630, n11631,
    n11632, n11633, n11634, n11635, n11636, n11637,
    n11638, n11639, n11640, n11641, n11642, n11643,
    n11644, n11645, n11646, n11647, n11648, n11649,
    n11650, n11651, n11652, n11653, n11654, n11655,
    n11656, n11657, n11658, n11659, n11660, n11661,
    n11662, n11663, n11664, n11665, n11666, n11667,
    n11668, n11669, n11670, n11671, n11672, n11673,
    n11674, n11675, n11676, n11677, n11678, n11679,
    n11680, n11681, n11682, n11683, n11684, n11685,
    n11686, n11687, n11688, n11689, n11690, n11691,
    n11692, n11693, n11694, n11695, n11696, n11697,
    n11698, n11699, n11700, n11701, n11702, n11703,
    n11704, n11705, n11706, n11707, n11708, n11709,
    n11710, n11711, n11712, n11713, n11714, n11715,
    n11716, n11717, n11718, n11719, n11720, n11721,
    n11722, n11723, n11724, n11725, n11726, n11727,
    n11728, n11729, n11731, n11732, n11733, n11734,
    n11735, n11736, n11737, n11738, n11739, n11740,
    n11741, n11742, n11743, n11744, n11745, n11746,
    n11747, n11748, n11749, n11750, n11751, n11752,
    n11753, n11754, n11755, n11756, n11757, n11758,
    n11759, n11760, n11761, n11762, n11763, n11764,
    n11765, n11766, n11767, n11768, n11769, n11770,
    n11771, n11772, n11773, n11774, n11775, n11776,
    n11777, n11778, n11779, n11780, n11781, n11782,
    n11783, n11784, n11785, n11786, n11787, n11788,
    n11789, n11790, n11791, n11792, n11793, n11794,
    n11795, n11796, n11797, n11798, n11799, n11800,
    n11801, n11802, n11803, n11804, n11805, n11806,
    n11807, n11808, n11809, n11810, n11811, n11812,
    n11813, n11814, n11815, n11816, n11817, n11818,
    n11819, n11820, n11821, n11822, n11823, n11824,
    n11825, n11826, n11827, n11828, n11829, n11830,
    n11831, n11832, n11833, n11834, n11835, n11836,
    n11837, n11838, n11839, n11840, n11841, n11842,
    n11843, n11844, n11845, n11846, n11847, n11848,
    n11849, n11850, n11851, n11852, n11853, n11854,
    n11855, n11856, n11857, n11858, n11859, n11860,
    n11861, n11862, n11863, n11864, n11865, n11866,
    n11867, n11868, n11869, n11870, n11871, n11872,
    n11873, n11874, n11875, n11876, n11877, n11878,
    n11879, n11880, n11881, n11882, n11883, n11884,
    n11885, n11886, n11887, n11888, n11889, n11890,
    n11891, n11892, n11893, n11894, n11895, n11896,
    n11897, n11898, n11899, n11900, n11901, n11902,
    n11903, n11904, n11905, n11906, n11907, n11908,
    n11909, n11910, n11911, n11912, n11913, n11914,
    n11915, n11916, n11917, n11918, n11919, n11920,
    n11921, n11922, n11923, n11924, n11925, n11926,
    n11927, n11928, n11929, n11930, n11931, n11932,
    n11933, n11934, n11935, n11936, n11937, n11938,
    n11939, n11940, n11941, n11942, n11943, n11944,
    n11945, n11946, n11947, n11948, n11949, n11950,
    n11951, n11952, n11953, n11954, n11955, n11956,
    n11957, n11958, n11959, n11960, n11961, n11962,
    n11963, n11964, n11965, n11966, n11967, n11968,
    n11969, n11970, n11971, n11972, n11973, n11974,
    n11975, n11976, n11977, n11978, n11979, n11980,
    n11981, n11982, n11983, n11984, n11985, n11986,
    n11987, n11988, n11989, n11990, n11991, n11992,
    n11993, n11994, n11995, n11996, n11997, n11998,
    n11999, n12000, n12001, n12002, n12003, n12004,
    n12005, n12006, n12007, n12008, n12009, n12010,
    n12011, n12012, n12013, n12014, n12015, n12016,
    n12017, n12018, n12019, n12020, n12021, n12022,
    n12023, n12024, n12025, n12026, n12027, n12028,
    n12029, n12030, n12031, n12032, n12033, n12034,
    n12035, n12036, n12037, n12038, n12039, n12040,
    n12041, n12042, n12043, n12044, n12045, n12046,
    n12047, n12048, n12049, n12050, n12051, n12052,
    n12053, n12054, n12055, n12056, n12057, n12058,
    n12059, n12060, n12061, n12062, n12063, n12064,
    n12065, n12066, n12067, n12068, n12069, n12070,
    n12071, n12072, n12073, n12074, n12075, n12076,
    n12077, n12078, n12079, n12080, n12081, n12082,
    n12083, n12084, n12085, n12086, n12087, n12088,
    n12089, n12090, n12091, n12092, n12093, n12094,
    n12095, n12096, n12097, n12098, n12099, n12100,
    n12101, n12102, n12103, n12104, n12105, n12106,
    n12107, n12108, n12109, n12110, n12111, n12112,
    n12113, n12114, n12115, n12116, n12117, n12118,
    n12119, n12120, n12121, n12122, n12123, n12124,
    n12125, n12126, n12127, n12128, n12129, n12130,
    n12131, n12132, n12133, n12134, n12135, n12136,
    n12137, n12138, n12139, n12140, n12141, n12142,
    n12143, n12144, n12145, n12146, n12147, n12148,
    n12149, n12150, n12151, n12152, n12153, n12154,
    n12155, n12156, n12157, n12158, n12159, n12160,
    n12161, n12162, n12163, n12164, n12165, n12166,
    n12167, n12168, n12169, n12170, n12171, n12172,
    n12173, n12174, n12175, n12176, n12177, n12178,
    n12179, n12180, n12181, n12182, n12183, n12184,
    n12185, n12186, n12187, n12188, n12189, n12190,
    n12191, n12192, n12193, n12194, n12195, n12196,
    n12197, n12198, n12199, n12200, n12201, n12202,
    n12203, n12204, n12205, n12206, n12207, n12208,
    n12209, n12210, n12211, n12212, n12213, n12214,
    n12215, n12216, n12217, n12218, n12219, n12220,
    n12221, n12222, n12223, n12224, n12225, n12226,
    n12227, n12229, n12230, n12231, n12232, n12233,
    n12234, n12235, n12236, n12237, n12238, n12239,
    n12240, n12241, n12242, n12243, n12244, n12245,
    n12246, n12247, n12248, n12249, n12250, n12251,
    n12252, n12253, n12254, n12255, n12256, n12257,
    n12258, n12259, n12260, n12261, n12262, n12263,
    n12264, n12265, n12266, n12267, n12268, n12269,
    n12270, n12271, n12272, n12273, n12274, n12275,
    n12276, n12277, n12278, n12279, n12280, n12281,
    n12282, n12283, n12284, n12285, n12286, n12287,
    n12288, n12289, n12290, n12291, n12292, n12293,
    n12294, n12295, n12296, n12297, n12298, n12299,
    n12300, n12301, n12302, n12303, n12304, n12305,
    n12306, n12307, n12308, n12309, n12310, n12311,
    n12312, n12313, n12314, n12315, n12316, n12317,
    n12318, n12319, n12320, n12321, n12322, n12323,
    n12324, n12325, n12326, n12327, n12328, n12329,
    n12330, n12331, n12332, n12333, n12334, n12335,
    n12336, n12337, n12338, n12339, n12340, n12341,
    n12342, n12343, n12344, n12345, n12346, n12347,
    n12348, n12349, n12350, n12351, n12352, n12353,
    n12354, n12355, n12356, n12357, n12358, n12359,
    n12360, n12361, n12362, n12363, n12364, n12365,
    n12366, n12367, n12368, n12369, n12370, n12371,
    n12372, n12373, n12374, n12375, n12376, n12377,
    n12378, n12379, n12380, n12381, n12382, n12383,
    n12384, n12385, n12386, n12387, n12388, n12389,
    n12390, n12391, n12392, n12393, n12394, n12395,
    n12396, n12397, n12398, n12399, n12400, n12401,
    n12402, n12403, n12404, n12405, n12406, n12407,
    n12408, n12409, n12410, n12411, n12412, n12413,
    n12414, n12415, n12416, n12417, n12418, n12419,
    n12420, n12421, n12422, n12423, n12424, n12425,
    n12426, n12427, n12428, n12429, n12430, n12431,
    n12432, n12433, n12434, n12435, n12436, n12437,
    n12438, n12439, n12440, n12441, n12442, n12443,
    n12444, n12445, n12446, n12447, n12448, n12449,
    n12450, n12451, n12452, n12453, n12454, n12455,
    n12456, n12457, n12458, n12459, n12460, n12461,
    n12462, n12463, n12464, n12465, n12466, n12467,
    n12468, n12469, n12470, n12471, n12472, n12473,
    n12474, n12475, n12476, n12477, n12478, n12479,
    n12480, n12481, n12482, n12483, n12484, n12485,
    n12486, n12487, n12488, n12489, n12490, n12491,
    n12492, n12493, n12494, n12495, n12496, n12497,
    n12498, n12499, n12500, n12501, n12502, n12503,
    n12504, n12505, n12506, n12507, n12508, n12509,
    n12510, n12511, n12512, n12513, n12514, n12515,
    n12516, n12517, n12518, n12519, n12520, n12521,
    n12522, n12523, n12524, n12525, n12526, n12527,
    n12528, n12529, n12530, n12531, n12532, n12533,
    n12534, n12535, n12536, n12537, n12538, n12539,
    n12540, n12541, n12542, n12543, n12544, n12545,
    n12546, n12547, n12548, n12549, n12550, n12551,
    n12552, n12553, n12554, n12555, n12556, n12557,
    n12558, n12559, n12560, n12561, n12562, n12563,
    n12564, n12565, n12566, n12567, n12568, n12569,
    n12570, n12571, n12572, n12573, n12574, n12575,
    n12576, n12577, n12578, n12579, n12580, n12581,
    n12582, n12583, n12584, n12585, n12586, n12587,
    n12588, n12589, n12590, n12591, n12592, n12593,
    n12594, n12595, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12604, n12605,
    n12606, n12607, n12608, n12609, n12610, n12611,
    n12612, n12613, n12614, n12615, n12616, n12617,
    n12618, n12619, n12620, n12621, n12622, n12623,
    n12624, n12625, n12626, n12627, n12628, n12629,
    n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641,
    n12642, n12643, n12644, n12645, n12646, n12647,
    n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659,
    n12660, n12661, n12662, n12663, n12664, n12665,
    n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677,
    n12678, n12679, n12680, n12681, n12682, n12683,
    n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12691, n12692, n12693, n12694, n12695,
    n12696, n12697, n12698, n12699, n12700, n12701,
    n12702, n12703, n12704, n12705, n12706, n12707,
    n12708, n12709, n12710, n12711, n12712, n12713,
    n12714, n12715, n12716, n12717, n12718, n12719,
    n12720, n12721, n12722, n12723, n12724, n12725,
    n12726, n12727, n12728, n12729, n12730, n12731,
    n12732, n12733, n12734, n12735, n12736, n12738,
    n12739, n12740, n12741, n12742, n12743, n12744,
    n12745, n12746, n12747, n12748, n12749, n12750,
    n12751, n12752, n12753, n12754, n12755, n12756,
    n12757, n12758, n12759, n12760, n12761, n12762,
    n12763, n12764, n12765, n12766, n12767, n12768,
    n12769, n12770, n12771, n12772, n12773, n12774,
    n12775, n12776, n12777, n12778, n12779, n12780,
    n12781, n12782, n12783, n12784, n12785, n12786,
    n12787, n12788, n12789, n12790, n12791, n12792,
    n12793, n12794, n12795, n12796, n12797, n12798,
    n12799, n12800, n12801, n12802, n12803, n12804,
    n12805, n12806, n12807, n12808, n12809, n12810,
    n12811, n12812, n12813, n12814, n12815, n12816,
    n12817, n12818, n12819, n12820, n12821, n12822,
    n12823, n12824, n12825, n12826, n12827, n12828,
    n12829, n12830, n12831, n12832, n12833, n12834,
    n12835, n12836, n12837, n12838, n12839, n12840,
    n12841, n12842, n12843, n12844, n12845, n12846,
    n12847, n12848, n12849, n12850, n12851, n12852,
    n12853, n12854, n12855, n12856, n12857, n12858,
    n12859, n12860, n12861, n12862, n12863, n12864,
    n12865, n12866, n12867, n12868, n12869, n12870,
    n12871, n12872, n12873, n12874, n12875, n12876,
    n12877, n12878, n12879, n12880, n12881, n12882,
    n12883, n12884, n12885, n12886, n12887, n12888,
    n12889, n12890, n12891, n12892, n12893, n12894,
    n12895, n12896, n12897, n12898, n12899, n12900,
    n12901, n12902, n12903, n12904, n12905, n12906,
    n12907, n12908, n12909, n12910, n12911, n12912,
    n12913, n12914, n12915, n12916, n12917, n12918,
    n12919, n12920, n12921, n12922, n12923, n12924,
    n12925, n12926, n12927, n12928, n12929, n12930,
    n12931, n12932, n12933, n12934, n12935, n12936,
    n12937, n12938, n12939, n12940, n12941, n12942,
    n12943, n12944, n12945, n12946, n12947, n12948,
    n12949, n12950, n12951, n12952, n12953, n12954,
    n12955, n12956, n12957, n12958, n12959, n12960,
    n12961, n12962, n12963, n12964, n12965, n12966,
    n12967, n12968, n12969, n12970, n12971, n12972,
    n12973, n12974, n12975, n12976, n12977, n12978,
    n12979, n12980, n12981, n12982, n12983, n12984,
    n12985, n12986, n12987, n12988, n12989, n12990,
    n12991, n12992, n12993, n12994, n12995, n12996,
    n12997, n12998, n12999, n13000, n13001, n13002,
    n13003, n13004, n13005, n13006, n13007, n13008,
    n13009, n13010, n13011, n13012, n13013, n13014,
    n13015, n13016, n13017, n13018, n13019, n13020,
    n13021, n13022, n13023, n13024, n13025, n13026,
    n13027, n13028, n13029, n13030, n13031, n13032,
    n13033, n13034, n13035, n13036, n13037, n13038,
    n13039, n13040, n13041, n13042, n13043, n13044,
    n13045, n13046, n13047, n13048, n13049, n13050,
    n13051, n13052, n13053, n13054, n13055, n13056,
    n13057, n13058, n13059, n13060, n13061, n13062,
    n13063, n13064, n13065, n13066, n13067, n13068,
    n13069, n13070, n13071, n13072, n13073, n13074,
    n13075, n13076, n13077, n13078, n13079, n13080,
    n13081, n13082, n13083, n13084, n13085, n13086,
    n13087, n13088, n13089, n13090, n13091, n13092,
    n13093, n13094, n13095, n13096, n13097, n13098,
    n13099, n13100, n13101, n13102, n13103, n13104,
    n13105, n13106, n13107, n13108, n13109, n13110,
    n13111, n13112, n13113, n13114, n13115, n13116,
    n13117, n13118, n13119, n13120, n13121, n13122,
    n13123, n13124, n13125, n13126, n13127, n13128,
    n13129, n13130, n13131, n13132, n13133, n13134,
    n13135, n13136, n13137, n13138, n13139, n13140,
    n13141, n13142, n13143, n13144, n13145, n13146,
    n13147, n13148, n13149, n13150, n13151, n13152,
    n13153, n13154, n13155, n13156, n13157, n13158,
    n13159, n13160, n13161, n13162, n13163, n13164,
    n13165, n13166, n13167, n13168, n13169, n13170,
    n13171, n13172, n13173, n13174, n13175, n13176,
    n13177, n13178, n13179, n13180, n13181, n13182,
    n13183, n13184, n13185, n13186, n13187, n13188,
    n13189, n13190, n13191, n13192, n13193, n13194,
    n13195, n13196, n13197, n13198, n13199, n13200,
    n13201, n13202, n13203, n13204, n13205, n13206,
    n13207, n13208, n13209, n13210, n13211, n13212,
    n13213, n13214, n13215, n13216, n13217, n13218,
    n13219, n13220, n13221, n13222, n13223, n13224,
    n13225, n13226, n13227, n13228, n13229, n13230,
    n13231, n13232, n13233, n13234, n13235, n13236,
    n13237, n13238, n13239, n13240, n13241, n13242,
    n13243, n13244, n13245, n13246, n13247, n13248,
    n13249, n13250, n13251, n13252, n13253, n13254,
    n13255, n13257, n13258, n13259, n13260, n13261,
    n13262, n13263, n13264, n13265, n13266, n13267,
    n13268, n13269, n13270, n13271, n13272, n13273,
    n13274, n13275, n13276, n13277, n13278, n13279,
    n13280, n13281, n13282, n13283, n13284, n13285,
    n13286, n13287, n13288, n13289, n13290, n13291,
    n13292, n13293, n13294, n13295, n13296, n13297,
    n13298, n13299, n13300, n13301, n13302, n13303,
    n13304, n13305, n13306, n13307, n13308, n13309,
    n13310, n13311, n13312, n13313, n13314, n13315,
    n13316, n13317, n13318, n13319, n13320, n13321,
    n13322, n13323, n13324, n13325, n13326, n13327,
    n13328, n13329, n13330, n13331, n13332, n13333,
    n13334, n13335, n13336, n13337, n13338, n13339,
    n13340, n13341, n13342, n13343, n13344, n13345,
    n13346, n13347, n13348, n13349, n13350, n13351,
    n13352, n13353, n13354, n13355, n13356, n13357,
    n13358, n13359, n13360, n13361, n13362, n13363,
    n13364, n13365, n13366, n13367, n13368, n13369,
    n13370, n13371, n13372, n13373, n13374, n13375,
    n13376, n13377, n13378, n13379, n13380, n13381,
    n13382, n13383, n13384, n13385, n13386, n13387,
    n13388, n13389, n13390, n13391, n13392, n13393,
    n13394, n13395, n13396, n13397, n13398, n13399,
    n13400, n13401, n13402, n13403, n13404, n13405,
    n13406, n13407, n13408, n13409, n13410, n13411,
    n13412, n13413, n13414, n13415, n13416, n13417,
    n13418, n13419, n13420, n13421, n13422, n13423,
    n13424, n13425, n13426, n13427, n13428, n13429,
    n13430, n13431, n13432, n13433, n13434, n13435,
    n13436, n13437, n13438, n13439, n13440, n13441,
    n13442, n13443, n13444, n13445, n13446, n13447,
    n13448, n13449, n13450, n13451, n13452, n13453,
    n13454, n13455, n13456, n13457, n13458, n13459,
    n13460, n13461, n13462, n13463, n13464, n13465,
    n13466, n13467, n13468, n13469, n13470, n13471,
    n13472, n13473, n13474, n13475, n13476, n13477,
    n13478, n13479, n13480, n13481, n13482, n13483,
    n13484, n13485, n13486, n13487, n13488, n13489,
    n13490, n13491, n13492, n13493, n13494, n13495,
    n13496, n13497, n13498, n13499, n13500, n13501,
    n13502, n13503, n13504, n13505, n13506, n13507,
    n13508, n13509, n13510, n13511, n13512, n13513,
    n13514, n13515, n13516, n13517, n13518, n13519,
    n13520, n13521, n13522, n13523, n13524, n13525,
    n13526, n13527, n13528, n13529, n13530, n13531,
    n13532, n13533, n13534, n13535, n13536, n13537,
    n13538, n13539, n13540, n13541, n13542, n13543,
    n13544, n13545, n13546, n13547, n13548, n13549,
    n13550, n13551, n13552, n13553, n13554, n13555,
    n13556, n13557, n13558, n13559, n13560, n13561,
    n13562, n13563, n13564, n13565, n13566, n13567,
    n13568, n13569, n13570, n13571, n13572, n13573,
    n13574, n13575, n13576, n13577, n13578, n13579,
    n13580, n13581, n13582, n13583, n13584, n13585,
    n13586, n13587, n13588, n13589, n13590, n13591,
    n13592, n13593, n13594, n13595, n13596, n13597,
    n13598, n13599, n13600, n13601, n13602, n13603,
    n13604, n13605, n13606, n13607, n13608, n13609,
    n13610, n13611, n13612, n13613, n13614, n13615,
    n13616, n13617, n13618, n13619, n13620, n13621,
    n13622, n13623, n13624, n13625, n13626, n13627,
    n13628, n13629, n13630, n13631, n13632, n13633,
    n13634, n13635, n13636, n13637, n13638, n13639,
    n13640, n13641, n13642, n13643, n13644, n13645,
    n13646, n13647, n13648, n13649, n13650, n13651,
    n13652, n13653, n13654, n13655, n13656, n13657,
    n13658, n13659, n13660, n13661, n13662, n13663,
    n13664, n13665, n13666, n13667, n13668, n13669,
    n13670, n13671, n13672, n13673, n13674, n13675,
    n13676, n13677, n13678, n13679, n13680, n13681,
    n13682, n13683, n13684, n13685, n13686, n13687,
    n13688, n13689, n13690, n13691, n13692, n13693,
    n13694, n13695, n13696, n13697, n13698, n13699,
    n13700, n13701, n13702, n13703, n13704, n13705,
    n13706, n13707, n13708, n13709, n13710, n13711,
    n13712, n13713, n13714, n13715, n13716, n13717,
    n13718, n13719, n13720, n13721, n13722, n13723,
    n13724, n13725, n13726, n13727, n13728, n13729,
    n13730, n13731, n13732, n13733, n13734, n13735,
    n13736, n13737, n13738, n13739, n13740, n13741,
    n13742, n13743, n13744, n13745, n13746, n13747,
    n13748, n13749, n13750, n13751, n13752, n13753,
    n13754, n13755, n13756, n13757, n13758, n13759,
    n13760, n13761, n13762, n13763, n13764, n13765,
    n13766, n13767, n13768, n13769, n13770, n13771,
    n13772, n13773, n13774, n13775, n13776, n13777,
    n13778, n13779, n13780, n13781, n13782, n13783,
    n13784, n13785, n13787, n13788, n13789, n13790,
    n13791, n13792, n13793, n13794, n13795, n13796,
    n13797, n13798, n13799, n13800, n13801, n13802,
    n13803, n13804, n13805, n13806, n13807, n13808,
    n13809, n13810, n13811, n13812, n13813, n13814,
    n13815, n13816, n13817, n13818, n13819, n13820,
    n13821, n13822, n13823, n13824, n13825, n13826,
    n13827, n13828, n13829, n13830, n13831, n13832,
    n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844,
    n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13862,
    n13863, n13864, n13865, n13866, n13867, n13868,
    n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880,
    n13881, n13882, n13883, n13884, n13885, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892,
    n13893, n13894, n13895, n13896, n13897, n13898,
    n13899, n13900, n13901, n13902, n13903, n13904,
    n13905, n13906, n13907, n13908, n13909, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916,
    n13917, n13918, n13919, n13920, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928,
    n13929, n13930, n13931, n13932, n13933, n13934,
    n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952,
    n13953, n13954, n13955, n13956, n13957, n13958,
    n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970,
    n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988,
    n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006,
    n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14041, n14042,
    n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054,
    n14055, n14056, n14057, n14058, n14059, n14060,
    n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078,
    n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14095, n14096,
    n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108,
    n14109, n14110, n14111, n14112, n14113, n14114,
    n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126,
    n14127, n14128, n14129, n14130, n14131, n14132,
    n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144,
    n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162,
    n14163, n14164, n14165, n14166, n14167, n14168,
    n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180,
    n14181, n14182, n14183, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198,
    n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216,
    n14217, n14218, n14219, n14220, n14221, n14222,
    n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240,
    n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252,
    n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14327, n14328, n14329, n14330, n14331,
    n14332, n14333, n14334, n14335, n14336, n14337,
    n14338, n14339, n14340, n14341, n14342, n14343,
    n14344, n14345, n14346, n14347, n14348, n14349,
    n14350, n14351, n14352, n14353, n14354, n14355,
    n14356, n14357, n14358, n14359, n14360, n14361,
    n14362, n14363, n14364, n14365, n14366, n14367,
    n14368, n14369, n14370, n14371, n14372, n14373,
    n14374, n14375, n14376, n14377, n14378, n14379,
    n14380, n14381, n14382, n14383, n14384, n14385,
    n14386, n14387, n14388, n14389, n14390, n14391,
    n14392, n14393, n14394, n14395, n14396, n14397,
    n14398, n14399, n14400, n14401, n14402, n14403,
    n14404, n14405, n14406, n14407, n14408, n14409,
    n14410, n14411, n14412, n14413, n14414, n14415,
    n14416, n14417, n14418, n14419, n14420, n14421,
    n14422, n14423, n14424, n14425, n14426, n14427,
    n14428, n14429, n14430, n14431, n14432, n14433,
    n14434, n14435, n14436, n14437, n14438, n14439,
    n14440, n14441, n14442, n14443, n14444, n14445,
    n14446, n14447, n14448, n14449, n14450, n14451,
    n14452, n14453, n14454, n14455, n14456, n14457,
    n14458, n14459, n14460, n14461, n14462, n14463,
    n14464, n14465, n14466, n14467, n14468, n14469,
    n14470, n14471, n14472, n14473, n14474, n14475,
    n14476, n14477, n14478, n14479, n14480, n14481,
    n14482, n14483, n14484, n14485, n14486, n14487,
    n14488, n14489, n14490, n14491, n14492, n14493,
    n14494, n14495, n14496, n14497, n14498, n14499,
    n14500, n14501, n14502, n14503, n14504, n14505,
    n14506, n14507, n14508, n14509, n14510, n14511,
    n14512, n14513, n14514, n14515, n14516, n14517,
    n14518, n14519, n14520, n14521, n14522, n14523,
    n14524, n14525, n14526, n14527, n14528, n14529,
    n14530, n14531, n14532, n14533, n14534, n14535,
    n14536, n14537, n14538, n14539, n14540, n14541,
    n14542, n14543, n14544, n14545, n14546, n14547,
    n14548, n14549, n14550, n14551, n14552, n14553,
    n14554, n14555, n14556, n14557, n14558, n14559,
    n14560, n14561, n14562, n14563, n14564, n14565,
    n14566, n14567, n14568, n14569, n14570, n14571,
    n14572, n14573, n14574, n14575, n14576, n14577,
    n14578, n14579, n14580, n14581, n14582, n14583,
    n14584, n14585, n14586, n14587, n14588, n14589,
    n14590, n14591, n14592, n14593, n14594, n14595,
    n14596, n14597, n14598, n14599, n14600, n14601,
    n14602, n14603, n14604, n14605, n14606, n14607,
    n14608, n14609, n14610, n14611, n14612, n14613,
    n14614, n14615, n14616, n14617, n14618, n14619,
    n14620, n14621, n14622, n14623, n14624, n14625,
    n14626, n14627, n14628, n14629, n14630, n14631,
    n14632, n14633, n14634, n14635, n14636, n14637,
    n14638, n14639, n14640, n14641, n14642, n14643,
    n14644, n14645, n14646, n14647, n14648, n14649,
    n14650, n14651, n14652, n14653, n14654, n14655,
    n14656, n14657, n14658, n14659, n14660, n14661,
    n14662, n14663, n14664, n14665, n14666, n14667,
    n14668, n14669, n14670, n14671, n14672, n14673,
    n14674, n14675, n14676, n14677, n14678, n14679,
    n14680, n14681, n14682, n14683, n14684, n14685,
    n14686, n14687, n14688, n14689, n14690, n14691,
    n14692, n14693, n14694, n14695, n14696, n14697,
    n14698, n14699, n14700, n14701, n14702, n14703,
    n14704, n14705, n14706, n14707, n14708, n14709,
    n14710, n14711, n14712, n14713, n14714, n14715,
    n14716, n14717, n14718, n14719, n14720, n14721,
    n14722, n14723, n14724, n14725, n14726, n14727,
    n14728, n14729, n14730, n14731, n14732, n14733,
    n14734, n14735, n14736, n14737, n14738, n14739,
    n14740, n14741, n14742, n14743, n14744, n14745,
    n14746, n14747, n14748, n14749, n14750, n14751,
    n14752, n14753, n14754, n14755, n14756, n14757,
    n14758, n14759, n14760, n14761, n14762, n14763,
    n14764, n14765, n14766, n14767, n14768, n14769,
    n14770, n14771, n14772, n14773, n14774, n14775,
    n14776, n14777, n14778, n14779, n14780, n14781,
    n14782, n14783, n14784, n14785, n14786, n14787,
    n14788, n14789, n14790, n14791, n14792, n14793,
    n14794, n14795, n14796, n14797, n14798, n14799,
    n14800, n14801, n14802, n14803, n14804, n14805,
    n14806, n14807, n14808, n14809, n14810, n14811,
    n14812, n14813, n14814, n14815, n14816, n14817,
    n14818, n14819, n14820, n14821, n14822, n14823,
    n14824, n14825, n14826, n14827, n14828, n14829,
    n14830, n14831, n14832, n14833, n14834, n14835,
    n14836, n14837, n14838, n14839, n14840, n14841,
    n14842, n14843, n14844, n14845, n14846, n14847,
    n14848, n14849, n14850, n14851, n14852, n14853,
    n14854, n14855, n14856, n14857, n14858, n14859,
    n14860, n14861, n14862, n14863, n14864, n14865,
    n14866, n14867, n14868, n14869, n14870, n14871,
    n14872, n14873, n14874, n14875, n14876, n14878,
    n14879, n14880, n14881, n14882, n14883, n14884,
    n14885, n14886, n14887, n14888, n14889, n14890,
    n14891, n14892, n14893, n14894, n14895, n14896,
    n14897, n14898, n14899, n14900, n14901, n14902,
    n14903, n14904, n14905, n14906, n14907, n14908,
    n14909, n14910, n14911, n14912, n14913, n14914,
    n14915, n14916, n14917, n14918, n14919, n14920,
    n14921, n14922, n14923, n14924, n14925, n14926,
    n14927, n14928, n14929, n14930, n14931, n14932,
    n14933, n14934, n14935, n14936, n14937, n14938,
    n14939, n14940, n14941, n14942, n14943, n14944,
    n14945, n14946, n14947, n14948, n14949, n14950,
    n14951, n14952, n14953, n14954, n14955, n14956,
    n14957, n14958, n14959, n14960, n14961, n14962,
    n14963, n14964, n14965, n14966, n14967, n14968,
    n14969, n14970, n14971, n14972, n14973, n14974,
    n14975, n14976, n14977, n14978, n14979, n14980,
    n14981, n14982, n14983, n14984, n14985, n14986,
    n14987, n14988, n14989, n14990, n14991, n14992,
    n14993, n14994, n14995, n14996, n14997, n14998,
    n14999, n15000, n15001, n15002, n15003, n15004,
    n15005, n15006, n15007, n15008, n15009, n15010,
    n15011, n15012, n15013, n15014, n15015, n15016,
    n15017, n15018, n15019, n15020, n15021, n15022,
    n15023, n15024, n15025, n15026, n15027, n15028,
    n15029, n15030, n15031, n15032, n15033, n15034,
    n15035, n15036, n15037, n15038, n15039, n15040,
    n15041, n15042, n15043, n15044, n15045, n15046,
    n15047, n15048, n15049, n15050, n15051, n15052,
    n15053, n15054, n15055, n15056, n15057, n15058,
    n15059, n15060, n15061, n15062, n15063, n15064,
    n15065, n15066, n15067, n15068, n15069, n15070,
    n15071, n15072, n15073, n15074, n15075, n15076,
    n15077, n15078, n15079, n15080, n15081, n15082,
    n15083, n15084, n15085, n15086, n15087, n15088,
    n15089, n15090, n15091, n15092, n15093, n15094,
    n15095, n15096, n15097, n15098, n15099, n15100,
    n15101, n15102, n15103, n15104, n15105, n15106,
    n15107, n15108, n15109, n15110, n15111, n15112,
    n15113, n15114, n15115, n15116, n15117, n15118,
    n15119, n15120, n15121, n15122, n15123, n15124,
    n15125, n15126, n15127, n15128, n15129, n15130,
    n15131, n15132, n15133, n15134, n15135, n15136,
    n15137, n15138, n15139, n15140, n15141, n15142,
    n15143, n15144, n15145, n15146, n15147, n15148,
    n15149, n15150, n15151, n15152, n15153, n15154,
    n15155, n15156, n15157, n15158, n15159, n15160,
    n15161, n15162, n15163, n15164, n15165, n15166,
    n15167, n15168, n15169, n15170, n15171, n15172,
    n15173, n15174, n15175, n15176, n15177, n15178,
    n15179, n15180, n15181, n15182, n15183, n15184,
    n15185, n15186, n15187, n15188, n15189, n15190,
    n15191, n15192, n15193, n15194, n15195, n15196,
    n15197, n15198, n15199, n15200, n15201, n15202,
    n15203, n15204, n15205, n15206, n15207, n15208,
    n15209, n15210, n15211, n15212, n15213, n15214,
    n15215, n15216, n15217, n15218, n15219, n15220,
    n15221, n15222, n15223, n15224, n15225, n15226,
    n15227, n15228, n15229, n15230, n15231, n15232,
    n15233, n15234, n15235, n15236, n15237, n15238,
    n15239, n15240, n15241, n15242, n15243, n15244,
    n15245, n15246, n15247, n15248, n15249, n15250,
    n15251, n15252, n15253, n15254, n15255, n15256,
    n15257, n15258, n15259, n15260, n15261, n15262,
    n15263, n15264, n15265, n15266, n15267, n15268,
    n15269, n15270, n15271, n15272, n15273, n15274,
    n15275, n15276, n15277, n15278, n15279, n15280,
    n15281, n15282, n15283, n15284, n15285, n15286,
    n15287, n15288, n15289, n15290, n15291, n15292,
    n15293, n15294, n15295, n15296, n15297, n15298,
    n15299, n15300, n15301, n15302, n15303, n15304,
    n15305, n15306, n15307, n15308, n15309, n15310,
    n15311, n15312, n15313, n15314, n15315, n15316,
    n15317, n15318, n15319, n15320, n15321, n15322,
    n15323, n15324, n15325, n15326, n15327, n15328,
    n15329, n15330, n15331, n15332, n15333, n15334,
    n15335, n15336, n15337, n15338, n15339, n15340,
    n15341, n15342, n15343, n15344, n15345, n15346,
    n15347, n15348, n15349, n15350, n15351, n15352,
    n15353, n15354, n15355, n15356, n15357, n15358,
    n15359, n15360, n15361, n15362, n15363, n15364,
    n15365, n15366, n15367, n15368, n15369, n15370,
    n15371, n15372, n15373, n15374, n15375, n15376,
    n15377, n15378, n15379, n15380, n15381, n15382,
    n15383, n15384, n15385, n15386, n15387, n15388,
    n15389, n15390, n15391, n15392, n15393, n15394,
    n15395, n15396, n15397, n15398, n15399, n15400,
    n15401, n15402, n15403, n15404, n15405, n15406,
    n15407, n15408, n15409, n15410, n15411, n15412,
    n15413, n15414, n15415, n15416, n15417, n15418,
    n15419, n15420, n15421, n15422, n15423, n15424,
    n15425, n15426, n15427, n15428, n15429, n15430,
    n15431, n15432, n15433, n15434, n15435, n15436,
    n15437, n15439, n15440, n15441, n15442, n15443,
    n15444, n15445, n15446, n15447, n15448, n15449,
    n15450, n15451, n15452, n15453, n15454, n15455,
    n15456, n15457, n15458, n15459, n15460, n15461,
    n15462, n15463, n15464, n15465, n15466, n15467,
    n15468, n15469, n15470, n15471, n15472, n15473,
    n15474, n15475, n15476, n15477, n15478, n15479,
    n15480, n15481, n15482, n15483, n15484, n15485,
    n15486, n15487, n15488, n15489, n15490, n15491,
    n15492, n15493, n15494, n15495, n15496, n15497,
    n15498, n15499, n15500, n15501, n15502, n15503,
    n15504, n15505, n15506, n15507, n15508, n15509,
    n15510, n15511, n15512, n15513, n15514, n15515,
    n15516, n15517, n15518, n15519, n15520, n15521,
    n15522, n15523, n15524, n15525, n15526, n15527,
    n15528, n15529, n15530, n15531, n15532, n15533,
    n15534, n15535, n15536, n15537, n15538, n15539,
    n15540, n15541, n15542, n15543, n15544, n15545,
    n15546, n15547, n15548, n15549, n15550, n15551,
    n15552, n15553, n15554, n15555, n15556, n15557,
    n15558, n15559, n15560, n15561, n15562, n15563,
    n15564, n15565, n15566, n15567, n15568, n15569,
    n15570, n15571, n15572, n15573, n15574, n15575,
    n15576, n15577, n15578, n15579, n15580, n15581,
    n15582, n15583, n15584, n15585, n15586, n15587,
    n15588, n15589, n15590, n15591, n15592, n15593,
    n15594, n15595, n15596, n15597, n15598, n15599,
    n15600, n15601, n15602, n15603, n15604, n15605,
    n15606, n15607, n15608, n15609, n15610, n15611,
    n15612, n15613, n15614, n15615, n15616, n15617,
    n15618, n15619, n15620, n15621, n15622, n15623,
    n15624, n15625, n15626, n15627, n15628, n15629,
    n15630, n15631, n15632, n15633, n15634, n15635,
    n15636, n15637, n15638, n15639, n15640, n15641,
    n15642, n15643, n15644, n15645, n15646, n15647,
    n15648, n15649, n15650, n15651, n15652, n15653,
    n15654, n15655, n15656, n15657, n15658, n15659,
    n15660, n15661, n15662, n15663, n15664, n15665,
    n15666, n15667, n15668, n15669, n15670, n15671,
    n15672, n15673, n15674, n15675, n15676, n15677,
    n15678, n15679, n15680, n15681, n15682, n15683,
    n15684, n15685, n15686, n15687, n15688, n15689,
    n15690, n15691, n15692, n15693, n15694, n15695,
    n15696, n15697, n15698, n15699, n15700, n15701,
    n15702, n15703, n15704, n15705, n15706, n15707,
    n15708, n15709, n15710, n15711, n15712, n15713,
    n15714, n15715, n15716, n15717, n15718, n15719,
    n15720, n15721, n15722, n15723, n15724, n15725,
    n15726, n15727, n15728, n15729, n15730, n15731,
    n15732, n15733, n15734, n15735, n15736, n15737,
    n15738, n15739, n15740, n15741, n15742, n15743,
    n15744, n15745, n15746, n15747, n15748, n15749,
    n15750, n15751, n15752, n15753, n15754, n15755,
    n15756, n15757, n15758, n15759, n15760, n15761,
    n15762, n15763, n15764, n15765, n15766, n15767,
    n15768, n15769, n15770, n15771, n15772, n15773,
    n15774, n15775, n15776, n15777, n15778, n15779,
    n15780, n15781, n15782, n15783, n15784, n15785,
    n15786, n15787, n15788, n15789, n15790, n15791,
    n15792, n15793, n15794, n15795, n15796, n15797,
    n15798, n15799, n15800, n15801, n15802, n15803,
    n15804, n15805, n15806, n15807, n15808, n15809,
    n15810, n15811, n15812, n15813, n15814, n15815,
    n15816, n15817, n15818, n15819, n15820, n15821,
    n15822, n15823, n15824, n15825, n15826, n15827,
    n15828, n15829, n15830, n15831, n15832, n15833,
    n15834, n15835, n15836, n15837, n15838, n15839,
    n15840, n15841, n15842, n15843, n15844, n15845,
    n15846, n15847, n15848, n15849, n15850, n15851,
    n15852, n15853, n15854, n15855, n15856, n15857,
    n15858, n15859, n15860, n15861, n15862, n15863,
    n15864, n15865, n15866, n15867, n15868, n15869,
    n15870, n15871, n15872, n15873, n15874, n15875,
    n15876, n15877, n15878, n15879, n15880, n15881,
    n15882, n15883, n15884, n15885, n15886, n15887,
    n15888, n15889, n15890, n15891, n15892, n15893,
    n15894, n15895, n15896, n15897, n15898, n15899,
    n15900, n15901, n15902, n15903, n15904, n15905,
    n15906, n15907, n15908, n15909, n15910, n15911,
    n15912, n15913, n15914, n15915, n15916, n15917,
    n15918, n15919, n15920, n15921, n15922, n15923,
    n15924, n15925, n15926, n15927, n15928, n15929,
    n15930, n15931, n15932, n15933, n15934, n15935,
    n15936, n15937, n15938, n15939, n15940, n15941,
    n15942, n15943, n15944, n15945, n15946, n15947,
    n15948, n15949, n15950, n15951, n15952, n15953,
    n15954, n15955, n15956, n15957, n15958, n15959,
    n15960, n15961, n15962, n15963, n15964, n15965,
    n15966, n15967, n15968, n15969, n15970, n15971,
    n15972, n15973, n15974, n15975, n15976, n15977,
    n15978, n15979, n15980, n15981, n15982, n15983,
    n15984, n15985, n15986, n15987, n15988, n15989,
    n15990, n15991, n15992, n15993, n15994, n15995,
    n15996, n15997, n15998, n15999, n16000, n16001,
    n16002, n16003, n16004, n16005, n16006, n16007,
    n16008, n16009, n16011, n16012, n16013, n16014,
    n16015, n16016, n16017, n16018, n16019, n16020,
    n16021, n16022, n16023, n16024, n16025, n16026,
    n16027, n16028, n16029, n16030, n16031, n16032,
    n16033, n16034, n16035, n16036, n16037, n16038,
    n16039, n16040, n16041, n16042, n16043, n16044,
    n16045, n16046, n16047, n16048, n16049, n16050,
    n16051, n16052, n16053, n16054, n16055, n16056,
    n16057, n16058, n16059, n16060, n16061, n16062,
    n16063, n16064, n16065, n16066, n16067, n16068,
    n16069, n16070, n16071, n16072, n16073, n16074,
    n16075, n16076, n16077, n16078, n16079, n16080,
    n16081, n16082, n16083, n16084, n16085, n16086,
    n16087, n16088, n16089, n16090, n16091, n16092,
    n16093, n16094, n16095, n16096, n16097, n16098,
    n16099, n16100, n16101, n16102, n16103, n16104,
    n16105, n16106, n16107, n16108, n16109, n16110,
    n16111, n16112, n16113, n16114, n16115, n16116,
    n16117, n16118, n16119, n16120, n16121, n16122,
    n16123, n16124, n16125, n16126, n16127, n16128,
    n16129, n16130, n16131, n16132, n16133, n16134,
    n16135, n16136, n16137, n16138, n16139, n16140,
    n16141, n16142, n16143, n16144, n16145, n16146,
    n16147, n16148, n16149, n16150, n16151, n16152,
    n16153, n16154, n16155, n16156, n16157, n16158,
    n16159, n16160, n16161, n16162, n16163, n16164,
    n16165, n16166, n16167, n16168, n16169, n16170,
    n16171, n16172, n16173, n16174, n16175, n16176,
    n16177, n16178, n16179, n16180, n16181, n16182,
    n16183, n16184, n16185, n16186, n16187, n16188,
    n16189, n16190, n16191, n16192, n16193, n16194,
    n16195, n16196, n16197, n16198, n16199, n16200,
    n16201, n16202, n16203, n16204, n16205, n16206,
    n16207, n16208, n16209, n16210, n16211, n16212,
    n16213, n16214, n16215, n16216, n16217, n16218,
    n16219, n16220, n16221, n16222, n16223, n16224,
    n16225, n16226, n16227, n16228, n16229, n16230,
    n16231, n16232, n16233, n16234, n16235, n16236,
    n16237, n16238, n16239, n16240, n16241, n16242,
    n16243, n16244, n16245, n16246, n16247, n16248,
    n16249, n16250, n16251, n16252, n16253, n16254,
    n16255, n16256, n16257, n16258, n16259, n16260,
    n16261, n16262, n16263, n16264, n16265, n16266,
    n16267, n16268, n16269, n16270, n16271, n16272,
    n16273, n16274, n16275, n16276, n16277, n16278,
    n16279, n16280, n16281, n16282, n16283, n16284,
    n16285, n16286, n16287, n16288, n16289, n16290,
    n16291, n16292, n16293, n16294, n16295, n16296,
    n16297, n16298, n16299, n16300, n16301, n16302,
    n16303, n16304, n16305, n16306, n16307, n16308,
    n16309, n16310, n16311, n16312, n16313, n16314,
    n16315, n16316, n16317, n16318, n16319, n16320,
    n16321, n16322, n16323, n16324, n16325, n16326,
    n16327, n16328, n16329, n16330, n16331, n16332,
    n16333, n16334, n16335, n16336, n16337, n16338,
    n16339, n16340, n16341, n16342, n16343, n16344,
    n16345, n16346, n16347, n16348, n16349, n16350,
    n16351, n16352, n16353, n16354, n16355, n16356,
    n16357, n16358, n16359, n16360, n16361, n16362,
    n16363, n16364, n16365, n16366, n16367, n16368,
    n16369, n16370, n16371, n16372, n16373, n16374,
    n16375, n16376, n16377, n16378, n16379, n16380,
    n16381, n16382, n16383, n16384, n16385, n16386,
    n16387, n16388, n16389, n16390, n16391, n16392,
    n16393, n16394, n16395, n16396, n16397, n16398,
    n16399, n16400, n16401, n16402, n16403, n16404,
    n16405, n16406, n16407, n16408, n16409, n16410,
    n16411, n16412, n16413, n16414, n16415, n16416,
    n16417, n16418, n16419, n16420, n16421, n16422,
    n16423, n16424, n16425, n16426, n16427, n16428,
    n16429, n16430, n16431, n16432, n16433, n16434,
    n16435, n16436, n16437, n16438, n16439, n16440,
    n16441, n16442, n16443, n16444, n16445, n16446,
    n16447, n16448, n16449, n16450, n16451, n16452,
    n16453, n16454, n16455, n16456, n16457, n16458,
    n16459, n16460, n16461, n16462, n16463, n16464,
    n16465, n16466, n16467, n16468, n16469, n16470,
    n16471, n16472, n16473, n16474, n16475, n16476,
    n16477, n16478, n16479, n16480, n16481, n16482,
    n16483, n16484, n16485, n16486, n16487, n16488,
    n16489, n16490, n16491, n16492, n16493, n16494,
    n16495, n16496, n16497, n16498, n16499, n16500,
    n16501, n16502, n16503, n16504, n16505, n16506,
    n16507, n16508, n16509, n16510, n16511, n16512,
    n16513, n16514, n16515, n16516, n16517, n16518,
    n16519, n16520, n16521, n16522, n16523, n16524,
    n16525, n16526, n16527, n16528, n16529, n16530,
    n16531, n16532, n16533, n16534, n16535, n16536,
    n16537, n16538, n16539, n16540, n16541, n16542,
    n16543, n16544, n16545, n16546, n16547, n16548,
    n16549, n16550, n16551, n16552, n16553, n16554,
    n16555, n16556, n16557, n16558, n16559, n16560,
    n16561, n16562, n16563, n16564, n16565, n16566,
    n16567, n16568, n16569, n16570, n16571, n16572,
    n16573, n16574, n16575, n16576, n16577, n16578,
    n16579, n16580, n16581, n16582, n16583, n16584,
    n16585, n16586, n16587, n16588, n16589, n16590,
    n16591, n16593, n16594, n16595, n16596, n16597,
    n16598, n16599, n16600, n16601, n16602, n16603,
    n16604, n16605, n16606, n16607, n16608, n16609,
    n16610, n16611, n16612, n16613, n16614, n16615,
    n16616, n16617, n16618, n16619, n16620, n16621,
    n16622, n16623, n16624, n16625, n16626, n16627,
    n16628, n16629, n16630, n16631, n16632, n16633,
    n16634, n16635, n16636, n16637, n16638, n16639,
    n16640, n16641, n16642, n16643, n16644, n16645,
    n16646, n16647, n16648, n16649, n16650, n16651,
    n16652, n16653, n16654, n16655, n16656, n16657,
    n16658, n16659, n16660, n16661, n16662, n16663,
    n16664, n16665, n16666, n16667, n16668, n16669,
    n16670, n16671, n16672, n16673, n16674, n16675,
    n16676, n16677, n16678, n16679, n16680, n16681,
    n16682, n16683, n16684, n16685, n16686, n16687,
    n16688, n16689, n16690, n16691, n16692, n16693,
    n16694, n16695, n16696, n16697, n16698, n16699,
    n16700, n16701, n16702, n16703, n16704, n16705,
    n16706, n16707, n16708, n16709, n16710, n16711,
    n16712, n16713, n16714, n16715, n16716, n16717,
    n16718, n16719, n16720, n16721, n16722, n16723,
    n16724, n16725, n16726, n16727, n16728, n16729,
    n16730, n16731, n16732, n16733, n16734, n16735,
    n16736, n16737, n16738, n16739, n16740, n16741,
    n16742, n16743, n16744, n16745, n16746, n16747,
    n16748, n16749, n16750, n16751, n16752, n16753,
    n16754, n16755, n16756, n16757, n16758, n16759,
    n16760, n16761, n16762, n16763, n16764, n16765,
    n16766, n16767, n16768, n16769, n16770, n16771,
    n16772, n16773, n16774, n16775, n16776, n16777,
    n16778, n16779, n16780, n16781, n16782, n16783,
    n16784, n16785, n16786, n16787, n16788, n16789,
    n16790, n16791, n16792, n16793, n16794, n16795,
    n16796, n16797, n16798, n16799, n16800, n16801,
    n16802, n16803, n16804, n16805, n16806, n16807,
    n16808, n16809, n16810, n16811, n16812, n16813,
    n16814, n16815, n16816, n16817, n16818, n16819,
    n16820, n16821, n16822, n16823, n16824, n16825,
    n16826, n16827, n16828, n16829, n16830, n16831,
    n16832, n16833, n16834, n16835, n16836, n16837,
    n16838, n16839, n16840, n16841, n16842, n16843,
    n16844, n16845, n16846, n16847, n16848, n16849,
    n16850, n16851, n16852, n16853, n16854, n16855,
    n16856, n16857, n16858, n16859, n16860, n16861,
    n16862, n16863, n16864, n16865, n16866, n16867,
    n16868, n16869, n16870, n16871, n16872, n16873,
    n16874, n16875, n16876, n16877, n16878, n16879,
    n16880, n16881, n16882, n16883, n16884, n16885,
    n16886, n16887, n16888, n16889, n16890, n16891,
    n16892, n16893, n16894, n16895, n16896, n16897,
    n16898, n16899, n16900, n16901, n16902, n16903,
    n16904, n16905, n16906, n16907, n16908, n16909,
    n16910, n16911, n16912, n16913, n16914, n16915,
    n16916, n16917, n16918, n16919, n16920, n16921,
    n16922, n16923, n16924, n16925, n16926, n16927,
    n16928, n16929, n16930, n16931, n16932, n16933,
    n16934, n16935, n16936, n16937, n16938, n16939,
    n16940, n16941, n16942, n16943, n16944, n16945,
    n16946, n16947, n16948, n16949, n16950, n16951,
    n16952, n16953, n16954, n16955, n16956, n16957,
    n16958, n16959, n16960, n16961, n16962, n16963,
    n16964, n16965, n16966, n16967, n16968, n16969,
    n16970, n16971, n16972, n16973, n16974, n16975,
    n16976, n16977, n16978, n16979, n16980, n16981,
    n16982, n16983, n16984, n16985, n16986, n16987,
    n16988, n16989, n16990, n16991, n16992, n16993,
    n16994, n16995, n16996, n16997, n16998, n16999,
    n17000, n17001, n17002, n17003, n17004, n17005,
    n17006, n17007, n17008, n17009, n17010, n17011,
    n17012, n17013, n17014, n17015, n17016, n17017,
    n17018, n17019, n17020, n17021, n17022, n17023,
    n17024, n17025, n17026, n17027, n17028, n17029,
    n17030, n17031, n17032, n17033, n17034, n17035,
    n17036, n17037, n17038, n17039, n17040, n17041,
    n17042, n17043, n17044, n17045, n17046, n17047,
    n17048, n17049, n17050, n17051, n17052, n17053,
    n17054, n17055, n17056, n17057, n17058, n17059,
    n17060, n17061, n17062, n17063, n17064, n17065,
    n17066, n17067, n17068, n17069, n17070, n17071,
    n17072, n17073, n17074, n17075, n17076, n17077,
    n17078, n17079, n17080, n17081, n17082, n17083,
    n17084, n17085, n17086, n17087, n17088, n17089,
    n17090, n17091, n17092, n17093, n17094, n17095,
    n17096, n17097, n17098, n17099, n17100, n17101,
    n17102, n17103, n17104, n17105, n17106, n17107,
    n17108, n17109, n17110, n17111, n17112, n17113,
    n17114, n17115, n17116, n17117, n17118, n17119,
    n17120, n17121, n17122, n17123, n17124, n17125,
    n17126, n17127, n17128, n17129, n17130, n17131,
    n17132, n17133, n17134, n17135, n17136, n17137,
    n17138, n17139, n17140, n17141, n17142, n17143,
    n17144, n17145, n17146, n17147, n17148, n17149,
    n17150, n17151, n17152, n17153, n17154, n17155,
    n17156, n17157, n17158, n17159, n17160, n17161,
    n17162, n17163, n17164, n17165, n17166, n17167,
    n17168, n17169, n17170, n17171, n17172, n17173,
    n17174, n17175, n17176, n17177, n17178, n17179,
    n17180, n17181, n17182, n17183, n17184, n17186,
    n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204,
    n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222,
    n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240,
    n17241, n17242, n17243, n17244, n17245, n17246,
    n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258,
    n17259, n17260, n17261, n17262, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276,
    n17277, n17278, n17279, n17280, n17281, n17282,
    n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294,
    n17295, n17296, n17297, n17298, n17299, n17300,
    n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312,
    n17313, n17314, n17315, n17316, n17317, n17318,
    n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330,
    n17331, n17332, n17333, n17334, n17335, n17336,
    n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348,
    n17349, n17350, n17351, n17352, n17353, n17354,
    n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366,
    n17367, n17368, n17369, n17370, n17371, n17372,
    n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384,
    n17385, n17386, n17387, n17388, n17389, n17390,
    n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402,
    n17403, n17404, n17405, n17406, n17407, n17408,
    n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420,
    n17421, n17422, n17423, n17424, n17425, n17426,
    n17427, n17428, n17429, n17430, n17431, n17432,
    n17433, n17434, n17435, n17436, n17437, n17438,
    n17439, n17440, n17441, n17442, n17443, n17444,
    n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17456,
    n17457, n17458, n17459, n17460, n17461, n17462,
    n17463, n17464, n17465, n17466, n17467, n17468,
    n17469, n17470, n17471, n17472, n17473, n17474,
    n17475, n17476, n17477, n17478, n17479, n17480,
    n17481, n17482, n17483, n17484, n17485, n17486,
    n17487, n17488, n17489, n17490, n17491, n17492,
    n17493, n17494, n17495, n17496, n17497, n17498,
    n17499, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510,
    n17511, n17512, n17513, n17514, n17515, n17516,
    n17517, n17518, n17519, n17520, n17521, n17522,
    n17523, n17524, n17525, n17526, n17527, n17528,
    n17529, n17530, n17531, n17532, n17533, n17534,
    n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546,
    n17547, n17548, n17549, n17550, n17551, n17552,
    n17553, n17554, n17555, n17556, n17557, n17558,
    n17559, n17560, n17561, n17562, n17563, n17564,
    n17565, n17566, n17567, n17568, n17569, n17570,
    n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582,
    n17583, n17584, n17585, n17586, n17587, n17588,
    n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600,
    n17601, n17602, n17603, n17604, n17605, n17606,
    n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618,
    n17619, n17620, n17621, n17622, n17623, n17624,
    n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636,
    n17637, n17638, n17639, n17640, n17641, n17642,
    n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654,
    n17655, n17656, n17657, n17658, n17659, n17660,
    n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672,
    n17673, n17674, n17675, n17676, n17677, n17678,
    n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690,
    n17691, n17692, n17693, n17694, n17695, n17696,
    n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708,
    n17709, n17710, n17711, n17712, n17713, n17714,
    n17715, n17716, n17717, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726,
    n17727, n17728, n17729, n17730, n17731, n17732,
    n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744,
    n17745, n17746, n17747, n17748, n17749, n17750,
    n17751, n17752, n17753, n17754, n17755, n17756,
    n17757, n17758, n17759, n17760, n17761, n17762,
    n17763, n17764, n17765, n17766, n17767, n17768,
    n17769, n17770, n17771, n17772, n17773, n17774,
    n17775, n17776, n17777, n17778, n17779, n17780,
    n17781, n17782, n17783, n17784, n17785, n17786,
    n17787, n17789, n17790, n17791, n17792, n17793,
    n17794, n17795, n17796, n17797, n17798, n17799,
    n17800, n17801, n17802, n17803, n17804, n17805,
    n17806, n17807, n17808, n17809, n17810, n17811,
    n17812, n17813, n17814, n17815, n17816, n17817,
    n17818, n17819, n17820, n17821, n17822, n17823,
    n17824, n17825, n17826, n17827, n17828, n17829,
    n17830, n17831, n17832, n17833, n17834, n17835,
    n17836, n17837, n17838, n17839, n17840, n17841,
    n17842, n17843, n17844, n17845, n17846, n17847,
    n17848, n17849, n17850, n17851, n17852, n17853,
    n17854, n17855, n17856, n17857, n17858, n17859,
    n17860, n17861, n17862, n17863, n17864, n17865,
    n17866, n17867, n17868, n17869, n17870, n17871,
    n17872, n17873, n17874, n17875, n17876, n17877,
    n17878, n17879, n17880, n17881, n17882, n17883,
    n17884, n17885, n17886, n17887, n17888, n17889,
    n17890, n17891, n17892, n17893, n17894, n17895,
    n17896, n17897, n17898, n17899, n17900, n17901,
    n17902, n17903, n17904, n17905, n17906, n17907,
    n17908, n17909, n17910, n17911, n17912, n17913,
    n17914, n17915, n17916, n17917, n17918, n17919,
    n17920, n17921, n17922, n17923, n17924, n17925,
    n17926, n17927, n17928, n17929, n17930, n17931,
    n17932, n17933, n17934, n17935, n17936, n17937,
    n17938, n17939, n17940, n17941, n17942, n17943,
    n17944, n17945, n17946, n17947, n17948, n17949,
    n17950, n17951, n17952, n17953, n17954, n17955,
    n17956, n17957, n17958, n17959, n17960, n17961,
    n17962, n17963, n17964, n17965, n17966, n17967,
    n17968, n17969, n17970, n17971, n17972, n17973,
    n17974, n17975, n17976, n17977, n17978, n17979,
    n17980, n17981, n17982, n17983, n17984, n17985,
    n17986, n17987, n17988, n17989, n17990, n17991,
    n17992, n17993, n17994, n17995, n17996, n17997,
    n17998, n17999, n18000, n18001, n18002, n18003,
    n18004, n18005, n18006, n18007, n18008, n18009,
    n18010, n18011, n18012, n18013, n18014, n18015,
    n18016, n18017, n18018, n18019, n18020, n18021,
    n18022, n18023, n18024, n18025, n18026, n18027,
    n18028, n18029, n18030, n18031, n18032, n18033,
    n18034, n18035, n18036, n18037, n18038, n18039,
    n18040, n18041, n18042, n18043, n18044, n18045,
    n18046, n18047, n18048, n18049, n18050, n18051,
    n18052, n18053, n18054, n18055, n18056, n18057,
    n18058, n18059, n18060, n18061, n18062, n18063,
    n18064, n18065, n18066, n18067, n18068, n18069,
    n18070, n18071, n18072, n18073, n18074, n18075,
    n18076, n18077, n18078, n18079, n18080, n18081,
    n18082, n18083, n18084, n18085, n18086, n18087,
    n18088, n18089, n18090, n18091, n18092, n18093,
    n18094, n18095, n18096, n18097, n18098, n18099,
    n18100, n18101, n18102, n18103, n18104, n18105,
    n18106, n18107, n18108, n18109, n18110, n18111,
    n18112, n18113, n18114, n18115, n18116, n18117,
    n18118, n18119, n18120, n18121, n18122, n18123,
    n18124, n18125, n18126, n18127, n18128, n18129,
    n18130, n18131, n18132, n18133, n18134, n18135,
    n18136, n18137, n18138, n18139, n18140, n18141,
    n18142, n18143, n18144, n18145, n18146, n18147,
    n18148, n18149, n18150, n18151, n18152, n18153,
    n18154, n18155, n18156, n18157, n18158, n18159,
    n18160, n18161, n18162, n18163, n18164, n18165,
    n18166, n18167, n18168, n18169, n18170, n18171,
    n18172, n18173, n18174, n18175, n18176, n18177,
    n18178, n18179, n18180, n18181, n18182, n18183,
    n18184, n18185, n18186, n18187, n18188, n18189,
    n18190, n18191, n18192, n18193, n18194, n18195,
    n18196, n18197, n18198, n18199, n18200, n18201,
    n18202, n18203, n18204, n18205, n18206, n18207,
    n18208, n18209, n18210, n18211, n18212, n18213,
    n18214, n18215, n18216, n18217, n18218, n18219,
    n18220, n18221, n18222, n18223, n18224, n18225,
    n18226, n18227, n18228, n18229, n18230, n18231,
    n18232, n18233, n18234, n18235, n18236, n18237,
    n18238, n18239, n18240, n18241, n18242, n18243,
    n18244, n18245, n18246, n18247, n18248, n18249,
    n18250, n18251, n18252, n18253, n18254, n18255,
    n18256, n18257, n18258, n18259, n18260, n18261,
    n18262, n18263, n18264, n18265, n18266, n18267,
    n18268, n18269, n18270, n18271, n18272, n18273,
    n18274, n18275, n18276, n18277, n18278, n18279,
    n18280, n18281, n18282, n18283, n18284, n18285,
    n18286, n18287, n18288, n18289, n18290, n18291,
    n18292, n18293, n18294, n18295, n18296, n18297,
    n18298, n18299, n18300, n18301, n18302, n18303,
    n18304, n18305, n18306, n18307, n18308, n18309,
    n18310, n18311, n18312, n18313, n18314, n18315,
    n18316, n18317, n18318, n18319, n18320, n18321,
    n18322, n18323, n18324, n18325, n18326, n18327,
    n18328, n18329, n18330, n18331, n18332, n18333,
    n18334, n18335, n18336, n18337, n18338, n18339,
    n18340, n18341, n18342, n18343, n18344, n18345,
    n18346, n18347, n18348, n18349, n18350, n18351,
    n18352, n18353, n18354, n18355, n18356, n18357,
    n18358, n18359, n18360, n18361, n18362, n18363,
    n18364, n18365, n18366, n18367, n18368, n18369,
    n18370, n18371, n18372, n18373, n18374, n18375,
    n18376, n18377, n18378, n18379, n18380, n18381,
    n18382, n18383, n18384, n18385, n18386, n18387,
    n18388, n18389, n18390, n18391, n18392, n18393,
    n18394, n18395, n18396, n18397, n18398, n18399,
    n18401, n18402, n18403, n18404, n18405, n18406,
    n18407, n18408, n18409, n18410, n18411, n18412,
    n18413, n18414, n18415, n18416, n18417, n18418,
    n18419, n18420, n18421, n18422, n18423, n18424,
    n18425, n18426, n18427, n18428, n18429, n18430,
    n18431, n18432, n18433, n18434, n18435, n18436,
    n18437, n18438, n18439, n18440, n18441, n18442,
    n18443, n18444, n18445, n18446, n18447, n18448,
    n18449, n18450, n18451, n18452, n18453, n18454,
    n18455, n18456, n18457, n18458, n18459, n18460,
    n18461, n18462, n18463, n18464, n18465, n18466,
    n18467, n18468, n18469, n18470, n18471, n18472,
    n18473, n18474, n18475, n18476, n18477, n18478,
    n18479, n18480, n18481, n18482, n18483, n18484,
    n18485, n18486, n18487, n18488, n18489, n18490,
    n18491, n18492, n18493, n18494, n18495, n18496,
    n18497, n18498, n18499, n18500, n18501, n18502,
    n18503, n18504, n18505, n18506, n18507, n18508,
    n18509, n18510, n18511, n18512, n18513, n18514,
    n18515, n18516, n18517, n18518, n18519, n18520,
    n18521, n18522, n18523, n18524, n18525, n18526,
    n18527, n18528, n18529, n18530, n18531, n18532,
    n18533, n18534, n18535, n18536, n18537, n18538,
    n18539, n18540, n18541, n18542, n18543, n18544,
    n18545, n18546, n18547, n18548, n18549, n18550,
    n18551, n18552, n18553, n18554, n18555, n18556,
    n18557, n18558, n18559, n18560, n18561, n18562,
    n18563, n18564, n18565, n18566, n18567, n18568,
    n18569, n18570, n18571, n18572, n18573, n18574,
    n18575, n18576, n18577, n18578, n18579, n18580,
    n18581, n18582, n18583, n18584, n18585, n18586,
    n18587, n18588, n18589, n18590, n18591, n18592,
    n18593, n18594, n18595, n18596, n18597, n18598,
    n18599, n18600, n18601, n18602, n18603, n18604,
    n18605, n18606, n18607, n18608, n18609, n18610,
    n18611, n18612, n18613, n18614, n18615, n18616,
    n18617, n18618, n18619, n18620, n18621, n18622,
    n18623, n18624, n18625, n18626, n18627, n18628,
    n18629, n18630, n18631, n18632, n18633, n18634,
    n18635, n18636, n18637, n18638, n18639, n18640,
    n18641, n18642, n18643, n18644, n18645, n18646,
    n18647, n18648, n18649, n18650, n18651, n18652,
    n18653, n18654, n18655, n18656, n18657, n18658,
    n18659, n18660, n18661, n18662, n18663, n18664,
    n18665, n18666, n18667, n18668, n18669, n18670,
    n18671, n18672, n18673, n18674, n18675, n18676,
    n18677, n18678, n18679, n18680, n18681, n18682,
    n18683, n18684, n18685, n18686, n18687, n18688,
    n18689, n18690, n18691, n18692, n18693, n18694,
    n18695, n18696, n18697, n18698, n18699, n18700,
    n18701, n18702, n18703, n18704, n18705, n18706,
    n18707, n18708, n18709, n18710, n18711, n18712,
    n18713, n18714, n18715, n18716, n18717, n18718,
    n18719, n18720, n18721, n18722, n18723, n18724,
    n18725, n18726, n18727, n18728, n18729, n18730,
    n18731, n18732, n18733, n18734, n18735, n18736,
    n18737, n18738, n18739, n18740, n18741, n18742,
    n18743, n18744, n18745, n18746, n18747, n18748,
    n18749, n18750, n18751, n18752, n18753, n18754,
    n18755, n18756, n18757, n18758, n18759, n18760,
    n18761, n18762, n18763, n18764, n18765, n18766,
    n18767, n18768, n18769, n18770, n18771, n18772,
    n18773, n18774, n18775, n18776, n18777, n18778,
    n18779, n18780, n18781, n18782, n18783, n18784,
    n18785, n18786, n18787, n18788, n18789, n18790,
    n18791, n18792, n18793, n18794, n18795, n18796,
    n18797, n18798, n18799, n18800, n18801, n18802,
    n18803, n18804, n18805, n18806, n18807, n18808,
    n18809, n18810, n18811, n18812, n18813, n18814,
    n18815, n18816, n18817, n18818, n18819, n18820,
    n18821, n18822, n18823, n18824, n18825, n18826,
    n18827, n18828, n18829, n18830, n18831, n18832,
    n18833, n18834, n18835, n18836, n18837, n18838,
    n18839, n18840, n18841, n18842, n18843, n18844,
    n18845, n18846, n18847, n18848, n18849, n18850,
    n18851, n18852, n18853, n18854, n18855, n18856,
    n18857, n18858, n18859, n18860, n18861, n18862,
    n18863, n18864, n18865, n18866, n18867, n18868,
    n18869, n18870, n18871, n18872, n18873, n18874,
    n18875, n18876, n18877, n18878, n18879, n18880,
    n18881, n18882, n18883, n18884, n18885, n18886,
    n18887, n18888, n18889, n18890, n18891, n18892,
    n18893, n18894, n18895, n18896, n18897, n18898,
    n18899, n18900, n18901, n18902, n18903, n18904,
    n18905, n18906, n18907, n18908, n18909, n18910,
    n18911, n18912, n18913, n18914, n18915, n18916,
    n18917, n18918, n18919, n18920, n18921, n18922,
    n18923, n18924, n18925, n18926, n18927, n18928,
    n18929, n18930, n18931, n18932, n18933, n18934,
    n18935, n18936, n18937, n18938, n18939, n18940,
    n18941, n18942, n18943, n18944, n18945, n18946,
    n18947, n18948, n18949, n18950, n18951, n18952,
    n18953, n18954, n18955, n18956, n18957, n18958,
    n18959, n18960, n18961, n18962, n18963, n18964,
    n18965, n18966, n18967, n18968, n18969, n18970,
    n18971, n18972, n18973, n18974, n18975, n18976,
    n18977, n18978, n18979, n18980, n18981, n18982,
    n18983, n18984, n18985, n18986, n18987, n18988,
    n18989, n18990, n18991, n18992, n18993, n18994,
    n18995, n18996, n18997, n18998, n18999, n19000,
    n19001, n19002, n19003, n19004, n19005, n19006,
    n19007, n19008, n19009, n19010, n19011, n19012,
    n19013, n19014, n19015, n19016, n19017, n19018,
    n19019, n19020, n19021, n19023, n19024, n19025,
    n19026, n19027, n19028, n19029, n19030, n19031,
    n19032, n19033, n19034, n19035, n19036, n19037,
    n19038, n19039, n19040, n19041, n19042, n19043,
    n19044, n19045, n19046, n19047, n19048, n19049,
    n19050, n19051, n19052, n19053, n19054, n19055,
    n19056, n19057, n19058, n19059, n19060, n19061,
    n19062, n19063, n19064, n19065, n19066, n19067,
    n19068, n19069, n19070, n19071, n19072, n19073,
    n19074, n19075, n19076, n19077, n19078, n19079,
    n19080, n19081, n19082, n19083, n19084, n19085,
    n19086, n19087, n19088, n19089, n19090, n19091,
    n19092, n19093, n19094, n19095, n19096, n19097,
    n19098, n19099, n19100, n19101, n19102, n19103,
    n19104, n19105, n19106, n19107, n19108, n19109,
    n19110, n19111, n19112, n19113, n19114, n19115,
    n19116, n19117, n19118, n19119, n19120, n19121,
    n19122, n19123, n19124, n19125, n19126, n19127,
    n19128, n19129, n19130, n19131, n19132, n19133,
    n19134, n19135, n19136, n19137, n19138, n19139,
    n19140, n19141, n19142, n19143, n19144, n19145,
    n19146, n19147, n19148, n19149, n19150, n19151,
    n19152, n19153, n19154, n19155, n19156, n19157,
    n19158, n19159, n19160, n19161, n19162, n19163,
    n19164, n19165, n19166, n19167, n19168, n19169,
    n19170, n19171, n19172, n19173, n19174, n19175,
    n19176, n19177, n19178, n19179, n19180, n19181,
    n19182, n19183, n19184, n19185, n19186, n19187,
    n19188, n19189, n19190, n19191, n19192, n19193,
    n19194, n19195, n19196, n19197, n19198, n19199,
    n19200, n19201, n19202, n19203, n19204, n19205,
    n19206, n19207, n19208, n19209, n19210, n19211,
    n19212, n19213, n19214, n19215, n19216, n19217,
    n19218, n19219, n19220, n19221, n19222, n19223,
    n19224, n19225, n19226, n19227, n19228, n19229,
    n19230, n19231, n19232, n19233, n19234, n19235,
    n19236, n19237, n19238, n19239, n19240, n19241,
    n19242, n19243, n19244, n19245, n19246, n19247,
    n19248, n19249, n19250, n19251, n19252, n19253,
    n19254, n19255, n19256, n19257, n19258, n19259,
    n19260, n19261, n19262, n19263, n19264, n19265,
    n19266, n19267, n19268, n19269, n19270, n19271,
    n19272, n19273, n19274, n19275, n19276, n19277,
    n19278, n19279, n19280, n19281, n19282, n19283,
    n19284, n19285, n19286, n19287, n19288, n19289,
    n19290, n19291, n19292, n19293, n19294, n19295,
    n19296, n19297, n19298, n19299, n19300, n19301,
    n19302, n19303, n19304, n19305, n19306, n19307,
    n19308, n19309, n19310, n19311, n19312, n19313,
    n19314, n19315, n19316, n19317, n19318, n19319,
    n19320, n19321, n19322, n19323, n19324, n19325,
    n19326, n19327, n19328, n19329, n19330, n19331,
    n19332, n19333, n19334, n19335, n19336, n19337,
    n19338, n19339, n19340, n19341, n19342, n19343,
    n19344, n19345, n19346, n19347, n19348, n19349,
    n19350, n19351, n19352, n19353, n19354, n19355,
    n19356, n19357, n19358, n19359, n19360, n19361,
    n19362, n19363, n19364, n19365, n19366, n19367,
    n19368, n19369, n19370, n19371, n19372, n19373,
    n19374, n19375, n19376, n19377, n19378, n19379,
    n19380, n19381, n19382, n19383, n19384, n19385,
    n19386, n19387, n19388, n19389, n19390, n19391,
    n19392, n19393, n19394, n19395, n19396, n19397,
    n19398, n19399, n19400, n19401, n19402, n19403,
    n19404, n19405, n19406, n19407, n19408, n19409,
    n19410, n19411, n19412, n19413, n19414, n19415,
    n19416, n19417, n19418, n19419, n19420, n19421,
    n19422, n19423, n19424, n19425, n19426, n19427,
    n19428, n19429, n19430, n19431, n19432, n19433,
    n19434, n19435, n19436, n19437, n19438, n19439,
    n19440, n19441, n19442, n19443, n19444, n19445,
    n19446, n19447, n19448, n19449, n19450, n19451,
    n19452, n19453, n19454, n19455, n19456, n19457,
    n19458, n19459, n19460, n19461, n19462, n19463,
    n19464, n19465, n19466, n19467, n19468, n19469,
    n19470, n19471, n19472, n19473, n19474, n19475,
    n19476, n19477, n19478, n19479, n19480, n19481,
    n19482, n19483, n19484, n19485, n19486, n19487,
    n19488, n19489, n19490, n19491, n19492, n19493,
    n19494, n19495, n19496, n19497, n19498, n19499,
    n19500, n19501, n19502, n19503, n19504, n19505,
    n19506, n19507, n19508, n19509, n19510, n19511,
    n19512, n19513, n19514, n19515, n19516, n19517,
    n19518, n19519, n19520, n19521, n19522, n19523,
    n19524, n19525, n19526, n19527, n19528, n19529,
    n19530, n19531, n19532, n19533, n19534, n19535,
    n19536, n19537, n19538, n19539, n19540, n19541,
    n19542, n19543, n19544, n19545, n19546, n19547,
    n19548, n19549, n19550, n19551, n19552, n19553,
    n19554, n19555, n19556, n19557, n19558, n19559,
    n19560, n19561, n19562, n19563, n19564, n19565,
    n19566, n19567, n19568, n19569, n19570, n19571,
    n19572, n19573, n19574, n19575, n19576, n19577,
    n19578, n19579, n19580, n19581, n19582, n19583,
    n19584, n19585, n19586, n19587, n19588, n19589,
    n19590, n19591, n19592, n19593, n19594, n19595,
    n19596, n19597, n19598, n19599, n19600, n19601,
    n19602, n19603, n19604, n19605, n19606, n19607,
    n19608, n19609, n19610, n19611, n19612, n19613,
    n19614, n19615, n19616, n19617, n19618, n19619,
    n19620, n19621, n19622, n19623, n19624, n19625,
    n19626, n19627, n19628, n19629, n19630, n19631,
    n19632, n19633, n19634, n19635, n19636, n19637,
    n19638, n19639, n19640, n19641, n19642, n19643,
    n19644, n19645, n19646, n19647, n19648, n19649,
    n19650, n19651, n19652, n19653, n19654, n19656,
    n19657, n19658, n19659, n19660, n19661, n19662,
    n19663, n19664, n19665, n19666, n19667, n19668,
    n19669, n19670, n19671, n19672, n19673, n19674,
    n19675, n19676, n19677, n19678, n19679, n19680,
    n19681, n19682, n19683, n19684, n19685, n19686,
    n19687, n19688, n19689, n19690, n19691, n19692,
    n19693, n19694, n19695, n19696, n19697, n19698,
    n19699, n19700, n19701, n19702, n19703, n19704,
    n19705, n19706, n19707, n19708, n19709, n19710,
    n19711, n19712, n19713, n19714, n19715, n19716,
    n19717, n19718, n19719, n19720, n19721, n19722,
    n19723, n19724, n19725, n19726, n19727, n19728,
    n19729, n19730, n19731, n19732, n19733, n19734,
    n19735, n19736, n19737, n19738, n19739, n19740,
    n19741, n19742, n19743, n19744, n19745, n19746,
    n19747, n19748, n19749, n19750, n19751, n19752,
    n19753, n19754, n19755, n19756, n19757, n19758,
    n19759, n19760, n19761, n19762, n19763, n19764,
    n19765, n19766, n19767, n19768, n19769, n19770,
    n19771, n19772, n19773, n19774, n19775, n19776,
    n19777, n19778, n19779, n19780, n19781, n19782,
    n19783, n19784, n19785, n19786, n19787, n19788,
    n19789, n19790, n19791, n19792, n19793, n19794,
    n19795, n19796, n19797, n19798, n19799, n19800,
    n19801, n19802, n19803, n19804, n19805, n19806,
    n19807, n19808, n19809, n19810, n19811, n19812,
    n19813, n19814, n19815, n19816, n19817, n19818,
    n19819, n19820, n19821, n19822, n19823, n19824,
    n19825, n19826, n19827, n19828, n19829, n19830,
    n19831, n19832, n19833, n19834, n19835, n19836,
    n19837, n19838, n19839, n19840, n19841, n19842,
    n19843, n19844, n19845, n19846, n19847, n19848,
    n19849, n19850, n19851, n19852, n19853, n19854,
    n19855, n19856, n19857, n19858, n19859, n19860,
    n19861, n19862, n19863, n19864, n19865, n19866,
    n19867, n19868, n19869, n19870, n19871, n19872,
    n19873, n19874, n19875, n19876, n19877, n19878,
    n19879, n19880, n19881, n19882, n19883, n19884,
    n19885, n19886, n19887, n19888, n19889, n19890,
    n19891, n19892, n19893, n19894, n19895, n19896,
    n19897, n19898, n19899, n19900, n19901, n19902,
    n19903, n19904, n19905, n19906, n19907, n19908,
    n19909, n19910, n19911, n19912, n19913, n19914,
    n19915, n19916, n19917, n19918, n19919, n19920,
    n19921, n19922, n19923, n19924, n19925, n19926,
    n19927, n19928, n19929, n19930, n19931, n19932,
    n19933, n19934, n19935, n19936, n19937, n19938,
    n19939, n19940, n19941, n19942, n19943, n19944,
    n19945, n19946, n19947, n19948, n19949, n19950,
    n19951, n19952, n19953, n19954, n19955, n19956,
    n19957, n19958, n19959, n19960, n19961, n19962,
    n19963, n19964, n19965, n19966, n19967, n19968,
    n19969, n19970, n19971, n19972, n19973, n19974,
    n19975, n19976, n19977, n19978, n19979, n19980,
    n19981, n19982, n19983, n19984, n19985, n19986,
    n19987, n19988, n19989, n19990, n19991, n19992,
    n19993, n19994, n19995, n19996, n19997, n19998,
    n19999, n20000, n20001, n20002, n20003, n20004,
    n20005, n20006, n20007, n20008, n20009, n20010,
    n20011, n20012, n20013, n20014, n20015, n20016,
    n20017, n20018, n20019, n20020, n20021, n20022,
    n20023, n20024, n20025, n20026, n20027, n20028,
    n20029, n20030, n20031, n20032, n20033, n20034,
    n20035, n20036, n20037, n20038, n20039, n20040,
    n20041, n20042, n20043, n20044, n20045, n20046,
    n20047, n20048, n20049, n20050, n20051, n20052,
    n20053, n20054, n20055, n20056, n20057, n20058,
    n20059, n20060, n20061, n20062, n20063, n20064,
    n20065, n20066, n20067, n20068, n20069, n20070,
    n20071, n20072, n20073, n20074, n20075, n20076,
    n20077, n20078, n20079, n20080, n20081, n20082,
    n20083, n20084, n20085, n20086, n20087, n20088,
    n20089, n20090, n20091, n20092, n20093, n20094,
    n20095, n20096, n20097, n20098, n20099, n20100,
    n20101, n20102, n20103, n20104, n20105, n20106,
    n20107, n20108, n20109, n20110, n20111, n20112,
    n20113, n20114, n20115, n20116, n20117, n20118,
    n20119, n20120, n20121, n20122, n20123, n20124,
    n20125, n20126, n20127, n20128, n20129, n20130,
    n20131, n20132, n20133, n20134, n20135, n20136,
    n20137, n20138, n20139, n20140, n20141, n20142,
    n20143, n20144, n20145, n20146, n20147, n20148,
    n20149, n20150, n20151, n20152, n20153, n20154,
    n20155, n20156, n20157, n20158, n20159, n20160,
    n20161, n20162, n20163, n20164, n20165, n20166,
    n20167, n20168, n20169, n20170, n20171, n20172,
    n20173, n20174, n20175, n20176, n20177, n20178,
    n20179, n20180, n20181, n20182, n20183, n20184,
    n20185, n20186, n20187, n20188, n20189, n20190,
    n20191, n20192, n20193, n20194, n20195, n20196,
    n20197, n20198, n20199, n20200, n20201, n20202,
    n20203, n20204, n20205, n20206, n20207, n20208,
    n20209, n20210, n20211, n20212, n20213, n20214,
    n20215, n20216, n20217, n20218, n20219, n20220,
    n20221, n20222, n20223, n20224, n20225, n20226,
    n20227, n20228, n20229, n20230, n20231, n20232,
    n20233, n20234, n20235, n20236, n20237, n20238,
    n20239, n20240, n20241, n20242, n20243, n20244,
    n20245, n20246, n20247, n20248, n20249, n20250,
    n20251, n20252, n20253, n20254, n20255, n20256,
    n20257, n20258, n20259, n20260, n20261, n20262,
    n20263, n20264, n20265, n20266, n20267, n20268,
    n20269, n20270, n20271, n20272, n20273, n20274,
    n20275, n20276, n20277, n20278, n20279, n20280,
    n20281, n20282, n20283, n20284, n20285, n20286,
    n20287, n20288, n20289, n20290, n20291, n20292,
    n20293, n20294, n20295, n20296, n20297, n20299,
    n20300, n20301, n20302, n20303, n20304, n20305,
    n20306, n20307, n20308, n20309, n20310, n20311,
    n20312, n20313, n20314, n20315, n20316, n20317,
    n20318, n20319, n20320, n20321, n20322, n20323,
    n20324, n20325, n20326, n20327, n20328, n20329,
    n20330, n20331, n20332, n20333, n20334, n20335,
    n20336, n20337, n20338, n20339, n20340, n20341,
    n20342, n20343, n20344, n20345, n20346, n20347,
    n20348, n20349, n20350, n20351, n20352, n20353,
    n20354, n20355, n20356, n20357, n20358, n20359,
    n20360, n20361, n20362, n20363, n20364, n20365,
    n20366, n20367, n20368, n20369, n20370, n20371,
    n20372, n20373, n20374, n20375, n20376, n20377,
    n20378, n20379, n20380, n20381, n20382, n20383,
    n20384, n20385, n20386, n20387, n20388, n20389,
    n20390, n20391, n20392, n20393, n20394, n20395,
    n20396, n20397, n20398, n20399, n20400, n20401,
    n20402, n20403, n20404, n20405, n20406, n20407,
    n20408, n20409, n20410, n20411, n20412, n20413,
    n20414, n20415, n20416, n20417, n20418, n20419,
    n20420, n20421, n20422, n20423, n20424, n20425,
    n20426, n20427, n20428, n20429, n20430, n20431,
    n20432, n20433, n20434, n20435, n20436, n20437,
    n20438, n20439, n20440, n20441, n20442, n20443,
    n20444, n20445, n20446, n20447, n20448, n20449,
    n20450, n20451, n20452, n20453, n20454, n20455,
    n20456, n20457, n20458, n20459, n20460, n20461,
    n20462, n20463, n20464, n20465, n20466, n20467,
    n20468, n20469, n20470, n20471, n20472, n20473,
    n20474, n20475, n20476, n20477, n20478, n20479,
    n20480, n20481, n20482, n20483, n20484, n20485,
    n20486, n20487, n20488, n20489, n20490, n20491,
    n20492, n20493, n20494, n20495, n20496, n20497,
    n20498, n20499, n20500, n20501, n20502, n20503,
    n20504, n20505, n20506, n20507, n20508, n20509,
    n20510, n20511, n20512, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521,
    n20522, n20523, n20524, n20525, n20526, n20527,
    n20528, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539,
    n20540, n20541, n20542, n20543, n20544, n20545,
    n20546, n20547, n20548, n20549, n20550, n20551,
    n20552, n20553, n20554, n20555, n20556, n20557,
    n20558, n20559, n20560, n20561, n20562, n20563,
    n20564, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581,
    n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599,
    n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617,
    n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20631, n20632, n20633, n20634, n20635,
    n20636, n20637, n20638, n20639, n20640, n20641,
    n20642, n20643, n20644, n20645, n20646, n20647,
    n20648, n20649, n20650, n20651, n20652, n20653,
    n20654, n20655, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665,
    n20666, n20667, n20668, n20669, n20670, n20671,
    n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683,
    n20684, n20685, n20686, n20687, n20688, n20689,
    n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701,
    n20702, n20703, n20704, n20705, n20706, n20707,
    n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719,
    n20720, n20721, n20722, n20723, n20724, n20725,
    n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737,
    n20738, n20739, n20740, n20741, n20742, n20743,
    n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755,
    n20756, n20757, n20758, n20759, n20760, n20761,
    n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773,
    n20774, n20775, n20776, n20777, n20778, n20779,
    n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20789, n20790, n20791,
    n20792, n20793, n20794, n20795, n20796, n20797,
    n20798, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809,
    n20810, n20811, n20812, n20813, n20814, n20815,
    n20816, n20817, n20818, n20819, n20820, n20821,
    n20822, n20823, n20824, n20825, n20826, n20827,
    n20828, n20829, n20830, n20831, n20832, n20833,
    n20834, n20835, n20836, n20837, n20838, n20839,
    n20840, n20841, n20842, n20843, n20844, n20845,
    n20846, n20847, n20848, n20849, n20850, n20851,
    n20852, n20853, n20854, n20855, n20856, n20857,
    n20858, n20859, n20860, n20861, n20862, n20863,
    n20864, n20865, n20866, n20867, n20868, n20869,
    n20870, n20871, n20872, n20873, n20874, n20875,
    n20876, n20877, n20878, n20879, n20880, n20881,
    n20882, n20883, n20884, n20885, n20886, n20887,
    n20888, n20889, n20890, n20891, n20892, n20893,
    n20894, n20895, n20896, n20897, n20898, n20899,
    n20900, n20901, n20902, n20903, n20904, n20905,
    n20906, n20907, n20908, n20909, n20910, n20911,
    n20912, n20913, n20914, n20915, n20916, n20917,
    n20918, n20919, n20920, n20921, n20922, n20923,
    n20924, n20925, n20926, n20927, n20928, n20929,
    n20930, n20931, n20932, n20933, n20934, n20935,
    n20936, n20937, n20938, n20939, n20940, n20941,
    n20942, n20943, n20944, n20945, n20946, n20947,
    n20948, n20949, n20950, n20951, n20953, n20954,
    n20955, n20956, n20957, n20958, n20959, n20960,
    n20961, n20962, n20963, n20964, n20965, n20966,
    n20967, n20968, n20969, n20970, n20971, n20972,
    n20973, n20974, n20975, n20976, n20977, n20978,
    n20979, n20980, n20981, n20982, n20983, n20984,
    n20985, n20986, n20987, n20988, n20989, n20990,
    n20991, n20992, n20993, n20994, n20995, n20996,
    n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21005, n21006, n21007, n21008,
    n21009, n21010, n21011, n21012, n21013, n21014,
    n21015, n21016, n21017, n21018, n21019, n21020,
    n21021, n21022, n21023, n21024, n21025, n21026,
    n21027, n21028, n21029, n21030, n21031, n21032,
    n21033, n21034, n21035, n21036, n21037, n21038,
    n21039, n21040, n21041, n21042, n21043, n21044,
    n21045, n21046, n21047, n21048, n21049, n21050,
    n21051, n21052, n21053, n21054, n21055, n21056,
    n21057, n21058, n21059, n21060, n21061, n21062,
    n21063, n21064, n21065, n21066, n21067, n21068,
    n21069, n21070, n21071, n21072, n21073, n21074,
    n21075, n21076, n21077, n21078, n21079, n21080,
    n21081, n21082, n21083, n21084, n21085, n21086,
    n21087, n21088, n21089, n21090, n21091, n21092,
    n21093, n21094, n21095, n21096, n21097, n21098,
    n21099, n21100, n21101, n21102, n21103, n21104,
    n21105, n21106, n21107, n21108, n21109, n21110,
    n21111, n21112, n21113, n21114, n21115, n21116,
    n21117, n21118, n21119, n21120, n21121, n21122,
    n21123, n21124, n21125, n21126, n21127, n21128,
    n21129, n21130, n21131, n21132, n21133, n21134,
    n21135, n21136, n21137, n21138, n21139, n21140,
    n21141, n21142, n21143, n21144, n21145, n21146,
    n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158,
    n21159, n21160, n21161, n21162, n21163, n21164,
    n21165, n21166, n21167, n21168, n21169, n21170,
    n21171, n21172, n21173, n21174, n21175, n21176,
    n21177, n21178, n21179, n21180, n21181, n21182,
    n21183, n21184, n21185, n21186, n21187, n21188,
    n21189, n21190, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200,
    n21201, n21202, n21203, n21204, n21205, n21206,
    n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218,
    n21219, n21220, n21221, n21222, n21223, n21224,
    n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236,
    n21237, n21238, n21239, n21240, n21241, n21242,
    n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254,
    n21255, n21256, n21257, n21258, n21259, n21260,
    n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21268, n21269, n21270, n21271, n21272,
    n21273, n21274, n21275, n21276, n21277, n21278,
    n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290,
    n21291, n21292, n21293, n21294, n21295, n21296,
    n21297, n21298, n21299, n21300, n21301, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308,
    n21309, n21310, n21311, n21312, n21313, n21314,
    n21315, n21316, n21317, n21318, n21319, n21320,
    n21321, n21322, n21323, n21324, n21325, n21326,
    n21327, n21328, n21329, n21330, n21331, n21332,
    n21333, n21334, n21335, n21336, n21337, n21338,
    n21339, n21340, n21341, n21342, n21343, n21344,
    n21345, n21346, n21347, n21348, n21349, n21350,
    n21351, n21352, n21353, n21354, n21355, n21356,
    n21357, n21358, n21359, n21360, n21361, n21362,
    n21363, n21364, n21365, n21366, n21367, n21368,
    n21369, n21370, n21371, n21372, n21373, n21374,
    n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386,
    n21387, n21388, n21389, n21390, n21391, n21392,
    n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410,
    n21411, n21412, n21413, n21414, n21415, n21416,
    n21417, n21418, n21419, n21420, n21421, n21422,
    n21423, n21424, n21425, n21426, n21427, n21428,
    n21429, n21430, n21431, n21432, n21433, n21434,
    n21435, n21436, n21437, n21438, n21439, n21440,
    n21441, n21442, n21443, n21444, n21445, n21446,
    n21447, n21448, n21449, n21450, n21451, n21452,
    n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21463, n21464,
    n21465, n21466, n21467, n21468, n21469, n21470,
    n21471, n21472, n21473, n21474, n21475, n21476,
    n21477, n21478, n21479, n21480, n21481, n21482,
    n21483, n21484, n21485, n21486, n21487, n21488,
    n21489, n21490, n21491, n21492, n21493, n21494,
    n21495, n21496, n21497, n21498, n21499, n21500,
    n21501, n21502, n21503, n21504, n21505, n21506,
    n21507, n21508, n21509, n21510, n21511, n21512,
    n21513, n21514, n21515, n21516, n21517, n21518,
    n21519, n21520, n21521, n21522, n21523, n21524,
    n21525, n21526, n21527, n21528, n21529, n21530,
    n21531, n21532, n21533, n21534, n21535, n21536,
    n21537, n21538, n21539, n21540, n21541, n21542,
    n21543, n21544, n21545, n21546, n21547, n21548,
    n21549, n21550, n21551, n21552, n21553, n21554,
    n21555, n21556, n21557, n21558, n21559, n21560,
    n21561, n21562, n21563, n21564, n21565, n21566,
    n21567, n21568, n21569, n21570, n21571, n21572,
    n21573, n21574, n21575, n21576, n21577, n21578,
    n21579, n21580, n21581, n21582, n21583, n21584,
    n21585, n21586, n21587, n21588, n21589, n21590,
    n21591, n21592, n21593, n21594, n21595, n21596,
    n21597, n21598, n21599, n21600, n21601, n21602,
    n21603, n21604, n21605, n21606, n21607, n21608,
    n21609, n21610, n21611, n21612, n21613, n21614,
    n21615;
  assign po63  = pi126  | pi127 ;
  assign n194 = pi126  & pi127 ;
  assign n195 = ~pi124  & ~pi125 ;
  assign n196 = ~pi126  & ~n195;
  assign po62  = n194 | n196;
  assign n198 = pi124  & po62 ;
  assign n199 = ~pi122  & ~pi123 ;
  assign n200 = ~pi124  & n199;
  assign n201 = ~n198 & ~n200;
  assign n202 = ~pi124  & po62 ;
  assign n203 = pi125  & ~n202;
  assign n204 = n195 & po62 ;
  assign n205 = ~n203 & ~n204;
  assign n206 = ~n201 & n205;
  assign n207 = ~po63  & ~n206;
  assign n208 = n201 & ~n205;
  assign n209 = pi126  & n195;
  assign n210 = pi127  & ~n196;
  assign n211 = ~n209 & n210;
  assign n212 = ~n208 & ~n211;
  assign po61  = n207 | ~n212;
  assign n214 = pi122  & po61 ;
  assign n215 = ~pi120  & ~pi121 ;
  assign n216 = ~pi122  & n215;
  assign n217 = ~po62  & ~n216;
  assign n218 = ~n214 & n217;
  assign n219 = n199 & po61 ;
  assign n220 = ~pi122  & po61 ;
  assign n221 = pi123  & ~n220;
  assign n222 = ~n219 & ~n221;
  assign n223 = ~n214 & ~n216;
  assign n224 = po62  & ~n223;
  assign n225 = ~n218 & ~n224;
  assign n226 = ~n222 & n225;
  assign n227 = ~n218 & ~n226;
  assign n228 = po62  & ~po61 ;
  assign n229 = ~n219 & ~n228;
  assign n230 = pi124  & ~n229;
  assign n231 = ~pi124  & n229;
  assign n232 = ~n230 & ~n231;
  assign n233 = n206 & po61 ;
  assign n234 = ~n208 & ~n233;
  assign n235 = ~n232 & n234;
  assign n236 = n227 & n235;
  assign n237 = ~po63  & ~n236;
  assign n238 = ~n227 & n232;
  assign n239 = n205 & po61 ;
  assign n240 = n201 & ~n239;
  assign n241 = po63  & ~n206;
  assign n242 = ~n240 & n241;
  assign n243 = ~n238 & ~n242;
  assign po60  = n237 | ~n243;
  assign n245 = pi120  & po60 ;
  assign n246 = ~pi118  & ~pi119 ;
  assign n247 = ~pi120  & n246;
  assign n248 = ~n245 & ~n247;
  assign n249 = po61  & ~n248;
  assign n250 = ~pi120  & po60 ;
  assign n251 = pi121  & ~n250;
  assign n252 = n215 & po60 ;
  assign n253 = ~n251 & ~n252;
  assign n254 = ~po61  & ~n247;
  assign n255 = ~n245 & n254;
  assign n256 = n253 & ~n255;
  assign n257 = ~n249 & ~n256;
  assign n258 = po62  & ~n257;
  assign n259 = ~po62  & ~n249;
  assign n260 = ~n256 & n259;
  assign n261 = po61  & ~po60 ;
  assign n262 = ~n252 & ~n261;
  assign n263 = pi122  & ~n262;
  assign n264 = ~pi122  & n262;
  assign n265 = ~n263 & ~n264;
  assign n266 = ~n260 & ~n265;
  assign n267 = ~n258 & ~n266;
  assign n268 = n226 & po60 ;
  assign n269 = n225 & po60 ;
  assign n270 = n222 & ~n269;
  assign n271 = ~n268 & ~n270;
  assign n272 = ~n227 & po60 ;
  assign n273 = ~n232 & ~n272;
  assign n274 = po60  & n273;
  assign n275 = ~n238 & ~n271;
  assign n276 = ~n274 & n275;
  assign n277 = ~n267 & n276;
  assign n278 = ~po63  & ~n277;
  assign n279 = po63  & ~n238;
  assign n280 = ~n273 & n279;
  assign n281 = n267 & n271;
  assign n282 = ~n280 & ~n281;
  assign po59  = n278 | ~n282;
  assign n284 = pi118  & po59 ;
  assign n285 = ~pi116  & ~pi117 ;
  assign n286 = ~pi118  & n285;
  assign n287 = ~n284 & ~n286;
  assign n288 = po60  & ~n287;
  assign n289 = ~po60  & ~n286;
  assign n290 = ~n284 & n289;
  assign n291 = ~pi118  & po59 ;
  assign n292 = pi119  & ~n291;
  assign n293 = n246 & po59 ;
  assign n294 = ~n292 & ~n293;
  assign n295 = ~n290 & n294;
  assign n296 = ~n288 & ~n295;
  assign n297 = po61  & ~n296;
  assign n298 = po60  & ~po59 ;
  assign n299 = ~n293 & ~n298;
  assign n300 = pi120  & ~n299;
  assign n301 = ~pi120  & n299;
  assign n302 = ~n300 & ~n301;
  assign n303 = ~po61  & n296;
  assign n304 = ~n302 & ~n303;
  assign n305 = ~n297 & ~n304;
  assign n306 = po62  & ~n305;
  assign n307 = ~po62  & ~n297;
  assign n308 = ~n304 & n307;
  assign n309 = ~n249 & ~n255;
  assign n310 = ~n253 & n309;
  assign n311 = po59  & n310;
  assign n312 = po59  & n309;
  assign n313 = n253 & ~n312;
  assign n314 = ~n311 & ~n313;
  assign n315 = ~n308 & ~n314;
  assign n316 = ~n306 & ~n315;
  assign n317 = ~n258 & ~n260;
  assign n318 = po59  & n317;
  assign n319 = ~n265 & ~n318;
  assign n320 = n265 & n318;
  assign n321 = ~n319 & ~n320;
  assign n322 = n267 & po59 ;
  assign n323 = ~n271 & ~n322;
  assign n324 = po59  & n323;
  assign n325 = ~n281 & ~n321;
  assign n326 = ~n324 & n325;
  assign n327 = ~n316 & n326;
  assign n328 = ~po63  & ~n327;
  assign n329 = po63  & ~n281;
  assign n330 = ~n323 & n329;
  assign n331 = n316 & n321;
  assign n332 = ~n330 & ~n331;
  assign po58  = n328 | ~n332;
  assign n334 = pi116  & po58 ;
  assign n335 = ~pi114  & ~pi115 ;
  assign n336 = ~pi116  & n335;
  assign n337 = ~n334 & ~n336;
  assign n338 = po59  & ~n337;
  assign n339 = ~n205 & ~po61 ;
  assign n340 = ~n230 & ~n339;
  assign n341 = ~n231 & n340;
  assign n342 = ~po60  & n341;
  assign n343 = ~n336 & ~n342;
  assign n344 = ~po59  & n343;
  assign n345 = ~n334 & n344;
  assign n346 = ~pi116  & po58 ;
  assign n347 = pi117  & ~n346;
  assign n348 = n285 & po58 ;
  assign n349 = ~n347 & ~n348;
  assign n350 = ~n345 & n349;
  assign n351 = ~n338 & ~n350;
  assign n352 = po60  & ~n351;
  assign n353 = ~po60  & ~n338;
  assign n354 = ~n350 & n353;
  assign n355 = po59  & ~n330;
  assign n356 = ~n331 & n355;
  assign n357 = ~n328 & n356;
  assign n358 = ~n348 & ~n357;
  assign n359 = pi118  & ~n358;
  assign n360 = ~pi118  & n358;
  assign n361 = ~n359 & ~n360;
  assign n362 = ~n354 & ~n361;
  assign n363 = ~n352 & ~n362;
  assign n364 = po61  & ~n363;
  assign n365 = ~n288 & ~n290;
  assign n366 = ~n294 & n365;
  assign n367 = po58  & n366;
  assign n368 = po58  & n365;
  assign n369 = n294 & ~n368;
  assign n370 = ~n367 & ~n369;
  assign n371 = ~po61  & n363;
  assign n372 = ~n370 & ~n371;
  assign n373 = ~n364 & ~n372;
  assign n374 = po62  & ~n373;
  assign n375 = ~n297 & ~n303;
  assign n376 = ~n304 & n375;
  assign n377 = po58  & n376;
  assign n378 = po58  & n375;
  assign n379 = ~n302 & ~n378;
  assign n380 = ~n377 & ~n379;
  assign n381 = ~po62  & ~n364;
  assign n382 = ~n372 & n381;
  assign n383 = ~n380 & ~n382;
  assign n384 = ~n374 & ~n383;
  assign n385 = ~n306 & ~n308;
  assign n386 = po58  & n385;
  assign n387 = ~n314 & ~n386;
  assign n388 = n314 & n386;
  assign n389 = ~n387 & ~n388;
  assign n390 = ~n316 & ~n321;
  assign n391 = po58  & n390;
  assign n392 = ~n331 & ~n391;
  assign n393 = ~n389 & n392;
  assign n394 = ~n384 & n393;
  assign n395 = ~po63  & ~n394;
  assign n396 = ~n321 & po58 ;
  assign n397 = n316 & ~n396;
  assign n398 = po63  & ~n390;
  assign n399 = ~n397 & n398;
  assign n400 = n271 & ~n342;
  assign n401 = ~n280 & n400;
  assign n402 = ~n281 & n401;
  assign n403 = ~n278 & n402;
  assign n404 = ~n319 & ~n403;
  assign n405 = ~n320 & n404;
  assign n406 = ~po58  & n405;
  assign n407 = ~n399 & ~n406;
  assign n408 = n384 & n389;
  assign n409 = n407 & ~n408;
  assign po57  = n395 | ~n409;
  assign n411 = pi114  & po57 ;
  assign n412 = ~pi112  & ~pi113 ;
  assign n413 = ~pi114  & n412;
  assign n414 = ~n411 & ~n413;
  assign n415 = po58  & ~n414;
  assign n416 = ~n330 & ~n413;
  assign n417 = ~n331 & n416;
  assign n418 = ~n328 & n417;
  assign n419 = ~n411 & n418;
  assign n420 = ~pi114  & po57 ;
  assign n421 = pi115  & ~n420;
  assign n422 = n335 & po57 ;
  assign n423 = ~n421 & ~n422;
  assign n424 = ~n419 & n423;
  assign n425 = ~n415 & ~n424;
  assign n426 = po59  & ~n425;
  assign n427 = po58  & ~n399;
  assign n428 = ~n408 & n427;
  assign n429 = ~n395 & n428;
  assign n430 = ~n422 & ~n429;
  assign n431 = pi116  & ~n430;
  assign n432 = ~pi116  & n430;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~po59  & n425;
  assign n435 = ~n433 & ~n434;
  assign n436 = ~n426 & ~n435;
  assign n437 = po60  & ~n436;
  assign n438 = ~n338 & ~n345;
  assign n439 = ~n349 & n438;
  assign n440 = po57  & n439;
  assign n441 = po57  & n438;
  assign n442 = n349 & ~n441;
  assign n443 = ~n440 & ~n442;
  assign n444 = ~po60  & ~n426;
  assign n445 = ~n435 & n444;
  assign n446 = ~n443 & ~n445;
  assign n447 = ~n437 & ~n446;
  assign n448 = po61  & ~n447;
  assign n449 = ~n352 & ~n354;
  assign n450 = ~n362 & n449;
  assign n451 = po57  & n450;
  assign n452 = po57  & n449;
  assign n453 = ~n361 & ~n452;
  assign n454 = ~n451 & ~n453;
  assign n455 = ~po61  & n447;
  assign n456 = ~n454 & ~n455;
  assign n457 = ~n448 & ~n456;
  assign n458 = po62  & ~n457;
  assign n459 = ~n364 & ~n371;
  assign n460 = n370 & n459;
  assign n461 = po57  & n460;
  assign n462 = po57  & n459;
  assign n463 = ~n370 & ~n462;
  assign n464 = ~n461 & ~n463;
  assign n465 = ~po62  & ~n448;
  assign n466 = ~n456 & n465;
  assign n467 = ~n464 & ~n466;
  assign n468 = ~n458 & ~n467;
  assign n469 = ~n374 & ~n382;
  assign n470 = po57  & n469;
  assign n471 = ~n380 & ~n470;
  assign n472 = n380 & n470;
  assign n473 = ~n471 & ~n472;
  assign n474 = ~n384 & ~n389;
  assign n475 = po57  & n474;
  assign n476 = ~n408 & ~n475;
  assign n477 = ~n473 & n476;
  assign n478 = ~n468 & n477;
  assign n479 = ~po63  & ~n478;
  assign n480 = ~n389 & po57 ;
  assign n481 = n384 & ~n480;
  assign n482 = po63  & ~n474;
  assign n483 = ~n481 & n482;
  assign n484 = n389 & ~po57 ;
  assign n485 = ~n483 & ~n484;
  assign n486 = n468 & n473;
  assign n487 = n485 & ~n486;
  assign po56  = n479 | ~n487;
  assign n489 = pi112  & po56 ;
  assign n490 = ~pi110  & ~pi111 ;
  assign n491 = ~pi112  & n490;
  assign n492 = ~n489 & ~n491;
  assign n493 = po57  & ~n492;
  assign n494 = ~pi112  & po56 ;
  assign n495 = pi113  & ~n494;
  assign n496 = n412 & po56 ;
  assign n497 = ~n495 & ~n496;
  assign n498 = n407 & ~n491;
  assign n499 = ~n408 & n498;
  assign n500 = ~n395 & n499;
  assign n501 = ~n489 & n500;
  assign n502 = n497 & ~n501;
  assign n503 = ~n493 & ~n502;
  assign n504 = po58  & ~n503;
  assign n505 = ~po58  & ~n493;
  assign n506 = ~n502 & n505;
  assign n507 = po57  & n485;
  assign n508 = ~n486 & n507;
  assign n509 = ~n479 & n508;
  assign n510 = ~n496 & ~n509;
  assign n511 = pi114  & ~n510;
  assign n512 = ~pi114  & n510;
  assign n513 = ~n511 & ~n512;
  assign n514 = ~n506 & ~n513;
  assign n515 = ~n504 & ~n514;
  assign n516 = po59  & ~n515;
  assign n517 = ~n415 & ~n419;
  assign n518 = ~n423 & n517;
  assign n519 = po56  & n518;
  assign n520 = po56  & n517;
  assign n521 = n423 & ~n520;
  assign n522 = ~n519 & ~n521;
  assign n523 = ~po59  & n515;
  assign n524 = ~n522 & ~n523;
  assign n525 = ~n516 & ~n524;
  assign n526 = po60  & ~n525;
  assign n527 = ~n426 & ~n434;
  assign n528 = n433 & n527;
  assign n529 = po56  & n528;
  assign n530 = po56  & n527;
  assign n531 = ~n433 & ~n530;
  assign n532 = ~n529 & ~n531;
  assign n533 = ~po60  & ~n516;
  assign n534 = ~n524 & n533;
  assign n535 = ~n532 & ~n534;
  assign n536 = ~n526 & ~n535;
  assign n537 = po61  & ~n536;
  assign n538 = ~n437 & ~n445;
  assign n539 = n443 & n538;
  assign n540 = po56  & n539;
  assign n541 = po56  & n538;
  assign n542 = ~n443 & ~n541;
  assign n543 = ~n540 & ~n542;
  assign n544 = ~po61  & n536;
  assign n545 = ~n543 & ~n544;
  assign n546 = ~n537 & ~n545;
  assign n547 = po62  & ~n546;
  assign n548 = ~n448 & ~n455;
  assign n549 = n454 & n548;
  assign n550 = po56  & n549;
  assign n551 = po56  & n548;
  assign n552 = ~n454 & ~n551;
  assign n553 = ~n550 & ~n552;
  assign n554 = ~po62  & ~n537;
  assign n555 = ~n545 & n554;
  assign n556 = ~n553 & ~n555;
  assign n557 = ~n547 & ~n556;
  assign n558 = ~n458 & ~n466;
  assign n559 = po56  & n558;
  assign n560 = ~n464 & ~n559;
  assign n561 = n464 & n559;
  assign n562 = ~n560 & ~n561;
  assign n563 = ~n468 & ~n473;
  assign n564 = po56  & n563;
  assign n565 = ~n486 & ~n564;
  assign n566 = ~n562 & n565;
  assign n567 = ~n557 & n566;
  assign n568 = ~po63  & ~n567;
  assign n569 = ~n473 & po56 ;
  assign n570 = n468 & ~n569;
  assign n571 = po63  & ~n563;
  assign n572 = ~n570 & n571;
  assign n573 = n473 & ~po56 ;
  assign n574 = ~n572 & ~n573;
  assign n575 = n557 & n562;
  assign n576 = n574 & ~n575;
  assign po55  = n568 | ~n576;
  assign n578 = pi110  & po55 ;
  assign n579 = ~pi108  & ~pi109 ;
  assign n580 = ~pi110  & n579;
  assign n581 = ~n578 & ~n580;
  assign n582 = po56  & ~n581;
  assign n583 = n485 & ~n580;
  assign n584 = ~n486 & n583;
  assign n585 = ~n479 & n584;
  assign n586 = ~n578 & n585;
  assign n587 = ~pi110  & po55 ;
  assign n588 = pi111  & ~n587;
  assign n589 = n490 & po55 ;
  assign n590 = ~n588 & ~n589;
  assign n591 = ~n586 & n590;
  assign n592 = ~n582 & ~n591;
  assign n593 = po57  & ~n592;
  assign n594 = po56  & n574;
  assign n595 = ~n575 & n594;
  assign n596 = ~n568 & n595;
  assign n597 = ~n589 & ~n596;
  assign n598 = pi112  & ~n597;
  assign n599 = ~pi112  & n597;
  assign n600 = ~n598 & ~n599;
  assign n601 = ~po57  & n592;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~n593 & ~n602;
  assign n604 = po58  & ~n603;
  assign n605 = ~po58  & ~n593;
  assign n606 = ~n602 & n605;
  assign n607 = ~n493 & ~n501;
  assign n608 = ~n497 & n607;
  assign n609 = po55  & n608;
  assign n610 = po55  & n607;
  assign n611 = n497 & ~n610;
  assign n612 = ~n609 & ~n611;
  assign n613 = ~n606 & ~n612;
  assign n614 = ~n604 & ~n613;
  assign n615 = po59  & ~n614;
  assign n616 = ~n504 & ~n506;
  assign n617 = n513 & n616;
  assign n618 = po55  & n617;
  assign n619 = po55  & n616;
  assign n620 = ~n513 & ~n619;
  assign n621 = ~n618 & ~n620;
  assign n622 = ~po59  & n614;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~n615 & ~n623;
  assign n625 = po60  & ~n624;
  assign n626 = ~n516 & ~n523;
  assign n627 = n522 & n626;
  assign n628 = po55  & n627;
  assign n629 = po55  & n626;
  assign n630 = ~n522 & ~n629;
  assign n631 = ~n628 & ~n630;
  assign n632 = ~po60  & ~n615;
  assign n633 = ~n623 & n632;
  assign n634 = ~n631 & ~n633;
  assign n635 = ~n625 & ~n634;
  assign n636 = po61  & ~n635;
  assign n637 = ~n526 & ~n534;
  assign n638 = n532 & n637;
  assign n639 = po55  & n638;
  assign n640 = po55  & n637;
  assign n641 = ~n532 & ~n640;
  assign n642 = ~n639 & ~n641;
  assign n643 = ~po61  & n635;
  assign n644 = ~n642 & ~n643;
  assign n645 = ~n636 & ~n644;
  assign n646 = po62  & ~n645;
  assign n647 = ~n537 & ~n544;
  assign n648 = n543 & n647;
  assign n649 = po55  & n648;
  assign n650 = po55  & n647;
  assign n651 = ~n543 & ~n650;
  assign n652 = ~n649 & ~n651;
  assign n653 = ~po62  & ~n636;
  assign n654 = ~n644 & n653;
  assign n655 = ~n652 & ~n654;
  assign n656 = ~n646 & ~n655;
  assign n657 = ~n547 & ~n555;
  assign n658 = po55  & n657;
  assign n659 = ~n553 & ~n658;
  assign n660 = n553 & n658;
  assign n661 = ~n659 & ~n660;
  assign n662 = ~n557 & ~n562;
  assign n663 = po55  & n662;
  assign n664 = ~n575 & ~n663;
  assign n665 = ~n661 & n664;
  assign n666 = ~n656 & n665;
  assign n667 = ~po63  & ~n666;
  assign n668 = ~n562 & po55 ;
  assign n669 = n557 & ~n668;
  assign n670 = po63  & ~n662;
  assign n671 = ~n669 & n670;
  assign n672 = n562 & ~po55 ;
  assign n673 = ~n671 & ~n672;
  assign n674 = n656 & n661;
  assign n675 = n673 & ~n674;
  assign po54  = n667 | ~n675;
  assign n677 = pi108  & po54 ;
  assign n678 = ~pi106  & ~pi107 ;
  assign n679 = ~pi108  & n678;
  assign n680 = ~n677 & ~n679;
  assign n681 = po55  & ~n680;
  assign n682 = n574 & ~n679;
  assign n683 = ~n575 & n682;
  assign n684 = ~n568 & n683;
  assign n685 = ~n677 & n684;
  assign n686 = ~pi108  & po54 ;
  assign n687 = pi109  & ~n686;
  assign n688 = n579 & po54 ;
  assign n689 = ~n687 & ~n688;
  assign n690 = ~n685 & n689;
  assign n691 = ~n681 & ~n690;
  assign n692 = po56  & ~n691;
  assign n693 = ~po56  & ~n681;
  assign n694 = ~n690 & n693;
  assign n695 = po55  & n673;
  assign n696 = ~n674 & n695;
  assign n697 = ~n667 & n696;
  assign n698 = ~n688 & ~n697;
  assign n699 = pi110  & ~n698;
  assign n700 = ~pi110  & n698;
  assign n701 = ~n699 & ~n700;
  assign n702 = ~n694 & ~n701;
  assign n703 = ~n692 & ~n702;
  assign n704 = po57  & ~n703;
  assign n705 = ~n582 & ~n586;
  assign n706 = ~n590 & n705;
  assign n707 = po54  & n706;
  assign n708 = po54  & n705;
  assign n709 = n590 & ~n708;
  assign n710 = ~n707 & ~n709;
  assign n711 = ~po57  & n703;
  assign n712 = ~n710 & ~n711;
  assign n713 = ~n704 & ~n712;
  assign n714 = po58  & ~n713;
  assign n715 = ~n593 & ~n601;
  assign n716 = n600 & n715;
  assign n717 = po54  & n716;
  assign n718 = po54  & n715;
  assign n719 = ~n600 & ~n718;
  assign n720 = ~n717 & ~n719;
  assign n721 = ~po58  & ~n704;
  assign n722 = ~n712 & n721;
  assign n723 = ~n720 & ~n722;
  assign n724 = ~n714 & ~n723;
  assign n725 = po59  & ~n724;
  assign n726 = ~n604 & ~n606;
  assign n727 = n612 & n726;
  assign n728 = po54  & n727;
  assign n729 = po54  & n726;
  assign n730 = ~n612 & ~n729;
  assign n731 = ~n728 & ~n730;
  assign n732 = ~po59  & n724;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~n725 & ~n733;
  assign n735 = po60  & ~n734;
  assign n736 = ~n615 & ~n622;
  assign n737 = n621 & n736;
  assign n738 = po54  & n737;
  assign n739 = po54  & n736;
  assign n740 = ~n621 & ~n739;
  assign n741 = ~n738 & ~n740;
  assign n742 = ~po60  & ~n725;
  assign n743 = ~n733 & n742;
  assign n744 = ~n741 & ~n743;
  assign n745 = ~n735 & ~n744;
  assign n746 = po61  & ~n745;
  assign n747 = ~n625 & ~n633;
  assign n748 = n631 & n747;
  assign n749 = po54  & n748;
  assign n750 = po54  & n747;
  assign n751 = ~n631 & ~n750;
  assign n752 = ~n749 & ~n751;
  assign n753 = ~po61  & n745;
  assign n754 = ~n752 & ~n753;
  assign n755 = ~n746 & ~n754;
  assign n756 = po62  & ~n755;
  assign n757 = ~n636 & ~n643;
  assign n758 = n642 & n757;
  assign n759 = po54  & n758;
  assign n760 = po54  & n757;
  assign n761 = ~n642 & ~n760;
  assign n762 = ~n759 & ~n761;
  assign n763 = ~po62  & ~n746;
  assign n764 = ~n754 & n763;
  assign n765 = ~n762 & ~n764;
  assign n766 = ~n756 & ~n765;
  assign n767 = ~n646 & ~n654;
  assign n768 = po54  & n767;
  assign n769 = ~n652 & ~n768;
  assign n770 = n652 & n768;
  assign n771 = ~n769 & ~n770;
  assign n772 = ~n656 & ~n661;
  assign n773 = po54  & n772;
  assign n774 = ~n674 & ~n773;
  assign n775 = ~n771 & n774;
  assign n776 = ~n766 & n775;
  assign n777 = ~po63  & ~n776;
  assign n778 = ~n661 & po54 ;
  assign n779 = n656 & ~n778;
  assign n780 = po63  & ~n772;
  assign n781 = ~n779 & n780;
  assign n782 = n661 & ~po54 ;
  assign n783 = ~n781 & ~n782;
  assign n784 = n766 & n771;
  assign n785 = n783 & ~n784;
  assign po53  = n777 | ~n785;
  assign n787 = pi106  & po53 ;
  assign n788 = ~pi104  & ~pi105 ;
  assign n789 = ~pi106  & n788;
  assign n790 = ~n787 & ~n789;
  assign n791 = po54  & ~n790;
  assign n792 = n673 & ~n789;
  assign n793 = ~n674 & n792;
  assign n794 = ~n667 & n793;
  assign n795 = ~n787 & n794;
  assign n796 = ~pi106  & po53 ;
  assign n797 = pi107  & ~n796;
  assign n798 = n678 & po53 ;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~n795 & n799;
  assign n801 = ~n791 & ~n800;
  assign n802 = po55  & ~n801;
  assign n803 = po54  & n783;
  assign n804 = ~n784 & n803;
  assign n805 = ~n777 & n804;
  assign n806 = ~n798 & ~n805;
  assign n807 = pi108  & ~n806;
  assign n808 = ~pi108  & n806;
  assign n809 = ~n807 & ~n808;
  assign n810 = ~po55  & n801;
  assign n811 = ~n809 & ~n810;
  assign n812 = ~n802 & ~n811;
  assign n813 = po56  & ~n812;
  assign n814 = ~n681 & ~n685;
  assign n815 = ~n689 & n814;
  assign n816 = po53  & n815;
  assign n817 = po53  & n814;
  assign n818 = n689 & ~n817;
  assign n819 = ~n816 & ~n818;
  assign n820 = ~po56  & ~n802;
  assign n821 = ~n811 & n820;
  assign n822 = ~n819 & ~n821;
  assign n823 = ~n813 & ~n822;
  assign n824 = po57  & ~n823;
  assign n825 = ~n692 & ~n694;
  assign n826 = n701 & n825;
  assign n827 = po53  & n826;
  assign n828 = po53  & n825;
  assign n829 = ~n701 & ~n828;
  assign n830 = ~n827 & ~n829;
  assign n831 = ~po57  & n823;
  assign n832 = ~n830 & ~n831;
  assign n833 = ~n824 & ~n832;
  assign n834 = po58  & ~n833;
  assign n835 = ~n704 & ~n711;
  assign n836 = n710 & n835;
  assign n837 = po53  & n836;
  assign n838 = po53  & n835;
  assign n839 = ~n710 & ~n838;
  assign n840 = ~n837 & ~n839;
  assign n841 = ~po58  & ~n824;
  assign n842 = ~n832 & n841;
  assign n843 = ~n840 & ~n842;
  assign n844 = ~n834 & ~n843;
  assign n845 = po59  & ~n844;
  assign n846 = ~n714 & ~n722;
  assign n847 = n720 & n846;
  assign n848 = po53  & n847;
  assign n849 = po53  & n846;
  assign n850 = ~n720 & ~n849;
  assign n851 = ~n848 & ~n850;
  assign n852 = ~po59  & n844;
  assign n853 = ~n851 & ~n852;
  assign n854 = ~n845 & ~n853;
  assign n855 = po60  & ~n854;
  assign n856 = ~po60  & ~n845;
  assign n857 = ~n853 & n856;
  assign n858 = ~n725 & ~n732;
  assign n859 = n731 & n858;
  assign n860 = po53  & n859;
  assign n861 = po53  & n858;
  assign n862 = ~n731 & ~n861;
  assign n863 = ~n860 & ~n862;
  assign n864 = ~n857 & ~n863;
  assign n865 = ~n855 & ~n864;
  assign n866 = po61  & ~n865;
  assign n867 = ~n735 & ~n743;
  assign n868 = n741 & n867;
  assign n869 = po53  & n868;
  assign n870 = po53  & n867;
  assign n871 = ~n741 & ~n870;
  assign n872 = ~n869 & ~n871;
  assign n873 = ~po61  & n865;
  assign n874 = ~n872 & ~n873;
  assign n875 = ~n866 & ~n874;
  assign n876 = po62  & ~n875;
  assign n877 = ~n746 & ~n753;
  assign n878 = n752 & n877;
  assign n879 = po53  & n878;
  assign n880 = po53  & n877;
  assign n881 = ~n752 & ~n880;
  assign n882 = ~n879 & ~n881;
  assign n883 = ~po62  & ~n866;
  assign n884 = ~n874 & n883;
  assign n885 = ~n882 & ~n884;
  assign n886 = ~n876 & ~n885;
  assign n887 = ~n756 & ~n764;
  assign n888 = po53  & n887;
  assign n889 = ~n762 & ~n888;
  assign n890 = n762 & n888;
  assign n891 = ~n889 & ~n890;
  assign n892 = ~n766 & ~n771;
  assign n893 = po53  & n892;
  assign n894 = ~n784 & ~n893;
  assign n895 = ~n891 & n894;
  assign n896 = ~n886 & n895;
  assign n897 = ~po63  & ~n896;
  assign n898 = ~n771 & po53 ;
  assign n899 = n766 & ~n898;
  assign n900 = po63  & ~n892;
  assign n901 = ~n899 & n900;
  assign n902 = n771 & ~po53 ;
  assign n903 = ~n901 & ~n902;
  assign n904 = n886 & n891;
  assign n905 = n903 & ~n904;
  assign po52  = n897 | ~n905;
  assign n907 = pi104  & po52 ;
  assign n908 = ~pi102  & ~pi103 ;
  assign n909 = ~pi104  & n908;
  assign n910 = ~n907 & ~n909;
  assign n911 = po53  & ~n910;
  assign n912 = n783 & ~n909;
  assign n913 = ~n784 & n912;
  assign n914 = ~n777 & n913;
  assign n915 = ~n907 & n914;
  assign n916 = ~pi104  & po52 ;
  assign n917 = pi105  & ~n916;
  assign n918 = n788 & po52 ;
  assign n919 = ~n917 & ~n918;
  assign n920 = ~n915 & n919;
  assign n921 = ~n911 & ~n920;
  assign n922 = po54  & ~n921;
  assign n923 = ~po54  & ~n911;
  assign n924 = ~n920 & n923;
  assign n925 = po53  & n903;
  assign n926 = ~n904 & n925;
  assign n927 = ~n897 & n926;
  assign n928 = ~n918 & ~n927;
  assign n929 = pi106  & ~n928;
  assign n930 = ~pi106  & n928;
  assign n931 = ~n929 & ~n930;
  assign n932 = ~n924 & ~n931;
  assign n933 = ~n922 & ~n932;
  assign n934 = po55  & ~n933;
  assign n935 = ~n791 & ~n795;
  assign n936 = ~n799 & n935;
  assign n937 = po52  & n936;
  assign n938 = po52  & n935;
  assign n939 = n799 & ~n938;
  assign n940 = ~n937 & ~n939;
  assign n941 = ~po55  & n933;
  assign n942 = ~n940 & ~n941;
  assign n943 = ~n934 & ~n942;
  assign n944 = po56  & ~n943;
  assign n945 = ~n802 & ~n810;
  assign n946 = n809 & n945;
  assign n947 = po52  & n946;
  assign n948 = po52  & n945;
  assign n949 = ~n809 & ~n948;
  assign n950 = ~n947 & ~n949;
  assign n951 = ~po56  & ~n934;
  assign n952 = ~n942 & n951;
  assign n953 = ~n950 & ~n952;
  assign n954 = ~n944 & ~n953;
  assign n955 = po57  & ~n954;
  assign n956 = ~n813 & ~n821;
  assign n957 = n819 & n956;
  assign n958 = po52  & n957;
  assign n959 = po52  & n956;
  assign n960 = ~n819 & ~n959;
  assign n961 = ~n958 & ~n960;
  assign n962 = ~po57  & n954;
  assign n963 = ~n961 & ~n962;
  assign n964 = ~n955 & ~n963;
  assign n965 = po58  & ~n964;
  assign n966 = ~n824 & ~n831;
  assign n967 = n830 & n966;
  assign n968 = po52  & n967;
  assign n969 = po52  & n966;
  assign n970 = ~n830 & ~n969;
  assign n971 = ~n968 & ~n970;
  assign n972 = ~po58  & ~n955;
  assign n973 = ~n963 & n972;
  assign n974 = ~n971 & ~n973;
  assign n975 = ~n965 & ~n974;
  assign n976 = po59  & ~n975;
  assign n977 = ~n834 & ~n842;
  assign n978 = n840 & n977;
  assign n979 = po52  & n978;
  assign n980 = po52  & n977;
  assign n981 = ~n840 & ~n980;
  assign n982 = ~n979 & ~n981;
  assign n983 = ~po59  & n975;
  assign n984 = ~n982 & ~n983;
  assign n985 = ~n976 & ~n984;
  assign n986 = po60  & ~n985;
  assign n987 = ~n845 & ~n852;
  assign n988 = n851 & n987;
  assign n989 = po52  & n988;
  assign n990 = po52  & n987;
  assign n991 = ~n851 & ~n990;
  assign n992 = ~n989 & ~n991;
  assign n993 = ~po60  & ~n976;
  assign n994 = ~n984 & n993;
  assign n995 = ~n992 & ~n994;
  assign n996 = ~n986 & ~n995;
  assign n997 = po61  & ~n996;
  assign n998 = ~n855 & ~n857;
  assign n999 = n863 & n998;
  assign n1000 = po52  & n999;
  assign n1001 = po52  & n998;
  assign n1002 = ~n863 & ~n1001;
  assign n1003 = ~n1000 & ~n1002;
  assign n1004 = ~po61  & n996;
  assign n1005 = ~n1003 & ~n1004;
  assign n1006 = ~n997 & ~n1005;
  assign n1007 = po62  & ~n1006;
  assign n1008 = ~n866 & ~n873;
  assign n1009 = n872 & n1008;
  assign n1010 = po52  & n1009;
  assign n1011 = po52  & n1008;
  assign n1012 = ~n872 & ~n1011;
  assign n1013 = ~n1010 & ~n1012;
  assign n1014 = ~po62  & ~n997;
  assign n1015 = ~n1005 & n1014;
  assign n1016 = ~n1013 & ~n1015;
  assign n1017 = ~n1007 & ~n1016;
  assign n1018 = ~n876 & ~n884;
  assign n1019 = po52  & n1018;
  assign n1020 = ~n882 & ~n1019;
  assign n1021 = n882 & n1019;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n886 & ~n891;
  assign n1024 = po52  & n1023;
  assign n1025 = ~n904 & ~n1024;
  assign n1026 = ~n1022 & n1025;
  assign n1027 = ~n1017 & n1026;
  assign n1028 = ~po63  & ~n1027;
  assign n1029 = ~n891 & po52 ;
  assign n1030 = n886 & ~n1029;
  assign n1031 = po63  & ~n1023;
  assign n1032 = ~n1030 & n1031;
  assign n1033 = n891 & ~po52 ;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = n1017 & n1022;
  assign n1036 = n1034 & ~n1035;
  assign po51  = n1028 | ~n1036;
  assign n1038 = pi102  & po51 ;
  assign n1039 = ~pi100  & ~pi101 ;
  assign n1040 = ~pi102  & n1039;
  assign n1041 = ~n1038 & ~n1040;
  assign n1042 = po52  & ~n1041;
  assign n1043 = n903 & ~n1040;
  assign n1044 = ~n904 & n1043;
  assign n1045 = ~n897 & n1044;
  assign n1046 = ~n1038 & n1045;
  assign n1047 = ~pi102  & po51 ;
  assign n1048 = pi103  & ~n1047;
  assign n1049 = n908 & po51 ;
  assign n1050 = ~n1048 & ~n1049;
  assign n1051 = ~n1046 & n1050;
  assign n1052 = ~n1042 & ~n1051;
  assign n1053 = po53  & ~n1052;
  assign n1054 = po52  & n1034;
  assign n1055 = ~n1035 & n1054;
  assign n1056 = ~n1028 & n1055;
  assign n1057 = ~n1049 & ~n1056;
  assign n1058 = pi104  & ~n1057;
  assign n1059 = ~pi104  & n1057;
  assign n1060 = ~n1058 & ~n1059;
  assign n1061 = ~po53  & n1052;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~n1053 & ~n1062;
  assign n1064 = po54  & ~n1063;
  assign n1065 = ~n911 & ~n915;
  assign n1066 = ~n919 & n1065;
  assign n1067 = po51  & n1066;
  assign n1068 = po51  & n1065;
  assign n1069 = n919 & ~n1068;
  assign n1070 = ~n1067 & ~n1069;
  assign n1071 = ~po54  & ~n1053;
  assign n1072 = ~n1062 & n1071;
  assign n1073 = ~n1070 & ~n1072;
  assign n1074 = ~n1064 & ~n1073;
  assign n1075 = po55  & ~n1074;
  assign n1076 = ~n922 & ~n924;
  assign n1077 = n931 & n1076;
  assign n1078 = po51  & n1077;
  assign n1079 = po51  & n1076;
  assign n1080 = ~n931 & ~n1079;
  assign n1081 = ~n1078 & ~n1080;
  assign n1082 = ~po55  & n1074;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = ~n1075 & ~n1083;
  assign n1085 = po56  & ~n1084;
  assign n1086 = ~n934 & ~n941;
  assign n1087 = n940 & n1086;
  assign n1088 = po51  & n1087;
  assign n1089 = po51  & n1086;
  assign n1090 = ~n940 & ~n1089;
  assign n1091 = ~n1088 & ~n1090;
  assign n1092 = ~po56  & ~n1075;
  assign n1093 = ~n1083 & n1092;
  assign n1094 = ~n1091 & ~n1093;
  assign n1095 = ~n1085 & ~n1094;
  assign n1096 = po57  & ~n1095;
  assign n1097 = ~n944 & ~n952;
  assign n1098 = n950 & n1097;
  assign n1099 = po51  & n1098;
  assign n1100 = po51  & n1097;
  assign n1101 = ~n950 & ~n1100;
  assign n1102 = ~n1099 & ~n1101;
  assign n1103 = ~po57  & n1095;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~n1096 & ~n1104;
  assign n1106 = po58  & ~n1105;
  assign n1107 = ~n955 & ~n962;
  assign n1108 = n961 & n1107;
  assign n1109 = po51  & n1108;
  assign n1110 = po51  & n1107;
  assign n1111 = ~n961 & ~n1110;
  assign n1112 = ~n1109 & ~n1111;
  assign n1113 = ~po58  & ~n1096;
  assign n1114 = ~n1104 & n1113;
  assign n1115 = ~n1112 & ~n1114;
  assign n1116 = ~n1106 & ~n1115;
  assign n1117 = po59  & ~n1116;
  assign n1118 = ~n965 & ~n973;
  assign n1119 = n971 & n1118;
  assign n1120 = po51  & n1119;
  assign n1121 = po51  & n1118;
  assign n1122 = ~n971 & ~n1121;
  assign n1123 = ~n1120 & ~n1122;
  assign n1124 = ~po59  & n1116;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~n1117 & ~n1125;
  assign n1127 = po60  & ~n1126;
  assign n1128 = ~n976 & ~n983;
  assign n1129 = n982 & n1128;
  assign n1130 = po51  & n1129;
  assign n1131 = po51  & n1128;
  assign n1132 = ~n982 & ~n1131;
  assign n1133 = ~n1130 & ~n1132;
  assign n1134 = ~po60  & ~n1117;
  assign n1135 = ~n1125 & n1134;
  assign n1136 = ~n1133 & ~n1135;
  assign n1137 = ~n1127 & ~n1136;
  assign n1138 = po61  & ~n1137;
  assign n1139 = ~n986 & ~n994;
  assign n1140 = n992 & n1139;
  assign n1141 = po51  & n1140;
  assign n1142 = po51  & n1139;
  assign n1143 = ~n992 & ~n1142;
  assign n1144 = ~n1141 & ~n1143;
  assign n1145 = ~po61  & n1137;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = ~n1138 & ~n1146;
  assign n1148 = po62  & ~n1147;
  assign n1149 = ~po62  & ~n1138;
  assign n1150 = ~n1146 & n1149;
  assign n1151 = ~n997 & ~n1004;
  assign n1152 = n1003 & n1151;
  assign n1153 = po51  & n1152;
  assign n1154 = po51  & n1151;
  assign n1155 = ~n1003 & ~n1154;
  assign n1156 = ~n1153 & ~n1155;
  assign n1157 = ~n1150 & ~n1156;
  assign n1158 = ~n1148 & ~n1157;
  assign n1159 = ~n1007 & ~n1015;
  assign n1160 = po51  & n1159;
  assign n1161 = ~n1013 & ~n1160;
  assign n1162 = n1013 & n1160;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = ~n1017 & ~n1022;
  assign n1165 = po51  & n1164;
  assign n1166 = ~n1035 & ~n1165;
  assign n1167 = ~n1163 & n1166;
  assign n1168 = ~n1158 & n1167;
  assign n1169 = ~po63  & ~n1168;
  assign n1170 = ~n1022 & po51 ;
  assign n1171 = n1017 & ~n1170;
  assign n1172 = po63  & ~n1164;
  assign n1173 = ~n1171 & n1172;
  assign n1174 = n1022 & ~po51 ;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = n1158 & n1163;
  assign n1177 = n1175 & ~n1176;
  assign po50  = n1169 | ~n1177;
  assign n1179 = pi100  & po50 ;
  assign n1180 = ~pi98  & ~pi99 ;
  assign n1181 = ~pi100  & n1180;
  assign n1182 = ~n1179 & ~n1181;
  assign n1183 = po51  & ~n1182;
  assign n1184 = n1034 & ~n1181;
  assign n1185 = ~n1035 & n1184;
  assign n1186 = ~n1028 & n1185;
  assign n1187 = ~n1179 & n1186;
  assign n1188 = ~pi100  & po50 ;
  assign n1189 = pi101  & ~n1188;
  assign n1190 = n1039 & po50 ;
  assign n1191 = ~n1189 & ~n1190;
  assign n1192 = ~n1187 & n1191;
  assign n1193 = ~n1183 & ~n1192;
  assign n1194 = po52  & ~n1193;
  assign n1195 = ~po52  & ~n1183;
  assign n1196 = ~n1192 & n1195;
  assign n1197 = po51  & n1175;
  assign n1198 = ~n1176 & n1197;
  assign n1199 = ~n1169 & n1198;
  assign n1200 = ~n1190 & ~n1199;
  assign n1201 = pi102  & ~n1200;
  assign n1202 = ~pi102  & n1200;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = ~n1196 & ~n1203;
  assign n1205 = ~n1194 & ~n1204;
  assign n1206 = po53  & ~n1205;
  assign n1207 = ~n1042 & ~n1046;
  assign n1208 = ~n1050 & n1207;
  assign n1209 = po50  & n1208;
  assign n1210 = po50  & n1207;
  assign n1211 = n1050 & ~n1210;
  assign n1212 = ~n1209 & ~n1211;
  assign n1213 = ~po53  & n1205;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = ~n1206 & ~n1214;
  assign n1216 = po54  & ~n1215;
  assign n1217 = ~n1053 & ~n1061;
  assign n1218 = n1060 & n1217;
  assign n1219 = po50  & n1218;
  assign n1220 = po50  & n1217;
  assign n1221 = ~n1060 & ~n1220;
  assign n1222 = ~n1219 & ~n1221;
  assign n1223 = ~po54  & ~n1206;
  assign n1224 = ~n1214 & n1223;
  assign n1225 = ~n1222 & ~n1224;
  assign n1226 = ~n1216 & ~n1225;
  assign n1227 = po55  & ~n1226;
  assign n1228 = ~n1064 & ~n1072;
  assign n1229 = n1070 & n1228;
  assign n1230 = po50  & n1229;
  assign n1231 = po50  & n1228;
  assign n1232 = ~n1070 & ~n1231;
  assign n1233 = ~n1230 & ~n1232;
  assign n1234 = ~po55  & n1226;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = ~n1227 & ~n1235;
  assign n1237 = po56  & ~n1236;
  assign n1238 = ~n1075 & ~n1082;
  assign n1239 = n1081 & n1238;
  assign n1240 = po50  & n1239;
  assign n1241 = po50  & n1238;
  assign n1242 = ~n1081 & ~n1241;
  assign n1243 = ~n1240 & ~n1242;
  assign n1244 = ~po56  & ~n1227;
  assign n1245 = ~n1235 & n1244;
  assign n1246 = ~n1243 & ~n1245;
  assign n1247 = ~n1237 & ~n1246;
  assign n1248 = po57  & ~n1247;
  assign n1249 = ~n1085 & ~n1093;
  assign n1250 = n1091 & n1249;
  assign n1251 = po50  & n1250;
  assign n1252 = po50  & n1249;
  assign n1253 = ~n1091 & ~n1252;
  assign n1254 = ~n1251 & ~n1253;
  assign n1255 = ~po57  & n1247;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = ~n1248 & ~n1256;
  assign n1258 = po58  & ~n1257;
  assign n1259 = ~n1096 & ~n1103;
  assign n1260 = n1102 & n1259;
  assign n1261 = po50  & n1260;
  assign n1262 = po50  & n1259;
  assign n1263 = ~n1102 & ~n1262;
  assign n1264 = ~n1261 & ~n1263;
  assign n1265 = ~po58  & ~n1248;
  assign n1266 = ~n1256 & n1265;
  assign n1267 = ~n1264 & ~n1266;
  assign n1268 = ~n1258 & ~n1267;
  assign n1269 = po59  & ~n1268;
  assign n1270 = ~n1106 & ~n1114;
  assign n1271 = n1112 & n1270;
  assign n1272 = po50  & n1271;
  assign n1273 = po50  & n1270;
  assign n1274 = ~n1112 & ~n1273;
  assign n1275 = ~n1272 & ~n1274;
  assign n1276 = ~po59  & n1268;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = ~n1269 & ~n1277;
  assign n1279 = po60  & ~n1278;
  assign n1280 = ~n1117 & ~n1124;
  assign n1281 = n1123 & n1280;
  assign n1282 = po50  & n1281;
  assign n1283 = po50  & n1280;
  assign n1284 = ~n1123 & ~n1283;
  assign n1285 = ~n1282 & ~n1284;
  assign n1286 = ~po60  & ~n1269;
  assign n1287 = ~n1277 & n1286;
  assign n1288 = ~n1285 & ~n1287;
  assign n1289 = ~n1279 & ~n1288;
  assign n1290 = po61  & ~n1289;
  assign n1291 = ~n1127 & ~n1135;
  assign n1292 = n1133 & n1291;
  assign n1293 = po50  & n1292;
  assign n1294 = po50  & n1291;
  assign n1295 = ~n1133 & ~n1294;
  assign n1296 = ~n1293 & ~n1295;
  assign n1297 = ~po61  & n1289;
  assign n1298 = ~n1296 & ~n1297;
  assign n1299 = ~n1290 & ~n1298;
  assign n1300 = po62  & ~n1299;
  assign n1301 = ~n1138 & ~n1145;
  assign n1302 = n1144 & n1301;
  assign n1303 = po50  & n1302;
  assign n1304 = po50  & n1301;
  assign n1305 = ~n1144 & ~n1304;
  assign n1306 = ~n1303 & ~n1305;
  assign n1307 = ~po62  & ~n1290;
  assign n1308 = ~n1298 & n1307;
  assign n1309 = ~n1306 & ~n1308;
  assign n1310 = ~n1300 & ~n1309;
  assign n1311 = ~n1148 & ~n1150;
  assign n1312 = po50  & n1311;
  assign n1313 = ~n1156 & ~n1312;
  assign n1314 = n1156 & n1312;
  assign n1315 = ~n1313 & ~n1314;
  assign n1316 = ~n1158 & ~n1163;
  assign n1317 = po50  & n1316;
  assign n1318 = ~n1176 & ~n1317;
  assign n1319 = ~n1315 & n1318;
  assign n1320 = ~n1310 & n1319;
  assign n1321 = ~po63  & ~n1320;
  assign n1322 = ~n1163 & po50 ;
  assign n1323 = n1158 & ~n1322;
  assign n1324 = po63  & ~n1316;
  assign n1325 = ~n1323 & n1324;
  assign n1326 = n1163 & ~po50 ;
  assign n1327 = ~n1325 & ~n1326;
  assign n1328 = n1310 & n1315;
  assign n1329 = n1327 & ~n1328;
  assign po49  = n1321 | ~n1329;
  assign n1331 = pi98  & po49 ;
  assign n1332 = ~pi96  & ~pi97 ;
  assign n1333 = ~pi98  & n1332;
  assign n1334 = ~n1331 & ~n1333;
  assign n1335 = po50  & ~n1334;
  assign n1336 = n1175 & ~n1333;
  assign n1337 = ~n1176 & n1336;
  assign n1338 = ~n1169 & n1337;
  assign n1339 = ~n1331 & n1338;
  assign n1340 = ~pi98  & po49 ;
  assign n1341 = pi99  & ~n1340;
  assign n1342 = n1180 & po49 ;
  assign n1343 = ~n1341 & ~n1342;
  assign n1344 = ~n1339 & n1343;
  assign n1345 = ~n1335 & ~n1344;
  assign n1346 = po51  & ~n1345;
  assign n1347 = po50  & n1327;
  assign n1348 = ~n1328 & n1347;
  assign n1349 = ~n1321 & n1348;
  assign n1350 = ~n1342 & ~n1349;
  assign n1351 = pi100  & ~n1350;
  assign n1352 = ~pi100  & n1350;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = ~po51  & n1345;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = ~n1346 & ~n1355;
  assign n1357 = po52  & ~n1356;
  assign n1358 = ~n1183 & ~n1187;
  assign n1359 = ~n1191 & n1358;
  assign n1360 = po49  & n1359;
  assign n1361 = po49  & n1358;
  assign n1362 = n1191 & ~n1361;
  assign n1363 = ~n1360 & ~n1362;
  assign n1364 = ~po52  & ~n1346;
  assign n1365 = ~n1355 & n1364;
  assign n1366 = ~n1363 & ~n1365;
  assign n1367 = ~n1357 & ~n1366;
  assign n1368 = po53  & ~n1367;
  assign n1369 = ~n1194 & ~n1196;
  assign n1370 = n1203 & n1369;
  assign n1371 = po49  & n1370;
  assign n1372 = po49  & n1369;
  assign n1373 = ~n1203 & ~n1372;
  assign n1374 = ~n1371 & ~n1373;
  assign n1375 = ~po53  & n1367;
  assign n1376 = ~n1374 & ~n1375;
  assign n1377 = ~n1368 & ~n1376;
  assign n1378 = po54  & ~n1377;
  assign n1379 = ~n1206 & ~n1213;
  assign n1380 = n1212 & n1379;
  assign n1381 = po49  & n1380;
  assign n1382 = po49  & n1379;
  assign n1383 = ~n1212 & ~n1382;
  assign n1384 = ~n1381 & ~n1383;
  assign n1385 = ~po54  & ~n1368;
  assign n1386 = ~n1376 & n1385;
  assign n1387 = ~n1384 & ~n1386;
  assign n1388 = ~n1378 & ~n1387;
  assign n1389 = po55  & ~n1388;
  assign n1390 = ~n1216 & ~n1224;
  assign n1391 = n1222 & n1390;
  assign n1392 = po49  & n1391;
  assign n1393 = po49  & n1390;
  assign n1394 = ~n1222 & ~n1393;
  assign n1395 = ~n1392 & ~n1394;
  assign n1396 = ~po55  & n1388;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = ~n1389 & ~n1397;
  assign n1399 = po56  & ~n1398;
  assign n1400 = ~n1227 & ~n1234;
  assign n1401 = n1233 & n1400;
  assign n1402 = po49  & n1401;
  assign n1403 = po49  & n1400;
  assign n1404 = ~n1233 & ~n1403;
  assign n1405 = ~n1402 & ~n1404;
  assign n1406 = ~po56  & ~n1389;
  assign n1407 = ~n1397 & n1406;
  assign n1408 = ~n1405 & ~n1407;
  assign n1409 = ~n1399 & ~n1408;
  assign n1410 = po57  & ~n1409;
  assign n1411 = ~n1237 & ~n1245;
  assign n1412 = n1243 & n1411;
  assign n1413 = po49  & n1412;
  assign n1414 = po49  & n1411;
  assign n1415 = ~n1243 & ~n1414;
  assign n1416 = ~n1413 & ~n1415;
  assign n1417 = ~po57  & n1409;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = ~n1410 & ~n1418;
  assign n1420 = po58  & ~n1419;
  assign n1421 = ~n1248 & ~n1255;
  assign n1422 = n1254 & n1421;
  assign n1423 = po49  & n1422;
  assign n1424 = po49  & n1421;
  assign n1425 = ~n1254 & ~n1424;
  assign n1426 = ~n1423 & ~n1425;
  assign n1427 = ~po58  & ~n1410;
  assign n1428 = ~n1418 & n1427;
  assign n1429 = ~n1426 & ~n1428;
  assign n1430 = ~n1420 & ~n1429;
  assign n1431 = po59  & ~n1430;
  assign n1432 = ~n1258 & ~n1266;
  assign n1433 = n1264 & n1432;
  assign n1434 = po49  & n1433;
  assign n1435 = po49  & n1432;
  assign n1436 = ~n1264 & ~n1435;
  assign n1437 = ~n1434 & ~n1436;
  assign n1438 = ~po59  & n1430;
  assign n1439 = ~n1437 & ~n1438;
  assign n1440 = ~n1431 & ~n1439;
  assign n1441 = po60  & ~n1440;
  assign n1442 = ~n1269 & ~n1276;
  assign n1443 = n1275 & n1442;
  assign n1444 = po49  & n1443;
  assign n1445 = po49  & n1442;
  assign n1446 = ~n1275 & ~n1445;
  assign n1447 = ~n1444 & ~n1446;
  assign n1448 = ~po60  & ~n1431;
  assign n1449 = ~n1439 & n1448;
  assign n1450 = ~n1447 & ~n1449;
  assign n1451 = ~n1441 & ~n1450;
  assign n1452 = po61  & ~n1451;
  assign n1453 = ~n1279 & ~n1287;
  assign n1454 = n1285 & n1453;
  assign n1455 = po49  & n1454;
  assign n1456 = po49  & n1453;
  assign n1457 = ~n1285 & ~n1456;
  assign n1458 = ~n1455 & ~n1457;
  assign n1459 = ~po61  & n1451;
  assign n1460 = ~n1458 & ~n1459;
  assign n1461 = ~n1452 & ~n1460;
  assign n1462 = po62  & ~n1461;
  assign n1463 = ~n1290 & ~n1297;
  assign n1464 = n1296 & n1463;
  assign n1465 = po49  & n1464;
  assign n1466 = po49  & n1463;
  assign n1467 = ~n1296 & ~n1466;
  assign n1468 = ~n1465 & ~n1467;
  assign n1469 = ~po62  & ~n1452;
  assign n1470 = ~n1460 & n1469;
  assign n1471 = ~n1468 & ~n1470;
  assign n1472 = ~n1462 & ~n1471;
  assign n1473 = ~n1300 & ~n1308;
  assign n1474 = po49  & n1473;
  assign n1475 = ~n1306 & ~n1474;
  assign n1476 = n1306 & n1474;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = ~n1310 & ~n1315;
  assign n1479 = po49  & n1478;
  assign n1480 = ~n1328 & ~n1479;
  assign n1481 = ~n1477 & n1480;
  assign n1482 = ~n1472 & n1481;
  assign n1483 = ~po63  & ~n1482;
  assign n1484 = ~n1315 & po49 ;
  assign n1485 = n1310 & ~n1484;
  assign n1486 = po63  & ~n1478;
  assign n1487 = ~n1485 & n1486;
  assign n1488 = n1315 & ~po49 ;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = n1472 & n1477;
  assign n1491 = n1489 & ~n1490;
  assign po48  = n1483 | ~n1491;
  assign n1493 = pi96  & po48 ;
  assign n1494 = ~pi94  & ~pi95 ;
  assign n1495 = ~pi96  & n1494;
  assign n1496 = ~n1493 & ~n1495;
  assign n1497 = po49  & ~n1496;
  assign n1498 = ~pi96  & po48 ;
  assign n1499 = pi97  & ~n1498;
  assign n1500 = n1332 & po48 ;
  assign n1501 = ~n1499 & ~n1500;
  assign n1502 = n1327 & ~n1495;
  assign n1503 = ~n1328 & n1502;
  assign n1504 = ~n1321 & n1503;
  assign n1505 = ~n1493 & n1504;
  assign n1506 = n1501 & ~n1505;
  assign n1507 = ~n1497 & ~n1506;
  assign n1508 = po50  & ~n1507;
  assign n1509 = ~po50  & ~n1497;
  assign n1510 = ~n1506 & n1509;
  assign n1511 = po49  & n1489;
  assign n1512 = ~n1490 & n1511;
  assign n1513 = ~n1483 & n1512;
  assign n1514 = ~n1500 & ~n1513;
  assign n1515 = pi98  & ~n1514;
  assign n1516 = ~pi98  & n1514;
  assign n1517 = ~n1515 & ~n1516;
  assign n1518 = ~n1510 & ~n1517;
  assign n1519 = ~n1508 & ~n1518;
  assign n1520 = po51  & ~n1519;
  assign n1521 = ~n1335 & ~n1339;
  assign n1522 = ~n1343 & n1521;
  assign n1523 = po48  & n1522;
  assign n1524 = po48  & n1521;
  assign n1525 = n1343 & ~n1524;
  assign n1526 = ~n1523 & ~n1525;
  assign n1527 = ~po51  & n1519;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = ~n1520 & ~n1528;
  assign n1530 = po52  & ~n1529;
  assign n1531 = ~n1346 & ~n1354;
  assign n1532 = n1353 & n1531;
  assign n1533 = po48  & n1532;
  assign n1534 = po48  & n1531;
  assign n1535 = ~n1353 & ~n1534;
  assign n1536 = ~n1533 & ~n1535;
  assign n1537 = ~po52  & ~n1520;
  assign n1538 = ~n1528 & n1537;
  assign n1539 = ~n1536 & ~n1538;
  assign n1540 = ~n1530 & ~n1539;
  assign n1541 = po53  & ~n1540;
  assign n1542 = ~n1357 & ~n1365;
  assign n1543 = n1363 & n1542;
  assign n1544 = po48  & n1543;
  assign n1545 = po48  & n1542;
  assign n1546 = ~n1363 & ~n1545;
  assign n1547 = ~n1544 & ~n1546;
  assign n1548 = ~po53  & n1540;
  assign n1549 = ~n1547 & ~n1548;
  assign n1550 = ~n1541 & ~n1549;
  assign n1551 = po54  & ~n1550;
  assign n1552 = ~n1368 & ~n1375;
  assign n1553 = n1374 & n1552;
  assign n1554 = po48  & n1553;
  assign n1555 = po48  & n1552;
  assign n1556 = ~n1374 & ~n1555;
  assign n1557 = ~n1554 & ~n1556;
  assign n1558 = ~po54  & ~n1541;
  assign n1559 = ~n1549 & n1558;
  assign n1560 = ~n1557 & ~n1559;
  assign n1561 = ~n1551 & ~n1560;
  assign n1562 = po55  & ~n1561;
  assign n1563 = ~n1378 & ~n1386;
  assign n1564 = n1384 & n1563;
  assign n1565 = po48  & n1564;
  assign n1566 = po48  & n1563;
  assign n1567 = ~n1384 & ~n1566;
  assign n1568 = ~n1565 & ~n1567;
  assign n1569 = ~po55  & n1561;
  assign n1570 = ~n1568 & ~n1569;
  assign n1571 = ~n1562 & ~n1570;
  assign n1572 = po56  & ~n1571;
  assign n1573 = ~n1389 & ~n1396;
  assign n1574 = n1395 & n1573;
  assign n1575 = po48  & n1574;
  assign n1576 = po48  & n1573;
  assign n1577 = ~n1395 & ~n1576;
  assign n1578 = ~n1575 & ~n1577;
  assign n1579 = ~po56  & ~n1562;
  assign n1580 = ~n1570 & n1579;
  assign n1581 = ~n1578 & ~n1580;
  assign n1582 = ~n1572 & ~n1581;
  assign n1583 = po57  & ~n1582;
  assign n1584 = ~n1399 & ~n1407;
  assign n1585 = n1405 & n1584;
  assign n1586 = po48  & n1585;
  assign n1587 = po48  & n1584;
  assign n1588 = ~n1405 & ~n1587;
  assign n1589 = ~n1586 & ~n1588;
  assign n1590 = ~po57  & n1582;
  assign n1591 = ~n1589 & ~n1590;
  assign n1592 = ~n1583 & ~n1591;
  assign n1593 = po58  & ~n1592;
  assign n1594 = ~n1410 & ~n1417;
  assign n1595 = n1416 & n1594;
  assign n1596 = po48  & n1595;
  assign n1597 = po48  & n1594;
  assign n1598 = ~n1416 & ~n1597;
  assign n1599 = ~n1596 & ~n1598;
  assign n1600 = ~po58  & ~n1583;
  assign n1601 = ~n1591 & n1600;
  assign n1602 = ~n1599 & ~n1601;
  assign n1603 = ~n1593 & ~n1602;
  assign n1604 = po59  & ~n1603;
  assign n1605 = ~n1420 & ~n1428;
  assign n1606 = n1426 & n1605;
  assign n1607 = po48  & n1606;
  assign n1608 = po48  & n1605;
  assign n1609 = ~n1426 & ~n1608;
  assign n1610 = ~n1607 & ~n1609;
  assign n1611 = ~po59  & n1603;
  assign n1612 = ~n1610 & ~n1611;
  assign n1613 = ~n1604 & ~n1612;
  assign n1614 = po60  & ~n1613;
  assign n1615 = ~n1431 & ~n1438;
  assign n1616 = n1437 & n1615;
  assign n1617 = po48  & n1616;
  assign n1618 = po48  & n1615;
  assign n1619 = ~n1437 & ~n1618;
  assign n1620 = ~n1617 & ~n1619;
  assign n1621 = ~po60  & ~n1604;
  assign n1622 = ~n1612 & n1621;
  assign n1623 = ~n1620 & ~n1622;
  assign n1624 = ~n1614 & ~n1623;
  assign n1625 = po61  & ~n1624;
  assign n1626 = ~n1441 & ~n1449;
  assign n1627 = n1447 & n1626;
  assign n1628 = po48  & n1627;
  assign n1629 = po48  & n1626;
  assign n1630 = ~n1447 & ~n1629;
  assign n1631 = ~n1628 & ~n1630;
  assign n1632 = ~po61  & n1624;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = ~n1625 & ~n1633;
  assign n1635 = po62  & ~n1634;
  assign n1636 = ~n1452 & ~n1459;
  assign n1637 = n1458 & n1636;
  assign n1638 = po48  & n1637;
  assign n1639 = po48  & n1636;
  assign n1640 = ~n1458 & ~n1639;
  assign n1641 = ~n1638 & ~n1640;
  assign n1642 = ~po62  & ~n1625;
  assign n1643 = ~n1633 & n1642;
  assign n1644 = ~n1641 & ~n1643;
  assign n1645 = ~n1635 & ~n1644;
  assign n1646 = ~n1462 & ~n1470;
  assign n1647 = po48  & n1646;
  assign n1648 = ~n1468 & ~n1647;
  assign n1649 = n1468 & n1647;
  assign n1650 = ~n1648 & ~n1649;
  assign n1651 = ~n1472 & ~n1477;
  assign n1652 = po48  & n1651;
  assign n1653 = ~n1490 & ~n1652;
  assign n1654 = ~n1650 & n1653;
  assign n1655 = ~n1645 & n1654;
  assign n1656 = ~po63  & ~n1655;
  assign n1657 = ~n1477 & po48 ;
  assign n1658 = n1472 & ~n1657;
  assign n1659 = po63  & ~n1651;
  assign n1660 = ~n1658 & n1659;
  assign n1661 = n1477 & ~po48 ;
  assign n1662 = ~n1660 & ~n1661;
  assign n1663 = n1645 & n1650;
  assign n1664 = n1662 & ~n1663;
  assign po47  = n1656 | ~n1664;
  assign n1666 = pi94  & po47 ;
  assign n1667 = ~pi92  & ~pi93 ;
  assign n1668 = ~pi94  & n1667;
  assign n1669 = ~n1666 & ~n1668;
  assign n1670 = po48  & ~n1669;
  assign n1671 = n1489 & ~n1668;
  assign n1672 = ~n1490 & n1671;
  assign n1673 = ~n1483 & n1672;
  assign n1674 = ~n1666 & n1673;
  assign n1675 = ~pi94  & po47 ;
  assign n1676 = pi95  & ~n1675;
  assign n1677 = n1494 & po47 ;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = ~n1674 & n1678;
  assign n1680 = ~n1670 & ~n1679;
  assign n1681 = po49  & ~n1680;
  assign n1682 = po48  & n1662;
  assign n1683 = ~n1663 & n1682;
  assign n1684 = ~n1656 & n1683;
  assign n1685 = ~n1677 & ~n1684;
  assign n1686 = pi96  & ~n1685;
  assign n1687 = ~pi96  & n1685;
  assign n1688 = ~n1686 & ~n1687;
  assign n1689 = ~po49  & n1680;
  assign n1690 = ~n1688 & ~n1689;
  assign n1691 = ~n1681 & ~n1690;
  assign n1692 = po50  & ~n1691;
  assign n1693 = ~po50  & ~n1681;
  assign n1694 = ~n1690 & n1693;
  assign n1695 = ~n1497 & ~n1505;
  assign n1696 = ~n1501 & n1695;
  assign n1697 = po47  & n1696;
  assign n1698 = po47  & n1695;
  assign n1699 = n1501 & ~n1698;
  assign n1700 = ~n1697 & ~n1699;
  assign n1701 = ~n1694 & ~n1700;
  assign n1702 = ~n1692 & ~n1701;
  assign n1703 = po51  & ~n1702;
  assign n1704 = ~n1508 & ~n1510;
  assign n1705 = n1517 & n1704;
  assign n1706 = po47  & n1705;
  assign n1707 = po47  & n1704;
  assign n1708 = ~n1517 & ~n1707;
  assign n1709 = ~n1706 & ~n1708;
  assign n1710 = ~po51  & n1702;
  assign n1711 = ~n1709 & ~n1710;
  assign n1712 = ~n1703 & ~n1711;
  assign n1713 = po52  & ~n1712;
  assign n1714 = ~n1520 & ~n1527;
  assign n1715 = n1526 & n1714;
  assign n1716 = po47  & n1715;
  assign n1717 = po47  & n1714;
  assign n1718 = ~n1526 & ~n1717;
  assign n1719 = ~n1716 & ~n1718;
  assign n1720 = ~po52  & ~n1703;
  assign n1721 = ~n1711 & n1720;
  assign n1722 = ~n1719 & ~n1721;
  assign n1723 = ~n1713 & ~n1722;
  assign n1724 = po53  & ~n1723;
  assign n1725 = ~n1530 & ~n1538;
  assign n1726 = n1536 & n1725;
  assign n1727 = po47  & n1726;
  assign n1728 = po47  & n1725;
  assign n1729 = ~n1536 & ~n1728;
  assign n1730 = ~n1727 & ~n1729;
  assign n1731 = ~po53  & n1723;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = ~n1724 & ~n1732;
  assign n1734 = po54  & ~n1733;
  assign n1735 = ~n1541 & ~n1548;
  assign n1736 = n1547 & n1735;
  assign n1737 = po47  & n1736;
  assign n1738 = po47  & n1735;
  assign n1739 = ~n1547 & ~n1738;
  assign n1740 = ~n1737 & ~n1739;
  assign n1741 = ~po54  & ~n1724;
  assign n1742 = ~n1732 & n1741;
  assign n1743 = ~n1740 & ~n1742;
  assign n1744 = ~n1734 & ~n1743;
  assign n1745 = po55  & ~n1744;
  assign n1746 = ~n1551 & ~n1559;
  assign n1747 = n1557 & n1746;
  assign n1748 = po47  & n1747;
  assign n1749 = po47  & n1746;
  assign n1750 = ~n1557 & ~n1749;
  assign n1751 = ~n1748 & ~n1750;
  assign n1752 = ~po55  & n1744;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = ~n1745 & ~n1753;
  assign n1755 = po56  & ~n1754;
  assign n1756 = ~n1562 & ~n1569;
  assign n1757 = n1568 & n1756;
  assign n1758 = po47  & n1757;
  assign n1759 = po47  & n1756;
  assign n1760 = ~n1568 & ~n1759;
  assign n1761 = ~n1758 & ~n1760;
  assign n1762 = ~po56  & ~n1745;
  assign n1763 = ~n1753 & n1762;
  assign n1764 = ~n1761 & ~n1763;
  assign n1765 = ~n1755 & ~n1764;
  assign n1766 = po57  & ~n1765;
  assign n1767 = ~n1572 & ~n1580;
  assign n1768 = n1578 & n1767;
  assign n1769 = po47  & n1768;
  assign n1770 = po47  & n1767;
  assign n1771 = ~n1578 & ~n1770;
  assign n1772 = ~n1769 & ~n1771;
  assign n1773 = ~po57  & n1765;
  assign n1774 = ~n1772 & ~n1773;
  assign n1775 = ~n1766 & ~n1774;
  assign n1776 = po58  & ~n1775;
  assign n1777 = ~n1583 & ~n1590;
  assign n1778 = n1589 & n1777;
  assign n1779 = po47  & n1778;
  assign n1780 = po47  & n1777;
  assign n1781 = ~n1589 & ~n1780;
  assign n1782 = ~n1779 & ~n1781;
  assign n1783 = ~po58  & ~n1766;
  assign n1784 = ~n1774 & n1783;
  assign n1785 = ~n1782 & ~n1784;
  assign n1786 = ~n1776 & ~n1785;
  assign n1787 = po59  & ~n1786;
  assign n1788 = ~n1593 & ~n1601;
  assign n1789 = n1599 & n1788;
  assign n1790 = po47  & n1789;
  assign n1791 = po47  & n1788;
  assign n1792 = ~n1599 & ~n1791;
  assign n1793 = ~n1790 & ~n1792;
  assign n1794 = ~po59  & n1786;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = ~n1787 & ~n1795;
  assign n1797 = po60  & ~n1796;
  assign n1798 = ~n1604 & ~n1611;
  assign n1799 = n1610 & n1798;
  assign n1800 = po47  & n1799;
  assign n1801 = po47  & n1798;
  assign n1802 = ~n1610 & ~n1801;
  assign n1803 = ~n1800 & ~n1802;
  assign n1804 = ~po60  & ~n1787;
  assign n1805 = ~n1795 & n1804;
  assign n1806 = ~n1803 & ~n1805;
  assign n1807 = ~n1797 & ~n1806;
  assign n1808 = po61  & ~n1807;
  assign n1809 = ~n1614 & ~n1622;
  assign n1810 = n1620 & n1809;
  assign n1811 = po47  & n1810;
  assign n1812 = po47  & n1809;
  assign n1813 = ~n1620 & ~n1812;
  assign n1814 = ~n1811 & ~n1813;
  assign n1815 = ~po61  & n1807;
  assign n1816 = ~n1814 & ~n1815;
  assign n1817 = ~n1808 & ~n1816;
  assign n1818 = po62  & ~n1817;
  assign n1819 = ~n1625 & ~n1632;
  assign n1820 = n1631 & n1819;
  assign n1821 = po47  & n1820;
  assign n1822 = po47  & n1819;
  assign n1823 = ~n1631 & ~n1822;
  assign n1824 = ~n1821 & ~n1823;
  assign n1825 = ~po62  & ~n1808;
  assign n1826 = ~n1816 & n1825;
  assign n1827 = ~n1824 & ~n1826;
  assign n1828 = ~n1818 & ~n1827;
  assign n1829 = ~n1635 & ~n1643;
  assign n1830 = po47  & n1829;
  assign n1831 = ~n1641 & ~n1830;
  assign n1832 = n1641 & n1830;
  assign n1833 = ~n1831 & ~n1832;
  assign n1834 = ~n1645 & ~n1650;
  assign n1835 = po47  & n1834;
  assign n1836 = ~n1663 & ~n1835;
  assign n1837 = ~n1833 & n1836;
  assign n1838 = ~n1828 & n1837;
  assign n1839 = ~po63  & ~n1838;
  assign n1840 = ~n1650 & po47 ;
  assign n1841 = n1645 & ~n1840;
  assign n1842 = po63  & ~n1834;
  assign n1843 = ~n1841 & n1842;
  assign n1844 = n1650 & ~po47 ;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = n1828 & n1833;
  assign n1847 = n1845 & ~n1846;
  assign po46  = n1839 | ~n1847;
  assign n1849 = pi92  & po46 ;
  assign n1850 = ~pi90  & ~pi91 ;
  assign n1851 = ~pi92  & n1850;
  assign n1852 = ~n1849 & ~n1851;
  assign n1853 = po47  & ~n1852;
  assign n1854 = n1662 & ~n1851;
  assign n1855 = ~n1663 & n1854;
  assign n1856 = ~n1656 & n1855;
  assign n1857 = ~n1849 & n1856;
  assign n1858 = ~pi92  & po46 ;
  assign n1859 = pi93  & ~n1858;
  assign n1860 = n1667 & po46 ;
  assign n1861 = ~n1859 & ~n1860;
  assign n1862 = ~n1857 & n1861;
  assign n1863 = ~n1853 & ~n1862;
  assign n1864 = po48  & ~n1863;
  assign n1865 = ~po48  & ~n1853;
  assign n1866 = ~n1862 & n1865;
  assign n1867 = po47  & n1845;
  assign n1868 = ~n1846 & n1867;
  assign n1869 = ~n1839 & n1868;
  assign n1870 = ~n1860 & ~n1869;
  assign n1871 = pi94  & ~n1870;
  assign n1872 = ~pi94  & n1870;
  assign n1873 = ~n1871 & ~n1872;
  assign n1874 = ~n1866 & ~n1873;
  assign n1875 = ~n1864 & ~n1874;
  assign n1876 = po49  & ~n1875;
  assign n1877 = ~n1670 & ~n1674;
  assign n1878 = ~n1678 & n1877;
  assign n1879 = po46  & n1878;
  assign n1880 = po46  & n1877;
  assign n1881 = n1678 & ~n1880;
  assign n1882 = ~n1879 & ~n1881;
  assign n1883 = ~po49  & n1875;
  assign n1884 = ~n1882 & ~n1883;
  assign n1885 = ~n1876 & ~n1884;
  assign n1886 = po50  & ~n1885;
  assign n1887 = ~n1681 & ~n1689;
  assign n1888 = n1688 & n1887;
  assign n1889 = po46  & n1888;
  assign n1890 = po46  & n1887;
  assign n1891 = ~n1688 & ~n1890;
  assign n1892 = ~n1889 & ~n1891;
  assign n1893 = ~po50  & ~n1876;
  assign n1894 = ~n1884 & n1893;
  assign n1895 = ~n1892 & ~n1894;
  assign n1896 = ~n1886 & ~n1895;
  assign n1897 = po51  & ~n1896;
  assign n1898 = ~n1692 & ~n1694;
  assign n1899 = n1700 & n1898;
  assign n1900 = po46  & n1899;
  assign n1901 = po46  & n1898;
  assign n1902 = ~n1700 & ~n1901;
  assign n1903 = ~n1900 & ~n1902;
  assign n1904 = ~po51  & n1896;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = ~n1897 & ~n1905;
  assign n1907 = po52  & ~n1906;
  assign n1908 = ~n1703 & ~n1710;
  assign n1909 = n1709 & n1908;
  assign n1910 = po46  & n1909;
  assign n1911 = po46  & n1908;
  assign n1912 = ~n1709 & ~n1911;
  assign n1913 = ~n1910 & ~n1912;
  assign n1914 = ~po52  & ~n1897;
  assign n1915 = ~n1905 & n1914;
  assign n1916 = ~n1913 & ~n1915;
  assign n1917 = ~n1907 & ~n1916;
  assign n1918 = po53  & ~n1917;
  assign n1919 = ~n1713 & ~n1721;
  assign n1920 = n1719 & n1919;
  assign n1921 = po46  & n1920;
  assign n1922 = po46  & n1919;
  assign n1923 = ~n1719 & ~n1922;
  assign n1924 = ~n1921 & ~n1923;
  assign n1925 = ~po53  & n1917;
  assign n1926 = ~n1924 & ~n1925;
  assign n1927 = ~n1918 & ~n1926;
  assign n1928 = po54  & ~n1927;
  assign n1929 = ~n1724 & ~n1731;
  assign n1930 = n1730 & n1929;
  assign n1931 = po46  & n1930;
  assign n1932 = po46  & n1929;
  assign n1933 = ~n1730 & ~n1932;
  assign n1934 = ~n1931 & ~n1933;
  assign n1935 = ~po54  & ~n1918;
  assign n1936 = ~n1926 & n1935;
  assign n1937 = ~n1934 & ~n1936;
  assign n1938 = ~n1928 & ~n1937;
  assign n1939 = po55  & ~n1938;
  assign n1940 = ~n1734 & ~n1742;
  assign n1941 = n1740 & n1940;
  assign n1942 = po46  & n1941;
  assign n1943 = po46  & n1940;
  assign n1944 = ~n1740 & ~n1943;
  assign n1945 = ~n1942 & ~n1944;
  assign n1946 = ~po55  & n1938;
  assign n1947 = ~n1945 & ~n1946;
  assign n1948 = ~n1939 & ~n1947;
  assign n1949 = po56  & ~n1948;
  assign n1950 = ~n1745 & ~n1752;
  assign n1951 = n1751 & n1950;
  assign n1952 = po46  & n1951;
  assign n1953 = po46  & n1950;
  assign n1954 = ~n1751 & ~n1953;
  assign n1955 = ~n1952 & ~n1954;
  assign n1956 = ~po56  & ~n1939;
  assign n1957 = ~n1947 & n1956;
  assign n1958 = ~n1955 & ~n1957;
  assign n1959 = ~n1949 & ~n1958;
  assign n1960 = po57  & ~n1959;
  assign n1961 = ~n1755 & ~n1763;
  assign n1962 = n1761 & n1961;
  assign n1963 = po46  & n1962;
  assign n1964 = po46  & n1961;
  assign n1965 = ~n1761 & ~n1964;
  assign n1966 = ~n1963 & ~n1965;
  assign n1967 = ~po57  & n1959;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = ~n1960 & ~n1968;
  assign n1970 = po58  & ~n1969;
  assign n1971 = ~n1766 & ~n1773;
  assign n1972 = n1772 & n1971;
  assign n1973 = po46  & n1972;
  assign n1974 = po46  & n1971;
  assign n1975 = ~n1772 & ~n1974;
  assign n1976 = ~n1973 & ~n1975;
  assign n1977 = ~po58  & ~n1960;
  assign n1978 = ~n1968 & n1977;
  assign n1979 = ~n1976 & ~n1978;
  assign n1980 = ~n1970 & ~n1979;
  assign n1981 = po59  & ~n1980;
  assign n1982 = ~n1776 & ~n1784;
  assign n1983 = n1782 & n1982;
  assign n1984 = po46  & n1983;
  assign n1985 = po46  & n1982;
  assign n1986 = ~n1782 & ~n1985;
  assign n1987 = ~n1984 & ~n1986;
  assign n1988 = ~po59  & n1980;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = ~n1981 & ~n1989;
  assign n1991 = po60  & ~n1990;
  assign n1992 = ~n1787 & ~n1794;
  assign n1993 = n1793 & n1992;
  assign n1994 = po46  & n1993;
  assign n1995 = po46  & n1992;
  assign n1996 = ~n1793 & ~n1995;
  assign n1997 = ~n1994 & ~n1996;
  assign n1998 = ~po60  & ~n1981;
  assign n1999 = ~n1989 & n1998;
  assign n2000 = ~n1997 & ~n1999;
  assign n2001 = ~n1991 & ~n2000;
  assign n2002 = po61  & ~n2001;
  assign n2003 = ~n1797 & ~n1805;
  assign n2004 = n1803 & n2003;
  assign n2005 = po46  & n2004;
  assign n2006 = po46  & n2003;
  assign n2007 = ~n1803 & ~n2006;
  assign n2008 = ~n2005 & ~n2007;
  assign n2009 = ~po61  & n2001;
  assign n2010 = ~n2008 & ~n2009;
  assign n2011 = ~n2002 & ~n2010;
  assign n2012 = po62  & ~n2011;
  assign n2013 = ~n1808 & ~n1815;
  assign n2014 = n1814 & n2013;
  assign n2015 = po46  & n2014;
  assign n2016 = po46  & n2013;
  assign n2017 = ~n1814 & ~n2016;
  assign n2018 = ~n2015 & ~n2017;
  assign n2019 = ~po62  & ~n2002;
  assign n2020 = ~n2010 & n2019;
  assign n2021 = ~n2018 & ~n2020;
  assign n2022 = ~n2012 & ~n2021;
  assign n2023 = ~n1818 & ~n1826;
  assign n2024 = po46  & n2023;
  assign n2025 = ~n1824 & ~n2024;
  assign n2026 = n1824 & n2024;
  assign n2027 = ~n2025 & ~n2026;
  assign n2028 = ~n1828 & ~n1833;
  assign n2029 = po46  & n2028;
  assign n2030 = ~n1846 & ~n2029;
  assign n2031 = ~n2027 & n2030;
  assign n2032 = ~n2022 & n2031;
  assign n2033 = ~po63  & ~n2032;
  assign n2034 = ~n1833 & po46 ;
  assign n2035 = n1828 & ~n2034;
  assign n2036 = po63  & ~n2028;
  assign n2037 = ~n2035 & n2036;
  assign n2038 = n1833 & ~po46 ;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = n2022 & n2027;
  assign n2041 = n2039 & ~n2040;
  assign po45  = n2033 | ~n2041;
  assign n2043 = pi90  & po45 ;
  assign n2044 = ~pi88  & ~pi89 ;
  assign n2045 = ~pi90  & n2044;
  assign n2046 = ~n2043 & ~n2045;
  assign n2047 = po46  & ~n2046;
  assign n2048 = n1845 & ~n2045;
  assign n2049 = ~n1846 & n2048;
  assign n2050 = ~n1839 & n2049;
  assign n2051 = ~n2043 & n2050;
  assign n2052 = ~pi90  & po45 ;
  assign n2053 = pi91  & ~n2052;
  assign n2054 = n1850 & po45 ;
  assign n2055 = ~n2053 & ~n2054;
  assign n2056 = ~n2051 & n2055;
  assign n2057 = ~n2047 & ~n2056;
  assign n2058 = po47  & ~n2057;
  assign n2059 = po46  & n2039;
  assign n2060 = ~n2040 & n2059;
  assign n2061 = ~n2033 & n2060;
  assign n2062 = ~n2054 & ~n2061;
  assign n2063 = pi92  & ~n2062;
  assign n2064 = ~pi92  & n2062;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = ~po47  & n2057;
  assign n2067 = ~n2065 & ~n2066;
  assign n2068 = ~n2058 & ~n2067;
  assign n2069 = po48  & ~n2068;
  assign n2070 = ~n1853 & ~n1857;
  assign n2071 = ~n1861 & n2070;
  assign n2072 = po45  & n2071;
  assign n2073 = po45  & n2070;
  assign n2074 = n1861 & ~n2073;
  assign n2075 = ~n2072 & ~n2074;
  assign n2076 = ~po48  & ~n2058;
  assign n2077 = ~n2067 & n2076;
  assign n2078 = ~n2075 & ~n2077;
  assign n2079 = ~n2069 & ~n2078;
  assign n2080 = po49  & ~n2079;
  assign n2081 = ~n1864 & ~n1866;
  assign n2082 = n1873 & n2081;
  assign n2083 = po45  & n2082;
  assign n2084 = po45  & n2081;
  assign n2085 = ~n1873 & ~n2084;
  assign n2086 = ~n2083 & ~n2085;
  assign n2087 = ~po49  & n2079;
  assign n2088 = ~n2086 & ~n2087;
  assign n2089 = ~n2080 & ~n2088;
  assign n2090 = po50  & ~n2089;
  assign n2091 = ~n1876 & ~n1883;
  assign n2092 = n1882 & n2091;
  assign n2093 = po45  & n2092;
  assign n2094 = po45  & n2091;
  assign n2095 = ~n1882 & ~n2094;
  assign n2096 = ~n2093 & ~n2095;
  assign n2097 = ~po50  & ~n2080;
  assign n2098 = ~n2088 & n2097;
  assign n2099 = ~n2096 & ~n2098;
  assign n2100 = ~n2090 & ~n2099;
  assign n2101 = po51  & ~n2100;
  assign n2102 = ~n1886 & ~n1894;
  assign n2103 = n1892 & n2102;
  assign n2104 = po45  & n2103;
  assign n2105 = po45  & n2102;
  assign n2106 = ~n1892 & ~n2105;
  assign n2107 = ~n2104 & ~n2106;
  assign n2108 = ~po51  & n2100;
  assign n2109 = ~n2107 & ~n2108;
  assign n2110 = ~n2101 & ~n2109;
  assign n2111 = po52  & ~n2110;
  assign n2112 = ~po52  & ~n2101;
  assign n2113 = ~n2109 & n2112;
  assign n2114 = ~n1897 & ~n1904;
  assign n2115 = n1903 & n2114;
  assign n2116 = po45  & n2115;
  assign n2117 = po45  & n2114;
  assign n2118 = ~n1903 & ~n2117;
  assign n2119 = ~n2116 & ~n2118;
  assign n2120 = ~n2113 & ~n2119;
  assign n2121 = ~n2111 & ~n2120;
  assign n2122 = po53  & ~n2121;
  assign n2123 = ~n1907 & ~n1915;
  assign n2124 = n1913 & n2123;
  assign n2125 = po45  & n2124;
  assign n2126 = po45  & n2123;
  assign n2127 = ~n1913 & ~n2126;
  assign n2128 = ~n2125 & ~n2127;
  assign n2129 = ~po53  & n2121;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = ~n2122 & ~n2130;
  assign n2132 = po54  & ~n2131;
  assign n2133 = ~n1918 & ~n1925;
  assign n2134 = n1924 & n2133;
  assign n2135 = po45  & n2134;
  assign n2136 = po45  & n2133;
  assign n2137 = ~n1924 & ~n2136;
  assign n2138 = ~n2135 & ~n2137;
  assign n2139 = ~po54  & ~n2122;
  assign n2140 = ~n2130 & n2139;
  assign n2141 = ~n2138 & ~n2140;
  assign n2142 = ~n2132 & ~n2141;
  assign n2143 = po55  & ~n2142;
  assign n2144 = ~n1928 & ~n1936;
  assign n2145 = n1934 & n2144;
  assign n2146 = po45  & n2145;
  assign n2147 = po45  & n2144;
  assign n2148 = ~n1934 & ~n2147;
  assign n2149 = ~n2146 & ~n2148;
  assign n2150 = ~po55  & n2142;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = ~n2143 & ~n2151;
  assign n2153 = po56  & ~n2152;
  assign n2154 = ~n1939 & ~n1946;
  assign n2155 = n1945 & n2154;
  assign n2156 = po45  & n2155;
  assign n2157 = po45  & n2154;
  assign n2158 = ~n1945 & ~n2157;
  assign n2159 = ~n2156 & ~n2158;
  assign n2160 = ~po56  & ~n2143;
  assign n2161 = ~n2151 & n2160;
  assign n2162 = ~n2159 & ~n2161;
  assign n2163 = ~n2153 & ~n2162;
  assign n2164 = po57  & ~n2163;
  assign n2165 = ~n1949 & ~n1957;
  assign n2166 = n1955 & n2165;
  assign n2167 = po45  & n2166;
  assign n2168 = po45  & n2165;
  assign n2169 = ~n1955 & ~n2168;
  assign n2170 = ~n2167 & ~n2169;
  assign n2171 = ~po57  & n2163;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173 = ~n2164 & ~n2172;
  assign n2174 = po58  & ~n2173;
  assign n2175 = ~n1960 & ~n1967;
  assign n2176 = n1966 & n2175;
  assign n2177 = po45  & n2176;
  assign n2178 = po45  & n2175;
  assign n2179 = ~n1966 & ~n2178;
  assign n2180 = ~n2177 & ~n2179;
  assign n2181 = ~po58  & ~n2164;
  assign n2182 = ~n2172 & n2181;
  assign n2183 = ~n2180 & ~n2182;
  assign n2184 = ~n2174 & ~n2183;
  assign n2185 = po59  & ~n2184;
  assign n2186 = ~n1970 & ~n1978;
  assign n2187 = n1976 & n2186;
  assign n2188 = po45  & n2187;
  assign n2189 = po45  & n2186;
  assign n2190 = ~n1976 & ~n2189;
  assign n2191 = ~n2188 & ~n2190;
  assign n2192 = ~po59  & n2184;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = ~n2185 & ~n2193;
  assign n2195 = po60  & ~n2194;
  assign n2196 = ~n1981 & ~n1988;
  assign n2197 = n1987 & n2196;
  assign n2198 = po45  & n2197;
  assign n2199 = po45  & n2196;
  assign n2200 = ~n1987 & ~n2199;
  assign n2201 = ~n2198 & ~n2200;
  assign n2202 = ~po60  & ~n2185;
  assign n2203 = ~n2193 & n2202;
  assign n2204 = ~n2201 & ~n2203;
  assign n2205 = ~n2195 & ~n2204;
  assign n2206 = po61  & ~n2205;
  assign n2207 = ~n1991 & ~n1999;
  assign n2208 = n1997 & n2207;
  assign n2209 = po45  & n2208;
  assign n2210 = po45  & n2207;
  assign n2211 = ~n1997 & ~n2210;
  assign n2212 = ~n2209 & ~n2211;
  assign n2213 = ~po61  & n2205;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = ~n2206 & ~n2214;
  assign n2216 = po62  & ~n2215;
  assign n2217 = ~n2002 & ~n2009;
  assign n2218 = n2008 & n2217;
  assign n2219 = po45  & n2218;
  assign n2220 = po45  & n2217;
  assign n2221 = ~n2008 & ~n2220;
  assign n2222 = ~n2219 & ~n2221;
  assign n2223 = ~po62  & ~n2206;
  assign n2224 = ~n2214 & n2223;
  assign n2225 = ~n2222 & ~n2224;
  assign n2226 = ~n2216 & ~n2225;
  assign n2227 = ~n2012 & ~n2020;
  assign n2228 = po45  & n2227;
  assign n2229 = ~n2018 & ~n2228;
  assign n2230 = n2018 & n2228;
  assign n2231 = ~n2229 & ~n2230;
  assign n2232 = ~n2022 & ~n2027;
  assign n2233 = po45  & n2232;
  assign n2234 = ~n2040 & ~n2233;
  assign n2235 = ~n2231 & n2234;
  assign n2236 = ~n2226 & n2235;
  assign n2237 = ~po63  & ~n2236;
  assign n2238 = ~n2027 & po45 ;
  assign n2239 = n2022 & ~n2238;
  assign n2240 = po63  & ~n2232;
  assign n2241 = ~n2239 & n2240;
  assign n2242 = n2027 & ~po45 ;
  assign n2243 = ~n2241 & ~n2242;
  assign n2244 = n2226 & n2231;
  assign n2245 = n2243 & ~n2244;
  assign po44  = n2237 | ~n2245;
  assign n2247 = pi88  & po44 ;
  assign n2248 = ~pi86  & ~pi87 ;
  assign n2249 = ~pi88  & n2248;
  assign n2250 = ~n2247 & ~n2249;
  assign n2251 = po45  & ~n2250;
  assign n2252 = n2039 & ~n2249;
  assign n2253 = ~n2040 & n2252;
  assign n2254 = ~n2033 & n2253;
  assign n2255 = ~n2247 & n2254;
  assign n2256 = ~pi88  & po44 ;
  assign n2257 = pi89  & ~n2256;
  assign n2258 = n2044 & po44 ;
  assign n2259 = ~n2257 & ~n2258;
  assign n2260 = ~n2255 & n2259;
  assign n2261 = ~n2251 & ~n2260;
  assign n2262 = po46  & ~n2261;
  assign n2263 = ~po46  & ~n2251;
  assign n2264 = ~n2260 & n2263;
  assign n2265 = po45  & n2243;
  assign n2266 = ~n2244 & n2265;
  assign n2267 = ~n2237 & n2266;
  assign n2268 = ~n2258 & ~n2267;
  assign n2269 = pi90  & ~n2268;
  assign n2270 = ~pi90  & n2268;
  assign n2271 = ~n2269 & ~n2270;
  assign n2272 = ~n2264 & ~n2271;
  assign n2273 = ~n2262 & ~n2272;
  assign n2274 = po47  & ~n2273;
  assign n2275 = ~n2047 & ~n2051;
  assign n2276 = ~n2055 & n2275;
  assign n2277 = po44  & n2276;
  assign n2278 = po44  & n2275;
  assign n2279 = n2055 & ~n2278;
  assign n2280 = ~n2277 & ~n2279;
  assign n2281 = ~po47  & n2273;
  assign n2282 = ~n2280 & ~n2281;
  assign n2283 = ~n2274 & ~n2282;
  assign n2284 = po48  & ~n2283;
  assign n2285 = ~n2058 & ~n2066;
  assign n2286 = n2065 & n2285;
  assign n2287 = po44  & n2286;
  assign n2288 = po44  & n2285;
  assign n2289 = ~n2065 & ~n2288;
  assign n2290 = ~n2287 & ~n2289;
  assign n2291 = ~po48  & ~n2274;
  assign n2292 = ~n2282 & n2291;
  assign n2293 = ~n2290 & ~n2292;
  assign n2294 = ~n2284 & ~n2293;
  assign n2295 = po49  & ~n2294;
  assign n2296 = ~n2069 & ~n2077;
  assign n2297 = n2075 & n2296;
  assign n2298 = po44  & n2297;
  assign n2299 = po44  & n2296;
  assign n2300 = ~n2075 & ~n2299;
  assign n2301 = ~n2298 & ~n2300;
  assign n2302 = ~po49  & n2294;
  assign n2303 = ~n2301 & ~n2302;
  assign n2304 = ~n2295 & ~n2303;
  assign n2305 = po50  & ~n2304;
  assign n2306 = ~n2080 & ~n2087;
  assign n2307 = n2086 & n2306;
  assign n2308 = po44  & n2307;
  assign n2309 = po44  & n2306;
  assign n2310 = ~n2086 & ~n2309;
  assign n2311 = ~n2308 & ~n2310;
  assign n2312 = ~po50  & ~n2295;
  assign n2313 = ~n2303 & n2312;
  assign n2314 = ~n2311 & ~n2313;
  assign n2315 = ~n2305 & ~n2314;
  assign n2316 = po51  & ~n2315;
  assign n2317 = ~n2090 & ~n2098;
  assign n2318 = n2096 & n2317;
  assign n2319 = po44  & n2318;
  assign n2320 = po44  & n2317;
  assign n2321 = ~n2096 & ~n2320;
  assign n2322 = ~n2319 & ~n2321;
  assign n2323 = ~po51  & n2315;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = ~n2316 & ~n2324;
  assign n2326 = po52  & ~n2325;
  assign n2327 = ~n2101 & ~n2108;
  assign n2328 = n2107 & n2327;
  assign n2329 = po44  & n2328;
  assign n2330 = po44  & n2327;
  assign n2331 = ~n2107 & ~n2330;
  assign n2332 = ~n2329 & ~n2331;
  assign n2333 = ~po52  & ~n2316;
  assign n2334 = ~n2324 & n2333;
  assign n2335 = ~n2332 & ~n2334;
  assign n2336 = ~n2326 & ~n2335;
  assign n2337 = po53  & ~n2336;
  assign n2338 = ~n2111 & ~n2113;
  assign n2339 = n2119 & n2338;
  assign n2340 = po44  & n2339;
  assign n2341 = po44  & n2338;
  assign n2342 = ~n2119 & ~n2341;
  assign n2343 = ~n2340 & ~n2342;
  assign n2344 = ~po53  & n2336;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = ~n2337 & ~n2345;
  assign n2347 = po54  & ~n2346;
  assign n2348 = ~n2122 & ~n2129;
  assign n2349 = n2128 & n2348;
  assign n2350 = po44  & n2349;
  assign n2351 = po44  & n2348;
  assign n2352 = ~n2128 & ~n2351;
  assign n2353 = ~n2350 & ~n2352;
  assign n2354 = ~po54  & ~n2337;
  assign n2355 = ~n2345 & n2354;
  assign n2356 = ~n2353 & ~n2355;
  assign n2357 = ~n2347 & ~n2356;
  assign n2358 = po55  & ~n2357;
  assign n2359 = ~n2132 & ~n2140;
  assign n2360 = n2138 & n2359;
  assign n2361 = po44  & n2360;
  assign n2362 = po44  & n2359;
  assign n2363 = ~n2138 & ~n2362;
  assign n2364 = ~n2361 & ~n2363;
  assign n2365 = ~po55  & n2357;
  assign n2366 = ~n2364 & ~n2365;
  assign n2367 = ~n2358 & ~n2366;
  assign n2368 = po56  & ~n2367;
  assign n2369 = ~n2143 & ~n2150;
  assign n2370 = n2149 & n2369;
  assign n2371 = po44  & n2370;
  assign n2372 = po44  & n2369;
  assign n2373 = ~n2149 & ~n2372;
  assign n2374 = ~n2371 & ~n2373;
  assign n2375 = ~po56  & ~n2358;
  assign n2376 = ~n2366 & n2375;
  assign n2377 = ~n2374 & ~n2376;
  assign n2378 = ~n2368 & ~n2377;
  assign n2379 = po57  & ~n2378;
  assign n2380 = ~n2153 & ~n2161;
  assign n2381 = n2159 & n2380;
  assign n2382 = po44  & n2381;
  assign n2383 = po44  & n2380;
  assign n2384 = ~n2159 & ~n2383;
  assign n2385 = ~n2382 & ~n2384;
  assign n2386 = ~po57  & n2378;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = ~n2379 & ~n2387;
  assign n2389 = po58  & ~n2388;
  assign n2390 = ~n2164 & ~n2171;
  assign n2391 = n2170 & n2390;
  assign n2392 = po44  & n2391;
  assign n2393 = po44  & n2390;
  assign n2394 = ~n2170 & ~n2393;
  assign n2395 = ~n2392 & ~n2394;
  assign n2396 = ~po58  & ~n2379;
  assign n2397 = ~n2387 & n2396;
  assign n2398 = ~n2395 & ~n2397;
  assign n2399 = ~n2389 & ~n2398;
  assign n2400 = po59  & ~n2399;
  assign n2401 = ~n2174 & ~n2182;
  assign n2402 = n2180 & n2401;
  assign n2403 = po44  & n2402;
  assign n2404 = po44  & n2401;
  assign n2405 = ~n2180 & ~n2404;
  assign n2406 = ~n2403 & ~n2405;
  assign n2407 = ~po59  & n2399;
  assign n2408 = ~n2406 & ~n2407;
  assign n2409 = ~n2400 & ~n2408;
  assign n2410 = po60  & ~n2409;
  assign n2411 = ~n2185 & ~n2192;
  assign n2412 = n2191 & n2411;
  assign n2413 = po44  & n2412;
  assign n2414 = po44  & n2411;
  assign n2415 = ~n2191 & ~n2414;
  assign n2416 = ~n2413 & ~n2415;
  assign n2417 = ~po60  & ~n2400;
  assign n2418 = ~n2408 & n2417;
  assign n2419 = ~n2416 & ~n2418;
  assign n2420 = ~n2410 & ~n2419;
  assign n2421 = po61  & ~n2420;
  assign n2422 = ~n2195 & ~n2203;
  assign n2423 = n2201 & n2422;
  assign n2424 = po44  & n2423;
  assign n2425 = po44  & n2422;
  assign n2426 = ~n2201 & ~n2425;
  assign n2427 = ~n2424 & ~n2426;
  assign n2428 = ~po61  & n2420;
  assign n2429 = ~n2427 & ~n2428;
  assign n2430 = ~n2421 & ~n2429;
  assign n2431 = po62  & ~n2430;
  assign n2432 = ~n2206 & ~n2213;
  assign n2433 = n2212 & n2432;
  assign n2434 = po44  & n2433;
  assign n2435 = po44  & n2432;
  assign n2436 = ~n2212 & ~n2435;
  assign n2437 = ~n2434 & ~n2436;
  assign n2438 = ~po62  & ~n2421;
  assign n2439 = ~n2429 & n2438;
  assign n2440 = ~n2437 & ~n2439;
  assign n2441 = ~n2431 & ~n2440;
  assign n2442 = ~n2216 & ~n2224;
  assign n2443 = po44  & n2442;
  assign n2444 = ~n2222 & ~n2443;
  assign n2445 = n2222 & n2443;
  assign n2446 = ~n2444 & ~n2445;
  assign n2447 = ~n2226 & ~n2231;
  assign n2448 = po44  & n2447;
  assign n2449 = ~n2244 & ~n2448;
  assign n2450 = ~n2446 & n2449;
  assign n2451 = ~n2441 & n2450;
  assign n2452 = ~po63  & ~n2451;
  assign n2453 = ~n2231 & po44 ;
  assign n2454 = n2226 & ~n2453;
  assign n2455 = po63  & ~n2447;
  assign n2456 = ~n2454 & n2455;
  assign n2457 = n2231 & ~po44 ;
  assign n2458 = ~n2456 & ~n2457;
  assign n2459 = n2441 & n2446;
  assign n2460 = n2458 & ~n2459;
  assign po43  = n2452 | ~n2460;
  assign n2462 = pi86  & po43 ;
  assign n2463 = ~pi84  & ~pi85 ;
  assign n2464 = ~pi86  & n2463;
  assign n2465 = ~n2462 & ~n2464;
  assign n2466 = po44  & ~n2465;
  assign n2467 = n2243 & ~n2464;
  assign n2468 = ~n2244 & n2467;
  assign n2469 = ~n2237 & n2468;
  assign n2470 = ~n2462 & n2469;
  assign n2471 = ~pi86  & po43 ;
  assign n2472 = pi87  & ~n2471;
  assign n2473 = n2248 & po43 ;
  assign n2474 = ~n2472 & ~n2473;
  assign n2475 = ~n2470 & n2474;
  assign n2476 = ~n2466 & ~n2475;
  assign n2477 = po45  & ~n2476;
  assign n2478 = po44  & n2458;
  assign n2479 = ~n2459 & n2478;
  assign n2480 = ~n2452 & n2479;
  assign n2481 = ~n2473 & ~n2480;
  assign n2482 = pi88  & ~n2481;
  assign n2483 = ~pi88  & n2481;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = ~po45  & n2476;
  assign n2486 = ~n2484 & ~n2485;
  assign n2487 = ~n2477 & ~n2486;
  assign n2488 = po46  & ~n2487;
  assign n2489 = ~n2251 & ~n2255;
  assign n2490 = ~n2259 & n2489;
  assign n2491 = po43  & n2490;
  assign n2492 = po43  & n2489;
  assign n2493 = n2259 & ~n2492;
  assign n2494 = ~n2491 & ~n2493;
  assign n2495 = ~po46  & ~n2477;
  assign n2496 = ~n2486 & n2495;
  assign n2497 = ~n2494 & ~n2496;
  assign n2498 = ~n2488 & ~n2497;
  assign n2499 = po47  & ~n2498;
  assign n2500 = ~n2262 & ~n2264;
  assign n2501 = n2271 & n2500;
  assign n2502 = po43  & n2501;
  assign n2503 = po43  & n2500;
  assign n2504 = ~n2271 & ~n2503;
  assign n2505 = ~n2502 & ~n2504;
  assign n2506 = ~po47  & n2498;
  assign n2507 = ~n2505 & ~n2506;
  assign n2508 = ~n2499 & ~n2507;
  assign n2509 = po48  & ~n2508;
  assign n2510 = ~n2274 & ~n2281;
  assign n2511 = n2280 & n2510;
  assign n2512 = po43  & n2511;
  assign n2513 = po43  & n2510;
  assign n2514 = ~n2280 & ~n2513;
  assign n2515 = ~n2512 & ~n2514;
  assign n2516 = ~po48  & ~n2499;
  assign n2517 = ~n2507 & n2516;
  assign n2518 = ~n2515 & ~n2517;
  assign n2519 = ~n2509 & ~n2518;
  assign n2520 = po49  & ~n2519;
  assign n2521 = ~n2284 & ~n2292;
  assign n2522 = n2290 & n2521;
  assign n2523 = po43  & n2522;
  assign n2524 = po43  & n2521;
  assign n2525 = ~n2290 & ~n2524;
  assign n2526 = ~n2523 & ~n2525;
  assign n2527 = ~po49  & n2519;
  assign n2528 = ~n2526 & ~n2527;
  assign n2529 = ~n2520 & ~n2528;
  assign n2530 = po50  & ~n2529;
  assign n2531 = ~n2295 & ~n2302;
  assign n2532 = n2301 & n2531;
  assign n2533 = po43  & n2532;
  assign n2534 = po43  & n2531;
  assign n2535 = ~n2301 & ~n2534;
  assign n2536 = ~n2533 & ~n2535;
  assign n2537 = ~po50  & ~n2520;
  assign n2538 = ~n2528 & n2537;
  assign n2539 = ~n2536 & ~n2538;
  assign n2540 = ~n2530 & ~n2539;
  assign n2541 = po51  & ~n2540;
  assign n2542 = ~n2305 & ~n2313;
  assign n2543 = n2311 & n2542;
  assign n2544 = po43  & n2543;
  assign n2545 = po43  & n2542;
  assign n2546 = ~n2311 & ~n2545;
  assign n2547 = ~n2544 & ~n2546;
  assign n2548 = ~po51  & n2540;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = ~n2541 & ~n2549;
  assign n2551 = po52  & ~n2550;
  assign n2552 = ~n2316 & ~n2323;
  assign n2553 = n2322 & n2552;
  assign n2554 = po43  & n2553;
  assign n2555 = po43  & n2552;
  assign n2556 = ~n2322 & ~n2555;
  assign n2557 = ~n2554 & ~n2556;
  assign n2558 = ~po52  & ~n2541;
  assign n2559 = ~n2549 & n2558;
  assign n2560 = ~n2557 & ~n2559;
  assign n2561 = ~n2551 & ~n2560;
  assign n2562 = po53  & ~n2561;
  assign n2563 = ~n2326 & ~n2334;
  assign n2564 = n2332 & n2563;
  assign n2565 = po43  & n2564;
  assign n2566 = po43  & n2563;
  assign n2567 = ~n2332 & ~n2566;
  assign n2568 = ~n2565 & ~n2567;
  assign n2569 = ~po53  & n2561;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = ~n2562 & ~n2570;
  assign n2572 = po54  & ~n2571;
  assign n2573 = ~po54  & ~n2562;
  assign n2574 = ~n2570 & n2573;
  assign n2575 = ~n2337 & ~n2344;
  assign n2576 = n2343 & n2575;
  assign n2577 = po43  & n2576;
  assign n2578 = po43  & n2575;
  assign n2579 = ~n2343 & ~n2578;
  assign n2580 = ~n2577 & ~n2579;
  assign n2581 = ~n2574 & ~n2580;
  assign n2582 = ~n2572 & ~n2581;
  assign n2583 = po55  & ~n2582;
  assign n2584 = ~n2347 & ~n2355;
  assign n2585 = n2353 & n2584;
  assign n2586 = po43  & n2585;
  assign n2587 = po43  & n2584;
  assign n2588 = ~n2353 & ~n2587;
  assign n2589 = ~n2586 & ~n2588;
  assign n2590 = ~po55  & n2582;
  assign n2591 = ~n2589 & ~n2590;
  assign n2592 = ~n2583 & ~n2591;
  assign n2593 = po56  & ~n2592;
  assign n2594 = ~n2358 & ~n2365;
  assign n2595 = n2364 & n2594;
  assign n2596 = po43  & n2595;
  assign n2597 = po43  & n2594;
  assign n2598 = ~n2364 & ~n2597;
  assign n2599 = ~n2596 & ~n2598;
  assign n2600 = ~po56  & ~n2583;
  assign n2601 = ~n2591 & n2600;
  assign n2602 = ~n2599 & ~n2601;
  assign n2603 = ~n2593 & ~n2602;
  assign n2604 = po57  & ~n2603;
  assign n2605 = ~n2368 & ~n2376;
  assign n2606 = n2374 & n2605;
  assign n2607 = po43  & n2606;
  assign n2608 = po43  & n2605;
  assign n2609 = ~n2374 & ~n2608;
  assign n2610 = ~n2607 & ~n2609;
  assign n2611 = ~po57  & n2603;
  assign n2612 = ~n2610 & ~n2611;
  assign n2613 = ~n2604 & ~n2612;
  assign n2614 = po58  & ~n2613;
  assign n2615 = ~n2379 & ~n2386;
  assign n2616 = n2385 & n2615;
  assign n2617 = po43  & n2616;
  assign n2618 = po43  & n2615;
  assign n2619 = ~n2385 & ~n2618;
  assign n2620 = ~n2617 & ~n2619;
  assign n2621 = ~po58  & ~n2604;
  assign n2622 = ~n2612 & n2621;
  assign n2623 = ~n2620 & ~n2622;
  assign n2624 = ~n2614 & ~n2623;
  assign n2625 = po59  & ~n2624;
  assign n2626 = ~n2389 & ~n2397;
  assign n2627 = n2395 & n2626;
  assign n2628 = po43  & n2627;
  assign n2629 = po43  & n2626;
  assign n2630 = ~n2395 & ~n2629;
  assign n2631 = ~n2628 & ~n2630;
  assign n2632 = ~po59  & n2624;
  assign n2633 = ~n2631 & ~n2632;
  assign n2634 = ~n2625 & ~n2633;
  assign n2635 = po60  & ~n2634;
  assign n2636 = ~n2400 & ~n2407;
  assign n2637 = n2406 & n2636;
  assign n2638 = po43  & n2637;
  assign n2639 = po43  & n2636;
  assign n2640 = ~n2406 & ~n2639;
  assign n2641 = ~n2638 & ~n2640;
  assign n2642 = ~po60  & ~n2625;
  assign n2643 = ~n2633 & n2642;
  assign n2644 = ~n2641 & ~n2643;
  assign n2645 = ~n2635 & ~n2644;
  assign n2646 = po61  & ~n2645;
  assign n2647 = ~n2410 & ~n2418;
  assign n2648 = n2416 & n2647;
  assign n2649 = po43  & n2648;
  assign n2650 = po43  & n2647;
  assign n2651 = ~n2416 & ~n2650;
  assign n2652 = ~n2649 & ~n2651;
  assign n2653 = ~po61  & n2645;
  assign n2654 = ~n2652 & ~n2653;
  assign n2655 = ~n2646 & ~n2654;
  assign n2656 = po62  & ~n2655;
  assign n2657 = ~n2421 & ~n2428;
  assign n2658 = n2427 & n2657;
  assign n2659 = po43  & n2658;
  assign n2660 = po43  & n2657;
  assign n2661 = ~n2427 & ~n2660;
  assign n2662 = ~n2659 & ~n2661;
  assign n2663 = ~po62  & ~n2646;
  assign n2664 = ~n2654 & n2663;
  assign n2665 = ~n2662 & ~n2664;
  assign n2666 = ~n2656 & ~n2665;
  assign n2667 = ~n2431 & ~n2439;
  assign n2668 = po43  & n2667;
  assign n2669 = ~n2437 & ~n2668;
  assign n2670 = n2437 & n2668;
  assign n2671 = ~n2669 & ~n2670;
  assign n2672 = ~n2441 & ~n2446;
  assign n2673 = po43  & n2672;
  assign n2674 = ~n2459 & ~n2673;
  assign n2675 = ~n2671 & n2674;
  assign n2676 = ~n2666 & n2675;
  assign n2677 = ~po63  & ~n2676;
  assign n2678 = ~n2446 & po43 ;
  assign n2679 = n2441 & ~n2678;
  assign n2680 = po63  & ~n2672;
  assign n2681 = ~n2679 & n2680;
  assign n2682 = n2446 & ~po43 ;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = n2666 & n2671;
  assign n2685 = n2683 & ~n2684;
  assign po42  = n2677 | ~n2685;
  assign n2687 = pi84  & po42 ;
  assign n2688 = ~pi82  & ~pi83 ;
  assign n2689 = ~pi84  & n2688;
  assign n2690 = ~n2687 & ~n2689;
  assign n2691 = po43  & ~n2690;
  assign n2692 = n2458 & ~n2689;
  assign n2693 = ~n2459 & n2692;
  assign n2694 = ~n2452 & n2693;
  assign n2695 = ~n2687 & n2694;
  assign n2696 = ~pi84  & po42 ;
  assign n2697 = pi85  & ~n2696;
  assign n2698 = n2463 & po42 ;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = ~n2695 & n2699;
  assign n2701 = ~n2691 & ~n2700;
  assign n2702 = po44  & ~n2701;
  assign n2703 = ~po44  & ~n2691;
  assign n2704 = ~n2700 & n2703;
  assign n2705 = po43  & n2683;
  assign n2706 = ~n2684 & n2705;
  assign n2707 = ~n2677 & n2706;
  assign n2708 = ~n2698 & ~n2707;
  assign n2709 = pi86  & ~n2708;
  assign n2710 = ~pi86  & n2708;
  assign n2711 = ~n2709 & ~n2710;
  assign n2712 = ~n2704 & ~n2711;
  assign n2713 = ~n2702 & ~n2712;
  assign n2714 = po45  & ~n2713;
  assign n2715 = ~n2466 & ~n2470;
  assign n2716 = ~n2474 & n2715;
  assign n2717 = po42  & n2716;
  assign n2718 = po42  & n2715;
  assign n2719 = n2474 & ~n2718;
  assign n2720 = ~n2717 & ~n2719;
  assign n2721 = ~po45  & n2713;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = ~n2714 & ~n2722;
  assign n2724 = po46  & ~n2723;
  assign n2725 = ~n2477 & ~n2485;
  assign n2726 = n2484 & n2725;
  assign n2727 = po42  & n2726;
  assign n2728 = po42  & n2725;
  assign n2729 = ~n2484 & ~n2728;
  assign n2730 = ~n2727 & ~n2729;
  assign n2731 = ~po46  & ~n2714;
  assign n2732 = ~n2722 & n2731;
  assign n2733 = ~n2730 & ~n2732;
  assign n2734 = ~n2724 & ~n2733;
  assign n2735 = po47  & ~n2734;
  assign n2736 = ~n2488 & ~n2496;
  assign n2737 = n2494 & n2736;
  assign n2738 = po42  & n2737;
  assign n2739 = po42  & n2736;
  assign n2740 = ~n2494 & ~n2739;
  assign n2741 = ~n2738 & ~n2740;
  assign n2742 = ~po47  & n2734;
  assign n2743 = ~n2741 & ~n2742;
  assign n2744 = ~n2735 & ~n2743;
  assign n2745 = po48  & ~n2744;
  assign n2746 = ~n2499 & ~n2506;
  assign n2747 = n2505 & n2746;
  assign n2748 = po42  & n2747;
  assign n2749 = po42  & n2746;
  assign n2750 = ~n2505 & ~n2749;
  assign n2751 = ~n2748 & ~n2750;
  assign n2752 = ~po48  & ~n2735;
  assign n2753 = ~n2743 & n2752;
  assign n2754 = ~n2751 & ~n2753;
  assign n2755 = ~n2745 & ~n2754;
  assign n2756 = po49  & ~n2755;
  assign n2757 = ~n2509 & ~n2517;
  assign n2758 = n2515 & n2757;
  assign n2759 = po42  & n2758;
  assign n2760 = po42  & n2757;
  assign n2761 = ~n2515 & ~n2760;
  assign n2762 = ~n2759 & ~n2761;
  assign n2763 = ~po49  & n2755;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = ~n2756 & ~n2764;
  assign n2766 = po50  & ~n2765;
  assign n2767 = ~n2520 & ~n2527;
  assign n2768 = n2526 & n2767;
  assign n2769 = po42  & n2768;
  assign n2770 = po42  & n2767;
  assign n2771 = ~n2526 & ~n2770;
  assign n2772 = ~n2769 & ~n2771;
  assign n2773 = ~po50  & ~n2756;
  assign n2774 = ~n2764 & n2773;
  assign n2775 = ~n2772 & ~n2774;
  assign n2776 = ~n2766 & ~n2775;
  assign n2777 = po51  & ~n2776;
  assign n2778 = ~n2530 & ~n2538;
  assign n2779 = n2536 & n2778;
  assign n2780 = po42  & n2779;
  assign n2781 = po42  & n2778;
  assign n2782 = ~n2536 & ~n2781;
  assign n2783 = ~n2780 & ~n2782;
  assign n2784 = ~po51  & n2776;
  assign n2785 = ~n2783 & ~n2784;
  assign n2786 = ~n2777 & ~n2785;
  assign n2787 = po52  & ~n2786;
  assign n2788 = ~n2541 & ~n2548;
  assign n2789 = n2547 & n2788;
  assign n2790 = po42  & n2789;
  assign n2791 = po42  & n2788;
  assign n2792 = ~n2547 & ~n2791;
  assign n2793 = ~n2790 & ~n2792;
  assign n2794 = ~po52  & ~n2777;
  assign n2795 = ~n2785 & n2794;
  assign n2796 = ~n2793 & ~n2795;
  assign n2797 = ~n2787 & ~n2796;
  assign n2798 = po53  & ~n2797;
  assign n2799 = ~n2551 & ~n2559;
  assign n2800 = n2557 & n2799;
  assign n2801 = po42  & n2800;
  assign n2802 = po42  & n2799;
  assign n2803 = ~n2557 & ~n2802;
  assign n2804 = ~n2801 & ~n2803;
  assign n2805 = ~po53  & n2797;
  assign n2806 = ~n2804 & ~n2805;
  assign n2807 = ~n2798 & ~n2806;
  assign n2808 = po54  & ~n2807;
  assign n2809 = ~n2562 & ~n2569;
  assign n2810 = n2568 & n2809;
  assign n2811 = po42  & n2810;
  assign n2812 = po42  & n2809;
  assign n2813 = ~n2568 & ~n2812;
  assign n2814 = ~n2811 & ~n2813;
  assign n2815 = ~po54  & ~n2798;
  assign n2816 = ~n2806 & n2815;
  assign n2817 = ~n2814 & ~n2816;
  assign n2818 = ~n2808 & ~n2817;
  assign n2819 = po55  & ~n2818;
  assign n2820 = ~n2572 & ~n2574;
  assign n2821 = n2580 & n2820;
  assign n2822 = po42  & n2821;
  assign n2823 = po42  & n2820;
  assign n2824 = ~n2580 & ~n2823;
  assign n2825 = ~n2822 & ~n2824;
  assign n2826 = ~po55  & n2818;
  assign n2827 = ~n2825 & ~n2826;
  assign n2828 = ~n2819 & ~n2827;
  assign n2829 = po56  & ~n2828;
  assign n2830 = ~n2583 & ~n2590;
  assign n2831 = n2589 & n2830;
  assign n2832 = po42  & n2831;
  assign n2833 = po42  & n2830;
  assign n2834 = ~n2589 & ~n2833;
  assign n2835 = ~n2832 & ~n2834;
  assign n2836 = ~po56  & ~n2819;
  assign n2837 = ~n2827 & n2836;
  assign n2838 = ~n2835 & ~n2837;
  assign n2839 = ~n2829 & ~n2838;
  assign n2840 = po57  & ~n2839;
  assign n2841 = ~n2593 & ~n2601;
  assign n2842 = n2599 & n2841;
  assign n2843 = po42  & n2842;
  assign n2844 = po42  & n2841;
  assign n2845 = ~n2599 & ~n2844;
  assign n2846 = ~n2843 & ~n2845;
  assign n2847 = ~po57  & n2839;
  assign n2848 = ~n2846 & ~n2847;
  assign n2849 = ~n2840 & ~n2848;
  assign n2850 = po58  & ~n2849;
  assign n2851 = ~n2604 & ~n2611;
  assign n2852 = n2610 & n2851;
  assign n2853 = po42  & n2852;
  assign n2854 = po42  & n2851;
  assign n2855 = ~n2610 & ~n2854;
  assign n2856 = ~n2853 & ~n2855;
  assign n2857 = ~po58  & ~n2840;
  assign n2858 = ~n2848 & n2857;
  assign n2859 = ~n2856 & ~n2858;
  assign n2860 = ~n2850 & ~n2859;
  assign n2861 = po59  & ~n2860;
  assign n2862 = ~n2614 & ~n2622;
  assign n2863 = n2620 & n2862;
  assign n2864 = po42  & n2863;
  assign n2865 = po42  & n2862;
  assign n2866 = ~n2620 & ~n2865;
  assign n2867 = ~n2864 & ~n2866;
  assign n2868 = ~po59  & n2860;
  assign n2869 = ~n2867 & ~n2868;
  assign n2870 = ~n2861 & ~n2869;
  assign n2871 = po60  & ~n2870;
  assign n2872 = ~n2625 & ~n2632;
  assign n2873 = n2631 & n2872;
  assign n2874 = po42  & n2873;
  assign n2875 = po42  & n2872;
  assign n2876 = ~n2631 & ~n2875;
  assign n2877 = ~n2874 & ~n2876;
  assign n2878 = ~po60  & ~n2861;
  assign n2879 = ~n2869 & n2878;
  assign n2880 = ~n2877 & ~n2879;
  assign n2881 = ~n2871 & ~n2880;
  assign n2882 = po61  & ~n2881;
  assign n2883 = ~n2635 & ~n2643;
  assign n2884 = n2641 & n2883;
  assign n2885 = po42  & n2884;
  assign n2886 = po42  & n2883;
  assign n2887 = ~n2641 & ~n2886;
  assign n2888 = ~n2885 & ~n2887;
  assign n2889 = ~po61  & n2881;
  assign n2890 = ~n2888 & ~n2889;
  assign n2891 = ~n2882 & ~n2890;
  assign n2892 = po62  & ~n2891;
  assign n2893 = ~n2646 & ~n2653;
  assign n2894 = n2652 & n2893;
  assign n2895 = po42  & n2894;
  assign n2896 = po42  & n2893;
  assign n2897 = ~n2652 & ~n2896;
  assign n2898 = ~n2895 & ~n2897;
  assign n2899 = ~po62  & ~n2882;
  assign n2900 = ~n2890 & n2899;
  assign n2901 = ~n2898 & ~n2900;
  assign n2902 = ~n2892 & ~n2901;
  assign n2903 = ~n2656 & ~n2664;
  assign n2904 = po42  & n2903;
  assign n2905 = ~n2662 & ~n2904;
  assign n2906 = n2662 & n2904;
  assign n2907 = ~n2905 & ~n2906;
  assign n2908 = ~n2666 & ~n2671;
  assign n2909 = po42  & n2908;
  assign n2910 = ~n2684 & ~n2909;
  assign n2911 = ~n2907 & n2910;
  assign n2912 = ~n2902 & n2911;
  assign n2913 = ~po63  & ~n2912;
  assign n2914 = ~n2671 & po42 ;
  assign n2915 = n2666 & ~n2914;
  assign n2916 = po63  & ~n2908;
  assign n2917 = ~n2915 & n2916;
  assign n2918 = n2671 & ~po42 ;
  assign n2919 = ~n2917 & ~n2918;
  assign n2920 = n2902 & n2907;
  assign n2921 = n2919 & ~n2920;
  assign po41  = n2913 | ~n2921;
  assign n2923 = pi82  & po41 ;
  assign n2924 = ~pi80  & ~pi81 ;
  assign n2925 = ~pi82  & n2924;
  assign n2926 = ~n2923 & ~n2925;
  assign n2927 = po42  & ~n2926;
  assign n2928 = n2683 & ~n2925;
  assign n2929 = ~n2684 & n2928;
  assign n2930 = ~n2677 & n2929;
  assign n2931 = ~n2923 & n2930;
  assign n2932 = ~pi82  & po41 ;
  assign n2933 = pi83  & ~n2932;
  assign n2934 = n2688 & po41 ;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = ~n2931 & n2935;
  assign n2937 = ~n2927 & ~n2936;
  assign n2938 = po43  & ~n2937;
  assign n2939 = po42  & n2919;
  assign n2940 = ~n2920 & n2939;
  assign n2941 = ~n2913 & n2940;
  assign n2942 = ~n2934 & ~n2941;
  assign n2943 = pi84  & ~n2942;
  assign n2944 = ~pi84  & n2942;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = ~po43  & n2937;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = ~n2938 & ~n2947;
  assign n2949 = po44  & ~n2948;
  assign n2950 = ~n2691 & ~n2695;
  assign n2951 = ~n2699 & n2950;
  assign n2952 = po41  & n2951;
  assign n2953 = po41  & n2950;
  assign n2954 = n2699 & ~n2953;
  assign n2955 = ~n2952 & ~n2954;
  assign n2956 = ~po44  & ~n2938;
  assign n2957 = ~n2947 & n2956;
  assign n2958 = ~n2955 & ~n2957;
  assign n2959 = ~n2949 & ~n2958;
  assign n2960 = po45  & ~n2959;
  assign n2961 = ~n2702 & ~n2704;
  assign n2962 = n2711 & n2961;
  assign n2963 = po41  & n2962;
  assign n2964 = po41  & n2961;
  assign n2965 = ~n2711 & ~n2964;
  assign n2966 = ~n2963 & ~n2965;
  assign n2967 = ~po45  & n2959;
  assign n2968 = ~n2966 & ~n2967;
  assign n2969 = ~n2960 & ~n2968;
  assign n2970 = po46  & ~n2969;
  assign n2971 = ~n2714 & ~n2721;
  assign n2972 = n2720 & n2971;
  assign n2973 = po41  & n2972;
  assign n2974 = po41  & n2971;
  assign n2975 = ~n2720 & ~n2974;
  assign n2976 = ~n2973 & ~n2975;
  assign n2977 = ~po46  & ~n2960;
  assign n2978 = ~n2968 & n2977;
  assign n2979 = ~n2976 & ~n2978;
  assign n2980 = ~n2970 & ~n2979;
  assign n2981 = po47  & ~n2980;
  assign n2982 = ~n2724 & ~n2732;
  assign n2983 = n2730 & n2982;
  assign n2984 = po41  & n2983;
  assign n2985 = po41  & n2982;
  assign n2986 = ~n2730 & ~n2985;
  assign n2987 = ~n2984 & ~n2986;
  assign n2988 = ~po47  & n2980;
  assign n2989 = ~n2987 & ~n2988;
  assign n2990 = ~n2981 & ~n2989;
  assign n2991 = po48  & ~n2990;
  assign n2992 = ~n2735 & ~n2742;
  assign n2993 = n2741 & n2992;
  assign n2994 = po41  & n2993;
  assign n2995 = po41  & n2992;
  assign n2996 = ~n2741 & ~n2995;
  assign n2997 = ~n2994 & ~n2996;
  assign n2998 = ~po48  & ~n2981;
  assign n2999 = ~n2989 & n2998;
  assign n3000 = ~n2997 & ~n2999;
  assign n3001 = ~n2991 & ~n3000;
  assign n3002 = po49  & ~n3001;
  assign n3003 = ~n2745 & ~n2753;
  assign n3004 = n2751 & n3003;
  assign n3005 = po41  & n3004;
  assign n3006 = po41  & n3003;
  assign n3007 = ~n2751 & ~n3006;
  assign n3008 = ~n3005 & ~n3007;
  assign n3009 = ~po49  & n3001;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = ~n3002 & ~n3010;
  assign n3012 = po50  & ~n3011;
  assign n3013 = ~n2756 & ~n2763;
  assign n3014 = n2762 & n3013;
  assign n3015 = po41  & n3014;
  assign n3016 = po41  & n3013;
  assign n3017 = ~n2762 & ~n3016;
  assign n3018 = ~n3015 & ~n3017;
  assign n3019 = ~po50  & ~n3002;
  assign n3020 = ~n3010 & n3019;
  assign n3021 = ~n3018 & ~n3020;
  assign n3022 = ~n3012 & ~n3021;
  assign n3023 = po51  & ~n3022;
  assign n3024 = ~n2766 & ~n2774;
  assign n3025 = n2772 & n3024;
  assign n3026 = po41  & n3025;
  assign n3027 = po41  & n3024;
  assign n3028 = ~n2772 & ~n3027;
  assign n3029 = ~n3026 & ~n3028;
  assign n3030 = ~po51  & n3022;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = ~n3023 & ~n3031;
  assign n3033 = po52  & ~n3032;
  assign n3034 = ~n2777 & ~n2784;
  assign n3035 = n2783 & n3034;
  assign n3036 = po41  & n3035;
  assign n3037 = po41  & n3034;
  assign n3038 = ~n2783 & ~n3037;
  assign n3039 = ~n3036 & ~n3038;
  assign n3040 = ~po52  & ~n3023;
  assign n3041 = ~n3031 & n3040;
  assign n3042 = ~n3039 & ~n3041;
  assign n3043 = ~n3033 & ~n3042;
  assign n3044 = po53  & ~n3043;
  assign n3045 = ~n2787 & ~n2795;
  assign n3046 = n2793 & n3045;
  assign n3047 = po41  & n3046;
  assign n3048 = po41  & n3045;
  assign n3049 = ~n2793 & ~n3048;
  assign n3050 = ~n3047 & ~n3049;
  assign n3051 = ~po53  & n3043;
  assign n3052 = ~n3050 & ~n3051;
  assign n3053 = ~n3044 & ~n3052;
  assign n3054 = po54  & ~n3053;
  assign n3055 = ~n2798 & ~n2805;
  assign n3056 = n2804 & n3055;
  assign n3057 = po41  & n3056;
  assign n3058 = po41  & n3055;
  assign n3059 = ~n2804 & ~n3058;
  assign n3060 = ~n3057 & ~n3059;
  assign n3061 = ~po54  & ~n3044;
  assign n3062 = ~n3052 & n3061;
  assign n3063 = ~n3060 & ~n3062;
  assign n3064 = ~n3054 & ~n3063;
  assign n3065 = po55  & ~n3064;
  assign n3066 = ~n2808 & ~n2816;
  assign n3067 = n2814 & n3066;
  assign n3068 = po41  & n3067;
  assign n3069 = po41  & n3066;
  assign n3070 = ~n2814 & ~n3069;
  assign n3071 = ~n3068 & ~n3070;
  assign n3072 = ~po55  & n3064;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = ~n3065 & ~n3073;
  assign n3075 = po56  & ~n3074;
  assign n3076 = ~po56  & ~n3065;
  assign n3077 = ~n3073 & n3076;
  assign n3078 = ~n2819 & ~n2826;
  assign n3079 = n2825 & n3078;
  assign n3080 = po41  & n3079;
  assign n3081 = po41  & n3078;
  assign n3082 = ~n2825 & ~n3081;
  assign n3083 = ~n3080 & ~n3082;
  assign n3084 = ~n3077 & ~n3083;
  assign n3085 = ~n3075 & ~n3084;
  assign n3086 = po57  & ~n3085;
  assign n3087 = ~n2829 & ~n2837;
  assign n3088 = n2835 & n3087;
  assign n3089 = po41  & n3088;
  assign n3090 = po41  & n3087;
  assign n3091 = ~n2835 & ~n3090;
  assign n3092 = ~n3089 & ~n3091;
  assign n3093 = ~po57  & n3085;
  assign n3094 = ~n3092 & ~n3093;
  assign n3095 = ~n3086 & ~n3094;
  assign n3096 = po58  & ~n3095;
  assign n3097 = ~n2840 & ~n2847;
  assign n3098 = n2846 & n3097;
  assign n3099 = po41  & n3098;
  assign n3100 = po41  & n3097;
  assign n3101 = ~n2846 & ~n3100;
  assign n3102 = ~n3099 & ~n3101;
  assign n3103 = ~po58  & ~n3086;
  assign n3104 = ~n3094 & n3103;
  assign n3105 = ~n3102 & ~n3104;
  assign n3106 = ~n3096 & ~n3105;
  assign n3107 = po59  & ~n3106;
  assign n3108 = ~n2850 & ~n2858;
  assign n3109 = n2856 & n3108;
  assign n3110 = po41  & n3109;
  assign n3111 = po41  & n3108;
  assign n3112 = ~n2856 & ~n3111;
  assign n3113 = ~n3110 & ~n3112;
  assign n3114 = ~po59  & n3106;
  assign n3115 = ~n3113 & ~n3114;
  assign n3116 = ~n3107 & ~n3115;
  assign n3117 = po60  & ~n3116;
  assign n3118 = ~n2861 & ~n2868;
  assign n3119 = n2867 & n3118;
  assign n3120 = po41  & n3119;
  assign n3121 = po41  & n3118;
  assign n3122 = ~n2867 & ~n3121;
  assign n3123 = ~n3120 & ~n3122;
  assign n3124 = ~po60  & ~n3107;
  assign n3125 = ~n3115 & n3124;
  assign n3126 = ~n3123 & ~n3125;
  assign n3127 = ~n3117 & ~n3126;
  assign n3128 = po61  & ~n3127;
  assign n3129 = ~n2871 & ~n2879;
  assign n3130 = n2877 & n3129;
  assign n3131 = po41  & n3130;
  assign n3132 = po41  & n3129;
  assign n3133 = ~n2877 & ~n3132;
  assign n3134 = ~n3131 & ~n3133;
  assign n3135 = ~po61  & n3127;
  assign n3136 = ~n3134 & ~n3135;
  assign n3137 = ~n3128 & ~n3136;
  assign n3138 = po62  & ~n3137;
  assign n3139 = ~n2882 & ~n2889;
  assign n3140 = n2888 & n3139;
  assign n3141 = po41  & n3140;
  assign n3142 = po41  & n3139;
  assign n3143 = ~n2888 & ~n3142;
  assign n3144 = ~n3141 & ~n3143;
  assign n3145 = ~po62  & ~n3128;
  assign n3146 = ~n3136 & n3145;
  assign n3147 = ~n3144 & ~n3146;
  assign n3148 = ~n3138 & ~n3147;
  assign n3149 = ~n2892 & ~n2900;
  assign n3150 = po41  & n3149;
  assign n3151 = ~n2898 & ~n3150;
  assign n3152 = n2898 & n3150;
  assign n3153 = ~n3151 & ~n3152;
  assign n3154 = ~n2902 & ~n2907;
  assign n3155 = po41  & n3154;
  assign n3156 = ~n2920 & ~n3155;
  assign n3157 = ~n3153 & n3156;
  assign n3158 = ~n3148 & n3157;
  assign n3159 = ~po63  & ~n3158;
  assign n3160 = ~n2907 & po41 ;
  assign n3161 = n2902 & ~n3160;
  assign n3162 = po63  & ~n3154;
  assign n3163 = ~n3161 & n3162;
  assign n3164 = n2907 & ~po41 ;
  assign n3165 = ~n3163 & ~n3164;
  assign n3166 = n3148 & n3153;
  assign n3167 = n3165 & ~n3166;
  assign po40  = n3159 | ~n3167;
  assign n3169 = pi80  & po40 ;
  assign n3170 = ~pi78  & ~pi79 ;
  assign n3171 = ~pi80  & n3170;
  assign n3172 = ~n3169 & ~n3171;
  assign n3173 = po41  & ~n3172;
  assign n3174 = n2919 & ~n3171;
  assign n3175 = ~n2920 & n3174;
  assign n3176 = ~n2913 & n3175;
  assign n3177 = ~n3169 & n3176;
  assign n3178 = ~pi80  & po40 ;
  assign n3179 = pi81  & ~n3178;
  assign n3180 = n2924 & po40 ;
  assign n3181 = ~n3179 & ~n3180;
  assign n3182 = ~n3177 & n3181;
  assign n3183 = ~n3173 & ~n3182;
  assign n3184 = po42  & ~n3183;
  assign n3185 = ~po42  & ~n3173;
  assign n3186 = ~n3182 & n3185;
  assign n3187 = po41  & n3165;
  assign n3188 = ~n3166 & n3187;
  assign n3189 = ~n3159 & n3188;
  assign n3190 = ~n3180 & ~n3189;
  assign n3191 = pi82  & ~n3190;
  assign n3192 = ~pi82  & n3190;
  assign n3193 = ~n3191 & ~n3192;
  assign n3194 = ~n3186 & ~n3193;
  assign n3195 = ~n3184 & ~n3194;
  assign n3196 = po43  & ~n3195;
  assign n3197 = ~n2927 & ~n2931;
  assign n3198 = ~n2935 & n3197;
  assign n3199 = po40  & n3198;
  assign n3200 = po40  & n3197;
  assign n3201 = n2935 & ~n3200;
  assign n3202 = ~n3199 & ~n3201;
  assign n3203 = ~po43  & n3195;
  assign n3204 = ~n3202 & ~n3203;
  assign n3205 = ~n3196 & ~n3204;
  assign n3206 = po44  & ~n3205;
  assign n3207 = ~n2938 & ~n2946;
  assign n3208 = n2945 & n3207;
  assign n3209 = po40  & n3208;
  assign n3210 = po40  & n3207;
  assign n3211 = ~n2945 & ~n3210;
  assign n3212 = ~n3209 & ~n3211;
  assign n3213 = ~po44  & ~n3196;
  assign n3214 = ~n3204 & n3213;
  assign n3215 = ~n3212 & ~n3214;
  assign n3216 = ~n3206 & ~n3215;
  assign n3217 = po45  & ~n3216;
  assign n3218 = ~n2949 & ~n2957;
  assign n3219 = n2955 & n3218;
  assign n3220 = po40  & n3219;
  assign n3221 = po40  & n3218;
  assign n3222 = ~n2955 & ~n3221;
  assign n3223 = ~n3220 & ~n3222;
  assign n3224 = ~po45  & n3216;
  assign n3225 = ~n3223 & ~n3224;
  assign n3226 = ~n3217 & ~n3225;
  assign n3227 = po46  & ~n3226;
  assign n3228 = ~n2960 & ~n2967;
  assign n3229 = n2966 & n3228;
  assign n3230 = po40  & n3229;
  assign n3231 = po40  & n3228;
  assign n3232 = ~n2966 & ~n3231;
  assign n3233 = ~n3230 & ~n3232;
  assign n3234 = ~po46  & ~n3217;
  assign n3235 = ~n3225 & n3234;
  assign n3236 = ~n3233 & ~n3235;
  assign n3237 = ~n3227 & ~n3236;
  assign n3238 = po47  & ~n3237;
  assign n3239 = ~n2970 & ~n2978;
  assign n3240 = n2976 & n3239;
  assign n3241 = po40  & n3240;
  assign n3242 = po40  & n3239;
  assign n3243 = ~n2976 & ~n3242;
  assign n3244 = ~n3241 & ~n3243;
  assign n3245 = ~po47  & n3237;
  assign n3246 = ~n3244 & ~n3245;
  assign n3247 = ~n3238 & ~n3246;
  assign n3248 = po48  & ~n3247;
  assign n3249 = ~n2981 & ~n2988;
  assign n3250 = n2987 & n3249;
  assign n3251 = po40  & n3250;
  assign n3252 = po40  & n3249;
  assign n3253 = ~n2987 & ~n3252;
  assign n3254 = ~n3251 & ~n3253;
  assign n3255 = ~po48  & ~n3238;
  assign n3256 = ~n3246 & n3255;
  assign n3257 = ~n3254 & ~n3256;
  assign n3258 = ~n3248 & ~n3257;
  assign n3259 = po49  & ~n3258;
  assign n3260 = ~n2991 & ~n2999;
  assign n3261 = n2997 & n3260;
  assign n3262 = po40  & n3261;
  assign n3263 = po40  & n3260;
  assign n3264 = ~n2997 & ~n3263;
  assign n3265 = ~n3262 & ~n3264;
  assign n3266 = ~po49  & n3258;
  assign n3267 = ~n3265 & ~n3266;
  assign n3268 = ~n3259 & ~n3267;
  assign n3269 = po50  & ~n3268;
  assign n3270 = ~n3002 & ~n3009;
  assign n3271 = n3008 & n3270;
  assign n3272 = po40  & n3271;
  assign n3273 = po40  & n3270;
  assign n3274 = ~n3008 & ~n3273;
  assign n3275 = ~n3272 & ~n3274;
  assign n3276 = ~po50  & ~n3259;
  assign n3277 = ~n3267 & n3276;
  assign n3278 = ~n3275 & ~n3277;
  assign n3279 = ~n3269 & ~n3278;
  assign n3280 = po51  & ~n3279;
  assign n3281 = ~n3012 & ~n3020;
  assign n3282 = n3018 & n3281;
  assign n3283 = po40  & n3282;
  assign n3284 = po40  & n3281;
  assign n3285 = ~n3018 & ~n3284;
  assign n3286 = ~n3283 & ~n3285;
  assign n3287 = ~po51  & n3279;
  assign n3288 = ~n3286 & ~n3287;
  assign n3289 = ~n3280 & ~n3288;
  assign n3290 = po52  & ~n3289;
  assign n3291 = ~n3023 & ~n3030;
  assign n3292 = n3029 & n3291;
  assign n3293 = po40  & n3292;
  assign n3294 = po40  & n3291;
  assign n3295 = ~n3029 & ~n3294;
  assign n3296 = ~n3293 & ~n3295;
  assign n3297 = ~po52  & ~n3280;
  assign n3298 = ~n3288 & n3297;
  assign n3299 = ~n3296 & ~n3298;
  assign n3300 = ~n3290 & ~n3299;
  assign n3301 = po53  & ~n3300;
  assign n3302 = ~n3033 & ~n3041;
  assign n3303 = n3039 & n3302;
  assign n3304 = po40  & n3303;
  assign n3305 = po40  & n3302;
  assign n3306 = ~n3039 & ~n3305;
  assign n3307 = ~n3304 & ~n3306;
  assign n3308 = ~po53  & n3300;
  assign n3309 = ~n3307 & ~n3308;
  assign n3310 = ~n3301 & ~n3309;
  assign n3311 = po54  & ~n3310;
  assign n3312 = ~n3044 & ~n3051;
  assign n3313 = n3050 & n3312;
  assign n3314 = po40  & n3313;
  assign n3315 = po40  & n3312;
  assign n3316 = ~n3050 & ~n3315;
  assign n3317 = ~n3314 & ~n3316;
  assign n3318 = ~po54  & ~n3301;
  assign n3319 = ~n3309 & n3318;
  assign n3320 = ~n3317 & ~n3319;
  assign n3321 = ~n3311 & ~n3320;
  assign n3322 = po55  & ~n3321;
  assign n3323 = ~n3054 & ~n3062;
  assign n3324 = n3060 & n3323;
  assign n3325 = po40  & n3324;
  assign n3326 = po40  & n3323;
  assign n3327 = ~n3060 & ~n3326;
  assign n3328 = ~n3325 & ~n3327;
  assign n3329 = ~po55  & n3321;
  assign n3330 = ~n3328 & ~n3329;
  assign n3331 = ~n3322 & ~n3330;
  assign n3332 = po56  & ~n3331;
  assign n3333 = ~n3065 & ~n3072;
  assign n3334 = n3071 & n3333;
  assign n3335 = po40  & n3334;
  assign n3336 = po40  & n3333;
  assign n3337 = ~n3071 & ~n3336;
  assign n3338 = ~n3335 & ~n3337;
  assign n3339 = ~po56  & ~n3322;
  assign n3340 = ~n3330 & n3339;
  assign n3341 = ~n3338 & ~n3340;
  assign n3342 = ~n3332 & ~n3341;
  assign n3343 = po57  & ~n3342;
  assign n3344 = ~n3075 & ~n3077;
  assign n3345 = n3083 & n3344;
  assign n3346 = po40  & n3345;
  assign n3347 = po40  & n3344;
  assign n3348 = ~n3083 & ~n3347;
  assign n3349 = ~n3346 & ~n3348;
  assign n3350 = ~po57  & n3342;
  assign n3351 = ~n3349 & ~n3350;
  assign n3352 = ~n3343 & ~n3351;
  assign n3353 = po58  & ~n3352;
  assign n3354 = ~n3086 & ~n3093;
  assign n3355 = n3092 & n3354;
  assign n3356 = po40  & n3355;
  assign n3357 = po40  & n3354;
  assign n3358 = ~n3092 & ~n3357;
  assign n3359 = ~n3356 & ~n3358;
  assign n3360 = ~po58  & ~n3343;
  assign n3361 = ~n3351 & n3360;
  assign n3362 = ~n3359 & ~n3361;
  assign n3363 = ~n3353 & ~n3362;
  assign n3364 = po59  & ~n3363;
  assign n3365 = ~n3096 & ~n3104;
  assign n3366 = n3102 & n3365;
  assign n3367 = po40  & n3366;
  assign n3368 = po40  & n3365;
  assign n3369 = ~n3102 & ~n3368;
  assign n3370 = ~n3367 & ~n3369;
  assign n3371 = ~po59  & n3363;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = ~n3364 & ~n3372;
  assign n3374 = po60  & ~n3373;
  assign n3375 = ~n3107 & ~n3114;
  assign n3376 = n3113 & n3375;
  assign n3377 = po40  & n3376;
  assign n3378 = po40  & n3375;
  assign n3379 = ~n3113 & ~n3378;
  assign n3380 = ~n3377 & ~n3379;
  assign n3381 = ~po60  & ~n3364;
  assign n3382 = ~n3372 & n3381;
  assign n3383 = ~n3380 & ~n3382;
  assign n3384 = ~n3374 & ~n3383;
  assign n3385 = po61  & ~n3384;
  assign n3386 = ~n3117 & ~n3125;
  assign n3387 = n3123 & n3386;
  assign n3388 = po40  & n3387;
  assign n3389 = po40  & n3386;
  assign n3390 = ~n3123 & ~n3389;
  assign n3391 = ~n3388 & ~n3390;
  assign n3392 = ~po61  & n3384;
  assign n3393 = ~n3391 & ~n3392;
  assign n3394 = ~n3385 & ~n3393;
  assign n3395 = po62  & ~n3394;
  assign n3396 = ~n3128 & ~n3135;
  assign n3397 = n3134 & n3396;
  assign n3398 = po40  & n3397;
  assign n3399 = po40  & n3396;
  assign n3400 = ~n3134 & ~n3399;
  assign n3401 = ~n3398 & ~n3400;
  assign n3402 = ~po62  & ~n3385;
  assign n3403 = ~n3393 & n3402;
  assign n3404 = ~n3401 & ~n3403;
  assign n3405 = ~n3395 & ~n3404;
  assign n3406 = ~n3138 & ~n3146;
  assign n3407 = po40  & n3406;
  assign n3408 = ~n3144 & ~n3407;
  assign n3409 = n3144 & n3407;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = ~n3148 & ~n3153;
  assign n3412 = po40  & n3411;
  assign n3413 = ~n3166 & ~n3412;
  assign n3414 = ~n3410 & n3413;
  assign n3415 = ~n3405 & n3414;
  assign n3416 = ~po63  & ~n3415;
  assign n3417 = ~n3153 & po40 ;
  assign n3418 = n3148 & ~n3417;
  assign n3419 = po63  & ~n3411;
  assign n3420 = ~n3418 & n3419;
  assign n3421 = n3153 & ~po40 ;
  assign n3422 = ~n3420 & ~n3421;
  assign n3423 = n3405 & n3410;
  assign n3424 = n3422 & ~n3423;
  assign po39  = n3416 | ~n3424;
  assign n3426 = pi78  & po39 ;
  assign n3427 = ~pi76  & ~pi77 ;
  assign n3428 = ~pi78  & n3427;
  assign n3429 = ~n3426 & ~n3428;
  assign n3430 = po40  & ~n3429;
  assign n3431 = n3165 & ~n3428;
  assign n3432 = ~n3166 & n3431;
  assign n3433 = ~n3159 & n3432;
  assign n3434 = ~n3426 & n3433;
  assign n3435 = ~pi78  & po39 ;
  assign n3436 = pi79  & ~n3435;
  assign n3437 = n3170 & po39 ;
  assign n3438 = ~n3436 & ~n3437;
  assign n3439 = ~n3434 & n3438;
  assign n3440 = ~n3430 & ~n3439;
  assign n3441 = po41  & ~n3440;
  assign n3442 = po40  & n3422;
  assign n3443 = ~n3423 & n3442;
  assign n3444 = ~n3416 & n3443;
  assign n3445 = ~n3437 & ~n3444;
  assign n3446 = pi80  & ~n3445;
  assign n3447 = ~pi80  & n3445;
  assign n3448 = ~n3446 & ~n3447;
  assign n3449 = ~po41  & n3440;
  assign n3450 = ~n3448 & ~n3449;
  assign n3451 = ~n3441 & ~n3450;
  assign n3452 = po42  & ~n3451;
  assign n3453 = ~n3173 & ~n3177;
  assign n3454 = ~n3181 & n3453;
  assign n3455 = po39  & n3454;
  assign n3456 = po39  & n3453;
  assign n3457 = n3181 & ~n3456;
  assign n3458 = ~n3455 & ~n3457;
  assign n3459 = ~po42  & ~n3441;
  assign n3460 = ~n3450 & n3459;
  assign n3461 = ~n3458 & ~n3460;
  assign n3462 = ~n3452 & ~n3461;
  assign n3463 = po43  & ~n3462;
  assign n3464 = ~n3184 & ~n3186;
  assign n3465 = n3193 & n3464;
  assign n3466 = po39  & n3465;
  assign n3467 = po39  & n3464;
  assign n3468 = ~n3193 & ~n3467;
  assign n3469 = ~n3466 & ~n3468;
  assign n3470 = ~po43  & n3462;
  assign n3471 = ~n3469 & ~n3470;
  assign n3472 = ~n3463 & ~n3471;
  assign n3473 = po44  & ~n3472;
  assign n3474 = ~n3196 & ~n3203;
  assign n3475 = n3202 & n3474;
  assign n3476 = po39  & n3475;
  assign n3477 = po39  & n3474;
  assign n3478 = ~n3202 & ~n3477;
  assign n3479 = ~n3476 & ~n3478;
  assign n3480 = ~po44  & ~n3463;
  assign n3481 = ~n3471 & n3480;
  assign n3482 = ~n3479 & ~n3481;
  assign n3483 = ~n3473 & ~n3482;
  assign n3484 = po45  & ~n3483;
  assign n3485 = ~n3206 & ~n3214;
  assign n3486 = n3212 & n3485;
  assign n3487 = po39  & n3486;
  assign n3488 = po39  & n3485;
  assign n3489 = ~n3212 & ~n3488;
  assign n3490 = ~n3487 & ~n3489;
  assign n3491 = ~po45  & n3483;
  assign n3492 = ~n3490 & ~n3491;
  assign n3493 = ~n3484 & ~n3492;
  assign n3494 = po46  & ~n3493;
  assign n3495 = ~n3217 & ~n3224;
  assign n3496 = n3223 & n3495;
  assign n3497 = po39  & n3496;
  assign n3498 = po39  & n3495;
  assign n3499 = ~n3223 & ~n3498;
  assign n3500 = ~n3497 & ~n3499;
  assign n3501 = ~po46  & ~n3484;
  assign n3502 = ~n3492 & n3501;
  assign n3503 = ~n3500 & ~n3502;
  assign n3504 = ~n3494 & ~n3503;
  assign n3505 = po47  & ~n3504;
  assign n3506 = ~n3227 & ~n3235;
  assign n3507 = n3233 & n3506;
  assign n3508 = po39  & n3507;
  assign n3509 = po39  & n3506;
  assign n3510 = ~n3233 & ~n3509;
  assign n3511 = ~n3508 & ~n3510;
  assign n3512 = ~po47  & n3504;
  assign n3513 = ~n3511 & ~n3512;
  assign n3514 = ~n3505 & ~n3513;
  assign n3515 = po48  & ~n3514;
  assign n3516 = ~n3238 & ~n3245;
  assign n3517 = n3244 & n3516;
  assign n3518 = po39  & n3517;
  assign n3519 = po39  & n3516;
  assign n3520 = ~n3244 & ~n3519;
  assign n3521 = ~n3518 & ~n3520;
  assign n3522 = ~po48  & ~n3505;
  assign n3523 = ~n3513 & n3522;
  assign n3524 = ~n3521 & ~n3523;
  assign n3525 = ~n3515 & ~n3524;
  assign n3526 = po49  & ~n3525;
  assign n3527 = ~n3248 & ~n3256;
  assign n3528 = n3254 & n3527;
  assign n3529 = po39  & n3528;
  assign n3530 = po39  & n3527;
  assign n3531 = ~n3254 & ~n3530;
  assign n3532 = ~n3529 & ~n3531;
  assign n3533 = ~po49  & n3525;
  assign n3534 = ~n3532 & ~n3533;
  assign n3535 = ~n3526 & ~n3534;
  assign n3536 = po50  & ~n3535;
  assign n3537 = ~n3259 & ~n3266;
  assign n3538 = n3265 & n3537;
  assign n3539 = po39  & n3538;
  assign n3540 = po39  & n3537;
  assign n3541 = ~n3265 & ~n3540;
  assign n3542 = ~n3539 & ~n3541;
  assign n3543 = ~po50  & ~n3526;
  assign n3544 = ~n3534 & n3543;
  assign n3545 = ~n3542 & ~n3544;
  assign n3546 = ~n3536 & ~n3545;
  assign n3547 = po51  & ~n3546;
  assign n3548 = ~n3269 & ~n3277;
  assign n3549 = n3275 & n3548;
  assign n3550 = po39  & n3549;
  assign n3551 = po39  & n3548;
  assign n3552 = ~n3275 & ~n3551;
  assign n3553 = ~n3550 & ~n3552;
  assign n3554 = ~po51  & n3546;
  assign n3555 = ~n3553 & ~n3554;
  assign n3556 = ~n3547 & ~n3555;
  assign n3557 = po52  & ~n3556;
  assign n3558 = ~n3280 & ~n3287;
  assign n3559 = n3286 & n3558;
  assign n3560 = po39  & n3559;
  assign n3561 = po39  & n3558;
  assign n3562 = ~n3286 & ~n3561;
  assign n3563 = ~n3560 & ~n3562;
  assign n3564 = ~po52  & ~n3547;
  assign n3565 = ~n3555 & n3564;
  assign n3566 = ~n3563 & ~n3565;
  assign n3567 = ~n3557 & ~n3566;
  assign n3568 = po53  & ~n3567;
  assign n3569 = ~n3290 & ~n3298;
  assign n3570 = n3296 & n3569;
  assign n3571 = po39  & n3570;
  assign n3572 = po39  & n3569;
  assign n3573 = ~n3296 & ~n3572;
  assign n3574 = ~n3571 & ~n3573;
  assign n3575 = ~po53  & n3567;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = ~n3568 & ~n3576;
  assign n3578 = po54  & ~n3577;
  assign n3579 = ~n3301 & ~n3308;
  assign n3580 = n3307 & n3579;
  assign n3581 = po39  & n3580;
  assign n3582 = po39  & n3579;
  assign n3583 = ~n3307 & ~n3582;
  assign n3584 = ~n3581 & ~n3583;
  assign n3585 = ~po54  & ~n3568;
  assign n3586 = ~n3576 & n3585;
  assign n3587 = ~n3584 & ~n3586;
  assign n3588 = ~n3578 & ~n3587;
  assign n3589 = po55  & ~n3588;
  assign n3590 = ~n3311 & ~n3319;
  assign n3591 = n3317 & n3590;
  assign n3592 = po39  & n3591;
  assign n3593 = po39  & n3590;
  assign n3594 = ~n3317 & ~n3593;
  assign n3595 = ~n3592 & ~n3594;
  assign n3596 = ~po55  & n3588;
  assign n3597 = ~n3595 & ~n3596;
  assign n3598 = ~n3589 & ~n3597;
  assign n3599 = po56  & ~n3598;
  assign n3600 = ~n3322 & ~n3329;
  assign n3601 = n3328 & n3600;
  assign n3602 = po39  & n3601;
  assign n3603 = po39  & n3600;
  assign n3604 = ~n3328 & ~n3603;
  assign n3605 = ~n3602 & ~n3604;
  assign n3606 = ~po56  & ~n3589;
  assign n3607 = ~n3597 & n3606;
  assign n3608 = ~n3605 & ~n3607;
  assign n3609 = ~n3599 & ~n3608;
  assign n3610 = po57  & ~n3609;
  assign n3611 = ~n3332 & ~n3340;
  assign n3612 = n3338 & n3611;
  assign n3613 = po39  & n3612;
  assign n3614 = po39  & n3611;
  assign n3615 = ~n3338 & ~n3614;
  assign n3616 = ~n3613 & ~n3615;
  assign n3617 = ~po57  & n3609;
  assign n3618 = ~n3616 & ~n3617;
  assign n3619 = ~n3610 & ~n3618;
  assign n3620 = po58  & ~n3619;
  assign n3621 = ~po58  & ~n3610;
  assign n3622 = ~n3618 & n3621;
  assign n3623 = ~n3343 & ~n3350;
  assign n3624 = n3349 & n3623;
  assign n3625 = po39  & n3624;
  assign n3626 = po39  & n3623;
  assign n3627 = ~n3349 & ~n3626;
  assign n3628 = ~n3625 & ~n3627;
  assign n3629 = ~n3622 & ~n3628;
  assign n3630 = ~n3620 & ~n3629;
  assign n3631 = po59  & ~n3630;
  assign n3632 = ~n3353 & ~n3361;
  assign n3633 = n3359 & n3632;
  assign n3634 = po39  & n3633;
  assign n3635 = po39  & n3632;
  assign n3636 = ~n3359 & ~n3635;
  assign n3637 = ~n3634 & ~n3636;
  assign n3638 = ~po59  & n3630;
  assign n3639 = ~n3637 & ~n3638;
  assign n3640 = ~n3631 & ~n3639;
  assign n3641 = po60  & ~n3640;
  assign n3642 = ~n3364 & ~n3371;
  assign n3643 = n3370 & n3642;
  assign n3644 = po39  & n3643;
  assign n3645 = po39  & n3642;
  assign n3646 = ~n3370 & ~n3645;
  assign n3647 = ~n3644 & ~n3646;
  assign n3648 = ~po60  & ~n3631;
  assign n3649 = ~n3639 & n3648;
  assign n3650 = ~n3647 & ~n3649;
  assign n3651 = ~n3641 & ~n3650;
  assign n3652 = po61  & ~n3651;
  assign n3653 = ~n3374 & ~n3382;
  assign n3654 = n3380 & n3653;
  assign n3655 = po39  & n3654;
  assign n3656 = po39  & n3653;
  assign n3657 = ~n3380 & ~n3656;
  assign n3658 = ~n3655 & ~n3657;
  assign n3659 = ~po61  & n3651;
  assign n3660 = ~n3658 & ~n3659;
  assign n3661 = ~n3652 & ~n3660;
  assign n3662 = po62  & ~n3661;
  assign n3663 = ~n3385 & ~n3392;
  assign n3664 = n3391 & n3663;
  assign n3665 = po39  & n3664;
  assign n3666 = po39  & n3663;
  assign n3667 = ~n3391 & ~n3666;
  assign n3668 = ~n3665 & ~n3667;
  assign n3669 = ~po62  & ~n3652;
  assign n3670 = ~n3660 & n3669;
  assign n3671 = ~n3668 & ~n3670;
  assign n3672 = ~n3662 & ~n3671;
  assign n3673 = ~n3395 & ~n3403;
  assign n3674 = po39  & n3673;
  assign n3675 = ~n3401 & ~n3674;
  assign n3676 = n3401 & n3674;
  assign n3677 = ~n3675 & ~n3676;
  assign n3678 = ~n3405 & ~n3410;
  assign n3679 = po39  & n3678;
  assign n3680 = ~n3423 & ~n3679;
  assign n3681 = ~n3677 & n3680;
  assign n3682 = ~n3672 & n3681;
  assign n3683 = ~po63  & ~n3682;
  assign n3684 = ~n3410 & po39 ;
  assign n3685 = n3405 & ~n3684;
  assign n3686 = po63  & ~n3678;
  assign n3687 = ~n3685 & n3686;
  assign n3688 = n3410 & ~po39 ;
  assign n3689 = ~n3687 & ~n3688;
  assign n3690 = n3672 & n3677;
  assign n3691 = n3689 & ~n3690;
  assign po38  = n3683 | ~n3691;
  assign n3693 = pi76  & po38 ;
  assign n3694 = ~pi74  & ~pi75 ;
  assign n3695 = ~pi76  & n3694;
  assign n3696 = ~n3693 & ~n3695;
  assign n3697 = po39  & ~n3696;
  assign n3698 = n3422 & ~n3695;
  assign n3699 = ~n3423 & n3698;
  assign n3700 = ~n3416 & n3699;
  assign n3701 = ~n3693 & n3700;
  assign n3702 = ~pi76  & po38 ;
  assign n3703 = pi77  & ~n3702;
  assign n3704 = n3427 & po38 ;
  assign n3705 = ~n3703 & ~n3704;
  assign n3706 = ~n3701 & n3705;
  assign n3707 = ~n3697 & ~n3706;
  assign n3708 = po40  & ~n3707;
  assign n3709 = ~po40  & ~n3697;
  assign n3710 = ~n3706 & n3709;
  assign n3711 = po39  & n3689;
  assign n3712 = ~n3690 & n3711;
  assign n3713 = ~n3683 & n3712;
  assign n3714 = ~n3704 & ~n3713;
  assign n3715 = pi78  & ~n3714;
  assign n3716 = ~pi78  & n3714;
  assign n3717 = ~n3715 & ~n3716;
  assign n3718 = ~n3710 & ~n3717;
  assign n3719 = ~n3708 & ~n3718;
  assign n3720 = po41  & ~n3719;
  assign n3721 = ~n3430 & ~n3434;
  assign n3722 = ~n3438 & n3721;
  assign n3723 = po38  & n3722;
  assign n3724 = po38  & n3721;
  assign n3725 = n3438 & ~n3724;
  assign n3726 = ~n3723 & ~n3725;
  assign n3727 = ~po41  & n3719;
  assign n3728 = ~n3726 & ~n3727;
  assign n3729 = ~n3720 & ~n3728;
  assign n3730 = po42  & ~n3729;
  assign n3731 = ~n3441 & ~n3449;
  assign n3732 = n3448 & n3731;
  assign n3733 = po38  & n3732;
  assign n3734 = po38  & n3731;
  assign n3735 = ~n3448 & ~n3734;
  assign n3736 = ~n3733 & ~n3735;
  assign n3737 = ~po42  & ~n3720;
  assign n3738 = ~n3728 & n3737;
  assign n3739 = ~n3736 & ~n3738;
  assign n3740 = ~n3730 & ~n3739;
  assign n3741 = po43  & ~n3740;
  assign n3742 = ~n3452 & ~n3460;
  assign n3743 = n3458 & n3742;
  assign n3744 = po38  & n3743;
  assign n3745 = po38  & n3742;
  assign n3746 = ~n3458 & ~n3745;
  assign n3747 = ~n3744 & ~n3746;
  assign n3748 = ~po43  & n3740;
  assign n3749 = ~n3747 & ~n3748;
  assign n3750 = ~n3741 & ~n3749;
  assign n3751 = po44  & ~n3750;
  assign n3752 = ~n3463 & ~n3470;
  assign n3753 = n3469 & n3752;
  assign n3754 = po38  & n3753;
  assign n3755 = po38  & n3752;
  assign n3756 = ~n3469 & ~n3755;
  assign n3757 = ~n3754 & ~n3756;
  assign n3758 = ~po44  & ~n3741;
  assign n3759 = ~n3749 & n3758;
  assign n3760 = ~n3757 & ~n3759;
  assign n3761 = ~n3751 & ~n3760;
  assign n3762 = po45  & ~n3761;
  assign n3763 = ~n3473 & ~n3481;
  assign n3764 = n3479 & n3763;
  assign n3765 = po38  & n3764;
  assign n3766 = po38  & n3763;
  assign n3767 = ~n3479 & ~n3766;
  assign n3768 = ~n3765 & ~n3767;
  assign n3769 = ~po45  & n3761;
  assign n3770 = ~n3768 & ~n3769;
  assign n3771 = ~n3762 & ~n3770;
  assign n3772 = po46  & ~n3771;
  assign n3773 = ~n3484 & ~n3491;
  assign n3774 = n3490 & n3773;
  assign n3775 = po38  & n3774;
  assign n3776 = po38  & n3773;
  assign n3777 = ~n3490 & ~n3776;
  assign n3778 = ~n3775 & ~n3777;
  assign n3779 = ~po46  & ~n3762;
  assign n3780 = ~n3770 & n3779;
  assign n3781 = ~n3778 & ~n3780;
  assign n3782 = ~n3772 & ~n3781;
  assign n3783 = po47  & ~n3782;
  assign n3784 = ~n3494 & ~n3502;
  assign n3785 = n3500 & n3784;
  assign n3786 = po38  & n3785;
  assign n3787 = po38  & n3784;
  assign n3788 = ~n3500 & ~n3787;
  assign n3789 = ~n3786 & ~n3788;
  assign n3790 = ~po47  & n3782;
  assign n3791 = ~n3789 & ~n3790;
  assign n3792 = ~n3783 & ~n3791;
  assign n3793 = po48  & ~n3792;
  assign n3794 = ~n3505 & ~n3512;
  assign n3795 = n3511 & n3794;
  assign n3796 = po38  & n3795;
  assign n3797 = po38  & n3794;
  assign n3798 = ~n3511 & ~n3797;
  assign n3799 = ~n3796 & ~n3798;
  assign n3800 = ~po48  & ~n3783;
  assign n3801 = ~n3791 & n3800;
  assign n3802 = ~n3799 & ~n3801;
  assign n3803 = ~n3793 & ~n3802;
  assign n3804 = po49  & ~n3803;
  assign n3805 = ~n3515 & ~n3523;
  assign n3806 = n3521 & n3805;
  assign n3807 = po38  & n3806;
  assign n3808 = po38  & n3805;
  assign n3809 = ~n3521 & ~n3808;
  assign n3810 = ~n3807 & ~n3809;
  assign n3811 = ~po49  & n3803;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = ~n3804 & ~n3812;
  assign n3814 = po50  & ~n3813;
  assign n3815 = ~n3526 & ~n3533;
  assign n3816 = n3532 & n3815;
  assign n3817 = po38  & n3816;
  assign n3818 = po38  & n3815;
  assign n3819 = ~n3532 & ~n3818;
  assign n3820 = ~n3817 & ~n3819;
  assign n3821 = ~po50  & ~n3804;
  assign n3822 = ~n3812 & n3821;
  assign n3823 = ~n3820 & ~n3822;
  assign n3824 = ~n3814 & ~n3823;
  assign n3825 = po51  & ~n3824;
  assign n3826 = ~n3536 & ~n3544;
  assign n3827 = n3542 & n3826;
  assign n3828 = po38  & n3827;
  assign n3829 = po38  & n3826;
  assign n3830 = ~n3542 & ~n3829;
  assign n3831 = ~n3828 & ~n3830;
  assign n3832 = ~po51  & n3824;
  assign n3833 = ~n3831 & ~n3832;
  assign n3834 = ~n3825 & ~n3833;
  assign n3835 = po52  & ~n3834;
  assign n3836 = ~n3547 & ~n3554;
  assign n3837 = n3553 & n3836;
  assign n3838 = po38  & n3837;
  assign n3839 = po38  & n3836;
  assign n3840 = ~n3553 & ~n3839;
  assign n3841 = ~n3838 & ~n3840;
  assign n3842 = ~po52  & ~n3825;
  assign n3843 = ~n3833 & n3842;
  assign n3844 = ~n3841 & ~n3843;
  assign n3845 = ~n3835 & ~n3844;
  assign n3846 = po53  & ~n3845;
  assign n3847 = ~n3557 & ~n3565;
  assign n3848 = n3563 & n3847;
  assign n3849 = po38  & n3848;
  assign n3850 = po38  & n3847;
  assign n3851 = ~n3563 & ~n3850;
  assign n3852 = ~n3849 & ~n3851;
  assign n3853 = ~po53  & n3845;
  assign n3854 = ~n3852 & ~n3853;
  assign n3855 = ~n3846 & ~n3854;
  assign n3856 = po54  & ~n3855;
  assign n3857 = ~n3568 & ~n3575;
  assign n3858 = n3574 & n3857;
  assign n3859 = po38  & n3858;
  assign n3860 = po38  & n3857;
  assign n3861 = ~n3574 & ~n3860;
  assign n3862 = ~n3859 & ~n3861;
  assign n3863 = ~po54  & ~n3846;
  assign n3864 = ~n3854 & n3863;
  assign n3865 = ~n3862 & ~n3864;
  assign n3866 = ~n3856 & ~n3865;
  assign n3867 = po55  & ~n3866;
  assign n3868 = ~n3578 & ~n3586;
  assign n3869 = n3584 & n3868;
  assign n3870 = po38  & n3869;
  assign n3871 = po38  & n3868;
  assign n3872 = ~n3584 & ~n3871;
  assign n3873 = ~n3870 & ~n3872;
  assign n3874 = ~po55  & n3866;
  assign n3875 = ~n3873 & ~n3874;
  assign n3876 = ~n3867 & ~n3875;
  assign n3877 = po56  & ~n3876;
  assign n3878 = ~n3589 & ~n3596;
  assign n3879 = n3595 & n3878;
  assign n3880 = po38  & n3879;
  assign n3881 = po38  & n3878;
  assign n3882 = ~n3595 & ~n3881;
  assign n3883 = ~n3880 & ~n3882;
  assign n3884 = ~po56  & ~n3867;
  assign n3885 = ~n3875 & n3884;
  assign n3886 = ~n3883 & ~n3885;
  assign n3887 = ~n3877 & ~n3886;
  assign n3888 = po57  & ~n3887;
  assign n3889 = ~n3599 & ~n3607;
  assign n3890 = n3605 & n3889;
  assign n3891 = po38  & n3890;
  assign n3892 = po38  & n3889;
  assign n3893 = ~n3605 & ~n3892;
  assign n3894 = ~n3891 & ~n3893;
  assign n3895 = ~po57  & n3887;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = ~n3888 & ~n3896;
  assign n3898 = po58  & ~n3897;
  assign n3899 = ~n3610 & ~n3617;
  assign n3900 = n3616 & n3899;
  assign n3901 = po38  & n3900;
  assign n3902 = po38  & n3899;
  assign n3903 = ~n3616 & ~n3902;
  assign n3904 = ~n3901 & ~n3903;
  assign n3905 = ~po58  & ~n3888;
  assign n3906 = ~n3896 & n3905;
  assign n3907 = ~n3904 & ~n3906;
  assign n3908 = ~n3898 & ~n3907;
  assign n3909 = po59  & ~n3908;
  assign n3910 = ~n3620 & ~n3622;
  assign n3911 = n3628 & n3910;
  assign n3912 = po38  & n3911;
  assign n3913 = po38  & n3910;
  assign n3914 = ~n3628 & ~n3913;
  assign n3915 = ~n3912 & ~n3914;
  assign n3916 = ~po59  & n3908;
  assign n3917 = ~n3915 & ~n3916;
  assign n3918 = ~n3909 & ~n3917;
  assign n3919 = po60  & ~n3918;
  assign n3920 = ~n3631 & ~n3638;
  assign n3921 = n3637 & n3920;
  assign n3922 = po38  & n3921;
  assign n3923 = po38  & n3920;
  assign n3924 = ~n3637 & ~n3923;
  assign n3925 = ~n3922 & ~n3924;
  assign n3926 = ~po60  & ~n3909;
  assign n3927 = ~n3917 & n3926;
  assign n3928 = ~n3925 & ~n3927;
  assign n3929 = ~n3919 & ~n3928;
  assign n3930 = po61  & ~n3929;
  assign n3931 = ~n3641 & ~n3649;
  assign n3932 = n3647 & n3931;
  assign n3933 = po38  & n3932;
  assign n3934 = po38  & n3931;
  assign n3935 = ~n3647 & ~n3934;
  assign n3936 = ~n3933 & ~n3935;
  assign n3937 = ~po61  & n3929;
  assign n3938 = ~n3936 & ~n3937;
  assign n3939 = ~n3930 & ~n3938;
  assign n3940 = po62  & ~n3939;
  assign n3941 = ~n3652 & ~n3659;
  assign n3942 = n3658 & n3941;
  assign n3943 = po38  & n3942;
  assign n3944 = po38  & n3941;
  assign n3945 = ~n3658 & ~n3944;
  assign n3946 = ~n3943 & ~n3945;
  assign n3947 = ~po62  & ~n3930;
  assign n3948 = ~n3938 & n3947;
  assign n3949 = ~n3946 & ~n3948;
  assign n3950 = ~n3940 & ~n3949;
  assign n3951 = ~n3662 & ~n3670;
  assign n3952 = po38  & n3951;
  assign n3953 = ~n3668 & ~n3952;
  assign n3954 = n3668 & n3952;
  assign n3955 = ~n3953 & ~n3954;
  assign n3956 = ~n3672 & ~n3677;
  assign n3957 = po38  & n3956;
  assign n3958 = ~n3690 & ~n3957;
  assign n3959 = ~n3955 & n3958;
  assign n3960 = ~n3950 & n3959;
  assign n3961 = ~po63  & ~n3960;
  assign n3962 = ~n3677 & po38 ;
  assign n3963 = n3672 & ~n3962;
  assign n3964 = po63  & ~n3956;
  assign n3965 = ~n3963 & n3964;
  assign n3966 = n3677 & ~po38 ;
  assign n3967 = ~n3965 & ~n3966;
  assign n3968 = n3950 & n3955;
  assign n3969 = n3967 & ~n3968;
  assign po37  = n3961 | ~n3969;
  assign n3971 = pi74  & po37 ;
  assign n3972 = ~pi72  & ~pi73 ;
  assign n3973 = ~pi74  & n3972;
  assign n3974 = ~n3971 & ~n3973;
  assign n3975 = po38  & ~n3974;
  assign n3976 = n3689 & ~n3973;
  assign n3977 = ~n3690 & n3976;
  assign n3978 = ~n3683 & n3977;
  assign n3979 = ~n3971 & n3978;
  assign n3980 = ~pi74  & po37 ;
  assign n3981 = pi75  & ~n3980;
  assign n3982 = n3694 & po37 ;
  assign n3983 = ~n3981 & ~n3982;
  assign n3984 = ~n3979 & n3983;
  assign n3985 = ~n3975 & ~n3984;
  assign n3986 = po39  & ~n3985;
  assign n3987 = po38  & n3967;
  assign n3988 = ~n3968 & n3987;
  assign n3989 = ~n3961 & n3988;
  assign n3990 = ~n3982 & ~n3989;
  assign n3991 = pi76  & ~n3990;
  assign n3992 = ~pi76  & n3990;
  assign n3993 = ~n3991 & ~n3992;
  assign n3994 = ~po39  & n3985;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = ~n3986 & ~n3995;
  assign n3997 = po40  & ~n3996;
  assign n3998 = ~n3697 & ~n3701;
  assign n3999 = ~n3705 & n3998;
  assign n4000 = po37  & n3999;
  assign n4001 = po37  & n3998;
  assign n4002 = n3705 & ~n4001;
  assign n4003 = ~n4000 & ~n4002;
  assign n4004 = ~po40  & ~n3986;
  assign n4005 = ~n3995 & n4004;
  assign n4006 = ~n4003 & ~n4005;
  assign n4007 = ~n3997 & ~n4006;
  assign n4008 = po41  & ~n4007;
  assign n4009 = ~n3708 & ~n3710;
  assign n4010 = n3717 & n4009;
  assign n4011 = po37  & n4010;
  assign n4012 = po37  & n4009;
  assign n4013 = ~n3717 & ~n4012;
  assign n4014 = ~n4011 & ~n4013;
  assign n4015 = ~po41  & n4007;
  assign n4016 = ~n4014 & ~n4015;
  assign n4017 = ~n4008 & ~n4016;
  assign n4018 = po42  & ~n4017;
  assign n4019 = ~n3720 & ~n3727;
  assign n4020 = n3726 & n4019;
  assign n4021 = po37  & n4020;
  assign n4022 = po37  & n4019;
  assign n4023 = ~n3726 & ~n4022;
  assign n4024 = ~n4021 & ~n4023;
  assign n4025 = ~po42  & ~n4008;
  assign n4026 = ~n4016 & n4025;
  assign n4027 = ~n4024 & ~n4026;
  assign n4028 = ~n4018 & ~n4027;
  assign n4029 = po43  & ~n4028;
  assign n4030 = ~n3730 & ~n3738;
  assign n4031 = n3736 & n4030;
  assign n4032 = po37  & n4031;
  assign n4033 = po37  & n4030;
  assign n4034 = ~n3736 & ~n4033;
  assign n4035 = ~n4032 & ~n4034;
  assign n4036 = ~po43  & n4028;
  assign n4037 = ~n4035 & ~n4036;
  assign n4038 = ~n4029 & ~n4037;
  assign n4039 = po44  & ~n4038;
  assign n4040 = ~n3741 & ~n3748;
  assign n4041 = n3747 & n4040;
  assign n4042 = po37  & n4041;
  assign n4043 = po37  & n4040;
  assign n4044 = ~n3747 & ~n4043;
  assign n4045 = ~n4042 & ~n4044;
  assign n4046 = ~po44  & ~n4029;
  assign n4047 = ~n4037 & n4046;
  assign n4048 = ~n4045 & ~n4047;
  assign n4049 = ~n4039 & ~n4048;
  assign n4050 = po45  & ~n4049;
  assign n4051 = ~n3751 & ~n3759;
  assign n4052 = n3757 & n4051;
  assign n4053 = po37  & n4052;
  assign n4054 = po37  & n4051;
  assign n4055 = ~n3757 & ~n4054;
  assign n4056 = ~n4053 & ~n4055;
  assign n4057 = ~po45  & n4049;
  assign n4058 = ~n4056 & ~n4057;
  assign n4059 = ~n4050 & ~n4058;
  assign n4060 = po46  & ~n4059;
  assign n4061 = ~n3762 & ~n3769;
  assign n4062 = n3768 & n4061;
  assign n4063 = po37  & n4062;
  assign n4064 = po37  & n4061;
  assign n4065 = ~n3768 & ~n4064;
  assign n4066 = ~n4063 & ~n4065;
  assign n4067 = ~po46  & ~n4050;
  assign n4068 = ~n4058 & n4067;
  assign n4069 = ~n4066 & ~n4068;
  assign n4070 = ~n4060 & ~n4069;
  assign n4071 = po47  & ~n4070;
  assign n4072 = ~n3772 & ~n3780;
  assign n4073 = n3778 & n4072;
  assign n4074 = po37  & n4073;
  assign n4075 = po37  & n4072;
  assign n4076 = ~n3778 & ~n4075;
  assign n4077 = ~n4074 & ~n4076;
  assign n4078 = ~po47  & n4070;
  assign n4079 = ~n4077 & ~n4078;
  assign n4080 = ~n4071 & ~n4079;
  assign n4081 = po48  & ~n4080;
  assign n4082 = ~n3783 & ~n3790;
  assign n4083 = n3789 & n4082;
  assign n4084 = po37  & n4083;
  assign n4085 = po37  & n4082;
  assign n4086 = ~n3789 & ~n4085;
  assign n4087 = ~n4084 & ~n4086;
  assign n4088 = ~po48  & ~n4071;
  assign n4089 = ~n4079 & n4088;
  assign n4090 = ~n4087 & ~n4089;
  assign n4091 = ~n4081 & ~n4090;
  assign n4092 = po49  & ~n4091;
  assign n4093 = ~n3793 & ~n3801;
  assign n4094 = n3799 & n4093;
  assign n4095 = po37  & n4094;
  assign n4096 = po37  & n4093;
  assign n4097 = ~n3799 & ~n4096;
  assign n4098 = ~n4095 & ~n4097;
  assign n4099 = ~po49  & n4091;
  assign n4100 = ~n4098 & ~n4099;
  assign n4101 = ~n4092 & ~n4100;
  assign n4102 = po50  & ~n4101;
  assign n4103 = ~n3804 & ~n3811;
  assign n4104 = n3810 & n4103;
  assign n4105 = po37  & n4104;
  assign n4106 = po37  & n4103;
  assign n4107 = ~n3810 & ~n4106;
  assign n4108 = ~n4105 & ~n4107;
  assign n4109 = ~po50  & ~n4092;
  assign n4110 = ~n4100 & n4109;
  assign n4111 = ~n4108 & ~n4110;
  assign n4112 = ~n4102 & ~n4111;
  assign n4113 = po51  & ~n4112;
  assign n4114 = ~n3814 & ~n3822;
  assign n4115 = n3820 & n4114;
  assign n4116 = po37  & n4115;
  assign n4117 = po37  & n4114;
  assign n4118 = ~n3820 & ~n4117;
  assign n4119 = ~n4116 & ~n4118;
  assign n4120 = ~po51  & n4112;
  assign n4121 = ~n4119 & ~n4120;
  assign n4122 = ~n4113 & ~n4121;
  assign n4123 = po52  & ~n4122;
  assign n4124 = ~n3825 & ~n3832;
  assign n4125 = n3831 & n4124;
  assign n4126 = po37  & n4125;
  assign n4127 = po37  & n4124;
  assign n4128 = ~n3831 & ~n4127;
  assign n4129 = ~n4126 & ~n4128;
  assign n4130 = ~po52  & ~n4113;
  assign n4131 = ~n4121 & n4130;
  assign n4132 = ~n4129 & ~n4131;
  assign n4133 = ~n4123 & ~n4132;
  assign n4134 = po53  & ~n4133;
  assign n4135 = ~n3835 & ~n3843;
  assign n4136 = n3841 & n4135;
  assign n4137 = po37  & n4136;
  assign n4138 = po37  & n4135;
  assign n4139 = ~n3841 & ~n4138;
  assign n4140 = ~n4137 & ~n4139;
  assign n4141 = ~po53  & n4133;
  assign n4142 = ~n4140 & ~n4141;
  assign n4143 = ~n4134 & ~n4142;
  assign n4144 = po54  & ~n4143;
  assign n4145 = ~n3846 & ~n3853;
  assign n4146 = n3852 & n4145;
  assign n4147 = po37  & n4146;
  assign n4148 = po37  & n4145;
  assign n4149 = ~n3852 & ~n4148;
  assign n4150 = ~n4147 & ~n4149;
  assign n4151 = ~po54  & ~n4134;
  assign n4152 = ~n4142 & n4151;
  assign n4153 = ~n4150 & ~n4152;
  assign n4154 = ~n4144 & ~n4153;
  assign n4155 = po55  & ~n4154;
  assign n4156 = ~n3856 & ~n3864;
  assign n4157 = n3862 & n4156;
  assign n4158 = po37  & n4157;
  assign n4159 = po37  & n4156;
  assign n4160 = ~n3862 & ~n4159;
  assign n4161 = ~n4158 & ~n4160;
  assign n4162 = ~po55  & n4154;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = ~n4155 & ~n4163;
  assign n4165 = po56  & ~n4164;
  assign n4166 = ~n3867 & ~n3874;
  assign n4167 = n3873 & n4166;
  assign n4168 = po37  & n4167;
  assign n4169 = po37  & n4166;
  assign n4170 = ~n3873 & ~n4169;
  assign n4171 = ~n4168 & ~n4170;
  assign n4172 = ~po56  & ~n4155;
  assign n4173 = ~n4163 & n4172;
  assign n4174 = ~n4171 & ~n4173;
  assign n4175 = ~n4165 & ~n4174;
  assign n4176 = po57  & ~n4175;
  assign n4177 = ~n3877 & ~n3885;
  assign n4178 = n3883 & n4177;
  assign n4179 = po37  & n4178;
  assign n4180 = po37  & n4177;
  assign n4181 = ~n3883 & ~n4180;
  assign n4182 = ~n4179 & ~n4181;
  assign n4183 = ~po57  & n4175;
  assign n4184 = ~n4182 & ~n4183;
  assign n4185 = ~n4176 & ~n4184;
  assign n4186 = po58  & ~n4185;
  assign n4187 = ~n3888 & ~n3895;
  assign n4188 = n3894 & n4187;
  assign n4189 = po37  & n4188;
  assign n4190 = po37  & n4187;
  assign n4191 = ~n3894 & ~n4190;
  assign n4192 = ~n4189 & ~n4191;
  assign n4193 = ~po58  & ~n4176;
  assign n4194 = ~n4184 & n4193;
  assign n4195 = ~n4192 & ~n4194;
  assign n4196 = ~n4186 & ~n4195;
  assign n4197 = po59  & ~n4196;
  assign n4198 = ~n3898 & ~n3906;
  assign n4199 = n3904 & n4198;
  assign n4200 = po37  & n4199;
  assign n4201 = po37  & n4198;
  assign n4202 = ~n3904 & ~n4201;
  assign n4203 = ~n4200 & ~n4202;
  assign n4204 = ~po59  & n4196;
  assign n4205 = ~n4203 & ~n4204;
  assign n4206 = ~n4197 & ~n4205;
  assign n4207 = po60  & ~n4206;
  assign n4208 = ~po60  & ~n4197;
  assign n4209 = ~n4205 & n4208;
  assign n4210 = ~n3909 & ~n3916;
  assign n4211 = n3915 & n4210;
  assign n4212 = po37  & n4211;
  assign n4213 = po37  & n4210;
  assign n4214 = ~n3915 & ~n4213;
  assign n4215 = ~n4212 & ~n4214;
  assign n4216 = ~n4209 & ~n4215;
  assign n4217 = ~n4207 & ~n4216;
  assign n4218 = po61  & ~n4217;
  assign n4219 = ~n3919 & ~n3927;
  assign n4220 = n3925 & n4219;
  assign n4221 = po37  & n4220;
  assign n4222 = po37  & n4219;
  assign n4223 = ~n3925 & ~n4222;
  assign n4224 = ~n4221 & ~n4223;
  assign n4225 = ~po61  & n4217;
  assign n4226 = ~n4224 & ~n4225;
  assign n4227 = ~n4218 & ~n4226;
  assign n4228 = po62  & ~n4227;
  assign n4229 = ~n3930 & ~n3937;
  assign n4230 = n3936 & n4229;
  assign n4231 = po37  & n4230;
  assign n4232 = po37  & n4229;
  assign n4233 = ~n3936 & ~n4232;
  assign n4234 = ~n4231 & ~n4233;
  assign n4235 = ~po62  & ~n4218;
  assign n4236 = ~n4226 & n4235;
  assign n4237 = ~n4234 & ~n4236;
  assign n4238 = ~n4228 & ~n4237;
  assign n4239 = ~n3940 & ~n3948;
  assign n4240 = po37  & n4239;
  assign n4241 = ~n3946 & ~n4240;
  assign n4242 = n3946 & n4240;
  assign n4243 = ~n4241 & ~n4242;
  assign n4244 = ~n3950 & ~n3955;
  assign n4245 = po37  & n4244;
  assign n4246 = ~n3968 & ~n4245;
  assign n4247 = ~n4243 & n4246;
  assign n4248 = ~n4238 & n4247;
  assign n4249 = ~po63  & ~n4248;
  assign n4250 = ~n3955 & po37 ;
  assign n4251 = n3950 & ~n4250;
  assign n4252 = po63  & ~n4244;
  assign n4253 = ~n4251 & n4252;
  assign n4254 = n3955 & ~po37 ;
  assign n4255 = ~n4253 & ~n4254;
  assign n4256 = n4238 & n4243;
  assign n4257 = n4255 & ~n4256;
  assign po36  = n4249 | ~n4257;
  assign n4259 = pi72  & po36 ;
  assign n4260 = ~pi70  & ~pi71 ;
  assign n4261 = ~pi72  & n4260;
  assign n4262 = ~n4259 & ~n4261;
  assign n4263 = po37  & ~n4262;
  assign n4264 = n3967 & ~n4261;
  assign n4265 = ~n3968 & n4264;
  assign n4266 = ~n3961 & n4265;
  assign n4267 = ~n4259 & n4266;
  assign n4268 = ~pi72  & po36 ;
  assign n4269 = pi73  & ~n4268;
  assign n4270 = n3972 & po36 ;
  assign n4271 = ~n4269 & ~n4270;
  assign n4272 = ~n4267 & n4271;
  assign n4273 = ~n4263 & ~n4272;
  assign n4274 = po38  & ~n4273;
  assign n4275 = ~po38  & ~n4263;
  assign n4276 = ~n4272 & n4275;
  assign n4277 = po37  & n4255;
  assign n4278 = ~n4256 & n4277;
  assign n4279 = ~n4249 & n4278;
  assign n4280 = ~n4270 & ~n4279;
  assign n4281 = pi74  & ~n4280;
  assign n4282 = ~pi74  & n4280;
  assign n4283 = ~n4281 & ~n4282;
  assign n4284 = ~n4276 & ~n4283;
  assign n4285 = ~n4274 & ~n4284;
  assign n4286 = po39  & ~n4285;
  assign n4287 = ~n3975 & ~n3979;
  assign n4288 = ~n3983 & n4287;
  assign n4289 = po36  & n4288;
  assign n4290 = po36  & n4287;
  assign n4291 = n3983 & ~n4290;
  assign n4292 = ~n4289 & ~n4291;
  assign n4293 = ~po39  & n4285;
  assign n4294 = ~n4292 & ~n4293;
  assign n4295 = ~n4286 & ~n4294;
  assign n4296 = po40  & ~n4295;
  assign n4297 = ~n3986 & ~n3994;
  assign n4298 = n3993 & n4297;
  assign n4299 = po36  & n4298;
  assign n4300 = po36  & n4297;
  assign n4301 = ~n3993 & ~n4300;
  assign n4302 = ~n4299 & ~n4301;
  assign n4303 = ~po40  & ~n4286;
  assign n4304 = ~n4294 & n4303;
  assign n4305 = ~n4302 & ~n4304;
  assign n4306 = ~n4296 & ~n4305;
  assign n4307 = po41  & ~n4306;
  assign n4308 = ~n3997 & ~n4005;
  assign n4309 = n4003 & n4308;
  assign n4310 = po36  & n4309;
  assign n4311 = po36  & n4308;
  assign n4312 = ~n4003 & ~n4311;
  assign n4313 = ~n4310 & ~n4312;
  assign n4314 = ~po41  & n4306;
  assign n4315 = ~n4313 & ~n4314;
  assign n4316 = ~n4307 & ~n4315;
  assign n4317 = po42  & ~n4316;
  assign n4318 = ~n4008 & ~n4015;
  assign n4319 = n4014 & n4318;
  assign n4320 = po36  & n4319;
  assign n4321 = po36  & n4318;
  assign n4322 = ~n4014 & ~n4321;
  assign n4323 = ~n4320 & ~n4322;
  assign n4324 = ~po42  & ~n4307;
  assign n4325 = ~n4315 & n4324;
  assign n4326 = ~n4323 & ~n4325;
  assign n4327 = ~n4317 & ~n4326;
  assign n4328 = po43  & ~n4327;
  assign n4329 = ~n4018 & ~n4026;
  assign n4330 = n4024 & n4329;
  assign n4331 = po36  & n4330;
  assign n4332 = po36  & n4329;
  assign n4333 = ~n4024 & ~n4332;
  assign n4334 = ~n4331 & ~n4333;
  assign n4335 = ~po43  & n4327;
  assign n4336 = ~n4334 & ~n4335;
  assign n4337 = ~n4328 & ~n4336;
  assign n4338 = po44  & ~n4337;
  assign n4339 = ~n4029 & ~n4036;
  assign n4340 = n4035 & n4339;
  assign n4341 = po36  & n4340;
  assign n4342 = po36  & n4339;
  assign n4343 = ~n4035 & ~n4342;
  assign n4344 = ~n4341 & ~n4343;
  assign n4345 = ~po44  & ~n4328;
  assign n4346 = ~n4336 & n4345;
  assign n4347 = ~n4344 & ~n4346;
  assign n4348 = ~n4338 & ~n4347;
  assign n4349 = po45  & ~n4348;
  assign n4350 = ~n4039 & ~n4047;
  assign n4351 = n4045 & n4350;
  assign n4352 = po36  & n4351;
  assign n4353 = po36  & n4350;
  assign n4354 = ~n4045 & ~n4353;
  assign n4355 = ~n4352 & ~n4354;
  assign n4356 = ~po45  & n4348;
  assign n4357 = ~n4355 & ~n4356;
  assign n4358 = ~n4349 & ~n4357;
  assign n4359 = po46  & ~n4358;
  assign n4360 = ~n4050 & ~n4057;
  assign n4361 = n4056 & n4360;
  assign n4362 = po36  & n4361;
  assign n4363 = po36  & n4360;
  assign n4364 = ~n4056 & ~n4363;
  assign n4365 = ~n4362 & ~n4364;
  assign n4366 = ~po46  & ~n4349;
  assign n4367 = ~n4357 & n4366;
  assign n4368 = ~n4365 & ~n4367;
  assign n4369 = ~n4359 & ~n4368;
  assign n4370 = po47  & ~n4369;
  assign n4371 = ~n4060 & ~n4068;
  assign n4372 = n4066 & n4371;
  assign n4373 = po36  & n4372;
  assign n4374 = po36  & n4371;
  assign n4375 = ~n4066 & ~n4374;
  assign n4376 = ~n4373 & ~n4375;
  assign n4377 = ~po47  & n4369;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = ~n4370 & ~n4378;
  assign n4380 = po48  & ~n4379;
  assign n4381 = ~n4071 & ~n4078;
  assign n4382 = n4077 & n4381;
  assign n4383 = po36  & n4382;
  assign n4384 = po36  & n4381;
  assign n4385 = ~n4077 & ~n4384;
  assign n4386 = ~n4383 & ~n4385;
  assign n4387 = ~po48  & ~n4370;
  assign n4388 = ~n4378 & n4387;
  assign n4389 = ~n4386 & ~n4388;
  assign n4390 = ~n4380 & ~n4389;
  assign n4391 = po49  & ~n4390;
  assign n4392 = ~n4081 & ~n4089;
  assign n4393 = n4087 & n4392;
  assign n4394 = po36  & n4393;
  assign n4395 = po36  & n4392;
  assign n4396 = ~n4087 & ~n4395;
  assign n4397 = ~n4394 & ~n4396;
  assign n4398 = ~po49  & n4390;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = ~n4391 & ~n4399;
  assign n4401 = po50  & ~n4400;
  assign n4402 = ~n4092 & ~n4099;
  assign n4403 = n4098 & n4402;
  assign n4404 = po36  & n4403;
  assign n4405 = po36  & n4402;
  assign n4406 = ~n4098 & ~n4405;
  assign n4407 = ~n4404 & ~n4406;
  assign n4408 = ~po50  & ~n4391;
  assign n4409 = ~n4399 & n4408;
  assign n4410 = ~n4407 & ~n4409;
  assign n4411 = ~n4401 & ~n4410;
  assign n4412 = po51  & ~n4411;
  assign n4413 = ~n4102 & ~n4110;
  assign n4414 = n4108 & n4413;
  assign n4415 = po36  & n4414;
  assign n4416 = po36  & n4413;
  assign n4417 = ~n4108 & ~n4416;
  assign n4418 = ~n4415 & ~n4417;
  assign n4419 = ~po51  & n4411;
  assign n4420 = ~n4418 & ~n4419;
  assign n4421 = ~n4412 & ~n4420;
  assign n4422 = po52  & ~n4421;
  assign n4423 = ~n4113 & ~n4120;
  assign n4424 = n4119 & n4423;
  assign n4425 = po36  & n4424;
  assign n4426 = po36  & n4423;
  assign n4427 = ~n4119 & ~n4426;
  assign n4428 = ~n4425 & ~n4427;
  assign n4429 = ~po52  & ~n4412;
  assign n4430 = ~n4420 & n4429;
  assign n4431 = ~n4428 & ~n4430;
  assign n4432 = ~n4422 & ~n4431;
  assign n4433 = po53  & ~n4432;
  assign n4434 = ~n4123 & ~n4131;
  assign n4435 = n4129 & n4434;
  assign n4436 = po36  & n4435;
  assign n4437 = po36  & n4434;
  assign n4438 = ~n4129 & ~n4437;
  assign n4439 = ~n4436 & ~n4438;
  assign n4440 = ~po53  & n4432;
  assign n4441 = ~n4439 & ~n4440;
  assign n4442 = ~n4433 & ~n4441;
  assign n4443 = po54  & ~n4442;
  assign n4444 = ~n4134 & ~n4141;
  assign n4445 = n4140 & n4444;
  assign n4446 = po36  & n4445;
  assign n4447 = po36  & n4444;
  assign n4448 = ~n4140 & ~n4447;
  assign n4449 = ~n4446 & ~n4448;
  assign n4450 = ~po54  & ~n4433;
  assign n4451 = ~n4441 & n4450;
  assign n4452 = ~n4449 & ~n4451;
  assign n4453 = ~n4443 & ~n4452;
  assign n4454 = po55  & ~n4453;
  assign n4455 = ~n4144 & ~n4152;
  assign n4456 = n4150 & n4455;
  assign n4457 = po36  & n4456;
  assign n4458 = po36  & n4455;
  assign n4459 = ~n4150 & ~n4458;
  assign n4460 = ~n4457 & ~n4459;
  assign n4461 = ~po55  & n4453;
  assign n4462 = ~n4460 & ~n4461;
  assign n4463 = ~n4454 & ~n4462;
  assign n4464 = po56  & ~n4463;
  assign n4465 = ~n4155 & ~n4162;
  assign n4466 = n4161 & n4465;
  assign n4467 = po36  & n4466;
  assign n4468 = po36  & n4465;
  assign n4469 = ~n4161 & ~n4468;
  assign n4470 = ~n4467 & ~n4469;
  assign n4471 = ~po56  & ~n4454;
  assign n4472 = ~n4462 & n4471;
  assign n4473 = ~n4470 & ~n4472;
  assign n4474 = ~n4464 & ~n4473;
  assign n4475 = po57  & ~n4474;
  assign n4476 = ~n4165 & ~n4173;
  assign n4477 = n4171 & n4476;
  assign n4478 = po36  & n4477;
  assign n4479 = po36  & n4476;
  assign n4480 = ~n4171 & ~n4479;
  assign n4481 = ~n4478 & ~n4480;
  assign n4482 = ~po57  & n4474;
  assign n4483 = ~n4481 & ~n4482;
  assign n4484 = ~n4475 & ~n4483;
  assign n4485 = po58  & ~n4484;
  assign n4486 = ~n4176 & ~n4183;
  assign n4487 = n4182 & n4486;
  assign n4488 = po36  & n4487;
  assign n4489 = po36  & n4486;
  assign n4490 = ~n4182 & ~n4489;
  assign n4491 = ~n4488 & ~n4490;
  assign n4492 = ~po58  & ~n4475;
  assign n4493 = ~n4483 & n4492;
  assign n4494 = ~n4491 & ~n4493;
  assign n4495 = ~n4485 & ~n4494;
  assign n4496 = po59  & ~n4495;
  assign n4497 = ~n4186 & ~n4194;
  assign n4498 = n4192 & n4497;
  assign n4499 = po36  & n4498;
  assign n4500 = po36  & n4497;
  assign n4501 = ~n4192 & ~n4500;
  assign n4502 = ~n4499 & ~n4501;
  assign n4503 = ~po59  & n4495;
  assign n4504 = ~n4502 & ~n4503;
  assign n4505 = ~n4496 & ~n4504;
  assign n4506 = po60  & ~n4505;
  assign n4507 = ~n4197 & ~n4204;
  assign n4508 = n4203 & n4507;
  assign n4509 = po36  & n4508;
  assign n4510 = po36  & n4507;
  assign n4511 = ~n4203 & ~n4510;
  assign n4512 = ~n4509 & ~n4511;
  assign n4513 = ~po60  & ~n4496;
  assign n4514 = ~n4504 & n4513;
  assign n4515 = ~n4512 & ~n4514;
  assign n4516 = ~n4506 & ~n4515;
  assign n4517 = po61  & ~n4516;
  assign n4518 = ~n4207 & ~n4209;
  assign n4519 = n4215 & n4518;
  assign n4520 = po36  & n4519;
  assign n4521 = po36  & n4518;
  assign n4522 = ~n4215 & ~n4521;
  assign n4523 = ~n4520 & ~n4522;
  assign n4524 = ~po61  & n4516;
  assign n4525 = ~n4523 & ~n4524;
  assign n4526 = ~n4517 & ~n4525;
  assign n4527 = po62  & ~n4526;
  assign n4528 = ~n4218 & ~n4225;
  assign n4529 = n4224 & n4528;
  assign n4530 = po36  & n4529;
  assign n4531 = po36  & n4528;
  assign n4532 = ~n4224 & ~n4531;
  assign n4533 = ~n4530 & ~n4532;
  assign n4534 = ~po62  & ~n4517;
  assign n4535 = ~n4525 & n4534;
  assign n4536 = ~n4533 & ~n4535;
  assign n4537 = ~n4527 & ~n4536;
  assign n4538 = ~n4228 & ~n4236;
  assign n4539 = po36  & n4538;
  assign n4540 = ~n4234 & ~n4539;
  assign n4541 = n4234 & n4539;
  assign n4542 = ~n4540 & ~n4541;
  assign n4543 = ~n4238 & ~n4243;
  assign n4544 = po36  & n4543;
  assign n4545 = ~n4256 & ~n4544;
  assign n4546 = ~n4542 & n4545;
  assign n4547 = ~n4537 & n4546;
  assign n4548 = ~po63  & ~n4547;
  assign n4549 = ~n4243 & po36 ;
  assign n4550 = n4238 & ~n4549;
  assign n4551 = po63  & ~n4543;
  assign n4552 = ~n4550 & n4551;
  assign n4553 = n4243 & ~po36 ;
  assign n4554 = ~n4552 & ~n4553;
  assign n4555 = n4537 & n4542;
  assign n4556 = n4554 & ~n4555;
  assign po35  = n4548 | ~n4556;
  assign n4558 = pi70  & po35 ;
  assign n4559 = ~pi68  & ~pi69 ;
  assign n4560 = ~pi70  & n4559;
  assign n4561 = ~n4558 & ~n4560;
  assign n4562 = po36  & ~n4561;
  assign n4563 = n4255 & ~n4560;
  assign n4564 = ~n4256 & n4563;
  assign n4565 = ~n4249 & n4564;
  assign n4566 = ~n4558 & n4565;
  assign n4567 = ~pi70  & po35 ;
  assign n4568 = pi71  & ~n4567;
  assign n4569 = n4260 & po35 ;
  assign n4570 = ~n4568 & ~n4569;
  assign n4571 = ~n4566 & n4570;
  assign n4572 = ~n4562 & ~n4571;
  assign n4573 = po37  & ~n4572;
  assign n4574 = po36  & n4554;
  assign n4575 = ~n4555 & n4574;
  assign n4576 = ~n4548 & n4575;
  assign n4577 = ~n4569 & ~n4576;
  assign n4578 = pi72  & ~n4577;
  assign n4579 = ~pi72  & n4577;
  assign n4580 = ~n4578 & ~n4579;
  assign n4581 = ~po37  & n4572;
  assign n4582 = ~n4580 & ~n4581;
  assign n4583 = ~n4573 & ~n4582;
  assign n4584 = po38  & ~n4583;
  assign n4585 = ~n4263 & ~n4267;
  assign n4586 = ~n4271 & n4585;
  assign n4587 = po35  & n4586;
  assign n4588 = po35  & n4585;
  assign n4589 = n4271 & ~n4588;
  assign n4590 = ~n4587 & ~n4589;
  assign n4591 = ~po38  & ~n4573;
  assign n4592 = ~n4582 & n4591;
  assign n4593 = ~n4590 & ~n4592;
  assign n4594 = ~n4584 & ~n4593;
  assign n4595 = po39  & ~n4594;
  assign n4596 = ~n4274 & ~n4276;
  assign n4597 = n4283 & n4596;
  assign n4598 = po35  & n4597;
  assign n4599 = po35  & n4596;
  assign n4600 = ~n4283 & ~n4599;
  assign n4601 = ~n4598 & ~n4600;
  assign n4602 = ~po39  & n4594;
  assign n4603 = ~n4601 & ~n4602;
  assign n4604 = ~n4595 & ~n4603;
  assign n4605 = po40  & ~n4604;
  assign n4606 = ~n4286 & ~n4293;
  assign n4607 = n4292 & n4606;
  assign n4608 = po35  & n4607;
  assign n4609 = po35  & n4606;
  assign n4610 = ~n4292 & ~n4609;
  assign n4611 = ~n4608 & ~n4610;
  assign n4612 = ~po40  & ~n4595;
  assign n4613 = ~n4603 & n4612;
  assign n4614 = ~n4611 & ~n4613;
  assign n4615 = ~n4605 & ~n4614;
  assign n4616 = po41  & ~n4615;
  assign n4617 = ~n4296 & ~n4304;
  assign n4618 = n4302 & n4617;
  assign n4619 = po35  & n4618;
  assign n4620 = po35  & n4617;
  assign n4621 = ~n4302 & ~n4620;
  assign n4622 = ~n4619 & ~n4621;
  assign n4623 = ~po41  & n4615;
  assign n4624 = ~n4622 & ~n4623;
  assign n4625 = ~n4616 & ~n4624;
  assign n4626 = po42  & ~n4625;
  assign n4627 = ~n4307 & ~n4314;
  assign n4628 = n4313 & n4627;
  assign n4629 = po35  & n4628;
  assign n4630 = po35  & n4627;
  assign n4631 = ~n4313 & ~n4630;
  assign n4632 = ~n4629 & ~n4631;
  assign n4633 = ~po42  & ~n4616;
  assign n4634 = ~n4624 & n4633;
  assign n4635 = ~n4632 & ~n4634;
  assign n4636 = ~n4626 & ~n4635;
  assign n4637 = po43  & ~n4636;
  assign n4638 = ~n4317 & ~n4325;
  assign n4639 = n4323 & n4638;
  assign n4640 = po35  & n4639;
  assign n4641 = po35  & n4638;
  assign n4642 = ~n4323 & ~n4641;
  assign n4643 = ~n4640 & ~n4642;
  assign n4644 = ~po43  & n4636;
  assign n4645 = ~n4643 & ~n4644;
  assign n4646 = ~n4637 & ~n4645;
  assign n4647 = po44  & ~n4646;
  assign n4648 = ~n4328 & ~n4335;
  assign n4649 = n4334 & n4648;
  assign n4650 = po35  & n4649;
  assign n4651 = po35  & n4648;
  assign n4652 = ~n4334 & ~n4651;
  assign n4653 = ~n4650 & ~n4652;
  assign n4654 = ~po44  & ~n4637;
  assign n4655 = ~n4645 & n4654;
  assign n4656 = ~n4653 & ~n4655;
  assign n4657 = ~n4647 & ~n4656;
  assign n4658 = po45  & ~n4657;
  assign n4659 = ~n4338 & ~n4346;
  assign n4660 = n4344 & n4659;
  assign n4661 = po35  & n4660;
  assign n4662 = po35  & n4659;
  assign n4663 = ~n4344 & ~n4662;
  assign n4664 = ~n4661 & ~n4663;
  assign n4665 = ~po45  & n4657;
  assign n4666 = ~n4664 & ~n4665;
  assign n4667 = ~n4658 & ~n4666;
  assign n4668 = po46  & ~n4667;
  assign n4669 = ~n4349 & ~n4356;
  assign n4670 = n4355 & n4669;
  assign n4671 = po35  & n4670;
  assign n4672 = po35  & n4669;
  assign n4673 = ~n4355 & ~n4672;
  assign n4674 = ~n4671 & ~n4673;
  assign n4675 = ~po46  & ~n4658;
  assign n4676 = ~n4666 & n4675;
  assign n4677 = ~n4674 & ~n4676;
  assign n4678 = ~n4668 & ~n4677;
  assign n4679 = po47  & ~n4678;
  assign n4680 = ~n4359 & ~n4367;
  assign n4681 = n4365 & n4680;
  assign n4682 = po35  & n4681;
  assign n4683 = po35  & n4680;
  assign n4684 = ~n4365 & ~n4683;
  assign n4685 = ~n4682 & ~n4684;
  assign n4686 = ~po47  & n4678;
  assign n4687 = ~n4685 & ~n4686;
  assign n4688 = ~n4679 & ~n4687;
  assign n4689 = po48  & ~n4688;
  assign n4690 = ~n4370 & ~n4377;
  assign n4691 = n4376 & n4690;
  assign n4692 = po35  & n4691;
  assign n4693 = po35  & n4690;
  assign n4694 = ~n4376 & ~n4693;
  assign n4695 = ~n4692 & ~n4694;
  assign n4696 = ~po48  & ~n4679;
  assign n4697 = ~n4687 & n4696;
  assign n4698 = ~n4695 & ~n4697;
  assign n4699 = ~n4689 & ~n4698;
  assign n4700 = po49  & ~n4699;
  assign n4701 = ~n4380 & ~n4388;
  assign n4702 = n4386 & n4701;
  assign n4703 = po35  & n4702;
  assign n4704 = po35  & n4701;
  assign n4705 = ~n4386 & ~n4704;
  assign n4706 = ~n4703 & ~n4705;
  assign n4707 = ~po49  & n4699;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = ~n4700 & ~n4708;
  assign n4710 = po50  & ~n4709;
  assign n4711 = ~n4391 & ~n4398;
  assign n4712 = n4397 & n4711;
  assign n4713 = po35  & n4712;
  assign n4714 = po35  & n4711;
  assign n4715 = ~n4397 & ~n4714;
  assign n4716 = ~n4713 & ~n4715;
  assign n4717 = ~po50  & ~n4700;
  assign n4718 = ~n4708 & n4717;
  assign n4719 = ~n4716 & ~n4718;
  assign n4720 = ~n4710 & ~n4719;
  assign n4721 = po51  & ~n4720;
  assign n4722 = ~n4401 & ~n4409;
  assign n4723 = n4407 & n4722;
  assign n4724 = po35  & n4723;
  assign n4725 = po35  & n4722;
  assign n4726 = ~n4407 & ~n4725;
  assign n4727 = ~n4724 & ~n4726;
  assign n4728 = ~po51  & n4720;
  assign n4729 = ~n4727 & ~n4728;
  assign n4730 = ~n4721 & ~n4729;
  assign n4731 = po52  & ~n4730;
  assign n4732 = ~n4412 & ~n4419;
  assign n4733 = n4418 & n4732;
  assign n4734 = po35  & n4733;
  assign n4735 = po35  & n4732;
  assign n4736 = ~n4418 & ~n4735;
  assign n4737 = ~n4734 & ~n4736;
  assign n4738 = ~po52  & ~n4721;
  assign n4739 = ~n4729 & n4738;
  assign n4740 = ~n4737 & ~n4739;
  assign n4741 = ~n4731 & ~n4740;
  assign n4742 = po53  & ~n4741;
  assign n4743 = ~n4422 & ~n4430;
  assign n4744 = n4428 & n4743;
  assign n4745 = po35  & n4744;
  assign n4746 = po35  & n4743;
  assign n4747 = ~n4428 & ~n4746;
  assign n4748 = ~n4745 & ~n4747;
  assign n4749 = ~po53  & n4741;
  assign n4750 = ~n4748 & ~n4749;
  assign n4751 = ~n4742 & ~n4750;
  assign n4752 = po54  & ~n4751;
  assign n4753 = ~n4433 & ~n4440;
  assign n4754 = n4439 & n4753;
  assign n4755 = po35  & n4754;
  assign n4756 = po35  & n4753;
  assign n4757 = ~n4439 & ~n4756;
  assign n4758 = ~n4755 & ~n4757;
  assign n4759 = ~po54  & ~n4742;
  assign n4760 = ~n4750 & n4759;
  assign n4761 = ~n4758 & ~n4760;
  assign n4762 = ~n4752 & ~n4761;
  assign n4763 = po55  & ~n4762;
  assign n4764 = ~n4443 & ~n4451;
  assign n4765 = n4449 & n4764;
  assign n4766 = po35  & n4765;
  assign n4767 = po35  & n4764;
  assign n4768 = ~n4449 & ~n4767;
  assign n4769 = ~n4766 & ~n4768;
  assign n4770 = ~po55  & n4762;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = ~n4763 & ~n4771;
  assign n4773 = po56  & ~n4772;
  assign n4774 = ~n4454 & ~n4461;
  assign n4775 = n4460 & n4774;
  assign n4776 = po35  & n4775;
  assign n4777 = po35  & n4774;
  assign n4778 = ~n4460 & ~n4777;
  assign n4779 = ~n4776 & ~n4778;
  assign n4780 = ~po56  & ~n4763;
  assign n4781 = ~n4771 & n4780;
  assign n4782 = ~n4779 & ~n4781;
  assign n4783 = ~n4773 & ~n4782;
  assign n4784 = po57  & ~n4783;
  assign n4785 = ~n4464 & ~n4472;
  assign n4786 = n4470 & n4785;
  assign n4787 = po35  & n4786;
  assign n4788 = po35  & n4785;
  assign n4789 = ~n4470 & ~n4788;
  assign n4790 = ~n4787 & ~n4789;
  assign n4791 = ~po57  & n4783;
  assign n4792 = ~n4790 & ~n4791;
  assign n4793 = ~n4784 & ~n4792;
  assign n4794 = po58  & ~n4793;
  assign n4795 = ~n4475 & ~n4482;
  assign n4796 = n4481 & n4795;
  assign n4797 = po35  & n4796;
  assign n4798 = po35  & n4795;
  assign n4799 = ~n4481 & ~n4798;
  assign n4800 = ~n4797 & ~n4799;
  assign n4801 = ~po58  & ~n4784;
  assign n4802 = ~n4792 & n4801;
  assign n4803 = ~n4800 & ~n4802;
  assign n4804 = ~n4794 & ~n4803;
  assign n4805 = po59  & ~n4804;
  assign n4806 = ~n4485 & ~n4493;
  assign n4807 = n4491 & n4806;
  assign n4808 = po35  & n4807;
  assign n4809 = po35  & n4806;
  assign n4810 = ~n4491 & ~n4809;
  assign n4811 = ~n4808 & ~n4810;
  assign n4812 = ~po59  & n4804;
  assign n4813 = ~n4811 & ~n4812;
  assign n4814 = ~n4805 & ~n4813;
  assign n4815 = po60  & ~n4814;
  assign n4816 = ~n4496 & ~n4503;
  assign n4817 = n4502 & n4816;
  assign n4818 = po35  & n4817;
  assign n4819 = po35  & n4816;
  assign n4820 = ~n4502 & ~n4819;
  assign n4821 = ~n4818 & ~n4820;
  assign n4822 = ~po60  & ~n4805;
  assign n4823 = ~n4813 & n4822;
  assign n4824 = ~n4821 & ~n4823;
  assign n4825 = ~n4815 & ~n4824;
  assign n4826 = po61  & ~n4825;
  assign n4827 = ~n4506 & ~n4514;
  assign n4828 = n4512 & n4827;
  assign n4829 = po35  & n4828;
  assign n4830 = po35  & n4827;
  assign n4831 = ~n4512 & ~n4830;
  assign n4832 = ~n4829 & ~n4831;
  assign n4833 = ~po61  & n4825;
  assign n4834 = ~n4832 & ~n4833;
  assign n4835 = ~n4826 & ~n4834;
  assign n4836 = po62  & ~n4835;
  assign n4837 = ~po62  & ~n4826;
  assign n4838 = ~n4834 & n4837;
  assign n4839 = ~n4517 & ~n4524;
  assign n4840 = n4523 & n4839;
  assign n4841 = po35  & n4840;
  assign n4842 = po35  & n4839;
  assign n4843 = ~n4523 & ~n4842;
  assign n4844 = ~n4841 & ~n4843;
  assign n4845 = ~n4838 & ~n4844;
  assign n4846 = ~n4836 & ~n4845;
  assign n4847 = ~n4527 & ~n4535;
  assign n4848 = po35  & n4847;
  assign n4849 = ~n4533 & ~n4848;
  assign n4850 = n4533 & n4848;
  assign n4851 = ~n4849 & ~n4850;
  assign n4852 = ~n4537 & ~n4542;
  assign n4853 = po35  & n4852;
  assign n4854 = ~n4555 & ~n4853;
  assign n4855 = ~n4851 & n4854;
  assign n4856 = ~n4846 & n4855;
  assign n4857 = ~po63  & ~n4856;
  assign n4858 = ~n4542 & po35 ;
  assign n4859 = n4537 & ~n4858;
  assign n4860 = po63  & ~n4852;
  assign n4861 = ~n4859 & n4860;
  assign n4862 = n4542 & ~po35 ;
  assign n4863 = ~n4861 & ~n4862;
  assign n4864 = n4846 & n4851;
  assign n4865 = n4863 & ~n4864;
  assign po34  = n4857 | ~n4865;
  assign n4867 = pi68  & po34 ;
  assign n4868 = ~pi66  & ~pi67 ;
  assign n4869 = ~pi68  & n4868;
  assign n4870 = ~n4867 & ~n4869;
  assign n4871 = po35  & ~n4870;
  assign n4872 = n4554 & ~n4869;
  assign n4873 = ~n4555 & n4872;
  assign n4874 = ~n4548 & n4873;
  assign n4875 = ~n4867 & n4874;
  assign n4876 = ~pi68  & po34 ;
  assign n4877 = pi69  & ~n4876;
  assign n4878 = n4559 & po34 ;
  assign n4879 = ~n4877 & ~n4878;
  assign n4880 = ~n4875 & n4879;
  assign n4881 = ~n4871 & ~n4880;
  assign n4882 = po36  & ~n4881;
  assign n4883 = ~po36  & ~n4871;
  assign n4884 = ~n4880 & n4883;
  assign n4885 = po35  & n4863;
  assign n4886 = ~n4864 & n4885;
  assign n4887 = ~n4857 & n4886;
  assign n4888 = ~n4878 & ~n4887;
  assign n4889 = pi70  & ~n4888;
  assign n4890 = ~pi70  & n4888;
  assign n4891 = ~n4889 & ~n4890;
  assign n4892 = ~n4884 & ~n4891;
  assign n4893 = ~n4882 & ~n4892;
  assign n4894 = po37  & ~n4893;
  assign n4895 = ~n4562 & ~n4566;
  assign n4896 = ~n4570 & n4895;
  assign n4897 = po34  & n4896;
  assign n4898 = po34  & n4895;
  assign n4899 = n4570 & ~n4898;
  assign n4900 = ~n4897 & ~n4899;
  assign n4901 = ~po37  & n4893;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = ~n4894 & ~n4902;
  assign n4904 = po38  & ~n4903;
  assign n4905 = ~n4573 & ~n4581;
  assign n4906 = n4580 & n4905;
  assign n4907 = po34  & n4906;
  assign n4908 = po34  & n4905;
  assign n4909 = ~n4580 & ~n4908;
  assign n4910 = ~n4907 & ~n4909;
  assign n4911 = ~po38  & ~n4894;
  assign n4912 = ~n4902 & n4911;
  assign n4913 = ~n4910 & ~n4912;
  assign n4914 = ~n4904 & ~n4913;
  assign n4915 = po39  & ~n4914;
  assign n4916 = ~n4584 & ~n4592;
  assign n4917 = n4590 & n4916;
  assign n4918 = po34  & n4917;
  assign n4919 = po34  & n4916;
  assign n4920 = ~n4590 & ~n4919;
  assign n4921 = ~n4918 & ~n4920;
  assign n4922 = ~po39  & n4914;
  assign n4923 = ~n4921 & ~n4922;
  assign n4924 = ~n4915 & ~n4923;
  assign n4925 = po40  & ~n4924;
  assign n4926 = ~n4595 & ~n4602;
  assign n4927 = n4601 & n4926;
  assign n4928 = po34  & n4927;
  assign n4929 = po34  & n4926;
  assign n4930 = ~n4601 & ~n4929;
  assign n4931 = ~n4928 & ~n4930;
  assign n4932 = ~po40  & ~n4915;
  assign n4933 = ~n4923 & n4932;
  assign n4934 = ~n4931 & ~n4933;
  assign n4935 = ~n4925 & ~n4934;
  assign n4936 = po41  & ~n4935;
  assign n4937 = ~n4605 & ~n4613;
  assign n4938 = n4611 & n4937;
  assign n4939 = po34  & n4938;
  assign n4940 = po34  & n4937;
  assign n4941 = ~n4611 & ~n4940;
  assign n4942 = ~n4939 & ~n4941;
  assign n4943 = ~po41  & n4935;
  assign n4944 = ~n4942 & ~n4943;
  assign n4945 = ~n4936 & ~n4944;
  assign n4946 = po42  & ~n4945;
  assign n4947 = ~n4616 & ~n4623;
  assign n4948 = n4622 & n4947;
  assign n4949 = po34  & n4948;
  assign n4950 = po34  & n4947;
  assign n4951 = ~n4622 & ~n4950;
  assign n4952 = ~n4949 & ~n4951;
  assign n4953 = ~po42  & ~n4936;
  assign n4954 = ~n4944 & n4953;
  assign n4955 = ~n4952 & ~n4954;
  assign n4956 = ~n4946 & ~n4955;
  assign n4957 = po43  & ~n4956;
  assign n4958 = ~n4626 & ~n4634;
  assign n4959 = n4632 & n4958;
  assign n4960 = po34  & n4959;
  assign n4961 = po34  & n4958;
  assign n4962 = ~n4632 & ~n4961;
  assign n4963 = ~n4960 & ~n4962;
  assign n4964 = ~po43  & n4956;
  assign n4965 = ~n4963 & ~n4964;
  assign n4966 = ~n4957 & ~n4965;
  assign n4967 = po44  & ~n4966;
  assign n4968 = ~n4637 & ~n4644;
  assign n4969 = n4643 & n4968;
  assign n4970 = po34  & n4969;
  assign n4971 = po34  & n4968;
  assign n4972 = ~n4643 & ~n4971;
  assign n4973 = ~n4970 & ~n4972;
  assign n4974 = ~po44  & ~n4957;
  assign n4975 = ~n4965 & n4974;
  assign n4976 = ~n4973 & ~n4975;
  assign n4977 = ~n4967 & ~n4976;
  assign n4978 = po45  & ~n4977;
  assign n4979 = ~n4647 & ~n4655;
  assign n4980 = n4653 & n4979;
  assign n4981 = po34  & n4980;
  assign n4982 = po34  & n4979;
  assign n4983 = ~n4653 & ~n4982;
  assign n4984 = ~n4981 & ~n4983;
  assign n4985 = ~po45  & n4977;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = ~n4978 & ~n4986;
  assign n4988 = po46  & ~n4987;
  assign n4989 = ~n4658 & ~n4665;
  assign n4990 = n4664 & n4989;
  assign n4991 = po34  & n4990;
  assign n4992 = po34  & n4989;
  assign n4993 = ~n4664 & ~n4992;
  assign n4994 = ~n4991 & ~n4993;
  assign n4995 = ~po46  & ~n4978;
  assign n4996 = ~n4986 & n4995;
  assign n4997 = ~n4994 & ~n4996;
  assign n4998 = ~n4988 & ~n4997;
  assign n4999 = po47  & ~n4998;
  assign n5000 = ~n4668 & ~n4676;
  assign n5001 = n4674 & n5000;
  assign n5002 = po34  & n5001;
  assign n5003 = po34  & n5000;
  assign n5004 = ~n4674 & ~n5003;
  assign n5005 = ~n5002 & ~n5004;
  assign n5006 = ~po47  & n4998;
  assign n5007 = ~n5005 & ~n5006;
  assign n5008 = ~n4999 & ~n5007;
  assign n5009 = po48  & ~n5008;
  assign n5010 = ~n4679 & ~n4686;
  assign n5011 = n4685 & n5010;
  assign n5012 = po34  & n5011;
  assign n5013 = po34  & n5010;
  assign n5014 = ~n4685 & ~n5013;
  assign n5015 = ~n5012 & ~n5014;
  assign n5016 = ~po48  & ~n4999;
  assign n5017 = ~n5007 & n5016;
  assign n5018 = ~n5015 & ~n5017;
  assign n5019 = ~n5009 & ~n5018;
  assign n5020 = po49  & ~n5019;
  assign n5021 = ~n4689 & ~n4697;
  assign n5022 = n4695 & n5021;
  assign n5023 = po34  & n5022;
  assign n5024 = po34  & n5021;
  assign n5025 = ~n4695 & ~n5024;
  assign n5026 = ~n5023 & ~n5025;
  assign n5027 = ~po49  & n5019;
  assign n5028 = ~n5026 & ~n5027;
  assign n5029 = ~n5020 & ~n5028;
  assign n5030 = po50  & ~n5029;
  assign n5031 = ~n4700 & ~n4707;
  assign n5032 = n4706 & n5031;
  assign n5033 = po34  & n5032;
  assign n5034 = po34  & n5031;
  assign n5035 = ~n4706 & ~n5034;
  assign n5036 = ~n5033 & ~n5035;
  assign n5037 = ~po50  & ~n5020;
  assign n5038 = ~n5028 & n5037;
  assign n5039 = ~n5036 & ~n5038;
  assign n5040 = ~n5030 & ~n5039;
  assign n5041 = po51  & ~n5040;
  assign n5042 = ~n4710 & ~n4718;
  assign n5043 = n4716 & n5042;
  assign n5044 = po34  & n5043;
  assign n5045 = po34  & n5042;
  assign n5046 = ~n4716 & ~n5045;
  assign n5047 = ~n5044 & ~n5046;
  assign n5048 = ~po51  & n5040;
  assign n5049 = ~n5047 & ~n5048;
  assign n5050 = ~n5041 & ~n5049;
  assign n5051 = po52  & ~n5050;
  assign n5052 = ~n4721 & ~n4728;
  assign n5053 = n4727 & n5052;
  assign n5054 = po34  & n5053;
  assign n5055 = po34  & n5052;
  assign n5056 = ~n4727 & ~n5055;
  assign n5057 = ~n5054 & ~n5056;
  assign n5058 = ~po52  & ~n5041;
  assign n5059 = ~n5049 & n5058;
  assign n5060 = ~n5057 & ~n5059;
  assign n5061 = ~n5051 & ~n5060;
  assign n5062 = po53  & ~n5061;
  assign n5063 = ~n4731 & ~n4739;
  assign n5064 = n4737 & n5063;
  assign n5065 = po34  & n5064;
  assign n5066 = po34  & n5063;
  assign n5067 = ~n4737 & ~n5066;
  assign n5068 = ~n5065 & ~n5067;
  assign n5069 = ~po53  & n5061;
  assign n5070 = ~n5068 & ~n5069;
  assign n5071 = ~n5062 & ~n5070;
  assign n5072 = po54  & ~n5071;
  assign n5073 = ~n4742 & ~n4749;
  assign n5074 = n4748 & n5073;
  assign n5075 = po34  & n5074;
  assign n5076 = po34  & n5073;
  assign n5077 = ~n4748 & ~n5076;
  assign n5078 = ~n5075 & ~n5077;
  assign n5079 = ~po54  & ~n5062;
  assign n5080 = ~n5070 & n5079;
  assign n5081 = ~n5078 & ~n5080;
  assign n5082 = ~n5072 & ~n5081;
  assign n5083 = po55  & ~n5082;
  assign n5084 = ~n4752 & ~n4760;
  assign n5085 = n4758 & n5084;
  assign n5086 = po34  & n5085;
  assign n5087 = po34  & n5084;
  assign n5088 = ~n4758 & ~n5087;
  assign n5089 = ~n5086 & ~n5088;
  assign n5090 = ~po55  & n5082;
  assign n5091 = ~n5089 & ~n5090;
  assign n5092 = ~n5083 & ~n5091;
  assign n5093 = po56  & ~n5092;
  assign n5094 = ~n4763 & ~n4770;
  assign n5095 = n4769 & n5094;
  assign n5096 = po34  & n5095;
  assign n5097 = po34  & n5094;
  assign n5098 = ~n4769 & ~n5097;
  assign n5099 = ~n5096 & ~n5098;
  assign n5100 = ~po56  & ~n5083;
  assign n5101 = ~n5091 & n5100;
  assign n5102 = ~n5099 & ~n5101;
  assign n5103 = ~n5093 & ~n5102;
  assign n5104 = po57  & ~n5103;
  assign n5105 = ~n4773 & ~n4781;
  assign n5106 = n4779 & n5105;
  assign n5107 = po34  & n5106;
  assign n5108 = po34  & n5105;
  assign n5109 = ~n4779 & ~n5108;
  assign n5110 = ~n5107 & ~n5109;
  assign n5111 = ~po57  & n5103;
  assign n5112 = ~n5110 & ~n5111;
  assign n5113 = ~n5104 & ~n5112;
  assign n5114 = po58  & ~n5113;
  assign n5115 = ~n4784 & ~n4791;
  assign n5116 = n4790 & n5115;
  assign n5117 = po34  & n5116;
  assign n5118 = po34  & n5115;
  assign n5119 = ~n4790 & ~n5118;
  assign n5120 = ~n5117 & ~n5119;
  assign n5121 = ~po58  & ~n5104;
  assign n5122 = ~n5112 & n5121;
  assign n5123 = ~n5120 & ~n5122;
  assign n5124 = ~n5114 & ~n5123;
  assign n5125 = po59  & ~n5124;
  assign n5126 = ~n4794 & ~n4802;
  assign n5127 = n4800 & n5126;
  assign n5128 = po34  & n5127;
  assign n5129 = po34  & n5126;
  assign n5130 = ~n4800 & ~n5129;
  assign n5131 = ~n5128 & ~n5130;
  assign n5132 = ~po59  & n5124;
  assign n5133 = ~n5131 & ~n5132;
  assign n5134 = ~n5125 & ~n5133;
  assign n5135 = po60  & ~n5134;
  assign n5136 = ~n4805 & ~n4812;
  assign n5137 = n4811 & n5136;
  assign n5138 = po34  & n5137;
  assign n5139 = po34  & n5136;
  assign n5140 = ~n4811 & ~n5139;
  assign n5141 = ~n5138 & ~n5140;
  assign n5142 = ~po60  & ~n5125;
  assign n5143 = ~n5133 & n5142;
  assign n5144 = ~n5141 & ~n5143;
  assign n5145 = ~n5135 & ~n5144;
  assign n5146 = po61  & ~n5145;
  assign n5147 = ~n4815 & ~n4823;
  assign n5148 = n4821 & n5147;
  assign n5149 = po34  & n5148;
  assign n5150 = po34  & n5147;
  assign n5151 = ~n4821 & ~n5150;
  assign n5152 = ~n5149 & ~n5151;
  assign n5153 = ~po61  & n5145;
  assign n5154 = ~n5152 & ~n5153;
  assign n5155 = ~n5146 & ~n5154;
  assign n5156 = po62  & ~n5155;
  assign n5157 = ~n4826 & ~n4833;
  assign n5158 = n4832 & n5157;
  assign n5159 = po34  & n5158;
  assign n5160 = po34  & n5157;
  assign n5161 = ~n4832 & ~n5160;
  assign n5162 = ~n5159 & ~n5161;
  assign n5163 = ~po62  & ~n5146;
  assign n5164 = ~n5154 & n5163;
  assign n5165 = ~n5162 & ~n5164;
  assign n5166 = ~n5156 & ~n5165;
  assign n5167 = ~n4836 & ~n4838;
  assign n5168 = po34  & n5167;
  assign n5169 = ~n4844 & ~n5168;
  assign n5170 = n4844 & n5168;
  assign n5171 = ~n5169 & ~n5170;
  assign n5172 = ~n4846 & ~n4851;
  assign n5173 = po34  & n5172;
  assign n5174 = ~n4864 & ~n5173;
  assign n5175 = ~n5171 & n5174;
  assign n5176 = ~n5166 & n5175;
  assign n5177 = ~po63  & ~n5176;
  assign n5178 = ~n4851 & po34 ;
  assign n5179 = n4846 & ~n5178;
  assign n5180 = po63  & ~n5172;
  assign n5181 = ~n5179 & n5180;
  assign n5182 = n4851 & ~po34 ;
  assign n5183 = ~n5181 & ~n5182;
  assign n5184 = n5166 & n5171;
  assign n5185 = n5183 & ~n5184;
  assign po33  = n5177 | ~n5185;
  assign n5187 = pi66  & po33 ;
  assign n5188 = ~pi64  & ~pi65 ;
  assign n5189 = ~pi66  & n5188;
  assign n5190 = ~n5187 & ~n5189;
  assign n5191 = po34  & ~n5190;
  assign n5192 = n4863 & ~n5189;
  assign n5193 = ~n4864 & n5192;
  assign n5194 = ~n4857 & n5193;
  assign n5195 = ~n5187 & n5194;
  assign n5196 = ~pi66  & po33 ;
  assign n5197 = pi67  & ~n5196;
  assign n5198 = n4868 & po33 ;
  assign n5199 = ~n5197 & ~n5198;
  assign n5200 = ~n5195 & n5199;
  assign n5201 = ~n5191 & ~n5200;
  assign n5202 = po35  & ~n5201;
  assign n5203 = po34  & n5183;
  assign n5204 = ~n5184 & n5203;
  assign n5205 = ~n5177 & n5204;
  assign n5206 = ~n5198 & ~n5205;
  assign n5207 = pi68  & ~n5206;
  assign n5208 = ~pi68  & n5206;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = ~po35  & n5201;
  assign n5211 = ~n5209 & ~n5210;
  assign n5212 = ~n5202 & ~n5211;
  assign n5213 = po36  & ~n5212;
  assign n5214 = ~n4871 & ~n4875;
  assign n5215 = ~n4879 & n5214;
  assign n5216 = po33  & n5215;
  assign n5217 = po33  & n5214;
  assign n5218 = n4879 & ~n5217;
  assign n5219 = ~n5216 & ~n5218;
  assign n5220 = ~po36  & ~n5202;
  assign n5221 = ~n5211 & n5220;
  assign n5222 = ~n5219 & ~n5221;
  assign n5223 = ~n5213 & ~n5222;
  assign n5224 = po37  & ~n5223;
  assign n5225 = ~n4882 & ~n4884;
  assign n5226 = n4891 & n5225;
  assign n5227 = po33  & n5226;
  assign n5228 = po33  & n5225;
  assign n5229 = ~n4891 & ~n5228;
  assign n5230 = ~n5227 & ~n5229;
  assign n5231 = ~po37  & n5223;
  assign n5232 = ~n5230 & ~n5231;
  assign n5233 = ~n5224 & ~n5232;
  assign n5234 = po38  & ~n5233;
  assign n5235 = ~n4894 & ~n4901;
  assign n5236 = n4900 & n5235;
  assign n5237 = po33  & n5236;
  assign n5238 = po33  & n5235;
  assign n5239 = ~n4900 & ~n5238;
  assign n5240 = ~n5237 & ~n5239;
  assign n5241 = ~po38  & ~n5224;
  assign n5242 = ~n5232 & n5241;
  assign n5243 = ~n5240 & ~n5242;
  assign n5244 = ~n5234 & ~n5243;
  assign n5245 = po39  & ~n5244;
  assign n5246 = ~n4904 & ~n4912;
  assign n5247 = n4910 & n5246;
  assign n5248 = po33  & n5247;
  assign n5249 = po33  & n5246;
  assign n5250 = ~n4910 & ~n5249;
  assign n5251 = ~n5248 & ~n5250;
  assign n5252 = ~po39  & n5244;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = ~n5245 & ~n5253;
  assign n5255 = po40  & ~n5254;
  assign n5256 = ~n4915 & ~n4922;
  assign n5257 = n4921 & n5256;
  assign n5258 = po33  & n5257;
  assign n5259 = po33  & n5256;
  assign n5260 = ~n4921 & ~n5259;
  assign n5261 = ~n5258 & ~n5260;
  assign n5262 = ~po40  & ~n5245;
  assign n5263 = ~n5253 & n5262;
  assign n5264 = ~n5261 & ~n5263;
  assign n5265 = ~n5255 & ~n5264;
  assign n5266 = po41  & ~n5265;
  assign n5267 = ~n4925 & ~n4933;
  assign n5268 = n4931 & n5267;
  assign n5269 = po33  & n5268;
  assign n5270 = po33  & n5267;
  assign n5271 = ~n4931 & ~n5270;
  assign n5272 = ~n5269 & ~n5271;
  assign n5273 = ~po41  & n5265;
  assign n5274 = ~n5272 & ~n5273;
  assign n5275 = ~n5266 & ~n5274;
  assign n5276 = po42  & ~n5275;
  assign n5277 = ~n4936 & ~n4943;
  assign n5278 = n4942 & n5277;
  assign n5279 = po33  & n5278;
  assign n5280 = po33  & n5277;
  assign n5281 = ~n4942 & ~n5280;
  assign n5282 = ~n5279 & ~n5281;
  assign n5283 = ~po42  & ~n5266;
  assign n5284 = ~n5274 & n5283;
  assign n5285 = ~n5282 & ~n5284;
  assign n5286 = ~n5276 & ~n5285;
  assign n5287 = po43  & ~n5286;
  assign n5288 = ~n4946 & ~n4954;
  assign n5289 = n4952 & n5288;
  assign n5290 = po33  & n5289;
  assign n5291 = po33  & n5288;
  assign n5292 = ~n4952 & ~n5291;
  assign n5293 = ~n5290 & ~n5292;
  assign n5294 = ~po43  & n5286;
  assign n5295 = ~n5293 & ~n5294;
  assign n5296 = ~n5287 & ~n5295;
  assign n5297 = po44  & ~n5296;
  assign n5298 = ~n4957 & ~n4964;
  assign n5299 = n4963 & n5298;
  assign n5300 = po33  & n5299;
  assign n5301 = po33  & n5298;
  assign n5302 = ~n4963 & ~n5301;
  assign n5303 = ~n5300 & ~n5302;
  assign n5304 = ~po44  & ~n5287;
  assign n5305 = ~n5295 & n5304;
  assign n5306 = ~n5303 & ~n5305;
  assign n5307 = ~n5297 & ~n5306;
  assign n5308 = po45  & ~n5307;
  assign n5309 = ~n4967 & ~n4975;
  assign n5310 = n4973 & n5309;
  assign n5311 = po33  & n5310;
  assign n5312 = po33  & n5309;
  assign n5313 = ~n4973 & ~n5312;
  assign n5314 = ~n5311 & ~n5313;
  assign n5315 = ~po45  & n5307;
  assign n5316 = ~n5314 & ~n5315;
  assign n5317 = ~n5308 & ~n5316;
  assign n5318 = po46  & ~n5317;
  assign n5319 = ~n4978 & ~n4985;
  assign n5320 = n4984 & n5319;
  assign n5321 = po33  & n5320;
  assign n5322 = po33  & n5319;
  assign n5323 = ~n4984 & ~n5322;
  assign n5324 = ~n5321 & ~n5323;
  assign n5325 = ~po46  & ~n5308;
  assign n5326 = ~n5316 & n5325;
  assign n5327 = ~n5324 & ~n5326;
  assign n5328 = ~n5318 & ~n5327;
  assign n5329 = po47  & ~n5328;
  assign n5330 = ~n4988 & ~n4996;
  assign n5331 = n4994 & n5330;
  assign n5332 = po33  & n5331;
  assign n5333 = po33  & n5330;
  assign n5334 = ~n4994 & ~n5333;
  assign n5335 = ~n5332 & ~n5334;
  assign n5336 = ~po47  & n5328;
  assign n5337 = ~n5335 & ~n5336;
  assign n5338 = ~n5329 & ~n5337;
  assign n5339 = po48  & ~n5338;
  assign n5340 = ~n4999 & ~n5006;
  assign n5341 = n5005 & n5340;
  assign n5342 = po33  & n5341;
  assign n5343 = po33  & n5340;
  assign n5344 = ~n5005 & ~n5343;
  assign n5345 = ~n5342 & ~n5344;
  assign n5346 = ~po48  & ~n5329;
  assign n5347 = ~n5337 & n5346;
  assign n5348 = ~n5345 & ~n5347;
  assign n5349 = ~n5339 & ~n5348;
  assign n5350 = po49  & ~n5349;
  assign n5351 = ~n5009 & ~n5017;
  assign n5352 = n5015 & n5351;
  assign n5353 = po33  & n5352;
  assign n5354 = po33  & n5351;
  assign n5355 = ~n5015 & ~n5354;
  assign n5356 = ~n5353 & ~n5355;
  assign n5357 = ~po49  & n5349;
  assign n5358 = ~n5356 & ~n5357;
  assign n5359 = ~n5350 & ~n5358;
  assign n5360 = po50  & ~n5359;
  assign n5361 = ~n5020 & ~n5027;
  assign n5362 = n5026 & n5361;
  assign n5363 = po33  & n5362;
  assign n5364 = po33  & n5361;
  assign n5365 = ~n5026 & ~n5364;
  assign n5366 = ~n5363 & ~n5365;
  assign n5367 = ~po50  & ~n5350;
  assign n5368 = ~n5358 & n5367;
  assign n5369 = ~n5366 & ~n5368;
  assign n5370 = ~n5360 & ~n5369;
  assign n5371 = po51  & ~n5370;
  assign n5372 = ~n5030 & ~n5038;
  assign n5373 = n5036 & n5372;
  assign n5374 = po33  & n5373;
  assign n5375 = po33  & n5372;
  assign n5376 = ~n5036 & ~n5375;
  assign n5377 = ~n5374 & ~n5376;
  assign n5378 = ~po51  & n5370;
  assign n5379 = ~n5377 & ~n5378;
  assign n5380 = ~n5371 & ~n5379;
  assign n5381 = po52  & ~n5380;
  assign n5382 = ~n5041 & ~n5048;
  assign n5383 = n5047 & n5382;
  assign n5384 = po33  & n5383;
  assign n5385 = po33  & n5382;
  assign n5386 = ~n5047 & ~n5385;
  assign n5387 = ~n5384 & ~n5386;
  assign n5388 = ~po52  & ~n5371;
  assign n5389 = ~n5379 & n5388;
  assign n5390 = ~n5387 & ~n5389;
  assign n5391 = ~n5381 & ~n5390;
  assign n5392 = po53  & ~n5391;
  assign n5393 = ~n5051 & ~n5059;
  assign n5394 = n5057 & n5393;
  assign n5395 = po33  & n5394;
  assign n5396 = po33  & n5393;
  assign n5397 = ~n5057 & ~n5396;
  assign n5398 = ~n5395 & ~n5397;
  assign n5399 = ~po53  & n5391;
  assign n5400 = ~n5398 & ~n5399;
  assign n5401 = ~n5392 & ~n5400;
  assign n5402 = po54  & ~n5401;
  assign n5403 = ~n5062 & ~n5069;
  assign n5404 = n5068 & n5403;
  assign n5405 = po33  & n5404;
  assign n5406 = po33  & n5403;
  assign n5407 = ~n5068 & ~n5406;
  assign n5408 = ~n5405 & ~n5407;
  assign n5409 = ~po54  & ~n5392;
  assign n5410 = ~n5400 & n5409;
  assign n5411 = ~n5408 & ~n5410;
  assign n5412 = ~n5402 & ~n5411;
  assign n5413 = po55  & ~n5412;
  assign n5414 = ~n5072 & ~n5080;
  assign n5415 = n5078 & n5414;
  assign n5416 = po33  & n5415;
  assign n5417 = po33  & n5414;
  assign n5418 = ~n5078 & ~n5417;
  assign n5419 = ~n5416 & ~n5418;
  assign n5420 = ~po55  & n5412;
  assign n5421 = ~n5419 & ~n5420;
  assign n5422 = ~n5413 & ~n5421;
  assign n5423 = po56  & ~n5422;
  assign n5424 = ~n5083 & ~n5090;
  assign n5425 = n5089 & n5424;
  assign n5426 = po33  & n5425;
  assign n5427 = po33  & n5424;
  assign n5428 = ~n5089 & ~n5427;
  assign n5429 = ~n5426 & ~n5428;
  assign n5430 = ~po56  & ~n5413;
  assign n5431 = ~n5421 & n5430;
  assign n5432 = ~n5429 & ~n5431;
  assign n5433 = ~n5423 & ~n5432;
  assign n5434 = po57  & ~n5433;
  assign n5435 = ~n5093 & ~n5101;
  assign n5436 = n5099 & n5435;
  assign n5437 = po33  & n5436;
  assign n5438 = po33  & n5435;
  assign n5439 = ~n5099 & ~n5438;
  assign n5440 = ~n5437 & ~n5439;
  assign n5441 = ~po57  & n5433;
  assign n5442 = ~n5440 & ~n5441;
  assign n5443 = ~n5434 & ~n5442;
  assign n5444 = po58  & ~n5443;
  assign n5445 = ~n5104 & ~n5111;
  assign n5446 = n5110 & n5445;
  assign n5447 = po33  & n5446;
  assign n5448 = po33  & n5445;
  assign n5449 = ~n5110 & ~n5448;
  assign n5450 = ~n5447 & ~n5449;
  assign n5451 = ~po58  & ~n5434;
  assign n5452 = ~n5442 & n5451;
  assign n5453 = ~n5450 & ~n5452;
  assign n5454 = ~n5444 & ~n5453;
  assign n5455 = po59  & ~n5454;
  assign n5456 = ~n5114 & ~n5122;
  assign n5457 = n5120 & n5456;
  assign n5458 = po33  & n5457;
  assign n5459 = po33  & n5456;
  assign n5460 = ~n5120 & ~n5459;
  assign n5461 = ~n5458 & ~n5460;
  assign n5462 = ~po59  & n5454;
  assign n5463 = ~n5461 & ~n5462;
  assign n5464 = ~n5455 & ~n5463;
  assign n5465 = po60  & ~n5464;
  assign n5466 = ~n5125 & ~n5132;
  assign n5467 = n5131 & n5466;
  assign n5468 = po33  & n5467;
  assign n5469 = po33  & n5466;
  assign n5470 = ~n5131 & ~n5469;
  assign n5471 = ~n5468 & ~n5470;
  assign n5472 = ~po60  & ~n5455;
  assign n5473 = ~n5463 & n5472;
  assign n5474 = ~n5471 & ~n5473;
  assign n5475 = ~n5465 & ~n5474;
  assign n5476 = po61  & ~n5475;
  assign n5477 = ~n5135 & ~n5143;
  assign n5478 = n5141 & n5477;
  assign n5479 = po33  & n5478;
  assign n5480 = po33  & n5477;
  assign n5481 = ~n5141 & ~n5480;
  assign n5482 = ~n5479 & ~n5481;
  assign n5483 = ~po61  & n5475;
  assign n5484 = ~n5482 & ~n5483;
  assign n5485 = ~n5476 & ~n5484;
  assign n5486 = po62  & ~n5485;
  assign n5487 = ~n5146 & ~n5153;
  assign n5488 = n5152 & n5487;
  assign n5489 = po33  & n5488;
  assign n5490 = po33  & n5487;
  assign n5491 = ~n5152 & ~n5490;
  assign n5492 = ~n5489 & ~n5491;
  assign n5493 = ~po62  & ~n5476;
  assign n5494 = ~n5484 & n5493;
  assign n5495 = ~n5492 & ~n5494;
  assign n5496 = ~n5486 & ~n5495;
  assign n5497 = ~n5156 & ~n5164;
  assign n5498 = po33  & n5497;
  assign n5499 = ~n5162 & ~n5498;
  assign n5500 = n5162 & n5498;
  assign n5501 = ~n5499 & ~n5500;
  assign n5502 = ~n5166 & ~n5171;
  assign n5503 = po33  & n5502;
  assign n5504 = ~n5184 & ~n5503;
  assign n5505 = ~n5501 & n5504;
  assign n5506 = ~n5496 & n5505;
  assign n5507 = ~po63  & ~n5506;
  assign n5508 = ~n5171 & po33 ;
  assign n5509 = n5166 & ~n5508;
  assign n5510 = po63  & ~n5502;
  assign n5511 = ~n5509 & n5510;
  assign n5512 = n5171 & ~po33 ;
  assign n5513 = ~n5511 & ~n5512;
  assign n5514 = n5496 & n5501;
  assign n5515 = n5513 & ~n5514;
  assign po32  = n5507 | ~n5515;
  assign n5517 = pi64  & po32 ;
  assign n5518 = ~pi62  & ~pi63 ;
  assign n5519 = ~pi64  & n5518;
  assign n5520 = ~n5517 & ~n5519;
  assign n5521 = po33  & ~n5520;
  assign n5522 = ~pi64  & po32 ;
  assign n5523 = pi65  & ~n5522;
  assign n5524 = n5188 & po32 ;
  assign n5525 = ~n5523 & ~n5524;
  assign n5526 = n5183 & ~n5519;
  assign n5527 = ~n5184 & n5526;
  assign n5528 = ~n5177 & n5527;
  assign n5529 = ~n5517 & n5528;
  assign n5530 = n5525 & ~n5529;
  assign n5531 = ~n5521 & ~n5530;
  assign n5532 = po34  & ~n5531;
  assign n5533 = ~po34  & ~n5521;
  assign n5534 = ~n5530 & n5533;
  assign n5535 = po33  & n5513;
  assign n5536 = ~n5514 & n5535;
  assign n5537 = ~n5507 & n5536;
  assign n5538 = ~n5524 & ~n5537;
  assign n5539 = pi66  & ~n5538;
  assign n5540 = ~pi66  & n5538;
  assign n5541 = ~n5539 & ~n5540;
  assign n5542 = ~n5534 & ~n5541;
  assign n5543 = ~n5532 & ~n5542;
  assign n5544 = po35  & ~n5543;
  assign n5545 = ~n5191 & ~n5195;
  assign n5546 = ~n5199 & n5545;
  assign n5547 = po32  & n5546;
  assign n5548 = po32  & n5545;
  assign n5549 = n5199 & ~n5548;
  assign n5550 = ~n5547 & ~n5549;
  assign n5551 = ~po35  & n5543;
  assign n5552 = ~n5550 & ~n5551;
  assign n5553 = ~n5544 & ~n5552;
  assign n5554 = po36  & ~n5553;
  assign n5555 = ~n5202 & ~n5210;
  assign n5556 = n5209 & n5555;
  assign n5557 = po32  & n5556;
  assign n5558 = po32  & n5555;
  assign n5559 = ~n5209 & ~n5558;
  assign n5560 = ~n5557 & ~n5559;
  assign n5561 = ~po36  & ~n5544;
  assign n5562 = ~n5552 & n5561;
  assign n5563 = ~n5560 & ~n5562;
  assign n5564 = ~n5554 & ~n5563;
  assign n5565 = po37  & ~n5564;
  assign n5566 = ~n5213 & ~n5221;
  assign n5567 = n5219 & n5566;
  assign n5568 = po32  & n5567;
  assign n5569 = po32  & n5566;
  assign n5570 = ~n5219 & ~n5569;
  assign n5571 = ~n5568 & ~n5570;
  assign n5572 = ~po37  & n5564;
  assign n5573 = ~n5571 & ~n5572;
  assign n5574 = ~n5565 & ~n5573;
  assign n5575 = po38  & ~n5574;
  assign n5576 = ~n5224 & ~n5231;
  assign n5577 = n5230 & n5576;
  assign n5578 = po32  & n5577;
  assign n5579 = po32  & n5576;
  assign n5580 = ~n5230 & ~n5579;
  assign n5581 = ~n5578 & ~n5580;
  assign n5582 = ~po38  & ~n5565;
  assign n5583 = ~n5573 & n5582;
  assign n5584 = ~n5581 & ~n5583;
  assign n5585 = ~n5575 & ~n5584;
  assign n5586 = po39  & ~n5585;
  assign n5587 = ~n5234 & ~n5242;
  assign n5588 = n5240 & n5587;
  assign n5589 = po32  & n5588;
  assign n5590 = po32  & n5587;
  assign n5591 = ~n5240 & ~n5590;
  assign n5592 = ~n5589 & ~n5591;
  assign n5593 = ~po39  & n5585;
  assign n5594 = ~n5592 & ~n5593;
  assign n5595 = ~n5586 & ~n5594;
  assign n5596 = po40  & ~n5595;
  assign n5597 = ~n5245 & ~n5252;
  assign n5598 = n5251 & n5597;
  assign n5599 = po32  & n5598;
  assign n5600 = po32  & n5597;
  assign n5601 = ~n5251 & ~n5600;
  assign n5602 = ~n5599 & ~n5601;
  assign n5603 = ~po40  & ~n5586;
  assign n5604 = ~n5594 & n5603;
  assign n5605 = ~n5602 & ~n5604;
  assign n5606 = ~n5596 & ~n5605;
  assign n5607 = po41  & ~n5606;
  assign n5608 = ~n5255 & ~n5263;
  assign n5609 = n5261 & n5608;
  assign n5610 = po32  & n5609;
  assign n5611 = po32  & n5608;
  assign n5612 = ~n5261 & ~n5611;
  assign n5613 = ~n5610 & ~n5612;
  assign n5614 = ~po41  & n5606;
  assign n5615 = ~n5613 & ~n5614;
  assign n5616 = ~n5607 & ~n5615;
  assign n5617 = po42  & ~n5616;
  assign n5618 = ~n5266 & ~n5273;
  assign n5619 = n5272 & n5618;
  assign n5620 = po32  & n5619;
  assign n5621 = po32  & n5618;
  assign n5622 = ~n5272 & ~n5621;
  assign n5623 = ~n5620 & ~n5622;
  assign n5624 = ~po42  & ~n5607;
  assign n5625 = ~n5615 & n5624;
  assign n5626 = ~n5623 & ~n5625;
  assign n5627 = ~n5617 & ~n5626;
  assign n5628 = po43  & ~n5627;
  assign n5629 = ~n5276 & ~n5284;
  assign n5630 = n5282 & n5629;
  assign n5631 = po32  & n5630;
  assign n5632 = po32  & n5629;
  assign n5633 = ~n5282 & ~n5632;
  assign n5634 = ~n5631 & ~n5633;
  assign n5635 = ~po43  & n5627;
  assign n5636 = ~n5634 & ~n5635;
  assign n5637 = ~n5628 & ~n5636;
  assign n5638 = po44  & ~n5637;
  assign n5639 = ~n5287 & ~n5294;
  assign n5640 = n5293 & n5639;
  assign n5641 = po32  & n5640;
  assign n5642 = po32  & n5639;
  assign n5643 = ~n5293 & ~n5642;
  assign n5644 = ~n5641 & ~n5643;
  assign n5645 = ~po44  & ~n5628;
  assign n5646 = ~n5636 & n5645;
  assign n5647 = ~n5644 & ~n5646;
  assign n5648 = ~n5638 & ~n5647;
  assign n5649 = po45  & ~n5648;
  assign n5650 = ~n5297 & ~n5305;
  assign n5651 = n5303 & n5650;
  assign n5652 = po32  & n5651;
  assign n5653 = po32  & n5650;
  assign n5654 = ~n5303 & ~n5653;
  assign n5655 = ~n5652 & ~n5654;
  assign n5656 = ~po45  & n5648;
  assign n5657 = ~n5655 & ~n5656;
  assign n5658 = ~n5649 & ~n5657;
  assign n5659 = po46  & ~n5658;
  assign n5660 = ~n5308 & ~n5315;
  assign n5661 = n5314 & n5660;
  assign n5662 = po32  & n5661;
  assign n5663 = po32  & n5660;
  assign n5664 = ~n5314 & ~n5663;
  assign n5665 = ~n5662 & ~n5664;
  assign n5666 = ~po46  & ~n5649;
  assign n5667 = ~n5657 & n5666;
  assign n5668 = ~n5665 & ~n5667;
  assign n5669 = ~n5659 & ~n5668;
  assign n5670 = po47  & ~n5669;
  assign n5671 = ~n5318 & ~n5326;
  assign n5672 = n5324 & n5671;
  assign n5673 = po32  & n5672;
  assign n5674 = po32  & n5671;
  assign n5675 = ~n5324 & ~n5674;
  assign n5676 = ~n5673 & ~n5675;
  assign n5677 = ~po47  & n5669;
  assign n5678 = ~n5676 & ~n5677;
  assign n5679 = ~n5670 & ~n5678;
  assign n5680 = po48  & ~n5679;
  assign n5681 = ~n5329 & ~n5336;
  assign n5682 = n5335 & n5681;
  assign n5683 = po32  & n5682;
  assign n5684 = po32  & n5681;
  assign n5685 = ~n5335 & ~n5684;
  assign n5686 = ~n5683 & ~n5685;
  assign n5687 = ~po48  & ~n5670;
  assign n5688 = ~n5678 & n5687;
  assign n5689 = ~n5686 & ~n5688;
  assign n5690 = ~n5680 & ~n5689;
  assign n5691 = po49  & ~n5690;
  assign n5692 = ~n5339 & ~n5347;
  assign n5693 = n5345 & n5692;
  assign n5694 = po32  & n5693;
  assign n5695 = po32  & n5692;
  assign n5696 = ~n5345 & ~n5695;
  assign n5697 = ~n5694 & ~n5696;
  assign n5698 = ~po49  & n5690;
  assign n5699 = ~n5697 & ~n5698;
  assign n5700 = ~n5691 & ~n5699;
  assign n5701 = po50  & ~n5700;
  assign n5702 = ~n5350 & ~n5357;
  assign n5703 = n5356 & n5702;
  assign n5704 = po32  & n5703;
  assign n5705 = po32  & n5702;
  assign n5706 = ~n5356 & ~n5705;
  assign n5707 = ~n5704 & ~n5706;
  assign n5708 = ~po50  & ~n5691;
  assign n5709 = ~n5699 & n5708;
  assign n5710 = ~n5707 & ~n5709;
  assign n5711 = ~n5701 & ~n5710;
  assign n5712 = po51  & ~n5711;
  assign n5713 = ~n5360 & ~n5368;
  assign n5714 = n5366 & n5713;
  assign n5715 = po32  & n5714;
  assign n5716 = po32  & n5713;
  assign n5717 = ~n5366 & ~n5716;
  assign n5718 = ~n5715 & ~n5717;
  assign n5719 = ~po51  & n5711;
  assign n5720 = ~n5718 & ~n5719;
  assign n5721 = ~n5712 & ~n5720;
  assign n5722 = po52  & ~n5721;
  assign n5723 = ~n5371 & ~n5378;
  assign n5724 = n5377 & n5723;
  assign n5725 = po32  & n5724;
  assign n5726 = po32  & n5723;
  assign n5727 = ~n5377 & ~n5726;
  assign n5728 = ~n5725 & ~n5727;
  assign n5729 = ~po52  & ~n5712;
  assign n5730 = ~n5720 & n5729;
  assign n5731 = ~n5728 & ~n5730;
  assign n5732 = ~n5722 & ~n5731;
  assign n5733 = po53  & ~n5732;
  assign n5734 = ~n5381 & ~n5389;
  assign n5735 = n5387 & n5734;
  assign n5736 = po32  & n5735;
  assign n5737 = po32  & n5734;
  assign n5738 = ~n5387 & ~n5737;
  assign n5739 = ~n5736 & ~n5738;
  assign n5740 = ~po53  & n5732;
  assign n5741 = ~n5739 & ~n5740;
  assign n5742 = ~n5733 & ~n5741;
  assign n5743 = po54  & ~n5742;
  assign n5744 = ~n5392 & ~n5399;
  assign n5745 = n5398 & n5744;
  assign n5746 = po32  & n5745;
  assign n5747 = po32  & n5744;
  assign n5748 = ~n5398 & ~n5747;
  assign n5749 = ~n5746 & ~n5748;
  assign n5750 = ~po54  & ~n5733;
  assign n5751 = ~n5741 & n5750;
  assign n5752 = ~n5749 & ~n5751;
  assign n5753 = ~n5743 & ~n5752;
  assign n5754 = po55  & ~n5753;
  assign n5755 = ~n5402 & ~n5410;
  assign n5756 = n5408 & n5755;
  assign n5757 = po32  & n5756;
  assign n5758 = po32  & n5755;
  assign n5759 = ~n5408 & ~n5758;
  assign n5760 = ~n5757 & ~n5759;
  assign n5761 = ~po55  & n5753;
  assign n5762 = ~n5760 & ~n5761;
  assign n5763 = ~n5754 & ~n5762;
  assign n5764 = po56  & ~n5763;
  assign n5765 = ~n5413 & ~n5420;
  assign n5766 = n5419 & n5765;
  assign n5767 = po32  & n5766;
  assign n5768 = po32  & n5765;
  assign n5769 = ~n5419 & ~n5768;
  assign n5770 = ~n5767 & ~n5769;
  assign n5771 = ~po56  & ~n5754;
  assign n5772 = ~n5762 & n5771;
  assign n5773 = ~n5770 & ~n5772;
  assign n5774 = ~n5764 & ~n5773;
  assign n5775 = po57  & ~n5774;
  assign n5776 = ~n5423 & ~n5431;
  assign n5777 = n5429 & n5776;
  assign n5778 = po32  & n5777;
  assign n5779 = po32  & n5776;
  assign n5780 = ~n5429 & ~n5779;
  assign n5781 = ~n5778 & ~n5780;
  assign n5782 = ~po57  & n5774;
  assign n5783 = ~n5781 & ~n5782;
  assign n5784 = ~n5775 & ~n5783;
  assign n5785 = po58  & ~n5784;
  assign n5786 = ~n5434 & ~n5441;
  assign n5787 = n5440 & n5786;
  assign n5788 = po32  & n5787;
  assign n5789 = po32  & n5786;
  assign n5790 = ~n5440 & ~n5789;
  assign n5791 = ~n5788 & ~n5790;
  assign n5792 = ~po58  & ~n5775;
  assign n5793 = ~n5783 & n5792;
  assign n5794 = ~n5791 & ~n5793;
  assign n5795 = ~n5785 & ~n5794;
  assign n5796 = po59  & ~n5795;
  assign n5797 = ~n5444 & ~n5452;
  assign n5798 = n5450 & n5797;
  assign n5799 = po32  & n5798;
  assign n5800 = po32  & n5797;
  assign n5801 = ~n5450 & ~n5800;
  assign n5802 = ~n5799 & ~n5801;
  assign n5803 = ~po59  & n5795;
  assign n5804 = ~n5802 & ~n5803;
  assign n5805 = ~n5796 & ~n5804;
  assign n5806 = po60  & ~n5805;
  assign n5807 = ~n5455 & ~n5462;
  assign n5808 = n5461 & n5807;
  assign n5809 = po32  & n5808;
  assign n5810 = po32  & n5807;
  assign n5811 = ~n5461 & ~n5810;
  assign n5812 = ~n5809 & ~n5811;
  assign n5813 = ~po60  & ~n5796;
  assign n5814 = ~n5804 & n5813;
  assign n5815 = ~n5812 & ~n5814;
  assign n5816 = ~n5806 & ~n5815;
  assign n5817 = po61  & ~n5816;
  assign n5818 = ~n5465 & ~n5473;
  assign n5819 = n5471 & n5818;
  assign n5820 = po32  & n5819;
  assign n5821 = po32  & n5818;
  assign n5822 = ~n5471 & ~n5821;
  assign n5823 = ~n5820 & ~n5822;
  assign n5824 = ~po61  & n5816;
  assign n5825 = ~n5823 & ~n5824;
  assign n5826 = ~n5817 & ~n5825;
  assign n5827 = po62  & ~n5826;
  assign n5828 = ~n5476 & ~n5483;
  assign n5829 = n5482 & n5828;
  assign n5830 = po32  & n5829;
  assign n5831 = po32  & n5828;
  assign n5832 = ~n5482 & ~n5831;
  assign n5833 = ~n5830 & ~n5832;
  assign n5834 = ~po62  & ~n5817;
  assign n5835 = ~n5825 & n5834;
  assign n5836 = ~n5833 & ~n5835;
  assign n5837 = ~n5827 & ~n5836;
  assign n5838 = ~n5486 & ~n5494;
  assign n5839 = po32  & n5838;
  assign n5840 = ~n5492 & ~n5839;
  assign n5841 = n5492 & n5839;
  assign n5842 = ~n5840 & ~n5841;
  assign n5843 = ~n5496 & ~n5501;
  assign n5844 = po32  & n5843;
  assign n5845 = ~n5514 & ~n5844;
  assign n5846 = ~n5842 & n5845;
  assign n5847 = ~n5837 & n5846;
  assign n5848 = ~po63  & ~n5847;
  assign n5849 = ~n5501 & po32 ;
  assign n5850 = n5496 & ~n5849;
  assign n5851 = po63  & ~n5843;
  assign n5852 = ~n5850 & n5851;
  assign n5853 = n5501 & ~po32 ;
  assign n5854 = ~n5852 & ~n5853;
  assign n5855 = n5837 & n5842;
  assign n5856 = n5854 & ~n5855;
  assign po31  = n5848 | ~n5856;
  assign n5858 = pi62  & po31 ;
  assign n5859 = ~pi60  & ~pi61 ;
  assign n5860 = ~pi62  & n5859;
  assign n5861 = ~n5858 & ~n5860;
  assign n5862 = po32  & ~n5861;
  assign n5863 = n5513 & ~n5860;
  assign n5864 = ~n5514 & n5863;
  assign n5865 = ~n5507 & n5864;
  assign n5866 = ~n5858 & n5865;
  assign n5867 = ~pi62  & po31 ;
  assign n5868 = pi63  & ~n5867;
  assign n5869 = n5518 & po31 ;
  assign n5870 = ~n5868 & ~n5869;
  assign n5871 = ~n5866 & n5870;
  assign n5872 = ~n5862 & ~n5871;
  assign n5873 = po33  & ~n5872;
  assign n5874 = po32  & n5854;
  assign n5875 = ~n5855 & n5874;
  assign n5876 = ~n5848 & n5875;
  assign n5877 = ~n5869 & ~n5876;
  assign n5878 = pi64  & ~n5877;
  assign n5879 = ~pi64  & n5877;
  assign n5880 = ~n5878 & ~n5879;
  assign n5881 = ~po33  & n5872;
  assign n5882 = ~n5880 & ~n5881;
  assign n5883 = ~n5873 & ~n5882;
  assign n5884 = po34  & ~n5883;
  assign n5885 = ~po34  & ~n5873;
  assign n5886 = ~n5882 & n5885;
  assign n5887 = ~n5521 & ~n5529;
  assign n5888 = ~n5525 & n5887;
  assign n5889 = po31  & n5888;
  assign n5890 = po31  & n5887;
  assign n5891 = n5525 & ~n5890;
  assign n5892 = ~n5889 & ~n5891;
  assign n5893 = ~n5886 & ~n5892;
  assign n5894 = ~n5884 & ~n5893;
  assign n5895 = po35  & ~n5894;
  assign n5896 = ~n5532 & ~n5534;
  assign n5897 = n5541 & n5896;
  assign n5898 = po31  & n5897;
  assign n5899 = po31  & n5896;
  assign n5900 = ~n5541 & ~n5899;
  assign n5901 = ~n5898 & ~n5900;
  assign n5902 = ~po35  & n5894;
  assign n5903 = ~n5901 & ~n5902;
  assign n5904 = ~n5895 & ~n5903;
  assign n5905 = po36  & ~n5904;
  assign n5906 = ~n5544 & ~n5551;
  assign n5907 = n5550 & n5906;
  assign n5908 = po31  & n5907;
  assign n5909 = po31  & n5906;
  assign n5910 = ~n5550 & ~n5909;
  assign n5911 = ~n5908 & ~n5910;
  assign n5912 = ~po36  & ~n5895;
  assign n5913 = ~n5903 & n5912;
  assign n5914 = ~n5911 & ~n5913;
  assign n5915 = ~n5905 & ~n5914;
  assign n5916 = po37  & ~n5915;
  assign n5917 = ~n5554 & ~n5562;
  assign n5918 = n5560 & n5917;
  assign n5919 = po31  & n5918;
  assign n5920 = po31  & n5917;
  assign n5921 = ~n5560 & ~n5920;
  assign n5922 = ~n5919 & ~n5921;
  assign n5923 = ~po37  & n5915;
  assign n5924 = ~n5922 & ~n5923;
  assign n5925 = ~n5916 & ~n5924;
  assign n5926 = po38  & ~n5925;
  assign n5927 = ~n5565 & ~n5572;
  assign n5928 = n5571 & n5927;
  assign n5929 = po31  & n5928;
  assign n5930 = po31  & n5927;
  assign n5931 = ~n5571 & ~n5930;
  assign n5932 = ~n5929 & ~n5931;
  assign n5933 = ~po38  & ~n5916;
  assign n5934 = ~n5924 & n5933;
  assign n5935 = ~n5932 & ~n5934;
  assign n5936 = ~n5926 & ~n5935;
  assign n5937 = po39  & ~n5936;
  assign n5938 = ~n5575 & ~n5583;
  assign n5939 = n5581 & n5938;
  assign n5940 = po31  & n5939;
  assign n5941 = po31  & n5938;
  assign n5942 = ~n5581 & ~n5941;
  assign n5943 = ~n5940 & ~n5942;
  assign n5944 = ~po39  & n5936;
  assign n5945 = ~n5943 & ~n5944;
  assign n5946 = ~n5937 & ~n5945;
  assign n5947 = po40  & ~n5946;
  assign n5948 = ~n5586 & ~n5593;
  assign n5949 = n5592 & n5948;
  assign n5950 = po31  & n5949;
  assign n5951 = po31  & n5948;
  assign n5952 = ~n5592 & ~n5951;
  assign n5953 = ~n5950 & ~n5952;
  assign n5954 = ~po40  & ~n5937;
  assign n5955 = ~n5945 & n5954;
  assign n5956 = ~n5953 & ~n5955;
  assign n5957 = ~n5947 & ~n5956;
  assign n5958 = po41  & ~n5957;
  assign n5959 = ~n5596 & ~n5604;
  assign n5960 = n5602 & n5959;
  assign n5961 = po31  & n5960;
  assign n5962 = po31  & n5959;
  assign n5963 = ~n5602 & ~n5962;
  assign n5964 = ~n5961 & ~n5963;
  assign n5965 = ~po41  & n5957;
  assign n5966 = ~n5964 & ~n5965;
  assign n5967 = ~n5958 & ~n5966;
  assign n5968 = po42  & ~n5967;
  assign n5969 = ~n5607 & ~n5614;
  assign n5970 = n5613 & n5969;
  assign n5971 = po31  & n5970;
  assign n5972 = po31  & n5969;
  assign n5973 = ~n5613 & ~n5972;
  assign n5974 = ~n5971 & ~n5973;
  assign n5975 = ~po42  & ~n5958;
  assign n5976 = ~n5966 & n5975;
  assign n5977 = ~n5974 & ~n5976;
  assign n5978 = ~n5968 & ~n5977;
  assign n5979 = po43  & ~n5978;
  assign n5980 = ~n5617 & ~n5625;
  assign n5981 = n5623 & n5980;
  assign n5982 = po31  & n5981;
  assign n5983 = po31  & n5980;
  assign n5984 = ~n5623 & ~n5983;
  assign n5985 = ~n5982 & ~n5984;
  assign n5986 = ~po43  & n5978;
  assign n5987 = ~n5985 & ~n5986;
  assign n5988 = ~n5979 & ~n5987;
  assign n5989 = po44  & ~n5988;
  assign n5990 = ~n5628 & ~n5635;
  assign n5991 = n5634 & n5990;
  assign n5992 = po31  & n5991;
  assign n5993 = po31  & n5990;
  assign n5994 = ~n5634 & ~n5993;
  assign n5995 = ~n5992 & ~n5994;
  assign n5996 = ~po44  & ~n5979;
  assign n5997 = ~n5987 & n5996;
  assign n5998 = ~n5995 & ~n5997;
  assign n5999 = ~n5989 & ~n5998;
  assign n6000 = po45  & ~n5999;
  assign n6001 = ~n5638 & ~n5646;
  assign n6002 = n5644 & n6001;
  assign n6003 = po31  & n6002;
  assign n6004 = po31  & n6001;
  assign n6005 = ~n5644 & ~n6004;
  assign n6006 = ~n6003 & ~n6005;
  assign n6007 = ~po45  & n5999;
  assign n6008 = ~n6006 & ~n6007;
  assign n6009 = ~n6000 & ~n6008;
  assign n6010 = po46  & ~n6009;
  assign n6011 = ~n5649 & ~n5656;
  assign n6012 = n5655 & n6011;
  assign n6013 = po31  & n6012;
  assign n6014 = po31  & n6011;
  assign n6015 = ~n5655 & ~n6014;
  assign n6016 = ~n6013 & ~n6015;
  assign n6017 = ~po46  & ~n6000;
  assign n6018 = ~n6008 & n6017;
  assign n6019 = ~n6016 & ~n6018;
  assign n6020 = ~n6010 & ~n6019;
  assign n6021 = po47  & ~n6020;
  assign n6022 = ~n5659 & ~n5667;
  assign n6023 = n5665 & n6022;
  assign n6024 = po31  & n6023;
  assign n6025 = po31  & n6022;
  assign n6026 = ~n5665 & ~n6025;
  assign n6027 = ~n6024 & ~n6026;
  assign n6028 = ~po47  & n6020;
  assign n6029 = ~n6027 & ~n6028;
  assign n6030 = ~n6021 & ~n6029;
  assign n6031 = po48  & ~n6030;
  assign n6032 = ~n5670 & ~n5677;
  assign n6033 = n5676 & n6032;
  assign n6034 = po31  & n6033;
  assign n6035 = po31  & n6032;
  assign n6036 = ~n5676 & ~n6035;
  assign n6037 = ~n6034 & ~n6036;
  assign n6038 = ~po48  & ~n6021;
  assign n6039 = ~n6029 & n6038;
  assign n6040 = ~n6037 & ~n6039;
  assign n6041 = ~n6031 & ~n6040;
  assign n6042 = po49  & ~n6041;
  assign n6043 = ~n5680 & ~n5688;
  assign n6044 = n5686 & n6043;
  assign n6045 = po31  & n6044;
  assign n6046 = po31  & n6043;
  assign n6047 = ~n5686 & ~n6046;
  assign n6048 = ~n6045 & ~n6047;
  assign n6049 = ~po49  & n6041;
  assign n6050 = ~n6048 & ~n6049;
  assign n6051 = ~n6042 & ~n6050;
  assign n6052 = po50  & ~n6051;
  assign n6053 = ~n5691 & ~n5698;
  assign n6054 = n5697 & n6053;
  assign n6055 = po31  & n6054;
  assign n6056 = po31  & n6053;
  assign n6057 = ~n5697 & ~n6056;
  assign n6058 = ~n6055 & ~n6057;
  assign n6059 = ~po50  & ~n6042;
  assign n6060 = ~n6050 & n6059;
  assign n6061 = ~n6058 & ~n6060;
  assign n6062 = ~n6052 & ~n6061;
  assign n6063 = po51  & ~n6062;
  assign n6064 = ~n5701 & ~n5709;
  assign n6065 = n5707 & n6064;
  assign n6066 = po31  & n6065;
  assign n6067 = po31  & n6064;
  assign n6068 = ~n5707 & ~n6067;
  assign n6069 = ~n6066 & ~n6068;
  assign n6070 = ~po51  & n6062;
  assign n6071 = ~n6069 & ~n6070;
  assign n6072 = ~n6063 & ~n6071;
  assign n6073 = po52  & ~n6072;
  assign n6074 = ~n5712 & ~n5719;
  assign n6075 = n5718 & n6074;
  assign n6076 = po31  & n6075;
  assign n6077 = po31  & n6074;
  assign n6078 = ~n5718 & ~n6077;
  assign n6079 = ~n6076 & ~n6078;
  assign n6080 = ~po52  & ~n6063;
  assign n6081 = ~n6071 & n6080;
  assign n6082 = ~n6079 & ~n6081;
  assign n6083 = ~n6073 & ~n6082;
  assign n6084 = po53  & ~n6083;
  assign n6085 = ~n5722 & ~n5730;
  assign n6086 = n5728 & n6085;
  assign n6087 = po31  & n6086;
  assign n6088 = po31  & n6085;
  assign n6089 = ~n5728 & ~n6088;
  assign n6090 = ~n6087 & ~n6089;
  assign n6091 = ~po53  & n6083;
  assign n6092 = ~n6090 & ~n6091;
  assign n6093 = ~n6084 & ~n6092;
  assign n6094 = po54  & ~n6093;
  assign n6095 = ~n5733 & ~n5740;
  assign n6096 = n5739 & n6095;
  assign n6097 = po31  & n6096;
  assign n6098 = po31  & n6095;
  assign n6099 = ~n5739 & ~n6098;
  assign n6100 = ~n6097 & ~n6099;
  assign n6101 = ~po54  & ~n6084;
  assign n6102 = ~n6092 & n6101;
  assign n6103 = ~n6100 & ~n6102;
  assign n6104 = ~n6094 & ~n6103;
  assign n6105 = po55  & ~n6104;
  assign n6106 = ~n5743 & ~n5751;
  assign n6107 = n5749 & n6106;
  assign n6108 = po31  & n6107;
  assign n6109 = po31  & n6106;
  assign n6110 = ~n5749 & ~n6109;
  assign n6111 = ~n6108 & ~n6110;
  assign n6112 = ~po55  & n6104;
  assign n6113 = ~n6111 & ~n6112;
  assign n6114 = ~n6105 & ~n6113;
  assign n6115 = po56  & ~n6114;
  assign n6116 = ~n5754 & ~n5761;
  assign n6117 = n5760 & n6116;
  assign n6118 = po31  & n6117;
  assign n6119 = po31  & n6116;
  assign n6120 = ~n5760 & ~n6119;
  assign n6121 = ~n6118 & ~n6120;
  assign n6122 = ~po56  & ~n6105;
  assign n6123 = ~n6113 & n6122;
  assign n6124 = ~n6121 & ~n6123;
  assign n6125 = ~n6115 & ~n6124;
  assign n6126 = po57  & ~n6125;
  assign n6127 = ~n5764 & ~n5772;
  assign n6128 = n5770 & n6127;
  assign n6129 = po31  & n6128;
  assign n6130 = po31  & n6127;
  assign n6131 = ~n5770 & ~n6130;
  assign n6132 = ~n6129 & ~n6131;
  assign n6133 = ~po57  & n6125;
  assign n6134 = ~n6132 & ~n6133;
  assign n6135 = ~n6126 & ~n6134;
  assign n6136 = po58  & ~n6135;
  assign n6137 = ~n5775 & ~n5782;
  assign n6138 = n5781 & n6137;
  assign n6139 = po31  & n6138;
  assign n6140 = po31  & n6137;
  assign n6141 = ~n5781 & ~n6140;
  assign n6142 = ~n6139 & ~n6141;
  assign n6143 = ~po58  & ~n6126;
  assign n6144 = ~n6134 & n6143;
  assign n6145 = ~n6142 & ~n6144;
  assign n6146 = ~n6136 & ~n6145;
  assign n6147 = po59  & ~n6146;
  assign n6148 = ~n5785 & ~n5793;
  assign n6149 = n5791 & n6148;
  assign n6150 = po31  & n6149;
  assign n6151 = po31  & n6148;
  assign n6152 = ~n5791 & ~n6151;
  assign n6153 = ~n6150 & ~n6152;
  assign n6154 = ~po59  & n6146;
  assign n6155 = ~n6153 & ~n6154;
  assign n6156 = ~n6147 & ~n6155;
  assign n6157 = po60  & ~n6156;
  assign n6158 = ~n5796 & ~n5803;
  assign n6159 = n5802 & n6158;
  assign n6160 = po31  & n6159;
  assign n6161 = po31  & n6158;
  assign n6162 = ~n5802 & ~n6161;
  assign n6163 = ~n6160 & ~n6162;
  assign n6164 = ~po60  & ~n6147;
  assign n6165 = ~n6155 & n6164;
  assign n6166 = ~n6163 & ~n6165;
  assign n6167 = ~n6157 & ~n6166;
  assign n6168 = po61  & ~n6167;
  assign n6169 = ~n5806 & ~n5814;
  assign n6170 = n5812 & n6169;
  assign n6171 = po31  & n6170;
  assign n6172 = po31  & n6169;
  assign n6173 = ~n5812 & ~n6172;
  assign n6174 = ~n6171 & ~n6173;
  assign n6175 = ~po61  & n6167;
  assign n6176 = ~n6174 & ~n6175;
  assign n6177 = ~n6168 & ~n6176;
  assign n6178 = po62  & ~n6177;
  assign n6179 = ~n5817 & ~n5824;
  assign n6180 = n5823 & n6179;
  assign n6181 = po31  & n6180;
  assign n6182 = po31  & n6179;
  assign n6183 = ~n5823 & ~n6182;
  assign n6184 = ~n6181 & ~n6183;
  assign n6185 = ~po62  & ~n6168;
  assign n6186 = ~n6176 & n6185;
  assign n6187 = ~n6184 & ~n6186;
  assign n6188 = ~n6178 & ~n6187;
  assign n6189 = ~n5827 & ~n5835;
  assign n6190 = po31  & n6189;
  assign n6191 = ~n5833 & ~n6190;
  assign n6192 = n5833 & n6190;
  assign n6193 = ~n6191 & ~n6192;
  assign n6194 = ~n5837 & ~n5842;
  assign n6195 = po31  & n6194;
  assign n6196 = ~n5855 & ~n6195;
  assign n6197 = ~n6193 & n6196;
  assign n6198 = ~n6188 & n6197;
  assign n6199 = ~po63  & ~n6198;
  assign n6200 = ~n5842 & po31 ;
  assign n6201 = n5837 & ~n6200;
  assign n6202 = po63  & ~n6194;
  assign n6203 = ~n6201 & n6202;
  assign n6204 = n5842 & ~po31 ;
  assign n6205 = ~n6203 & ~n6204;
  assign n6206 = n6188 & n6193;
  assign n6207 = n6205 & ~n6206;
  assign po30  = n6199 | ~n6207;
  assign n6209 = pi60  & po30 ;
  assign n6210 = ~pi58  & ~pi59 ;
  assign n6211 = ~pi60  & n6210;
  assign n6212 = ~n6209 & ~n6211;
  assign n6213 = po31  & ~n6212;
  assign n6214 = n5854 & ~n6211;
  assign n6215 = ~n5855 & n6214;
  assign n6216 = ~n5848 & n6215;
  assign n6217 = ~n6209 & n6216;
  assign n6218 = ~pi60  & po30 ;
  assign n6219 = pi61  & ~n6218;
  assign n6220 = n5859 & po30 ;
  assign n6221 = ~n6219 & ~n6220;
  assign n6222 = ~n6217 & n6221;
  assign n6223 = ~n6213 & ~n6222;
  assign n6224 = po32  & ~n6223;
  assign n6225 = ~po32  & ~n6213;
  assign n6226 = ~n6222 & n6225;
  assign n6227 = po31  & n6205;
  assign n6228 = ~n6206 & n6227;
  assign n6229 = ~n6199 & n6228;
  assign n6230 = ~n6220 & ~n6229;
  assign n6231 = pi62  & ~n6230;
  assign n6232 = ~pi62  & n6230;
  assign n6233 = ~n6231 & ~n6232;
  assign n6234 = ~n6226 & ~n6233;
  assign n6235 = ~n6224 & ~n6234;
  assign n6236 = po33  & ~n6235;
  assign n6237 = ~n5862 & ~n5866;
  assign n6238 = ~n5870 & n6237;
  assign n6239 = po30  & n6238;
  assign n6240 = po30  & n6237;
  assign n6241 = n5870 & ~n6240;
  assign n6242 = ~n6239 & ~n6241;
  assign n6243 = ~po33  & n6235;
  assign n6244 = ~n6242 & ~n6243;
  assign n6245 = ~n6236 & ~n6244;
  assign n6246 = po34  & ~n6245;
  assign n6247 = ~n5873 & ~n5881;
  assign n6248 = n5880 & n6247;
  assign n6249 = po30  & n6248;
  assign n6250 = po30  & n6247;
  assign n6251 = ~n5880 & ~n6250;
  assign n6252 = ~n6249 & ~n6251;
  assign n6253 = ~po34  & ~n6236;
  assign n6254 = ~n6244 & n6253;
  assign n6255 = ~n6252 & ~n6254;
  assign n6256 = ~n6246 & ~n6255;
  assign n6257 = po35  & ~n6256;
  assign n6258 = ~n5884 & ~n5886;
  assign n6259 = n5892 & n6258;
  assign n6260 = po30  & n6259;
  assign n6261 = po30  & n6258;
  assign n6262 = ~n5892 & ~n6261;
  assign n6263 = ~n6260 & ~n6262;
  assign n6264 = ~po35  & n6256;
  assign n6265 = ~n6263 & ~n6264;
  assign n6266 = ~n6257 & ~n6265;
  assign n6267 = po36  & ~n6266;
  assign n6268 = ~n5895 & ~n5902;
  assign n6269 = n5901 & n6268;
  assign n6270 = po30  & n6269;
  assign n6271 = po30  & n6268;
  assign n6272 = ~n5901 & ~n6271;
  assign n6273 = ~n6270 & ~n6272;
  assign n6274 = ~po36  & ~n6257;
  assign n6275 = ~n6265 & n6274;
  assign n6276 = ~n6273 & ~n6275;
  assign n6277 = ~n6267 & ~n6276;
  assign n6278 = po37  & ~n6277;
  assign n6279 = ~n5905 & ~n5913;
  assign n6280 = n5911 & n6279;
  assign n6281 = po30  & n6280;
  assign n6282 = po30  & n6279;
  assign n6283 = ~n5911 & ~n6282;
  assign n6284 = ~n6281 & ~n6283;
  assign n6285 = ~po37  & n6277;
  assign n6286 = ~n6284 & ~n6285;
  assign n6287 = ~n6278 & ~n6286;
  assign n6288 = po38  & ~n6287;
  assign n6289 = ~n5916 & ~n5923;
  assign n6290 = n5922 & n6289;
  assign n6291 = po30  & n6290;
  assign n6292 = po30  & n6289;
  assign n6293 = ~n5922 & ~n6292;
  assign n6294 = ~n6291 & ~n6293;
  assign n6295 = ~po38  & ~n6278;
  assign n6296 = ~n6286 & n6295;
  assign n6297 = ~n6294 & ~n6296;
  assign n6298 = ~n6288 & ~n6297;
  assign n6299 = po39  & ~n6298;
  assign n6300 = ~n5926 & ~n5934;
  assign n6301 = n5932 & n6300;
  assign n6302 = po30  & n6301;
  assign n6303 = po30  & n6300;
  assign n6304 = ~n5932 & ~n6303;
  assign n6305 = ~n6302 & ~n6304;
  assign n6306 = ~po39  & n6298;
  assign n6307 = ~n6305 & ~n6306;
  assign n6308 = ~n6299 & ~n6307;
  assign n6309 = po40  & ~n6308;
  assign n6310 = ~n5937 & ~n5944;
  assign n6311 = n5943 & n6310;
  assign n6312 = po30  & n6311;
  assign n6313 = po30  & n6310;
  assign n6314 = ~n5943 & ~n6313;
  assign n6315 = ~n6312 & ~n6314;
  assign n6316 = ~po40  & ~n6299;
  assign n6317 = ~n6307 & n6316;
  assign n6318 = ~n6315 & ~n6317;
  assign n6319 = ~n6309 & ~n6318;
  assign n6320 = po41  & ~n6319;
  assign n6321 = ~n5947 & ~n5955;
  assign n6322 = n5953 & n6321;
  assign n6323 = po30  & n6322;
  assign n6324 = po30  & n6321;
  assign n6325 = ~n5953 & ~n6324;
  assign n6326 = ~n6323 & ~n6325;
  assign n6327 = ~po41  & n6319;
  assign n6328 = ~n6326 & ~n6327;
  assign n6329 = ~n6320 & ~n6328;
  assign n6330 = po42  & ~n6329;
  assign n6331 = ~n5958 & ~n5965;
  assign n6332 = n5964 & n6331;
  assign n6333 = po30  & n6332;
  assign n6334 = po30  & n6331;
  assign n6335 = ~n5964 & ~n6334;
  assign n6336 = ~n6333 & ~n6335;
  assign n6337 = ~po42  & ~n6320;
  assign n6338 = ~n6328 & n6337;
  assign n6339 = ~n6336 & ~n6338;
  assign n6340 = ~n6330 & ~n6339;
  assign n6341 = po43  & ~n6340;
  assign n6342 = ~n5968 & ~n5976;
  assign n6343 = n5974 & n6342;
  assign n6344 = po30  & n6343;
  assign n6345 = po30  & n6342;
  assign n6346 = ~n5974 & ~n6345;
  assign n6347 = ~n6344 & ~n6346;
  assign n6348 = ~po43  & n6340;
  assign n6349 = ~n6347 & ~n6348;
  assign n6350 = ~n6341 & ~n6349;
  assign n6351 = po44  & ~n6350;
  assign n6352 = ~n5979 & ~n5986;
  assign n6353 = n5985 & n6352;
  assign n6354 = po30  & n6353;
  assign n6355 = po30  & n6352;
  assign n6356 = ~n5985 & ~n6355;
  assign n6357 = ~n6354 & ~n6356;
  assign n6358 = ~po44  & ~n6341;
  assign n6359 = ~n6349 & n6358;
  assign n6360 = ~n6357 & ~n6359;
  assign n6361 = ~n6351 & ~n6360;
  assign n6362 = po45  & ~n6361;
  assign n6363 = ~n5989 & ~n5997;
  assign n6364 = n5995 & n6363;
  assign n6365 = po30  & n6364;
  assign n6366 = po30  & n6363;
  assign n6367 = ~n5995 & ~n6366;
  assign n6368 = ~n6365 & ~n6367;
  assign n6369 = ~po45  & n6361;
  assign n6370 = ~n6368 & ~n6369;
  assign n6371 = ~n6362 & ~n6370;
  assign n6372 = po46  & ~n6371;
  assign n6373 = ~n6000 & ~n6007;
  assign n6374 = n6006 & n6373;
  assign n6375 = po30  & n6374;
  assign n6376 = po30  & n6373;
  assign n6377 = ~n6006 & ~n6376;
  assign n6378 = ~n6375 & ~n6377;
  assign n6379 = ~po46  & ~n6362;
  assign n6380 = ~n6370 & n6379;
  assign n6381 = ~n6378 & ~n6380;
  assign n6382 = ~n6372 & ~n6381;
  assign n6383 = po47  & ~n6382;
  assign n6384 = ~n6010 & ~n6018;
  assign n6385 = n6016 & n6384;
  assign n6386 = po30  & n6385;
  assign n6387 = po30  & n6384;
  assign n6388 = ~n6016 & ~n6387;
  assign n6389 = ~n6386 & ~n6388;
  assign n6390 = ~po47  & n6382;
  assign n6391 = ~n6389 & ~n6390;
  assign n6392 = ~n6383 & ~n6391;
  assign n6393 = po48  & ~n6392;
  assign n6394 = ~n6021 & ~n6028;
  assign n6395 = n6027 & n6394;
  assign n6396 = po30  & n6395;
  assign n6397 = po30  & n6394;
  assign n6398 = ~n6027 & ~n6397;
  assign n6399 = ~n6396 & ~n6398;
  assign n6400 = ~po48  & ~n6383;
  assign n6401 = ~n6391 & n6400;
  assign n6402 = ~n6399 & ~n6401;
  assign n6403 = ~n6393 & ~n6402;
  assign n6404 = po49  & ~n6403;
  assign n6405 = ~n6031 & ~n6039;
  assign n6406 = n6037 & n6405;
  assign n6407 = po30  & n6406;
  assign n6408 = po30  & n6405;
  assign n6409 = ~n6037 & ~n6408;
  assign n6410 = ~n6407 & ~n6409;
  assign n6411 = ~po49  & n6403;
  assign n6412 = ~n6410 & ~n6411;
  assign n6413 = ~n6404 & ~n6412;
  assign n6414 = po50  & ~n6413;
  assign n6415 = ~n6042 & ~n6049;
  assign n6416 = n6048 & n6415;
  assign n6417 = po30  & n6416;
  assign n6418 = po30  & n6415;
  assign n6419 = ~n6048 & ~n6418;
  assign n6420 = ~n6417 & ~n6419;
  assign n6421 = ~po50  & ~n6404;
  assign n6422 = ~n6412 & n6421;
  assign n6423 = ~n6420 & ~n6422;
  assign n6424 = ~n6414 & ~n6423;
  assign n6425 = po51  & ~n6424;
  assign n6426 = ~n6052 & ~n6060;
  assign n6427 = n6058 & n6426;
  assign n6428 = po30  & n6427;
  assign n6429 = po30  & n6426;
  assign n6430 = ~n6058 & ~n6429;
  assign n6431 = ~n6428 & ~n6430;
  assign n6432 = ~po51  & n6424;
  assign n6433 = ~n6431 & ~n6432;
  assign n6434 = ~n6425 & ~n6433;
  assign n6435 = po52  & ~n6434;
  assign n6436 = ~n6063 & ~n6070;
  assign n6437 = n6069 & n6436;
  assign n6438 = po30  & n6437;
  assign n6439 = po30  & n6436;
  assign n6440 = ~n6069 & ~n6439;
  assign n6441 = ~n6438 & ~n6440;
  assign n6442 = ~po52  & ~n6425;
  assign n6443 = ~n6433 & n6442;
  assign n6444 = ~n6441 & ~n6443;
  assign n6445 = ~n6435 & ~n6444;
  assign n6446 = po53  & ~n6445;
  assign n6447 = ~n6073 & ~n6081;
  assign n6448 = n6079 & n6447;
  assign n6449 = po30  & n6448;
  assign n6450 = po30  & n6447;
  assign n6451 = ~n6079 & ~n6450;
  assign n6452 = ~n6449 & ~n6451;
  assign n6453 = ~po53  & n6445;
  assign n6454 = ~n6452 & ~n6453;
  assign n6455 = ~n6446 & ~n6454;
  assign n6456 = po54  & ~n6455;
  assign n6457 = ~n6084 & ~n6091;
  assign n6458 = n6090 & n6457;
  assign n6459 = po30  & n6458;
  assign n6460 = po30  & n6457;
  assign n6461 = ~n6090 & ~n6460;
  assign n6462 = ~n6459 & ~n6461;
  assign n6463 = ~po54  & ~n6446;
  assign n6464 = ~n6454 & n6463;
  assign n6465 = ~n6462 & ~n6464;
  assign n6466 = ~n6456 & ~n6465;
  assign n6467 = po55  & ~n6466;
  assign n6468 = ~n6094 & ~n6102;
  assign n6469 = n6100 & n6468;
  assign n6470 = po30  & n6469;
  assign n6471 = po30  & n6468;
  assign n6472 = ~n6100 & ~n6471;
  assign n6473 = ~n6470 & ~n6472;
  assign n6474 = ~po55  & n6466;
  assign n6475 = ~n6473 & ~n6474;
  assign n6476 = ~n6467 & ~n6475;
  assign n6477 = po56  & ~n6476;
  assign n6478 = ~n6105 & ~n6112;
  assign n6479 = n6111 & n6478;
  assign n6480 = po30  & n6479;
  assign n6481 = po30  & n6478;
  assign n6482 = ~n6111 & ~n6481;
  assign n6483 = ~n6480 & ~n6482;
  assign n6484 = ~po56  & ~n6467;
  assign n6485 = ~n6475 & n6484;
  assign n6486 = ~n6483 & ~n6485;
  assign n6487 = ~n6477 & ~n6486;
  assign n6488 = po57  & ~n6487;
  assign n6489 = ~n6115 & ~n6123;
  assign n6490 = n6121 & n6489;
  assign n6491 = po30  & n6490;
  assign n6492 = po30  & n6489;
  assign n6493 = ~n6121 & ~n6492;
  assign n6494 = ~n6491 & ~n6493;
  assign n6495 = ~po57  & n6487;
  assign n6496 = ~n6494 & ~n6495;
  assign n6497 = ~n6488 & ~n6496;
  assign n6498 = po58  & ~n6497;
  assign n6499 = ~n6126 & ~n6133;
  assign n6500 = n6132 & n6499;
  assign n6501 = po30  & n6500;
  assign n6502 = po30  & n6499;
  assign n6503 = ~n6132 & ~n6502;
  assign n6504 = ~n6501 & ~n6503;
  assign n6505 = ~po58  & ~n6488;
  assign n6506 = ~n6496 & n6505;
  assign n6507 = ~n6504 & ~n6506;
  assign n6508 = ~n6498 & ~n6507;
  assign n6509 = po59  & ~n6508;
  assign n6510 = ~n6136 & ~n6144;
  assign n6511 = n6142 & n6510;
  assign n6512 = po30  & n6511;
  assign n6513 = po30  & n6510;
  assign n6514 = ~n6142 & ~n6513;
  assign n6515 = ~n6512 & ~n6514;
  assign n6516 = ~po59  & n6508;
  assign n6517 = ~n6515 & ~n6516;
  assign n6518 = ~n6509 & ~n6517;
  assign n6519 = po60  & ~n6518;
  assign n6520 = ~n6147 & ~n6154;
  assign n6521 = n6153 & n6520;
  assign n6522 = po30  & n6521;
  assign n6523 = po30  & n6520;
  assign n6524 = ~n6153 & ~n6523;
  assign n6525 = ~n6522 & ~n6524;
  assign n6526 = ~po60  & ~n6509;
  assign n6527 = ~n6517 & n6526;
  assign n6528 = ~n6525 & ~n6527;
  assign n6529 = ~n6519 & ~n6528;
  assign n6530 = po61  & ~n6529;
  assign n6531 = ~n6157 & ~n6165;
  assign n6532 = n6163 & n6531;
  assign n6533 = po30  & n6532;
  assign n6534 = po30  & n6531;
  assign n6535 = ~n6163 & ~n6534;
  assign n6536 = ~n6533 & ~n6535;
  assign n6537 = ~po61  & n6529;
  assign n6538 = ~n6536 & ~n6537;
  assign n6539 = ~n6530 & ~n6538;
  assign n6540 = po62  & ~n6539;
  assign n6541 = ~n6168 & ~n6175;
  assign n6542 = n6174 & n6541;
  assign n6543 = po30  & n6542;
  assign n6544 = po30  & n6541;
  assign n6545 = ~n6174 & ~n6544;
  assign n6546 = ~n6543 & ~n6545;
  assign n6547 = ~po62  & ~n6530;
  assign n6548 = ~n6538 & n6547;
  assign n6549 = ~n6546 & ~n6548;
  assign n6550 = ~n6540 & ~n6549;
  assign n6551 = ~n6178 & ~n6186;
  assign n6552 = po30  & n6551;
  assign n6553 = ~n6184 & ~n6552;
  assign n6554 = n6184 & n6552;
  assign n6555 = ~n6553 & ~n6554;
  assign n6556 = ~n6188 & ~n6193;
  assign n6557 = po30  & n6556;
  assign n6558 = ~n6206 & ~n6557;
  assign n6559 = ~n6555 & n6558;
  assign n6560 = ~n6550 & n6559;
  assign n6561 = ~po63  & ~n6560;
  assign n6562 = ~n6193 & po30 ;
  assign n6563 = n6188 & ~n6562;
  assign n6564 = po63  & ~n6556;
  assign n6565 = ~n6563 & n6564;
  assign n6566 = n6193 & ~po30 ;
  assign n6567 = ~n6565 & ~n6566;
  assign n6568 = n6550 & n6555;
  assign n6569 = n6567 & ~n6568;
  assign po29  = n6561 | ~n6569;
  assign n6571 = pi58  & po29 ;
  assign n6572 = ~pi56  & ~pi57 ;
  assign n6573 = ~pi58  & n6572;
  assign n6574 = ~n6571 & ~n6573;
  assign n6575 = po30  & ~n6574;
  assign n6576 = n6205 & ~n6573;
  assign n6577 = ~n6206 & n6576;
  assign n6578 = ~n6199 & n6577;
  assign n6579 = ~n6571 & n6578;
  assign n6580 = ~pi58  & po29 ;
  assign n6581 = pi59  & ~n6580;
  assign n6582 = n6210 & po29 ;
  assign n6583 = ~n6581 & ~n6582;
  assign n6584 = ~n6579 & n6583;
  assign n6585 = ~n6575 & ~n6584;
  assign n6586 = po31  & ~n6585;
  assign n6587 = po30  & n6567;
  assign n6588 = ~n6568 & n6587;
  assign n6589 = ~n6561 & n6588;
  assign n6590 = ~n6582 & ~n6589;
  assign n6591 = pi60  & ~n6590;
  assign n6592 = ~pi60  & n6590;
  assign n6593 = ~n6591 & ~n6592;
  assign n6594 = ~po31  & n6585;
  assign n6595 = ~n6593 & ~n6594;
  assign n6596 = ~n6586 & ~n6595;
  assign n6597 = po32  & ~n6596;
  assign n6598 = ~n6213 & ~n6217;
  assign n6599 = ~n6221 & n6598;
  assign n6600 = po29  & n6599;
  assign n6601 = po29  & n6598;
  assign n6602 = n6221 & ~n6601;
  assign n6603 = ~n6600 & ~n6602;
  assign n6604 = ~po32  & ~n6586;
  assign n6605 = ~n6595 & n6604;
  assign n6606 = ~n6603 & ~n6605;
  assign n6607 = ~n6597 & ~n6606;
  assign n6608 = po33  & ~n6607;
  assign n6609 = ~n6224 & ~n6226;
  assign n6610 = n6233 & n6609;
  assign n6611 = po29  & n6610;
  assign n6612 = po29  & n6609;
  assign n6613 = ~n6233 & ~n6612;
  assign n6614 = ~n6611 & ~n6613;
  assign n6615 = ~po33  & n6607;
  assign n6616 = ~n6614 & ~n6615;
  assign n6617 = ~n6608 & ~n6616;
  assign n6618 = po34  & ~n6617;
  assign n6619 = ~n6236 & ~n6243;
  assign n6620 = n6242 & n6619;
  assign n6621 = po29  & n6620;
  assign n6622 = po29  & n6619;
  assign n6623 = ~n6242 & ~n6622;
  assign n6624 = ~n6621 & ~n6623;
  assign n6625 = ~po34  & ~n6608;
  assign n6626 = ~n6616 & n6625;
  assign n6627 = ~n6624 & ~n6626;
  assign n6628 = ~n6618 & ~n6627;
  assign n6629 = po35  & ~n6628;
  assign n6630 = ~n6246 & ~n6254;
  assign n6631 = n6252 & n6630;
  assign n6632 = po29  & n6631;
  assign n6633 = po29  & n6630;
  assign n6634 = ~n6252 & ~n6633;
  assign n6635 = ~n6632 & ~n6634;
  assign n6636 = ~po35  & n6628;
  assign n6637 = ~n6635 & ~n6636;
  assign n6638 = ~n6629 & ~n6637;
  assign n6639 = po36  & ~n6638;
  assign n6640 = ~po36  & ~n6629;
  assign n6641 = ~n6637 & n6640;
  assign n6642 = ~n6257 & ~n6264;
  assign n6643 = n6263 & n6642;
  assign n6644 = po29  & n6643;
  assign n6645 = po29  & n6642;
  assign n6646 = ~n6263 & ~n6645;
  assign n6647 = ~n6644 & ~n6646;
  assign n6648 = ~n6641 & ~n6647;
  assign n6649 = ~n6639 & ~n6648;
  assign n6650 = po37  & ~n6649;
  assign n6651 = ~n6267 & ~n6275;
  assign n6652 = n6273 & n6651;
  assign n6653 = po29  & n6652;
  assign n6654 = po29  & n6651;
  assign n6655 = ~n6273 & ~n6654;
  assign n6656 = ~n6653 & ~n6655;
  assign n6657 = ~po37  & n6649;
  assign n6658 = ~n6656 & ~n6657;
  assign n6659 = ~n6650 & ~n6658;
  assign n6660 = po38  & ~n6659;
  assign n6661 = ~n6278 & ~n6285;
  assign n6662 = n6284 & n6661;
  assign n6663 = po29  & n6662;
  assign n6664 = po29  & n6661;
  assign n6665 = ~n6284 & ~n6664;
  assign n6666 = ~n6663 & ~n6665;
  assign n6667 = ~po38  & ~n6650;
  assign n6668 = ~n6658 & n6667;
  assign n6669 = ~n6666 & ~n6668;
  assign n6670 = ~n6660 & ~n6669;
  assign n6671 = po39  & ~n6670;
  assign n6672 = ~n6288 & ~n6296;
  assign n6673 = n6294 & n6672;
  assign n6674 = po29  & n6673;
  assign n6675 = po29  & n6672;
  assign n6676 = ~n6294 & ~n6675;
  assign n6677 = ~n6674 & ~n6676;
  assign n6678 = ~po39  & n6670;
  assign n6679 = ~n6677 & ~n6678;
  assign n6680 = ~n6671 & ~n6679;
  assign n6681 = po40  & ~n6680;
  assign n6682 = ~n6299 & ~n6306;
  assign n6683 = n6305 & n6682;
  assign n6684 = po29  & n6683;
  assign n6685 = po29  & n6682;
  assign n6686 = ~n6305 & ~n6685;
  assign n6687 = ~n6684 & ~n6686;
  assign n6688 = ~po40  & ~n6671;
  assign n6689 = ~n6679 & n6688;
  assign n6690 = ~n6687 & ~n6689;
  assign n6691 = ~n6681 & ~n6690;
  assign n6692 = po41  & ~n6691;
  assign n6693 = ~n6309 & ~n6317;
  assign n6694 = n6315 & n6693;
  assign n6695 = po29  & n6694;
  assign n6696 = po29  & n6693;
  assign n6697 = ~n6315 & ~n6696;
  assign n6698 = ~n6695 & ~n6697;
  assign n6699 = ~po41  & n6691;
  assign n6700 = ~n6698 & ~n6699;
  assign n6701 = ~n6692 & ~n6700;
  assign n6702 = po42  & ~n6701;
  assign n6703 = ~n6320 & ~n6327;
  assign n6704 = n6326 & n6703;
  assign n6705 = po29  & n6704;
  assign n6706 = po29  & n6703;
  assign n6707 = ~n6326 & ~n6706;
  assign n6708 = ~n6705 & ~n6707;
  assign n6709 = ~po42  & ~n6692;
  assign n6710 = ~n6700 & n6709;
  assign n6711 = ~n6708 & ~n6710;
  assign n6712 = ~n6702 & ~n6711;
  assign n6713 = po43  & ~n6712;
  assign n6714 = ~n6330 & ~n6338;
  assign n6715 = n6336 & n6714;
  assign n6716 = po29  & n6715;
  assign n6717 = po29  & n6714;
  assign n6718 = ~n6336 & ~n6717;
  assign n6719 = ~n6716 & ~n6718;
  assign n6720 = ~po43  & n6712;
  assign n6721 = ~n6719 & ~n6720;
  assign n6722 = ~n6713 & ~n6721;
  assign n6723 = po44  & ~n6722;
  assign n6724 = ~n6341 & ~n6348;
  assign n6725 = n6347 & n6724;
  assign n6726 = po29  & n6725;
  assign n6727 = po29  & n6724;
  assign n6728 = ~n6347 & ~n6727;
  assign n6729 = ~n6726 & ~n6728;
  assign n6730 = ~po44  & ~n6713;
  assign n6731 = ~n6721 & n6730;
  assign n6732 = ~n6729 & ~n6731;
  assign n6733 = ~n6723 & ~n6732;
  assign n6734 = po45  & ~n6733;
  assign n6735 = ~n6351 & ~n6359;
  assign n6736 = n6357 & n6735;
  assign n6737 = po29  & n6736;
  assign n6738 = po29  & n6735;
  assign n6739 = ~n6357 & ~n6738;
  assign n6740 = ~n6737 & ~n6739;
  assign n6741 = ~po45  & n6733;
  assign n6742 = ~n6740 & ~n6741;
  assign n6743 = ~n6734 & ~n6742;
  assign n6744 = po46  & ~n6743;
  assign n6745 = ~n6362 & ~n6369;
  assign n6746 = n6368 & n6745;
  assign n6747 = po29  & n6746;
  assign n6748 = po29  & n6745;
  assign n6749 = ~n6368 & ~n6748;
  assign n6750 = ~n6747 & ~n6749;
  assign n6751 = ~po46  & ~n6734;
  assign n6752 = ~n6742 & n6751;
  assign n6753 = ~n6750 & ~n6752;
  assign n6754 = ~n6744 & ~n6753;
  assign n6755 = po47  & ~n6754;
  assign n6756 = ~n6372 & ~n6380;
  assign n6757 = n6378 & n6756;
  assign n6758 = po29  & n6757;
  assign n6759 = po29  & n6756;
  assign n6760 = ~n6378 & ~n6759;
  assign n6761 = ~n6758 & ~n6760;
  assign n6762 = ~po47  & n6754;
  assign n6763 = ~n6761 & ~n6762;
  assign n6764 = ~n6755 & ~n6763;
  assign n6765 = po48  & ~n6764;
  assign n6766 = ~n6383 & ~n6390;
  assign n6767 = n6389 & n6766;
  assign n6768 = po29  & n6767;
  assign n6769 = po29  & n6766;
  assign n6770 = ~n6389 & ~n6769;
  assign n6771 = ~n6768 & ~n6770;
  assign n6772 = ~po48  & ~n6755;
  assign n6773 = ~n6763 & n6772;
  assign n6774 = ~n6771 & ~n6773;
  assign n6775 = ~n6765 & ~n6774;
  assign n6776 = po49  & ~n6775;
  assign n6777 = ~n6393 & ~n6401;
  assign n6778 = n6399 & n6777;
  assign n6779 = po29  & n6778;
  assign n6780 = po29  & n6777;
  assign n6781 = ~n6399 & ~n6780;
  assign n6782 = ~n6779 & ~n6781;
  assign n6783 = ~po49  & n6775;
  assign n6784 = ~n6782 & ~n6783;
  assign n6785 = ~n6776 & ~n6784;
  assign n6786 = po50  & ~n6785;
  assign n6787 = ~n6404 & ~n6411;
  assign n6788 = n6410 & n6787;
  assign n6789 = po29  & n6788;
  assign n6790 = po29  & n6787;
  assign n6791 = ~n6410 & ~n6790;
  assign n6792 = ~n6789 & ~n6791;
  assign n6793 = ~po50  & ~n6776;
  assign n6794 = ~n6784 & n6793;
  assign n6795 = ~n6792 & ~n6794;
  assign n6796 = ~n6786 & ~n6795;
  assign n6797 = po51  & ~n6796;
  assign n6798 = ~n6414 & ~n6422;
  assign n6799 = n6420 & n6798;
  assign n6800 = po29  & n6799;
  assign n6801 = po29  & n6798;
  assign n6802 = ~n6420 & ~n6801;
  assign n6803 = ~n6800 & ~n6802;
  assign n6804 = ~po51  & n6796;
  assign n6805 = ~n6803 & ~n6804;
  assign n6806 = ~n6797 & ~n6805;
  assign n6807 = po52  & ~n6806;
  assign n6808 = ~n6425 & ~n6432;
  assign n6809 = n6431 & n6808;
  assign n6810 = po29  & n6809;
  assign n6811 = po29  & n6808;
  assign n6812 = ~n6431 & ~n6811;
  assign n6813 = ~n6810 & ~n6812;
  assign n6814 = ~po52  & ~n6797;
  assign n6815 = ~n6805 & n6814;
  assign n6816 = ~n6813 & ~n6815;
  assign n6817 = ~n6807 & ~n6816;
  assign n6818 = po53  & ~n6817;
  assign n6819 = ~n6435 & ~n6443;
  assign n6820 = n6441 & n6819;
  assign n6821 = po29  & n6820;
  assign n6822 = po29  & n6819;
  assign n6823 = ~n6441 & ~n6822;
  assign n6824 = ~n6821 & ~n6823;
  assign n6825 = ~po53  & n6817;
  assign n6826 = ~n6824 & ~n6825;
  assign n6827 = ~n6818 & ~n6826;
  assign n6828 = po54  & ~n6827;
  assign n6829 = ~n6446 & ~n6453;
  assign n6830 = n6452 & n6829;
  assign n6831 = po29  & n6830;
  assign n6832 = po29  & n6829;
  assign n6833 = ~n6452 & ~n6832;
  assign n6834 = ~n6831 & ~n6833;
  assign n6835 = ~po54  & ~n6818;
  assign n6836 = ~n6826 & n6835;
  assign n6837 = ~n6834 & ~n6836;
  assign n6838 = ~n6828 & ~n6837;
  assign n6839 = po55  & ~n6838;
  assign n6840 = ~n6456 & ~n6464;
  assign n6841 = n6462 & n6840;
  assign n6842 = po29  & n6841;
  assign n6843 = po29  & n6840;
  assign n6844 = ~n6462 & ~n6843;
  assign n6845 = ~n6842 & ~n6844;
  assign n6846 = ~po55  & n6838;
  assign n6847 = ~n6845 & ~n6846;
  assign n6848 = ~n6839 & ~n6847;
  assign n6849 = po56  & ~n6848;
  assign n6850 = ~n6467 & ~n6474;
  assign n6851 = n6473 & n6850;
  assign n6852 = po29  & n6851;
  assign n6853 = po29  & n6850;
  assign n6854 = ~n6473 & ~n6853;
  assign n6855 = ~n6852 & ~n6854;
  assign n6856 = ~po56  & ~n6839;
  assign n6857 = ~n6847 & n6856;
  assign n6858 = ~n6855 & ~n6857;
  assign n6859 = ~n6849 & ~n6858;
  assign n6860 = po57  & ~n6859;
  assign n6861 = ~n6477 & ~n6485;
  assign n6862 = n6483 & n6861;
  assign n6863 = po29  & n6862;
  assign n6864 = po29  & n6861;
  assign n6865 = ~n6483 & ~n6864;
  assign n6866 = ~n6863 & ~n6865;
  assign n6867 = ~po57  & n6859;
  assign n6868 = ~n6866 & ~n6867;
  assign n6869 = ~n6860 & ~n6868;
  assign n6870 = po58  & ~n6869;
  assign n6871 = ~n6488 & ~n6495;
  assign n6872 = n6494 & n6871;
  assign n6873 = po29  & n6872;
  assign n6874 = po29  & n6871;
  assign n6875 = ~n6494 & ~n6874;
  assign n6876 = ~n6873 & ~n6875;
  assign n6877 = ~po58  & ~n6860;
  assign n6878 = ~n6868 & n6877;
  assign n6879 = ~n6876 & ~n6878;
  assign n6880 = ~n6870 & ~n6879;
  assign n6881 = po59  & ~n6880;
  assign n6882 = ~n6498 & ~n6506;
  assign n6883 = n6504 & n6882;
  assign n6884 = po29  & n6883;
  assign n6885 = po29  & n6882;
  assign n6886 = ~n6504 & ~n6885;
  assign n6887 = ~n6884 & ~n6886;
  assign n6888 = ~po59  & n6880;
  assign n6889 = ~n6887 & ~n6888;
  assign n6890 = ~n6881 & ~n6889;
  assign n6891 = po60  & ~n6890;
  assign n6892 = ~n6509 & ~n6516;
  assign n6893 = n6515 & n6892;
  assign n6894 = po29  & n6893;
  assign n6895 = po29  & n6892;
  assign n6896 = ~n6515 & ~n6895;
  assign n6897 = ~n6894 & ~n6896;
  assign n6898 = ~po60  & ~n6881;
  assign n6899 = ~n6889 & n6898;
  assign n6900 = ~n6897 & ~n6899;
  assign n6901 = ~n6891 & ~n6900;
  assign n6902 = po61  & ~n6901;
  assign n6903 = ~n6519 & ~n6527;
  assign n6904 = n6525 & n6903;
  assign n6905 = po29  & n6904;
  assign n6906 = po29  & n6903;
  assign n6907 = ~n6525 & ~n6906;
  assign n6908 = ~n6905 & ~n6907;
  assign n6909 = ~po61  & n6901;
  assign n6910 = ~n6908 & ~n6909;
  assign n6911 = ~n6902 & ~n6910;
  assign n6912 = po62  & ~n6911;
  assign n6913 = ~n6530 & ~n6537;
  assign n6914 = n6536 & n6913;
  assign n6915 = po29  & n6914;
  assign n6916 = po29  & n6913;
  assign n6917 = ~n6536 & ~n6916;
  assign n6918 = ~n6915 & ~n6917;
  assign n6919 = ~po62  & ~n6902;
  assign n6920 = ~n6910 & n6919;
  assign n6921 = ~n6918 & ~n6920;
  assign n6922 = ~n6912 & ~n6921;
  assign n6923 = ~n6540 & ~n6548;
  assign n6924 = po29  & n6923;
  assign n6925 = ~n6546 & ~n6924;
  assign n6926 = n6546 & n6924;
  assign n6927 = ~n6925 & ~n6926;
  assign n6928 = ~n6550 & ~n6555;
  assign n6929 = po29  & n6928;
  assign n6930 = ~n6568 & ~n6929;
  assign n6931 = ~n6927 & n6930;
  assign n6932 = ~n6922 & n6931;
  assign n6933 = ~po63  & ~n6932;
  assign n6934 = ~n6555 & po29 ;
  assign n6935 = n6550 & ~n6934;
  assign n6936 = po63  & ~n6928;
  assign n6937 = ~n6935 & n6936;
  assign n6938 = n6555 & ~po29 ;
  assign n6939 = ~n6937 & ~n6938;
  assign n6940 = n6922 & n6927;
  assign n6941 = n6939 & ~n6940;
  assign po28  = n6933 | ~n6941;
  assign n6943 = pi56  & po28 ;
  assign n6944 = ~pi54  & ~pi55 ;
  assign n6945 = ~pi56  & n6944;
  assign n6946 = ~n6943 & ~n6945;
  assign n6947 = po29  & ~n6946;
  assign n6948 = n6567 & ~n6945;
  assign n6949 = ~n6568 & n6948;
  assign n6950 = ~n6561 & n6949;
  assign n6951 = ~n6943 & n6950;
  assign n6952 = ~pi56  & po28 ;
  assign n6953 = pi57  & ~n6952;
  assign n6954 = n6572 & po28 ;
  assign n6955 = ~n6953 & ~n6954;
  assign n6956 = ~n6951 & n6955;
  assign n6957 = ~n6947 & ~n6956;
  assign n6958 = po30  & ~n6957;
  assign n6959 = ~po30  & ~n6947;
  assign n6960 = ~n6956 & n6959;
  assign n6961 = po29  & n6939;
  assign n6962 = ~n6940 & n6961;
  assign n6963 = ~n6933 & n6962;
  assign n6964 = ~n6954 & ~n6963;
  assign n6965 = pi58  & ~n6964;
  assign n6966 = ~pi58  & n6964;
  assign n6967 = ~n6965 & ~n6966;
  assign n6968 = ~n6960 & ~n6967;
  assign n6969 = ~n6958 & ~n6968;
  assign n6970 = po31  & ~n6969;
  assign n6971 = ~n6575 & ~n6579;
  assign n6972 = ~n6583 & n6971;
  assign n6973 = po28  & n6972;
  assign n6974 = po28  & n6971;
  assign n6975 = n6583 & ~n6974;
  assign n6976 = ~n6973 & ~n6975;
  assign n6977 = ~po31  & n6969;
  assign n6978 = ~n6976 & ~n6977;
  assign n6979 = ~n6970 & ~n6978;
  assign n6980 = po32  & ~n6979;
  assign n6981 = ~n6586 & ~n6594;
  assign n6982 = n6593 & n6981;
  assign n6983 = po28  & n6982;
  assign n6984 = po28  & n6981;
  assign n6985 = ~n6593 & ~n6984;
  assign n6986 = ~n6983 & ~n6985;
  assign n6987 = ~po32  & ~n6970;
  assign n6988 = ~n6978 & n6987;
  assign n6989 = ~n6986 & ~n6988;
  assign n6990 = ~n6980 & ~n6989;
  assign n6991 = po33  & ~n6990;
  assign n6992 = ~n6597 & ~n6605;
  assign n6993 = n6603 & n6992;
  assign n6994 = po28  & n6993;
  assign n6995 = po28  & n6992;
  assign n6996 = ~n6603 & ~n6995;
  assign n6997 = ~n6994 & ~n6996;
  assign n6998 = ~po33  & n6990;
  assign n6999 = ~n6997 & ~n6998;
  assign n7000 = ~n6991 & ~n6999;
  assign n7001 = po34  & ~n7000;
  assign n7002 = ~n6608 & ~n6615;
  assign n7003 = n6614 & n7002;
  assign n7004 = po28  & n7003;
  assign n7005 = po28  & n7002;
  assign n7006 = ~n6614 & ~n7005;
  assign n7007 = ~n7004 & ~n7006;
  assign n7008 = ~po34  & ~n6991;
  assign n7009 = ~n6999 & n7008;
  assign n7010 = ~n7007 & ~n7009;
  assign n7011 = ~n7001 & ~n7010;
  assign n7012 = po35  & ~n7011;
  assign n7013 = ~n6618 & ~n6626;
  assign n7014 = n6624 & n7013;
  assign n7015 = po28  & n7014;
  assign n7016 = po28  & n7013;
  assign n7017 = ~n6624 & ~n7016;
  assign n7018 = ~n7015 & ~n7017;
  assign n7019 = ~po35  & n7011;
  assign n7020 = ~n7018 & ~n7019;
  assign n7021 = ~n7012 & ~n7020;
  assign n7022 = po36  & ~n7021;
  assign n7023 = ~n6629 & ~n6636;
  assign n7024 = n6635 & n7023;
  assign n7025 = po28  & n7024;
  assign n7026 = po28  & n7023;
  assign n7027 = ~n6635 & ~n7026;
  assign n7028 = ~n7025 & ~n7027;
  assign n7029 = ~po36  & ~n7012;
  assign n7030 = ~n7020 & n7029;
  assign n7031 = ~n7028 & ~n7030;
  assign n7032 = ~n7022 & ~n7031;
  assign n7033 = po37  & ~n7032;
  assign n7034 = ~n6639 & ~n6641;
  assign n7035 = n6647 & n7034;
  assign n7036 = po28  & n7035;
  assign n7037 = po28  & n7034;
  assign n7038 = ~n6647 & ~n7037;
  assign n7039 = ~n7036 & ~n7038;
  assign n7040 = ~po37  & n7032;
  assign n7041 = ~n7039 & ~n7040;
  assign n7042 = ~n7033 & ~n7041;
  assign n7043 = po38  & ~n7042;
  assign n7044 = ~n6650 & ~n6657;
  assign n7045 = n6656 & n7044;
  assign n7046 = po28  & n7045;
  assign n7047 = po28  & n7044;
  assign n7048 = ~n6656 & ~n7047;
  assign n7049 = ~n7046 & ~n7048;
  assign n7050 = ~po38  & ~n7033;
  assign n7051 = ~n7041 & n7050;
  assign n7052 = ~n7049 & ~n7051;
  assign n7053 = ~n7043 & ~n7052;
  assign n7054 = po39  & ~n7053;
  assign n7055 = ~n6660 & ~n6668;
  assign n7056 = n6666 & n7055;
  assign n7057 = po28  & n7056;
  assign n7058 = po28  & n7055;
  assign n7059 = ~n6666 & ~n7058;
  assign n7060 = ~n7057 & ~n7059;
  assign n7061 = ~po39  & n7053;
  assign n7062 = ~n7060 & ~n7061;
  assign n7063 = ~n7054 & ~n7062;
  assign n7064 = po40  & ~n7063;
  assign n7065 = ~n6671 & ~n6678;
  assign n7066 = n6677 & n7065;
  assign n7067 = po28  & n7066;
  assign n7068 = po28  & n7065;
  assign n7069 = ~n6677 & ~n7068;
  assign n7070 = ~n7067 & ~n7069;
  assign n7071 = ~po40  & ~n7054;
  assign n7072 = ~n7062 & n7071;
  assign n7073 = ~n7070 & ~n7072;
  assign n7074 = ~n7064 & ~n7073;
  assign n7075 = po41  & ~n7074;
  assign n7076 = ~n6681 & ~n6689;
  assign n7077 = n6687 & n7076;
  assign n7078 = po28  & n7077;
  assign n7079 = po28  & n7076;
  assign n7080 = ~n6687 & ~n7079;
  assign n7081 = ~n7078 & ~n7080;
  assign n7082 = ~po41  & n7074;
  assign n7083 = ~n7081 & ~n7082;
  assign n7084 = ~n7075 & ~n7083;
  assign n7085 = po42  & ~n7084;
  assign n7086 = ~n6692 & ~n6699;
  assign n7087 = n6698 & n7086;
  assign n7088 = po28  & n7087;
  assign n7089 = po28  & n7086;
  assign n7090 = ~n6698 & ~n7089;
  assign n7091 = ~n7088 & ~n7090;
  assign n7092 = ~po42  & ~n7075;
  assign n7093 = ~n7083 & n7092;
  assign n7094 = ~n7091 & ~n7093;
  assign n7095 = ~n7085 & ~n7094;
  assign n7096 = po43  & ~n7095;
  assign n7097 = ~n6702 & ~n6710;
  assign n7098 = n6708 & n7097;
  assign n7099 = po28  & n7098;
  assign n7100 = po28  & n7097;
  assign n7101 = ~n6708 & ~n7100;
  assign n7102 = ~n7099 & ~n7101;
  assign n7103 = ~po43  & n7095;
  assign n7104 = ~n7102 & ~n7103;
  assign n7105 = ~n7096 & ~n7104;
  assign n7106 = po44  & ~n7105;
  assign n7107 = ~n6713 & ~n6720;
  assign n7108 = n6719 & n7107;
  assign n7109 = po28  & n7108;
  assign n7110 = po28  & n7107;
  assign n7111 = ~n6719 & ~n7110;
  assign n7112 = ~n7109 & ~n7111;
  assign n7113 = ~po44  & ~n7096;
  assign n7114 = ~n7104 & n7113;
  assign n7115 = ~n7112 & ~n7114;
  assign n7116 = ~n7106 & ~n7115;
  assign n7117 = po45  & ~n7116;
  assign n7118 = ~n6723 & ~n6731;
  assign n7119 = n6729 & n7118;
  assign n7120 = po28  & n7119;
  assign n7121 = po28  & n7118;
  assign n7122 = ~n6729 & ~n7121;
  assign n7123 = ~n7120 & ~n7122;
  assign n7124 = ~po45  & n7116;
  assign n7125 = ~n7123 & ~n7124;
  assign n7126 = ~n7117 & ~n7125;
  assign n7127 = po46  & ~n7126;
  assign n7128 = ~n6734 & ~n6741;
  assign n7129 = n6740 & n7128;
  assign n7130 = po28  & n7129;
  assign n7131 = po28  & n7128;
  assign n7132 = ~n6740 & ~n7131;
  assign n7133 = ~n7130 & ~n7132;
  assign n7134 = ~po46  & ~n7117;
  assign n7135 = ~n7125 & n7134;
  assign n7136 = ~n7133 & ~n7135;
  assign n7137 = ~n7127 & ~n7136;
  assign n7138 = po47  & ~n7137;
  assign n7139 = ~n6744 & ~n6752;
  assign n7140 = n6750 & n7139;
  assign n7141 = po28  & n7140;
  assign n7142 = po28  & n7139;
  assign n7143 = ~n6750 & ~n7142;
  assign n7144 = ~n7141 & ~n7143;
  assign n7145 = ~po47  & n7137;
  assign n7146 = ~n7144 & ~n7145;
  assign n7147 = ~n7138 & ~n7146;
  assign n7148 = po48  & ~n7147;
  assign n7149 = ~n6755 & ~n6762;
  assign n7150 = n6761 & n7149;
  assign n7151 = po28  & n7150;
  assign n7152 = po28  & n7149;
  assign n7153 = ~n6761 & ~n7152;
  assign n7154 = ~n7151 & ~n7153;
  assign n7155 = ~po48  & ~n7138;
  assign n7156 = ~n7146 & n7155;
  assign n7157 = ~n7154 & ~n7156;
  assign n7158 = ~n7148 & ~n7157;
  assign n7159 = po49  & ~n7158;
  assign n7160 = ~n6765 & ~n6773;
  assign n7161 = n6771 & n7160;
  assign n7162 = po28  & n7161;
  assign n7163 = po28  & n7160;
  assign n7164 = ~n6771 & ~n7163;
  assign n7165 = ~n7162 & ~n7164;
  assign n7166 = ~po49  & n7158;
  assign n7167 = ~n7165 & ~n7166;
  assign n7168 = ~n7159 & ~n7167;
  assign n7169 = po50  & ~n7168;
  assign n7170 = ~n6776 & ~n6783;
  assign n7171 = n6782 & n7170;
  assign n7172 = po28  & n7171;
  assign n7173 = po28  & n7170;
  assign n7174 = ~n6782 & ~n7173;
  assign n7175 = ~n7172 & ~n7174;
  assign n7176 = ~po50  & ~n7159;
  assign n7177 = ~n7167 & n7176;
  assign n7178 = ~n7175 & ~n7177;
  assign n7179 = ~n7169 & ~n7178;
  assign n7180 = po51  & ~n7179;
  assign n7181 = ~n6786 & ~n6794;
  assign n7182 = n6792 & n7181;
  assign n7183 = po28  & n7182;
  assign n7184 = po28  & n7181;
  assign n7185 = ~n6792 & ~n7184;
  assign n7186 = ~n7183 & ~n7185;
  assign n7187 = ~po51  & n7179;
  assign n7188 = ~n7186 & ~n7187;
  assign n7189 = ~n7180 & ~n7188;
  assign n7190 = po52  & ~n7189;
  assign n7191 = ~n6797 & ~n6804;
  assign n7192 = n6803 & n7191;
  assign n7193 = po28  & n7192;
  assign n7194 = po28  & n7191;
  assign n7195 = ~n6803 & ~n7194;
  assign n7196 = ~n7193 & ~n7195;
  assign n7197 = ~po52  & ~n7180;
  assign n7198 = ~n7188 & n7197;
  assign n7199 = ~n7196 & ~n7198;
  assign n7200 = ~n7190 & ~n7199;
  assign n7201 = po53  & ~n7200;
  assign n7202 = ~n6807 & ~n6815;
  assign n7203 = n6813 & n7202;
  assign n7204 = po28  & n7203;
  assign n7205 = po28  & n7202;
  assign n7206 = ~n6813 & ~n7205;
  assign n7207 = ~n7204 & ~n7206;
  assign n7208 = ~po53  & n7200;
  assign n7209 = ~n7207 & ~n7208;
  assign n7210 = ~n7201 & ~n7209;
  assign n7211 = po54  & ~n7210;
  assign n7212 = ~n6818 & ~n6825;
  assign n7213 = n6824 & n7212;
  assign n7214 = po28  & n7213;
  assign n7215 = po28  & n7212;
  assign n7216 = ~n6824 & ~n7215;
  assign n7217 = ~n7214 & ~n7216;
  assign n7218 = ~po54  & ~n7201;
  assign n7219 = ~n7209 & n7218;
  assign n7220 = ~n7217 & ~n7219;
  assign n7221 = ~n7211 & ~n7220;
  assign n7222 = po55  & ~n7221;
  assign n7223 = ~n6828 & ~n6836;
  assign n7224 = n6834 & n7223;
  assign n7225 = po28  & n7224;
  assign n7226 = po28  & n7223;
  assign n7227 = ~n6834 & ~n7226;
  assign n7228 = ~n7225 & ~n7227;
  assign n7229 = ~po55  & n7221;
  assign n7230 = ~n7228 & ~n7229;
  assign n7231 = ~n7222 & ~n7230;
  assign n7232 = po56  & ~n7231;
  assign n7233 = ~n6839 & ~n6846;
  assign n7234 = n6845 & n7233;
  assign n7235 = po28  & n7234;
  assign n7236 = po28  & n7233;
  assign n7237 = ~n6845 & ~n7236;
  assign n7238 = ~n7235 & ~n7237;
  assign n7239 = ~po56  & ~n7222;
  assign n7240 = ~n7230 & n7239;
  assign n7241 = ~n7238 & ~n7240;
  assign n7242 = ~n7232 & ~n7241;
  assign n7243 = po57  & ~n7242;
  assign n7244 = ~n6849 & ~n6857;
  assign n7245 = n6855 & n7244;
  assign n7246 = po28  & n7245;
  assign n7247 = po28  & n7244;
  assign n7248 = ~n6855 & ~n7247;
  assign n7249 = ~n7246 & ~n7248;
  assign n7250 = ~po57  & n7242;
  assign n7251 = ~n7249 & ~n7250;
  assign n7252 = ~n7243 & ~n7251;
  assign n7253 = po58  & ~n7252;
  assign n7254 = ~n6860 & ~n6867;
  assign n7255 = n6866 & n7254;
  assign n7256 = po28  & n7255;
  assign n7257 = po28  & n7254;
  assign n7258 = ~n6866 & ~n7257;
  assign n7259 = ~n7256 & ~n7258;
  assign n7260 = ~po58  & ~n7243;
  assign n7261 = ~n7251 & n7260;
  assign n7262 = ~n7259 & ~n7261;
  assign n7263 = ~n7253 & ~n7262;
  assign n7264 = po59  & ~n7263;
  assign n7265 = ~n6870 & ~n6878;
  assign n7266 = n6876 & n7265;
  assign n7267 = po28  & n7266;
  assign n7268 = po28  & n7265;
  assign n7269 = ~n6876 & ~n7268;
  assign n7270 = ~n7267 & ~n7269;
  assign n7271 = ~po59  & n7263;
  assign n7272 = ~n7270 & ~n7271;
  assign n7273 = ~n7264 & ~n7272;
  assign n7274 = po60  & ~n7273;
  assign n7275 = ~n6881 & ~n6888;
  assign n7276 = n6887 & n7275;
  assign n7277 = po28  & n7276;
  assign n7278 = po28  & n7275;
  assign n7279 = ~n6887 & ~n7278;
  assign n7280 = ~n7277 & ~n7279;
  assign n7281 = ~po60  & ~n7264;
  assign n7282 = ~n7272 & n7281;
  assign n7283 = ~n7280 & ~n7282;
  assign n7284 = ~n7274 & ~n7283;
  assign n7285 = po61  & ~n7284;
  assign n7286 = ~n6891 & ~n6899;
  assign n7287 = n6897 & n7286;
  assign n7288 = po28  & n7287;
  assign n7289 = po28  & n7286;
  assign n7290 = ~n6897 & ~n7289;
  assign n7291 = ~n7288 & ~n7290;
  assign n7292 = ~po61  & n7284;
  assign n7293 = ~n7291 & ~n7292;
  assign n7294 = ~n7285 & ~n7293;
  assign n7295 = po62  & ~n7294;
  assign n7296 = ~n6902 & ~n6909;
  assign n7297 = n6908 & n7296;
  assign n7298 = po28  & n7297;
  assign n7299 = po28  & n7296;
  assign n7300 = ~n6908 & ~n7299;
  assign n7301 = ~n7298 & ~n7300;
  assign n7302 = ~po62  & ~n7285;
  assign n7303 = ~n7293 & n7302;
  assign n7304 = ~n7301 & ~n7303;
  assign n7305 = ~n7295 & ~n7304;
  assign n7306 = ~n6912 & ~n6920;
  assign n7307 = po28  & n7306;
  assign n7308 = ~n6918 & ~n7307;
  assign n7309 = n6918 & n7307;
  assign n7310 = ~n7308 & ~n7309;
  assign n7311 = ~n6922 & ~n6927;
  assign n7312 = po28  & n7311;
  assign n7313 = ~n6940 & ~n7312;
  assign n7314 = ~n7310 & n7313;
  assign n7315 = ~n7305 & n7314;
  assign n7316 = ~po63  & ~n7315;
  assign n7317 = ~n6927 & po28 ;
  assign n7318 = n6922 & ~n7317;
  assign n7319 = po63  & ~n7311;
  assign n7320 = ~n7318 & n7319;
  assign n7321 = n6927 & ~po28 ;
  assign n7322 = ~n7320 & ~n7321;
  assign n7323 = n7305 & n7310;
  assign n7324 = n7322 & ~n7323;
  assign po27  = n7316 | ~n7324;
  assign n7326 = pi54  & po27 ;
  assign n7327 = ~pi52  & ~pi53 ;
  assign n7328 = ~pi54  & n7327;
  assign n7329 = ~n7326 & ~n7328;
  assign n7330 = po28  & ~n7329;
  assign n7331 = n6939 & ~n7328;
  assign n7332 = ~n6940 & n7331;
  assign n7333 = ~n6933 & n7332;
  assign n7334 = ~n7326 & n7333;
  assign n7335 = ~pi54  & po27 ;
  assign n7336 = pi55  & ~n7335;
  assign n7337 = n6944 & po27 ;
  assign n7338 = ~n7336 & ~n7337;
  assign n7339 = ~n7334 & n7338;
  assign n7340 = ~n7330 & ~n7339;
  assign n7341 = po29  & ~n7340;
  assign n7342 = po28  & n7322;
  assign n7343 = ~n7323 & n7342;
  assign n7344 = ~n7316 & n7343;
  assign n7345 = ~n7337 & ~n7344;
  assign n7346 = pi56  & ~n7345;
  assign n7347 = ~pi56  & n7345;
  assign n7348 = ~n7346 & ~n7347;
  assign n7349 = ~po29  & n7340;
  assign n7350 = ~n7348 & ~n7349;
  assign n7351 = ~n7341 & ~n7350;
  assign n7352 = po30  & ~n7351;
  assign n7353 = ~n6947 & ~n6951;
  assign n7354 = ~n6955 & n7353;
  assign n7355 = po27  & n7354;
  assign n7356 = po27  & n7353;
  assign n7357 = n6955 & ~n7356;
  assign n7358 = ~n7355 & ~n7357;
  assign n7359 = ~po30  & ~n7341;
  assign n7360 = ~n7350 & n7359;
  assign n7361 = ~n7358 & ~n7360;
  assign n7362 = ~n7352 & ~n7361;
  assign n7363 = po31  & ~n7362;
  assign n7364 = ~n6958 & ~n6960;
  assign n7365 = n6967 & n7364;
  assign n7366 = po27  & n7365;
  assign n7367 = po27  & n7364;
  assign n7368 = ~n6967 & ~n7367;
  assign n7369 = ~n7366 & ~n7368;
  assign n7370 = ~po31  & n7362;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = ~n7363 & ~n7371;
  assign n7373 = po32  & ~n7372;
  assign n7374 = ~n6970 & ~n6977;
  assign n7375 = n6976 & n7374;
  assign n7376 = po27  & n7375;
  assign n7377 = po27  & n7374;
  assign n7378 = ~n6976 & ~n7377;
  assign n7379 = ~n7376 & ~n7378;
  assign n7380 = ~po32  & ~n7363;
  assign n7381 = ~n7371 & n7380;
  assign n7382 = ~n7379 & ~n7381;
  assign n7383 = ~n7373 & ~n7382;
  assign n7384 = po33  & ~n7383;
  assign n7385 = ~n6980 & ~n6988;
  assign n7386 = n6986 & n7385;
  assign n7387 = po27  & n7386;
  assign n7388 = po27  & n7385;
  assign n7389 = ~n6986 & ~n7388;
  assign n7390 = ~n7387 & ~n7389;
  assign n7391 = ~po33  & n7383;
  assign n7392 = ~n7390 & ~n7391;
  assign n7393 = ~n7384 & ~n7392;
  assign n7394 = po34  & ~n7393;
  assign n7395 = ~n6991 & ~n6998;
  assign n7396 = n6997 & n7395;
  assign n7397 = po27  & n7396;
  assign n7398 = po27  & n7395;
  assign n7399 = ~n6997 & ~n7398;
  assign n7400 = ~n7397 & ~n7399;
  assign n7401 = ~po34  & ~n7384;
  assign n7402 = ~n7392 & n7401;
  assign n7403 = ~n7400 & ~n7402;
  assign n7404 = ~n7394 & ~n7403;
  assign n7405 = po35  & ~n7404;
  assign n7406 = ~n7001 & ~n7009;
  assign n7407 = n7007 & n7406;
  assign n7408 = po27  & n7407;
  assign n7409 = po27  & n7406;
  assign n7410 = ~n7007 & ~n7409;
  assign n7411 = ~n7408 & ~n7410;
  assign n7412 = ~po35  & n7404;
  assign n7413 = ~n7411 & ~n7412;
  assign n7414 = ~n7405 & ~n7413;
  assign n7415 = po36  & ~n7414;
  assign n7416 = ~n7012 & ~n7019;
  assign n7417 = n7018 & n7416;
  assign n7418 = po27  & n7417;
  assign n7419 = po27  & n7416;
  assign n7420 = ~n7018 & ~n7419;
  assign n7421 = ~n7418 & ~n7420;
  assign n7422 = ~po36  & ~n7405;
  assign n7423 = ~n7413 & n7422;
  assign n7424 = ~n7421 & ~n7423;
  assign n7425 = ~n7415 & ~n7424;
  assign n7426 = po37  & ~n7425;
  assign n7427 = ~n7022 & ~n7030;
  assign n7428 = n7028 & n7427;
  assign n7429 = po27  & n7428;
  assign n7430 = po27  & n7427;
  assign n7431 = ~n7028 & ~n7430;
  assign n7432 = ~n7429 & ~n7431;
  assign n7433 = ~po37  & n7425;
  assign n7434 = ~n7432 & ~n7433;
  assign n7435 = ~n7426 & ~n7434;
  assign n7436 = po38  & ~n7435;
  assign n7437 = ~po38  & ~n7426;
  assign n7438 = ~n7434 & n7437;
  assign n7439 = ~n7033 & ~n7040;
  assign n7440 = n7039 & n7439;
  assign n7441 = po27  & n7440;
  assign n7442 = po27  & n7439;
  assign n7443 = ~n7039 & ~n7442;
  assign n7444 = ~n7441 & ~n7443;
  assign n7445 = ~n7438 & ~n7444;
  assign n7446 = ~n7436 & ~n7445;
  assign n7447 = po39  & ~n7446;
  assign n7448 = ~n7043 & ~n7051;
  assign n7449 = n7049 & n7448;
  assign n7450 = po27  & n7449;
  assign n7451 = po27  & n7448;
  assign n7452 = ~n7049 & ~n7451;
  assign n7453 = ~n7450 & ~n7452;
  assign n7454 = ~po39  & n7446;
  assign n7455 = ~n7453 & ~n7454;
  assign n7456 = ~n7447 & ~n7455;
  assign n7457 = po40  & ~n7456;
  assign n7458 = ~n7054 & ~n7061;
  assign n7459 = n7060 & n7458;
  assign n7460 = po27  & n7459;
  assign n7461 = po27  & n7458;
  assign n7462 = ~n7060 & ~n7461;
  assign n7463 = ~n7460 & ~n7462;
  assign n7464 = ~po40  & ~n7447;
  assign n7465 = ~n7455 & n7464;
  assign n7466 = ~n7463 & ~n7465;
  assign n7467 = ~n7457 & ~n7466;
  assign n7468 = po41  & ~n7467;
  assign n7469 = ~n7064 & ~n7072;
  assign n7470 = n7070 & n7469;
  assign n7471 = po27  & n7470;
  assign n7472 = po27  & n7469;
  assign n7473 = ~n7070 & ~n7472;
  assign n7474 = ~n7471 & ~n7473;
  assign n7475 = ~po41  & n7467;
  assign n7476 = ~n7474 & ~n7475;
  assign n7477 = ~n7468 & ~n7476;
  assign n7478 = po42  & ~n7477;
  assign n7479 = ~n7075 & ~n7082;
  assign n7480 = n7081 & n7479;
  assign n7481 = po27  & n7480;
  assign n7482 = po27  & n7479;
  assign n7483 = ~n7081 & ~n7482;
  assign n7484 = ~n7481 & ~n7483;
  assign n7485 = ~po42  & ~n7468;
  assign n7486 = ~n7476 & n7485;
  assign n7487 = ~n7484 & ~n7486;
  assign n7488 = ~n7478 & ~n7487;
  assign n7489 = po43  & ~n7488;
  assign n7490 = ~n7085 & ~n7093;
  assign n7491 = n7091 & n7490;
  assign n7492 = po27  & n7491;
  assign n7493 = po27  & n7490;
  assign n7494 = ~n7091 & ~n7493;
  assign n7495 = ~n7492 & ~n7494;
  assign n7496 = ~po43  & n7488;
  assign n7497 = ~n7495 & ~n7496;
  assign n7498 = ~n7489 & ~n7497;
  assign n7499 = po44  & ~n7498;
  assign n7500 = ~n7096 & ~n7103;
  assign n7501 = n7102 & n7500;
  assign n7502 = po27  & n7501;
  assign n7503 = po27  & n7500;
  assign n7504 = ~n7102 & ~n7503;
  assign n7505 = ~n7502 & ~n7504;
  assign n7506 = ~po44  & ~n7489;
  assign n7507 = ~n7497 & n7506;
  assign n7508 = ~n7505 & ~n7507;
  assign n7509 = ~n7499 & ~n7508;
  assign n7510 = po45  & ~n7509;
  assign n7511 = ~n7106 & ~n7114;
  assign n7512 = n7112 & n7511;
  assign n7513 = po27  & n7512;
  assign n7514 = po27  & n7511;
  assign n7515 = ~n7112 & ~n7514;
  assign n7516 = ~n7513 & ~n7515;
  assign n7517 = ~po45  & n7509;
  assign n7518 = ~n7516 & ~n7517;
  assign n7519 = ~n7510 & ~n7518;
  assign n7520 = po46  & ~n7519;
  assign n7521 = ~n7117 & ~n7124;
  assign n7522 = n7123 & n7521;
  assign n7523 = po27  & n7522;
  assign n7524 = po27  & n7521;
  assign n7525 = ~n7123 & ~n7524;
  assign n7526 = ~n7523 & ~n7525;
  assign n7527 = ~po46  & ~n7510;
  assign n7528 = ~n7518 & n7527;
  assign n7529 = ~n7526 & ~n7528;
  assign n7530 = ~n7520 & ~n7529;
  assign n7531 = po47  & ~n7530;
  assign n7532 = ~n7127 & ~n7135;
  assign n7533 = n7133 & n7532;
  assign n7534 = po27  & n7533;
  assign n7535 = po27  & n7532;
  assign n7536 = ~n7133 & ~n7535;
  assign n7537 = ~n7534 & ~n7536;
  assign n7538 = ~po47  & n7530;
  assign n7539 = ~n7537 & ~n7538;
  assign n7540 = ~n7531 & ~n7539;
  assign n7541 = po48  & ~n7540;
  assign n7542 = ~n7138 & ~n7145;
  assign n7543 = n7144 & n7542;
  assign n7544 = po27  & n7543;
  assign n7545 = po27  & n7542;
  assign n7546 = ~n7144 & ~n7545;
  assign n7547 = ~n7544 & ~n7546;
  assign n7548 = ~po48  & ~n7531;
  assign n7549 = ~n7539 & n7548;
  assign n7550 = ~n7547 & ~n7549;
  assign n7551 = ~n7541 & ~n7550;
  assign n7552 = po49  & ~n7551;
  assign n7553 = ~n7148 & ~n7156;
  assign n7554 = n7154 & n7553;
  assign n7555 = po27  & n7554;
  assign n7556 = po27  & n7553;
  assign n7557 = ~n7154 & ~n7556;
  assign n7558 = ~n7555 & ~n7557;
  assign n7559 = ~po49  & n7551;
  assign n7560 = ~n7558 & ~n7559;
  assign n7561 = ~n7552 & ~n7560;
  assign n7562 = po50  & ~n7561;
  assign n7563 = ~n7159 & ~n7166;
  assign n7564 = n7165 & n7563;
  assign n7565 = po27  & n7564;
  assign n7566 = po27  & n7563;
  assign n7567 = ~n7165 & ~n7566;
  assign n7568 = ~n7565 & ~n7567;
  assign n7569 = ~po50  & ~n7552;
  assign n7570 = ~n7560 & n7569;
  assign n7571 = ~n7568 & ~n7570;
  assign n7572 = ~n7562 & ~n7571;
  assign n7573 = po51  & ~n7572;
  assign n7574 = ~n7169 & ~n7177;
  assign n7575 = n7175 & n7574;
  assign n7576 = po27  & n7575;
  assign n7577 = po27  & n7574;
  assign n7578 = ~n7175 & ~n7577;
  assign n7579 = ~n7576 & ~n7578;
  assign n7580 = ~po51  & n7572;
  assign n7581 = ~n7579 & ~n7580;
  assign n7582 = ~n7573 & ~n7581;
  assign n7583 = po52  & ~n7582;
  assign n7584 = ~n7180 & ~n7187;
  assign n7585 = n7186 & n7584;
  assign n7586 = po27  & n7585;
  assign n7587 = po27  & n7584;
  assign n7588 = ~n7186 & ~n7587;
  assign n7589 = ~n7586 & ~n7588;
  assign n7590 = ~po52  & ~n7573;
  assign n7591 = ~n7581 & n7590;
  assign n7592 = ~n7589 & ~n7591;
  assign n7593 = ~n7583 & ~n7592;
  assign n7594 = po53  & ~n7593;
  assign n7595 = ~n7190 & ~n7198;
  assign n7596 = n7196 & n7595;
  assign n7597 = po27  & n7596;
  assign n7598 = po27  & n7595;
  assign n7599 = ~n7196 & ~n7598;
  assign n7600 = ~n7597 & ~n7599;
  assign n7601 = ~po53  & n7593;
  assign n7602 = ~n7600 & ~n7601;
  assign n7603 = ~n7594 & ~n7602;
  assign n7604 = po54  & ~n7603;
  assign n7605 = ~n7201 & ~n7208;
  assign n7606 = n7207 & n7605;
  assign n7607 = po27  & n7606;
  assign n7608 = po27  & n7605;
  assign n7609 = ~n7207 & ~n7608;
  assign n7610 = ~n7607 & ~n7609;
  assign n7611 = ~po54  & ~n7594;
  assign n7612 = ~n7602 & n7611;
  assign n7613 = ~n7610 & ~n7612;
  assign n7614 = ~n7604 & ~n7613;
  assign n7615 = po55  & ~n7614;
  assign n7616 = ~n7211 & ~n7219;
  assign n7617 = n7217 & n7616;
  assign n7618 = po27  & n7617;
  assign n7619 = po27  & n7616;
  assign n7620 = ~n7217 & ~n7619;
  assign n7621 = ~n7618 & ~n7620;
  assign n7622 = ~po55  & n7614;
  assign n7623 = ~n7621 & ~n7622;
  assign n7624 = ~n7615 & ~n7623;
  assign n7625 = po56  & ~n7624;
  assign n7626 = ~n7222 & ~n7229;
  assign n7627 = n7228 & n7626;
  assign n7628 = po27  & n7627;
  assign n7629 = po27  & n7626;
  assign n7630 = ~n7228 & ~n7629;
  assign n7631 = ~n7628 & ~n7630;
  assign n7632 = ~po56  & ~n7615;
  assign n7633 = ~n7623 & n7632;
  assign n7634 = ~n7631 & ~n7633;
  assign n7635 = ~n7625 & ~n7634;
  assign n7636 = po57  & ~n7635;
  assign n7637 = ~n7232 & ~n7240;
  assign n7638 = n7238 & n7637;
  assign n7639 = po27  & n7638;
  assign n7640 = po27  & n7637;
  assign n7641 = ~n7238 & ~n7640;
  assign n7642 = ~n7639 & ~n7641;
  assign n7643 = ~po57  & n7635;
  assign n7644 = ~n7642 & ~n7643;
  assign n7645 = ~n7636 & ~n7644;
  assign n7646 = po58  & ~n7645;
  assign n7647 = ~n7243 & ~n7250;
  assign n7648 = n7249 & n7647;
  assign n7649 = po27  & n7648;
  assign n7650 = po27  & n7647;
  assign n7651 = ~n7249 & ~n7650;
  assign n7652 = ~n7649 & ~n7651;
  assign n7653 = ~po58  & ~n7636;
  assign n7654 = ~n7644 & n7653;
  assign n7655 = ~n7652 & ~n7654;
  assign n7656 = ~n7646 & ~n7655;
  assign n7657 = po59  & ~n7656;
  assign n7658 = ~n7253 & ~n7261;
  assign n7659 = n7259 & n7658;
  assign n7660 = po27  & n7659;
  assign n7661 = po27  & n7658;
  assign n7662 = ~n7259 & ~n7661;
  assign n7663 = ~n7660 & ~n7662;
  assign n7664 = ~po59  & n7656;
  assign n7665 = ~n7663 & ~n7664;
  assign n7666 = ~n7657 & ~n7665;
  assign n7667 = po60  & ~n7666;
  assign n7668 = ~n7264 & ~n7271;
  assign n7669 = n7270 & n7668;
  assign n7670 = po27  & n7669;
  assign n7671 = po27  & n7668;
  assign n7672 = ~n7270 & ~n7671;
  assign n7673 = ~n7670 & ~n7672;
  assign n7674 = ~po60  & ~n7657;
  assign n7675 = ~n7665 & n7674;
  assign n7676 = ~n7673 & ~n7675;
  assign n7677 = ~n7667 & ~n7676;
  assign n7678 = po61  & ~n7677;
  assign n7679 = ~n7274 & ~n7282;
  assign n7680 = n7280 & n7679;
  assign n7681 = po27  & n7680;
  assign n7682 = po27  & n7679;
  assign n7683 = ~n7280 & ~n7682;
  assign n7684 = ~n7681 & ~n7683;
  assign n7685 = ~po61  & n7677;
  assign n7686 = ~n7684 & ~n7685;
  assign n7687 = ~n7678 & ~n7686;
  assign n7688 = po62  & ~n7687;
  assign n7689 = ~n7285 & ~n7292;
  assign n7690 = n7291 & n7689;
  assign n7691 = po27  & n7690;
  assign n7692 = po27  & n7689;
  assign n7693 = ~n7291 & ~n7692;
  assign n7694 = ~n7691 & ~n7693;
  assign n7695 = ~po62  & ~n7678;
  assign n7696 = ~n7686 & n7695;
  assign n7697 = ~n7694 & ~n7696;
  assign n7698 = ~n7688 & ~n7697;
  assign n7699 = ~n7295 & ~n7303;
  assign n7700 = po27  & n7699;
  assign n7701 = ~n7301 & ~n7700;
  assign n7702 = n7301 & n7700;
  assign n7703 = ~n7701 & ~n7702;
  assign n7704 = ~n7305 & ~n7310;
  assign n7705 = po27  & n7704;
  assign n7706 = ~n7323 & ~n7705;
  assign n7707 = ~n7703 & n7706;
  assign n7708 = ~n7698 & n7707;
  assign n7709 = ~po63  & ~n7708;
  assign n7710 = ~n7310 & po27 ;
  assign n7711 = n7305 & ~n7710;
  assign n7712 = po63  & ~n7704;
  assign n7713 = ~n7711 & n7712;
  assign n7714 = n7310 & ~po27 ;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = n7698 & n7703;
  assign n7717 = n7715 & ~n7716;
  assign po26  = n7709 | ~n7717;
  assign n7719 = pi52  & po26 ;
  assign n7720 = ~pi50  & ~pi51 ;
  assign n7721 = ~pi52  & n7720;
  assign n7722 = ~n7719 & ~n7721;
  assign n7723 = po27  & ~n7722;
  assign n7724 = n7322 & ~n7721;
  assign n7725 = ~n7323 & n7724;
  assign n7726 = ~n7316 & n7725;
  assign n7727 = ~n7719 & n7726;
  assign n7728 = ~pi52  & po26 ;
  assign n7729 = pi53  & ~n7728;
  assign n7730 = n7327 & po26 ;
  assign n7731 = ~n7729 & ~n7730;
  assign n7732 = ~n7727 & n7731;
  assign n7733 = ~n7723 & ~n7732;
  assign n7734 = po28  & ~n7733;
  assign n7735 = ~po28  & ~n7723;
  assign n7736 = ~n7732 & n7735;
  assign n7737 = po27  & n7715;
  assign n7738 = ~n7716 & n7737;
  assign n7739 = ~n7709 & n7738;
  assign n7740 = ~n7730 & ~n7739;
  assign n7741 = pi54  & ~n7740;
  assign n7742 = ~pi54  & n7740;
  assign n7743 = ~n7741 & ~n7742;
  assign n7744 = ~n7736 & ~n7743;
  assign n7745 = ~n7734 & ~n7744;
  assign n7746 = po29  & ~n7745;
  assign n7747 = ~n7330 & ~n7334;
  assign n7748 = ~n7338 & n7747;
  assign n7749 = po26  & n7748;
  assign n7750 = po26  & n7747;
  assign n7751 = n7338 & ~n7750;
  assign n7752 = ~n7749 & ~n7751;
  assign n7753 = ~po29  & n7745;
  assign n7754 = ~n7752 & ~n7753;
  assign n7755 = ~n7746 & ~n7754;
  assign n7756 = po30  & ~n7755;
  assign n7757 = ~n7341 & ~n7349;
  assign n7758 = n7348 & n7757;
  assign n7759 = po26  & n7758;
  assign n7760 = po26  & n7757;
  assign n7761 = ~n7348 & ~n7760;
  assign n7762 = ~n7759 & ~n7761;
  assign n7763 = ~po30  & ~n7746;
  assign n7764 = ~n7754 & n7763;
  assign n7765 = ~n7762 & ~n7764;
  assign n7766 = ~n7756 & ~n7765;
  assign n7767 = po31  & ~n7766;
  assign n7768 = ~n7352 & ~n7360;
  assign n7769 = n7358 & n7768;
  assign n7770 = po26  & n7769;
  assign n7771 = po26  & n7768;
  assign n7772 = ~n7358 & ~n7771;
  assign n7773 = ~n7770 & ~n7772;
  assign n7774 = ~po31  & n7766;
  assign n7775 = ~n7773 & ~n7774;
  assign n7776 = ~n7767 & ~n7775;
  assign n7777 = po32  & ~n7776;
  assign n7778 = ~n7363 & ~n7370;
  assign n7779 = n7369 & n7778;
  assign n7780 = po26  & n7779;
  assign n7781 = po26  & n7778;
  assign n7782 = ~n7369 & ~n7781;
  assign n7783 = ~n7780 & ~n7782;
  assign n7784 = ~po32  & ~n7767;
  assign n7785 = ~n7775 & n7784;
  assign n7786 = ~n7783 & ~n7785;
  assign n7787 = ~n7777 & ~n7786;
  assign n7788 = po33  & ~n7787;
  assign n7789 = ~n7373 & ~n7381;
  assign n7790 = n7379 & n7789;
  assign n7791 = po26  & n7790;
  assign n7792 = po26  & n7789;
  assign n7793 = ~n7379 & ~n7792;
  assign n7794 = ~n7791 & ~n7793;
  assign n7795 = ~po33  & n7787;
  assign n7796 = ~n7794 & ~n7795;
  assign n7797 = ~n7788 & ~n7796;
  assign n7798 = po34  & ~n7797;
  assign n7799 = ~n7384 & ~n7391;
  assign n7800 = n7390 & n7799;
  assign n7801 = po26  & n7800;
  assign n7802 = po26  & n7799;
  assign n7803 = ~n7390 & ~n7802;
  assign n7804 = ~n7801 & ~n7803;
  assign n7805 = ~po34  & ~n7788;
  assign n7806 = ~n7796 & n7805;
  assign n7807 = ~n7804 & ~n7806;
  assign n7808 = ~n7798 & ~n7807;
  assign n7809 = po35  & ~n7808;
  assign n7810 = ~n7394 & ~n7402;
  assign n7811 = n7400 & n7810;
  assign n7812 = po26  & n7811;
  assign n7813 = po26  & n7810;
  assign n7814 = ~n7400 & ~n7813;
  assign n7815 = ~n7812 & ~n7814;
  assign n7816 = ~po35  & n7808;
  assign n7817 = ~n7815 & ~n7816;
  assign n7818 = ~n7809 & ~n7817;
  assign n7819 = po36  & ~n7818;
  assign n7820 = ~n7405 & ~n7412;
  assign n7821 = n7411 & n7820;
  assign n7822 = po26  & n7821;
  assign n7823 = po26  & n7820;
  assign n7824 = ~n7411 & ~n7823;
  assign n7825 = ~n7822 & ~n7824;
  assign n7826 = ~po36  & ~n7809;
  assign n7827 = ~n7817 & n7826;
  assign n7828 = ~n7825 & ~n7827;
  assign n7829 = ~n7819 & ~n7828;
  assign n7830 = po37  & ~n7829;
  assign n7831 = ~n7415 & ~n7423;
  assign n7832 = n7421 & n7831;
  assign n7833 = po26  & n7832;
  assign n7834 = po26  & n7831;
  assign n7835 = ~n7421 & ~n7834;
  assign n7836 = ~n7833 & ~n7835;
  assign n7837 = ~po37  & n7829;
  assign n7838 = ~n7836 & ~n7837;
  assign n7839 = ~n7830 & ~n7838;
  assign n7840 = po38  & ~n7839;
  assign n7841 = ~n7426 & ~n7433;
  assign n7842 = n7432 & n7841;
  assign n7843 = po26  & n7842;
  assign n7844 = po26  & n7841;
  assign n7845 = ~n7432 & ~n7844;
  assign n7846 = ~n7843 & ~n7845;
  assign n7847 = ~po38  & ~n7830;
  assign n7848 = ~n7838 & n7847;
  assign n7849 = ~n7846 & ~n7848;
  assign n7850 = ~n7840 & ~n7849;
  assign n7851 = po39  & ~n7850;
  assign n7852 = ~n7436 & ~n7438;
  assign n7853 = n7444 & n7852;
  assign n7854 = po26  & n7853;
  assign n7855 = po26  & n7852;
  assign n7856 = ~n7444 & ~n7855;
  assign n7857 = ~n7854 & ~n7856;
  assign n7858 = ~po39  & n7850;
  assign n7859 = ~n7857 & ~n7858;
  assign n7860 = ~n7851 & ~n7859;
  assign n7861 = po40  & ~n7860;
  assign n7862 = ~n7447 & ~n7454;
  assign n7863 = n7453 & n7862;
  assign n7864 = po26  & n7863;
  assign n7865 = po26  & n7862;
  assign n7866 = ~n7453 & ~n7865;
  assign n7867 = ~n7864 & ~n7866;
  assign n7868 = ~po40  & ~n7851;
  assign n7869 = ~n7859 & n7868;
  assign n7870 = ~n7867 & ~n7869;
  assign n7871 = ~n7861 & ~n7870;
  assign n7872 = po41  & ~n7871;
  assign n7873 = ~n7457 & ~n7465;
  assign n7874 = n7463 & n7873;
  assign n7875 = po26  & n7874;
  assign n7876 = po26  & n7873;
  assign n7877 = ~n7463 & ~n7876;
  assign n7878 = ~n7875 & ~n7877;
  assign n7879 = ~po41  & n7871;
  assign n7880 = ~n7878 & ~n7879;
  assign n7881 = ~n7872 & ~n7880;
  assign n7882 = po42  & ~n7881;
  assign n7883 = ~n7468 & ~n7475;
  assign n7884 = n7474 & n7883;
  assign n7885 = po26  & n7884;
  assign n7886 = po26  & n7883;
  assign n7887 = ~n7474 & ~n7886;
  assign n7888 = ~n7885 & ~n7887;
  assign n7889 = ~po42  & ~n7872;
  assign n7890 = ~n7880 & n7889;
  assign n7891 = ~n7888 & ~n7890;
  assign n7892 = ~n7882 & ~n7891;
  assign n7893 = po43  & ~n7892;
  assign n7894 = ~n7478 & ~n7486;
  assign n7895 = n7484 & n7894;
  assign n7896 = po26  & n7895;
  assign n7897 = po26  & n7894;
  assign n7898 = ~n7484 & ~n7897;
  assign n7899 = ~n7896 & ~n7898;
  assign n7900 = ~po43  & n7892;
  assign n7901 = ~n7899 & ~n7900;
  assign n7902 = ~n7893 & ~n7901;
  assign n7903 = po44  & ~n7902;
  assign n7904 = ~n7489 & ~n7496;
  assign n7905 = n7495 & n7904;
  assign n7906 = po26  & n7905;
  assign n7907 = po26  & n7904;
  assign n7908 = ~n7495 & ~n7907;
  assign n7909 = ~n7906 & ~n7908;
  assign n7910 = ~po44  & ~n7893;
  assign n7911 = ~n7901 & n7910;
  assign n7912 = ~n7909 & ~n7911;
  assign n7913 = ~n7903 & ~n7912;
  assign n7914 = po45  & ~n7913;
  assign n7915 = ~n7499 & ~n7507;
  assign n7916 = n7505 & n7915;
  assign n7917 = po26  & n7916;
  assign n7918 = po26  & n7915;
  assign n7919 = ~n7505 & ~n7918;
  assign n7920 = ~n7917 & ~n7919;
  assign n7921 = ~po45  & n7913;
  assign n7922 = ~n7920 & ~n7921;
  assign n7923 = ~n7914 & ~n7922;
  assign n7924 = po46  & ~n7923;
  assign n7925 = ~n7510 & ~n7517;
  assign n7926 = n7516 & n7925;
  assign n7927 = po26  & n7926;
  assign n7928 = po26  & n7925;
  assign n7929 = ~n7516 & ~n7928;
  assign n7930 = ~n7927 & ~n7929;
  assign n7931 = ~po46  & ~n7914;
  assign n7932 = ~n7922 & n7931;
  assign n7933 = ~n7930 & ~n7932;
  assign n7934 = ~n7924 & ~n7933;
  assign n7935 = po47  & ~n7934;
  assign n7936 = ~n7520 & ~n7528;
  assign n7937 = n7526 & n7936;
  assign n7938 = po26  & n7937;
  assign n7939 = po26  & n7936;
  assign n7940 = ~n7526 & ~n7939;
  assign n7941 = ~n7938 & ~n7940;
  assign n7942 = ~po47  & n7934;
  assign n7943 = ~n7941 & ~n7942;
  assign n7944 = ~n7935 & ~n7943;
  assign n7945 = po48  & ~n7944;
  assign n7946 = ~n7531 & ~n7538;
  assign n7947 = n7537 & n7946;
  assign n7948 = po26  & n7947;
  assign n7949 = po26  & n7946;
  assign n7950 = ~n7537 & ~n7949;
  assign n7951 = ~n7948 & ~n7950;
  assign n7952 = ~po48  & ~n7935;
  assign n7953 = ~n7943 & n7952;
  assign n7954 = ~n7951 & ~n7953;
  assign n7955 = ~n7945 & ~n7954;
  assign n7956 = po49  & ~n7955;
  assign n7957 = ~n7541 & ~n7549;
  assign n7958 = n7547 & n7957;
  assign n7959 = po26  & n7958;
  assign n7960 = po26  & n7957;
  assign n7961 = ~n7547 & ~n7960;
  assign n7962 = ~n7959 & ~n7961;
  assign n7963 = ~po49  & n7955;
  assign n7964 = ~n7962 & ~n7963;
  assign n7965 = ~n7956 & ~n7964;
  assign n7966 = po50  & ~n7965;
  assign n7967 = ~n7552 & ~n7559;
  assign n7968 = n7558 & n7967;
  assign n7969 = po26  & n7968;
  assign n7970 = po26  & n7967;
  assign n7971 = ~n7558 & ~n7970;
  assign n7972 = ~n7969 & ~n7971;
  assign n7973 = ~po50  & ~n7956;
  assign n7974 = ~n7964 & n7973;
  assign n7975 = ~n7972 & ~n7974;
  assign n7976 = ~n7966 & ~n7975;
  assign n7977 = po51  & ~n7976;
  assign n7978 = ~n7562 & ~n7570;
  assign n7979 = n7568 & n7978;
  assign n7980 = po26  & n7979;
  assign n7981 = po26  & n7978;
  assign n7982 = ~n7568 & ~n7981;
  assign n7983 = ~n7980 & ~n7982;
  assign n7984 = ~po51  & n7976;
  assign n7985 = ~n7983 & ~n7984;
  assign n7986 = ~n7977 & ~n7985;
  assign n7987 = po52  & ~n7986;
  assign n7988 = ~n7573 & ~n7580;
  assign n7989 = n7579 & n7988;
  assign n7990 = po26  & n7989;
  assign n7991 = po26  & n7988;
  assign n7992 = ~n7579 & ~n7991;
  assign n7993 = ~n7990 & ~n7992;
  assign n7994 = ~po52  & ~n7977;
  assign n7995 = ~n7985 & n7994;
  assign n7996 = ~n7993 & ~n7995;
  assign n7997 = ~n7987 & ~n7996;
  assign n7998 = po53  & ~n7997;
  assign n7999 = ~n7583 & ~n7591;
  assign n8000 = n7589 & n7999;
  assign n8001 = po26  & n8000;
  assign n8002 = po26  & n7999;
  assign n8003 = ~n7589 & ~n8002;
  assign n8004 = ~n8001 & ~n8003;
  assign n8005 = ~po53  & n7997;
  assign n8006 = ~n8004 & ~n8005;
  assign n8007 = ~n7998 & ~n8006;
  assign n8008 = po54  & ~n8007;
  assign n8009 = ~n7594 & ~n7601;
  assign n8010 = n7600 & n8009;
  assign n8011 = po26  & n8010;
  assign n8012 = po26  & n8009;
  assign n8013 = ~n7600 & ~n8012;
  assign n8014 = ~n8011 & ~n8013;
  assign n8015 = ~po54  & ~n7998;
  assign n8016 = ~n8006 & n8015;
  assign n8017 = ~n8014 & ~n8016;
  assign n8018 = ~n8008 & ~n8017;
  assign n8019 = po55  & ~n8018;
  assign n8020 = ~n7604 & ~n7612;
  assign n8021 = n7610 & n8020;
  assign n8022 = po26  & n8021;
  assign n8023 = po26  & n8020;
  assign n8024 = ~n7610 & ~n8023;
  assign n8025 = ~n8022 & ~n8024;
  assign n8026 = ~po55  & n8018;
  assign n8027 = ~n8025 & ~n8026;
  assign n8028 = ~n8019 & ~n8027;
  assign n8029 = po56  & ~n8028;
  assign n8030 = ~n7615 & ~n7622;
  assign n8031 = n7621 & n8030;
  assign n8032 = po26  & n8031;
  assign n8033 = po26  & n8030;
  assign n8034 = ~n7621 & ~n8033;
  assign n8035 = ~n8032 & ~n8034;
  assign n8036 = ~po56  & ~n8019;
  assign n8037 = ~n8027 & n8036;
  assign n8038 = ~n8035 & ~n8037;
  assign n8039 = ~n8029 & ~n8038;
  assign n8040 = po57  & ~n8039;
  assign n8041 = ~n7625 & ~n7633;
  assign n8042 = n7631 & n8041;
  assign n8043 = po26  & n8042;
  assign n8044 = po26  & n8041;
  assign n8045 = ~n7631 & ~n8044;
  assign n8046 = ~n8043 & ~n8045;
  assign n8047 = ~po57  & n8039;
  assign n8048 = ~n8046 & ~n8047;
  assign n8049 = ~n8040 & ~n8048;
  assign n8050 = po58  & ~n8049;
  assign n8051 = ~n7636 & ~n7643;
  assign n8052 = n7642 & n8051;
  assign n8053 = po26  & n8052;
  assign n8054 = po26  & n8051;
  assign n8055 = ~n7642 & ~n8054;
  assign n8056 = ~n8053 & ~n8055;
  assign n8057 = ~po58  & ~n8040;
  assign n8058 = ~n8048 & n8057;
  assign n8059 = ~n8056 & ~n8058;
  assign n8060 = ~n8050 & ~n8059;
  assign n8061 = po59  & ~n8060;
  assign n8062 = ~n7646 & ~n7654;
  assign n8063 = n7652 & n8062;
  assign n8064 = po26  & n8063;
  assign n8065 = po26  & n8062;
  assign n8066 = ~n7652 & ~n8065;
  assign n8067 = ~n8064 & ~n8066;
  assign n8068 = ~po59  & n8060;
  assign n8069 = ~n8067 & ~n8068;
  assign n8070 = ~n8061 & ~n8069;
  assign n8071 = po60  & ~n8070;
  assign n8072 = ~n7657 & ~n7664;
  assign n8073 = n7663 & n8072;
  assign n8074 = po26  & n8073;
  assign n8075 = po26  & n8072;
  assign n8076 = ~n7663 & ~n8075;
  assign n8077 = ~n8074 & ~n8076;
  assign n8078 = ~po60  & ~n8061;
  assign n8079 = ~n8069 & n8078;
  assign n8080 = ~n8077 & ~n8079;
  assign n8081 = ~n8071 & ~n8080;
  assign n8082 = po61  & ~n8081;
  assign n8083 = ~n7667 & ~n7675;
  assign n8084 = n7673 & n8083;
  assign n8085 = po26  & n8084;
  assign n8086 = po26  & n8083;
  assign n8087 = ~n7673 & ~n8086;
  assign n8088 = ~n8085 & ~n8087;
  assign n8089 = ~po61  & n8081;
  assign n8090 = ~n8088 & ~n8089;
  assign n8091 = ~n8082 & ~n8090;
  assign n8092 = po62  & ~n8091;
  assign n8093 = ~n7678 & ~n7685;
  assign n8094 = n7684 & n8093;
  assign n8095 = po26  & n8094;
  assign n8096 = po26  & n8093;
  assign n8097 = ~n7684 & ~n8096;
  assign n8098 = ~n8095 & ~n8097;
  assign n8099 = ~po62  & ~n8082;
  assign n8100 = ~n8090 & n8099;
  assign n8101 = ~n8098 & ~n8100;
  assign n8102 = ~n8092 & ~n8101;
  assign n8103 = ~n7688 & ~n7696;
  assign n8104 = po26  & n8103;
  assign n8105 = ~n7694 & ~n8104;
  assign n8106 = n7694 & n8104;
  assign n8107 = ~n8105 & ~n8106;
  assign n8108 = ~n7698 & ~n7703;
  assign n8109 = po26  & n8108;
  assign n8110 = ~n7716 & ~n8109;
  assign n8111 = ~n8107 & n8110;
  assign n8112 = ~n8102 & n8111;
  assign n8113 = ~po63  & ~n8112;
  assign n8114 = ~n7703 & po26 ;
  assign n8115 = n7698 & ~n8114;
  assign n8116 = po63  & ~n8108;
  assign n8117 = ~n8115 & n8116;
  assign n8118 = n7703 & ~po26 ;
  assign n8119 = ~n8117 & ~n8118;
  assign n8120 = n8102 & n8107;
  assign n8121 = n8119 & ~n8120;
  assign po25  = n8113 | ~n8121;
  assign n8123 = pi50  & po25 ;
  assign n8124 = ~pi48  & ~pi49 ;
  assign n8125 = ~pi50  & n8124;
  assign n8126 = ~n8123 & ~n8125;
  assign n8127 = po26  & ~n8126;
  assign n8128 = n7715 & ~n8125;
  assign n8129 = ~n7716 & n8128;
  assign n8130 = ~n7709 & n8129;
  assign n8131 = ~n8123 & n8130;
  assign n8132 = ~pi50  & po25 ;
  assign n8133 = pi51  & ~n8132;
  assign n8134 = n7720 & po25 ;
  assign n8135 = ~n8133 & ~n8134;
  assign n8136 = ~n8131 & n8135;
  assign n8137 = ~n8127 & ~n8136;
  assign n8138 = po27  & ~n8137;
  assign n8139 = po26  & n8119;
  assign n8140 = ~n8120 & n8139;
  assign n8141 = ~n8113 & n8140;
  assign n8142 = ~n8134 & ~n8141;
  assign n8143 = pi52  & ~n8142;
  assign n8144 = ~pi52  & n8142;
  assign n8145 = ~n8143 & ~n8144;
  assign n8146 = ~po27  & n8137;
  assign n8147 = ~n8145 & ~n8146;
  assign n8148 = ~n8138 & ~n8147;
  assign n8149 = po28  & ~n8148;
  assign n8150 = ~n7723 & ~n7727;
  assign n8151 = ~n7731 & n8150;
  assign n8152 = po25  & n8151;
  assign n8153 = po25  & n8150;
  assign n8154 = n7731 & ~n8153;
  assign n8155 = ~n8152 & ~n8154;
  assign n8156 = ~po28  & ~n8138;
  assign n8157 = ~n8147 & n8156;
  assign n8158 = ~n8155 & ~n8157;
  assign n8159 = ~n8149 & ~n8158;
  assign n8160 = po29  & ~n8159;
  assign n8161 = ~n7734 & ~n7736;
  assign n8162 = n7743 & n8161;
  assign n8163 = po25  & n8162;
  assign n8164 = po25  & n8161;
  assign n8165 = ~n7743 & ~n8164;
  assign n8166 = ~n8163 & ~n8165;
  assign n8167 = ~po29  & n8159;
  assign n8168 = ~n8166 & ~n8167;
  assign n8169 = ~n8160 & ~n8168;
  assign n8170 = po30  & ~n8169;
  assign n8171 = ~n7746 & ~n7753;
  assign n8172 = n7752 & n8171;
  assign n8173 = po25  & n8172;
  assign n8174 = po25  & n8171;
  assign n8175 = ~n7752 & ~n8174;
  assign n8176 = ~n8173 & ~n8175;
  assign n8177 = ~po30  & ~n8160;
  assign n8178 = ~n8168 & n8177;
  assign n8179 = ~n8176 & ~n8178;
  assign n8180 = ~n8170 & ~n8179;
  assign n8181 = po31  & ~n8180;
  assign n8182 = ~n7756 & ~n7764;
  assign n8183 = n7762 & n8182;
  assign n8184 = po25  & n8183;
  assign n8185 = po25  & n8182;
  assign n8186 = ~n7762 & ~n8185;
  assign n8187 = ~n8184 & ~n8186;
  assign n8188 = ~po31  & n8180;
  assign n8189 = ~n8187 & ~n8188;
  assign n8190 = ~n8181 & ~n8189;
  assign n8191 = po32  & ~n8190;
  assign n8192 = ~n7767 & ~n7774;
  assign n8193 = n7773 & n8192;
  assign n8194 = po25  & n8193;
  assign n8195 = po25  & n8192;
  assign n8196 = ~n7773 & ~n8195;
  assign n8197 = ~n8194 & ~n8196;
  assign n8198 = ~po32  & ~n8181;
  assign n8199 = ~n8189 & n8198;
  assign n8200 = ~n8197 & ~n8199;
  assign n8201 = ~n8191 & ~n8200;
  assign n8202 = po33  & ~n8201;
  assign n8203 = ~n7777 & ~n7785;
  assign n8204 = n7783 & n8203;
  assign n8205 = po25  & n8204;
  assign n8206 = po25  & n8203;
  assign n8207 = ~n7783 & ~n8206;
  assign n8208 = ~n8205 & ~n8207;
  assign n8209 = ~po33  & n8201;
  assign n8210 = ~n8208 & ~n8209;
  assign n8211 = ~n8202 & ~n8210;
  assign n8212 = po34  & ~n8211;
  assign n8213 = ~n7788 & ~n7795;
  assign n8214 = n7794 & n8213;
  assign n8215 = po25  & n8214;
  assign n8216 = po25  & n8213;
  assign n8217 = ~n7794 & ~n8216;
  assign n8218 = ~n8215 & ~n8217;
  assign n8219 = ~po34  & ~n8202;
  assign n8220 = ~n8210 & n8219;
  assign n8221 = ~n8218 & ~n8220;
  assign n8222 = ~n8212 & ~n8221;
  assign n8223 = po35  & ~n8222;
  assign n8224 = ~n7798 & ~n7806;
  assign n8225 = n7804 & n8224;
  assign n8226 = po25  & n8225;
  assign n8227 = po25  & n8224;
  assign n8228 = ~n7804 & ~n8227;
  assign n8229 = ~n8226 & ~n8228;
  assign n8230 = ~po35  & n8222;
  assign n8231 = ~n8229 & ~n8230;
  assign n8232 = ~n8223 & ~n8231;
  assign n8233 = po36  & ~n8232;
  assign n8234 = ~n7809 & ~n7816;
  assign n8235 = n7815 & n8234;
  assign n8236 = po25  & n8235;
  assign n8237 = po25  & n8234;
  assign n8238 = ~n7815 & ~n8237;
  assign n8239 = ~n8236 & ~n8238;
  assign n8240 = ~po36  & ~n8223;
  assign n8241 = ~n8231 & n8240;
  assign n8242 = ~n8239 & ~n8241;
  assign n8243 = ~n8233 & ~n8242;
  assign n8244 = po37  & ~n8243;
  assign n8245 = ~n7819 & ~n7827;
  assign n8246 = n7825 & n8245;
  assign n8247 = po25  & n8246;
  assign n8248 = po25  & n8245;
  assign n8249 = ~n7825 & ~n8248;
  assign n8250 = ~n8247 & ~n8249;
  assign n8251 = ~po37  & n8243;
  assign n8252 = ~n8250 & ~n8251;
  assign n8253 = ~n8244 & ~n8252;
  assign n8254 = po38  & ~n8253;
  assign n8255 = ~n7830 & ~n7837;
  assign n8256 = n7836 & n8255;
  assign n8257 = po25  & n8256;
  assign n8258 = po25  & n8255;
  assign n8259 = ~n7836 & ~n8258;
  assign n8260 = ~n8257 & ~n8259;
  assign n8261 = ~po38  & ~n8244;
  assign n8262 = ~n8252 & n8261;
  assign n8263 = ~n8260 & ~n8262;
  assign n8264 = ~n8254 & ~n8263;
  assign n8265 = po39  & ~n8264;
  assign n8266 = ~n7840 & ~n7848;
  assign n8267 = n7846 & n8266;
  assign n8268 = po25  & n8267;
  assign n8269 = po25  & n8266;
  assign n8270 = ~n7846 & ~n8269;
  assign n8271 = ~n8268 & ~n8270;
  assign n8272 = ~po39  & n8264;
  assign n8273 = ~n8271 & ~n8272;
  assign n8274 = ~n8265 & ~n8273;
  assign n8275 = po40  & ~n8274;
  assign n8276 = ~po40  & ~n8265;
  assign n8277 = ~n8273 & n8276;
  assign n8278 = ~n7851 & ~n7858;
  assign n8279 = n7857 & n8278;
  assign n8280 = po25  & n8279;
  assign n8281 = po25  & n8278;
  assign n8282 = ~n7857 & ~n8281;
  assign n8283 = ~n8280 & ~n8282;
  assign n8284 = ~n8277 & ~n8283;
  assign n8285 = ~n8275 & ~n8284;
  assign n8286 = po41  & ~n8285;
  assign n8287 = ~n7861 & ~n7869;
  assign n8288 = n7867 & n8287;
  assign n8289 = po25  & n8288;
  assign n8290 = po25  & n8287;
  assign n8291 = ~n7867 & ~n8290;
  assign n8292 = ~n8289 & ~n8291;
  assign n8293 = ~po41  & n8285;
  assign n8294 = ~n8292 & ~n8293;
  assign n8295 = ~n8286 & ~n8294;
  assign n8296 = po42  & ~n8295;
  assign n8297 = ~n7872 & ~n7879;
  assign n8298 = n7878 & n8297;
  assign n8299 = po25  & n8298;
  assign n8300 = po25  & n8297;
  assign n8301 = ~n7878 & ~n8300;
  assign n8302 = ~n8299 & ~n8301;
  assign n8303 = ~po42  & ~n8286;
  assign n8304 = ~n8294 & n8303;
  assign n8305 = ~n8302 & ~n8304;
  assign n8306 = ~n8296 & ~n8305;
  assign n8307 = po43  & ~n8306;
  assign n8308 = ~n7882 & ~n7890;
  assign n8309 = n7888 & n8308;
  assign n8310 = po25  & n8309;
  assign n8311 = po25  & n8308;
  assign n8312 = ~n7888 & ~n8311;
  assign n8313 = ~n8310 & ~n8312;
  assign n8314 = ~po43  & n8306;
  assign n8315 = ~n8313 & ~n8314;
  assign n8316 = ~n8307 & ~n8315;
  assign n8317 = po44  & ~n8316;
  assign n8318 = ~n7893 & ~n7900;
  assign n8319 = n7899 & n8318;
  assign n8320 = po25  & n8319;
  assign n8321 = po25  & n8318;
  assign n8322 = ~n7899 & ~n8321;
  assign n8323 = ~n8320 & ~n8322;
  assign n8324 = ~po44  & ~n8307;
  assign n8325 = ~n8315 & n8324;
  assign n8326 = ~n8323 & ~n8325;
  assign n8327 = ~n8317 & ~n8326;
  assign n8328 = po45  & ~n8327;
  assign n8329 = ~n7903 & ~n7911;
  assign n8330 = n7909 & n8329;
  assign n8331 = po25  & n8330;
  assign n8332 = po25  & n8329;
  assign n8333 = ~n7909 & ~n8332;
  assign n8334 = ~n8331 & ~n8333;
  assign n8335 = ~po45  & n8327;
  assign n8336 = ~n8334 & ~n8335;
  assign n8337 = ~n8328 & ~n8336;
  assign n8338 = po46  & ~n8337;
  assign n8339 = ~n7914 & ~n7921;
  assign n8340 = n7920 & n8339;
  assign n8341 = po25  & n8340;
  assign n8342 = po25  & n8339;
  assign n8343 = ~n7920 & ~n8342;
  assign n8344 = ~n8341 & ~n8343;
  assign n8345 = ~po46  & ~n8328;
  assign n8346 = ~n8336 & n8345;
  assign n8347 = ~n8344 & ~n8346;
  assign n8348 = ~n8338 & ~n8347;
  assign n8349 = po47  & ~n8348;
  assign n8350 = ~n7924 & ~n7932;
  assign n8351 = n7930 & n8350;
  assign n8352 = po25  & n8351;
  assign n8353 = po25  & n8350;
  assign n8354 = ~n7930 & ~n8353;
  assign n8355 = ~n8352 & ~n8354;
  assign n8356 = ~po47  & n8348;
  assign n8357 = ~n8355 & ~n8356;
  assign n8358 = ~n8349 & ~n8357;
  assign n8359 = po48  & ~n8358;
  assign n8360 = ~n7935 & ~n7942;
  assign n8361 = n7941 & n8360;
  assign n8362 = po25  & n8361;
  assign n8363 = po25  & n8360;
  assign n8364 = ~n7941 & ~n8363;
  assign n8365 = ~n8362 & ~n8364;
  assign n8366 = ~po48  & ~n8349;
  assign n8367 = ~n8357 & n8366;
  assign n8368 = ~n8365 & ~n8367;
  assign n8369 = ~n8359 & ~n8368;
  assign n8370 = po49  & ~n8369;
  assign n8371 = ~n7945 & ~n7953;
  assign n8372 = n7951 & n8371;
  assign n8373 = po25  & n8372;
  assign n8374 = po25  & n8371;
  assign n8375 = ~n7951 & ~n8374;
  assign n8376 = ~n8373 & ~n8375;
  assign n8377 = ~po49  & n8369;
  assign n8378 = ~n8376 & ~n8377;
  assign n8379 = ~n8370 & ~n8378;
  assign n8380 = po50  & ~n8379;
  assign n8381 = ~n7956 & ~n7963;
  assign n8382 = n7962 & n8381;
  assign n8383 = po25  & n8382;
  assign n8384 = po25  & n8381;
  assign n8385 = ~n7962 & ~n8384;
  assign n8386 = ~n8383 & ~n8385;
  assign n8387 = ~po50  & ~n8370;
  assign n8388 = ~n8378 & n8387;
  assign n8389 = ~n8386 & ~n8388;
  assign n8390 = ~n8380 & ~n8389;
  assign n8391 = po51  & ~n8390;
  assign n8392 = ~n7966 & ~n7974;
  assign n8393 = n7972 & n8392;
  assign n8394 = po25  & n8393;
  assign n8395 = po25  & n8392;
  assign n8396 = ~n7972 & ~n8395;
  assign n8397 = ~n8394 & ~n8396;
  assign n8398 = ~po51  & n8390;
  assign n8399 = ~n8397 & ~n8398;
  assign n8400 = ~n8391 & ~n8399;
  assign n8401 = po52  & ~n8400;
  assign n8402 = ~n7977 & ~n7984;
  assign n8403 = n7983 & n8402;
  assign n8404 = po25  & n8403;
  assign n8405 = po25  & n8402;
  assign n8406 = ~n7983 & ~n8405;
  assign n8407 = ~n8404 & ~n8406;
  assign n8408 = ~po52  & ~n8391;
  assign n8409 = ~n8399 & n8408;
  assign n8410 = ~n8407 & ~n8409;
  assign n8411 = ~n8401 & ~n8410;
  assign n8412 = po53  & ~n8411;
  assign n8413 = ~n7987 & ~n7995;
  assign n8414 = n7993 & n8413;
  assign n8415 = po25  & n8414;
  assign n8416 = po25  & n8413;
  assign n8417 = ~n7993 & ~n8416;
  assign n8418 = ~n8415 & ~n8417;
  assign n8419 = ~po53  & n8411;
  assign n8420 = ~n8418 & ~n8419;
  assign n8421 = ~n8412 & ~n8420;
  assign n8422 = po54  & ~n8421;
  assign n8423 = ~n7998 & ~n8005;
  assign n8424 = n8004 & n8423;
  assign n8425 = po25  & n8424;
  assign n8426 = po25  & n8423;
  assign n8427 = ~n8004 & ~n8426;
  assign n8428 = ~n8425 & ~n8427;
  assign n8429 = ~po54  & ~n8412;
  assign n8430 = ~n8420 & n8429;
  assign n8431 = ~n8428 & ~n8430;
  assign n8432 = ~n8422 & ~n8431;
  assign n8433 = po55  & ~n8432;
  assign n8434 = ~n8008 & ~n8016;
  assign n8435 = n8014 & n8434;
  assign n8436 = po25  & n8435;
  assign n8437 = po25  & n8434;
  assign n8438 = ~n8014 & ~n8437;
  assign n8439 = ~n8436 & ~n8438;
  assign n8440 = ~po55  & n8432;
  assign n8441 = ~n8439 & ~n8440;
  assign n8442 = ~n8433 & ~n8441;
  assign n8443 = po56  & ~n8442;
  assign n8444 = ~n8019 & ~n8026;
  assign n8445 = n8025 & n8444;
  assign n8446 = po25  & n8445;
  assign n8447 = po25  & n8444;
  assign n8448 = ~n8025 & ~n8447;
  assign n8449 = ~n8446 & ~n8448;
  assign n8450 = ~po56  & ~n8433;
  assign n8451 = ~n8441 & n8450;
  assign n8452 = ~n8449 & ~n8451;
  assign n8453 = ~n8443 & ~n8452;
  assign n8454 = po57  & ~n8453;
  assign n8455 = ~n8029 & ~n8037;
  assign n8456 = n8035 & n8455;
  assign n8457 = po25  & n8456;
  assign n8458 = po25  & n8455;
  assign n8459 = ~n8035 & ~n8458;
  assign n8460 = ~n8457 & ~n8459;
  assign n8461 = ~po57  & n8453;
  assign n8462 = ~n8460 & ~n8461;
  assign n8463 = ~n8454 & ~n8462;
  assign n8464 = po58  & ~n8463;
  assign n8465 = ~n8040 & ~n8047;
  assign n8466 = n8046 & n8465;
  assign n8467 = po25  & n8466;
  assign n8468 = po25  & n8465;
  assign n8469 = ~n8046 & ~n8468;
  assign n8470 = ~n8467 & ~n8469;
  assign n8471 = ~po58  & ~n8454;
  assign n8472 = ~n8462 & n8471;
  assign n8473 = ~n8470 & ~n8472;
  assign n8474 = ~n8464 & ~n8473;
  assign n8475 = po59  & ~n8474;
  assign n8476 = ~n8050 & ~n8058;
  assign n8477 = n8056 & n8476;
  assign n8478 = po25  & n8477;
  assign n8479 = po25  & n8476;
  assign n8480 = ~n8056 & ~n8479;
  assign n8481 = ~n8478 & ~n8480;
  assign n8482 = ~po59  & n8474;
  assign n8483 = ~n8481 & ~n8482;
  assign n8484 = ~n8475 & ~n8483;
  assign n8485 = po60  & ~n8484;
  assign n8486 = ~n8061 & ~n8068;
  assign n8487 = n8067 & n8486;
  assign n8488 = po25  & n8487;
  assign n8489 = po25  & n8486;
  assign n8490 = ~n8067 & ~n8489;
  assign n8491 = ~n8488 & ~n8490;
  assign n8492 = ~po60  & ~n8475;
  assign n8493 = ~n8483 & n8492;
  assign n8494 = ~n8491 & ~n8493;
  assign n8495 = ~n8485 & ~n8494;
  assign n8496 = po61  & ~n8495;
  assign n8497 = ~n8071 & ~n8079;
  assign n8498 = n8077 & n8497;
  assign n8499 = po25  & n8498;
  assign n8500 = po25  & n8497;
  assign n8501 = ~n8077 & ~n8500;
  assign n8502 = ~n8499 & ~n8501;
  assign n8503 = ~po61  & n8495;
  assign n8504 = ~n8502 & ~n8503;
  assign n8505 = ~n8496 & ~n8504;
  assign n8506 = po62  & ~n8505;
  assign n8507 = ~n8082 & ~n8089;
  assign n8508 = n8088 & n8507;
  assign n8509 = po25  & n8508;
  assign n8510 = po25  & n8507;
  assign n8511 = ~n8088 & ~n8510;
  assign n8512 = ~n8509 & ~n8511;
  assign n8513 = ~po62  & ~n8496;
  assign n8514 = ~n8504 & n8513;
  assign n8515 = ~n8512 & ~n8514;
  assign n8516 = ~n8506 & ~n8515;
  assign n8517 = ~n8092 & ~n8100;
  assign n8518 = po25  & n8517;
  assign n8519 = ~n8098 & ~n8518;
  assign n8520 = n8098 & n8518;
  assign n8521 = ~n8519 & ~n8520;
  assign n8522 = ~n8102 & ~n8107;
  assign n8523 = po25  & n8522;
  assign n8524 = ~n8120 & ~n8523;
  assign n8525 = ~n8521 & n8524;
  assign n8526 = ~n8516 & n8525;
  assign n8527 = ~po63  & ~n8526;
  assign n8528 = ~n8107 & po25 ;
  assign n8529 = n8102 & ~n8528;
  assign n8530 = po63  & ~n8522;
  assign n8531 = ~n8529 & n8530;
  assign n8532 = n8107 & ~po25 ;
  assign n8533 = ~n8531 & ~n8532;
  assign n8534 = n8516 & n8521;
  assign n8535 = n8533 & ~n8534;
  assign po24  = n8527 | ~n8535;
  assign n8537 = pi48  & po24 ;
  assign n8538 = ~pi46  & ~pi47 ;
  assign n8539 = ~pi48  & n8538;
  assign n8540 = ~n8537 & ~n8539;
  assign n8541 = po25  & ~n8540;
  assign n8542 = n8119 & ~n8539;
  assign n8543 = ~n8120 & n8542;
  assign n8544 = ~n8113 & n8543;
  assign n8545 = ~n8537 & n8544;
  assign n8546 = ~pi48  & po24 ;
  assign n8547 = pi49  & ~n8546;
  assign n8548 = n8124 & po24 ;
  assign n8549 = ~n8547 & ~n8548;
  assign n8550 = ~n8545 & n8549;
  assign n8551 = ~n8541 & ~n8550;
  assign n8552 = po26  & ~n8551;
  assign n8553 = ~po26  & ~n8541;
  assign n8554 = ~n8550 & n8553;
  assign n8555 = po25  & n8533;
  assign n8556 = ~n8534 & n8555;
  assign n8557 = ~n8527 & n8556;
  assign n8558 = ~n8548 & ~n8557;
  assign n8559 = pi50  & ~n8558;
  assign n8560 = ~pi50  & n8558;
  assign n8561 = ~n8559 & ~n8560;
  assign n8562 = ~n8554 & ~n8561;
  assign n8563 = ~n8552 & ~n8562;
  assign n8564 = po27  & ~n8563;
  assign n8565 = ~n8127 & ~n8131;
  assign n8566 = ~n8135 & n8565;
  assign n8567 = po24  & n8566;
  assign n8568 = po24  & n8565;
  assign n8569 = n8135 & ~n8568;
  assign n8570 = ~n8567 & ~n8569;
  assign n8571 = ~po27  & n8563;
  assign n8572 = ~n8570 & ~n8571;
  assign n8573 = ~n8564 & ~n8572;
  assign n8574 = po28  & ~n8573;
  assign n8575 = ~n8138 & ~n8146;
  assign n8576 = n8145 & n8575;
  assign n8577 = po24  & n8576;
  assign n8578 = po24  & n8575;
  assign n8579 = ~n8145 & ~n8578;
  assign n8580 = ~n8577 & ~n8579;
  assign n8581 = ~po28  & ~n8564;
  assign n8582 = ~n8572 & n8581;
  assign n8583 = ~n8580 & ~n8582;
  assign n8584 = ~n8574 & ~n8583;
  assign n8585 = po29  & ~n8584;
  assign n8586 = ~n8149 & ~n8157;
  assign n8587 = n8155 & n8586;
  assign n8588 = po24  & n8587;
  assign n8589 = po24  & n8586;
  assign n8590 = ~n8155 & ~n8589;
  assign n8591 = ~n8588 & ~n8590;
  assign n8592 = ~po29  & n8584;
  assign n8593 = ~n8591 & ~n8592;
  assign n8594 = ~n8585 & ~n8593;
  assign n8595 = po30  & ~n8594;
  assign n8596 = ~n8160 & ~n8167;
  assign n8597 = n8166 & n8596;
  assign n8598 = po24  & n8597;
  assign n8599 = po24  & n8596;
  assign n8600 = ~n8166 & ~n8599;
  assign n8601 = ~n8598 & ~n8600;
  assign n8602 = ~po30  & ~n8585;
  assign n8603 = ~n8593 & n8602;
  assign n8604 = ~n8601 & ~n8603;
  assign n8605 = ~n8595 & ~n8604;
  assign n8606 = po31  & ~n8605;
  assign n8607 = ~n8170 & ~n8178;
  assign n8608 = n8176 & n8607;
  assign n8609 = po24  & n8608;
  assign n8610 = po24  & n8607;
  assign n8611 = ~n8176 & ~n8610;
  assign n8612 = ~n8609 & ~n8611;
  assign n8613 = ~po31  & n8605;
  assign n8614 = ~n8612 & ~n8613;
  assign n8615 = ~n8606 & ~n8614;
  assign n8616 = po32  & ~n8615;
  assign n8617 = ~n8181 & ~n8188;
  assign n8618 = n8187 & n8617;
  assign n8619 = po24  & n8618;
  assign n8620 = po24  & n8617;
  assign n8621 = ~n8187 & ~n8620;
  assign n8622 = ~n8619 & ~n8621;
  assign n8623 = ~po32  & ~n8606;
  assign n8624 = ~n8614 & n8623;
  assign n8625 = ~n8622 & ~n8624;
  assign n8626 = ~n8616 & ~n8625;
  assign n8627 = po33  & ~n8626;
  assign n8628 = ~n8191 & ~n8199;
  assign n8629 = n8197 & n8628;
  assign n8630 = po24  & n8629;
  assign n8631 = po24  & n8628;
  assign n8632 = ~n8197 & ~n8631;
  assign n8633 = ~n8630 & ~n8632;
  assign n8634 = ~po33  & n8626;
  assign n8635 = ~n8633 & ~n8634;
  assign n8636 = ~n8627 & ~n8635;
  assign n8637 = po34  & ~n8636;
  assign n8638 = ~n8202 & ~n8209;
  assign n8639 = n8208 & n8638;
  assign n8640 = po24  & n8639;
  assign n8641 = po24  & n8638;
  assign n8642 = ~n8208 & ~n8641;
  assign n8643 = ~n8640 & ~n8642;
  assign n8644 = ~po34  & ~n8627;
  assign n8645 = ~n8635 & n8644;
  assign n8646 = ~n8643 & ~n8645;
  assign n8647 = ~n8637 & ~n8646;
  assign n8648 = po35  & ~n8647;
  assign n8649 = ~n8212 & ~n8220;
  assign n8650 = n8218 & n8649;
  assign n8651 = po24  & n8650;
  assign n8652 = po24  & n8649;
  assign n8653 = ~n8218 & ~n8652;
  assign n8654 = ~n8651 & ~n8653;
  assign n8655 = ~po35  & n8647;
  assign n8656 = ~n8654 & ~n8655;
  assign n8657 = ~n8648 & ~n8656;
  assign n8658 = po36  & ~n8657;
  assign n8659 = ~n8223 & ~n8230;
  assign n8660 = n8229 & n8659;
  assign n8661 = po24  & n8660;
  assign n8662 = po24  & n8659;
  assign n8663 = ~n8229 & ~n8662;
  assign n8664 = ~n8661 & ~n8663;
  assign n8665 = ~po36  & ~n8648;
  assign n8666 = ~n8656 & n8665;
  assign n8667 = ~n8664 & ~n8666;
  assign n8668 = ~n8658 & ~n8667;
  assign n8669 = po37  & ~n8668;
  assign n8670 = ~n8233 & ~n8241;
  assign n8671 = n8239 & n8670;
  assign n8672 = po24  & n8671;
  assign n8673 = po24  & n8670;
  assign n8674 = ~n8239 & ~n8673;
  assign n8675 = ~n8672 & ~n8674;
  assign n8676 = ~po37  & n8668;
  assign n8677 = ~n8675 & ~n8676;
  assign n8678 = ~n8669 & ~n8677;
  assign n8679 = po38  & ~n8678;
  assign n8680 = ~n8244 & ~n8251;
  assign n8681 = n8250 & n8680;
  assign n8682 = po24  & n8681;
  assign n8683 = po24  & n8680;
  assign n8684 = ~n8250 & ~n8683;
  assign n8685 = ~n8682 & ~n8684;
  assign n8686 = ~po38  & ~n8669;
  assign n8687 = ~n8677 & n8686;
  assign n8688 = ~n8685 & ~n8687;
  assign n8689 = ~n8679 & ~n8688;
  assign n8690 = po39  & ~n8689;
  assign n8691 = ~n8254 & ~n8262;
  assign n8692 = n8260 & n8691;
  assign n8693 = po24  & n8692;
  assign n8694 = po24  & n8691;
  assign n8695 = ~n8260 & ~n8694;
  assign n8696 = ~n8693 & ~n8695;
  assign n8697 = ~po39  & n8689;
  assign n8698 = ~n8696 & ~n8697;
  assign n8699 = ~n8690 & ~n8698;
  assign n8700 = po40  & ~n8699;
  assign n8701 = ~n8265 & ~n8272;
  assign n8702 = n8271 & n8701;
  assign n8703 = po24  & n8702;
  assign n8704 = po24  & n8701;
  assign n8705 = ~n8271 & ~n8704;
  assign n8706 = ~n8703 & ~n8705;
  assign n8707 = ~po40  & ~n8690;
  assign n8708 = ~n8698 & n8707;
  assign n8709 = ~n8706 & ~n8708;
  assign n8710 = ~n8700 & ~n8709;
  assign n8711 = po41  & ~n8710;
  assign n8712 = ~n8275 & ~n8277;
  assign n8713 = n8283 & n8712;
  assign n8714 = po24  & n8713;
  assign n8715 = po24  & n8712;
  assign n8716 = ~n8283 & ~n8715;
  assign n8717 = ~n8714 & ~n8716;
  assign n8718 = ~po41  & n8710;
  assign n8719 = ~n8717 & ~n8718;
  assign n8720 = ~n8711 & ~n8719;
  assign n8721 = po42  & ~n8720;
  assign n8722 = ~n8286 & ~n8293;
  assign n8723 = n8292 & n8722;
  assign n8724 = po24  & n8723;
  assign n8725 = po24  & n8722;
  assign n8726 = ~n8292 & ~n8725;
  assign n8727 = ~n8724 & ~n8726;
  assign n8728 = ~po42  & ~n8711;
  assign n8729 = ~n8719 & n8728;
  assign n8730 = ~n8727 & ~n8729;
  assign n8731 = ~n8721 & ~n8730;
  assign n8732 = po43  & ~n8731;
  assign n8733 = ~n8296 & ~n8304;
  assign n8734 = n8302 & n8733;
  assign n8735 = po24  & n8734;
  assign n8736 = po24  & n8733;
  assign n8737 = ~n8302 & ~n8736;
  assign n8738 = ~n8735 & ~n8737;
  assign n8739 = ~po43  & n8731;
  assign n8740 = ~n8738 & ~n8739;
  assign n8741 = ~n8732 & ~n8740;
  assign n8742 = po44  & ~n8741;
  assign n8743 = ~n8307 & ~n8314;
  assign n8744 = n8313 & n8743;
  assign n8745 = po24  & n8744;
  assign n8746 = po24  & n8743;
  assign n8747 = ~n8313 & ~n8746;
  assign n8748 = ~n8745 & ~n8747;
  assign n8749 = ~po44  & ~n8732;
  assign n8750 = ~n8740 & n8749;
  assign n8751 = ~n8748 & ~n8750;
  assign n8752 = ~n8742 & ~n8751;
  assign n8753 = po45  & ~n8752;
  assign n8754 = ~n8317 & ~n8325;
  assign n8755 = n8323 & n8754;
  assign n8756 = po24  & n8755;
  assign n8757 = po24  & n8754;
  assign n8758 = ~n8323 & ~n8757;
  assign n8759 = ~n8756 & ~n8758;
  assign n8760 = ~po45  & n8752;
  assign n8761 = ~n8759 & ~n8760;
  assign n8762 = ~n8753 & ~n8761;
  assign n8763 = po46  & ~n8762;
  assign n8764 = ~n8328 & ~n8335;
  assign n8765 = n8334 & n8764;
  assign n8766 = po24  & n8765;
  assign n8767 = po24  & n8764;
  assign n8768 = ~n8334 & ~n8767;
  assign n8769 = ~n8766 & ~n8768;
  assign n8770 = ~po46  & ~n8753;
  assign n8771 = ~n8761 & n8770;
  assign n8772 = ~n8769 & ~n8771;
  assign n8773 = ~n8763 & ~n8772;
  assign n8774 = po47  & ~n8773;
  assign n8775 = ~n8338 & ~n8346;
  assign n8776 = n8344 & n8775;
  assign n8777 = po24  & n8776;
  assign n8778 = po24  & n8775;
  assign n8779 = ~n8344 & ~n8778;
  assign n8780 = ~n8777 & ~n8779;
  assign n8781 = ~po47  & n8773;
  assign n8782 = ~n8780 & ~n8781;
  assign n8783 = ~n8774 & ~n8782;
  assign n8784 = po48  & ~n8783;
  assign n8785 = ~n8349 & ~n8356;
  assign n8786 = n8355 & n8785;
  assign n8787 = po24  & n8786;
  assign n8788 = po24  & n8785;
  assign n8789 = ~n8355 & ~n8788;
  assign n8790 = ~n8787 & ~n8789;
  assign n8791 = ~po48  & ~n8774;
  assign n8792 = ~n8782 & n8791;
  assign n8793 = ~n8790 & ~n8792;
  assign n8794 = ~n8784 & ~n8793;
  assign n8795 = po49  & ~n8794;
  assign n8796 = ~n8359 & ~n8367;
  assign n8797 = n8365 & n8796;
  assign n8798 = po24  & n8797;
  assign n8799 = po24  & n8796;
  assign n8800 = ~n8365 & ~n8799;
  assign n8801 = ~n8798 & ~n8800;
  assign n8802 = ~po49  & n8794;
  assign n8803 = ~n8801 & ~n8802;
  assign n8804 = ~n8795 & ~n8803;
  assign n8805 = po50  & ~n8804;
  assign n8806 = ~n8370 & ~n8377;
  assign n8807 = n8376 & n8806;
  assign n8808 = po24  & n8807;
  assign n8809 = po24  & n8806;
  assign n8810 = ~n8376 & ~n8809;
  assign n8811 = ~n8808 & ~n8810;
  assign n8812 = ~po50  & ~n8795;
  assign n8813 = ~n8803 & n8812;
  assign n8814 = ~n8811 & ~n8813;
  assign n8815 = ~n8805 & ~n8814;
  assign n8816 = po51  & ~n8815;
  assign n8817 = ~n8380 & ~n8388;
  assign n8818 = n8386 & n8817;
  assign n8819 = po24  & n8818;
  assign n8820 = po24  & n8817;
  assign n8821 = ~n8386 & ~n8820;
  assign n8822 = ~n8819 & ~n8821;
  assign n8823 = ~po51  & n8815;
  assign n8824 = ~n8822 & ~n8823;
  assign n8825 = ~n8816 & ~n8824;
  assign n8826 = po52  & ~n8825;
  assign n8827 = ~n8391 & ~n8398;
  assign n8828 = n8397 & n8827;
  assign n8829 = po24  & n8828;
  assign n8830 = po24  & n8827;
  assign n8831 = ~n8397 & ~n8830;
  assign n8832 = ~n8829 & ~n8831;
  assign n8833 = ~po52  & ~n8816;
  assign n8834 = ~n8824 & n8833;
  assign n8835 = ~n8832 & ~n8834;
  assign n8836 = ~n8826 & ~n8835;
  assign n8837 = po53  & ~n8836;
  assign n8838 = ~n8401 & ~n8409;
  assign n8839 = n8407 & n8838;
  assign n8840 = po24  & n8839;
  assign n8841 = po24  & n8838;
  assign n8842 = ~n8407 & ~n8841;
  assign n8843 = ~n8840 & ~n8842;
  assign n8844 = ~po53  & n8836;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = ~n8837 & ~n8845;
  assign n8847 = po54  & ~n8846;
  assign n8848 = ~n8412 & ~n8419;
  assign n8849 = n8418 & n8848;
  assign n8850 = po24  & n8849;
  assign n8851 = po24  & n8848;
  assign n8852 = ~n8418 & ~n8851;
  assign n8853 = ~n8850 & ~n8852;
  assign n8854 = ~po54  & ~n8837;
  assign n8855 = ~n8845 & n8854;
  assign n8856 = ~n8853 & ~n8855;
  assign n8857 = ~n8847 & ~n8856;
  assign n8858 = po55  & ~n8857;
  assign n8859 = ~n8422 & ~n8430;
  assign n8860 = n8428 & n8859;
  assign n8861 = po24  & n8860;
  assign n8862 = po24  & n8859;
  assign n8863 = ~n8428 & ~n8862;
  assign n8864 = ~n8861 & ~n8863;
  assign n8865 = ~po55  & n8857;
  assign n8866 = ~n8864 & ~n8865;
  assign n8867 = ~n8858 & ~n8866;
  assign n8868 = po56  & ~n8867;
  assign n8869 = ~n8433 & ~n8440;
  assign n8870 = n8439 & n8869;
  assign n8871 = po24  & n8870;
  assign n8872 = po24  & n8869;
  assign n8873 = ~n8439 & ~n8872;
  assign n8874 = ~n8871 & ~n8873;
  assign n8875 = ~po56  & ~n8858;
  assign n8876 = ~n8866 & n8875;
  assign n8877 = ~n8874 & ~n8876;
  assign n8878 = ~n8868 & ~n8877;
  assign n8879 = po57  & ~n8878;
  assign n8880 = ~n8443 & ~n8451;
  assign n8881 = n8449 & n8880;
  assign n8882 = po24  & n8881;
  assign n8883 = po24  & n8880;
  assign n8884 = ~n8449 & ~n8883;
  assign n8885 = ~n8882 & ~n8884;
  assign n8886 = ~po57  & n8878;
  assign n8887 = ~n8885 & ~n8886;
  assign n8888 = ~n8879 & ~n8887;
  assign n8889 = po58  & ~n8888;
  assign n8890 = ~n8454 & ~n8461;
  assign n8891 = n8460 & n8890;
  assign n8892 = po24  & n8891;
  assign n8893 = po24  & n8890;
  assign n8894 = ~n8460 & ~n8893;
  assign n8895 = ~n8892 & ~n8894;
  assign n8896 = ~po58  & ~n8879;
  assign n8897 = ~n8887 & n8896;
  assign n8898 = ~n8895 & ~n8897;
  assign n8899 = ~n8889 & ~n8898;
  assign n8900 = po59  & ~n8899;
  assign n8901 = ~n8464 & ~n8472;
  assign n8902 = n8470 & n8901;
  assign n8903 = po24  & n8902;
  assign n8904 = po24  & n8901;
  assign n8905 = ~n8470 & ~n8904;
  assign n8906 = ~n8903 & ~n8905;
  assign n8907 = ~po59  & n8899;
  assign n8908 = ~n8906 & ~n8907;
  assign n8909 = ~n8900 & ~n8908;
  assign n8910 = po60  & ~n8909;
  assign n8911 = ~n8475 & ~n8482;
  assign n8912 = n8481 & n8911;
  assign n8913 = po24  & n8912;
  assign n8914 = po24  & n8911;
  assign n8915 = ~n8481 & ~n8914;
  assign n8916 = ~n8913 & ~n8915;
  assign n8917 = ~po60  & ~n8900;
  assign n8918 = ~n8908 & n8917;
  assign n8919 = ~n8916 & ~n8918;
  assign n8920 = ~n8910 & ~n8919;
  assign n8921 = po61  & ~n8920;
  assign n8922 = ~n8485 & ~n8493;
  assign n8923 = n8491 & n8922;
  assign n8924 = po24  & n8923;
  assign n8925 = po24  & n8922;
  assign n8926 = ~n8491 & ~n8925;
  assign n8927 = ~n8924 & ~n8926;
  assign n8928 = ~po61  & n8920;
  assign n8929 = ~n8927 & ~n8928;
  assign n8930 = ~n8921 & ~n8929;
  assign n8931 = po62  & ~n8930;
  assign n8932 = ~n8496 & ~n8503;
  assign n8933 = n8502 & n8932;
  assign n8934 = po24  & n8933;
  assign n8935 = po24  & n8932;
  assign n8936 = ~n8502 & ~n8935;
  assign n8937 = ~n8934 & ~n8936;
  assign n8938 = ~po62  & ~n8921;
  assign n8939 = ~n8929 & n8938;
  assign n8940 = ~n8937 & ~n8939;
  assign n8941 = ~n8931 & ~n8940;
  assign n8942 = ~n8506 & ~n8514;
  assign n8943 = po24  & n8942;
  assign n8944 = ~n8512 & ~n8943;
  assign n8945 = n8512 & n8943;
  assign n8946 = ~n8944 & ~n8945;
  assign n8947 = ~n8516 & ~n8521;
  assign n8948 = po24  & n8947;
  assign n8949 = ~n8534 & ~n8948;
  assign n8950 = ~n8946 & n8949;
  assign n8951 = ~n8941 & n8950;
  assign n8952 = ~po63  & ~n8951;
  assign n8953 = ~n8521 & po24 ;
  assign n8954 = n8516 & ~n8953;
  assign n8955 = po63  & ~n8947;
  assign n8956 = ~n8954 & n8955;
  assign n8957 = n8521 & ~po24 ;
  assign n8958 = ~n8956 & ~n8957;
  assign n8959 = n8941 & n8946;
  assign n8960 = n8958 & ~n8959;
  assign po23  = n8952 | ~n8960;
  assign n8962 = pi46  & po23 ;
  assign n8963 = ~pi44  & ~pi45 ;
  assign n8964 = ~pi46  & n8963;
  assign n8965 = ~n8962 & ~n8964;
  assign n8966 = po24  & ~n8965;
  assign n8967 = n8533 & ~n8964;
  assign n8968 = ~n8534 & n8967;
  assign n8969 = ~n8527 & n8968;
  assign n8970 = ~n8962 & n8969;
  assign n8971 = ~pi46  & po23 ;
  assign n8972 = pi47  & ~n8971;
  assign n8973 = n8538 & po23 ;
  assign n8974 = ~n8972 & ~n8973;
  assign n8975 = ~n8970 & n8974;
  assign n8976 = ~n8966 & ~n8975;
  assign n8977 = po25  & ~n8976;
  assign n8978 = po24  & n8958;
  assign n8979 = ~n8959 & n8978;
  assign n8980 = ~n8952 & n8979;
  assign n8981 = ~n8973 & ~n8980;
  assign n8982 = pi48  & ~n8981;
  assign n8983 = ~pi48  & n8981;
  assign n8984 = ~n8982 & ~n8983;
  assign n8985 = ~po25  & n8976;
  assign n8986 = ~n8984 & ~n8985;
  assign n8987 = ~n8977 & ~n8986;
  assign n8988 = po26  & ~n8987;
  assign n8989 = ~n8541 & ~n8545;
  assign n8990 = ~n8549 & n8989;
  assign n8991 = po23  & n8990;
  assign n8992 = po23  & n8989;
  assign n8993 = n8549 & ~n8992;
  assign n8994 = ~n8991 & ~n8993;
  assign n8995 = ~po26  & ~n8977;
  assign n8996 = ~n8986 & n8995;
  assign n8997 = ~n8994 & ~n8996;
  assign n8998 = ~n8988 & ~n8997;
  assign n8999 = po27  & ~n8998;
  assign n9000 = ~n8552 & ~n8554;
  assign n9001 = n8561 & n9000;
  assign n9002 = po23  & n9001;
  assign n9003 = po23  & n9000;
  assign n9004 = ~n8561 & ~n9003;
  assign n9005 = ~n9002 & ~n9004;
  assign n9006 = ~po27  & n8998;
  assign n9007 = ~n9005 & ~n9006;
  assign n9008 = ~n8999 & ~n9007;
  assign n9009 = po28  & ~n9008;
  assign n9010 = ~n8564 & ~n8571;
  assign n9011 = n8570 & n9010;
  assign n9012 = po23  & n9011;
  assign n9013 = po23  & n9010;
  assign n9014 = ~n8570 & ~n9013;
  assign n9015 = ~n9012 & ~n9014;
  assign n9016 = ~po28  & ~n8999;
  assign n9017 = ~n9007 & n9016;
  assign n9018 = ~n9015 & ~n9017;
  assign n9019 = ~n9009 & ~n9018;
  assign n9020 = po29  & ~n9019;
  assign n9021 = ~n8574 & ~n8582;
  assign n9022 = n8580 & n9021;
  assign n9023 = po23  & n9022;
  assign n9024 = po23  & n9021;
  assign n9025 = ~n8580 & ~n9024;
  assign n9026 = ~n9023 & ~n9025;
  assign n9027 = ~po29  & n9019;
  assign n9028 = ~n9026 & ~n9027;
  assign n9029 = ~n9020 & ~n9028;
  assign n9030 = po30  & ~n9029;
  assign n9031 = ~n8585 & ~n8592;
  assign n9032 = n8591 & n9031;
  assign n9033 = po23  & n9032;
  assign n9034 = po23  & n9031;
  assign n9035 = ~n8591 & ~n9034;
  assign n9036 = ~n9033 & ~n9035;
  assign n9037 = ~po30  & ~n9020;
  assign n9038 = ~n9028 & n9037;
  assign n9039 = ~n9036 & ~n9038;
  assign n9040 = ~n9030 & ~n9039;
  assign n9041 = po31  & ~n9040;
  assign n9042 = ~n8595 & ~n8603;
  assign n9043 = n8601 & n9042;
  assign n9044 = po23  & n9043;
  assign n9045 = po23  & n9042;
  assign n9046 = ~n8601 & ~n9045;
  assign n9047 = ~n9044 & ~n9046;
  assign n9048 = ~po31  & n9040;
  assign n9049 = ~n9047 & ~n9048;
  assign n9050 = ~n9041 & ~n9049;
  assign n9051 = po32  & ~n9050;
  assign n9052 = ~n8606 & ~n8613;
  assign n9053 = n8612 & n9052;
  assign n9054 = po23  & n9053;
  assign n9055 = po23  & n9052;
  assign n9056 = ~n8612 & ~n9055;
  assign n9057 = ~n9054 & ~n9056;
  assign n9058 = ~po32  & ~n9041;
  assign n9059 = ~n9049 & n9058;
  assign n9060 = ~n9057 & ~n9059;
  assign n9061 = ~n9051 & ~n9060;
  assign n9062 = po33  & ~n9061;
  assign n9063 = ~n8616 & ~n8624;
  assign n9064 = n8622 & n9063;
  assign n9065 = po23  & n9064;
  assign n9066 = po23  & n9063;
  assign n9067 = ~n8622 & ~n9066;
  assign n9068 = ~n9065 & ~n9067;
  assign n9069 = ~po33  & n9061;
  assign n9070 = ~n9068 & ~n9069;
  assign n9071 = ~n9062 & ~n9070;
  assign n9072 = po34  & ~n9071;
  assign n9073 = ~n8627 & ~n8634;
  assign n9074 = n8633 & n9073;
  assign n9075 = po23  & n9074;
  assign n9076 = po23  & n9073;
  assign n9077 = ~n8633 & ~n9076;
  assign n9078 = ~n9075 & ~n9077;
  assign n9079 = ~po34  & ~n9062;
  assign n9080 = ~n9070 & n9079;
  assign n9081 = ~n9078 & ~n9080;
  assign n9082 = ~n9072 & ~n9081;
  assign n9083 = po35  & ~n9082;
  assign n9084 = ~n8637 & ~n8645;
  assign n9085 = n8643 & n9084;
  assign n9086 = po23  & n9085;
  assign n9087 = po23  & n9084;
  assign n9088 = ~n8643 & ~n9087;
  assign n9089 = ~n9086 & ~n9088;
  assign n9090 = ~po35  & n9082;
  assign n9091 = ~n9089 & ~n9090;
  assign n9092 = ~n9083 & ~n9091;
  assign n9093 = po36  & ~n9092;
  assign n9094 = ~n8648 & ~n8655;
  assign n9095 = n8654 & n9094;
  assign n9096 = po23  & n9095;
  assign n9097 = po23  & n9094;
  assign n9098 = ~n8654 & ~n9097;
  assign n9099 = ~n9096 & ~n9098;
  assign n9100 = ~po36  & ~n9083;
  assign n9101 = ~n9091 & n9100;
  assign n9102 = ~n9099 & ~n9101;
  assign n9103 = ~n9093 & ~n9102;
  assign n9104 = po37  & ~n9103;
  assign n9105 = ~n8658 & ~n8666;
  assign n9106 = n8664 & n9105;
  assign n9107 = po23  & n9106;
  assign n9108 = po23  & n9105;
  assign n9109 = ~n8664 & ~n9108;
  assign n9110 = ~n9107 & ~n9109;
  assign n9111 = ~po37  & n9103;
  assign n9112 = ~n9110 & ~n9111;
  assign n9113 = ~n9104 & ~n9112;
  assign n9114 = po38  & ~n9113;
  assign n9115 = ~n8669 & ~n8676;
  assign n9116 = n8675 & n9115;
  assign n9117 = po23  & n9116;
  assign n9118 = po23  & n9115;
  assign n9119 = ~n8675 & ~n9118;
  assign n9120 = ~n9117 & ~n9119;
  assign n9121 = ~po38  & ~n9104;
  assign n9122 = ~n9112 & n9121;
  assign n9123 = ~n9120 & ~n9122;
  assign n9124 = ~n9114 & ~n9123;
  assign n9125 = po39  & ~n9124;
  assign n9126 = ~n8679 & ~n8687;
  assign n9127 = n8685 & n9126;
  assign n9128 = po23  & n9127;
  assign n9129 = po23  & n9126;
  assign n9130 = ~n8685 & ~n9129;
  assign n9131 = ~n9128 & ~n9130;
  assign n9132 = ~po39  & n9124;
  assign n9133 = ~n9131 & ~n9132;
  assign n9134 = ~n9125 & ~n9133;
  assign n9135 = po40  & ~n9134;
  assign n9136 = ~n8690 & ~n8697;
  assign n9137 = n8696 & n9136;
  assign n9138 = po23  & n9137;
  assign n9139 = po23  & n9136;
  assign n9140 = ~n8696 & ~n9139;
  assign n9141 = ~n9138 & ~n9140;
  assign n9142 = ~po40  & ~n9125;
  assign n9143 = ~n9133 & n9142;
  assign n9144 = ~n9141 & ~n9143;
  assign n9145 = ~n9135 & ~n9144;
  assign n9146 = po41  & ~n9145;
  assign n9147 = ~n8700 & ~n8708;
  assign n9148 = n8706 & n9147;
  assign n9149 = po23  & n9148;
  assign n9150 = po23  & n9147;
  assign n9151 = ~n8706 & ~n9150;
  assign n9152 = ~n9149 & ~n9151;
  assign n9153 = ~po41  & n9145;
  assign n9154 = ~n9152 & ~n9153;
  assign n9155 = ~n9146 & ~n9154;
  assign n9156 = po42  & ~n9155;
  assign n9157 = ~po42  & ~n9146;
  assign n9158 = ~n9154 & n9157;
  assign n9159 = ~n8711 & ~n8718;
  assign n9160 = n8717 & n9159;
  assign n9161 = po23  & n9160;
  assign n9162 = po23  & n9159;
  assign n9163 = ~n8717 & ~n9162;
  assign n9164 = ~n9161 & ~n9163;
  assign n9165 = ~n9158 & ~n9164;
  assign n9166 = ~n9156 & ~n9165;
  assign n9167 = po43  & ~n9166;
  assign n9168 = ~n8721 & ~n8729;
  assign n9169 = n8727 & n9168;
  assign n9170 = po23  & n9169;
  assign n9171 = po23  & n9168;
  assign n9172 = ~n8727 & ~n9171;
  assign n9173 = ~n9170 & ~n9172;
  assign n9174 = ~po43  & n9166;
  assign n9175 = ~n9173 & ~n9174;
  assign n9176 = ~n9167 & ~n9175;
  assign n9177 = po44  & ~n9176;
  assign n9178 = ~n8732 & ~n8739;
  assign n9179 = n8738 & n9178;
  assign n9180 = po23  & n9179;
  assign n9181 = po23  & n9178;
  assign n9182 = ~n8738 & ~n9181;
  assign n9183 = ~n9180 & ~n9182;
  assign n9184 = ~po44  & ~n9167;
  assign n9185 = ~n9175 & n9184;
  assign n9186 = ~n9183 & ~n9185;
  assign n9187 = ~n9177 & ~n9186;
  assign n9188 = po45  & ~n9187;
  assign n9189 = ~n8742 & ~n8750;
  assign n9190 = n8748 & n9189;
  assign n9191 = po23  & n9190;
  assign n9192 = po23  & n9189;
  assign n9193 = ~n8748 & ~n9192;
  assign n9194 = ~n9191 & ~n9193;
  assign n9195 = ~po45  & n9187;
  assign n9196 = ~n9194 & ~n9195;
  assign n9197 = ~n9188 & ~n9196;
  assign n9198 = po46  & ~n9197;
  assign n9199 = ~n8753 & ~n8760;
  assign n9200 = n8759 & n9199;
  assign n9201 = po23  & n9200;
  assign n9202 = po23  & n9199;
  assign n9203 = ~n8759 & ~n9202;
  assign n9204 = ~n9201 & ~n9203;
  assign n9205 = ~po46  & ~n9188;
  assign n9206 = ~n9196 & n9205;
  assign n9207 = ~n9204 & ~n9206;
  assign n9208 = ~n9198 & ~n9207;
  assign n9209 = po47  & ~n9208;
  assign n9210 = ~n8763 & ~n8771;
  assign n9211 = n8769 & n9210;
  assign n9212 = po23  & n9211;
  assign n9213 = po23  & n9210;
  assign n9214 = ~n8769 & ~n9213;
  assign n9215 = ~n9212 & ~n9214;
  assign n9216 = ~po47  & n9208;
  assign n9217 = ~n9215 & ~n9216;
  assign n9218 = ~n9209 & ~n9217;
  assign n9219 = po48  & ~n9218;
  assign n9220 = ~n8774 & ~n8781;
  assign n9221 = n8780 & n9220;
  assign n9222 = po23  & n9221;
  assign n9223 = po23  & n9220;
  assign n9224 = ~n8780 & ~n9223;
  assign n9225 = ~n9222 & ~n9224;
  assign n9226 = ~po48  & ~n9209;
  assign n9227 = ~n9217 & n9226;
  assign n9228 = ~n9225 & ~n9227;
  assign n9229 = ~n9219 & ~n9228;
  assign n9230 = po49  & ~n9229;
  assign n9231 = ~n8784 & ~n8792;
  assign n9232 = n8790 & n9231;
  assign n9233 = po23  & n9232;
  assign n9234 = po23  & n9231;
  assign n9235 = ~n8790 & ~n9234;
  assign n9236 = ~n9233 & ~n9235;
  assign n9237 = ~po49  & n9229;
  assign n9238 = ~n9236 & ~n9237;
  assign n9239 = ~n9230 & ~n9238;
  assign n9240 = po50  & ~n9239;
  assign n9241 = ~n8795 & ~n8802;
  assign n9242 = n8801 & n9241;
  assign n9243 = po23  & n9242;
  assign n9244 = po23  & n9241;
  assign n9245 = ~n8801 & ~n9244;
  assign n9246 = ~n9243 & ~n9245;
  assign n9247 = ~po50  & ~n9230;
  assign n9248 = ~n9238 & n9247;
  assign n9249 = ~n9246 & ~n9248;
  assign n9250 = ~n9240 & ~n9249;
  assign n9251 = po51  & ~n9250;
  assign n9252 = ~n8805 & ~n8813;
  assign n9253 = n8811 & n9252;
  assign n9254 = po23  & n9253;
  assign n9255 = po23  & n9252;
  assign n9256 = ~n8811 & ~n9255;
  assign n9257 = ~n9254 & ~n9256;
  assign n9258 = ~po51  & n9250;
  assign n9259 = ~n9257 & ~n9258;
  assign n9260 = ~n9251 & ~n9259;
  assign n9261 = po52  & ~n9260;
  assign n9262 = ~n8816 & ~n8823;
  assign n9263 = n8822 & n9262;
  assign n9264 = po23  & n9263;
  assign n9265 = po23  & n9262;
  assign n9266 = ~n8822 & ~n9265;
  assign n9267 = ~n9264 & ~n9266;
  assign n9268 = ~po52  & ~n9251;
  assign n9269 = ~n9259 & n9268;
  assign n9270 = ~n9267 & ~n9269;
  assign n9271 = ~n9261 & ~n9270;
  assign n9272 = po53  & ~n9271;
  assign n9273 = ~n8826 & ~n8834;
  assign n9274 = n8832 & n9273;
  assign n9275 = po23  & n9274;
  assign n9276 = po23  & n9273;
  assign n9277 = ~n8832 & ~n9276;
  assign n9278 = ~n9275 & ~n9277;
  assign n9279 = ~po53  & n9271;
  assign n9280 = ~n9278 & ~n9279;
  assign n9281 = ~n9272 & ~n9280;
  assign n9282 = po54  & ~n9281;
  assign n9283 = ~n8837 & ~n8844;
  assign n9284 = n8843 & n9283;
  assign n9285 = po23  & n9284;
  assign n9286 = po23  & n9283;
  assign n9287 = ~n8843 & ~n9286;
  assign n9288 = ~n9285 & ~n9287;
  assign n9289 = ~po54  & ~n9272;
  assign n9290 = ~n9280 & n9289;
  assign n9291 = ~n9288 & ~n9290;
  assign n9292 = ~n9282 & ~n9291;
  assign n9293 = po55  & ~n9292;
  assign n9294 = ~n8847 & ~n8855;
  assign n9295 = n8853 & n9294;
  assign n9296 = po23  & n9295;
  assign n9297 = po23  & n9294;
  assign n9298 = ~n8853 & ~n9297;
  assign n9299 = ~n9296 & ~n9298;
  assign n9300 = ~po55  & n9292;
  assign n9301 = ~n9299 & ~n9300;
  assign n9302 = ~n9293 & ~n9301;
  assign n9303 = po56  & ~n9302;
  assign n9304 = ~n8858 & ~n8865;
  assign n9305 = n8864 & n9304;
  assign n9306 = po23  & n9305;
  assign n9307 = po23  & n9304;
  assign n9308 = ~n8864 & ~n9307;
  assign n9309 = ~n9306 & ~n9308;
  assign n9310 = ~po56  & ~n9293;
  assign n9311 = ~n9301 & n9310;
  assign n9312 = ~n9309 & ~n9311;
  assign n9313 = ~n9303 & ~n9312;
  assign n9314 = po57  & ~n9313;
  assign n9315 = ~n8868 & ~n8876;
  assign n9316 = n8874 & n9315;
  assign n9317 = po23  & n9316;
  assign n9318 = po23  & n9315;
  assign n9319 = ~n8874 & ~n9318;
  assign n9320 = ~n9317 & ~n9319;
  assign n9321 = ~po57  & n9313;
  assign n9322 = ~n9320 & ~n9321;
  assign n9323 = ~n9314 & ~n9322;
  assign n9324 = po58  & ~n9323;
  assign n9325 = ~n8879 & ~n8886;
  assign n9326 = n8885 & n9325;
  assign n9327 = po23  & n9326;
  assign n9328 = po23  & n9325;
  assign n9329 = ~n8885 & ~n9328;
  assign n9330 = ~n9327 & ~n9329;
  assign n9331 = ~po58  & ~n9314;
  assign n9332 = ~n9322 & n9331;
  assign n9333 = ~n9330 & ~n9332;
  assign n9334 = ~n9324 & ~n9333;
  assign n9335 = po59  & ~n9334;
  assign n9336 = ~n8889 & ~n8897;
  assign n9337 = n8895 & n9336;
  assign n9338 = po23  & n9337;
  assign n9339 = po23  & n9336;
  assign n9340 = ~n8895 & ~n9339;
  assign n9341 = ~n9338 & ~n9340;
  assign n9342 = ~po59  & n9334;
  assign n9343 = ~n9341 & ~n9342;
  assign n9344 = ~n9335 & ~n9343;
  assign n9345 = po60  & ~n9344;
  assign n9346 = ~n8900 & ~n8907;
  assign n9347 = n8906 & n9346;
  assign n9348 = po23  & n9347;
  assign n9349 = po23  & n9346;
  assign n9350 = ~n8906 & ~n9349;
  assign n9351 = ~n9348 & ~n9350;
  assign n9352 = ~po60  & ~n9335;
  assign n9353 = ~n9343 & n9352;
  assign n9354 = ~n9351 & ~n9353;
  assign n9355 = ~n9345 & ~n9354;
  assign n9356 = po61  & ~n9355;
  assign n9357 = ~n8910 & ~n8918;
  assign n9358 = n8916 & n9357;
  assign n9359 = po23  & n9358;
  assign n9360 = po23  & n9357;
  assign n9361 = ~n8916 & ~n9360;
  assign n9362 = ~n9359 & ~n9361;
  assign n9363 = ~po61  & n9355;
  assign n9364 = ~n9362 & ~n9363;
  assign n9365 = ~n9356 & ~n9364;
  assign n9366 = po62  & ~n9365;
  assign n9367 = ~n8921 & ~n8928;
  assign n9368 = n8927 & n9367;
  assign n9369 = po23  & n9368;
  assign n9370 = po23  & n9367;
  assign n9371 = ~n8927 & ~n9370;
  assign n9372 = ~n9369 & ~n9371;
  assign n9373 = ~po62  & ~n9356;
  assign n9374 = ~n9364 & n9373;
  assign n9375 = ~n9372 & ~n9374;
  assign n9376 = ~n9366 & ~n9375;
  assign n9377 = ~n8931 & ~n8939;
  assign n9378 = po23  & n9377;
  assign n9379 = ~n8937 & ~n9378;
  assign n9380 = n8937 & n9378;
  assign n9381 = ~n9379 & ~n9380;
  assign n9382 = ~n8941 & ~n8946;
  assign n9383 = po23  & n9382;
  assign n9384 = ~n8959 & ~n9383;
  assign n9385 = ~n9381 & n9384;
  assign n9386 = ~n9376 & n9385;
  assign n9387 = ~po63  & ~n9386;
  assign n9388 = ~n8946 & po23 ;
  assign n9389 = n8941 & ~n9388;
  assign n9390 = po63  & ~n9382;
  assign n9391 = ~n9389 & n9390;
  assign n9392 = n8946 & ~po23 ;
  assign n9393 = ~n9391 & ~n9392;
  assign n9394 = n9376 & n9381;
  assign n9395 = n9393 & ~n9394;
  assign po22  = n9387 | ~n9395;
  assign n9397 = pi44  & po22 ;
  assign n9398 = ~pi42  & ~pi43 ;
  assign n9399 = ~pi44  & n9398;
  assign n9400 = ~n9397 & ~n9399;
  assign n9401 = po23  & ~n9400;
  assign n9402 = n8958 & ~n9399;
  assign n9403 = ~n8959 & n9402;
  assign n9404 = ~n8952 & n9403;
  assign n9405 = ~n9397 & n9404;
  assign n9406 = ~pi44  & po22 ;
  assign n9407 = pi45  & ~n9406;
  assign n9408 = n8963 & po22 ;
  assign n9409 = ~n9407 & ~n9408;
  assign n9410 = ~n9405 & n9409;
  assign n9411 = ~n9401 & ~n9410;
  assign n9412 = po24  & ~n9411;
  assign n9413 = ~po24  & ~n9401;
  assign n9414 = ~n9410 & n9413;
  assign n9415 = po23  & n9393;
  assign n9416 = ~n9394 & n9415;
  assign n9417 = ~n9387 & n9416;
  assign n9418 = ~n9408 & ~n9417;
  assign n9419 = pi46  & ~n9418;
  assign n9420 = ~pi46  & n9418;
  assign n9421 = ~n9419 & ~n9420;
  assign n9422 = ~n9414 & ~n9421;
  assign n9423 = ~n9412 & ~n9422;
  assign n9424 = po25  & ~n9423;
  assign n9425 = ~n8966 & ~n8970;
  assign n9426 = ~n8974 & n9425;
  assign n9427 = po22  & n9426;
  assign n9428 = po22  & n9425;
  assign n9429 = n8974 & ~n9428;
  assign n9430 = ~n9427 & ~n9429;
  assign n9431 = ~po25  & n9423;
  assign n9432 = ~n9430 & ~n9431;
  assign n9433 = ~n9424 & ~n9432;
  assign n9434 = po26  & ~n9433;
  assign n9435 = ~n8977 & ~n8985;
  assign n9436 = n8984 & n9435;
  assign n9437 = po22  & n9436;
  assign n9438 = po22  & n9435;
  assign n9439 = ~n8984 & ~n9438;
  assign n9440 = ~n9437 & ~n9439;
  assign n9441 = ~po26  & ~n9424;
  assign n9442 = ~n9432 & n9441;
  assign n9443 = ~n9440 & ~n9442;
  assign n9444 = ~n9434 & ~n9443;
  assign n9445 = po27  & ~n9444;
  assign n9446 = ~n8988 & ~n8996;
  assign n9447 = n8994 & n9446;
  assign n9448 = po22  & n9447;
  assign n9449 = po22  & n9446;
  assign n9450 = ~n8994 & ~n9449;
  assign n9451 = ~n9448 & ~n9450;
  assign n9452 = ~po27  & n9444;
  assign n9453 = ~n9451 & ~n9452;
  assign n9454 = ~n9445 & ~n9453;
  assign n9455 = po28  & ~n9454;
  assign n9456 = ~n8999 & ~n9006;
  assign n9457 = n9005 & n9456;
  assign n9458 = po22  & n9457;
  assign n9459 = po22  & n9456;
  assign n9460 = ~n9005 & ~n9459;
  assign n9461 = ~n9458 & ~n9460;
  assign n9462 = ~po28  & ~n9445;
  assign n9463 = ~n9453 & n9462;
  assign n9464 = ~n9461 & ~n9463;
  assign n9465 = ~n9455 & ~n9464;
  assign n9466 = po29  & ~n9465;
  assign n9467 = ~n9009 & ~n9017;
  assign n9468 = n9015 & n9467;
  assign n9469 = po22  & n9468;
  assign n9470 = po22  & n9467;
  assign n9471 = ~n9015 & ~n9470;
  assign n9472 = ~n9469 & ~n9471;
  assign n9473 = ~po29  & n9465;
  assign n9474 = ~n9472 & ~n9473;
  assign n9475 = ~n9466 & ~n9474;
  assign n9476 = po30  & ~n9475;
  assign n9477 = ~n9020 & ~n9027;
  assign n9478 = n9026 & n9477;
  assign n9479 = po22  & n9478;
  assign n9480 = po22  & n9477;
  assign n9481 = ~n9026 & ~n9480;
  assign n9482 = ~n9479 & ~n9481;
  assign n9483 = ~po30  & ~n9466;
  assign n9484 = ~n9474 & n9483;
  assign n9485 = ~n9482 & ~n9484;
  assign n9486 = ~n9476 & ~n9485;
  assign n9487 = po31  & ~n9486;
  assign n9488 = ~n9030 & ~n9038;
  assign n9489 = n9036 & n9488;
  assign n9490 = po22  & n9489;
  assign n9491 = po22  & n9488;
  assign n9492 = ~n9036 & ~n9491;
  assign n9493 = ~n9490 & ~n9492;
  assign n9494 = ~po31  & n9486;
  assign n9495 = ~n9493 & ~n9494;
  assign n9496 = ~n9487 & ~n9495;
  assign n9497 = po32  & ~n9496;
  assign n9498 = ~n9041 & ~n9048;
  assign n9499 = n9047 & n9498;
  assign n9500 = po22  & n9499;
  assign n9501 = po22  & n9498;
  assign n9502 = ~n9047 & ~n9501;
  assign n9503 = ~n9500 & ~n9502;
  assign n9504 = ~po32  & ~n9487;
  assign n9505 = ~n9495 & n9504;
  assign n9506 = ~n9503 & ~n9505;
  assign n9507 = ~n9497 & ~n9506;
  assign n9508 = po33  & ~n9507;
  assign n9509 = ~n9051 & ~n9059;
  assign n9510 = n9057 & n9509;
  assign n9511 = po22  & n9510;
  assign n9512 = po22  & n9509;
  assign n9513 = ~n9057 & ~n9512;
  assign n9514 = ~n9511 & ~n9513;
  assign n9515 = ~po33  & n9507;
  assign n9516 = ~n9514 & ~n9515;
  assign n9517 = ~n9508 & ~n9516;
  assign n9518 = po34  & ~n9517;
  assign n9519 = ~n9062 & ~n9069;
  assign n9520 = n9068 & n9519;
  assign n9521 = po22  & n9520;
  assign n9522 = po22  & n9519;
  assign n9523 = ~n9068 & ~n9522;
  assign n9524 = ~n9521 & ~n9523;
  assign n9525 = ~po34  & ~n9508;
  assign n9526 = ~n9516 & n9525;
  assign n9527 = ~n9524 & ~n9526;
  assign n9528 = ~n9518 & ~n9527;
  assign n9529 = po35  & ~n9528;
  assign n9530 = ~n9072 & ~n9080;
  assign n9531 = n9078 & n9530;
  assign n9532 = po22  & n9531;
  assign n9533 = po22  & n9530;
  assign n9534 = ~n9078 & ~n9533;
  assign n9535 = ~n9532 & ~n9534;
  assign n9536 = ~po35  & n9528;
  assign n9537 = ~n9535 & ~n9536;
  assign n9538 = ~n9529 & ~n9537;
  assign n9539 = po36  & ~n9538;
  assign n9540 = ~n9083 & ~n9090;
  assign n9541 = n9089 & n9540;
  assign n9542 = po22  & n9541;
  assign n9543 = po22  & n9540;
  assign n9544 = ~n9089 & ~n9543;
  assign n9545 = ~n9542 & ~n9544;
  assign n9546 = ~po36  & ~n9529;
  assign n9547 = ~n9537 & n9546;
  assign n9548 = ~n9545 & ~n9547;
  assign n9549 = ~n9539 & ~n9548;
  assign n9550 = po37  & ~n9549;
  assign n9551 = ~n9093 & ~n9101;
  assign n9552 = n9099 & n9551;
  assign n9553 = po22  & n9552;
  assign n9554 = po22  & n9551;
  assign n9555 = ~n9099 & ~n9554;
  assign n9556 = ~n9553 & ~n9555;
  assign n9557 = ~po37  & n9549;
  assign n9558 = ~n9556 & ~n9557;
  assign n9559 = ~n9550 & ~n9558;
  assign n9560 = po38  & ~n9559;
  assign n9561 = ~n9104 & ~n9111;
  assign n9562 = n9110 & n9561;
  assign n9563 = po22  & n9562;
  assign n9564 = po22  & n9561;
  assign n9565 = ~n9110 & ~n9564;
  assign n9566 = ~n9563 & ~n9565;
  assign n9567 = ~po38  & ~n9550;
  assign n9568 = ~n9558 & n9567;
  assign n9569 = ~n9566 & ~n9568;
  assign n9570 = ~n9560 & ~n9569;
  assign n9571 = po39  & ~n9570;
  assign n9572 = ~n9114 & ~n9122;
  assign n9573 = n9120 & n9572;
  assign n9574 = po22  & n9573;
  assign n9575 = po22  & n9572;
  assign n9576 = ~n9120 & ~n9575;
  assign n9577 = ~n9574 & ~n9576;
  assign n9578 = ~po39  & n9570;
  assign n9579 = ~n9577 & ~n9578;
  assign n9580 = ~n9571 & ~n9579;
  assign n9581 = po40  & ~n9580;
  assign n9582 = ~n9125 & ~n9132;
  assign n9583 = n9131 & n9582;
  assign n9584 = po22  & n9583;
  assign n9585 = po22  & n9582;
  assign n9586 = ~n9131 & ~n9585;
  assign n9587 = ~n9584 & ~n9586;
  assign n9588 = ~po40  & ~n9571;
  assign n9589 = ~n9579 & n9588;
  assign n9590 = ~n9587 & ~n9589;
  assign n9591 = ~n9581 & ~n9590;
  assign n9592 = po41  & ~n9591;
  assign n9593 = ~n9135 & ~n9143;
  assign n9594 = n9141 & n9593;
  assign n9595 = po22  & n9594;
  assign n9596 = po22  & n9593;
  assign n9597 = ~n9141 & ~n9596;
  assign n9598 = ~n9595 & ~n9597;
  assign n9599 = ~po41  & n9591;
  assign n9600 = ~n9598 & ~n9599;
  assign n9601 = ~n9592 & ~n9600;
  assign n9602 = po42  & ~n9601;
  assign n9603 = ~n9146 & ~n9153;
  assign n9604 = n9152 & n9603;
  assign n9605 = po22  & n9604;
  assign n9606 = po22  & n9603;
  assign n9607 = ~n9152 & ~n9606;
  assign n9608 = ~n9605 & ~n9607;
  assign n9609 = ~po42  & ~n9592;
  assign n9610 = ~n9600 & n9609;
  assign n9611 = ~n9608 & ~n9610;
  assign n9612 = ~n9602 & ~n9611;
  assign n9613 = po43  & ~n9612;
  assign n9614 = ~n9156 & ~n9158;
  assign n9615 = n9164 & n9614;
  assign n9616 = po22  & n9615;
  assign n9617 = po22  & n9614;
  assign n9618 = ~n9164 & ~n9617;
  assign n9619 = ~n9616 & ~n9618;
  assign n9620 = ~po43  & n9612;
  assign n9621 = ~n9619 & ~n9620;
  assign n9622 = ~n9613 & ~n9621;
  assign n9623 = po44  & ~n9622;
  assign n9624 = ~n9167 & ~n9174;
  assign n9625 = n9173 & n9624;
  assign n9626 = po22  & n9625;
  assign n9627 = po22  & n9624;
  assign n9628 = ~n9173 & ~n9627;
  assign n9629 = ~n9626 & ~n9628;
  assign n9630 = ~po44  & ~n9613;
  assign n9631 = ~n9621 & n9630;
  assign n9632 = ~n9629 & ~n9631;
  assign n9633 = ~n9623 & ~n9632;
  assign n9634 = po45  & ~n9633;
  assign n9635 = ~n9177 & ~n9185;
  assign n9636 = n9183 & n9635;
  assign n9637 = po22  & n9636;
  assign n9638 = po22  & n9635;
  assign n9639 = ~n9183 & ~n9638;
  assign n9640 = ~n9637 & ~n9639;
  assign n9641 = ~po45  & n9633;
  assign n9642 = ~n9640 & ~n9641;
  assign n9643 = ~n9634 & ~n9642;
  assign n9644 = po46  & ~n9643;
  assign n9645 = ~n9188 & ~n9195;
  assign n9646 = n9194 & n9645;
  assign n9647 = po22  & n9646;
  assign n9648 = po22  & n9645;
  assign n9649 = ~n9194 & ~n9648;
  assign n9650 = ~n9647 & ~n9649;
  assign n9651 = ~po46  & ~n9634;
  assign n9652 = ~n9642 & n9651;
  assign n9653 = ~n9650 & ~n9652;
  assign n9654 = ~n9644 & ~n9653;
  assign n9655 = po47  & ~n9654;
  assign n9656 = ~n9198 & ~n9206;
  assign n9657 = n9204 & n9656;
  assign n9658 = po22  & n9657;
  assign n9659 = po22  & n9656;
  assign n9660 = ~n9204 & ~n9659;
  assign n9661 = ~n9658 & ~n9660;
  assign n9662 = ~po47  & n9654;
  assign n9663 = ~n9661 & ~n9662;
  assign n9664 = ~n9655 & ~n9663;
  assign n9665 = po48  & ~n9664;
  assign n9666 = ~n9209 & ~n9216;
  assign n9667 = n9215 & n9666;
  assign n9668 = po22  & n9667;
  assign n9669 = po22  & n9666;
  assign n9670 = ~n9215 & ~n9669;
  assign n9671 = ~n9668 & ~n9670;
  assign n9672 = ~po48  & ~n9655;
  assign n9673 = ~n9663 & n9672;
  assign n9674 = ~n9671 & ~n9673;
  assign n9675 = ~n9665 & ~n9674;
  assign n9676 = po49  & ~n9675;
  assign n9677 = ~n9219 & ~n9227;
  assign n9678 = n9225 & n9677;
  assign n9679 = po22  & n9678;
  assign n9680 = po22  & n9677;
  assign n9681 = ~n9225 & ~n9680;
  assign n9682 = ~n9679 & ~n9681;
  assign n9683 = ~po49  & n9675;
  assign n9684 = ~n9682 & ~n9683;
  assign n9685 = ~n9676 & ~n9684;
  assign n9686 = po50  & ~n9685;
  assign n9687 = ~n9230 & ~n9237;
  assign n9688 = n9236 & n9687;
  assign n9689 = po22  & n9688;
  assign n9690 = po22  & n9687;
  assign n9691 = ~n9236 & ~n9690;
  assign n9692 = ~n9689 & ~n9691;
  assign n9693 = ~po50  & ~n9676;
  assign n9694 = ~n9684 & n9693;
  assign n9695 = ~n9692 & ~n9694;
  assign n9696 = ~n9686 & ~n9695;
  assign n9697 = po51  & ~n9696;
  assign n9698 = ~n9240 & ~n9248;
  assign n9699 = n9246 & n9698;
  assign n9700 = po22  & n9699;
  assign n9701 = po22  & n9698;
  assign n9702 = ~n9246 & ~n9701;
  assign n9703 = ~n9700 & ~n9702;
  assign n9704 = ~po51  & n9696;
  assign n9705 = ~n9703 & ~n9704;
  assign n9706 = ~n9697 & ~n9705;
  assign n9707 = po52  & ~n9706;
  assign n9708 = ~n9251 & ~n9258;
  assign n9709 = n9257 & n9708;
  assign n9710 = po22  & n9709;
  assign n9711 = po22  & n9708;
  assign n9712 = ~n9257 & ~n9711;
  assign n9713 = ~n9710 & ~n9712;
  assign n9714 = ~po52  & ~n9697;
  assign n9715 = ~n9705 & n9714;
  assign n9716 = ~n9713 & ~n9715;
  assign n9717 = ~n9707 & ~n9716;
  assign n9718 = po53  & ~n9717;
  assign n9719 = ~n9261 & ~n9269;
  assign n9720 = n9267 & n9719;
  assign n9721 = po22  & n9720;
  assign n9722 = po22  & n9719;
  assign n9723 = ~n9267 & ~n9722;
  assign n9724 = ~n9721 & ~n9723;
  assign n9725 = ~po53  & n9717;
  assign n9726 = ~n9724 & ~n9725;
  assign n9727 = ~n9718 & ~n9726;
  assign n9728 = po54  & ~n9727;
  assign n9729 = ~n9272 & ~n9279;
  assign n9730 = n9278 & n9729;
  assign n9731 = po22  & n9730;
  assign n9732 = po22  & n9729;
  assign n9733 = ~n9278 & ~n9732;
  assign n9734 = ~n9731 & ~n9733;
  assign n9735 = ~po54  & ~n9718;
  assign n9736 = ~n9726 & n9735;
  assign n9737 = ~n9734 & ~n9736;
  assign n9738 = ~n9728 & ~n9737;
  assign n9739 = po55  & ~n9738;
  assign n9740 = ~n9282 & ~n9290;
  assign n9741 = n9288 & n9740;
  assign n9742 = po22  & n9741;
  assign n9743 = po22  & n9740;
  assign n9744 = ~n9288 & ~n9743;
  assign n9745 = ~n9742 & ~n9744;
  assign n9746 = ~po55  & n9738;
  assign n9747 = ~n9745 & ~n9746;
  assign n9748 = ~n9739 & ~n9747;
  assign n9749 = po56  & ~n9748;
  assign n9750 = ~n9293 & ~n9300;
  assign n9751 = n9299 & n9750;
  assign n9752 = po22  & n9751;
  assign n9753 = po22  & n9750;
  assign n9754 = ~n9299 & ~n9753;
  assign n9755 = ~n9752 & ~n9754;
  assign n9756 = ~po56  & ~n9739;
  assign n9757 = ~n9747 & n9756;
  assign n9758 = ~n9755 & ~n9757;
  assign n9759 = ~n9749 & ~n9758;
  assign n9760 = po57  & ~n9759;
  assign n9761 = ~n9303 & ~n9311;
  assign n9762 = n9309 & n9761;
  assign n9763 = po22  & n9762;
  assign n9764 = po22  & n9761;
  assign n9765 = ~n9309 & ~n9764;
  assign n9766 = ~n9763 & ~n9765;
  assign n9767 = ~po57  & n9759;
  assign n9768 = ~n9766 & ~n9767;
  assign n9769 = ~n9760 & ~n9768;
  assign n9770 = po58  & ~n9769;
  assign n9771 = ~n9314 & ~n9321;
  assign n9772 = n9320 & n9771;
  assign n9773 = po22  & n9772;
  assign n9774 = po22  & n9771;
  assign n9775 = ~n9320 & ~n9774;
  assign n9776 = ~n9773 & ~n9775;
  assign n9777 = ~po58  & ~n9760;
  assign n9778 = ~n9768 & n9777;
  assign n9779 = ~n9776 & ~n9778;
  assign n9780 = ~n9770 & ~n9779;
  assign n9781 = po59  & ~n9780;
  assign n9782 = ~n9324 & ~n9332;
  assign n9783 = n9330 & n9782;
  assign n9784 = po22  & n9783;
  assign n9785 = po22  & n9782;
  assign n9786 = ~n9330 & ~n9785;
  assign n9787 = ~n9784 & ~n9786;
  assign n9788 = ~po59  & n9780;
  assign n9789 = ~n9787 & ~n9788;
  assign n9790 = ~n9781 & ~n9789;
  assign n9791 = po60  & ~n9790;
  assign n9792 = ~n9335 & ~n9342;
  assign n9793 = n9341 & n9792;
  assign n9794 = po22  & n9793;
  assign n9795 = po22  & n9792;
  assign n9796 = ~n9341 & ~n9795;
  assign n9797 = ~n9794 & ~n9796;
  assign n9798 = ~po60  & ~n9781;
  assign n9799 = ~n9789 & n9798;
  assign n9800 = ~n9797 & ~n9799;
  assign n9801 = ~n9791 & ~n9800;
  assign n9802 = po61  & ~n9801;
  assign n9803 = ~n9345 & ~n9353;
  assign n9804 = n9351 & n9803;
  assign n9805 = po22  & n9804;
  assign n9806 = po22  & n9803;
  assign n9807 = ~n9351 & ~n9806;
  assign n9808 = ~n9805 & ~n9807;
  assign n9809 = ~po61  & n9801;
  assign n9810 = ~n9808 & ~n9809;
  assign n9811 = ~n9802 & ~n9810;
  assign n9812 = po62  & ~n9811;
  assign n9813 = ~n9356 & ~n9363;
  assign n9814 = n9362 & n9813;
  assign n9815 = po22  & n9814;
  assign n9816 = po22  & n9813;
  assign n9817 = ~n9362 & ~n9816;
  assign n9818 = ~n9815 & ~n9817;
  assign n9819 = ~po62  & ~n9802;
  assign n9820 = ~n9810 & n9819;
  assign n9821 = ~n9818 & ~n9820;
  assign n9822 = ~n9812 & ~n9821;
  assign n9823 = ~n9366 & ~n9374;
  assign n9824 = po22  & n9823;
  assign n9825 = ~n9372 & ~n9824;
  assign n9826 = n9372 & n9824;
  assign n9827 = ~n9825 & ~n9826;
  assign n9828 = ~n9376 & ~n9381;
  assign n9829 = po22  & n9828;
  assign n9830 = ~n9394 & ~n9829;
  assign n9831 = ~n9827 & n9830;
  assign n9832 = ~n9822 & n9831;
  assign n9833 = ~po63  & ~n9832;
  assign n9834 = ~n9381 & po22 ;
  assign n9835 = n9376 & ~n9834;
  assign n9836 = po63  & ~n9828;
  assign n9837 = ~n9835 & n9836;
  assign n9838 = n9381 & ~po22 ;
  assign n9839 = ~n9837 & ~n9838;
  assign n9840 = n9822 & n9827;
  assign n9841 = n9839 & ~n9840;
  assign po21  = n9833 | ~n9841;
  assign n9843 = pi42  & po21 ;
  assign n9844 = ~pi40  & ~pi41 ;
  assign n9845 = ~pi42  & n9844;
  assign n9846 = ~n9843 & ~n9845;
  assign n9847 = po22  & ~n9846;
  assign n9848 = n9393 & ~n9845;
  assign n9849 = ~n9394 & n9848;
  assign n9850 = ~n9387 & n9849;
  assign n9851 = ~n9843 & n9850;
  assign n9852 = ~pi42  & po21 ;
  assign n9853 = pi43  & ~n9852;
  assign n9854 = n9398 & po21 ;
  assign n9855 = ~n9853 & ~n9854;
  assign n9856 = ~n9851 & n9855;
  assign n9857 = ~n9847 & ~n9856;
  assign n9858 = po23  & ~n9857;
  assign n9859 = po22  & n9839;
  assign n9860 = ~n9840 & n9859;
  assign n9861 = ~n9833 & n9860;
  assign n9862 = ~n9854 & ~n9861;
  assign n9863 = pi44  & ~n9862;
  assign n9864 = ~pi44  & n9862;
  assign n9865 = ~n9863 & ~n9864;
  assign n9866 = ~po23  & n9857;
  assign n9867 = ~n9865 & ~n9866;
  assign n9868 = ~n9858 & ~n9867;
  assign n9869 = po24  & ~n9868;
  assign n9870 = ~n9401 & ~n9405;
  assign n9871 = ~n9409 & n9870;
  assign n9872 = po21  & n9871;
  assign n9873 = po21  & n9870;
  assign n9874 = n9409 & ~n9873;
  assign n9875 = ~n9872 & ~n9874;
  assign n9876 = ~po24  & ~n9858;
  assign n9877 = ~n9867 & n9876;
  assign n9878 = ~n9875 & ~n9877;
  assign n9879 = ~n9869 & ~n9878;
  assign n9880 = po25  & ~n9879;
  assign n9881 = ~n9412 & ~n9414;
  assign n9882 = n9421 & n9881;
  assign n9883 = po21  & n9882;
  assign n9884 = po21  & n9881;
  assign n9885 = ~n9421 & ~n9884;
  assign n9886 = ~n9883 & ~n9885;
  assign n9887 = ~po25  & n9879;
  assign n9888 = ~n9886 & ~n9887;
  assign n9889 = ~n9880 & ~n9888;
  assign n9890 = po26  & ~n9889;
  assign n9891 = ~n9424 & ~n9431;
  assign n9892 = n9430 & n9891;
  assign n9893 = po21  & n9892;
  assign n9894 = po21  & n9891;
  assign n9895 = ~n9430 & ~n9894;
  assign n9896 = ~n9893 & ~n9895;
  assign n9897 = ~po26  & ~n9880;
  assign n9898 = ~n9888 & n9897;
  assign n9899 = ~n9896 & ~n9898;
  assign n9900 = ~n9890 & ~n9899;
  assign n9901 = po27  & ~n9900;
  assign n9902 = ~n9434 & ~n9442;
  assign n9903 = n9440 & n9902;
  assign n9904 = po21  & n9903;
  assign n9905 = po21  & n9902;
  assign n9906 = ~n9440 & ~n9905;
  assign n9907 = ~n9904 & ~n9906;
  assign n9908 = ~po27  & n9900;
  assign n9909 = ~n9907 & ~n9908;
  assign n9910 = ~n9901 & ~n9909;
  assign n9911 = po28  & ~n9910;
  assign n9912 = ~n9445 & ~n9452;
  assign n9913 = n9451 & n9912;
  assign n9914 = po21  & n9913;
  assign n9915 = po21  & n9912;
  assign n9916 = ~n9451 & ~n9915;
  assign n9917 = ~n9914 & ~n9916;
  assign n9918 = ~po28  & ~n9901;
  assign n9919 = ~n9909 & n9918;
  assign n9920 = ~n9917 & ~n9919;
  assign n9921 = ~n9911 & ~n9920;
  assign n9922 = po29  & ~n9921;
  assign n9923 = ~n9455 & ~n9463;
  assign n9924 = n9461 & n9923;
  assign n9925 = po21  & n9924;
  assign n9926 = po21  & n9923;
  assign n9927 = ~n9461 & ~n9926;
  assign n9928 = ~n9925 & ~n9927;
  assign n9929 = ~po29  & n9921;
  assign n9930 = ~n9928 & ~n9929;
  assign n9931 = ~n9922 & ~n9930;
  assign n9932 = po30  & ~n9931;
  assign n9933 = ~n9466 & ~n9473;
  assign n9934 = n9472 & n9933;
  assign n9935 = po21  & n9934;
  assign n9936 = po21  & n9933;
  assign n9937 = ~n9472 & ~n9936;
  assign n9938 = ~n9935 & ~n9937;
  assign n9939 = ~po30  & ~n9922;
  assign n9940 = ~n9930 & n9939;
  assign n9941 = ~n9938 & ~n9940;
  assign n9942 = ~n9932 & ~n9941;
  assign n9943 = po31  & ~n9942;
  assign n9944 = ~n9476 & ~n9484;
  assign n9945 = n9482 & n9944;
  assign n9946 = po21  & n9945;
  assign n9947 = po21  & n9944;
  assign n9948 = ~n9482 & ~n9947;
  assign n9949 = ~n9946 & ~n9948;
  assign n9950 = ~po31  & n9942;
  assign n9951 = ~n9949 & ~n9950;
  assign n9952 = ~n9943 & ~n9951;
  assign n9953 = po32  & ~n9952;
  assign n9954 = ~n9487 & ~n9494;
  assign n9955 = n9493 & n9954;
  assign n9956 = po21  & n9955;
  assign n9957 = po21  & n9954;
  assign n9958 = ~n9493 & ~n9957;
  assign n9959 = ~n9956 & ~n9958;
  assign n9960 = ~po32  & ~n9943;
  assign n9961 = ~n9951 & n9960;
  assign n9962 = ~n9959 & ~n9961;
  assign n9963 = ~n9953 & ~n9962;
  assign n9964 = po33  & ~n9963;
  assign n9965 = ~n9497 & ~n9505;
  assign n9966 = n9503 & n9965;
  assign n9967 = po21  & n9966;
  assign n9968 = po21  & n9965;
  assign n9969 = ~n9503 & ~n9968;
  assign n9970 = ~n9967 & ~n9969;
  assign n9971 = ~po33  & n9963;
  assign n9972 = ~n9970 & ~n9971;
  assign n9973 = ~n9964 & ~n9972;
  assign n9974 = po34  & ~n9973;
  assign n9975 = ~n9508 & ~n9515;
  assign n9976 = n9514 & n9975;
  assign n9977 = po21  & n9976;
  assign n9978 = po21  & n9975;
  assign n9979 = ~n9514 & ~n9978;
  assign n9980 = ~n9977 & ~n9979;
  assign n9981 = ~po34  & ~n9964;
  assign n9982 = ~n9972 & n9981;
  assign n9983 = ~n9980 & ~n9982;
  assign n9984 = ~n9974 & ~n9983;
  assign n9985 = po35  & ~n9984;
  assign n9986 = ~n9518 & ~n9526;
  assign n9987 = n9524 & n9986;
  assign n9988 = po21  & n9987;
  assign n9989 = po21  & n9986;
  assign n9990 = ~n9524 & ~n9989;
  assign n9991 = ~n9988 & ~n9990;
  assign n9992 = ~po35  & n9984;
  assign n9993 = ~n9991 & ~n9992;
  assign n9994 = ~n9985 & ~n9993;
  assign n9995 = po36  & ~n9994;
  assign n9996 = ~n9529 & ~n9536;
  assign n9997 = n9535 & n9996;
  assign n9998 = po21  & n9997;
  assign n9999 = po21  & n9996;
  assign n10000 = ~n9535 & ~n9999;
  assign n10001 = ~n9998 & ~n10000;
  assign n10002 = ~po36  & ~n9985;
  assign n10003 = ~n9993 & n10002;
  assign n10004 = ~n10001 & ~n10003;
  assign n10005 = ~n9995 & ~n10004;
  assign n10006 = po37  & ~n10005;
  assign n10007 = ~n9539 & ~n9547;
  assign n10008 = n9545 & n10007;
  assign n10009 = po21  & n10008;
  assign n10010 = po21  & n10007;
  assign n10011 = ~n9545 & ~n10010;
  assign n10012 = ~n10009 & ~n10011;
  assign n10013 = ~po37  & n10005;
  assign n10014 = ~n10012 & ~n10013;
  assign n10015 = ~n10006 & ~n10014;
  assign n10016 = po38  & ~n10015;
  assign n10017 = ~n9550 & ~n9557;
  assign n10018 = n9556 & n10017;
  assign n10019 = po21  & n10018;
  assign n10020 = po21  & n10017;
  assign n10021 = ~n9556 & ~n10020;
  assign n10022 = ~n10019 & ~n10021;
  assign n10023 = ~po38  & ~n10006;
  assign n10024 = ~n10014 & n10023;
  assign n10025 = ~n10022 & ~n10024;
  assign n10026 = ~n10016 & ~n10025;
  assign n10027 = po39  & ~n10026;
  assign n10028 = ~n9560 & ~n9568;
  assign n10029 = n9566 & n10028;
  assign n10030 = po21  & n10029;
  assign n10031 = po21  & n10028;
  assign n10032 = ~n9566 & ~n10031;
  assign n10033 = ~n10030 & ~n10032;
  assign n10034 = ~po39  & n10026;
  assign n10035 = ~n10033 & ~n10034;
  assign n10036 = ~n10027 & ~n10035;
  assign n10037 = po40  & ~n10036;
  assign n10038 = ~n9571 & ~n9578;
  assign n10039 = n9577 & n10038;
  assign n10040 = po21  & n10039;
  assign n10041 = po21  & n10038;
  assign n10042 = ~n9577 & ~n10041;
  assign n10043 = ~n10040 & ~n10042;
  assign n10044 = ~po40  & ~n10027;
  assign n10045 = ~n10035 & n10044;
  assign n10046 = ~n10043 & ~n10045;
  assign n10047 = ~n10037 & ~n10046;
  assign n10048 = po41  & ~n10047;
  assign n10049 = ~n9581 & ~n9589;
  assign n10050 = n9587 & n10049;
  assign n10051 = po21  & n10050;
  assign n10052 = po21  & n10049;
  assign n10053 = ~n9587 & ~n10052;
  assign n10054 = ~n10051 & ~n10053;
  assign n10055 = ~po41  & n10047;
  assign n10056 = ~n10054 & ~n10055;
  assign n10057 = ~n10048 & ~n10056;
  assign n10058 = po42  & ~n10057;
  assign n10059 = ~n9592 & ~n9599;
  assign n10060 = n9598 & n10059;
  assign n10061 = po21  & n10060;
  assign n10062 = po21  & n10059;
  assign n10063 = ~n9598 & ~n10062;
  assign n10064 = ~n10061 & ~n10063;
  assign n10065 = ~po42  & ~n10048;
  assign n10066 = ~n10056 & n10065;
  assign n10067 = ~n10064 & ~n10066;
  assign n10068 = ~n10058 & ~n10067;
  assign n10069 = po43  & ~n10068;
  assign n10070 = ~n9602 & ~n9610;
  assign n10071 = n9608 & n10070;
  assign n10072 = po21  & n10071;
  assign n10073 = po21  & n10070;
  assign n10074 = ~n9608 & ~n10073;
  assign n10075 = ~n10072 & ~n10074;
  assign n10076 = ~po43  & n10068;
  assign n10077 = ~n10075 & ~n10076;
  assign n10078 = ~n10069 & ~n10077;
  assign n10079 = po44  & ~n10078;
  assign n10080 = ~po44  & ~n10069;
  assign n10081 = ~n10077 & n10080;
  assign n10082 = ~n9613 & ~n9620;
  assign n10083 = n9619 & n10082;
  assign n10084 = po21  & n10083;
  assign n10085 = po21  & n10082;
  assign n10086 = ~n9619 & ~n10085;
  assign n10087 = ~n10084 & ~n10086;
  assign n10088 = ~n10081 & ~n10087;
  assign n10089 = ~n10079 & ~n10088;
  assign n10090 = po45  & ~n10089;
  assign n10091 = ~n9623 & ~n9631;
  assign n10092 = n9629 & n10091;
  assign n10093 = po21  & n10092;
  assign n10094 = po21  & n10091;
  assign n10095 = ~n9629 & ~n10094;
  assign n10096 = ~n10093 & ~n10095;
  assign n10097 = ~po45  & n10089;
  assign n10098 = ~n10096 & ~n10097;
  assign n10099 = ~n10090 & ~n10098;
  assign n10100 = po46  & ~n10099;
  assign n10101 = ~n9634 & ~n9641;
  assign n10102 = n9640 & n10101;
  assign n10103 = po21  & n10102;
  assign n10104 = po21  & n10101;
  assign n10105 = ~n9640 & ~n10104;
  assign n10106 = ~n10103 & ~n10105;
  assign n10107 = ~po46  & ~n10090;
  assign n10108 = ~n10098 & n10107;
  assign n10109 = ~n10106 & ~n10108;
  assign n10110 = ~n10100 & ~n10109;
  assign n10111 = po47  & ~n10110;
  assign n10112 = ~n9644 & ~n9652;
  assign n10113 = n9650 & n10112;
  assign n10114 = po21  & n10113;
  assign n10115 = po21  & n10112;
  assign n10116 = ~n9650 & ~n10115;
  assign n10117 = ~n10114 & ~n10116;
  assign n10118 = ~po47  & n10110;
  assign n10119 = ~n10117 & ~n10118;
  assign n10120 = ~n10111 & ~n10119;
  assign n10121 = po48  & ~n10120;
  assign n10122 = ~n9655 & ~n9662;
  assign n10123 = n9661 & n10122;
  assign n10124 = po21  & n10123;
  assign n10125 = po21  & n10122;
  assign n10126 = ~n9661 & ~n10125;
  assign n10127 = ~n10124 & ~n10126;
  assign n10128 = ~po48  & ~n10111;
  assign n10129 = ~n10119 & n10128;
  assign n10130 = ~n10127 & ~n10129;
  assign n10131 = ~n10121 & ~n10130;
  assign n10132 = po49  & ~n10131;
  assign n10133 = ~n9665 & ~n9673;
  assign n10134 = n9671 & n10133;
  assign n10135 = po21  & n10134;
  assign n10136 = po21  & n10133;
  assign n10137 = ~n9671 & ~n10136;
  assign n10138 = ~n10135 & ~n10137;
  assign n10139 = ~po49  & n10131;
  assign n10140 = ~n10138 & ~n10139;
  assign n10141 = ~n10132 & ~n10140;
  assign n10142 = po50  & ~n10141;
  assign n10143 = ~n9676 & ~n9683;
  assign n10144 = n9682 & n10143;
  assign n10145 = po21  & n10144;
  assign n10146 = po21  & n10143;
  assign n10147 = ~n9682 & ~n10146;
  assign n10148 = ~n10145 & ~n10147;
  assign n10149 = ~po50  & ~n10132;
  assign n10150 = ~n10140 & n10149;
  assign n10151 = ~n10148 & ~n10150;
  assign n10152 = ~n10142 & ~n10151;
  assign n10153 = po51  & ~n10152;
  assign n10154 = ~n9686 & ~n9694;
  assign n10155 = n9692 & n10154;
  assign n10156 = po21  & n10155;
  assign n10157 = po21  & n10154;
  assign n10158 = ~n9692 & ~n10157;
  assign n10159 = ~n10156 & ~n10158;
  assign n10160 = ~po51  & n10152;
  assign n10161 = ~n10159 & ~n10160;
  assign n10162 = ~n10153 & ~n10161;
  assign n10163 = po52  & ~n10162;
  assign n10164 = ~n9697 & ~n9704;
  assign n10165 = n9703 & n10164;
  assign n10166 = po21  & n10165;
  assign n10167 = po21  & n10164;
  assign n10168 = ~n9703 & ~n10167;
  assign n10169 = ~n10166 & ~n10168;
  assign n10170 = ~po52  & ~n10153;
  assign n10171 = ~n10161 & n10170;
  assign n10172 = ~n10169 & ~n10171;
  assign n10173 = ~n10163 & ~n10172;
  assign n10174 = po53  & ~n10173;
  assign n10175 = ~n9707 & ~n9715;
  assign n10176 = n9713 & n10175;
  assign n10177 = po21  & n10176;
  assign n10178 = po21  & n10175;
  assign n10179 = ~n9713 & ~n10178;
  assign n10180 = ~n10177 & ~n10179;
  assign n10181 = ~po53  & n10173;
  assign n10182 = ~n10180 & ~n10181;
  assign n10183 = ~n10174 & ~n10182;
  assign n10184 = po54  & ~n10183;
  assign n10185 = ~n9718 & ~n9725;
  assign n10186 = n9724 & n10185;
  assign n10187 = po21  & n10186;
  assign n10188 = po21  & n10185;
  assign n10189 = ~n9724 & ~n10188;
  assign n10190 = ~n10187 & ~n10189;
  assign n10191 = ~po54  & ~n10174;
  assign n10192 = ~n10182 & n10191;
  assign n10193 = ~n10190 & ~n10192;
  assign n10194 = ~n10184 & ~n10193;
  assign n10195 = po55  & ~n10194;
  assign n10196 = ~n9728 & ~n9736;
  assign n10197 = n9734 & n10196;
  assign n10198 = po21  & n10197;
  assign n10199 = po21  & n10196;
  assign n10200 = ~n9734 & ~n10199;
  assign n10201 = ~n10198 & ~n10200;
  assign n10202 = ~po55  & n10194;
  assign n10203 = ~n10201 & ~n10202;
  assign n10204 = ~n10195 & ~n10203;
  assign n10205 = po56  & ~n10204;
  assign n10206 = ~n9739 & ~n9746;
  assign n10207 = n9745 & n10206;
  assign n10208 = po21  & n10207;
  assign n10209 = po21  & n10206;
  assign n10210 = ~n9745 & ~n10209;
  assign n10211 = ~n10208 & ~n10210;
  assign n10212 = ~po56  & ~n10195;
  assign n10213 = ~n10203 & n10212;
  assign n10214 = ~n10211 & ~n10213;
  assign n10215 = ~n10205 & ~n10214;
  assign n10216 = po57  & ~n10215;
  assign n10217 = ~n9749 & ~n9757;
  assign n10218 = n9755 & n10217;
  assign n10219 = po21  & n10218;
  assign n10220 = po21  & n10217;
  assign n10221 = ~n9755 & ~n10220;
  assign n10222 = ~n10219 & ~n10221;
  assign n10223 = ~po57  & n10215;
  assign n10224 = ~n10222 & ~n10223;
  assign n10225 = ~n10216 & ~n10224;
  assign n10226 = po58  & ~n10225;
  assign n10227 = ~n9760 & ~n9767;
  assign n10228 = n9766 & n10227;
  assign n10229 = po21  & n10228;
  assign n10230 = po21  & n10227;
  assign n10231 = ~n9766 & ~n10230;
  assign n10232 = ~n10229 & ~n10231;
  assign n10233 = ~po58  & ~n10216;
  assign n10234 = ~n10224 & n10233;
  assign n10235 = ~n10232 & ~n10234;
  assign n10236 = ~n10226 & ~n10235;
  assign n10237 = po59  & ~n10236;
  assign n10238 = ~n9770 & ~n9778;
  assign n10239 = n9776 & n10238;
  assign n10240 = po21  & n10239;
  assign n10241 = po21  & n10238;
  assign n10242 = ~n9776 & ~n10241;
  assign n10243 = ~n10240 & ~n10242;
  assign n10244 = ~po59  & n10236;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = ~n10237 & ~n10245;
  assign n10247 = po60  & ~n10246;
  assign n10248 = ~n9781 & ~n9788;
  assign n10249 = n9787 & n10248;
  assign n10250 = po21  & n10249;
  assign n10251 = po21  & n10248;
  assign n10252 = ~n9787 & ~n10251;
  assign n10253 = ~n10250 & ~n10252;
  assign n10254 = ~po60  & ~n10237;
  assign n10255 = ~n10245 & n10254;
  assign n10256 = ~n10253 & ~n10255;
  assign n10257 = ~n10247 & ~n10256;
  assign n10258 = po61  & ~n10257;
  assign n10259 = ~n9791 & ~n9799;
  assign n10260 = n9797 & n10259;
  assign n10261 = po21  & n10260;
  assign n10262 = po21  & n10259;
  assign n10263 = ~n9797 & ~n10262;
  assign n10264 = ~n10261 & ~n10263;
  assign n10265 = ~po61  & n10257;
  assign n10266 = ~n10264 & ~n10265;
  assign n10267 = ~n10258 & ~n10266;
  assign n10268 = po62  & ~n10267;
  assign n10269 = ~n9802 & ~n9809;
  assign n10270 = n9808 & n10269;
  assign n10271 = po21  & n10270;
  assign n10272 = po21  & n10269;
  assign n10273 = ~n9808 & ~n10272;
  assign n10274 = ~n10271 & ~n10273;
  assign n10275 = ~po62  & ~n10258;
  assign n10276 = ~n10266 & n10275;
  assign n10277 = ~n10274 & ~n10276;
  assign n10278 = ~n10268 & ~n10277;
  assign n10279 = ~n9812 & ~n9820;
  assign n10280 = po21  & n10279;
  assign n10281 = ~n9818 & ~n10280;
  assign n10282 = n9818 & n10280;
  assign n10283 = ~n10281 & ~n10282;
  assign n10284 = ~n9822 & ~n9827;
  assign n10285 = po21  & n10284;
  assign n10286 = ~n9840 & ~n10285;
  assign n10287 = ~n10283 & n10286;
  assign n10288 = ~n10278 & n10287;
  assign n10289 = ~po63  & ~n10288;
  assign n10290 = ~n9827 & po21 ;
  assign n10291 = n9822 & ~n10290;
  assign n10292 = po63  & ~n10284;
  assign n10293 = ~n10291 & n10292;
  assign n10294 = n9827 & ~po21 ;
  assign n10295 = ~n10293 & ~n10294;
  assign n10296 = n10278 & n10283;
  assign n10297 = n10295 & ~n10296;
  assign po20  = n10289 | ~n10297;
  assign n10299 = pi40  & po20 ;
  assign n10300 = ~pi38  & ~pi39 ;
  assign n10301 = ~pi40  & n10300;
  assign n10302 = ~n10299 & ~n10301;
  assign n10303 = po21  & ~n10302;
  assign n10304 = n9839 & ~n10301;
  assign n10305 = ~n9840 & n10304;
  assign n10306 = ~n9833 & n10305;
  assign n10307 = ~n10299 & n10306;
  assign n10308 = ~pi40  & po20 ;
  assign n10309 = pi41  & ~n10308;
  assign n10310 = n9844 & po20 ;
  assign n10311 = ~n10309 & ~n10310;
  assign n10312 = ~n10307 & n10311;
  assign n10313 = ~n10303 & ~n10312;
  assign n10314 = po22  & ~n10313;
  assign n10315 = ~po22  & ~n10303;
  assign n10316 = ~n10312 & n10315;
  assign n10317 = po21  & n10295;
  assign n10318 = ~n10296 & n10317;
  assign n10319 = ~n10289 & n10318;
  assign n10320 = ~n10310 & ~n10319;
  assign n10321 = pi42  & ~n10320;
  assign n10322 = ~pi42  & n10320;
  assign n10323 = ~n10321 & ~n10322;
  assign n10324 = ~n10316 & ~n10323;
  assign n10325 = ~n10314 & ~n10324;
  assign n10326 = po23  & ~n10325;
  assign n10327 = ~n9847 & ~n9851;
  assign n10328 = ~n9855 & n10327;
  assign n10329 = po20  & n10328;
  assign n10330 = po20  & n10327;
  assign n10331 = n9855 & ~n10330;
  assign n10332 = ~n10329 & ~n10331;
  assign n10333 = ~po23  & n10325;
  assign n10334 = ~n10332 & ~n10333;
  assign n10335 = ~n10326 & ~n10334;
  assign n10336 = po24  & ~n10335;
  assign n10337 = ~n9858 & ~n9866;
  assign n10338 = n9865 & n10337;
  assign n10339 = po20  & n10338;
  assign n10340 = po20  & n10337;
  assign n10341 = ~n9865 & ~n10340;
  assign n10342 = ~n10339 & ~n10341;
  assign n10343 = ~po24  & ~n10326;
  assign n10344 = ~n10334 & n10343;
  assign n10345 = ~n10342 & ~n10344;
  assign n10346 = ~n10336 & ~n10345;
  assign n10347 = po25  & ~n10346;
  assign n10348 = ~n9869 & ~n9877;
  assign n10349 = n9875 & n10348;
  assign n10350 = po20  & n10349;
  assign n10351 = po20  & n10348;
  assign n10352 = ~n9875 & ~n10351;
  assign n10353 = ~n10350 & ~n10352;
  assign n10354 = ~po25  & n10346;
  assign n10355 = ~n10353 & ~n10354;
  assign n10356 = ~n10347 & ~n10355;
  assign n10357 = po26  & ~n10356;
  assign n10358 = ~n9880 & ~n9887;
  assign n10359 = n9886 & n10358;
  assign n10360 = po20  & n10359;
  assign n10361 = po20  & n10358;
  assign n10362 = ~n9886 & ~n10361;
  assign n10363 = ~n10360 & ~n10362;
  assign n10364 = ~po26  & ~n10347;
  assign n10365 = ~n10355 & n10364;
  assign n10366 = ~n10363 & ~n10365;
  assign n10367 = ~n10357 & ~n10366;
  assign n10368 = po27  & ~n10367;
  assign n10369 = ~n9890 & ~n9898;
  assign n10370 = n9896 & n10369;
  assign n10371 = po20  & n10370;
  assign n10372 = po20  & n10369;
  assign n10373 = ~n9896 & ~n10372;
  assign n10374 = ~n10371 & ~n10373;
  assign n10375 = ~po27  & n10367;
  assign n10376 = ~n10374 & ~n10375;
  assign n10377 = ~n10368 & ~n10376;
  assign n10378 = po28  & ~n10377;
  assign n10379 = ~n9901 & ~n9908;
  assign n10380 = n9907 & n10379;
  assign n10381 = po20  & n10380;
  assign n10382 = po20  & n10379;
  assign n10383 = ~n9907 & ~n10382;
  assign n10384 = ~n10381 & ~n10383;
  assign n10385 = ~po28  & ~n10368;
  assign n10386 = ~n10376 & n10385;
  assign n10387 = ~n10384 & ~n10386;
  assign n10388 = ~n10378 & ~n10387;
  assign n10389 = po29  & ~n10388;
  assign n10390 = ~n9911 & ~n9919;
  assign n10391 = n9917 & n10390;
  assign n10392 = po20  & n10391;
  assign n10393 = po20  & n10390;
  assign n10394 = ~n9917 & ~n10393;
  assign n10395 = ~n10392 & ~n10394;
  assign n10396 = ~po29  & n10388;
  assign n10397 = ~n10395 & ~n10396;
  assign n10398 = ~n10389 & ~n10397;
  assign n10399 = po30  & ~n10398;
  assign n10400 = ~n9922 & ~n9929;
  assign n10401 = n9928 & n10400;
  assign n10402 = po20  & n10401;
  assign n10403 = po20  & n10400;
  assign n10404 = ~n9928 & ~n10403;
  assign n10405 = ~n10402 & ~n10404;
  assign n10406 = ~po30  & ~n10389;
  assign n10407 = ~n10397 & n10406;
  assign n10408 = ~n10405 & ~n10407;
  assign n10409 = ~n10399 & ~n10408;
  assign n10410 = po31  & ~n10409;
  assign n10411 = ~n9932 & ~n9940;
  assign n10412 = n9938 & n10411;
  assign n10413 = po20  & n10412;
  assign n10414 = po20  & n10411;
  assign n10415 = ~n9938 & ~n10414;
  assign n10416 = ~n10413 & ~n10415;
  assign n10417 = ~po31  & n10409;
  assign n10418 = ~n10416 & ~n10417;
  assign n10419 = ~n10410 & ~n10418;
  assign n10420 = po32  & ~n10419;
  assign n10421 = ~n9943 & ~n9950;
  assign n10422 = n9949 & n10421;
  assign n10423 = po20  & n10422;
  assign n10424 = po20  & n10421;
  assign n10425 = ~n9949 & ~n10424;
  assign n10426 = ~n10423 & ~n10425;
  assign n10427 = ~po32  & ~n10410;
  assign n10428 = ~n10418 & n10427;
  assign n10429 = ~n10426 & ~n10428;
  assign n10430 = ~n10420 & ~n10429;
  assign n10431 = po33  & ~n10430;
  assign n10432 = ~n9953 & ~n9961;
  assign n10433 = n9959 & n10432;
  assign n10434 = po20  & n10433;
  assign n10435 = po20  & n10432;
  assign n10436 = ~n9959 & ~n10435;
  assign n10437 = ~n10434 & ~n10436;
  assign n10438 = ~po33  & n10430;
  assign n10439 = ~n10437 & ~n10438;
  assign n10440 = ~n10431 & ~n10439;
  assign n10441 = po34  & ~n10440;
  assign n10442 = ~n9964 & ~n9971;
  assign n10443 = n9970 & n10442;
  assign n10444 = po20  & n10443;
  assign n10445 = po20  & n10442;
  assign n10446 = ~n9970 & ~n10445;
  assign n10447 = ~n10444 & ~n10446;
  assign n10448 = ~po34  & ~n10431;
  assign n10449 = ~n10439 & n10448;
  assign n10450 = ~n10447 & ~n10449;
  assign n10451 = ~n10441 & ~n10450;
  assign n10452 = po35  & ~n10451;
  assign n10453 = ~n9974 & ~n9982;
  assign n10454 = n9980 & n10453;
  assign n10455 = po20  & n10454;
  assign n10456 = po20  & n10453;
  assign n10457 = ~n9980 & ~n10456;
  assign n10458 = ~n10455 & ~n10457;
  assign n10459 = ~po35  & n10451;
  assign n10460 = ~n10458 & ~n10459;
  assign n10461 = ~n10452 & ~n10460;
  assign n10462 = po36  & ~n10461;
  assign n10463 = ~n9985 & ~n9992;
  assign n10464 = n9991 & n10463;
  assign n10465 = po20  & n10464;
  assign n10466 = po20  & n10463;
  assign n10467 = ~n9991 & ~n10466;
  assign n10468 = ~n10465 & ~n10467;
  assign n10469 = ~po36  & ~n10452;
  assign n10470 = ~n10460 & n10469;
  assign n10471 = ~n10468 & ~n10470;
  assign n10472 = ~n10462 & ~n10471;
  assign n10473 = po37  & ~n10472;
  assign n10474 = ~n9995 & ~n10003;
  assign n10475 = n10001 & n10474;
  assign n10476 = po20  & n10475;
  assign n10477 = po20  & n10474;
  assign n10478 = ~n10001 & ~n10477;
  assign n10479 = ~n10476 & ~n10478;
  assign n10480 = ~po37  & n10472;
  assign n10481 = ~n10479 & ~n10480;
  assign n10482 = ~n10473 & ~n10481;
  assign n10483 = po38  & ~n10482;
  assign n10484 = ~n10006 & ~n10013;
  assign n10485 = n10012 & n10484;
  assign n10486 = po20  & n10485;
  assign n10487 = po20  & n10484;
  assign n10488 = ~n10012 & ~n10487;
  assign n10489 = ~n10486 & ~n10488;
  assign n10490 = ~po38  & ~n10473;
  assign n10491 = ~n10481 & n10490;
  assign n10492 = ~n10489 & ~n10491;
  assign n10493 = ~n10483 & ~n10492;
  assign n10494 = po39  & ~n10493;
  assign n10495 = ~n10016 & ~n10024;
  assign n10496 = n10022 & n10495;
  assign n10497 = po20  & n10496;
  assign n10498 = po20  & n10495;
  assign n10499 = ~n10022 & ~n10498;
  assign n10500 = ~n10497 & ~n10499;
  assign n10501 = ~po39  & n10493;
  assign n10502 = ~n10500 & ~n10501;
  assign n10503 = ~n10494 & ~n10502;
  assign n10504 = po40  & ~n10503;
  assign n10505 = ~n10027 & ~n10034;
  assign n10506 = n10033 & n10505;
  assign n10507 = po20  & n10506;
  assign n10508 = po20  & n10505;
  assign n10509 = ~n10033 & ~n10508;
  assign n10510 = ~n10507 & ~n10509;
  assign n10511 = ~po40  & ~n10494;
  assign n10512 = ~n10502 & n10511;
  assign n10513 = ~n10510 & ~n10512;
  assign n10514 = ~n10504 & ~n10513;
  assign n10515 = po41  & ~n10514;
  assign n10516 = ~n10037 & ~n10045;
  assign n10517 = n10043 & n10516;
  assign n10518 = po20  & n10517;
  assign n10519 = po20  & n10516;
  assign n10520 = ~n10043 & ~n10519;
  assign n10521 = ~n10518 & ~n10520;
  assign n10522 = ~po41  & n10514;
  assign n10523 = ~n10521 & ~n10522;
  assign n10524 = ~n10515 & ~n10523;
  assign n10525 = po42  & ~n10524;
  assign n10526 = ~n10048 & ~n10055;
  assign n10527 = n10054 & n10526;
  assign n10528 = po20  & n10527;
  assign n10529 = po20  & n10526;
  assign n10530 = ~n10054 & ~n10529;
  assign n10531 = ~n10528 & ~n10530;
  assign n10532 = ~po42  & ~n10515;
  assign n10533 = ~n10523 & n10532;
  assign n10534 = ~n10531 & ~n10533;
  assign n10535 = ~n10525 & ~n10534;
  assign n10536 = po43  & ~n10535;
  assign n10537 = ~n10058 & ~n10066;
  assign n10538 = n10064 & n10537;
  assign n10539 = po20  & n10538;
  assign n10540 = po20  & n10537;
  assign n10541 = ~n10064 & ~n10540;
  assign n10542 = ~n10539 & ~n10541;
  assign n10543 = ~po43  & n10535;
  assign n10544 = ~n10542 & ~n10543;
  assign n10545 = ~n10536 & ~n10544;
  assign n10546 = po44  & ~n10545;
  assign n10547 = ~n10069 & ~n10076;
  assign n10548 = n10075 & n10547;
  assign n10549 = po20  & n10548;
  assign n10550 = po20  & n10547;
  assign n10551 = ~n10075 & ~n10550;
  assign n10552 = ~n10549 & ~n10551;
  assign n10553 = ~po44  & ~n10536;
  assign n10554 = ~n10544 & n10553;
  assign n10555 = ~n10552 & ~n10554;
  assign n10556 = ~n10546 & ~n10555;
  assign n10557 = po45  & ~n10556;
  assign n10558 = ~n10079 & ~n10081;
  assign n10559 = n10087 & n10558;
  assign n10560 = po20  & n10559;
  assign n10561 = po20  & n10558;
  assign n10562 = ~n10087 & ~n10561;
  assign n10563 = ~n10560 & ~n10562;
  assign n10564 = ~po45  & n10556;
  assign n10565 = ~n10563 & ~n10564;
  assign n10566 = ~n10557 & ~n10565;
  assign n10567 = po46  & ~n10566;
  assign n10568 = ~n10090 & ~n10097;
  assign n10569 = n10096 & n10568;
  assign n10570 = po20  & n10569;
  assign n10571 = po20  & n10568;
  assign n10572 = ~n10096 & ~n10571;
  assign n10573 = ~n10570 & ~n10572;
  assign n10574 = ~po46  & ~n10557;
  assign n10575 = ~n10565 & n10574;
  assign n10576 = ~n10573 & ~n10575;
  assign n10577 = ~n10567 & ~n10576;
  assign n10578 = po47  & ~n10577;
  assign n10579 = ~n10100 & ~n10108;
  assign n10580 = n10106 & n10579;
  assign n10581 = po20  & n10580;
  assign n10582 = po20  & n10579;
  assign n10583 = ~n10106 & ~n10582;
  assign n10584 = ~n10581 & ~n10583;
  assign n10585 = ~po47  & n10577;
  assign n10586 = ~n10584 & ~n10585;
  assign n10587 = ~n10578 & ~n10586;
  assign n10588 = po48  & ~n10587;
  assign n10589 = ~n10111 & ~n10118;
  assign n10590 = n10117 & n10589;
  assign n10591 = po20  & n10590;
  assign n10592 = po20  & n10589;
  assign n10593 = ~n10117 & ~n10592;
  assign n10594 = ~n10591 & ~n10593;
  assign n10595 = ~po48  & ~n10578;
  assign n10596 = ~n10586 & n10595;
  assign n10597 = ~n10594 & ~n10596;
  assign n10598 = ~n10588 & ~n10597;
  assign n10599 = po49  & ~n10598;
  assign n10600 = ~n10121 & ~n10129;
  assign n10601 = n10127 & n10600;
  assign n10602 = po20  & n10601;
  assign n10603 = po20  & n10600;
  assign n10604 = ~n10127 & ~n10603;
  assign n10605 = ~n10602 & ~n10604;
  assign n10606 = ~po49  & n10598;
  assign n10607 = ~n10605 & ~n10606;
  assign n10608 = ~n10599 & ~n10607;
  assign n10609 = po50  & ~n10608;
  assign n10610 = ~n10132 & ~n10139;
  assign n10611 = n10138 & n10610;
  assign n10612 = po20  & n10611;
  assign n10613 = po20  & n10610;
  assign n10614 = ~n10138 & ~n10613;
  assign n10615 = ~n10612 & ~n10614;
  assign n10616 = ~po50  & ~n10599;
  assign n10617 = ~n10607 & n10616;
  assign n10618 = ~n10615 & ~n10617;
  assign n10619 = ~n10609 & ~n10618;
  assign n10620 = po51  & ~n10619;
  assign n10621 = ~n10142 & ~n10150;
  assign n10622 = n10148 & n10621;
  assign n10623 = po20  & n10622;
  assign n10624 = po20  & n10621;
  assign n10625 = ~n10148 & ~n10624;
  assign n10626 = ~n10623 & ~n10625;
  assign n10627 = ~po51  & n10619;
  assign n10628 = ~n10626 & ~n10627;
  assign n10629 = ~n10620 & ~n10628;
  assign n10630 = po52  & ~n10629;
  assign n10631 = ~n10153 & ~n10160;
  assign n10632 = n10159 & n10631;
  assign n10633 = po20  & n10632;
  assign n10634 = po20  & n10631;
  assign n10635 = ~n10159 & ~n10634;
  assign n10636 = ~n10633 & ~n10635;
  assign n10637 = ~po52  & ~n10620;
  assign n10638 = ~n10628 & n10637;
  assign n10639 = ~n10636 & ~n10638;
  assign n10640 = ~n10630 & ~n10639;
  assign n10641 = po53  & ~n10640;
  assign n10642 = ~n10163 & ~n10171;
  assign n10643 = n10169 & n10642;
  assign n10644 = po20  & n10643;
  assign n10645 = po20  & n10642;
  assign n10646 = ~n10169 & ~n10645;
  assign n10647 = ~n10644 & ~n10646;
  assign n10648 = ~po53  & n10640;
  assign n10649 = ~n10647 & ~n10648;
  assign n10650 = ~n10641 & ~n10649;
  assign n10651 = po54  & ~n10650;
  assign n10652 = ~n10174 & ~n10181;
  assign n10653 = n10180 & n10652;
  assign n10654 = po20  & n10653;
  assign n10655 = po20  & n10652;
  assign n10656 = ~n10180 & ~n10655;
  assign n10657 = ~n10654 & ~n10656;
  assign n10658 = ~po54  & ~n10641;
  assign n10659 = ~n10649 & n10658;
  assign n10660 = ~n10657 & ~n10659;
  assign n10661 = ~n10651 & ~n10660;
  assign n10662 = po55  & ~n10661;
  assign n10663 = ~n10184 & ~n10192;
  assign n10664 = n10190 & n10663;
  assign n10665 = po20  & n10664;
  assign n10666 = po20  & n10663;
  assign n10667 = ~n10190 & ~n10666;
  assign n10668 = ~n10665 & ~n10667;
  assign n10669 = ~po55  & n10661;
  assign n10670 = ~n10668 & ~n10669;
  assign n10671 = ~n10662 & ~n10670;
  assign n10672 = po56  & ~n10671;
  assign n10673 = ~n10195 & ~n10202;
  assign n10674 = n10201 & n10673;
  assign n10675 = po20  & n10674;
  assign n10676 = po20  & n10673;
  assign n10677 = ~n10201 & ~n10676;
  assign n10678 = ~n10675 & ~n10677;
  assign n10679 = ~po56  & ~n10662;
  assign n10680 = ~n10670 & n10679;
  assign n10681 = ~n10678 & ~n10680;
  assign n10682 = ~n10672 & ~n10681;
  assign n10683 = po57  & ~n10682;
  assign n10684 = ~n10205 & ~n10213;
  assign n10685 = n10211 & n10684;
  assign n10686 = po20  & n10685;
  assign n10687 = po20  & n10684;
  assign n10688 = ~n10211 & ~n10687;
  assign n10689 = ~n10686 & ~n10688;
  assign n10690 = ~po57  & n10682;
  assign n10691 = ~n10689 & ~n10690;
  assign n10692 = ~n10683 & ~n10691;
  assign n10693 = po58  & ~n10692;
  assign n10694 = ~n10216 & ~n10223;
  assign n10695 = n10222 & n10694;
  assign n10696 = po20  & n10695;
  assign n10697 = po20  & n10694;
  assign n10698 = ~n10222 & ~n10697;
  assign n10699 = ~n10696 & ~n10698;
  assign n10700 = ~po58  & ~n10683;
  assign n10701 = ~n10691 & n10700;
  assign n10702 = ~n10699 & ~n10701;
  assign n10703 = ~n10693 & ~n10702;
  assign n10704 = po59  & ~n10703;
  assign n10705 = ~n10226 & ~n10234;
  assign n10706 = n10232 & n10705;
  assign n10707 = po20  & n10706;
  assign n10708 = po20  & n10705;
  assign n10709 = ~n10232 & ~n10708;
  assign n10710 = ~n10707 & ~n10709;
  assign n10711 = ~po59  & n10703;
  assign n10712 = ~n10710 & ~n10711;
  assign n10713 = ~n10704 & ~n10712;
  assign n10714 = po60  & ~n10713;
  assign n10715 = ~n10237 & ~n10244;
  assign n10716 = n10243 & n10715;
  assign n10717 = po20  & n10716;
  assign n10718 = po20  & n10715;
  assign n10719 = ~n10243 & ~n10718;
  assign n10720 = ~n10717 & ~n10719;
  assign n10721 = ~po60  & ~n10704;
  assign n10722 = ~n10712 & n10721;
  assign n10723 = ~n10720 & ~n10722;
  assign n10724 = ~n10714 & ~n10723;
  assign n10725 = po61  & ~n10724;
  assign n10726 = ~n10247 & ~n10255;
  assign n10727 = n10253 & n10726;
  assign n10728 = po20  & n10727;
  assign n10729 = po20  & n10726;
  assign n10730 = ~n10253 & ~n10729;
  assign n10731 = ~n10728 & ~n10730;
  assign n10732 = ~po61  & n10724;
  assign n10733 = ~n10731 & ~n10732;
  assign n10734 = ~n10725 & ~n10733;
  assign n10735 = po62  & ~n10734;
  assign n10736 = ~n10258 & ~n10265;
  assign n10737 = n10264 & n10736;
  assign n10738 = po20  & n10737;
  assign n10739 = po20  & n10736;
  assign n10740 = ~n10264 & ~n10739;
  assign n10741 = ~n10738 & ~n10740;
  assign n10742 = ~po62  & ~n10725;
  assign n10743 = ~n10733 & n10742;
  assign n10744 = ~n10741 & ~n10743;
  assign n10745 = ~n10735 & ~n10744;
  assign n10746 = ~n10268 & ~n10276;
  assign n10747 = po20  & n10746;
  assign n10748 = ~n10274 & ~n10747;
  assign n10749 = n10274 & n10747;
  assign n10750 = ~n10748 & ~n10749;
  assign n10751 = ~n10278 & ~n10283;
  assign n10752 = po20  & n10751;
  assign n10753 = ~n10296 & ~n10752;
  assign n10754 = ~n10750 & n10753;
  assign n10755 = ~n10745 & n10754;
  assign n10756 = ~po63  & ~n10755;
  assign n10757 = ~n10283 & po20 ;
  assign n10758 = n10278 & ~n10757;
  assign n10759 = po63  & ~n10751;
  assign n10760 = ~n10758 & n10759;
  assign n10761 = n10283 & ~po20 ;
  assign n10762 = ~n10760 & ~n10761;
  assign n10763 = n10745 & n10750;
  assign n10764 = n10762 & ~n10763;
  assign po19  = n10756 | ~n10764;
  assign n10766 = pi38  & po19 ;
  assign n10767 = ~pi36  & ~pi37 ;
  assign n10768 = ~pi38  & n10767;
  assign n10769 = ~n10766 & ~n10768;
  assign n10770 = po20  & ~n10769;
  assign n10771 = n10295 & ~n10768;
  assign n10772 = ~n10296 & n10771;
  assign n10773 = ~n10289 & n10772;
  assign n10774 = ~n10766 & n10773;
  assign n10775 = ~pi38  & po19 ;
  assign n10776 = pi39  & ~n10775;
  assign n10777 = n10300 & po19 ;
  assign n10778 = ~n10776 & ~n10777;
  assign n10779 = ~n10774 & n10778;
  assign n10780 = ~n10770 & ~n10779;
  assign n10781 = po21  & ~n10780;
  assign n10782 = po20  & n10762;
  assign n10783 = ~n10763 & n10782;
  assign n10784 = ~n10756 & n10783;
  assign n10785 = ~n10777 & ~n10784;
  assign n10786 = pi40  & ~n10785;
  assign n10787 = ~pi40  & n10785;
  assign n10788 = ~n10786 & ~n10787;
  assign n10789 = ~po21  & n10780;
  assign n10790 = ~n10788 & ~n10789;
  assign n10791 = ~n10781 & ~n10790;
  assign n10792 = po22  & ~n10791;
  assign n10793 = ~n10303 & ~n10307;
  assign n10794 = ~n10311 & n10793;
  assign n10795 = po19  & n10794;
  assign n10796 = po19  & n10793;
  assign n10797 = n10311 & ~n10796;
  assign n10798 = ~n10795 & ~n10797;
  assign n10799 = ~po22  & ~n10781;
  assign n10800 = ~n10790 & n10799;
  assign n10801 = ~n10798 & ~n10800;
  assign n10802 = ~n10792 & ~n10801;
  assign n10803 = po23  & ~n10802;
  assign n10804 = ~n10314 & ~n10316;
  assign n10805 = n10323 & n10804;
  assign n10806 = po19  & n10805;
  assign n10807 = po19  & n10804;
  assign n10808 = ~n10323 & ~n10807;
  assign n10809 = ~n10806 & ~n10808;
  assign n10810 = ~po23  & n10802;
  assign n10811 = ~n10809 & ~n10810;
  assign n10812 = ~n10803 & ~n10811;
  assign n10813 = po24  & ~n10812;
  assign n10814 = ~n10326 & ~n10333;
  assign n10815 = n10332 & n10814;
  assign n10816 = po19  & n10815;
  assign n10817 = po19  & n10814;
  assign n10818 = ~n10332 & ~n10817;
  assign n10819 = ~n10816 & ~n10818;
  assign n10820 = ~po24  & ~n10803;
  assign n10821 = ~n10811 & n10820;
  assign n10822 = ~n10819 & ~n10821;
  assign n10823 = ~n10813 & ~n10822;
  assign n10824 = po25  & ~n10823;
  assign n10825 = ~n10336 & ~n10344;
  assign n10826 = n10342 & n10825;
  assign n10827 = po19  & n10826;
  assign n10828 = po19  & n10825;
  assign n10829 = ~n10342 & ~n10828;
  assign n10830 = ~n10827 & ~n10829;
  assign n10831 = ~po25  & n10823;
  assign n10832 = ~n10830 & ~n10831;
  assign n10833 = ~n10824 & ~n10832;
  assign n10834 = po26  & ~n10833;
  assign n10835 = ~n10347 & ~n10354;
  assign n10836 = n10353 & n10835;
  assign n10837 = po19  & n10836;
  assign n10838 = po19  & n10835;
  assign n10839 = ~n10353 & ~n10838;
  assign n10840 = ~n10837 & ~n10839;
  assign n10841 = ~po26  & ~n10824;
  assign n10842 = ~n10832 & n10841;
  assign n10843 = ~n10840 & ~n10842;
  assign n10844 = ~n10834 & ~n10843;
  assign n10845 = po27  & ~n10844;
  assign n10846 = ~n10357 & ~n10365;
  assign n10847 = n10363 & n10846;
  assign n10848 = po19  & n10847;
  assign n10849 = po19  & n10846;
  assign n10850 = ~n10363 & ~n10849;
  assign n10851 = ~n10848 & ~n10850;
  assign n10852 = ~po27  & n10844;
  assign n10853 = ~n10851 & ~n10852;
  assign n10854 = ~n10845 & ~n10853;
  assign n10855 = po28  & ~n10854;
  assign n10856 = ~n10368 & ~n10375;
  assign n10857 = n10374 & n10856;
  assign n10858 = po19  & n10857;
  assign n10859 = po19  & n10856;
  assign n10860 = ~n10374 & ~n10859;
  assign n10861 = ~n10858 & ~n10860;
  assign n10862 = ~po28  & ~n10845;
  assign n10863 = ~n10853 & n10862;
  assign n10864 = ~n10861 & ~n10863;
  assign n10865 = ~n10855 & ~n10864;
  assign n10866 = po29  & ~n10865;
  assign n10867 = ~n10378 & ~n10386;
  assign n10868 = n10384 & n10867;
  assign n10869 = po19  & n10868;
  assign n10870 = po19  & n10867;
  assign n10871 = ~n10384 & ~n10870;
  assign n10872 = ~n10869 & ~n10871;
  assign n10873 = ~po29  & n10865;
  assign n10874 = ~n10872 & ~n10873;
  assign n10875 = ~n10866 & ~n10874;
  assign n10876 = po30  & ~n10875;
  assign n10877 = ~n10389 & ~n10396;
  assign n10878 = n10395 & n10877;
  assign n10879 = po19  & n10878;
  assign n10880 = po19  & n10877;
  assign n10881 = ~n10395 & ~n10880;
  assign n10882 = ~n10879 & ~n10881;
  assign n10883 = ~po30  & ~n10866;
  assign n10884 = ~n10874 & n10883;
  assign n10885 = ~n10882 & ~n10884;
  assign n10886 = ~n10876 & ~n10885;
  assign n10887 = po31  & ~n10886;
  assign n10888 = ~n10399 & ~n10407;
  assign n10889 = n10405 & n10888;
  assign n10890 = po19  & n10889;
  assign n10891 = po19  & n10888;
  assign n10892 = ~n10405 & ~n10891;
  assign n10893 = ~n10890 & ~n10892;
  assign n10894 = ~po31  & n10886;
  assign n10895 = ~n10893 & ~n10894;
  assign n10896 = ~n10887 & ~n10895;
  assign n10897 = po32  & ~n10896;
  assign n10898 = ~n10410 & ~n10417;
  assign n10899 = n10416 & n10898;
  assign n10900 = po19  & n10899;
  assign n10901 = po19  & n10898;
  assign n10902 = ~n10416 & ~n10901;
  assign n10903 = ~n10900 & ~n10902;
  assign n10904 = ~po32  & ~n10887;
  assign n10905 = ~n10895 & n10904;
  assign n10906 = ~n10903 & ~n10905;
  assign n10907 = ~n10897 & ~n10906;
  assign n10908 = po33  & ~n10907;
  assign n10909 = ~n10420 & ~n10428;
  assign n10910 = n10426 & n10909;
  assign n10911 = po19  & n10910;
  assign n10912 = po19  & n10909;
  assign n10913 = ~n10426 & ~n10912;
  assign n10914 = ~n10911 & ~n10913;
  assign n10915 = ~po33  & n10907;
  assign n10916 = ~n10914 & ~n10915;
  assign n10917 = ~n10908 & ~n10916;
  assign n10918 = po34  & ~n10917;
  assign n10919 = ~n10431 & ~n10438;
  assign n10920 = n10437 & n10919;
  assign n10921 = po19  & n10920;
  assign n10922 = po19  & n10919;
  assign n10923 = ~n10437 & ~n10922;
  assign n10924 = ~n10921 & ~n10923;
  assign n10925 = ~po34  & ~n10908;
  assign n10926 = ~n10916 & n10925;
  assign n10927 = ~n10924 & ~n10926;
  assign n10928 = ~n10918 & ~n10927;
  assign n10929 = po35  & ~n10928;
  assign n10930 = ~n10441 & ~n10449;
  assign n10931 = n10447 & n10930;
  assign n10932 = po19  & n10931;
  assign n10933 = po19  & n10930;
  assign n10934 = ~n10447 & ~n10933;
  assign n10935 = ~n10932 & ~n10934;
  assign n10936 = ~po35  & n10928;
  assign n10937 = ~n10935 & ~n10936;
  assign n10938 = ~n10929 & ~n10937;
  assign n10939 = po36  & ~n10938;
  assign n10940 = ~n10452 & ~n10459;
  assign n10941 = n10458 & n10940;
  assign n10942 = po19  & n10941;
  assign n10943 = po19  & n10940;
  assign n10944 = ~n10458 & ~n10943;
  assign n10945 = ~n10942 & ~n10944;
  assign n10946 = ~po36  & ~n10929;
  assign n10947 = ~n10937 & n10946;
  assign n10948 = ~n10945 & ~n10947;
  assign n10949 = ~n10939 & ~n10948;
  assign n10950 = po37  & ~n10949;
  assign n10951 = ~n10462 & ~n10470;
  assign n10952 = n10468 & n10951;
  assign n10953 = po19  & n10952;
  assign n10954 = po19  & n10951;
  assign n10955 = ~n10468 & ~n10954;
  assign n10956 = ~n10953 & ~n10955;
  assign n10957 = ~po37  & n10949;
  assign n10958 = ~n10956 & ~n10957;
  assign n10959 = ~n10950 & ~n10958;
  assign n10960 = po38  & ~n10959;
  assign n10961 = ~n10473 & ~n10480;
  assign n10962 = n10479 & n10961;
  assign n10963 = po19  & n10962;
  assign n10964 = po19  & n10961;
  assign n10965 = ~n10479 & ~n10964;
  assign n10966 = ~n10963 & ~n10965;
  assign n10967 = ~po38  & ~n10950;
  assign n10968 = ~n10958 & n10967;
  assign n10969 = ~n10966 & ~n10968;
  assign n10970 = ~n10960 & ~n10969;
  assign n10971 = po39  & ~n10970;
  assign n10972 = ~n10483 & ~n10491;
  assign n10973 = n10489 & n10972;
  assign n10974 = po19  & n10973;
  assign n10975 = po19  & n10972;
  assign n10976 = ~n10489 & ~n10975;
  assign n10977 = ~n10974 & ~n10976;
  assign n10978 = ~po39  & n10970;
  assign n10979 = ~n10977 & ~n10978;
  assign n10980 = ~n10971 & ~n10979;
  assign n10981 = po40  & ~n10980;
  assign n10982 = ~n10494 & ~n10501;
  assign n10983 = n10500 & n10982;
  assign n10984 = po19  & n10983;
  assign n10985 = po19  & n10982;
  assign n10986 = ~n10500 & ~n10985;
  assign n10987 = ~n10984 & ~n10986;
  assign n10988 = ~po40  & ~n10971;
  assign n10989 = ~n10979 & n10988;
  assign n10990 = ~n10987 & ~n10989;
  assign n10991 = ~n10981 & ~n10990;
  assign n10992 = po41  & ~n10991;
  assign n10993 = ~n10504 & ~n10512;
  assign n10994 = n10510 & n10993;
  assign n10995 = po19  & n10994;
  assign n10996 = po19  & n10993;
  assign n10997 = ~n10510 & ~n10996;
  assign n10998 = ~n10995 & ~n10997;
  assign n10999 = ~po41  & n10991;
  assign n11000 = ~n10998 & ~n10999;
  assign n11001 = ~n10992 & ~n11000;
  assign n11002 = po42  & ~n11001;
  assign n11003 = ~n10515 & ~n10522;
  assign n11004 = n10521 & n11003;
  assign n11005 = po19  & n11004;
  assign n11006 = po19  & n11003;
  assign n11007 = ~n10521 & ~n11006;
  assign n11008 = ~n11005 & ~n11007;
  assign n11009 = ~po42  & ~n10992;
  assign n11010 = ~n11000 & n11009;
  assign n11011 = ~n11008 & ~n11010;
  assign n11012 = ~n11002 & ~n11011;
  assign n11013 = po43  & ~n11012;
  assign n11014 = ~n10525 & ~n10533;
  assign n11015 = n10531 & n11014;
  assign n11016 = po19  & n11015;
  assign n11017 = po19  & n11014;
  assign n11018 = ~n10531 & ~n11017;
  assign n11019 = ~n11016 & ~n11018;
  assign n11020 = ~po43  & n11012;
  assign n11021 = ~n11019 & ~n11020;
  assign n11022 = ~n11013 & ~n11021;
  assign n11023 = po44  & ~n11022;
  assign n11024 = ~n10536 & ~n10543;
  assign n11025 = n10542 & n11024;
  assign n11026 = po19  & n11025;
  assign n11027 = po19  & n11024;
  assign n11028 = ~n10542 & ~n11027;
  assign n11029 = ~n11026 & ~n11028;
  assign n11030 = ~po44  & ~n11013;
  assign n11031 = ~n11021 & n11030;
  assign n11032 = ~n11029 & ~n11031;
  assign n11033 = ~n11023 & ~n11032;
  assign n11034 = po45  & ~n11033;
  assign n11035 = ~n10546 & ~n10554;
  assign n11036 = n10552 & n11035;
  assign n11037 = po19  & n11036;
  assign n11038 = po19  & n11035;
  assign n11039 = ~n10552 & ~n11038;
  assign n11040 = ~n11037 & ~n11039;
  assign n11041 = ~po45  & n11033;
  assign n11042 = ~n11040 & ~n11041;
  assign n11043 = ~n11034 & ~n11042;
  assign n11044 = po46  & ~n11043;
  assign n11045 = ~po46  & ~n11034;
  assign n11046 = ~n11042 & n11045;
  assign n11047 = ~n10557 & ~n10564;
  assign n11048 = n10563 & n11047;
  assign n11049 = po19  & n11048;
  assign n11050 = po19  & n11047;
  assign n11051 = ~n10563 & ~n11050;
  assign n11052 = ~n11049 & ~n11051;
  assign n11053 = ~n11046 & ~n11052;
  assign n11054 = ~n11044 & ~n11053;
  assign n11055 = po47  & ~n11054;
  assign n11056 = ~n10567 & ~n10575;
  assign n11057 = n10573 & n11056;
  assign n11058 = po19  & n11057;
  assign n11059 = po19  & n11056;
  assign n11060 = ~n10573 & ~n11059;
  assign n11061 = ~n11058 & ~n11060;
  assign n11062 = ~po47  & n11054;
  assign n11063 = ~n11061 & ~n11062;
  assign n11064 = ~n11055 & ~n11063;
  assign n11065 = po48  & ~n11064;
  assign n11066 = ~n10578 & ~n10585;
  assign n11067 = n10584 & n11066;
  assign n11068 = po19  & n11067;
  assign n11069 = po19  & n11066;
  assign n11070 = ~n10584 & ~n11069;
  assign n11071 = ~n11068 & ~n11070;
  assign n11072 = ~po48  & ~n11055;
  assign n11073 = ~n11063 & n11072;
  assign n11074 = ~n11071 & ~n11073;
  assign n11075 = ~n11065 & ~n11074;
  assign n11076 = po49  & ~n11075;
  assign n11077 = ~n10588 & ~n10596;
  assign n11078 = n10594 & n11077;
  assign n11079 = po19  & n11078;
  assign n11080 = po19  & n11077;
  assign n11081 = ~n10594 & ~n11080;
  assign n11082 = ~n11079 & ~n11081;
  assign n11083 = ~po49  & n11075;
  assign n11084 = ~n11082 & ~n11083;
  assign n11085 = ~n11076 & ~n11084;
  assign n11086 = po50  & ~n11085;
  assign n11087 = ~n10599 & ~n10606;
  assign n11088 = n10605 & n11087;
  assign n11089 = po19  & n11088;
  assign n11090 = po19  & n11087;
  assign n11091 = ~n10605 & ~n11090;
  assign n11092 = ~n11089 & ~n11091;
  assign n11093 = ~po50  & ~n11076;
  assign n11094 = ~n11084 & n11093;
  assign n11095 = ~n11092 & ~n11094;
  assign n11096 = ~n11086 & ~n11095;
  assign n11097 = po51  & ~n11096;
  assign n11098 = ~n10609 & ~n10617;
  assign n11099 = n10615 & n11098;
  assign n11100 = po19  & n11099;
  assign n11101 = po19  & n11098;
  assign n11102 = ~n10615 & ~n11101;
  assign n11103 = ~n11100 & ~n11102;
  assign n11104 = ~po51  & n11096;
  assign n11105 = ~n11103 & ~n11104;
  assign n11106 = ~n11097 & ~n11105;
  assign n11107 = po52  & ~n11106;
  assign n11108 = ~n10620 & ~n10627;
  assign n11109 = n10626 & n11108;
  assign n11110 = po19  & n11109;
  assign n11111 = po19  & n11108;
  assign n11112 = ~n10626 & ~n11111;
  assign n11113 = ~n11110 & ~n11112;
  assign n11114 = ~po52  & ~n11097;
  assign n11115 = ~n11105 & n11114;
  assign n11116 = ~n11113 & ~n11115;
  assign n11117 = ~n11107 & ~n11116;
  assign n11118 = po53  & ~n11117;
  assign n11119 = ~n10630 & ~n10638;
  assign n11120 = n10636 & n11119;
  assign n11121 = po19  & n11120;
  assign n11122 = po19  & n11119;
  assign n11123 = ~n10636 & ~n11122;
  assign n11124 = ~n11121 & ~n11123;
  assign n11125 = ~po53  & n11117;
  assign n11126 = ~n11124 & ~n11125;
  assign n11127 = ~n11118 & ~n11126;
  assign n11128 = po54  & ~n11127;
  assign n11129 = ~n10641 & ~n10648;
  assign n11130 = n10647 & n11129;
  assign n11131 = po19  & n11130;
  assign n11132 = po19  & n11129;
  assign n11133 = ~n10647 & ~n11132;
  assign n11134 = ~n11131 & ~n11133;
  assign n11135 = ~po54  & ~n11118;
  assign n11136 = ~n11126 & n11135;
  assign n11137 = ~n11134 & ~n11136;
  assign n11138 = ~n11128 & ~n11137;
  assign n11139 = po55  & ~n11138;
  assign n11140 = ~n10651 & ~n10659;
  assign n11141 = n10657 & n11140;
  assign n11142 = po19  & n11141;
  assign n11143 = po19  & n11140;
  assign n11144 = ~n10657 & ~n11143;
  assign n11145 = ~n11142 & ~n11144;
  assign n11146 = ~po55  & n11138;
  assign n11147 = ~n11145 & ~n11146;
  assign n11148 = ~n11139 & ~n11147;
  assign n11149 = po56  & ~n11148;
  assign n11150 = ~n10662 & ~n10669;
  assign n11151 = n10668 & n11150;
  assign n11152 = po19  & n11151;
  assign n11153 = po19  & n11150;
  assign n11154 = ~n10668 & ~n11153;
  assign n11155 = ~n11152 & ~n11154;
  assign n11156 = ~po56  & ~n11139;
  assign n11157 = ~n11147 & n11156;
  assign n11158 = ~n11155 & ~n11157;
  assign n11159 = ~n11149 & ~n11158;
  assign n11160 = po57  & ~n11159;
  assign n11161 = ~n10672 & ~n10680;
  assign n11162 = n10678 & n11161;
  assign n11163 = po19  & n11162;
  assign n11164 = po19  & n11161;
  assign n11165 = ~n10678 & ~n11164;
  assign n11166 = ~n11163 & ~n11165;
  assign n11167 = ~po57  & n11159;
  assign n11168 = ~n11166 & ~n11167;
  assign n11169 = ~n11160 & ~n11168;
  assign n11170 = po58  & ~n11169;
  assign n11171 = ~n10683 & ~n10690;
  assign n11172 = n10689 & n11171;
  assign n11173 = po19  & n11172;
  assign n11174 = po19  & n11171;
  assign n11175 = ~n10689 & ~n11174;
  assign n11176 = ~n11173 & ~n11175;
  assign n11177 = ~po58  & ~n11160;
  assign n11178 = ~n11168 & n11177;
  assign n11179 = ~n11176 & ~n11178;
  assign n11180 = ~n11170 & ~n11179;
  assign n11181 = po59  & ~n11180;
  assign n11182 = ~n10693 & ~n10701;
  assign n11183 = n10699 & n11182;
  assign n11184 = po19  & n11183;
  assign n11185 = po19  & n11182;
  assign n11186 = ~n10699 & ~n11185;
  assign n11187 = ~n11184 & ~n11186;
  assign n11188 = ~po59  & n11180;
  assign n11189 = ~n11187 & ~n11188;
  assign n11190 = ~n11181 & ~n11189;
  assign n11191 = po60  & ~n11190;
  assign n11192 = ~n10704 & ~n10711;
  assign n11193 = n10710 & n11192;
  assign n11194 = po19  & n11193;
  assign n11195 = po19  & n11192;
  assign n11196 = ~n10710 & ~n11195;
  assign n11197 = ~n11194 & ~n11196;
  assign n11198 = ~po60  & ~n11181;
  assign n11199 = ~n11189 & n11198;
  assign n11200 = ~n11197 & ~n11199;
  assign n11201 = ~n11191 & ~n11200;
  assign n11202 = po61  & ~n11201;
  assign n11203 = ~n10714 & ~n10722;
  assign n11204 = n10720 & n11203;
  assign n11205 = po19  & n11204;
  assign n11206 = po19  & n11203;
  assign n11207 = ~n10720 & ~n11206;
  assign n11208 = ~n11205 & ~n11207;
  assign n11209 = ~po61  & n11201;
  assign n11210 = ~n11208 & ~n11209;
  assign n11211 = ~n11202 & ~n11210;
  assign n11212 = po62  & ~n11211;
  assign n11213 = ~n10725 & ~n10732;
  assign n11214 = n10731 & n11213;
  assign n11215 = po19  & n11214;
  assign n11216 = po19  & n11213;
  assign n11217 = ~n10731 & ~n11216;
  assign n11218 = ~n11215 & ~n11217;
  assign n11219 = ~po62  & ~n11202;
  assign n11220 = ~n11210 & n11219;
  assign n11221 = ~n11218 & ~n11220;
  assign n11222 = ~n11212 & ~n11221;
  assign n11223 = ~n10735 & ~n10743;
  assign n11224 = po19  & n11223;
  assign n11225 = ~n10741 & ~n11224;
  assign n11226 = n10741 & n11224;
  assign n11227 = ~n11225 & ~n11226;
  assign n11228 = ~n10745 & ~n10750;
  assign n11229 = po19  & n11228;
  assign n11230 = ~n10763 & ~n11229;
  assign n11231 = ~n11227 & n11230;
  assign n11232 = ~n11222 & n11231;
  assign n11233 = ~po63  & ~n11232;
  assign n11234 = ~n10750 & po19 ;
  assign n11235 = n10745 & ~n11234;
  assign n11236 = po63  & ~n11228;
  assign n11237 = ~n11235 & n11236;
  assign n11238 = n10750 & ~po19 ;
  assign n11239 = ~n11237 & ~n11238;
  assign n11240 = n11222 & n11227;
  assign n11241 = n11239 & ~n11240;
  assign po18  = n11233 | ~n11241;
  assign n11243 = pi36  & po18 ;
  assign n11244 = ~pi34  & ~pi35 ;
  assign n11245 = ~pi36  & n11244;
  assign n11246 = ~n11243 & ~n11245;
  assign n11247 = po19  & ~n11246;
  assign n11248 = n10762 & ~n11245;
  assign n11249 = ~n10763 & n11248;
  assign n11250 = ~n10756 & n11249;
  assign n11251 = ~n11243 & n11250;
  assign n11252 = ~pi36  & po18 ;
  assign n11253 = pi37  & ~n11252;
  assign n11254 = n10767 & po18 ;
  assign n11255 = ~n11253 & ~n11254;
  assign n11256 = ~n11251 & n11255;
  assign n11257 = ~n11247 & ~n11256;
  assign n11258 = po20  & ~n11257;
  assign n11259 = ~po20  & ~n11247;
  assign n11260 = ~n11256 & n11259;
  assign n11261 = po19  & n11239;
  assign n11262 = ~n11240 & n11261;
  assign n11263 = ~n11233 & n11262;
  assign n11264 = ~n11254 & ~n11263;
  assign n11265 = pi38  & ~n11264;
  assign n11266 = ~pi38  & n11264;
  assign n11267 = ~n11265 & ~n11266;
  assign n11268 = ~n11260 & ~n11267;
  assign n11269 = ~n11258 & ~n11268;
  assign n11270 = po21  & ~n11269;
  assign n11271 = ~n10770 & ~n10774;
  assign n11272 = ~n10778 & n11271;
  assign n11273 = po18  & n11272;
  assign n11274 = po18  & n11271;
  assign n11275 = n10778 & ~n11274;
  assign n11276 = ~n11273 & ~n11275;
  assign n11277 = ~po21  & n11269;
  assign n11278 = ~n11276 & ~n11277;
  assign n11279 = ~n11270 & ~n11278;
  assign n11280 = po22  & ~n11279;
  assign n11281 = ~n10781 & ~n10789;
  assign n11282 = n10788 & n11281;
  assign n11283 = po18  & n11282;
  assign n11284 = po18  & n11281;
  assign n11285 = ~n10788 & ~n11284;
  assign n11286 = ~n11283 & ~n11285;
  assign n11287 = ~po22  & ~n11270;
  assign n11288 = ~n11278 & n11287;
  assign n11289 = ~n11286 & ~n11288;
  assign n11290 = ~n11280 & ~n11289;
  assign n11291 = po23  & ~n11290;
  assign n11292 = ~n10792 & ~n10800;
  assign n11293 = n10798 & n11292;
  assign n11294 = po18  & n11293;
  assign n11295 = po18  & n11292;
  assign n11296 = ~n10798 & ~n11295;
  assign n11297 = ~n11294 & ~n11296;
  assign n11298 = ~po23  & n11290;
  assign n11299 = ~n11297 & ~n11298;
  assign n11300 = ~n11291 & ~n11299;
  assign n11301 = po24  & ~n11300;
  assign n11302 = ~n10803 & ~n10810;
  assign n11303 = n10809 & n11302;
  assign n11304 = po18  & n11303;
  assign n11305 = po18  & n11302;
  assign n11306 = ~n10809 & ~n11305;
  assign n11307 = ~n11304 & ~n11306;
  assign n11308 = ~po24  & ~n11291;
  assign n11309 = ~n11299 & n11308;
  assign n11310 = ~n11307 & ~n11309;
  assign n11311 = ~n11301 & ~n11310;
  assign n11312 = po25  & ~n11311;
  assign n11313 = ~n10813 & ~n10821;
  assign n11314 = n10819 & n11313;
  assign n11315 = po18  & n11314;
  assign n11316 = po18  & n11313;
  assign n11317 = ~n10819 & ~n11316;
  assign n11318 = ~n11315 & ~n11317;
  assign n11319 = ~po25  & n11311;
  assign n11320 = ~n11318 & ~n11319;
  assign n11321 = ~n11312 & ~n11320;
  assign n11322 = po26  & ~n11321;
  assign n11323 = ~n10824 & ~n10831;
  assign n11324 = n10830 & n11323;
  assign n11325 = po18  & n11324;
  assign n11326 = po18  & n11323;
  assign n11327 = ~n10830 & ~n11326;
  assign n11328 = ~n11325 & ~n11327;
  assign n11329 = ~po26  & ~n11312;
  assign n11330 = ~n11320 & n11329;
  assign n11331 = ~n11328 & ~n11330;
  assign n11332 = ~n11322 & ~n11331;
  assign n11333 = po27  & ~n11332;
  assign n11334 = ~n10834 & ~n10842;
  assign n11335 = n10840 & n11334;
  assign n11336 = po18  & n11335;
  assign n11337 = po18  & n11334;
  assign n11338 = ~n10840 & ~n11337;
  assign n11339 = ~n11336 & ~n11338;
  assign n11340 = ~po27  & n11332;
  assign n11341 = ~n11339 & ~n11340;
  assign n11342 = ~n11333 & ~n11341;
  assign n11343 = po28  & ~n11342;
  assign n11344 = ~n10845 & ~n10852;
  assign n11345 = n10851 & n11344;
  assign n11346 = po18  & n11345;
  assign n11347 = po18  & n11344;
  assign n11348 = ~n10851 & ~n11347;
  assign n11349 = ~n11346 & ~n11348;
  assign n11350 = ~po28  & ~n11333;
  assign n11351 = ~n11341 & n11350;
  assign n11352 = ~n11349 & ~n11351;
  assign n11353 = ~n11343 & ~n11352;
  assign n11354 = po29  & ~n11353;
  assign n11355 = ~n10855 & ~n10863;
  assign n11356 = n10861 & n11355;
  assign n11357 = po18  & n11356;
  assign n11358 = po18  & n11355;
  assign n11359 = ~n10861 & ~n11358;
  assign n11360 = ~n11357 & ~n11359;
  assign n11361 = ~po29  & n11353;
  assign n11362 = ~n11360 & ~n11361;
  assign n11363 = ~n11354 & ~n11362;
  assign n11364 = po30  & ~n11363;
  assign n11365 = ~n10866 & ~n10873;
  assign n11366 = n10872 & n11365;
  assign n11367 = po18  & n11366;
  assign n11368 = po18  & n11365;
  assign n11369 = ~n10872 & ~n11368;
  assign n11370 = ~n11367 & ~n11369;
  assign n11371 = ~po30  & ~n11354;
  assign n11372 = ~n11362 & n11371;
  assign n11373 = ~n11370 & ~n11372;
  assign n11374 = ~n11364 & ~n11373;
  assign n11375 = po31  & ~n11374;
  assign n11376 = ~n10876 & ~n10884;
  assign n11377 = n10882 & n11376;
  assign n11378 = po18  & n11377;
  assign n11379 = po18  & n11376;
  assign n11380 = ~n10882 & ~n11379;
  assign n11381 = ~n11378 & ~n11380;
  assign n11382 = ~po31  & n11374;
  assign n11383 = ~n11381 & ~n11382;
  assign n11384 = ~n11375 & ~n11383;
  assign n11385 = po32  & ~n11384;
  assign n11386 = ~n10887 & ~n10894;
  assign n11387 = n10893 & n11386;
  assign n11388 = po18  & n11387;
  assign n11389 = po18  & n11386;
  assign n11390 = ~n10893 & ~n11389;
  assign n11391 = ~n11388 & ~n11390;
  assign n11392 = ~po32  & ~n11375;
  assign n11393 = ~n11383 & n11392;
  assign n11394 = ~n11391 & ~n11393;
  assign n11395 = ~n11385 & ~n11394;
  assign n11396 = po33  & ~n11395;
  assign n11397 = ~n10897 & ~n10905;
  assign n11398 = n10903 & n11397;
  assign n11399 = po18  & n11398;
  assign n11400 = po18  & n11397;
  assign n11401 = ~n10903 & ~n11400;
  assign n11402 = ~n11399 & ~n11401;
  assign n11403 = ~po33  & n11395;
  assign n11404 = ~n11402 & ~n11403;
  assign n11405 = ~n11396 & ~n11404;
  assign n11406 = po34  & ~n11405;
  assign n11407 = ~n10908 & ~n10915;
  assign n11408 = n10914 & n11407;
  assign n11409 = po18  & n11408;
  assign n11410 = po18  & n11407;
  assign n11411 = ~n10914 & ~n11410;
  assign n11412 = ~n11409 & ~n11411;
  assign n11413 = ~po34  & ~n11396;
  assign n11414 = ~n11404 & n11413;
  assign n11415 = ~n11412 & ~n11414;
  assign n11416 = ~n11406 & ~n11415;
  assign n11417 = po35  & ~n11416;
  assign n11418 = ~n10918 & ~n10926;
  assign n11419 = n10924 & n11418;
  assign n11420 = po18  & n11419;
  assign n11421 = po18  & n11418;
  assign n11422 = ~n10924 & ~n11421;
  assign n11423 = ~n11420 & ~n11422;
  assign n11424 = ~po35  & n11416;
  assign n11425 = ~n11423 & ~n11424;
  assign n11426 = ~n11417 & ~n11425;
  assign n11427 = po36  & ~n11426;
  assign n11428 = ~n10929 & ~n10936;
  assign n11429 = n10935 & n11428;
  assign n11430 = po18  & n11429;
  assign n11431 = po18  & n11428;
  assign n11432 = ~n10935 & ~n11431;
  assign n11433 = ~n11430 & ~n11432;
  assign n11434 = ~po36  & ~n11417;
  assign n11435 = ~n11425 & n11434;
  assign n11436 = ~n11433 & ~n11435;
  assign n11437 = ~n11427 & ~n11436;
  assign n11438 = po37  & ~n11437;
  assign n11439 = ~n10939 & ~n10947;
  assign n11440 = n10945 & n11439;
  assign n11441 = po18  & n11440;
  assign n11442 = po18  & n11439;
  assign n11443 = ~n10945 & ~n11442;
  assign n11444 = ~n11441 & ~n11443;
  assign n11445 = ~po37  & n11437;
  assign n11446 = ~n11444 & ~n11445;
  assign n11447 = ~n11438 & ~n11446;
  assign n11448 = po38  & ~n11447;
  assign n11449 = ~n10950 & ~n10957;
  assign n11450 = n10956 & n11449;
  assign n11451 = po18  & n11450;
  assign n11452 = po18  & n11449;
  assign n11453 = ~n10956 & ~n11452;
  assign n11454 = ~n11451 & ~n11453;
  assign n11455 = ~po38  & ~n11438;
  assign n11456 = ~n11446 & n11455;
  assign n11457 = ~n11454 & ~n11456;
  assign n11458 = ~n11448 & ~n11457;
  assign n11459 = po39  & ~n11458;
  assign n11460 = ~n10960 & ~n10968;
  assign n11461 = n10966 & n11460;
  assign n11462 = po18  & n11461;
  assign n11463 = po18  & n11460;
  assign n11464 = ~n10966 & ~n11463;
  assign n11465 = ~n11462 & ~n11464;
  assign n11466 = ~po39  & n11458;
  assign n11467 = ~n11465 & ~n11466;
  assign n11468 = ~n11459 & ~n11467;
  assign n11469 = po40  & ~n11468;
  assign n11470 = ~n10971 & ~n10978;
  assign n11471 = n10977 & n11470;
  assign n11472 = po18  & n11471;
  assign n11473 = po18  & n11470;
  assign n11474 = ~n10977 & ~n11473;
  assign n11475 = ~n11472 & ~n11474;
  assign n11476 = ~po40  & ~n11459;
  assign n11477 = ~n11467 & n11476;
  assign n11478 = ~n11475 & ~n11477;
  assign n11479 = ~n11469 & ~n11478;
  assign n11480 = po41  & ~n11479;
  assign n11481 = ~n10981 & ~n10989;
  assign n11482 = n10987 & n11481;
  assign n11483 = po18  & n11482;
  assign n11484 = po18  & n11481;
  assign n11485 = ~n10987 & ~n11484;
  assign n11486 = ~n11483 & ~n11485;
  assign n11487 = ~po41  & n11479;
  assign n11488 = ~n11486 & ~n11487;
  assign n11489 = ~n11480 & ~n11488;
  assign n11490 = po42  & ~n11489;
  assign n11491 = ~n10992 & ~n10999;
  assign n11492 = n10998 & n11491;
  assign n11493 = po18  & n11492;
  assign n11494 = po18  & n11491;
  assign n11495 = ~n10998 & ~n11494;
  assign n11496 = ~n11493 & ~n11495;
  assign n11497 = ~po42  & ~n11480;
  assign n11498 = ~n11488 & n11497;
  assign n11499 = ~n11496 & ~n11498;
  assign n11500 = ~n11490 & ~n11499;
  assign n11501 = po43  & ~n11500;
  assign n11502 = ~n11002 & ~n11010;
  assign n11503 = n11008 & n11502;
  assign n11504 = po18  & n11503;
  assign n11505 = po18  & n11502;
  assign n11506 = ~n11008 & ~n11505;
  assign n11507 = ~n11504 & ~n11506;
  assign n11508 = ~po43  & n11500;
  assign n11509 = ~n11507 & ~n11508;
  assign n11510 = ~n11501 & ~n11509;
  assign n11511 = po44  & ~n11510;
  assign n11512 = ~n11013 & ~n11020;
  assign n11513 = n11019 & n11512;
  assign n11514 = po18  & n11513;
  assign n11515 = po18  & n11512;
  assign n11516 = ~n11019 & ~n11515;
  assign n11517 = ~n11514 & ~n11516;
  assign n11518 = ~po44  & ~n11501;
  assign n11519 = ~n11509 & n11518;
  assign n11520 = ~n11517 & ~n11519;
  assign n11521 = ~n11511 & ~n11520;
  assign n11522 = po45  & ~n11521;
  assign n11523 = ~n11023 & ~n11031;
  assign n11524 = n11029 & n11523;
  assign n11525 = po18  & n11524;
  assign n11526 = po18  & n11523;
  assign n11527 = ~n11029 & ~n11526;
  assign n11528 = ~n11525 & ~n11527;
  assign n11529 = ~po45  & n11521;
  assign n11530 = ~n11528 & ~n11529;
  assign n11531 = ~n11522 & ~n11530;
  assign n11532 = po46  & ~n11531;
  assign n11533 = ~n11034 & ~n11041;
  assign n11534 = n11040 & n11533;
  assign n11535 = po18  & n11534;
  assign n11536 = po18  & n11533;
  assign n11537 = ~n11040 & ~n11536;
  assign n11538 = ~n11535 & ~n11537;
  assign n11539 = ~po46  & ~n11522;
  assign n11540 = ~n11530 & n11539;
  assign n11541 = ~n11538 & ~n11540;
  assign n11542 = ~n11532 & ~n11541;
  assign n11543 = po47  & ~n11542;
  assign n11544 = ~n11044 & ~n11046;
  assign n11545 = n11052 & n11544;
  assign n11546 = po18  & n11545;
  assign n11547 = po18  & n11544;
  assign n11548 = ~n11052 & ~n11547;
  assign n11549 = ~n11546 & ~n11548;
  assign n11550 = ~po47  & n11542;
  assign n11551 = ~n11549 & ~n11550;
  assign n11552 = ~n11543 & ~n11551;
  assign n11553 = po48  & ~n11552;
  assign n11554 = ~n11055 & ~n11062;
  assign n11555 = n11061 & n11554;
  assign n11556 = po18  & n11555;
  assign n11557 = po18  & n11554;
  assign n11558 = ~n11061 & ~n11557;
  assign n11559 = ~n11556 & ~n11558;
  assign n11560 = ~po48  & ~n11543;
  assign n11561 = ~n11551 & n11560;
  assign n11562 = ~n11559 & ~n11561;
  assign n11563 = ~n11553 & ~n11562;
  assign n11564 = po49  & ~n11563;
  assign n11565 = ~n11065 & ~n11073;
  assign n11566 = n11071 & n11565;
  assign n11567 = po18  & n11566;
  assign n11568 = po18  & n11565;
  assign n11569 = ~n11071 & ~n11568;
  assign n11570 = ~n11567 & ~n11569;
  assign n11571 = ~po49  & n11563;
  assign n11572 = ~n11570 & ~n11571;
  assign n11573 = ~n11564 & ~n11572;
  assign n11574 = po50  & ~n11573;
  assign n11575 = ~n11076 & ~n11083;
  assign n11576 = n11082 & n11575;
  assign n11577 = po18  & n11576;
  assign n11578 = po18  & n11575;
  assign n11579 = ~n11082 & ~n11578;
  assign n11580 = ~n11577 & ~n11579;
  assign n11581 = ~po50  & ~n11564;
  assign n11582 = ~n11572 & n11581;
  assign n11583 = ~n11580 & ~n11582;
  assign n11584 = ~n11574 & ~n11583;
  assign n11585 = po51  & ~n11584;
  assign n11586 = ~n11086 & ~n11094;
  assign n11587 = n11092 & n11586;
  assign n11588 = po18  & n11587;
  assign n11589 = po18  & n11586;
  assign n11590 = ~n11092 & ~n11589;
  assign n11591 = ~n11588 & ~n11590;
  assign n11592 = ~po51  & n11584;
  assign n11593 = ~n11591 & ~n11592;
  assign n11594 = ~n11585 & ~n11593;
  assign n11595 = po52  & ~n11594;
  assign n11596 = ~n11097 & ~n11104;
  assign n11597 = n11103 & n11596;
  assign n11598 = po18  & n11597;
  assign n11599 = po18  & n11596;
  assign n11600 = ~n11103 & ~n11599;
  assign n11601 = ~n11598 & ~n11600;
  assign n11602 = ~po52  & ~n11585;
  assign n11603 = ~n11593 & n11602;
  assign n11604 = ~n11601 & ~n11603;
  assign n11605 = ~n11595 & ~n11604;
  assign n11606 = po53  & ~n11605;
  assign n11607 = ~n11107 & ~n11115;
  assign n11608 = n11113 & n11607;
  assign n11609 = po18  & n11608;
  assign n11610 = po18  & n11607;
  assign n11611 = ~n11113 & ~n11610;
  assign n11612 = ~n11609 & ~n11611;
  assign n11613 = ~po53  & n11605;
  assign n11614 = ~n11612 & ~n11613;
  assign n11615 = ~n11606 & ~n11614;
  assign n11616 = po54  & ~n11615;
  assign n11617 = ~n11118 & ~n11125;
  assign n11618 = n11124 & n11617;
  assign n11619 = po18  & n11618;
  assign n11620 = po18  & n11617;
  assign n11621 = ~n11124 & ~n11620;
  assign n11622 = ~n11619 & ~n11621;
  assign n11623 = ~po54  & ~n11606;
  assign n11624 = ~n11614 & n11623;
  assign n11625 = ~n11622 & ~n11624;
  assign n11626 = ~n11616 & ~n11625;
  assign n11627 = po55  & ~n11626;
  assign n11628 = ~n11128 & ~n11136;
  assign n11629 = n11134 & n11628;
  assign n11630 = po18  & n11629;
  assign n11631 = po18  & n11628;
  assign n11632 = ~n11134 & ~n11631;
  assign n11633 = ~n11630 & ~n11632;
  assign n11634 = ~po55  & n11626;
  assign n11635 = ~n11633 & ~n11634;
  assign n11636 = ~n11627 & ~n11635;
  assign n11637 = po56  & ~n11636;
  assign n11638 = ~n11139 & ~n11146;
  assign n11639 = n11145 & n11638;
  assign n11640 = po18  & n11639;
  assign n11641 = po18  & n11638;
  assign n11642 = ~n11145 & ~n11641;
  assign n11643 = ~n11640 & ~n11642;
  assign n11644 = ~po56  & ~n11627;
  assign n11645 = ~n11635 & n11644;
  assign n11646 = ~n11643 & ~n11645;
  assign n11647 = ~n11637 & ~n11646;
  assign n11648 = po57  & ~n11647;
  assign n11649 = ~n11149 & ~n11157;
  assign n11650 = n11155 & n11649;
  assign n11651 = po18  & n11650;
  assign n11652 = po18  & n11649;
  assign n11653 = ~n11155 & ~n11652;
  assign n11654 = ~n11651 & ~n11653;
  assign n11655 = ~po57  & n11647;
  assign n11656 = ~n11654 & ~n11655;
  assign n11657 = ~n11648 & ~n11656;
  assign n11658 = po58  & ~n11657;
  assign n11659 = ~n11160 & ~n11167;
  assign n11660 = n11166 & n11659;
  assign n11661 = po18  & n11660;
  assign n11662 = po18  & n11659;
  assign n11663 = ~n11166 & ~n11662;
  assign n11664 = ~n11661 & ~n11663;
  assign n11665 = ~po58  & ~n11648;
  assign n11666 = ~n11656 & n11665;
  assign n11667 = ~n11664 & ~n11666;
  assign n11668 = ~n11658 & ~n11667;
  assign n11669 = po59  & ~n11668;
  assign n11670 = ~n11170 & ~n11178;
  assign n11671 = n11176 & n11670;
  assign n11672 = po18  & n11671;
  assign n11673 = po18  & n11670;
  assign n11674 = ~n11176 & ~n11673;
  assign n11675 = ~n11672 & ~n11674;
  assign n11676 = ~po59  & n11668;
  assign n11677 = ~n11675 & ~n11676;
  assign n11678 = ~n11669 & ~n11677;
  assign n11679 = po60  & ~n11678;
  assign n11680 = ~n11181 & ~n11188;
  assign n11681 = n11187 & n11680;
  assign n11682 = po18  & n11681;
  assign n11683 = po18  & n11680;
  assign n11684 = ~n11187 & ~n11683;
  assign n11685 = ~n11682 & ~n11684;
  assign n11686 = ~po60  & ~n11669;
  assign n11687 = ~n11677 & n11686;
  assign n11688 = ~n11685 & ~n11687;
  assign n11689 = ~n11679 & ~n11688;
  assign n11690 = po61  & ~n11689;
  assign n11691 = ~n11191 & ~n11199;
  assign n11692 = n11197 & n11691;
  assign n11693 = po18  & n11692;
  assign n11694 = po18  & n11691;
  assign n11695 = ~n11197 & ~n11694;
  assign n11696 = ~n11693 & ~n11695;
  assign n11697 = ~po61  & n11689;
  assign n11698 = ~n11696 & ~n11697;
  assign n11699 = ~n11690 & ~n11698;
  assign n11700 = po62  & ~n11699;
  assign n11701 = ~n11202 & ~n11209;
  assign n11702 = n11208 & n11701;
  assign n11703 = po18  & n11702;
  assign n11704 = po18  & n11701;
  assign n11705 = ~n11208 & ~n11704;
  assign n11706 = ~n11703 & ~n11705;
  assign n11707 = ~po62  & ~n11690;
  assign n11708 = ~n11698 & n11707;
  assign n11709 = ~n11706 & ~n11708;
  assign n11710 = ~n11700 & ~n11709;
  assign n11711 = ~n11212 & ~n11220;
  assign n11712 = po18  & n11711;
  assign n11713 = ~n11218 & ~n11712;
  assign n11714 = n11218 & n11712;
  assign n11715 = ~n11713 & ~n11714;
  assign n11716 = ~n11222 & ~n11227;
  assign n11717 = po18  & n11716;
  assign n11718 = ~n11240 & ~n11717;
  assign n11719 = ~n11715 & n11718;
  assign n11720 = ~n11710 & n11719;
  assign n11721 = ~po63  & ~n11720;
  assign n11722 = ~n11227 & po18 ;
  assign n11723 = n11222 & ~n11722;
  assign n11724 = po63  & ~n11716;
  assign n11725 = ~n11723 & n11724;
  assign n11726 = n11227 & ~po18 ;
  assign n11727 = ~n11725 & ~n11726;
  assign n11728 = n11710 & n11715;
  assign n11729 = n11727 & ~n11728;
  assign po17  = n11721 | ~n11729;
  assign n11731 = pi34  & po17 ;
  assign n11732 = ~pi32  & ~pi33 ;
  assign n11733 = ~pi34  & n11732;
  assign n11734 = ~n11731 & ~n11733;
  assign n11735 = po18  & ~n11734;
  assign n11736 = n11239 & ~n11733;
  assign n11737 = ~n11240 & n11736;
  assign n11738 = ~n11233 & n11737;
  assign n11739 = ~n11731 & n11738;
  assign n11740 = ~pi34  & po17 ;
  assign n11741 = pi35  & ~n11740;
  assign n11742 = n11244 & po17 ;
  assign n11743 = ~n11741 & ~n11742;
  assign n11744 = ~n11739 & n11743;
  assign n11745 = ~n11735 & ~n11744;
  assign n11746 = po19  & ~n11745;
  assign n11747 = po18  & n11727;
  assign n11748 = ~n11728 & n11747;
  assign n11749 = ~n11721 & n11748;
  assign n11750 = ~n11742 & ~n11749;
  assign n11751 = pi36  & ~n11750;
  assign n11752 = ~pi36  & n11750;
  assign n11753 = ~n11751 & ~n11752;
  assign n11754 = ~po19  & n11745;
  assign n11755 = ~n11753 & ~n11754;
  assign n11756 = ~n11746 & ~n11755;
  assign n11757 = po20  & ~n11756;
  assign n11758 = ~n11247 & ~n11251;
  assign n11759 = ~n11255 & n11758;
  assign n11760 = po17  & n11759;
  assign n11761 = po17  & n11758;
  assign n11762 = n11255 & ~n11761;
  assign n11763 = ~n11760 & ~n11762;
  assign n11764 = ~po20  & ~n11746;
  assign n11765 = ~n11755 & n11764;
  assign n11766 = ~n11763 & ~n11765;
  assign n11767 = ~n11757 & ~n11766;
  assign n11768 = po21  & ~n11767;
  assign n11769 = ~n11258 & ~n11260;
  assign n11770 = n11267 & n11769;
  assign n11771 = po17  & n11770;
  assign n11772 = po17  & n11769;
  assign n11773 = ~n11267 & ~n11772;
  assign n11774 = ~n11771 & ~n11773;
  assign n11775 = ~po21  & n11767;
  assign n11776 = ~n11774 & ~n11775;
  assign n11777 = ~n11768 & ~n11776;
  assign n11778 = po22  & ~n11777;
  assign n11779 = ~n11270 & ~n11277;
  assign n11780 = n11276 & n11779;
  assign n11781 = po17  & n11780;
  assign n11782 = po17  & n11779;
  assign n11783 = ~n11276 & ~n11782;
  assign n11784 = ~n11781 & ~n11783;
  assign n11785 = ~po22  & ~n11768;
  assign n11786 = ~n11776 & n11785;
  assign n11787 = ~n11784 & ~n11786;
  assign n11788 = ~n11778 & ~n11787;
  assign n11789 = po23  & ~n11788;
  assign n11790 = ~n11280 & ~n11288;
  assign n11791 = n11286 & n11790;
  assign n11792 = po17  & n11791;
  assign n11793 = po17  & n11790;
  assign n11794 = ~n11286 & ~n11793;
  assign n11795 = ~n11792 & ~n11794;
  assign n11796 = ~po23  & n11788;
  assign n11797 = ~n11795 & ~n11796;
  assign n11798 = ~n11789 & ~n11797;
  assign n11799 = po24  & ~n11798;
  assign n11800 = ~n11291 & ~n11298;
  assign n11801 = n11297 & n11800;
  assign n11802 = po17  & n11801;
  assign n11803 = po17  & n11800;
  assign n11804 = ~n11297 & ~n11803;
  assign n11805 = ~n11802 & ~n11804;
  assign n11806 = ~po24  & ~n11789;
  assign n11807 = ~n11797 & n11806;
  assign n11808 = ~n11805 & ~n11807;
  assign n11809 = ~n11799 & ~n11808;
  assign n11810 = po25  & ~n11809;
  assign n11811 = ~n11301 & ~n11309;
  assign n11812 = n11307 & n11811;
  assign n11813 = po17  & n11812;
  assign n11814 = po17  & n11811;
  assign n11815 = ~n11307 & ~n11814;
  assign n11816 = ~n11813 & ~n11815;
  assign n11817 = ~po25  & n11809;
  assign n11818 = ~n11816 & ~n11817;
  assign n11819 = ~n11810 & ~n11818;
  assign n11820 = po26  & ~n11819;
  assign n11821 = ~n11312 & ~n11319;
  assign n11822 = n11318 & n11821;
  assign n11823 = po17  & n11822;
  assign n11824 = po17  & n11821;
  assign n11825 = ~n11318 & ~n11824;
  assign n11826 = ~n11823 & ~n11825;
  assign n11827 = ~po26  & ~n11810;
  assign n11828 = ~n11818 & n11827;
  assign n11829 = ~n11826 & ~n11828;
  assign n11830 = ~n11820 & ~n11829;
  assign n11831 = po27  & ~n11830;
  assign n11832 = ~n11322 & ~n11330;
  assign n11833 = n11328 & n11832;
  assign n11834 = po17  & n11833;
  assign n11835 = po17  & n11832;
  assign n11836 = ~n11328 & ~n11835;
  assign n11837 = ~n11834 & ~n11836;
  assign n11838 = ~po27  & n11830;
  assign n11839 = ~n11837 & ~n11838;
  assign n11840 = ~n11831 & ~n11839;
  assign n11841 = po28  & ~n11840;
  assign n11842 = ~n11333 & ~n11340;
  assign n11843 = n11339 & n11842;
  assign n11844 = po17  & n11843;
  assign n11845 = po17  & n11842;
  assign n11846 = ~n11339 & ~n11845;
  assign n11847 = ~n11844 & ~n11846;
  assign n11848 = ~po28  & ~n11831;
  assign n11849 = ~n11839 & n11848;
  assign n11850 = ~n11847 & ~n11849;
  assign n11851 = ~n11841 & ~n11850;
  assign n11852 = po29  & ~n11851;
  assign n11853 = ~n11343 & ~n11351;
  assign n11854 = n11349 & n11853;
  assign n11855 = po17  & n11854;
  assign n11856 = po17  & n11853;
  assign n11857 = ~n11349 & ~n11856;
  assign n11858 = ~n11855 & ~n11857;
  assign n11859 = ~po29  & n11851;
  assign n11860 = ~n11858 & ~n11859;
  assign n11861 = ~n11852 & ~n11860;
  assign n11862 = po30  & ~n11861;
  assign n11863 = ~n11354 & ~n11361;
  assign n11864 = n11360 & n11863;
  assign n11865 = po17  & n11864;
  assign n11866 = po17  & n11863;
  assign n11867 = ~n11360 & ~n11866;
  assign n11868 = ~n11865 & ~n11867;
  assign n11869 = ~po30  & ~n11852;
  assign n11870 = ~n11860 & n11869;
  assign n11871 = ~n11868 & ~n11870;
  assign n11872 = ~n11862 & ~n11871;
  assign n11873 = po31  & ~n11872;
  assign n11874 = ~n11364 & ~n11372;
  assign n11875 = n11370 & n11874;
  assign n11876 = po17  & n11875;
  assign n11877 = po17  & n11874;
  assign n11878 = ~n11370 & ~n11877;
  assign n11879 = ~n11876 & ~n11878;
  assign n11880 = ~po31  & n11872;
  assign n11881 = ~n11879 & ~n11880;
  assign n11882 = ~n11873 & ~n11881;
  assign n11883 = po32  & ~n11882;
  assign n11884 = ~n11375 & ~n11382;
  assign n11885 = n11381 & n11884;
  assign n11886 = po17  & n11885;
  assign n11887 = po17  & n11884;
  assign n11888 = ~n11381 & ~n11887;
  assign n11889 = ~n11886 & ~n11888;
  assign n11890 = ~po32  & ~n11873;
  assign n11891 = ~n11881 & n11890;
  assign n11892 = ~n11889 & ~n11891;
  assign n11893 = ~n11883 & ~n11892;
  assign n11894 = po33  & ~n11893;
  assign n11895 = ~n11385 & ~n11393;
  assign n11896 = n11391 & n11895;
  assign n11897 = po17  & n11896;
  assign n11898 = po17  & n11895;
  assign n11899 = ~n11391 & ~n11898;
  assign n11900 = ~n11897 & ~n11899;
  assign n11901 = ~po33  & n11893;
  assign n11902 = ~n11900 & ~n11901;
  assign n11903 = ~n11894 & ~n11902;
  assign n11904 = po34  & ~n11903;
  assign n11905 = ~n11396 & ~n11403;
  assign n11906 = n11402 & n11905;
  assign n11907 = po17  & n11906;
  assign n11908 = po17  & n11905;
  assign n11909 = ~n11402 & ~n11908;
  assign n11910 = ~n11907 & ~n11909;
  assign n11911 = ~po34  & ~n11894;
  assign n11912 = ~n11902 & n11911;
  assign n11913 = ~n11910 & ~n11912;
  assign n11914 = ~n11904 & ~n11913;
  assign n11915 = po35  & ~n11914;
  assign n11916 = ~n11406 & ~n11414;
  assign n11917 = n11412 & n11916;
  assign n11918 = po17  & n11917;
  assign n11919 = po17  & n11916;
  assign n11920 = ~n11412 & ~n11919;
  assign n11921 = ~n11918 & ~n11920;
  assign n11922 = ~po35  & n11914;
  assign n11923 = ~n11921 & ~n11922;
  assign n11924 = ~n11915 & ~n11923;
  assign n11925 = po36  & ~n11924;
  assign n11926 = ~n11417 & ~n11424;
  assign n11927 = n11423 & n11926;
  assign n11928 = po17  & n11927;
  assign n11929 = po17  & n11926;
  assign n11930 = ~n11423 & ~n11929;
  assign n11931 = ~n11928 & ~n11930;
  assign n11932 = ~po36  & ~n11915;
  assign n11933 = ~n11923 & n11932;
  assign n11934 = ~n11931 & ~n11933;
  assign n11935 = ~n11925 & ~n11934;
  assign n11936 = po37  & ~n11935;
  assign n11937 = ~n11427 & ~n11435;
  assign n11938 = n11433 & n11937;
  assign n11939 = po17  & n11938;
  assign n11940 = po17  & n11937;
  assign n11941 = ~n11433 & ~n11940;
  assign n11942 = ~n11939 & ~n11941;
  assign n11943 = ~po37  & n11935;
  assign n11944 = ~n11942 & ~n11943;
  assign n11945 = ~n11936 & ~n11944;
  assign n11946 = po38  & ~n11945;
  assign n11947 = ~n11438 & ~n11445;
  assign n11948 = n11444 & n11947;
  assign n11949 = po17  & n11948;
  assign n11950 = po17  & n11947;
  assign n11951 = ~n11444 & ~n11950;
  assign n11952 = ~n11949 & ~n11951;
  assign n11953 = ~po38  & ~n11936;
  assign n11954 = ~n11944 & n11953;
  assign n11955 = ~n11952 & ~n11954;
  assign n11956 = ~n11946 & ~n11955;
  assign n11957 = po39  & ~n11956;
  assign n11958 = ~n11448 & ~n11456;
  assign n11959 = n11454 & n11958;
  assign n11960 = po17  & n11959;
  assign n11961 = po17  & n11958;
  assign n11962 = ~n11454 & ~n11961;
  assign n11963 = ~n11960 & ~n11962;
  assign n11964 = ~po39  & n11956;
  assign n11965 = ~n11963 & ~n11964;
  assign n11966 = ~n11957 & ~n11965;
  assign n11967 = po40  & ~n11966;
  assign n11968 = ~n11459 & ~n11466;
  assign n11969 = n11465 & n11968;
  assign n11970 = po17  & n11969;
  assign n11971 = po17  & n11968;
  assign n11972 = ~n11465 & ~n11971;
  assign n11973 = ~n11970 & ~n11972;
  assign n11974 = ~po40  & ~n11957;
  assign n11975 = ~n11965 & n11974;
  assign n11976 = ~n11973 & ~n11975;
  assign n11977 = ~n11967 & ~n11976;
  assign n11978 = po41  & ~n11977;
  assign n11979 = ~n11469 & ~n11477;
  assign n11980 = n11475 & n11979;
  assign n11981 = po17  & n11980;
  assign n11982 = po17  & n11979;
  assign n11983 = ~n11475 & ~n11982;
  assign n11984 = ~n11981 & ~n11983;
  assign n11985 = ~po41  & n11977;
  assign n11986 = ~n11984 & ~n11985;
  assign n11987 = ~n11978 & ~n11986;
  assign n11988 = po42  & ~n11987;
  assign n11989 = ~n11480 & ~n11487;
  assign n11990 = n11486 & n11989;
  assign n11991 = po17  & n11990;
  assign n11992 = po17  & n11989;
  assign n11993 = ~n11486 & ~n11992;
  assign n11994 = ~n11991 & ~n11993;
  assign n11995 = ~po42  & ~n11978;
  assign n11996 = ~n11986 & n11995;
  assign n11997 = ~n11994 & ~n11996;
  assign n11998 = ~n11988 & ~n11997;
  assign n11999 = po43  & ~n11998;
  assign n12000 = ~n11490 & ~n11498;
  assign n12001 = n11496 & n12000;
  assign n12002 = po17  & n12001;
  assign n12003 = po17  & n12000;
  assign n12004 = ~n11496 & ~n12003;
  assign n12005 = ~n12002 & ~n12004;
  assign n12006 = ~po43  & n11998;
  assign n12007 = ~n12005 & ~n12006;
  assign n12008 = ~n11999 & ~n12007;
  assign n12009 = po44  & ~n12008;
  assign n12010 = ~n11501 & ~n11508;
  assign n12011 = n11507 & n12010;
  assign n12012 = po17  & n12011;
  assign n12013 = po17  & n12010;
  assign n12014 = ~n11507 & ~n12013;
  assign n12015 = ~n12012 & ~n12014;
  assign n12016 = ~po44  & ~n11999;
  assign n12017 = ~n12007 & n12016;
  assign n12018 = ~n12015 & ~n12017;
  assign n12019 = ~n12009 & ~n12018;
  assign n12020 = po45  & ~n12019;
  assign n12021 = ~n11511 & ~n11519;
  assign n12022 = n11517 & n12021;
  assign n12023 = po17  & n12022;
  assign n12024 = po17  & n12021;
  assign n12025 = ~n11517 & ~n12024;
  assign n12026 = ~n12023 & ~n12025;
  assign n12027 = ~po45  & n12019;
  assign n12028 = ~n12026 & ~n12027;
  assign n12029 = ~n12020 & ~n12028;
  assign n12030 = po46  & ~n12029;
  assign n12031 = ~n11522 & ~n11529;
  assign n12032 = n11528 & n12031;
  assign n12033 = po17  & n12032;
  assign n12034 = po17  & n12031;
  assign n12035 = ~n11528 & ~n12034;
  assign n12036 = ~n12033 & ~n12035;
  assign n12037 = ~po46  & ~n12020;
  assign n12038 = ~n12028 & n12037;
  assign n12039 = ~n12036 & ~n12038;
  assign n12040 = ~n12030 & ~n12039;
  assign n12041 = po47  & ~n12040;
  assign n12042 = ~n11532 & ~n11540;
  assign n12043 = n11538 & n12042;
  assign n12044 = po17  & n12043;
  assign n12045 = po17  & n12042;
  assign n12046 = ~n11538 & ~n12045;
  assign n12047 = ~n12044 & ~n12046;
  assign n12048 = ~po47  & n12040;
  assign n12049 = ~n12047 & ~n12048;
  assign n12050 = ~n12041 & ~n12049;
  assign n12051 = po48  & ~n12050;
  assign n12052 = ~po48  & ~n12041;
  assign n12053 = ~n12049 & n12052;
  assign n12054 = ~n11543 & ~n11550;
  assign n12055 = n11549 & n12054;
  assign n12056 = po17  & n12055;
  assign n12057 = po17  & n12054;
  assign n12058 = ~n11549 & ~n12057;
  assign n12059 = ~n12056 & ~n12058;
  assign n12060 = ~n12053 & ~n12059;
  assign n12061 = ~n12051 & ~n12060;
  assign n12062 = po49  & ~n12061;
  assign n12063 = ~n11553 & ~n11561;
  assign n12064 = n11559 & n12063;
  assign n12065 = po17  & n12064;
  assign n12066 = po17  & n12063;
  assign n12067 = ~n11559 & ~n12066;
  assign n12068 = ~n12065 & ~n12067;
  assign n12069 = ~po49  & n12061;
  assign n12070 = ~n12068 & ~n12069;
  assign n12071 = ~n12062 & ~n12070;
  assign n12072 = po50  & ~n12071;
  assign n12073 = ~n11564 & ~n11571;
  assign n12074 = n11570 & n12073;
  assign n12075 = po17  & n12074;
  assign n12076 = po17  & n12073;
  assign n12077 = ~n11570 & ~n12076;
  assign n12078 = ~n12075 & ~n12077;
  assign n12079 = ~po50  & ~n12062;
  assign n12080 = ~n12070 & n12079;
  assign n12081 = ~n12078 & ~n12080;
  assign n12082 = ~n12072 & ~n12081;
  assign n12083 = po51  & ~n12082;
  assign n12084 = ~n11574 & ~n11582;
  assign n12085 = n11580 & n12084;
  assign n12086 = po17  & n12085;
  assign n12087 = po17  & n12084;
  assign n12088 = ~n11580 & ~n12087;
  assign n12089 = ~n12086 & ~n12088;
  assign n12090 = ~po51  & n12082;
  assign n12091 = ~n12089 & ~n12090;
  assign n12092 = ~n12083 & ~n12091;
  assign n12093 = po52  & ~n12092;
  assign n12094 = ~n11585 & ~n11592;
  assign n12095 = n11591 & n12094;
  assign n12096 = po17  & n12095;
  assign n12097 = po17  & n12094;
  assign n12098 = ~n11591 & ~n12097;
  assign n12099 = ~n12096 & ~n12098;
  assign n12100 = ~po52  & ~n12083;
  assign n12101 = ~n12091 & n12100;
  assign n12102 = ~n12099 & ~n12101;
  assign n12103 = ~n12093 & ~n12102;
  assign n12104 = po53  & ~n12103;
  assign n12105 = ~n11595 & ~n11603;
  assign n12106 = n11601 & n12105;
  assign n12107 = po17  & n12106;
  assign n12108 = po17  & n12105;
  assign n12109 = ~n11601 & ~n12108;
  assign n12110 = ~n12107 & ~n12109;
  assign n12111 = ~po53  & n12103;
  assign n12112 = ~n12110 & ~n12111;
  assign n12113 = ~n12104 & ~n12112;
  assign n12114 = po54  & ~n12113;
  assign n12115 = ~n11606 & ~n11613;
  assign n12116 = n11612 & n12115;
  assign n12117 = po17  & n12116;
  assign n12118 = po17  & n12115;
  assign n12119 = ~n11612 & ~n12118;
  assign n12120 = ~n12117 & ~n12119;
  assign n12121 = ~po54  & ~n12104;
  assign n12122 = ~n12112 & n12121;
  assign n12123 = ~n12120 & ~n12122;
  assign n12124 = ~n12114 & ~n12123;
  assign n12125 = po55  & ~n12124;
  assign n12126 = ~n11616 & ~n11624;
  assign n12127 = n11622 & n12126;
  assign n12128 = po17  & n12127;
  assign n12129 = po17  & n12126;
  assign n12130 = ~n11622 & ~n12129;
  assign n12131 = ~n12128 & ~n12130;
  assign n12132 = ~po55  & n12124;
  assign n12133 = ~n12131 & ~n12132;
  assign n12134 = ~n12125 & ~n12133;
  assign n12135 = po56  & ~n12134;
  assign n12136 = ~n11627 & ~n11634;
  assign n12137 = n11633 & n12136;
  assign n12138 = po17  & n12137;
  assign n12139 = po17  & n12136;
  assign n12140 = ~n11633 & ~n12139;
  assign n12141 = ~n12138 & ~n12140;
  assign n12142 = ~po56  & ~n12125;
  assign n12143 = ~n12133 & n12142;
  assign n12144 = ~n12141 & ~n12143;
  assign n12145 = ~n12135 & ~n12144;
  assign n12146 = po57  & ~n12145;
  assign n12147 = ~n11637 & ~n11645;
  assign n12148 = n11643 & n12147;
  assign n12149 = po17  & n12148;
  assign n12150 = po17  & n12147;
  assign n12151 = ~n11643 & ~n12150;
  assign n12152 = ~n12149 & ~n12151;
  assign n12153 = ~po57  & n12145;
  assign n12154 = ~n12152 & ~n12153;
  assign n12155 = ~n12146 & ~n12154;
  assign n12156 = po58  & ~n12155;
  assign n12157 = ~n11648 & ~n11655;
  assign n12158 = n11654 & n12157;
  assign n12159 = po17  & n12158;
  assign n12160 = po17  & n12157;
  assign n12161 = ~n11654 & ~n12160;
  assign n12162 = ~n12159 & ~n12161;
  assign n12163 = ~po58  & ~n12146;
  assign n12164 = ~n12154 & n12163;
  assign n12165 = ~n12162 & ~n12164;
  assign n12166 = ~n12156 & ~n12165;
  assign n12167 = po59  & ~n12166;
  assign n12168 = ~n11658 & ~n11666;
  assign n12169 = n11664 & n12168;
  assign n12170 = po17  & n12169;
  assign n12171 = po17  & n12168;
  assign n12172 = ~n11664 & ~n12171;
  assign n12173 = ~n12170 & ~n12172;
  assign n12174 = ~po59  & n12166;
  assign n12175 = ~n12173 & ~n12174;
  assign n12176 = ~n12167 & ~n12175;
  assign n12177 = po60  & ~n12176;
  assign n12178 = ~n11669 & ~n11676;
  assign n12179 = n11675 & n12178;
  assign n12180 = po17  & n12179;
  assign n12181 = po17  & n12178;
  assign n12182 = ~n11675 & ~n12181;
  assign n12183 = ~n12180 & ~n12182;
  assign n12184 = ~po60  & ~n12167;
  assign n12185 = ~n12175 & n12184;
  assign n12186 = ~n12183 & ~n12185;
  assign n12187 = ~n12177 & ~n12186;
  assign n12188 = po61  & ~n12187;
  assign n12189 = ~n11679 & ~n11687;
  assign n12190 = n11685 & n12189;
  assign n12191 = po17  & n12190;
  assign n12192 = po17  & n12189;
  assign n12193 = ~n11685 & ~n12192;
  assign n12194 = ~n12191 & ~n12193;
  assign n12195 = ~po61  & n12187;
  assign n12196 = ~n12194 & ~n12195;
  assign n12197 = ~n12188 & ~n12196;
  assign n12198 = po62  & ~n12197;
  assign n12199 = ~n11690 & ~n11697;
  assign n12200 = n11696 & n12199;
  assign n12201 = po17  & n12200;
  assign n12202 = po17  & n12199;
  assign n12203 = ~n11696 & ~n12202;
  assign n12204 = ~n12201 & ~n12203;
  assign n12205 = ~po62  & ~n12188;
  assign n12206 = ~n12196 & n12205;
  assign n12207 = ~n12204 & ~n12206;
  assign n12208 = ~n12198 & ~n12207;
  assign n12209 = ~n11700 & ~n11708;
  assign n12210 = po17  & n12209;
  assign n12211 = ~n11706 & ~n12210;
  assign n12212 = n11706 & n12210;
  assign n12213 = ~n12211 & ~n12212;
  assign n12214 = ~n11710 & ~n11715;
  assign n12215 = po17  & n12214;
  assign n12216 = ~n11728 & ~n12215;
  assign n12217 = ~n12213 & n12216;
  assign n12218 = ~n12208 & n12217;
  assign n12219 = ~po63  & ~n12218;
  assign n12220 = ~n11715 & po17 ;
  assign n12221 = n11710 & ~n12220;
  assign n12222 = po63  & ~n12214;
  assign n12223 = ~n12221 & n12222;
  assign n12224 = n11715 & ~po17 ;
  assign n12225 = ~n12223 & ~n12224;
  assign n12226 = n12208 & n12213;
  assign n12227 = n12225 & ~n12226;
  assign po16  = n12219 | ~n12227;
  assign n12229 = pi32  & po16 ;
  assign n12230 = ~pi30  & ~pi31 ;
  assign n12231 = ~pi32  & n12230;
  assign n12232 = ~n12229 & ~n12231;
  assign n12233 = po17  & ~n12232;
  assign n12234 = n11727 & ~n12231;
  assign n12235 = ~n11728 & n12234;
  assign n12236 = ~n11721 & n12235;
  assign n12237 = ~n12229 & n12236;
  assign n12238 = ~pi32  & po16 ;
  assign n12239 = pi33  & ~n12238;
  assign n12240 = n11732 & po16 ;
  assign n12241 = ~n12239 & ~n12240;
  assign n12242 = ~n12237 & n12241;
  assign n12243 = ~n12233 & ~n12242;
  assign n12244 = po18  & ~n12243;
  assign n12245 = ~po18  & ~n12233;
  assign n12246 = ~n12242 & n12245;
  assign n12247 = po17  & n12225;
  assign n12248 = ~n12226 & n12247;
  assign n12249 = ~n12219 & n12248;
  assign n12250 = ~n12240 & ~n12249;
  assign n12251 = pi34  & ~n12250;
  assign n12252 = ~pi34  & n12250;
  assign n12253 = ~n12251 & ~n12252;
  assign n12254 = ~n12246 & ~n12253;
  assign n12255 = ~n12244 & ~n12254;
  assign n12256 = po19  & ~n12255;
  assign n12257 = ~n11735 & ~n11739;
  assign n12258 = ~n11743 & n12257;
  assign n12259 = po16  & n12258;
  assign n12260 = po16  & n12257;
  assign n12261 = n11743 & ~n12260;
  assign n12262 = ~n12259 & ~n12261;
  assign n12263 = ~po19  & n12255;
  assign n12264 = ~n12262 & ~n12263;
  assign n12265 = ~n12256 & ~n12264;
  assign n12266 = po20  & ~n12265;
  assign n12267 = ~n11746 & ~n11754;
  assign n12268 = n11753 & n12267;
  assign n12269 = po16  & n12268;
  assign n12270 = po16  & n12267;
  assign n12271 = ~n11753 & ~n12270;
  assign n12272 = ~n12269 & ~n12271;
  assign n12273 = ~po20  & ~n12256;
  assign n12274 = ~n12264 & n12273;
  assign n12275 = ~n12272 & ~n12274;
  assign n12276 = ~n12266 & ~n12275;
  assign n12277 = po21  & ~n12276;
  assign n12278 = ~n11757 & ~n11765;
  assign n12279 = n11763 & n12278;
  assign n12280 = po16  & n12279;
  assign n12281 = po16  & n12278;
  assign n12282 = ~n11763 & ~n12281;
  assign n12283 = ~n12280 & ~n12282;
  assign n12284 = ~po21  & n12276;
  assign n12285 = ~n12283 & ~n12284;
  assign n12286 = ~n12277 & ~n12285;
  assign n12287 = po22  & ~n12286;
  assign n12288 = ~n11768 & ~n11775;
  assign n12289 = n11774 & n12288;
  assign n12290 = po16  & n12289;
  assign n12291 = po16  & n12288;
  assign n12292 = ~n11774 & ~n12291;
  assign n12293 = ~n12290 & ~n12292;
  assign n12294 = ~po22  & ~n12277;
  assign n12295 = ~n12285 & n12294;
  assign n12296 = ~n12293 & ~n12295;
  assign n12297 = ~n12287 & ~n12296;
  assign n12298 = po23  & ~n12297;
  assign n12299 = ~n11778 & ~n11786;
  assign n12300 = n11784 & n12299;
  assign n12301 = po16  & n12300;
  assign n12302 = po16  & n12299;
  assign n12303 = ~n11784 & ~n12302;
  assign n12304 = ~n12301 & ~n12303;
  assign n12305 = ~po23  & n12297;
  assign n12306 = ~n12304 & ~n12305;
  assign n12307 = ~n12298 & ~n12306;
  assign n12308 = po24  & ~n12307;
  assign n12309 = ~n11789 & ~n11796;
  assign n12310 = n11795 & n12309;
  assign n12311 = po16  & n12310;
  assign n12312 = po16  & n12309;
  assign n12313 = ~n11795 & ~n12312;
  assign n12314 = ~n12311 & ~n12313;
  assign n12315 = ~po24  & ~n12298;
  assign n12316 = ~n12306 & n12315;
  assign n12317 = ~n12314 & ~n12316;
  assign n12318 = ~n12308 & ~n12317;
  assign n12319 = po25  & ~n12318;
  assign n12320 = ~n11799 & ~n11807;
  assign n12321 = n11805 & n12320;
  assign n12322 = po16  & n12321;
  assign n12323 = po16  & n12320;
  assign n12324 = ~n11805 & ~n12323;
  assign n12325 = ~n12322 & ~n12324;
  assign n12326 = ~po25  & n12318;
  assign n12327 = ~n12325 & ~n12326;
  assign n12328 = ~n12319 & ~n12327;
  assign n12329 = po26  & ~n12328;
  assign n12330 = ~n11810 & ~n11817;
  assign n12331 = n11816 & n12330;
  assign n12332 = po16  & n12331;
  assign n12333 = po16  & n12330;
  assign n12334 = ~n11816 & ~n12333;
  assign n12335 = ~n12332 & ~n12334;
  assign n12336 = ~po26  & ~n12319;
  assign n12337 = ~n12327 & n12336;
  assign n12338 = ~n12335 & ~n12337;
  assign n12339 = ~n12329 & ~n12338;
  assign n12340 = po27  & ~n12339;
  assign n12341 = ~n11820 & ~n11828;
  assign n12342 = n11826 & n12341;
  assign n12343 = po16  & n12342;
  assign n12344 = po16  & n12341;
  assign n12345 = ~n11826 & ~n12344;
  assign n12346 = ~n12343 & ~n12345;
  assign n12347 = ~po27  & n12339;
  assign n12348 = ~n12346 & ~n12347;
  assign n12349 = ~n12340 & ~n12348;
  assign n12350 = po28  & ~n12349;
  assign n12351 = ~n11831 & ~n11838;
  assign n12352 = n11837 & n12351;
  assign n12353 = po16  & n12352;
  assign n12354 = po16  & n12351;
  assign n12355 = ~n11837 & ~n12354;
  assign n12356 = ~n12353 & ~n12355;
  assign n12357 = ~po28  & ~n12340;
  assign n12358 = ~n12348 & n12357;
  assign n12359 = ~n12356 & ~n12358;
  assign n12360 = ~n12350 & ~n12359;
  assign n12361 = po29  & ~n12360;
  assign n12362 = ~n11841 & ~n11849;
  assign n12363 = n11847 & n12362;
  assign n12364 = po16  & n12363;
  assign n12365 = po16  & n12362;
  assign n12366 = ~n11847 & ~n12365;
  assign n12367 = ~n12364 & ~n12366;
  assign n12368 = ~po29  & n12360;
  assign n12369 = ~n12367 & ~n12368;
  assign n12370 = ~n12361 & ~n12369;
  assign n12371 = po30  & ~n12370;
  assign n12372 = ~n11852 & ~n11859;
  assign n12373 = n11858 & n12372;
  assign n12374 = po16  & n12373;
  assign n12375 = po16  & n12372;
  assign n12376 = ~n11858 & ~n12375;
  assign n12377 = ~n12374 & ~n12376;
  assign n12378 = ~po30  & ~n12361;
  assign n12379 = ~n12369 & n12378;
  assign n12380 = ~n12377 & ~n12379;
  assign n12381 = ~n12371 & ~n12380;
  assign n12382 = po31  & ~n12381;
  assign n12383 = ~n11862 & ~n11870;
  assign n12384 = n11868 & n12383;
  assign n12385 = po16  & n12384;
  assign n12386 = po16  & n12383;
  assign n12387 = ~n11868 & ~n12386;
  assign n12388 = ~n12385 & ~n12387;
  assign n12389 = ~po31  & n12381;
  assign n12390 = ~n12388 & ~n12389;
  assign n12391 = ~n12382 & ~n12390;
  assign n12392 = po32  & ~n12391;
  assign n12393 = ~n11873 & ~n11880;
  assign n12394 = n11879 & n12393;
  assign n12395 = po16  & n12394;
  assign n12396 = po16  & n12393;
  assign n12397 = ~n11879 & ~n12396;
  assign n12398 = ~n12395 & ~n12397;
  assign n12399 = ~po32  & ~n12382;
  assign n12400 = ~n12390 & n12399;
  assign n12401 = ~n12398 & ~n12400;
  assign n12402 = ~n12392 & ~n12401;
  assign n12403 = po33  & ~n12402;
  assign n12404 = ~n11883 & ~n11891;
  assign n12405 = n11889 & n12404;
  assign n12406 = po16  & n12405;
  assign n12407 = po16  & n12404;
  assign n12408 = ~n11889 & ~n12407;
  assign n12409 = ~n12406 & ~n12408;
  assign n12410 = ~po33  & n12402;
  assign n12411 = ~n12409 & ~n12410;
  assign n12412 = ~n12403 & ~n12411;
  assign n12413 = po34  & ~n12412;
  assign n12414 = ~n11894 & ~n11901;
  assign n12415 = n11900 & n12414;
  assign n12416 = po16  & n12415;
  assign n12417 = po16  & n12414;
  assign n12418 = ~n11900 & ~n12417;
  assign n12419 = ~n12416 & ~n12418;
  assign n12420 = ~po34  & ~n12403;
  assign n12421 = ~n12411 & n12420;
  assign n12422 = ~n12419 & ~n12421;
  assign n12423 = ~n12413 & ~n12422;
  assign n12424 = po35  & ~n12423;
  assign n12425 = ~n11904 & ~n11912;
  assign n12426 = n11910 & n12425;
  assign n12427 = po16  & n12426;
  assign n12428 = po16  & n12425;
  assign n12429 = ~n11910 & ~n12428;
  assign n12430 = ~n12427 & ~n12429;
  assign n12431 = ~po35  & n12423;
  assign n12432 = ~n12430 & ~n12431;
  assign n12433 = ~n12424 & ~n12432;
  assign n12434 = po36  & ~n12433;
  assign n12435 = ~n11915 & ~n11922;
  assign n12436 = n11921 & n12435;
  assign n12437 = po16  & n12436;
  assign n12438 = po16  & n12435;
  assign n12439 = ~n11921 & ~n12438;
  assign n12440 = ~n12437 & ~n12439;
  assign n12441 = ~po36  & ~n12424;
  assign n12442 = ~n12432 & n12441;
  assign n12443 = ~n12440 & ~n12442;
  assign n12444 = ~n12434 & ~n12443;
  assign n12445 = po37  & ~n12444;
  assign n12446 = ~n11925 & ~n11933;
  assign n12447 = n11931 & n12446;
  assign n12448 = po16  & n12447;
  assign n12449 = po16  & n12446;
  assign n12450 = ~n11931 & ~n12449;
  assign n12451 = ~n12448 & ~n12450;
  assign n12452 = ~po37  & n12444;
  assign n12453 = ~n12451 & ~n12452;
  assign n12454 = ~n12445 & ~n12453;
  assign n12455 = po38  & ~n12454;
  assign n12456 = ~n11936 & ~n11943;
  assign n12457 = n11942 & n12456;
  assign n12458 = po16  & n12457;
  assign n12459 = po16  & n12456;
  assign n12460 = ~n11942 & ~n12459;
  assign n12461 = ~n12458 & ~n12460;
  assign n12462 = ~po38  & ~n12445;
  assign n12463 = ~n12453 & n12462;
  assign n12464 = ~n12461 & ~n12463;
  assign n12465 = ~n12455 & ~n12464;
  assign n12466 = po39  & ~n12465;
  assign n12467 = ~n11946 & ~n11954;
  assign n12468 = n11952 & n12467;
  assign n12469 = po16  & n12468;
  assign n12470 = po16  & n12467;
  assign n12471 = ~n11952 & ~n12470;
  assign n12472 = ~n12469 & ~n12471;
  assign n12473 = ~po39  & n12465;
  assign n12474 = ~n12472 & ~n12473;
  assign n12475 = ~n12466 & ~n12474;
  assign n12476 = po40  & ~n12475;
  assign n12477 = ~n11957 & ~n11964;
  assign n12478 = n11963 & n12477;
  assign n12479 = po16  & n12478;
  assign n12480 = po16  & n12477;
  assign n12481 = ~n11963 & ~n12480;
  assign n12482 = ~n12479 & ~n12481;
  assign n12483 = ~po40  & ~n12466;
  assign n12484 = ~n12474 & n12483;
  assign n12485 = ~n12482 & ~n12484;
  assign n12486 = ~n12476 & ~n12485;
  assign n12487 = po41  & ~n12486;
  assign n12488 = ~n11967 & ~n11975;
  assign n12489 = n11973 & n12488;
  assign n12490 = po16  & n12489;
  assign n12491 = po16  & n12488;
  assign n12492 = ~n11973 & ~n12491;
  assign n12493 = ~n12490 & ~n12492;
  assign n12494 = ~po41  & n12486;
  assign n12495 = ~n12493 & ~n12494;
  assign n12496 = ~n12487 & ~n12495;
  assign n12497 = po42  & ~n12496;
  assign n12498 = ~n11978 & ~n11985;
  assign n12499 = n11984 & n12498;
  assign n12500 = po16  & n12499;
  assign n12501 = po16  & n12498;
  assign n12502 = ~n11984 & ~n12501;
  assign n12503 = ~n12500 & ~n12502;
  assign n12504 = ~po42  & ~n12487;
  assign n12505 = ~n12495 & n12504;
  assign n12506 = ~n12503 & ~n12505;
  assign n12507 = ~n12497 & ~n12506;
  assign n12508 = po43  & ~n12507;
  assign n12509 = ~n11988 & ~n11996;
  assign n12510 = n11994 & n12509;
  assign n12511 = po16  & n12510;
  assign n12512 = po16  & n12509;
  assign n12513 = ~n11994 & ~n12512;
  assign n12514 = ~n12511 & ~n12513;
  assign n12515 = ~po43  & n12507;
  assign n12516 = ~n12514 & ~n12515;
  assign n12517 = ~n12508 & ~n12516;
  assign n12518 = po44  & ~n12517;
  assign n12519 = ~n11999 & ~n12006;
  assign n12520 = n12005 & n12519;
  assign n12521 = po16  & n12520;
  assign n12522 = po16  & n12519;
  assign n12523 = ~n12005 & ~n12522;
  assign n12524 = ~n12521 & ~n12523;
  assign n12525 = ~po44  & ~n12508;
  assign n12526 = ~n12516 & n12525;
  assign n12527 = ~n12524 & ~n12526;
  assign n12528 = ~n12518 & ~n12527;
  assign n12529 = po45  & ~n12528;
  assign n12530 = ~n12009 & ~n12017;
  assign n12531 = n12015 & n12530;
  assign n12532 = po16  & n12531;
  assign n12533 = po16  & n12530;
  assign n12534 = ~n12015 & ~n12533;
  assign n12535 = ~n12532 & ~n12534;
  assign n12536 = ~po45  & n12528;
  assign n12537 = ~n12535 & ~n12536;
  assign n12538 = ~n12529 & ~n12537;
  assign n12539 = po46  & ~n12538;
  assign n12540 = ~n12020 & ~n12027;
  assign n12541 = n12026 & n12540;
  assign n12542 = po16  & n12541;
  assign n12543 = po16  & n12540;
  assign n12544 = ~n12026 & ~n12543;
  assign n12545 = ~n12542 & ~n12544;
  assign n12546 = ~po46  & ~n12529;
  assign n12547 = ~n12537 & n12546;
  assign n12548 = ~n12545 & ~n12547;
  assign n12549 = ~n12539 & ~n12548;
  assign n12550 = po47  & ~n12549;
  assign n12551 = ~n12030 & ~n12038;
  assign n12552 = n12036 & n12551;
  assign n12553 = po16  & n12552;
  assign n12554 = po16  & n12551;
  assign n12555 = ~n12036 & ~n12554;
  assign n12556 = ~n12553 & ~n12555;
  assign n12557 = ~po47  & n12549;
  assign n12558 = ~n12556 & ~n12557;
  assign n12559 = ~n12550 & ~n12558;
  assign n12560 = po48  & ~n12559;
  assign n12561 = ~n12041 & ~n12048;
  assign n12562 = n12047 & n12561;
  assign n12563 = po16  & n12562;
  assign n12564 = po16  & n12561;
  assign n12565 = ~n12047 & ~n12564;
  assign n12566 = ~n12563 & ~n12565;
  assign n12567 = ~po48  & ~n12550;
  assign n12568 = ~n12558 & n12567;
  assign n12569 = ~n12566 & ~n12568;
  assign n12570 = ~n12560 & ~n12569;
  assign n12571 = po49  & ~n12570;
  assign n12572 = ~n12051 & ~n12053;
  assign n12573 = n12059 & n12572;
  assign n12574 = po16  & n12573;
  assign n12575 = po16  & n12572;
  assign n12576 = ~n12059 & ~n12575;
  assign n12577 = ~n12574 & ~n12576;
  assign n12578 = ~po49  & n12570;
  assign n12579 = ~n12577 & ~n12578;
  assign n12580 = ~n12571 & ~n12579;
  assign n12581 = po50  & ~n12580;
  assign n12582 = ~n12062 & ~n12069;
  assign n12583 = n12068 & n12582;
  assign n12584 = po16  & n12583;
  assign n12585 = po16  & n12582;
  assign n12586 = ~n12068 & ~n12585;
  assign n12587 = ~n12584 & ~n12586;
  assign n12588 = ~po50  & ~n12571;
  assign n12589 = ~n12579 & n12588;
  assign n12590 = ~n12587 & ~n12589;
  assign n12591 = ~n12581 & ~n12590;
  assign n12592 = po51  & ~n12591;
  assign n12593 = ~n12072 & ~n12080;
  assign n12594 = n12078 & n12593;
  assign n12595 = po16  & n12594;
  assign n12596 = po16  & n12593;
  assign n12597 = ~n12078 & ~n12596;
  assign n12598 = ~n12595 & ~n12597;
  assign n12599 = ~po51  & n12591;
  assign n12600 = ~n12598 & ~n12599;
  assign n12601 = ~n12592 & ~n12600;
  assign n12602 = po52  & ~n12601;
  assign n12603 = ~n12083 & ~n12090;
  assign n12604 = n12089 & n12603;
  assign n12605 = po16  & n12604;
  assign n12606 = po16  & n12603;
  assign n12607 = ~n12089 & ~n12606;
  assign n12608 = ~n12605 & ~n12607;
  assign n12609 = ~po52  & ~n12592;
  assign n12610 = ~n12600 & n12609;
  assign n12611 = ~n12608 & ~n12610;
  assign n12612 = ~n12602 & ~n12611;
  assign n12613 = po53  & ~n12612;
  assign n12614 = ~n12093 & ~n12101;
  assign n12615 = n12099 & n12614;
  assign n12616 = po16  & n12615;
  assign n12617 = po16  & n12614;
  assign n12618 = ~n12099 & ~n12617;
  assign n12619 = ~n12616 & ~n12618;
  assign n12620 = ~po53  & n12612;
  assign n12621 = ~n12619 & ~n12620;
  assign n12622 = ~n12613 & ~n12621;
  assign n12623 = po54  & ~n12622;
  assign n12624 = ~n12104 & ~n12111;
  assign n12625 = n12110 & n12624;
  assign n12626 = po16  & n12625;
  assign n12627 = po16  & n12624;
  assign n12628 = ~n12110 & ~n12627;
  assign n12629 = ~n12626 & ~n12628;
  assign n12630 = ~po54  & ~n12613;
  assign n12631 = ~n12621 & n12630;
  assign n12632 = ~n12629 & ~n12631;
  assign n12633 = ~n12623 & ~n12632;
  assign n12634 = po55  & ~n12633;
  assign n12635 = ~n12114 & ~n12122;
  assign n12636 = n12120 & n12635;
  assign n12637 = po16  & n12636;
  assign n12638 = po16  & n12635;
  assign n12639 = ~n12120 & ~n12638;
  assign n12640 = ~n12637 & ~n12639;
  assign n12641 = ~po55  & n12633;
  assign n12642 = ~n12640 & ~n12641;
  assign n12643 = ~n12634 & ~n12642;
  assign n12644 = po56  & ~n12643;
  assign n12645 = ~n12125 & ~n12132;
  assign n12646 = n12131 & n12645;
  assign n12647 = po16  & n12646;
  assign n12648 = po16  & n12645;
  assign n12649 = ~n12131 & ~n12648;
  assign n12650 = ~n12647 & ~n12649;
  assign n12651 = ~po56  & ~n12634;
  assign n12652 = ~n12642 & n12651;
  assign n12653 = ~n12650 & ~n12652;
  assign n12654 = ~n12644 & ~n12653;
  assign n12655 = po57  & ~n12654;
  assign n12656 = ~n12135 & ~n12143;
  assign n12657 = n12141 & n12656;
  assign n12658 = po16  & n12657;
  assign n12659 = po16  & n12656;
  assign n12660 = ~n12141 & ~n12659;
  assign n12661 = ~n12658 & ~n12660;
  assign n12662 = ~po57  & n12654;
  assign n12663 = ~n12661 & ~n12662;
  assign n12664 = ~n12655 & ~n12663;
  assign n12665 = po58  & ~n12664;
  assign n12666 = ~n12146 & ~n12153;
  assign n12667 = n12152 & n12666;
  assign n12668 = po16  & n12667;
  assign n12669 = po16  & n12666;
  assign n12670 = ~n12152 & ~n12669;
  assign n12671 = ~n12668 & ~n12670;
  assign n12672 = ~po58  & ~n12655;
  assign n12673 = ~n12663 & n12672;
  assign n12674 = ~n12671 & ~n12673;
  assign n12675 = ~n12665 & ~n12674;
  assign n12676 = po59  & ~n12675;
  assign n12677 = ~n12156 & ~n12164;
  assign n12678 = n12162 & n12677;
  assign n12679 = po16  & n12678;
  assign n12680 = po16  & n12677;
  assign n12681 = ~n12162 & ~n12680;
  assign n12682 = ~n12679 & ~n12681;
  assign n12683 = ~po59  & n12675;
  assign n12684 = ~n12682 & ~n12683;
  assign n12685 = ~n12676 & ~n12684;
  assign n12686 = po60  & ~n12685;
  assign n12687 = ~n12167 & ~n12174;
  assign n12688 = n12173 & n12687;
  assign n12689 = po16  & n12688;
  assign n12690 = po16  & n12687;
  assign n12691 = ~n12173 & ~n12690;
  assign n12692 = ~n12689 & ~n12691;
  assign n12693 = ~po60  & ~n12676;
  assign n12694 = ~n12684 & n12693;
  assign n12695 = ~n12692 & ~n12694;
  assign n12696 = ~n12686 & ~n12695;
  assign n12697 = po61  & ~n12696;
  assign n12698 = ~n12177 & ~n12185;
  assign n12699 = n12183 & n12698;
  assign n12700 = po16  & n12699;
  assign n12701 = po16  & n12698;
  assign n12702 = ~n12183 & ~n12701;
  assign n12703 = ~n12700 & ~n12702;
  assign n12704 = ~po61  & n12696;
  assign n12705 = ~n12703 & ~n12704;
  assign n12706 = ~n12697 & ~n12705;
  assign n12707 = po62  & ~n12706;
  assign n12708 = ~n12188 & ~n12195;
  assign n12709 = n12194 & n12708;
  assign n12710 = po16  & n12709;
  assign n12711 = po16  & n12708;
  assign n12712 = ~n12194 & ~n12711;
  assign n12713 = ~n12710 & ~n12712;
  assign n12714 = ~po62  & ~n12697;
  assign n12715 = ~n12705 & n12714;
  assign n12716 = ~n12713 & ~n12715;
  assign n12717 = ~n12707 & ~n12716;
  assign n12718 = ~n12198 & ~n12206;
  assign n12719 = po16  & n12718;
  assign n12720 = ~n12204 & ~n12719;
  assign n12721 = n12204 & n12719;
  assign n12722 = ~n12720 & ~n12721;
  assign n12723 = ~n12208 & ~n12213;
  assign n12724 = po16  & n12723;
  assign n12725 = ~n12226 & ~n12724;
  assign n12726 = ~n12722 & n12725;
  assign n12727 = ~n12717 & n12726;
  assign n12728 = ~po63  & ~n12727;
  assign n12729 = ~n12213 & po16 ;
  assign n12730 = n12208 & ~n12729;
  assign n12731 = po63  & ~n12723;
  assign n12732 = ~n12730 & n12731;
  assign n12733 = n12213 & ~po16 ;
  assign n12734 = ~n12732 & ~n12733;
  assign n12735 = n12717 & n12722;
  assign n12736 = n12734 & ~n12735;
  assign po15  = n12728 | ~n12736;
  assign n12738 = pi30  & po15 ;
  assign n12739 = ~pi28  & ~pi29 ;
  assign n12740 = ~pi30  & n12739;
  assign n12741 = ~n12738 & ~n12740;
  assign n12742 = po16  & ~n12741;
  assign n12743 = n12225 & ~n12740;
  assign n12744 = ~n12226 & n12743;
  assign n12745 = ~n12219 & n12744;
  assign n12746 = ~n12738 & n12745;
  assign n12747 = ~pi30  & po15 ;
  assign n12748 = pi31  & ~n12747;
  assign n12749 = n12230 & po15 ;
  assign n12750 = ~n12748 & ~n12749;
  assign n12751 = ~n12746 & n12750;
  assign n12752 = ~n12742 & ~n12751;
  assign n12753 = po17  & ~n12752;
  assign n12754 = po16  & n12734;
  assign n12755 = ~n12735 & n12754;
  assign n12756 = ~n12728 & n12755;
  assign n12757 = ~n12749 & ~n12756;
  assign n12758 = pi32  & ~n12757;
  assign n12759 = ~pi32  & n12757;
  assign n12760 = ~n12758 & ~n12759;
  assign n12761 = ~po17  & n12752;
  assign n12762 = ~n12760 & ~n12761;
  assign n12763 = ~n12753 & ~n12762;
  assign n12764 = po18  & ~n12763;
  assign n12765 = ~n12233 & ~n12237;
  assign n12766 = ~n12241 & n12765;
  assign n12767 = po15  & n12766;
  assign n12768 = po15  & n12765;
  assign n12769 = n12241 & ~n12768;
  assign n12770 = ~n12767 & ~n12769;
  assign n12771 = ~po18  & ~n12753;
  assign n12772 = ~n12762 & n12771;
  assign n12773 = ~n12770 & ~n12772;
  assign n12774 = ~n12764 & ~n12773;
  assign n12775 = po19  & ~n12774;
  assign n12776 = ~n12244 & ~n12246;
  assign n12777 = n12253 & n12776;
  assign n12778 = po15  & n12777;
  assign n12779 = po15  & n12776;
  assign n12780 = ~n12253 & ~n12779;
  assign n12781 = ~n12778 & ~n12780;
  assign n12782 = ~po19  & n12774;
  assign n12783 = ~n12781 & ~n12782;
  assign n12784 = ~n12775 & ~n12783;
  assign n12785 = po20  & ~n12784;
  assign n12786 = ~n12256 & ~n12263;
  assign n12787 = n12262 & n12786;
  assign n12788 = po15  & n12787;
  assign n12789 = po15  & n12786;
  assign n12790 = ~n12262 & ~n12789;
  assign n12791 = ~n12788 & ~n12790;
  assign n12792 = ~po20  & ~n12775;
  assign n12793 = ~n12783 & n12792;
  assign n12794 = ~n12791 & ~n12793;
  assign n12795 = ~n12785 & ~n12794;
  assign n12796 = po21  & ~n12795;
  assign n12797 = ~n12266 & ~n12274;
  assign n12798 = n12272 & n12797;
  assign n12799 = po15  & n12798;
  assign n12800 = po15  & n12797;
  assign n12801 = ~n12272 & ~n12800;
  assign n12802 = ~n12799 & ~n12801;
  assign n12803 = ~po21  & n12795;
  assign n12804 = ~n12802 & ~n12803;
  assign n12805 = ~n12796 & ~n12804;
  assign n12806 = po22  & ~n12805;
  assign n12807 = ~n12277 & ~n12284;
  assign n12808 = n12283 & n12807;
  assign n12809 = po15  & n12808;
  assign n12810 = po15  & n12807;
  assign n12811 = ~n12283 & ~n12810;
  assign n12812 = ~n12809 & ~n12811;
  assign n12813 = ~po22  & ~n12796;
  assign n12814 = ~n12804 & n12813;
  assign n12815 = ~n12812 & ~n12814;
  assign n12816 = ~n12806 & ~n12815;
  assign n12817 = po23  & ~n12816;
  assign n12818 = ~n12287 & ~n12295;
  assign n12819 = n12293 & n12818;
  assign n12820 = po15  & n12819;
  assign n12821 = po15  & n12818;
  assign n12822 = ~n12293 & ~n12821;
  assign n12823 = ~n12820 & ~n12822;
  assign n12824 = ~po23  & n12816;
  assign n12825 = ~n12823 & ~n12824;
  assign n12826 = ~n12817 & ~n12825;
  assign n12827 = po24  & ~n12826;
  assign n12828 = ~n12298 & ~n12305;
  assign n12829 = n12304 & n12828;
  assign n12830 = po15  & n12829;
  assign n12831 = po15  & n12828;
  assign n12832 = ~n12304 & ~n12831;
  assign n12833 = ~n12830 & ~n12832;
  assign n12834 = ~po24  & ~n12817;
  assign n12835 = ~n12825 & n12834;
  assign n12836 = ~n12833 & ~n12835;
  assign n12837 = ~n12827 & ~n12836;
  assign n12838 = po25  & ~n12837;
  assign n12839 = ~n12308 & ~n12316;
  assign n12840 = n12314 & n12839;
  assign n12841 = po15  & n12840;
  assign n12842 = po15  & n12839;
  assign n12843 = ~n12314 & ~n12842;
  assign n12844 = ~n12841 & ~n12843;
  assign n12845 = ~po25  & n12837;
  assign n12846 = ~n12844 & ~n12845;
  assign n12847 = ~n12838 & ~n12846;
  assign n12848 = po26  & ~n12847;
  assign n12849 = ~n12319 & ~n12326;
  assign n12850 = n12325 & n12849;
  assign n12851 = po15  & n12850;
  assign n12852 = po15  & n12849;
  assign n12853 = ~n12325 & ~n12852;
  assign n12854 = ~n12851 & ~n12853;
  assign n12855 = ~po26  & ~n12838;
  assign n12856 = ~n12846 & n12855;
  assign n12857 = ~n12854 & ~n12856;
  assign n12858 = ~n12848 & ~n12857;
  assign n12859 = po27  & ~n12858;
  assign n12860 = ~n12329 & ~n12337;
  assign n12861 = n12335 & n12860;
  assign n12862 = po15  & n12861;
  assign n12863 = po15  & n12860;
  assign n12864 = ~n12335 & ~n12863;
  assign n12865 = ~n12862 & ~n12864;
  assign n12866 = ~po27  & n12858;
  assign n12867 = ~n12865 & ~n12866;
  assign n12868 = ~n12859 & ~n12867;
  assign n12869 = po28  & ~n12868;
  assign n12870 = ~n12340 & ~n12347;
  assign n12871 = n12346 & n12870;
  assign n12872 = po15  & n12871;
  assign n12873 = po15  & n12870;
  assign n12874 = ~n12346 & ~n12873;
  assign n12875 = ~n12872 & ~n12874;
  assign n12876 = ~po28  & ~n12859;
  assign n12877 = ~n12867 & n12876;
  assign n12878 = ~n12875 & ~n12877;
  assign n12879 = ~n12869 & ~n12878;
  assign n12880 = po29  & ~n12879;
  assign n12881 = ~n12350 & ~n12358;
  assign n12882 = n12356 & n12881;
  assign n12883 = po15  & n12882;
  assign n12884 = po15  & n12881;
  assign n12885 = ~n12356 & ~n12884;
  assign n12886 = ~n12883 & ~n12885;
  assign n12887 = ~po29  & n12879;
  assign n12888 = ~n12886 & ~n12887;
  assign n12889 = ~n12880 & ~n12888;
  assign n12890 = po30  & ~n12889;
  assign n12891 = ~n12361 & ~n12368;
  assign n12892 = n12367 & n12891;
  assign n12893 = po15  & n12892;
  assign n12894 = po15  & n12891;
  assign n12895 = ~n12367 & ~n12894;
  assign n12896 = ~n12893 & ~n12895;
  assign n12897 = ~po30  & ~n12880;
  assign n12898 = ~n12888 & n12897;
  assign n12899 = ~n12896 & ~n12898;
  assign n12900 = ~n12890 & ~n12899;
  assign n12901 = po31  & ~n12900;
  assign n12902 = ~n12371 & ~n12379;
  assign n12903 = n12377 & n12902;
  assign n12904 = po15  & n12903;
  assign n12905 = po15  & n12902;
  assign n12906 = ~n12377 & ~n12905;
  assign n12907 = ~n12904 & ~n12906;
  assign n12908 = ~po31  & n12900;
  assign n12909 = ~n12907 & ~n12908;
  assign n12910 = ~n12901 & ~n12909;
  assign n12911 = po32  & ~n12910;
  assign n12912 = ~n12382 & ~n12389;
  assign n12913 = n12388 & n12912;
  assign n12914 = po15  & n12913;
  assign n12915 = po15  & n12912;
  assign n12916 = ~n12388 & ~n12915;
  assign n12917 = ~n12914 & ~n12916;
  assign n12918 = ~po32  & ~n12901;
  assign n12919 = ~n12909 & n12918;
  assign n12920 = ~n12917 & ~n12919;
  assign n12921 = ~n12911 & ~n12920;
  assign n12922 = po33  & ~n12921;
  assign n12923 = ~n12392 & ~n12400;
  assign n12924 = n12398 & n12923;
  assign n12925 = po15  & n12924;
  assign n12926 = po15  & n12923;
  assign n12927 = ~n12398 & ~n12926;
  assign n12928 = ~n12925 & ~n12927;
  assign n12929 = ~po33  & n12921;
  assign n12930 = ~n12928 & ~n12929;
  assign n12931 = ~n12922 & ~n12930;
  assign n12932 = po34  & ~n12931;
  assign n12933 = ~n12403 & ~n12410;
  assign n12934 = n12409 & n12933;
  assign n12935 = po15  & n12934;
  assign n12936 = po15  & n12933;
  assign n12937 = ~n12409 & ~n12936;
  assign n12938 = ~n12935 & ~n12937;
  assign n12939 = ~po34  & ~n12922;
  assign n12940 = ~n12930 & n12939;
  assign n12941 = ~n12938 & ~n12940;
  assign n12942 = ~n12932 & ~n12941;
  assign n12943 = po35  & ~n12942;
  assign n12944 = ~n12413 & ~n12421;
  assign n12945 = n12419 & n12944;
  assign n12946 = po15  & n12945;
  assign n12947 = po15  & n12944;
  assign n12948 = ~n12419 & ~n12947;
  assign n12949 = ~n12946 & ~n12948;
  assign n12950 = ~po35  & n12942;
  assign n12951 = ~n12949 & ~n12950;
  assign n12952 = ~n12943 & ~n12951;
  assign n12953 = po36  & ~n12952;
  assign n12954 = ~n12424 & ~n12431;
  assign n12955 = n12430 & n12954;
  assign n12956 = po15  & n12955;
  assign n12957 = po15  & n12954;
  assign n12958 = ~n12430 & ~n12957;
  assign n12959 = ~n12956 & ~n12958;
  assign n12960 = ~po36  & ~n12943;
  assign n12961 = ~n12951 & n12960;
  assign n12962 = ~n12959 & ~n12961;
  assign n12963 = ~n12953 & ~n12962;
  assign n12964 = po37  & ~n12963;
  assign n12965 = ~n12434 & ~n12442;
  assign n12966 = n12440 & n12965;
  assign n12967 = po15  & n12966;
  assign n12968 = po15  & n12965;
  assign n12969 = ~n12440 & ~n12968;
  assign n12970 = ~n12967 & ~n12969;
  assign n12971 = ~po37  & n12963;
  assign n12972 = ~n12970 & ~n12971;
  assign n12973 = ~n12964 & ~n12972;
  assign n12974 = po38  & ~n12973;
  assign n12975 = ~n12445 & ~n12452;
  assign n12976 = n12451 & n12975;
  assign n12977 = po15  & n12976;
  assign n12978 = po15  & n12975;
  assign n12979 = ~n12451 & ~n12978;
  assign n12980 = ~n12977 & ~n12979;
  assign n12981 = ~po38  & ~n12964;
  assign n12982 = ~n12972 & n12981;
  assign n12983 = ~n12980 & ~n12982;
  assign n12984 = ~n12974 & ~n12983;
  assign n12985 = po39  & ~n12984;
  assign n12986 = ~n12455 & ~n12463;
  assign n12987 = n12461 & n12986;
  assign n12988 = po15  & n12987;
  assign n12989 = po15  & n12986;
  assign n12990 = ~n12461 & ~n12989;
  assign n12991 = ~n12988 & ~n12990;
  assign n12992 = ~po39  & n12984;
  assign n12993 = ~n12991 & ~n12992;
  assign n12994 = ~n12985 & ~n12993;
  assign n12995 = po40  & ~n12994;
  assign n12996 = ~n12466 & ~n12473;
  assign n12997 = n12472 & n12996;
  assign n12998 = po15  & n12997;
  assign n12999 = po15  & n12996;
  assign n13000 = ~n12472 & ~n12999;
  assign n13001 = ~n12998 & ~n13000;
  assign n13002 = ~po40  & ~n12985;
  assign n13003 = ~n12993 & n13002;
  assign n13004 = ~n13001 & ~n13003;
  assign n13005 = ~n12995 & ~n13004;
  assign n13006 = po41  & ~n13005;
  assign n13007 = ~n12476 & ~n12484;
  assign n13008 = n12482 & n13007;
  assign n13009 = po15  & n13008;
  assign n13010 = po15  & n13007;
  assign n13011 = ~n12482 & ~n13010;
  assign n13012 = ~n13009 & ~n13011;
  assign n13013 = ~po41  & n13005;
  assign n13014 = ~n13012 & ~n13013;
  assign n13015 = ~n13006 & ~n13014;
  assign n13016 = po42  & ~n13015;
  assign n13017 = ~n12487 & ~n12494;
  assign n13018 = n12493 & n13017;
  assign n13019 = po15  & n13018;
  assign n13020 = po15  & n13017;
  assign n13021 = ~n12493 & ~n13020;
  assign n13022 = ~n13019 & ~n13021;
  assign n13023 = ~po42  & ~n13006;
  assign n13024 = ~n13014 & n13023;
  assign n13025 = ~n13022 & ~n13024;
  assign n13026 = ~n13016 & ~n13025;
  assign n13027 = po43  & ~n13026;
  assign n13028 = ~n12497 & ~n12505;
  assign n13029 = n12503 & n13028;
  assign n13030 = po15  & n13029;
  assign n13031 = po15  & n13028;
  assign n13032 = ~n12503 & ~n13031;
  assign n13033 = ~n13030 & ~n13032;
  assign n13034 = ~po43  & n13026;
  assign n13035 = ~n13033 & ~n13034;
  assign n13036 = ~n13027 & ~n13035;
  assign n13037 = po44  & ~n13036;
  assign n13038 = ~n12508 & ~n12515;
  assign n13039 = n12514 & n13038;
  assign n13040 = po15  & n13039;
  assign n13041 = po15  & n13038;
  assign n13042 = ~n12514 & ~n13041;
  assign n13043 = ~n13040 & ~n13042;
  assign n13044 = ~po44  & ~n13027;
  assign n13045 = ~n13035 & n13044;
  assign n13046 = ~n13043 & ~n13045;
  assign n13047 = ~n13037 & ~n13046;
  assign n13048 = po45  & ~n13047;
  assign n13049 = ~n12518 & ~n12526;
  assign n13050 = n12524 & n13049;
  assign n13051 = po15  & n13050;
  assign n13052 = po15  & n13049;
  assign n13053 = ~n12524 & ~n13052;
  assign n13054 = ~n13051 & ~n13053;
  assign n13055 = ~po45  & n13047;
  assign n13056 = ~n13054 & ~n13055;
  assign n13057 = ~n13048 & ~n13056;
  assign n13058 = po46  & ~n13057;
  assign n13059 = ~n12529 & ~n12536;
  assign n13060 = n12535 & n13059;
  assign n13061 = po15  & n13060;
  assign n13062 = po15  & n13059;
  assign n13063 = ~n12535 & ~n13062;
  assign n13064 = ~n13061 & ~n13063;
  assign n13065 = ~po46  & ~n13048;
  assign n13066 = ~n13056 & n13065;
  assign n13067 = ~n13064 & ~n13066;
  assign n13068 = ~n13058 & ~n13067;
  assign n13069 = po47  & ~n13068;
  assign n13070 = ~n12539 & ~n12547;
  assign n13071 = n12545 & n13070;
  assign n13072 = po15  & n13071;
  assign n13073 = po15  & n13070;
  assign n13074 = ~n12545 & ~n13073;
  assign n13075 = ~n13072 & ~n13074;
  assign n13076 = ~po47  & n13068;
  assign n13077 = ~n13075 & ~n13076;
  assign n13078 = ~n13069 & ~n13077;
  assign n13079 = po48  & ~n13078;
  assign n13080 = ~n12550 & ~n12557;
  assign n13081 = n12556 & n13080;
  assign n13082 = po15  & n13081;
  assign n13083 = po15  & n13080;
  assign n13084 = ~n12556 & ~n13083;
  assign n13085 = ~n13082 & ~n13084;
  assign n13086 = ~po48  & ~n13069;
  assign n13087 = ~n13077 & n13086;
  assign n13088 = ~n13085 & ~n13087;
  assign n13089 = ~n13079 & ~n13088;
  assign n13090 = po49  & ~n13089;
  assign n13091 = ~n12560 & ~n12568;
  assign n13092 = n12566 & n13091;
  assign n13093 = po15  & n13092;
  assign n13094 = po15  & n13091;
  assign n13095 = ~n12566 & ~n13094;
  assign n13096 = ~n13093 & ~n13095;
  assign n13097 = ~po49  & n13089;
  assign n13098 = ~n13096 & ~n13097;
  assign n13099 = ~n13090 & ~n13098;
  assign n13100 = po50  & ~n13099;
  assign n13101 = ~po50  & ~n13090;
  assign n13102 = ~n13098 & n13101;
  assign n13103 = ~n12571 & ~n12578;
  assign n13104 = n12577 & n13103;
  assign n13105 = po15  & n13104;
  assign n13106 = po15  & n13103;
  assign n13107 = ~n12577 & ~n13106;
  assign n13108 = ~n13105 & ~n13107;
  assign n13109 = ~n13102 & ~n13108;
  assign n13110 = ~n13100 & ~n13109;
  assign n13111 = po51  & ~n13110;
  assign n13112 = ~n12581 & ~n12589;
  assign n13113 = n12587 & n13112;
  assign n13114 = po15  & n13113;
  assign n13115 = po15  & n13112;
  assign n13116 = ~n12587 & ~n13115;
  assign n13117 = ~n13114 & ~n13116;
  assign n13118 = ~po51  & n13110;
  assign n13119 = ~n13117 & ~n13118;
  assign n13120 = ~n13111 & ~n13119;
  assign n13121 = po52  & ~n13120;
  assign n13122 = ~n12592 & ~n12599;
  assign n13123 = n12598 & n13122;
  assign n13124 = po15  & n13123;
  assign n13125 = po15  & n13122;
  assign n13126 = ~n12598 & ~n13125;
  assign n13127 = ~n13124 & ~n13126;
  assign n13128 = ~po52  & ~n13111;
  assign n13129 = ~n13119 & n13128;
  assign n13130 = ~n13127 & ~n13129;
  assign n13131 = ~n13121 & ~n13130;
  assign n13132 = po53  & ~n13131;
  assign n13133 = ~n12602 & ~n12610;
  assign n13134 = n12608 & n13133;
  assign n13135 = po15  & n13134;
  assign n13136 = po15  & n13133;
  assign n13137 = ~n12608 & ~n13136;
  assign n13138 = ~n13135 & ~n13137;
  assign n13139 = ~po53  & n13131;
  assign n13140 = ~n13138 & ~n13139;
  assign n13141 = ~n13132 & ~n13140;
  assign n13142 = po54  & ~n13141;
  assign n13143 = ~n12613 & ~n12620;
  assign n13144 = n12619 & n13143;
  assign n13145 = po15  & n13144;
  assign n13146 = po15  & n13143;
  assign n13147 = ~n12619 & ~n13146;
  assign n13148 = ~n13145 & ~n13147;
  assign n13149 = ~po54  & ~n13132;
  assign n13150 = ~n13140 & n13149;
  assign n13151 = ~n13148 & ~n13150;
  assign n13152 = ~n13142 & ~n13151;
  assign n13153 = po55  & ~n13152;
  assign n13154 = ~n12623 & ~n12631;
  assign n13155 = n12629 & n13154;
  assign n13156 = po15  & n13155;
  assign n13157 = po15  & n13154;
  assign n13158 = ~n12629 & ~n13157;
  assign n13159 = ~n13156 & ~n13158;
  assign n13160 = ~po55  & n13152;
  assign n13161 = ~n13159 & ~n13160;
  assign n13162 = ~n13153 & ~n13161;
  assign n13163 = po56  & ~n13162;
  assign n13164 = ~n12634 & ~n12641;
  assign n13165 = n12640 & n13164;
  assign n13166 = po15  & n13165;
  assign n13167 = po15  & n13164;
  assign n13168 = ~n12640 & ~n13167;
  assign n13169 = ~n13166 & ~n13168;
  assign n13170 = ~po56  & ~n13153;
  assign n13171 = ~n13161 & n13170;
  assign n13172 = ~n13169 & ~n13171;
  assign n13173 = ~n13163 & ~n13172;
  assign n13174 = po57  & ~n13173;
  assign n13175 = ~n12644 & ~n12652;
  assign n13176 = n12650 & n13175;
  assign n13177 = po15  & n13176;
  assign n13178 = po15  & n13175;
  assign n13179 = ~n12650 & ~n13178;
  assign n13180 = ~n13177 & ~n13179;
  assign n13181 = ~po57  & n13173;
  assign n13182 = ~n13180 & ~n13181;
  assign n13183 = ~n13174 & ~n13182;
  assign n13184 = po58  & ~n13183;
  assign n13185 = ~n12655 & ~n12662;
  assign n13186 = n12661 & n13185;
  assign n13187 = po15  & n13186;
  assign n13188 = po15  & n13185;
  assign n13189 = ~n12661 & ~n13188;
  assign n13190 = ~n13187 & ~n13189;
  assign n13191 = ~po58  & ~n13174;
  assign n13192 = ~n13182 & n13191;
  assign n13193 = ~n13190 & ~n13192;
  assign n13194 = ~n13184 & ~n13193;
  assign n13195 = po59  & ~n13194;
  assign n13196 = ~n12665 & ~n12673;
  assign n13197 = n12671 & n13196;
  assign n13198 = po15  & n13197;
  assign n13199 = po15  & n13196;
  assign n13200 = ~n12671 & ~n13199;
  assign n13201 = ~n13198 & ~n13200;
  assign n13202 = ~po59  & n13194;
  assign n13203 = ~n13201 & ~n13202;
  assign n13204 = ~n13195 & ~n13203;
  assign n13205 = po60  & ~n13204;
  assign n13206 = ~n12676 & ~n12683;
  assign n13207 = n12682 & n13206;
  assign n13208 = po15  & n13207;
  assign n13209 = po15  & n13206;
  assign n13210 = ~n12682 & ~n13209;
  assign n13211 = ~n13208 & ~n13210;
  assign n13212 = ~po60  & ~n13195;
  assign n13213 = ~n13203 & n13212;
  assign n13214 = ~n13211 & ~n13213;
  assign n13215 = ~n13205 & ~n13214;
  assign n13216 = po61  & ~n13215;
  assign n13217 = ~n12686 & ~n12694;
  assign n13218 = n12692 & n13217;
  assign n13219 = po15  & n13218;
  assign n13220 = po15  & n13217;
  assign n13221 = ~n12692 & ~n13220;
  assign n13222 = ~n13219 & ~n13221;
  assign n13223 = ~po61  & n13215;
  assign n13224 = ~n13222 & ~n13223;
  assign n13225 = ~n13216 & ~n13224;
  assign n13226 = po62  & ~n13225;
  assign n13227 = ~n12697 & ~n12704;
  assign n13228 = n12703 & n13227;
  assign n13229 = po15  & n13228;
  assign n13230 = po15  & n13227;
  assign n13231 = ~n12703 & ~n13230;
  assign n13232 = ~n13229 & ~n13231;
  assign n13233 = ~po62  & ~n13216;
  assign n13234 = ~n13224 & n13233;
  assign n13235 = ~n13232 & ~n13234;
  assign n13236 = ~n13226 & ~n13235;
  assign n13237 = ~n12707 & ~n12715;
  assign n13238 = po15  & n13237;
  assign n13239 = ~n12713 & ~n13238;
  assign n13240 = n12713 & n13238;
  assign n13241 = ~n13239 & ~n13240;
  assign n13242 = ~n12717 & ~n12722;
  assign n13243 = po15  & n13242;
  assign n13244 = ~n12735 & ~n13243;
  assign n13245 = ~n13241 & n13244;
  assign n13246 = ~n13236 & n13245;
  assign n13247 = ~po63  & ~n13246;
  assign n13248 = ~n12722 & po15 ;
  assign n13249 = n12717 & ~n13248;
  assign n13250 = po63  & ~n13242;
  assign n13251 = ~n13249 & n13250;
  assign n13252 = n12722 & ~po15 ;
  assign n13253 = ~n13251 & ~n13252;
  assign n13254 = n13236 & n13241;
  assign n13255 = n13253 & ~n13254;
  assign po14  = n13247 | ~n13255;
  assign n13257 = pi28  & po14 ;
  assign n13258 = ~pi26  & ~pi27 ;
  assign n13259 = ~pi28  & n13258;
  assign n13260 = ~n13257 & ~n13259;
  assign n13261 = po15  & ~n13260;
  assign n13262 = n12734 & ~n13259;
  assign n13263 = ~n12735 & n13262;
  assign n13264 = ~n12728 & n13263;
  assign n13265 = ~n13257 & n13264;
  assign n13266 = ~pi28  & po14 ;
  assign n13267 = pi29  & ~n13266;
  assign n13268 = n12739 & po14 ;
  assign n13269 = ~n13267 & ~n13268;
  assign n13270 = ~n13265 & n13269;
  assign n13271 = ~n13261 & ~n13270;
  assign n13272 = po16  & ~n13271;
  assign n13273 = ~po16  & ~n13261;
  assign n13274 = ~n13270 & n13273;
  assign n13275 = po15  & n13253;
  assign n13276 = ~n13254 & n13275;
  assign n13277 = ~n13247 & n13276;
  assign n13278 = ~n13268 & ~n13277;
  assign n13279 = pi30  & ~n13278;
  assign n13280 = ~pi30  & n13278;
  assign n13281 = ~n13279 & ~n13280;
  assign n13282 = ~n13274 & ~n13281;
  assign n13283 = ~n13272 & ~n13282;
  assign n13284 = po17  & ~n13283;
  assign n13285 = ~n12742 & ~n12746;
  assign n13286 = ~n12750 & n13285;
  assign n13287 = po14  & n13286;
  assign n13288 = po14  & n13285;
  assign n13289 = n12750 & ~n13288;
  assign n13290 = ~n13287 & ~n13289;
  assign n13291 = ~po17  & n13283;
  assign n13292 = ~n13290 & ~n13291;
  assign n13293 = ~n13284 & ~n13292;
  assign n13294 = po18  & ~n13293;
  assign n13295 = ~n12753 & ~n12761;
  assign n13296 = n12760 & n13295;
  assign n13297 = po14  & n13296;
  assign n13298 = po14  & n13295;
  assign n13299 = ~n12760 & ~n13298;
  assign n13300 = ~n13297 & ~n13299;
  assign n13301 = ~po18  & ~n13284;
  assign n13302 = ~n13292 & n13301;
  assign n13303 = ~n13300 & ~n13302;
  assign n13304 = ~n13294 & ~n13303;
  assign n13305 = po19  & ~n13304;
  assign n13306 = ~n12764 & ~n12772;
  assign n13307 = n12770 & n13306;
  assign n13308 = po14  & n13307;
  assign n13309 = po14  & n13306;
  assign n13310 = ~n12770 & ~n13309;
  assign n13311 = ~n13308 & ~n13310;
  assign n13312 = ~po19  & n13304;
  assign n13313 = ~n13311 & ~n13312;
  assign n13314 = ~n13305 & ~n13313;
  assign n13315 = po20  & ~n13314;
  assign n13316 = ~n12775 & ~n12782;
  assign n13317 = n12781 & n13316;
  assign n13318 = po14  & n13317;
  assign n13319 = po14  & n13316;
  assign n13320 = ~n12781 & ~n13319;
  assign n13321 = ~n13318 & ~n13320;
  assign n13322 = ~po20  & ~n13305;
  assign n13323 = ~n13313 & n13322;
  assign n13324 = ~n13321 & ~n13323;
  assign n13325 = ~n13315 & ~n13324;
  assign n13326 = po21  & ~n13325;
  assign n13327 = ~n12785 & ~n12793;
  assign n13328 = n12791 & n13327;
  assign n13329 = po14  & n13328;
  assign n13330 = po14  & n13327;
  assign n13331 = ~n12791 & ~n13330;
  assign n13332 = ~n13329 & ~n13331;
  assign n13333 = ~po21  & n13325;
  assign n13334 = ~n13332 & ~n13333;
  assign n13335 = ~n13326 & ~n13334;
  assign n13336 = po22  & ~n13335;
  assign n13337 = ~n12796 & ~n12803;
  assign n13338 = n12802 & n13337;
  assign n13339 = po14  & n13338;
  assign n13340 = po14  & n13337;
  assign n13341 = ~n12802 & ~n13340;
  assign n13342 = ~n13339 & ~n13341;
  assign n13343 = ~po22  & ~n13326;
  assign n13344 = ~n13334 & n13343;
  assign n13345 = ~n13342 & ~n13344;
  assign n13346 = ~n13336 & ~n13345;
  assign n13347 = po23  & ~n13346;
  assign n13348 = ~n12806 & ~n12814;
  assign n13349 = n12812 & n13348;
  assign n13350 = po14  & n13349;
  assign n13351 = po14  & n13348;
  assign n13352 = ~n12812 & ~n13351;
  assign n13353 = ~n13350 & ~n13352;
  assign n13354 = ~po23  & n13346;
  assign n13355 = ~n13353 & ~n13354;
  assign n13356 = ~n13347 & ~n13355;
  assign n13357 = po24  & ~n13356;
  assign n13358 = ~n12817 & ~n12824;
  assign n13359 = n12823 & n13358;
  assign n13360 = po14  & n13359;
  assign n13361 = po14  & n13358;
  assign n13362 = ~n12823 & ~n13361;
  assign n13363 = ~n13360 & ~n13362;
  assign n13364 = ~po24  & ~n13347;
  assign n13365 = ~n13355 & n13364;
  assign n13366 = ~n13363 & ~n13365;
  assign n13367 = ~n13357 & ~n13366;
  assign n13368 = po25  & ~n13367;
  assign n13369 = ~n12827 & ~n12835;
  assign n13370 = n12833 & n13369;
  assign n13371 = po14  & n13370;
  assign n13372 = po14  & n13369;
  assign n13373 = ~n12833 & ~n13372;
  assign n13374 = ~n13371 & ~n13373;
  assign n13375 = ~po25  & n13367;
  assign n13376 = ~n13374 & ~n13375;
  assign n13377 = ~n13368 & ~n13376;
  assign n13378 = po26  & ~n13377;
  assign n13379 = ~n12838 & ~n12845;
  assign n13380 = n12844 & n13379;
  assign n13381 = po14  & n13380;
  assign n13382 = po14  & n13379;
  assign n13383 = ~n12844 & ~n13382;
  assign n13384 = ~n13381 & ~n13383;
  assign n13385 = ~po26  & ~n13368;
  assign n13386 = ~n13376 & n13385;
  assign n13387 = ~n13384 & ~n13386;
  assign n13388 = ~n13378 & ~n13387;
  assign n13389 = po27  & ~n13388;
  assign n13390 = ~n12848 & ~n12856;
  assign n13391 = n12854 & n13390;
  assign n13392 = po14  & n13391;
  assign n13393 = po14  & n13390;
  assign n13394 = ~n12854 & ~n13393;
  assign n13395 = ~n13392 & ~n13394;
  assign n13396 = ~po27  & n13388;
  assign n13397 = ~n13395 & ~n13396;
  assign n13398 = ~n13389 & ~n13397;
  assign n13399 = po28  & ~n13398;
  assign n13400 = ~n12859 & ~n12866;
  assign n13401 = n12865 & n13400;
  assign n13402 = po14  & n13401;
  assign n13403 = po14  & n13400;
  assign n13404 = ~n12865 & ~n13403;
  assign n13405 = ~n13402 & ~n13404;
  assign n13406 = ~po28  & ~n13389;
  assign n13407 = ~n13397 & n13406;
  assign n13408 = ~n13405 & ~n13407;
  assign n13409 = ~n13399 & ~n13408;
  assign n13410 = po29  & ~n13409;
  assign n13411 = ~n12869 & ~n12877;
  assign n13412 = n12875 & n13411;
  assign n13413 = po14  & n13412;
  assign n13414 = po14  & n13411;
  assign n13415 = ~n12875 & ~n13414;
  assign n13416 = ~n13413 & ~n13415;
  assign n13417 = ~po29  & n13409;
  assign n13418 = ~n13416 & ~n13417;
  assign n13419 = ~n13410 & ~n13418;
  assign n13420 = po30  & ~n13419;
  assign n13421 = ~n12880 & ~n12887;
  assign n13422 = n12886 & n13421;
  assign n13423 = po14  & n13422;
  assign n13424 = po14  & n13421;
  assign n13425 = ~n12886 & ~n13424;
  assign n13426 = ~n13423 & ~n13425;
  assign n13427 = ~po30  & ~n13410;
  assign n13428 = ~n13418 & n13427;
  assign n13429 = ~n13426 & ~n13428;
  assign n13430 = ~n13420 & ~n13429;
  assign n13431 = po31  & ~n13430;
  assign n13432 = ~n12890 & ~n12898;
  assign n13433 = n12896 & n13432;
  assign n13434 = po14  & n13433;
  assign n13435 = po14  & n13432;
  assign n13436 = ~n12896 & ~n13435;
  assign n13437 = ~n13434 & ~n13436;
  assign n13438 = ~po31  & n13430;
  assign n13439 = ~n13437 & ~n13438;
  assign n13440 = ~n13431 & ~n13439;
  assign n13441 = po32  & ~n13440;
  assign n13442 = ~n12901 & ~n12908;
  assign n13443 = n12907 & n13442;
  assign n13444 = po14  & n13443;
  assign n13445 = po14  & n13442;
  assign n13446 = ~n12907 & ~n13445;
  assign n13447 = ~n13444 & ~n13446;
  assign n13448 = ~po32  & ~n13431;
  assign n13449 = ~n13439 & n13448;
  assign n13450 = ~n13447 & ~n13449;
  assign n13451 = ~n13441 & ~n13450;
  assign n13452 = po33  & ~n13451;
  assign n13453 = ~n12911 & ~n12919;
  assign n13454 = n12917 & n13453;
  assign n13455 = po14  & n13454;
  assign n13456 = po14  & n13453;
  assign n13457 = ~n12917 & ~n13456;
  assign n13458 = ~n13455 & ~n13457;
  assign n13459 = ~po33  & n13451;
  assign n13460 = ~n13458 & ~n13459;
  assign n13461 = ~n13452 & ~n13460;
  assign n13462 = po34  & ~n13461;
  assign n13463 = ~n12922 & ~n12929;
  assign n13464 = n12928 & n13463;
  assign n13465 = po14  & n13464;
  assign n13466 = po14  & n13463;
  assign n13467 = ~n12928 & ~n13466;
  assign n13468 = ~n13465 & ~n13467;
  assign n13469 = ~po34  & ~n13452;
  assign n13470 = ~n13460 & n13469;
  assign n13471 = ~n13468 & ~n13470;
  assign n13472 = ~n13462 & ~n13471;
  assign n13473 = po35  & ~n13472;
  assign n13474 = ~n12932 & ~n12940;
  assign n13475 = n12938 & n13474;
  assign n13476 = po14  & n13475;
  assign n13477 = po14  & n13474;
  assign n13478 = ~n12938 & ~n13477;
  assign n13479 = ~n13476 & ~n13478;
  assign n13480 = ~po35  & n13472;
  assign n13481 = ~n13479 & ~n13480;
  assign n13482 = ~n13473 & ~n13481;
  assign n13483 = po36  & ~n13482;
  assign n13484 = ~n12943 & ~n12950;
  assign n13485 = n12949 & n13484;
  assign n13486 = po14  & n13485;
  assign n13487 = po14  & n13484;
  assign n13488 = ~n12949 & ~n13487;
  assign n13489 = ~n13486 & ~n13488;
  assign n13490 = ~po36  & ~n13473;
  assign n13491 = ~n13481 & n13490;
  assign n13492 = ~n13489 & ~n13491;
  assign n13493 = ~n13483 & ~n13492;
  assign n13494 = po37  & ~n13493;
  assign n13495 = ~n12953 & ~n12961;
  assign n13496 = n12959 & n13495;
  assign n13497 = po14  & n13496;
  assign n13498 = po14  & n13495;
  assign n13499 = ~n12959 & ~n13498;
  assign n13500 = ~n13497 & ~n13499;
  assign n13501 = ~po37  & n13493;
  assign n13502 = ~n13500 & ~n13501;
  assign n13503 = ~n13494 & ~n13502;
  assign n13504 = po38  & ~n13503;
  assign n13505 = ~n12964 & ~n12971;
  assign n13506 = n12970 & n13505;
  assign n13507 = po14  & n13506;
  assign n13508 = po14  & n13505;
  assign n13509 = ~n12970 & ~n13508;
  assign n13510 = ~n13507 & ~n13509;
  assign n13511 = ~po38  & ~n13494;
  assign n13512 = ~n13502 & n13511;
  assign n13513 = ~n13510 & ~n13512;
  assign n13514 = ~n13504 & ~n13513;
  assign n13515 = po39  & ~n13514;
  assign n13516 = ~n12974 & ~n12982;
  assign n13517 = n12980 & n13516;
  assign n13518 = po14  & n13517;
  assign n13519 = po14  & n13516;
  assign n13520 = ~n12980 & ~n13519;
  assign n13521 = ~n13518 & ~n13520;
  assign n13522 = ~po39  & n13514;
  assign n13523 = ~n13521 & ~n13522;
  assign n13524 = ~n13515 & ~n13523;
  assign n13525 = po40  & ~n13524;
  assign n13526 = ~n12985 & ~n12992;
  assign n13527 = n12991 & n13526;
  assign n13528 = po14  & n13527;
  assign n13529 = po14  & n13526;
  assign n13530 = ~n12991 & ~n13529;
  assign n13531 = ~n13528 & ~n13530;
  assign n13532 = ~po40  & ~n13515;
  assign n13533 = ~n13523 & n13532;
  assign n13534 = ~n13531 & ~n13533;
  assign n13535 = ~n13525 & ~n13534;
  assign n13536 = po41  & ~n13535;
  assign n13537 = ~n12995 & ~n13003;
  assign n13538 = n13001 & n13537;
  assign n13539 = po14  & n13538;
  assign n13540 = po14  & n13537;
  assign n13541 = ~n13001 & ~n13540;
  assign n13542 = ~n13539 & ~n13541;
  assign n13543 = ~po41  & n13535;
  assign n13544 = ~n13542 & ~n13543;
  assign n13545 = ~n13536 & ~n13544;
  assign n13546 = po42  & ~n13545;
  assign n13547 = ~n13006 & ~n13013;
  assign n13548 = n13012 & n13547;
  assign n13549 = po14  & n13548;
  assign n13550 = po14  & n13547;
  assign n13551 = ~n13012 & ~n13550;
  assign n13552 = ~n13549 & ~n13551;
  assign n13553 = ~po42  & ~n13536;
  assign n13554 = ~n13544 & n13553;
  assign n13555 = ~n13552 & ~n13554;
  assign n13556 = ~n13546 & ~n13555;
  assign n13557 = po43  & ~n13556;
  assign n13558 = ~n13016 & ~n13024;
  assign n13559 = n13022 & n13558;
  assign n13560 = po14  & n13559;
  assign n13561 = po14  & n13558;
  assign n13562 = ~n13022 & ~n13561;
  assign n13563 = ~n13560 & ~n13562;
  assign n13564 = ~po43  & n13556;
  assign n13565 = ~n13563 & ~n13564;
  assign n13566 = ~n13557 & ~n13565;
  assign n13567 = po44  & ~n13566;
  assign n13568 = ~n13027 & ~n13034;
  assign n13569 = n13033 & n13568;
  assign n13570 = po14  & n13569;
  assign n13571 = po14  & n13568;
  assign n13572 = ~n13033 & ~n13571;
  assign n13573 = ~n13570 & ~n13572;
  assign n13574 = ~po44  & ~n13557;
  assign n13575 = ~n13565 & n13574;
  assign n13576 = ~n13573 & ~n13575;
  assign n13577 = ~n13567 & ~n13576;
  assign n13578 = po45  & ~n13577;
  assign n13579 = ~n13037 & ~n13045;
  assign n13580 = n13043 & n13579;
  assign n13581 = po14  & n13580;
  assign n13582 = po14  & n13579;
  assign n13583 = ~n13043 & ~n13582;
  assign n13584 = ~n13581 & ~n13583;
  assign n13585 = ~po45  & n13577;
  assign n13586 = ~n13584 & ~n13585;
  assign n13587 = ~n13578 & ~n13586;
  assign n13588 = po46  & ~n13587;
  assign n13589 = ~n13048 & ~n13055;
  assign n13590 = n13054 & n13589;
  assign n13591 = po14  & n13590;
  assign n13592 = po14  & n13589;
  assign n13593 = ~n13054 & ~n13592;
  assign n13594 = ~n13591 & ~n13593;
  assign n13595 = ~po46  & ~n13578;
  assign n13596 = ~n13586 & n13595;
  assign n13597 = ~n13594 & ~n13596;
  assign n13598 = ~n13588 & ~n13597;
  assign n13599 = po47  & ~n13598;
  assign n13600 = ~n13058 & ~n13066;
  assign n13601 = n13064 & n13600;
  assign n13602 = po14  & n13601;
  assign n13603 = po14  & n13600;
  assign n13604 = ~n13064 & ~n13603;
  assign n13605 = ~n13602 & ~n13604;
  assign n13606 = ~po47  & n13598;
  assign n13607 = ~n13605 & ~n13606;
  assign n13608 = ~n13599 & ~n13607;
  assign n13609 = po48  & ~n13608;
  assign n13610 = ~n13069 & ~n13076;
  assign n13611 = n13075 & n13610;
  assign n13612 = po14  & n13611;
  assign n13613 = po14  & n13610;
  assign n13614 = ~n13075 & ~n13613;
  assign n13615 = ~n13612 & ~n13614;
  assign n13616 = ~po48  & ~n13599;
  assign n13617 = ~n13607 & n13616;
  assign n13618 = ~n13615 & ~n13617;
  assign n13619 = ~n13609 & ~n13618;
  assign n13620 = po49  & ~n13619;
  assign n13621 = ~n13079 & ~n13087;
  assign n13622 = n13085 & n13621;
  assign n13623 = po14  & n13622;
  assign n13624 = po14  & n13621;
  assign n13625 = ~n13085 & ~n13624;
  assign n13626 = ~n13623 & ~n13625;
  assign n13627 = ~po49  & n13619;
  assign n13628 = ~n13626 & ~n13627;
  assign n13629 = ~n13620 & ~n13628;
  assign n13630 = po50  & ~n13629;
  assign n13631 = ~n13090 & ~n13097;
  assign n13632 = n13096 & n13631;
  assign n13633 = po14  & n13632;
  assign n13634 = po14  & n13631;
  assign n13635 = ~n13096 & ~n13634;
  assign n13636 = ~n13633 & ~n13635;
  assign n13637 = ~po50  & ~n13620;
  assign n13638 = ~n13628 & n13637;
  assign n13639 = ~n13636 & ~n13638;
  assign n13640 = ~n13630 & ~n13639;
  assign n13641 = po51  & ~n13640;
  assign n13642 = ~n13100 & ~n13102;
  assign n13643 = n13108 & n13642;
  assign n13644 = po14  & n13643;
  assign n13645 = po14  & n13642;
  assign n13646 = ~n13108 & ~n13645;
  assign n13647 = ~n13644 & ~n13646;
  assign n13648 = ~po51  & n13640;
  assign n13649 = ~n13647 & ~n13648;
  assign n13650 = ~n13641 & ~n13649;
  assign n13651 = po52  & ~n13650;
  assign n13652 = ~n13111 & ~n13118;
  assign n13653 = n13117 & n13652;
  assign n13654 = po14  & n13653;
  assign n13655 = po14  & n13652;
  assign n13656 = ~n13117 & ~n13655;
  assign n13657 = ~n13654 & ~n13656;
  assign n13658 = ~po52  & ~n13641;
  assign n13659 = ~n13649 & n13658;
  assign n13660 = ~n13657 & ~n13659;
  assign n13661 = ~n13651 & ~n13660;
  assign n13662 = po53  & ~n13661;
  assign n13663 = ~n13121 & ~n13129;
  assign n13664 = n13127 & n13663;
  assign n13665 = po14  & n13664;
  assign n13666 = po14  & n13663;
  assign n13667 = ~n13127 & ~n13666;
  assign n13668 = ~n13665 & ~n13667;
  assign n13669 = ~po53  & n13661;
  assign n13670 = ~n13668 & ~n13669;
  assign n13671 = ~n13662 & ~n13670;
  assign n13672 = po54  & ~n13671;
  assign n13673 = ~n13132 & ~n13139;
  assign n13674 = n13138 & n13673;
  assign n13675 = po14  & n13674;
  assign n13676 = po14  & n13673;
  assign n13677 = ~n13138 & ~n13676;
  assign n13678 = ~n13675 & ~n13677;
  assign n13679 = ~po54  & ~n13662;
  assign n13680 = ~n13670 & n13679;
  assign n13681 = ~n13678 & ~n13680;
  assign n13682 = ~n13672 & ~n13681;
  assign n13683 = po55  & ~n13682;
  assign n13684 = ~n13142 & ~n13150;
  assign n13685 = n13148 & n13684;
  assign n13686 = po14  & n13685;
  assign n13687 = po14  & n13684;
  assign n13688 = ~n13148 & ~n13687;
  assign n13689 = ~n13686 & ~n13688;
  assign n13690 = ~po55  & n13682;
  assign n13691 = ~n13689 & ~n13690;
  assign n13692 = ~n13683 & ~n13691;
  assign n13693 = po56  & ~n13692;
  assign n13694 = ~n13153 & ~n13160;
  assign n13695 = n13159 & n13694;
  assign n13696 = po14  & n13695;
  assign n13697 = po14  & n13694;
  assign n13698 = ~n13159 & ~n13697;
  assign n13699 = ~n13696 & ~n13698;
  assign n13700 = ~po56  & ~n13683;
  assign n13701 = ~n13691 & n13700;
  assign n13702 = ~n13699 & ~n13701;
  assign n13703 = ~n13693 & ~n13702;
  assign n13704 = po57  & ~n13703;
  assign n13705 = ~n13163 & ~n13171;
  assign n13706 = n13169 & n13705;
  assign n13707 = po14  & n13706;
  assign n13708 = po14  & n13705;
  assign n13709 = ~n13169 & ~n13708;
  assign n13710 = ~n13707 & ~n13709;
  assign n13711 = ~po57  & n13703;
  assign n13712 = ~n13710 & ~n13711;
  assign n13713 = ~n13704 & ~n13712;
  assign n13714 = po58  & ~n13713;
  assign n13715 = ~n13174 & ~n13181;
  assign n13716 = n13180 & n13715;
  assign n13717 = po14  & n13716;
  assign n13718 = po14  & n13715;
  assign n13719 = ~n13180 & ~n13718;
  assign n13720 = ~n13717 & ~n13719;
  assign n13721 = ~po58  & ~n13704;
  assign n13722 = ~n13712 & n13721;
  assign n13723 = ~n13720 & ~n13722;
  assign n13724 = ~n13714 & ~n13723;
  assign n13725 = po59  & ~n13724;
  assign n13726 = ~n13184 & ~n13192;
  assign n13727 = n13190 & n13726;
  assign n13728 = po14  & n13727;
  assign n13729 = po14  & n13726;
  assign n13730 = ~n13190 & ~n13729;
  assign n13731 = ~n13728 & ~n13730;
  assign n13732 = ~po59  & n13724;
  assign n13733 = ~n13731 & ~n13732;
  assign n13734 = ~n13725 & ~n13733;
  assign n13735 = po60  & ~n13734;
  assign n13736 = ~n13195 & ~n13202;
  assign n13737 = n13201 & n13736;
  assign n13738 = po14  & n13737;
  assign n13739 = po14  & n13736;
  assign n13740 = ~n13201 & ~n13739;
  assign n13741 = ~n13738 & ~n13740;
  assign n13742 = ~po60  & ~n13725;
  assign n13743 = ~n13733 & n13742;
  assign n13744 = ~n13741 & ~n13743;
  assign n13745 = ~n13735 & ~n13744;
  assign n13746 = po61  & ~n13745;
  assign n13747 = ~n13205 & ~n13213;
  assign n13748 = n13211 & n13747;
  assign n13749 = po14  & n13748;
  assign n13750 = po14  & n13747;
  assign n13751 = ~n13211 & ~n13750;
  assign n13752 = ~n13749 & ~n13751;
  assign n13753 = ~po61  & n13745;
  assign n13754 = ~n13752 & ~n13753;
  assign n13755 = ~n13746 & ~n13754;
  assign n13756 = po62  & ~n13755;
  assign n13757 = ~n13216 & ~n13223;
  assign n13758 = n13222 & n13757;
  assign n13759 = po14  & n13758;
  assign n13760 = po14  & n13757;
  assign n13761 = ~n13222 & ~n13760;
  assign n13762 = ~n13759 & ~n13761;
  assign n13763 = ~po62  & ~n13746;
  assign n13764 = ~n13754 & n13763;
  assign n13765 = ~n13762 & ~n13764;
  assign n13766 = ~n13756 & ~n13765;
  assign n13767 = ~n13226 & ~n13234;
  assign n13768 = po14  & n13767;
  assign n13769 = ~n13232 & ~n13768;
  assign n13770 = n13232 & n13768;
  assign n13771 = ~n13769 & ~n13770;
  assign n13772 = ~n13236 & ~n13241;
  assign n13773 = po14  & n13772;
  assign n13774 = ~n13254 & ~n13773;
  assign n13775 = ~n13771 & n13774;
  assign n13776 = ~n13766 & n13775;
  assign n13777 = ~po63  & ~n13776;
  assign n13778 = ~n13241 & po14 ;
  assign n13779 = n13236 & ~n13778;
  assign n13780 = po63  & ~n13772;
  assign n13781 = ~n13779 & n13780;
  assign n13782 = n13241 & ~po14 ;
  assign n13783 = ~n13781 & ~n13782;
  assign n13784 = n13766 & n13771;
  assign n13785 = n13783 & ~n13784;
  assign po13  = n13777 | ~n13785;
  assign n13787 = pi26  & po13 ;
  assign n13788 = ~pi24  & ~pi25 ;
  assign n13789 = ~pi26  & n13788;
  assign n13790 = ~n13787 & ~n13789;
  assign n13791 = po14  & ~n13790;
  assign n13792 = n13253 & ~n13789;
  assign n13793 = ~n13254 & n13792;
  assign n13794 = ~n13247 & n13793;
  assign n13795 = ~n13787 & n13794;
  assign n13796 = ~pi26  & po13 ;
  assign n13797 = pi27  & ~n13796;
  assign n13798 = n13258 & po13 ;
  assign n13799 = ~n13797 & ~n13798;
  assign n13800 = ~n13795 & n13799;
  assign n13801 = ~n13791 & ~n13800;
  assign n13802 = po15  & ~n13801;
  assign n13803 = po14  & n13783;
  assign n13804 = ~n13784 & n13803;
  assign n13805 = ~n13777 & n13804;
  assign n13806 = ~n13798 & ~n13805;
  assign n13807 = pi28  & ~n13806;
  assign n13808 = ~pi28  & n13806;
  assign n13809 = ~n13807 & ~n13808;
  assign n13810 = ~po15  & n13801;
  assign n13811 = ~n13809 & ~n13810;
  assign n13812 = ~n13802 & ~n13811;
  assign n13813 = po16  & ~n13812;
  assign n13814 = ~n13261 & ~n13265;
  assign n13815 = ~n13269 & n13814;
  assign n13816 = po13  & n13815;
  assign n13817 = po13  & n13814;
  assign n13818 = n13269 & ~n13817;
  assign n13819 = ~n13816 & ~n13818;
  assign n13820 = ~po16  & ~n13802;
  assign n13821 = ~n13811 & n13820;
  assign n13822 = ~n13819 & ~n13821;
  assign n13823 = ~n13813 & ~n13822;
  assign n13824 = po17  & ~n13823;
  assign n13825 = ~n13272 & ~n13274;
  assign n13826 = n13281 & n13825;
  assign n13827 = po13  & n13826;
  assign n13828 = po13  & n13825;
  assign n13829 = ~n13281 & ~n13828;
  assign n13830 = ~n13827 & ~n13829;
  assign n13831 = ~po17  & n13823;
  assign n13832 = ~n13830 & ~n13831;
  assign n13833 = ~n13824 & ~n13832;
  assign n13834 = po18  & ~n13833;
  assign n13835 = ~n13284 & ~n13291;
  assign n13836 = n13290 & n13835;
  assign n13837 = po13  & n13836;
  assign n13838 = po13  & n13835;
  assign n13839 = ~n13290 & ~n13838;
  assign n13840 = ~n13837 & ~n13839;
  assign n13841 = ~po18  & ~n13824;
  assign n13842 = ~n13832 & n13841;
  assign n13843 = ~n13840 & ~n13842;
  assign n13844 = ~n13834 & ~n13843;
  assign n13845 = po19  & ~n13844;
  assign n13846 = ~n13294 & ~n13302;
  assign n13847 = n13300 & n13846;
  assign n13848 = po13  & n13847;
  assign n13849 = po13  & n13846;
  assign n13850 = ~n13300 & ~n13849;
  assign n13851 = ~n13848 & ~n13850;
  assign n13852 = ~po19  & n13844;
  assign n13853 = ~n13851 & ~n13852;
  assign n13854 = ~n13845 & ~n13853;
  assign n13855 = po20  & ~n13854;
  assign n13856 = ~n13305 & ~n13312;
  assign n13857 = n13311 & n13856;
  assign n13858 = po13  & n13857;
  assign n13859 = po13  & n13856;
  assign n13860 = ~n13311 & ~n13859;
  assign n13861 = ~n13858 & ~n13860;
  assign n13862 = ~po20  & ~n13845;
  assign n13863 = ~n13853 & n13862;
  assign n13864 = ~n13861 & ~n13863;
  assign n13865 = ~n13855 & ~n13864;
  assign n13866 = po21  & ~n13865;
  assign n13867 = ~n13315 & ~n13323;
  assign n13868 = n13321 & n13867;
  assign n13869 = po13  & n13868;
  assign n13870 = po13  & n13867;
  assign n13871 = ~n13321 & ~n13870;
  assign n13872 = ~n13869 & ~n13871;
  assign n13873 = ~po21  & n13865;
  assign n13874 = ~n13872 & ~n13873;
  assign n13875 = ~n13866 & ~n13874;
  assign n13876 = po22  & ~n13875;
  assign n13877 = ~n13326 & ~n13333;
  assign n13878 = n13332 & n13877;
  assign n13879 = po13  & n13878;
  assign n13880 = po13  & n13877;
  assign n13881 = ~n13332 & ~n13880;
  assign n13882 = ~n13879 & ~n13881;
  assign n13883 = ~po22  & ~n13866;
  assign n13884 = ~n13874 & n13883;
  assign n13885 = ~n13882 & ~n13884;
  assign n13886 = ~n13876 & ~n13885;
  assign n13887 = po23  & ~n13886;
  assign n13888 = ~n13336 & ~n13344;
  assign n13889 = n13342 & n13888;
  assign n13890 = po13  & n13889;
  assign n13891 = po13  & n13888;
  assign n13892 = ~n13342 & ~n13891;
  assign n13893 = ~n13890 & ~n13892;
  assign n13894 = ~po23  & n13886;
  assign n13895 = ~n13893 & ~n13894;
  assign n13896 = ~n13887 & ~n13895;
  assign n13897 = po24  & ~n13896;
  assign n13898 = ~n13347 & ~n13354;
  assign n13899 = n13353 & n13898;
  assign n13900 = po13  & n13899;
  assign n13901 = po13  & n13898;
  assign n13902 = ~n13353 & ~n13901;
  assign n13903 = ~n13900 & ~n13902;
  assign n13904 = ~po24  & ~n13887;
  assign n13905 = ~n13895 & n13904;
  assign n13906 = ~n13903 & ~n13905;
  assign n13907 = ~n13897 & ~n13906;
  assign n13908 = po25  & ~n13907;
  assign n13909 = ~n13357 & ~n13365;
  assign n13910 = n13363 & n13909;
  assign n13911 = po13  & n13910;
  assign n13912 = po13  & n13909;
  assign n13913 = ~n13363 & ~n13912;
  assign n13914 = ~n13911 & ~n13913;
  assign n13915 = ~po25  & n13907;
  assign n13916 = ~n13914 & ~n13915;
  assign n13917 = ~n13908 & ~n13916;
  assign n13918 = po26  & ~n13917;
  assign n13919 = ~n13368 & ~n13375;
  assign n13920 = n13374 & n13919;
  assign n13921 = po13  & n13920;
  assign n13922 = po13  & n13919;
  assign n13923 = ~n13374 & ~n13922;
  assign n13924 = ~n13921 & ~n13923;
  assign n13925 = ~po26  & ~n13908;
  assign n13926 = ~n13916 & n13925;
  assign n13927 = ~n13924 & ~n13926;
  assign n13928 = ~n13918 & ~n13927;
  assign n13929 = po27  & ~n13928;
  assign n13930 = ~n13378 & ~n13386;
  assign n13931 = n13384 & n13930;
  assign n13932 = po13  & n13931;
  assign n13933 = po13  & n13930;
  assign n13934 = ~n13384 & ~n13933;
  assign n13935 = ~n13932 & ~n13934;
  assign n13936 = ~po27  & n13928;
  assign n13937 = ~n13935 & ~n13936;
  assign n13938 = ~n13929 & ~n13937;
  assign n13939 = po28  & ~n13938;
  assign n13940 = ~n13389 & ~n13396;
  assign n13941 = n13395 & n13940;
  assign n13942 = po13  & n13941;
  assign n13943 = po13  & n13940;
  assign n13944 = ~n13395 & ~n13943;
  assign n13945 = ~n13942 & ~n13944;
  assign n13946 = ~po28  & ~n13929;
  assign n13947 = ~n13937 & n13946;
  assign n13948 = ~n13945 & ~n13947;
  assign n13949 = ~n13939 & ~n13948;
  assign n13950 = po29  & ~n13949;
  assign n13951 = ~n13399 & ~n13407;
  assign n13952 = n13405 & n13951;
  assign n13953 = po13  & n13952;
  assign n13954 = po13  & n13951;
  assign n13955 = ~n13405 & ~n13954;
  assign n13956 = ~n13953 & ~n13955;
  assign n13957 = ~po29  & n13949;
  assign n13958 = ~n13956 & ~n13957;
  assign n13959 = ~n13950 & ~n13958;
  assign n13960 = po30  & ~n13959;
  assign n13961 = ~n13410 & ~n13417;
  assign n13962 = n13416 & n13961;
  assign n13963 = po13  & n13962;
  assign n13964 = po13  & n13961;
  assign n13965 = ~n13416 & ~n13964;
  assign n13966 = ~n13963 & ~n13965;
  assign n13967 = ~po30  & ~n13950;
  assign n13968 = ~n13958 & n13967;
  assign n13969 = ~n13966 & ~n13968;
  assign n13970 = ~n13960 & ~n13969;
  assign n13971 = po31  & ~n13970;
  assign n13972 = ~n13420 & ~n13428;
  assign n13973 = n13426 & n13972;
  assign n13974 = po13  & n13973;
  assign n13975 = po13  & n13972;
  assign n13976 = ~n13426 & ~n13975;
  assign n13977 = ~n13974 & ~n13976;
  assign n13978 = ~po31  & n13970;
  assign n13979 = ~n13977 & ~n13978;
  assign n13980 = ~n13971 & ~n13979;
  assign n13981 = po32  & ~n13980;
  assign n13982 = ~n13431 & ~n13438;
  assign n13983 = n13437 & n13982;
  assign n13984 = po13  & n13983;
  assign n13985 = po13  & n13982;
  assign n13986 = ~n13437 & ~n13985;
  assign n13987 = ~n13984 & ~n13986;
  assign n13988 = ~po32  & ~n13971;
  assign n13989 = ~n13979 & n13988;
  assign n13990 = ~n13987 & ~n13989;
  assign n13991 = ~n13981 & ~n13990;
  assign n13992 = po33  & ~n13991;
  assign n13993 = ~n13441 & ~n13449;
  assign n13994 = n13447 & n13993;
  assign n13995 = po13  & n13994;
  assign n13996 = po13  & n13993;
  assign n13997 = ~n13447 & ~n13996;
  assign n13998 = ~n13995 & ~n13997;
  assign n13999 = ~po33  & n13991;
  assign n14000 = ~n13998 & ~n13999;
  assign n14001 = ~n13992 & ~n14000;
  assign n14002 = po34  & ~n14001;
  assign n14003 = ~n13452 & ~n13459;
  assign n14004 = n13458 & n14003;
  assign n14005 = po13  & n14004;
  assign n14006 = po13  & n14003;
  assign n14007 = ~n13458 & ~n14006;
  assign n14008 = ~n14005 & ~n14007;
  assign n14009 = ~po34  & ~n13992;
  assign n14010 = ~n14000 & n14009;
  assign n14011 = ~n14008 & ~n14010;
  assign n14012 = ~n14002 & ~n14011;
  assign n14013 = po35  & ~n14012;
  assign n14014 = ~n13462 & ~n13470;
  assign n14015 = n13468 & n14014;
  assign n14016 = po13  & n14015;
  assign n14017 = po13  & n14014;
  assign n14018 = ~n13468 & ~n14017;
  assign n14019 = ~n14016 & ~n14018;
  assign n14020 = ~po35  & n14012;
  assign n14021 = ~n14019 & ~n14020;
  assign n14022 = ~n14013 & ~n14021;
  assign n14023 = po36  & ~n14022;
  assign n14024 = ~n13473 & ~n13480;
  assign n14025 = n13479 & n14024;
  assign n14026 = po13  & n14025;
  assign n14027 = po13  & n14024;
  assign n14028 = ~n13479 & ~n14027;
  assign n14029 = ~n14026 & ~n14028;
  assign n14030 = ~po36  & ~n14013;
  assign n14031 = ~n14021 & n14030;
  assign n14032 = ~n14029 & ~n14031;
  assign n14033 = ~n14023 & ~n14032;
  assign n14034 = po37  & ~n14033;
  assign n14035 = ~n13483 & ~n13491;
  assign n14036 = n13489 & n14035;
  assign n14037 = po13  & n14036;
  assign n14038 = po13  & n14035;
  assign n14039 = ~n13489 & ~n14038;
  assign n14040 = ~n14037 & ~n14039;
  assign n14041 = ~po37  & n14033;
  assign n14042 = ~n14040 & ~n14041;
  assign n14043 = ~n14034 & ~n14042;
  assign n14044 = po38  & ~n14043;
  assign n14045 = ~n13494 & ~n13501;
  assign n14046 = n13500 & n14045;
  assign n14047 = po13  & n14046;
  assign n14048 = po13  & n14045;
  assign n14049 = ~n13500 & ~n14048;
  assign n14050 = ~n14047 & ~n14049;
  assign n14051 = ~po38  & ~n14034;
  assign n14052 = ~n14042 & n14051;
  assign n14053 = ~n14050 & ~n14052;
  assign n14054 = ~n14044 & ~n14053;
  assign n14055 = po39  & ~n14054;
  assign n14056 = ~n13504 & ~n13512;
  assign n14057 = n13510 & n14056;
  assign n14058 = po13  & n14057;
  assign n14059 = po13  & n14056;
  assign n14060 = ~n13510 & ~n14059;
  assign n14061 = ~n14058 & ~n14060;
  assign n14062 = ~po39  & n14054;
  assign n14063 = ~n14061 & ~n14062;
  assign n14064 = ~n14055 & ~n14063;
  assign n14065 = po40  & ~n14064;
  assign n14066 = ~n13515 & ~n13522;
  assign n14067 = n13521 & n14066;
  assign n14068 = po13  & n14067;
  assign n14069 = po13  & n14066;
  assign n14070 = ~n13521 & ~n14069;
  assign n14071 = ~n14068 & ~n14070;
  assign n14072 = ~po40  & ~n14055;
  assign n14073 = ~n14063 & n14072;
  assign n14074 = ~n14071 & ~n14073;
  assign n14075 = ~n14065 & ~n14074;
  assign n14076 = po41  & ~n14075;
  assign n14077 = ~n13525 & ~n13533;
  assign n14078 = n13531 & n14077;
  assign n14079 = po13  & n14078;
  assign n14080 = po13  & n14077;
  assign n14081 = ~n13531 & ~n14080;
  assign n14082 = ~n14079 & ~n14081;
  assign n14083 = ~po41  & n14075;
  assign n14084 = ~n14082 & ~n14083;
  assign n14085 = ~n14076 & ~n14084;
  assign n14086 = po42  & ~n14085;
  assign n14087 = ~n13536 & ~n13543;
  assign n14088 = n13542 & n14087;
  assign n14089 = po13  & n14088;
  assign n14090 = po13  & n14087;
  assign n14091 = ~n13542 & ~n14090;
  assign n14092 = ~n14089 & ~n14091;
  assign n14093 = ~po42  & ~n14076;
  assign n14094 = ~n14084 & n14093;
  assign n14095 = ~n14092 & ~n14094;
  assign n14096 = ~n14086 & ~n14095;
  assign n14097 = po43  & ~n14096;
  assign n14098 = ~n13546 & ~n13554;
  assign n14099 = n13552 & n14098;
  assign n14100 = po13  & n14099;
  assign n14101 = po13  & n14098;
  assign n14102 = ~n13552 & ~n14101;
  assign n14103 = ~n14100 & ~n14102;
  assign n14104 = ~po43  & n14096;
  assign n14105 = ~n14103 & ~n14104;
  assign n14106 = ~n14097 & ~n14105;
  assign n14107 = po44  & ~n14106;
  assign n14108 = ~n13557 & ~n13564;
  assign n14109 = n13563 & n14108;
  assign n14110 = po13  & n14109;
  assign n14111 = po13  & n14108;
  assign n14112 = ~n13563 & ~n14111;
  assign n14113 = ~n14110 & ~n14112;
  assign n14114 = ~po44  & ~n14097;
  assign n14115 = ~n14105 & n14114;
  assign n14116 = ~n14113 & ~n14115;
  assign n14117 = ~n14107 & ~n14116;
  assign n14118 = po45  & ~n14117;
  assign n14119 = ~n13567 & ~n13575;
  assign n14120 = n13573 & n14119;
  assign n14121 = po13  & n14120;
  assign n14122 = po13  & n14119;
  assign n14123 = ~n13573 & ~n14122;
  assign n14124 = ~n14121 & ~n14123;
  assign n14125 = ~po45  & n14117;
  assign n14126 = ~n14124 & ~n14125;
  assign n14127 = ~n14118 & ~n14126;
  assign n14128 = po46  & ~n14127;
  assign n14129 = ~n13578 & ~n13585;
  assign n14130 = n13584 & n14129;
  assign n14131 = po13  & n14130;
  assign n14132 = po13  & n14129;
  assign n14133 = ~n13584 & ~n14132;
  assign n14134 = ~n14131 & ~n14133;
  assign n14135 = ~po46  & ~n14118;
  assign n14136 = ~n14126 & n14135;
  assign n14137 = ~n14134 & ~n14136;
  assign n14138 = ~n14128 & ~n14137;
  assign n14139 = po47  & ~n14138;
  assign n14140 = ~n13588 & ~n13596;
  assign n14141 = n13594 & n14140;
  assign n14142 = po13  & n14141;
  assign n14143 = po13  & n14140;
  assign n14144 = ~n13594 & ~n14143;
  assign n14145 = ~n14142 & ~n14144;
  assign n14146 = ~po47  & n14138;
  assign n14147 = ~n14145 & ~n14146;
  assign n14148 = ~n14139 & ~n14147;
  assign n14149 = po48  & ~n14148;
  assign n14150 = ~n13599 & ~n13606;
  assign n14151 = n13605 & n14150;
  assign n14152 = po13  & n14151;
  assign n14153 = po13  & n14150;
  assign n14154 = ~n13605 & ~n14153;
  assign n14155 = ~n14152 & ~n14154;
  assign n14156 = ~po48  & ~n14139;
  assign n14157 = ~n14147 & n14156;
  assign n14158 = ~n14155 & ~n14157;
  assign n14159 = ~n14149 & ~n14158;
  assign n14160 = po49  & ~n14159;
  assign n14161 = ~n13609 & ~n13617;
  assign n14162 = n13615 & n14161;
  assign n14163 = po13  & n14162;
  assign n14164 = po13  & n14161;
  assign n14165 = ~n13615 & ~n14164;
  assign n14166 = ~n14163 & ~n14165;
  assign n14167 = ~po49  & n14159;
  assign n14168 = ~n14166 & ~n14167;
  assign n14169 = ~n14160 & ~n14168;
  assign n14170 = po50  & ~n14169;
  assign n14171 = ~n13620 & ~n13627;
  assign n14172 = n13626 & n14171;
  assign n14173 = po13  & n14172;
  assign n14174 = po13  & n14171;
  assign n14175 = ~n13626 & ~n14174;
  assign n14176 = ~n14173 & ~n14175;
  assign n14177 = ~po50  & ~n14160;
  assign n14178 = ~n14168 & n14177;
  assign n14179 = ~n14176 & ~n14178;
  assign n14180 = ~n14170 & ~n14179;
  assign n14181 = po51  & ~n14180;
  assign n14182 = ~n13630 & ~n13638;
  assign n14183 = n13636 & n14182;
  assign n14184 = po13  & n14183;
  assign n14185 = po13  & n14182;
  assign n14186 = ~n13636 & ~n14185;
  assign n14187 = ~n14184 & ~n14186;
  assign n14188 = ~po51  & n14180;
  assign n14189 = ~n14187 & ~n14188;
  assign n14190 = ~n14181 & ~n14189;
  assign n14191 = po52  & ~n14190;
  assign n14192 = ~po52  & ~n14181;
  assign n14193 = ~n14189 & n14192;
  assign n14194 = ~n13641 & ~n13648;
  assign n14195 = n13647 & n14194;
  assign n14196 = po13  & n14195;
  assign n14197 = po13  & n14194;
  assign n14198 = ~n13647 & ~n14197;
  assign n14199 = ~n14196 & ~n14198;
  assign n14200 = ~n14193 & ~n14199;
  assign n14201 = ~n14191 & ~n14200;
  assign n14202 = po53  & ~n14201;
  assign n14203 = ~n13651 & ~n13659;
  assign n14204 = n13657 & n14203;
  assign n14205 = po13  & n14204;
  assign n14206 = po13  & n14203;
  assign n14207 = ~n13657 & ~n14206;
  assign n14208 = ~n14205 & ~n14207;
  assign n14209 = ~po53  & n14201;
  assign n14210 = ~n14208 & ~n14209;
  assign n14211 = ~n14202 & ~n14210;
  assign n14212 = po54  & ~n14211;
  assign n14213 = ~n13662 & ~n13669;
  assign n14214 = n13668 & n14213;
  assign n14215 = po13  & n14214;
  assign n14216 = po13  & n14213;
  assign n14217 = ~n13668 & ~n14216;
  assign n14218 = ~n14215 & ~n14217;
  assign n14219 = ~po54  & ~n14202;
  assign n14220 = ~n14210 & n14219;
  assign n14221 = ~n14218 & ~n14220;
  assign n14222 = ~n14212 & ~n14221;
  assign n14223 = po55  & ~n14222;
  assign n14224 = ~n13672 & ~n13680;
  assign n14225 = n13678 & n14224;
  assign n14226 = po13  & n14225;
  assign n14227 = po13  & n14224;
  assign n14228 = ~n13678 & ~n14227;
  assign n14229 = ~n14226 & ~n14228;
  assign n14230 = ~po55  & n14222;
  assign n14231 = ~n14229 & ~n14230;
  assign n14232 = ~n14223 & ~n14231;
  assign n14233 = po56  & ~n14232;
  assign n14234 = ~n13683 & ~n13690;
  assign n14235 = n13689 & n14234;
  assign n14236 = po13  & n14235;
  assign n14237 = po13  & n14234;
  assign n14238 = ~n13689 & ~n14237;
  assign n14239 = ~n14236 & ~n14238;
  assign n14240 = ~po56  & ~n14223;
  assign n14241 = ~n14231 & n14240;
  assign n14242 = ~n14239 & ~n14241;
  assign n14243 = ~n14233 & ~n14242;
  assign n14244 = po57  & ~n14243;
  assign n14245 = ~n13693 & ~n13701;
  assign n14246 = n13699 & n14245;
  assign n14247 = po13  & n14246;
  assign n14248 = po13  & n14245;
  assign n14249 = ~n13699 & ~n14248;
  assign n14250 = ~n14247 & ~n14249;
  assign n14251 = ~po57  & n14243;
  assign n14252 = ~n14250 & ~n14251;
  assign n14253 = ~n14244 & ~n14252;
  assign n14254 = po58  & ~n14253;
  assign n14255 = ~n13704 & ~n13711;
  assign n14256 = n13710 & n14255;
  assign n14257 = po13  & n14256;
  assign n14258 = po13  & n14255;
  assign n14259 = ~n13710 & ~n14258;
  assign n14260 = ~n14257 & ~n14259;
  assign n14261 = ~po58  & ~n14244;
  assign n14262 = ~n14252 & n14261;
  assign n14263 = ~n14260 & ~n14262;
  assign n14264 = ~n14254 & ~n14263;
  assign n14265 = po59  & ~n14264;
  assign n14266 = ~n13714 & ~n13722;
  assign n14267 = n13720 & n14266;
  assign n14268 = po13  & n14267;
  assign n14269 = po13  & n14266;
  assign n14270 = ~n13720 & ~n14269;
  assign n14271 = ~n14268 & ~n14270;
  assign n14272 = ~po59  & n14264;
  assign n14273 = ~n14271 & ~n14272;
  assign n14274 = ~n14265 & ~n14273;
  assign n14275 = po60  & ~n14274;
  assign n14276 = ~n13725 & ~n13732;
  assign n14277 = n13731 & n14276;
  assign n14278 = po13  & n14277;
  assign n14279 = po13  & n14276;
  assign n14280 = ~n13731 & ~n14279;
  assign n14281 = ~n14278 & ~n14280;
  assign n14282 = ~po60  & ~n14265;
  assign n14283 = ~n14273 & n14282;
  assign n14284 = ~n14281 & ~n14283;
  assign n14285 = ~n14275 & ~n14284;
  assign n14286 = po61  & ~n14285;
  assign n14287 = ~n13735 & ~n13743;
  assign n14288 = n13741 & n14287;
  assign n14289 = po13  & n14288;
  assign n14290 = po13  & n14287;
  assign n14291 = ~n13741 & ~n14290;
  assign n14292 = ~n14289 & ~n14291;
  assign n14293 = ~po61  & n14285;
  assign n14294 = ~n14292 & ~n14293;
  assign n14295 = ~n14286 & ~n14294;
  assign n14296 = po62  & ~n14295;
  assign n14297 = ~n13746 & ~n13753;
  assign n14298 = n13752 & n14297;
  assign n14299 = po13  & n14298;
  assign n14300 = po13  & n14297;
  assign n14301 = ~n13752 & ~n14300;
  assign n14302 = ~n14299 & ~n14301;
  assign n14303 = ~po62  & ~n14286;
  assign n14304 = ~n14294 & n14303;
  assign n14305 = ~n14302 & ~n14304;
  assign n14306 = ~n14296 & ~n14305;
  assign n14307 = ~n13756 & ~n13764;
  assign n14308 = po13  & n14307;
  assign n14309 = ~n13762 & ~n14308;
  assign n14310 = n13762 & n14308;
  assign n14311 = ~n14309 & ~n14310;
  assign n14312 = ~n13766 & ~n13771;
  assign n14313 = po13  & n14312;
  assign n14314 = ~n13784 & ~n14313;
  assign n14315 = ~n14311 & n14314;
  assign n14316 = ~n14306 & n14315;
  assign n14317 = ~po63  & ~n14316;
  assign n14318 = ~n13771 & po13 ;
  assign n14319 = n13766 & ~n14318;
  assign n14320 = po63  & ~n14312;
  assign n14321 = ~n14319 & n14320;
  assign n14322 = n13771 & ~po13 ;
  assign n14323 = ~n14321 & ~n14322;
  assign n14324 = n14306 & n14311;
  assign n14325 = n14323 & ~n14324;
  assign po12  = n14317 | ~n14325;
  assign n14327 = pi24  & po12 ;
  assign n14328 = ~pi22  & ~pi23 ;
  assign n14329 = ~pi24  & n14328;
  assign n14330 = ~n14327 & ~n14329;
  assign n14331 = po13  & ~n14330;
  assign n14332 = n13783 & ~n14329;
  assign n14333 = ~n13784 & n14332;
  assign n14334 = ~n13777 & n14333;
  assign n14335 = ~n14327 & n14334;
  assign n14336 = ~pi24  & po12 ;
  assign n14337 = pi25  & ~n14336;
  assign n14338 = n13788 & po12 ;
  assign n14339 = ~n14337 & ~n14338;
  assign n14340 = ~n14335 & n14339;
  assign n14341 = ~n14331 & ~n14340;
  assign n14342 = po14  & ~n14341;
  assign n14343 = ~po14  & ~n14331;
  assign n14344 = ~n14340 & n14343;
  assign n14345 = po13  & n14323;
  assign n14346 = ~n14324 & n14345;
  assign n14347 = ~n14317 & n14346;
  assign n14348 = ~n14338 & ~n14347;
  assign n14349 = pi26  & ~n14348;
  assign n14350 = ~pi26  & n14348;
  assign n14351 = ~n14349 & ~n14350;
  assign n14352 = ~n14344 & ~n14351;
  assign n14353 = ~n14342 & ~n14352;
  assign n14354 = po15  & ~n14353;
  assign n14355 = ~n13791 & ~n13795;
  assign n14356 = ~n13799 & n14355;
  assign n14357 = po12  & n14356;
  assign n14358 = po12  & n14355;
  assign n14359 = n13799 & ~n14358;
  assign n14360 = ~n14357 & ~n14359;
  assign n14361 = ~po15  & n14353;
  assign n14362 = ~n14360 & ~n14361;
  assign n14363 = ~n14354 & ~n14362;
  assign n14364 = po16  & ~n14363;
  assign n14365 = ~n13802 & ~n13810;
  assign n14366 = n13809 & n14365;
  assign n14367 = po12  & n14366;
  assign n14368 = po12  & n14365;
  assign n14369 = ~n13809 & ~n14368;
  assign n14370 = ~n14367 & ~n14369;
  assign n14371 = ~po16  & ~n14354;
  assign n14372 = ~n14362 & n14371;
  assign n14373 = ~n14370 & ~n14372;
  assign n14374 = ~n14364 & ~n14373;
  assign n14375 = po17  & ~n14374;
  assign n14376 = ~n13813 & ~n13821;
  assign n14377 = n13819 & n14376;
  assign n14378 = po12  & n14377;
  assign n14379 = po12  & n14376;
  assign n14380 = ~n13819 & ~n14379;
  assign n14381 = ~n14378 & ~n14380;
  assign n14382 = ~po17  & n14374;
  assign n14383 = ~n14381 & ~n14382;
  assign n14384 = ~n14375 & ~n14383;
  assign n14385 = po18  & ~n14384;
  assign n14386 = ~n13824 & ~n13831;
  assign n14387 = n13830 & n14386;
  assign n14388 = po12  & n14387;
  assign n14389 = po12  & n14386;
  assign n14390 = ~n13830 & ~n14389;
  assign n14391 = ~n14388 & ~n14390;
  assign n14392 = ~po18  & ~n14375;
  assign n14393 = ~n14383 & n14392;
  assign n14394 = ~n14391 & ~n14393;
  assign n14395 = ~n14385 & ~n14394;
  assign n14396 = po19  & ~n14395;
  assign n14397 = ~n13834 & ~n13842;
  assign n14398 = n13840 & n14397;
  assign n14399 = po12  & n14398;
  assign n14400 = po12  & n14397;
  assign n14401 = ~n13840 & ~n14400;
  assign n14402 = ~n14399 & ~n14401;
  assign n14403 = ~po19  & n14395;
  assign n14404 = ~n14402 & ~n14403;
  assign n14405 = ~n14396 & ~n14404;
  assign n14406 = po20  & ~n14405;
  assign n14407 = ~n13845 & ~n13852;
  assign n14408 = n13851 & n14407;
  assign n14409 = po12  & n14408;
  assign n14410 = po12  & n14407;
  assign n14411 = ~n13851 & ~n14410;
  assign n14412 = ~n14409 & ~n14411;
  assign n14413 = ~po20  & ~n14396;
  assign n14414 = ~n14404 & n14413;
  assign n14415 = ~n14412 & ~n14414;
  assign n14416 = ~n14406 & ~n14415;
  assign n14417 = po21  & ~n14416;
  assign n14418 = ~n13855 & ~n13863;
  assign n14419 = n13861 & n14418;
  assign n14420 = po12  & n14419;
  assign n14421 = po12  & n14418;
  assign n14422 = ~n13861 & ~n14421;
  assign n14423 = ~n14420 & ~n14422;
  assign n14424 = ~po21  & n14416;
  assign n14425 = ~n14423 & ~n14424;
  assign n14426 = ~n14417 & ~n14425;
  assign n14427 = po22  & ~n14426;
  assign n14428 = ~n13866 & ~n13873;
  assign n14429 = n13872 & n14428;
  assign n14430 = po12  & n14429;
  assign n14431 = po12  & n14428;
  assign n14432 = ~n13872 & ~n14431;
  assign n14433 = ~n14430 & ~n14432;
  assign n14434 = ~po22  & ~n14417;
  assign n14435 = ~n14425 & n14434;
  assign n14436 = ~n14433 & ~n14435;
  assign n14437 = ~n14427 & ~n14436;
  assign n14438 = po23  & ~n14437;
  assign n14439 = ~n13876 & ~n13884;
  assign n14440 = n13882 & n14439;
  assign n14441 = po12  & n14440;
  assign n14442 = po12  & n14439;
  assign n14443 = ~n13882 & ~n14442;
  assign n14444 = ~n14441 & ~n14443;
  assign n14445 = ~po23  & n14437;
  assign n14446 = ~n14444 & ~n14445;
  assign n14447 = ~n14438 & ~n14446;
  assign n14448 = po24  & ~n14447;
  assign n14449 = ~n13887 & ~n13894;
  assign n14450 = n13893 & n14449;
  assign n14451 = po12  & n14450;
  assign n14452 = po12  & n14449;
  assign n14453 = ~n13893 & ~n14452;
  assign n14454 = ~n14451 & ~n14453;
  assign n14455 = ~po24  & ~n14438;
  assign n14456 = ~n14446 & n14455;
  assign n14457 = ~n14454 & ~n14456;
  assign n14458 = ~n14448 & ~n14457;
  assign n14459 = po25  & ~n14458;
  assign n14460 = ~n13897 & ~n13905;
  assign n14461 = n13903 & n14460;
  assign n14462 = po12  & n14461;
  assign n14463 = po12  & n14460;
  assign n14464 = ~n13903 & ~n14463;
  assign n14465 = ~n14462 & ~n14464;
  assign n14466 = ~po25  & n14458;
  assign n14467 = ~n14465 & ~n14466;
  assign n14468 = ~n14459 & ~n14467;
  assign n14469 = po26  & ~n14468;
  assign n14470 = ~n13908 & ~n13915;
  assign n14471 = n13914 & n14470;
  assign n14472 = po12  & n14471;
  assign n14473 = po12  & n14470;
  assign n14474 = ~n13914 & ~n14473;
  assign n14475 = ~n14472 & ~n14474;
  assign n14476 = ~po26  & ~n14459;
  assign n14477 = ~n14467 & n14476;
  assign n14478 = ~n14475 & ~n14477;
  assign n14479 = ~n14469 & ~n14478;
  assign n14480 = po27  & ~n14479;
  assign n14481 = ~n13918 & ~n13926;
  assign n14482 = n13924 & n14481;
  assign n14483 = po12  & n14482;
  assign n14484 = po12  & n14481;
  assign n14485 = ~n13924 & ~n14484;
  assign n14486 = ~n14483 & ~n14485;
  assign n14487 = ~po27  & n14479;
  assign n14488 = ~n14486 & ~n14487;
  assign n14489 = ~n14480 & ~n14488;
  assign n14490 = po28  & ~n14489;
  assign n14491 = ~n13929 & ~n13936;
  assign n14492 = n13935 & n14491;
  assign n14493 = po12  & n14492;
  assign n14494 = po12  & n14491;
  assign n14495 = ~n13935 & ~n14494;
  assign n14496 = ~n14493 & ~n14495;
  assign n14497 = ~po28  & ~n14480;
  assign n14498 = ~n14488 & n14497;
  assign n14499 = ~n14496 & ~n14498;
  assign n14500 = ~n14490 & ~n14499;
  assign n14501 = po29  & ~n14500;
  assign n14502 = ~n13939 & ~n13947;
  assign n14503 = n13945 & n14502;
  assign n14504 = po12  & n14503;
  assign n14505 = po12  & n14502;
  assign n14506 = ~n13945 & ~n14505;
  assign n14507 = ~n14504 & ~n14506;
  assign n14508 = ~po29  & n14500;
  assign n14509 = ~n14507 & ~n14508;
  assign n14510 = ~n14501 & ~n14509;
  assign n14511 = po30  & ~n14510;
  assign n14512 = ~n13950 & ~n13957;
  assign n14513 = n13956 & n14512;
  assign n14514 = po12  & n14513;
  assign n14515 = po12  & n14512;
  assign n14516 = ~n13956 & ~n14515;
  assign n14517 = ~n14514 & ~n14516;
  assign n14518 = ~po30  & ~n14501;
  assign n14519 = ~n14509 & n14518;
  assign n14520 = ~n14517 & ~n14519;
  assign n14521 = ~n14511 & ~n14520;
  assign n14522 = po31  & ~n14521;
  assign n14523 = ~n13960 & ~n13968;
  assign n14524 = n13966 & n14523;
  assign n14525 = po12  & n14524;
  assign n14526 = po12  & n14523;
  assign n14527 = ~n13966 & ~n14526;
  assign n14528 = ~n14525 & ~n14527;
  assign n14529 = ~po31  & n14521;
  assign n14530 = ~n14528 & ~n14529;
  assign n14531 = ~n14522 & ~n14530;
  assign n14532 = po32  & ~n14531;
  assign n14533 = ~n13971 & ~n13978;
  assign n14534 = n13977 & n14533;
  assign n14535 = po12  & n14534;
  assign n14536 = po12  & n14533;
  assign n14537 = ~n13977 & ~n14536;
  assign n14538 = ~n14535 & ~n14537;
  assign n14539 = ~po32  & ~n14522;
  assign n14540 = ~n14530 & n14539;
  assign n14541 = ~n14538 & ~n14540;
  assign n14542 = ~n14532 & ~n14541;
  assign n14543 = po33  & ~n14542;
  assign n14544 = ~n13981 & ~n13989;
  assign n14545 = n13987 & n14544;
  assign n14546 = po12  & n14545;
  assign n14547 = po12  & n14544;
  assign n14548 = ~n13987 & ~n14547;
  assign n14549 = ~n14546 & ~n14548;
  assign n14550 = ~po33  & n14542;
  assign n14551 = ~n14549 & ~n14550;
  assign n14552 = ~n14543 & ~n14551;
  assign n14553 = po34  & ~n14552;
  assign n14554 = ~n13992 & ~n13999;
  assign n14555 = n13998 & n14554;
  assign n14556 = po12  & n14555;
  assign n14557 = po12  & n14554;
  assign n14558 = ~n13998 & ~n14557;
  assign n14559 = ~n14556 & ~n14558;
  assign n14560 = ~po34  & ~n14543;
  assign n14561 = ~n14551 & n14560;
  assign n14562 = ~n14559 & ~n14561;
  assign n14563 = ~n14553 & ~n14562;
  assign n14564 = po35  & ~n14563;
  assign n14565 = ~n14002 & ~n14010;
  assign n14566 = n14008 & n14565;
  assign n14567 = po12  & n14566;
  assign n14568 = po12  & n14565;
  assign n14569 = ~n14008 & ~n14568;
  assign n14570 = ~n14567 & ~n14569;
  assign n14571 = ~po35  & n14563;
  assign n14572 = ~n14570 & ~n14571;
  assign n14573 = ~n14564 & ~n14572;
  assign n14574 = po36  & ~n14573;
  assign n14575 = ~n14013 & ~n14020;
  assign n14576 = n14019 & n14575;
  assign n14577 = po12  & n14576;
  assign n14578 = po12  & n14575;
  assign n14579 = ~n14019 & ~n14578;
  assign n14580 = ~n14577 & ~n14579;
  assign n14581 = ~po36  & ~n14564;
  assign n14582 = ~n14572 & n14581;
  assign n14583 = ~n14580 & ~n14582;
  assign n14584 = ~n14574 & ~n14583;
  assign n14585 = po37  & ~n14584;
  assign n14586 = ~n14023 & ~n14031;
  assign n14587 = n14029 & n14586;
  assign n14588 = po12  & n14587;
  assign n14589 = po12  & n14586;
  assign n14590 = ~n14029 & ~n14589;
  assign n14591 = ~n14588 & ~n14590;
  assign n14592 = ~po37  & n14584;
  assign n14593 = ~n14591 & ~n14592;
  assign n14594 = ~n14585 & ~n14593;
  assign n14595 = po38  & ~n14594;
  assign n14596 = ~n14034 & ~n14041;
  assign n14597 = n14040 & n14596;
  assign n14598 = po12  & n14597;
  assign n14599 = po12  & n14596;
  assign n14600 = ~n14040 & ~n14599;
  assign n14601 = ~n14598 & ~n14600;
  assign n14602 = ~po38  & ~n14585;
  assign n14603 = ~n14593 & n14602;
  assign n14604 = ~n14601 & ~n14603;
  assign n14605 = ~n14595 & ~n14604;
  assign n14606 = po39  & ~n14605;
  assign n14607 = ~n14044 & ~n14052;
  assign n14608 = n14050 & n14607;
  assign n14609 = po12  & n14608;
  assign n14610 = po12  & n14607;
  assign n14611 = ~n14050 & ~n14610;
  assign n14612 = ~n14609 & ~n14611;
  assign n14613 = ~po39  & n14605;
  assign n14614 = ~n14612 & ~n14613;
  assign n14615 = ~n14606 & ~n14614;
  assign n14616 = po40  & ~n14615;
  assign n14617 = ~n14055 & ~n14062;
  assign n14618 = n14061 & n14617;
  assign n14619 = po12  & n14618;
  assign n14620 = po12  & n14617;
  assign n14621 = ~n14061 & ~n14620;
  assign n14622 = ~n14619 & ~n14621;
  assign n14623 = ~po40  & ~n14606;
  assign n14624 = ~n14614 & n14623;
  assign n14625 = ~n14622 & ~n14624;
  assign n14626 = ~n14616 & ~n14625;
  assign n14627 = po41  & ~n14626;
  assign n14628 = ~n14065 & ~n14073;
  assign n14629 = n14071 & n14628;
  assign n14630 = po12  & n14629;
  assign n14631 = po12  & n14628;
  assign n14632 = ~n14071 & ~n14631;
  assign n14633 = ~n14630 & ~n14632;
  assign n14634 = ~po41  & n14626;
  assign n14635 = ~n14633 & ~n14634;
  assign n14636 = ~n14627 & ~n14635;
  assign n14637 = po42  & ~n14636;
  assign n14638 = ~n14076 & ~n14083;
  assign n14639 = n14082 & n14638;
  assign n14640 = po12  & n14639;
  assign n14641 = po12  & n14638;
  assign n14642 = ~n14082 & ~n14641;
  assign n14643 = ~n14640 & ~n14642;
  assign n14644 = ~po42  & ~n14627;
  assign n14645 = ~n14635 & n14644;
  assign n14646 = ~n14643 & ~n14645;
  assign n14647 = ~n14637 & ~n14646;
  assign n14648 = po43  & ~n14647;
  assign n14649 = ~n14086 & ~n14094;
  assign n14650 = n14092 & n14649;
  assign n14651 = po12  & n14650;
  assign n14652 = po12  & n14649;
  assign n14653 = ~n14092 & ~n14652;
  assign n14654 = ~n14651 & ~n14653;
  assign n14655 = ~po43  & n14647;
  assign n14656 = ~n14654 & ~n14655;
  assign n14657 = ~n14648 & ~n14656;
  assign n14658 = po44  & ~n14657;
  assign n14659 = ~n14097 & ~n14104;
  assign n14660 = n14103 & n14659;
  assign n14661 = po12  & n14660;
  assign n14662 = po12  & n14659;
  assign n14663 = ~n14103 & ~n14662;
  assign n14664 = ~n14661 & ~n14663;
  assign n14665 = ~po44  & ~n14648;
  assign n14666 = ~n14656 & n14665;
  assign n14667 = ~n14664 & ~n14666;
  assign n14668 = ~n14658 & ~n14667;
  assign n14669 = po45  & ~n14668;
  assign n14670 = ~n14107 & ~n14115;
  assign n14671 = n14113 & n14670;
  assign n14672 = po12  & n14671;
  assign n14673 = po12  & n14670;
  assign n14674 = ~n14113 & ~n14673;
  assign n14675 = ~n14672 & ~n14674;
  assign n14676 = ~po45  & n14668;
  assign n14677 = ~n14675 & ~n14676;
  assign n14678 = ~n14669 & ~n14677;
  assign n14679 = po46  & ~n14678;
  assign n14680 = ~n14118 & ~n14125;
  assign n14681 = n14124 & n14680;
  assign n14682 = po12  & n14681;
  assign n14683 = po12  & n14680;
  assign n14684 = ~n14124 & ~n14683;
  assign n14685 = ~n14682 & ~n14684;
  assign n14686 = ~po46  & ~n14669;
  assign n14687 = ~n14677 & n14686;
  assign n14688 = ~n14685 & ~n14687;
  assign n14689 = ~n14679 & ~n14688;
  assign n14690 = po47  & ~n14689;
  assign n14691 = ~n14128 & ~n14136;
  assign n14692 = n14134 & n14691;
  assign n14693 = po12  & n14692;
  assign n14694 = po12  & n14691;
  assign n14695 = ~n14134 & ~n14694;
  assign n14696 = ~n14693 & ~n14695;
  assign n14697 = ~po47  & n14689;
  assign n14698 = ~n14696 & ~n14697;
  assign n14699 = ~n14690 & ~n14698;
  assign n14700 = po48  & ~n14699;
  assign n14701 = ~n14139 & ~n14146;
  assign n14702 = n14145 & n14701;
  assign n14703 = po12  & n14702;
  assign n14704 = po12  & n14701;
  assign n14705 = ~n14145 & ~n14704;
  assign n14706 = ~n14703 & ~n14705;
  assign n14707 = ~po48  & ~n14690;
  assign n14708 = ~n14698 & n14707;
  assign n14709 = ~n14706 & ~n14708;
  assign n14710 = ~n14700 & ~n14709;
  assign n14711 = po49  & ~n14710;
  assign n14712 = ~n14149 & ~n14157;
  assign n14713 = n14155 & n14712;
  assign n14714 = po12  & n14713;
  assign n14715 = po12  & n14712;
  assign n14716 = ~n14155 & ~n14715;
  assign n14717 = ~n14714 & ~n14716;
  assign n14718 = ~po49  & n14710;
  assign n14719 = ~n14717 & ~n14718;
  assign n14720 = ~n14711 & ~n14719;
  assign n14721 = po50  & ~n14720;
  assign n14722 = ~n14160 & ~n14167;
  assign n14723 = n14166 & n14722;
  assign n14724 = po12  & n14723;
  assign n14725 = po12  & n14722;
  assign n14726 = ~n14166 & ~n14725;
  assign n14727 = ~n14724 & ~n14726;
  assign n14728 = ~po50  & ~n14711;
  assign n14729 = ~n14719 & n14728;
  assign n14730 = ~n14727 & ~n14729;
  assign n14731 = ~n14721 & ~n14730;
  assign n14732 = po51  & ~n14731;
  assign n14733 = ~n14170 & ~n14178;
  assign n14734 = n14176 & n14733;
  assign n14735 = po12  & n14734;
  assign n14736 = po12  & n14733;
  assign n14737 = ~n14176 & ~n14736;
  assign n14738 = ~n14735 & ~n14737;
  assign n14739 = ~po51  & n14731;
  assign n14740 = ~n14738 & ~n14739;
  assign n14741 = ~n14732 & ~n14740;
  assign n14742 = po52  & ~n14741;
  assign n14743 = ~n14181 & ~n14188;
  assign n14744 = n14187 & n14743;
  assign n14745 = po12  & n14744;
  assign n14746 = po12  & n14743;
  assign n14747 = ~n14187 & ~n14746;
  assign n14748 = ~n14745 & ~n14747;
  assign n14749 = ~po52  & ~n14732;
  assign n14750 = ~n14740 & n14749;
  assign n14751 = ~n14748 & ~n14750;
  assign n14752 = ~n14742 & ~n14751;
  assign n14753 = po53  & ~n14752;
  assign n14754 = ~n14191 & ~n14193;
  assign n14755 = n14199 & n14754;
  assign n14756 = po12  & n14755;
  assign n14757 = po12  & n14754;
  assign n14758 = ~n14199 & ~n14757;
  assign n14759 = ~n14756 & ~n14758;
  assign n14760 = ~po53  & n14752;
  assign n14761 = ~n14759 & ~n14760;
  assign n14762 = ~n14753 & ~n14761;
  assign n14763 = po54  & ~n14762;
  assign n14764 = ~n14202 & ~n14209;
  assign n14765 = n14208 & n14764;
  assign n14766 = po12  & n14765;
  assign n14767 = po12  & n14764;
  assign n14768 = ~n14208 & ~n14767;
  assign n14769 = ~n14766 & ~n14768;
  assign n14770 = ~po54  & ~n14753;
  assign n14771 = ~n14761 & n14770;
  assign n14772 = ~n14769 & ~n14771;
  assign n14773 = ~n14763 & ~n14772;
  assign n14774 = po55  & ~n14773;
  assign n14775 = ~n14212 & ~n14220;
  assign n14776 = n14218 & n14775;
  assign n14777 = po12  & n14776;
  assign n14778 = po12  & n14775;
  assign n14779 = ~n14218 & ~n14778;
  assign n14780 = ~n14777 & ~n14779;
  assign n14781 = ~po55  & n14773;
  assign n14782 = ~n14780 & ~n14781;
  assign n14783 = ~n14774 & ~n14782;
  assign n14784 = po56  & ~n14783;
  assign n14785 = ~n14223 & ~n14230;
  assign n14786 = n14229 & n14785;
  assign n14787 = po12  & n14786;
  assign n14788 = po12  & n14785;
  assign n14789 = ~n14229 & ~n14788;
  assign n14790 = ~n14787 & ~n14789;
  assign n14791 = ~po56  & ~n14774;
  assign n14792 = ~n14782 & n14791;
  assign n14793 = ~n14790 & ~n14792;
  assign n14794 = ~n14784 & ~n14793;
  assign n14795 = po57  & ~n14794;
  assign n14796 = ~n14233 & ~n14241;
  assign n14797 = n14239 & n14796;
  assign n14798 = po12  & n14797;
  assign n14799 = po12  & n14796;
  assign n14800 = ~n14239 & ~n14799;
  assign n14801 = ~n14798 & ~n14800;
  assign n14802 = ~po57  & n14794;
  assign n14803 = ~n14801 & ~n14802;
  assign n14804 = ~n14795 & ~n14803;
  assign n14805 = po58  & ~n14804;
  assign n14806 = ~n14244 & ~n14251;
  assign n14807 = n14250 & n14806;
  assign n14808 = po12  & n14807;
  assign n14809 = po12  & n14806;
  assign n14810 = ~n14250 & ~n14809;
  assign n14811 = ~n14808 & ~n14810;
  assign n14812 = ~po58  & ~n14795;
  assign n14813 = ~n14803 & n14812;
  assign n14814 = ~n14811 & ~n14813;
  assign n14815 = ~n14805 & ~n14814;
  assign n14816 = po59  & ~n14815;
  assign n14817 = ~n14254 & ~n14262;
  assign n14818 = n14260 & n14817;
  assign n14819 = po12  & n14818;
  assign n14820 = po12  & n14817;
  assign n14821 = ~n14260 & ~n14820;
  assign n14822 = ~n14819 & ~n14821;
  assign n14823 = ~po59  & n14815;
  assign n14824 = ~n14822 & ~n14823;
  assign n14825 = ~n14816 & ~n14824;
  assign n14826 = po60  & ~n14825;
  assign n14827 = ~n14265 & ~n14272;
  assign n14828 = n14271 & n14827;
  assign n14829 = po12  & n14828;
  assign n14830 = po12  & n14827;
  assign n14831 = ~n14271 & ~n14830;
  assign n14832 = ~n14829 & ~n14831;
  assign n14833 = ~po60  & ~n14816;
  assign n14834 = ~n14824 & n14833;
  assign n14835 = ~n14832 & ~n14834;
  assign n14836 = ~n14826 & ~n14835;
  assign n14837 = po61  & ~n14836;
  assign n14838 = ~n14275 & ~n14283;
  assign n14839 = n14281 & n14838;
  assign n14840 = po12  & n14839;
  assign n14841 = po12  & n14838;
  assign n14842 = ~n14281 & ~n14841;
  assign n14843 = ~n14840 & ~n14842;
  assign n14844 = ~po61  & n14836;
  assign n14845 = ~n14843 & ~n14844;
  assign n14846 = ~n14837 & ~n14845;
  assign n14847 = po62  & ~n14846;
  assign n14848 = ~n14286 & ~n14293;
  assign n14849 = n14292 & n14848;
  assign n14850 = po12  & n14849;
  assign n14851 = po12  & n14848;
  assign n14852 = ~n14292 & ~n14851;
  assign n14853 = ~n14850 & ~n14852;
  assign n14854 = ~po62  & ~n14837;
  assign n14855 = ~n14845 & n14854;
  assign n14856 = ~n14853 & ~n14855;
  assign n14857 = ~n14847 & ~n14856;
  assign n14858 = ~n14296 & ~n14304;
  assign n14859 = po12  & n14858;
  assign n14860 = ~n14302 & ~n14859;
  assign n14861 = n14302 & n14859;
  assign n14862 = ~n14860 & ~n14861;
  assign n14863 = ~n14306 & ~n14311;
  assign n14864 = po12  & n14863;
  assign n14865 = ~n14324 & ~n14864;
  assign n14866 = ~n14862 & n14865;
  assign n14867 = ~n14857 & n14866;
  assign n14868 = ~po63  & ~n14867;
  assign n14869 = ~n14311 & po12 ;
  assign n14870 = n14306 & ~n14869;
  assign n14871 = po63  & ~n14863;
  assign n14872 = ~n14870 & n14871;
  assign n14873 = n14311 & ~po12 ;
  assign n14874 = ~n14872 & ~n14873;
  assign n14875 = n14857 & n14862;
  assign n14876 = n14874 & ~n14875;
  assign po11  = n14868 | ~n14876;
  assign n14878 = pi22  & po11 ;
  assign n14879 = ~pi20  & ~pi21 ;
  assign n14880 = ~pi22  & n14879;
  assign n14881 = ~n14878 & ~n14880;
  assign n14882 = po12  & ~n14881;
  assign n14883 = n14323 & ~n14880;
  assign n14884 = ~n14324 & n14883;
  assign n14885 = ~n14317 & n14884;
  assign n14886 = ~n14878 & n14885;
  assign n14887 = ~pi22  & po11 ;
  assign n14888 = pi23  & ~n14887;
  assign n14889 = n14328 & po11 ;
  assign n14890 = ~n14888 & ~n14889;
  assign n14891 = ~n14886 & n14890;
  assign n14892 = ~n14882 & ~n14891;
  assign n14893 = po13  & ~n14892;
  assign n14894 = po12  & n14874;
  assign n14895 = ~n14875 & n14894;
  assign n14896 = ~n14868 & n14895;
  assign n14897 = ~n14889 & ~n14896;
  assign n14898 = pi24  & ~n14897;
  assign n14899 = ~pi24  & n14897;
  assign n14900 = ~n14898 & ~n14899;
  assign n14901 = ~po13  & n14892;
  assign n14902 = ~n14900 & ~n14901;
  assign n14903 = ~n14893 & ~n14902;
  assign n14904 = po14  & ~n14903;
  assign n14905 = ~n14331 & ~n14335;
  assign n14906 = ~n14339 & n14905;
  assign n14907 = po11  & n14906;
  assign n14908 = po11  & n14905;
  assign n14909 = n14339 & ~n14908;
  assign n14910 = ~n14907 & ~n14909;
  assign n14911 = ~po14  & ~n14893;
  assign n14912 = ~n14902 & n14911;
  assign n14913 = ~n14910 & ~n14912;
  assign n14914 = ~n14904 & ~n14913;
  assign n14915 = po15  & ~n14914;
  assign n14916 = ~n14342 & ~n14344;
  assign n14917 = n14351 & n14916;
  assign n14918 = po11  & n14917;
  assign n14919 = po11  & n14916;
  assign n14920 = ~n14351 & ~n14919;
  assign n14921 = ~n14918 & ~n14920;
  assign n14922 = ~po15  & n14914;
  assign n14923 = ~n14921 & ~n14922;
  assign n14924 = ~n14915 & ~n14923;
  assign n14925 = po16  & ~n14924;
  assign n14926 = ~n14354 & ~n14361;
  assign n14927 = n14360 & n14926;
  assign n14928 = po11  & n14927;
  assign n14929 = po11  & n14926;
  assign n14930 = ~n14360 & ~n14929;
  assign n14931 = ~n14928 & ~n14930;
  assign n14932 = ~po16  & ~n14915;
  assign n14933 = ~n14923 & n14932;
  assign n14934 = ~n14931 & ~n14933;
  assign n14935 = ~n14925 & ~n14934;
  assign n14936 = po17  & ~n14935;
  assign n14937 = ~n14364 & ~n14372;
  assign n14938 = n14370 & n14937;
  assign n14939 = po11  & n14938;
  assign n14940 = po11  & n14937;
  assign n14941 = ~n14370 & ~n14940;
  assign n14942 = ~n14939 & ~n14941;
  assign n14943 = ~po17  & n14935;
  assign n14944 = ~n14942 & ~n14943;
  assign n14945 = ~n14936 & ~n14944;
  assign n14946 = po18  & ~n14945;
  assign n14947 = ~n14375 & ~n14382;
  assign n14948 = n14381 & n14947;
  assign n14949 = po11  & n14948;
  assign n14950 = po11  & n14947;
  assign n14951 = ~n14381 & ~n14950;
  assign n14952 = ~n14949 & ~n14951;
  assign n14953 = ~po18  & ~n14936;
  assign n14954 = ~n14944 & n14953;
  assign n14955 = ~n14952 & ~n14954;
  assign n14956 = ~n14946 & ~n14955;
  assign n14957 = po19  & ~n14956;
  assign n14958 = ~n14385 & ~n14393;
  assign n14959 = n14391 & n14958;
  assign n14960 = po11  & n14959;
  assign n14961 = po11  & n14958;
  assign n14962 = ~n14391 & ~n14961;
  assign n14963 = ~n14960 & ~n14962;
  assign n14964 = ~po19  & n14956;
  assign n14965 = ~n14963 & ~n14964;
  assign n14966 = ~n14957 & ~n14965;
  assign n14967 = po20  & ~n14966;
  assign n14968 = ~n14396 & ~n14403;
  assign n14969 = n14402 & n14968;
  assign n14970 = po11  & n14969;
  assign n14971 = po11  & n14968;
  assign n14972 = ~n14402 & ~n14971;
  assign n14973 = ~n14970 & ~n14972;
  assign n14974 = ~po20  & ~n14957;
  assign n14975 = ~n14965 & n14974;
  assign n14976 = ~n14973 & ~n14975;
  assign n14977 = ~n14967 & ~n14976;
  assign n14978 = po21  & ~n14977;
  assign n14979 = ~n14406 & ~n14414;
  assign n14980 = n14412 & n14979;
  assign n14981 = po11  & n14980;
  assign n14982 = po11  & n14979;
  assign n14983 = ~n14412 & ~n14982;
  assign n14984 = ~n14981 & ~n14983;
  assign n14985 = ~po21  & n14977;
  assign n14986 = ~n14984 & ~n14985;
  assign n14987 = ~n14978 & ~n14986;
  assign n14988 = po22  & ~n14987;
  assign n14989 = ~n14417 & ~n14424;
  assign n14990 = n14423 & n14989;
  assign n14991 = po11  & n14990;
  assign n14992 = po11  & n14989;
  assign n14993 = ~n14423 & ~n14992;
  assign n14994 = ~n14991 & ~n14993;
  assign n14995 = ~po22  & ~n14978;
  assign n14996 = ~n14986 & n14995;
  assign n14997 = ~n14994 & ~n14996;
  assign n14998 = ~n14988 & ~n14997;
  assign n14999 = po23  & ~n14998;
  assign n15000 = ~n14427 & ~n14435;
  assign n15001 = n14433 & n15000;
  assign n15002 = po11  & n15001;
  assign n15003 = po11  & n15000;
  assign n15004 = ~n14433 & ~n15003;
  assign n15005 = ~n15002 & ~n15004;
  assign n15006 = ~po23  & n14998;
  assign n15007 = ~n15005 & ~n15006;
  assign n15008 = ~n14999 & ~n15007;
  assign n15009 = po24  & ~n15008;
  assign n15010 = ~n14438 & ~n14445;
  assign n15011 = n14444 & n15010;
  assign n15012 = po11  & n15011;
  assign n15013 = po11  & n15010;
  assign n15014 = ~n14444 & ~n15013;
  assign n15015 = ~n15012 & ~n15014;
  assign n15016 = ~po24  & ~n14999;
  assign n15017 = ~n15007 & n15016;
  assign n15018 = ~n15015 & ~n15017;
  assign n15019 = ~n15009 & ~n15018;
  assign n15020 = po25  & ~n15019;
  assign n15021 = ~n14448 & ~n14456;
  assign n15022 = n14454 & n15021;
  assign n15023 = po11  & n15022;
  assign n15024 = po11  & n15021;
  assign n15025 = ~n14454 & ~n15024;
  assign n15026 = ~n15023 & ~n15025;
  assign n15027 = ~po25  & n15019;
  assign n15028 = ~n15026 & ~n15027;
  assign n15029 = ~n15020 & ~n15028;
  assign n15030 = po26  & ~n15029;
  assign n15031 = ~n14459 & ~n14466;
  assign n15032 = n14465 & n15031;
  assign n15033 = po11  & n15032;
  assign n15034 = po11  & n15031;
  assign n15035 = ~n14465 & ~n15034;
  assign n15036 = ~n15033 & ~n15035;
  assign n15037 = ~po26  & ~n15020;
  assign n15038 = ~n15028 & n15037;
  assign n15039 = ~n15036 & ~n15038;
  assign n15040 = ~n15030 & ~n15039;
  assign n15041 = po27  & ~n15040;
  assign n15042 = ~n14469 & ~n14477;
  assign n15043 = n14475 & n15042;
  assign n15044 = po11  & n15043;
  assign n15045 = po11  & n15042;
  assign n15046 = ~n14475 & ~n15045;
  assign n15047 = ~n15044 & ~n15046;
  assign n15048 = ~po27  & n15040;
  assign n15049 = ~n15047 & ~n15048;
  assign n15050 = ~n15041 & ~n15049;
  assign n15051 = po28  & ~n15050;
  assign n15052 = ~n14480 & ~n14487;
  assign n15053 = n14486 & n15052;
  assign n15054 = po11  & n15053;
  assign n15055 = po11  & n15052;
  assign n15056 = ~n14486 & ~n15055;
  assign n15057 = ~n15054 & ~n15056;
  assign n15058 = ~po28  & ~n15041;
  assign n15059 = ~n15049 & n15058;
  assign n15060 = ~n15057 & ~n15059;
  assign n15061 = ~n15051 & ~n15060;
  assign n15062 = po29  & ~n15061;
  assign n15063 = ~n14490 & ~n14498;
  assign n15064 = n14496 & n15063;
  assign n15065 = po11  & n15064;
  assign n15066 = po11  & n15063;
  assign n15067 = ~n14496 & ~n15066;
  assign n15068 = ~n15065 & ~n15067;
  assign n15069 = ~po29  & n15061;
  assign n15070 = ~n15068 & ~n15069;
  assign n15071 = ~n15062 & ~n15070;
  assign n15072 = po30  & ~n15071;
  assign n15073 = ~n14501 & ~n14508;
  assign n15074 = n14507 & n15073;
  assign n15075 = po11  & n15074;
  assign n15076 = po11  & n15073;
  assign n15077 = ~n14507 & ~n15076;
  assign n15078 = ~n15075 & ~n15077;
  assign n15079 = ~po30  & ~n15062;
  assign n15080 = ~n15070 & n15079;
  assign n15081 = ~n15078 & ~n15080;
  assign n15082 = ~n15072 & ~n15081;
  assign n15083 = po31  & ~n15082;
  assign n15084 = ~n14511 & ~n14519;
  assign n15085 = n14517 & n15084;
  assign n15086 = po11  & n15085;
  assign n15087 = po11  & n15084;
  assign n15088 = ~n14517 & ~n15087;
  assign n15089 = ~n15086 & ~n15088;
  assign n15090 = ~po31  & n15082;
  assign n15091 = ~n15089 & ~n15090;
  assign n15092 = ~n15083 & ~n15091;
  assign n15093 = po32  & ~n15092;
  assign n15094 = ~n14522 & ~n14529;
  assign n15095 = n14528 & n15094;
  assign n15096 = po11  & n15095;
  assign n15097 = po11  & n15094;
  assign n15098 = ~n14528 & ~n15097;
  assign n15099 = ~n15096 & ~n15098;
  assign n15100 = ~po32  & ~n15083;
  assign n15101 = ~n15091 & n15100;
  assign n15102 = ~n15099 & ~n15101;
  assign n15103 = ~n15093 & ~n15102;
  assign n15104 = po33  & ~n15103;
  assign n15105 = ~n14532 & ~n14540;
  assign n15106 = n14538 & n15105;
  assign n15107 = po11  & n15106;
  assign n15108 = po11  & n15105;
  assign n15109 = ~n14538 & ~n15108;
  assign n15110 = ~n15107 & ~n15109;
  assign n15111 = ~po33  & n15103;
  assign n15112 = ~n15110 & ~n15111;
  assign n15113 = ~n15104 & ~n15112;
  assign n15114 = po34  & ~n15113;
  assign n15115 = ~n14543 & ~n14550;
  assign n15116 = n14549 & n15115;
  assign n15117 = po11  & n15116;
  assign n15118 = po11  & n15115;
  assign n15119 = ~n14549 & ~n15118;
  assign n15120 = ~n15117 & ~n15119;
  assign n15121 = ~po34  & ~n15104;
  assign n15122 = ~n15112 & n15121;
  assign n15123 = ~n15120 & ~n15122;
  assign n15124 = ~n15114 & ~n15123;
  assign n15125 = po35  & ~n15124;
  assign n15126 = ~n14553 & ~n14561;
  assign n15127 = n14559 & n15126;
  assign n15128 = po11  & n15127;
  assign n15129 = po11  & n15126;
  assign n15130 = ~n14559 & ~n15129;
  assign n15131 = ~n15128 & ~n15130;
  assign n15132 = ~po35  & n15124;
  assign n15133 = ~n15131 & ~n15132;
  assign n15134 = ~n15125 & ~n15133;
  assign n15135 = po36  & ~n15134;
  assign n15136 = ~n14564 & ~n14571;
  assign n15137 = n14570 & n15136;
  assign n15138 = po11  & n15137;
  assign n15139 = po11  & n15136;
  assign n15140 = ~n14570 & ~n15139;
  assign n15141 = ~n15138 & ~n15140;
  assign n15142 = ~po36  & ~n15125;
  assign n15143 = ~n15133 & n15142;
  assign n15144 = ~n15141 & ~n15143;
  assign n15145 = ~n15135 & ~n15144;
  assign n15146 = po37  & ~n15145;
  assign n15147 = ~n14574 & ~n14582;
  assign n15148 = n14580 & n15147;
  assign n15149 = po11  & n15148;
  assign n15150 = po11  & n15147;
  assign n15151 = ~n14580 & ~n15150;
  assign n15152 = ~n15149 & ~n15151;
  assign n15153 = ~po37  & n15145;
  assign n15154 = ~n15152 & ~n15153;
  assign n15155 = ~n15146 & ~n15154;
  assign n15156 = po38  & ~n15155;
  assign n15157 = ~n14585 & ~n14592;
  assign n15158 = n14591 & n15157;
  assign n15159 = po11  & n15158;
  assign n15160 = po11  & n15157;
  assign n15161 = ~n14591 & ~n15160;
  assign n15162 = ~n15159 & ~n15161;
  assign n15163 = ~po38  & ~n15146;
  assign n15164 = ~n15154 & n15163;
  assign n15165 = ~n15162 & ~n15164;
  assign n15166 = ~n15156 & ~n15165;
  assign n15167 = po39  & ~n15166;
  assign n15168 = ~n14595 & ~n14603;
  assign n15169 = n14601 & n15168;
  assign n15170 = po11  & n15169;
  assign n15171 = po11  & n15168;
  assign n15172 = ~n14601 & ~n15171;
  assign n15173 = ~n15170 & ~n15172;
  assign n15174 = ~po39  & n15166;
  assign n15175 = ~n15173 & ~n15174;
  assign n15176 = ~n15167 & ~n15175;
  assign n15177 = po40  & ~n15176;
  assign n15178 = ~n14606 & ~n14613;
  assign n15179 = n14612 & n15178;
  assign n15180 = po11  & n15179;
  assign n15181 = po11  & n15178;
  assign n15182 = ~n14612 & ~n15181;
  assign n15183 = ~n15180 & ~n15182;
  assign n15184 = ~po40  & ~n15167;
  assign n15185 = ~n15175 & n15184;
  assign n15186 = ~n15183 & ~n15185;
  assign n15187 = ~n15177 & ~n15186;
  assign n15188 = po41  & ~n15187;
  assign n15189 = ~n14616 & ~n14624;
  assign n15190 = n14622 & n15189;
  assign n15191 = po11  & n15190;
  assign n15192 = po11  & n15189;
  assign n15193 = ~n14622 & ~n15192;
  assign n15194 = ~n15191 & ~n15193;
  assign n15195 = ~po41  & n15187;
  assign n15196 = ~n15194 & ~n15195;
  assign n15197 = ~n15188 & ~n15196;
  assign n15198 = po42  & ~n15197;
  assign n15199 = ~n14627 & ~n14634;
  assign n15200 = n14633 & n15199;
  assign n15201 = po11  & n15200;
  assign n15202 = po11  & n15199;
  assign n15203 = ~n14633 & ~n15202;
  assign n15204 = ~n15201 & ~n15203;
  assign n15205 = ~po42  & ~n15188;
  assign n15206 = ~n15196 & n15205;
  assign n15207 = ~n15204 & ~n15206;
  assign n15208 = ~n15198 & ~n15207;
  assign n15209 = po43  & ~n15208;
  assign n15210 = ~n14637 & ~n14645;
  assign n15211 = n14643 & n15210;
  assign n15212 = po11  & n15211;
  assign n15213 = po11  & n15210;
  assign n15214 = ~n14643 & ~n15213;
  assign n15215 = ~n15212 & ~n15214;
  assign n15216 = ~po43  & n15208;
  assign n15217 = ~n15215 & ~n15216;
  assign n15218 = ~n15209 & ~n15217;
  assign n15219 = po44  & ~n15218;
  assign n15220 = ~n14648 & ~n14655;
  assign n15221 = n14654 & n15220;
  assign n15222 = po11  & n15221;
  assign n15223 = po11  & n15220;
  assign n15224 = ~n14654 & ~n15223;
  assign n15225 = ~n15222 & ~n15224;
  assign n15226 = ~po44  & ~n15209;
  assign n15227 = ~n15217 & n15226;
  assign n15228 = ~n15225 & ~n15227;
  assign n15229 = ~n15219 & ~n15228;
  assign n15230 = po45  & ~n15229;
  assign n15231 = ~n14658 & ~n14666;
  assign n15232 = n14664 & n15231;
  assign n15233 = po11  & n15232;
  assign n15234 = po11  & n15231;
  assign n15235 = ~n14664 & ~n15234;
  assign n15236 = ~n15233 & ~n15235;
  assign n15237 = ~po45  & n15229;
  assign n15238 = ~n15236 & ~n15237;
  assign n15239 = ~n15230 & ~n15238;
  assign n15240 = po46  & ~n15239;
  assign n15241 = ~n14669 & ~n14676;
  assign n15242 = n14675 & n15241;
  assign n15243 = po11  & n15242;
  assign n15244 = po11  & n15241;
  assign n15245 = ~n14675 & ~n15244;
  assign n15246 = ~n15243 & ~n15245;
  assign n15247 = ~po46  & ~n15230;
  assign n15248 = ~n15238 & n15247;
  assign n15249 = ~n15246 & ~n15248;
  assign n15250 = ~n15240 & ~n15249;
  assign n15251 = po47  & ~n15250;
  assign n15252 = ~n14679 & ~n14687;
  assign n15253 = n14685 & n15252;
  assign n15254 = po11  & n15253;
  assign n15255 = po11  & n15252;
  assign n15256 = ~n14685 & ~n15255;
  assign n15257 = ~n15254 & ~n15256;
  assign n15258 = ~po47  & n15250;
  assign n15259 = ~n15257 & ~n15258;
  assign n15260 = ~n15251 & ~n15259;
  assign n15261 = po48  & ~n15260;
  assign n15262 = ~n14690 & ~n14697;
  assign n15263 = n14696 & n15262;
  assign n15264 = po11  & n15263;
  assign n15265 = po11  & n15262;
  assign n15266 = ~n14696 & ~n15265;
  assign n15267 = ~n15264 & ~n15266;
  assign n15268 = ~po48  & ~n15251;
  assign n15269 = ~n15259 & n15268;
  assign n15270 = ~n15267 & ~n15269;
  assign n15271 = ~n15261 & ~n15270;
  assign n15272 = po49  & ~n15271;
  assign n15273 = ~n14700 & ~n14708;
  assign n15274 = n14706 & n15273;
  assign n15275 = po11  & n15274;
  assign n15276 = po11  & n15273;
  assign n15277 = ~n14706 & ~n15276;
  assign n15278 = ~n15275 & ~n15277;
  assign n15279 = ~po49  & n15271;
  assign n15280 = ~n15278 & ~n15279;
  assign n15281 = ~n15272 & ~n15280;
  assign n15282 = po50  & ~n15281;
  assign n15283 = ~n14711 & ~n14718;
  assign n15284 = n14717 & n15283;
  assign n15285 = po11  & n15284;
  assign n15286 = po11  & n15283;
  assign n15287 = ~n14717 & ~n15286;
  assign n15288 = ~n15285 & ~n15287;
  assign n15289 = ~po50  & ~n15272;
  assign n15290 = ~n15280 & n15289;
  assign n15291 = ~n15288 & ~n15290;
  assign n15292 = ~n15282 & ~n15291;
  assign n15293 = po51  & ~n15292;
  assign n15294 = ~n14721 & ~n14729;
  assign n15295 = n14727 & n15294;
  assign n15296 = po11  & n15295;
  assign n15297 = po11  & n15294;
  assign n15298 = ~n14727 & ~n15297;
  assign n15299 = ~n15296 & ~n15298;
  assign n15300 = ~po51  & n15292;
  assign n15301 = ~n15299 & ~n15300;
  assign n15302 = ~n15293 & ~n15301;
  assign n15303 = po52  & ~n15302;
  assign n15304 = ~n14732 & ~n14739;
  assign n15305 = n14738 & n15304;
  assign n15306 = po11  & n15305;
  assign n15307 = po11  & n15304;
  assign n15308 = ~n14738 & ~n15307;
  assign n15309 = ~n15306 & ~n15308;
  assign n15310 = ~po52  & ~n15293;
  assign n15311 = ~n15301 & n15310;
  assign n15312 = ~n15309 & ~n15311;
  assign n15313 = ~n15303 & ~n15312;
  assign n15314 = po53  & ~n15313;
  assign n15315 = ~n14742 & ~n14750;
  assign n15316 = n14748 & n15315;
  assign n15317 = po11  & n15316;
  assign n15318 = po11  & n15315;
  assign n15319 = ~n14748 & ~n15318;
  assign n15320 = ~n15317 & ~n15319;
  assign n15321 = ~po53  & n15313;
  assign n15322 = ~n15320 & ~n15321;
  assign n15323 = ~n15314 & ~n15322;
  assign n15324 = po54  & ~n15323;
  assign n15325 = ~po54  & ~n15314;
  assign n15326 = ~n15322 & n15325;
  assign n15327 = ~n14753 & ~n14760;
  assign n15328 = n14759 & n15327;
  assign n15329 = po11  & n15328;
  assign n15330 = po11  & n15327;
  assign n15331 = ~n14759 & ~n15330;
  assign n15332 = ~n15329 & ~n15331;
  assign n15333 = ~n15326 & ~n15332;
  assign n15334 = ~n15324 & ~n15333;
  assign n15335 = po55  & ~n15334;
  assign n15336 = ~n14763 & ~n14771;
  assign n15337 = n14769 & n15336;
  assign n15338 = po11  & n15337;
  assign n15339 = po11  & n15336;
  assign n15340 = ~n14769 & ~n15339;
  assign n15341 = ~n15338 & ~n15340;
  assign n15342 = ~po55  & n15334;
  assign n15343 = ~n15341 & ~n15342;
  assign n15344 = ~n15335 & ~n15343;
  assign n15345 = po56  & ~n15344;
  assign n15346 = ~n14774 & ~n14781;
  assign n15347 = n14780 & n15346;
  assign n15348 = po11  & n15347;
  assign n15349 = po11  & n15346;
  assign n15350 = ~n14780 & ~n15349;
  assign n15351 = ~n15348 & ~n15350;
  assign n15352 = ~po56  & ~n15335;
  assign n15353 = ~n15343 & n15352;
  assign n15354 = ~n15351 & ~n15353;
  assign n15355 = ~n15345 & ~n15354;
  assign n15356 = po57  & ~n15355;
  assign n15357 = ~n14784 & ~n14792;
  assign n15358 = n14790 & n15357;
  assign n15359 = po11  & n15358;
  assign n15360 = po11  & n15357;
  assign n15361 = ~n14790 & ~n15360;
  assign n15362 = ~n15359 & ~n15361;
  assign n15363 = ~po57  & n15355;
  assign n15364 = ~n15362 & ~n15363;
  assign n15365 = ~n15356 & ~n15364;
  assign n15366 = po58  & ~n15365;
  assign n15367 = ~n14795 & ~n14802;
  assign n15368 = n14801 & n15367;
  assign n15369 = po11  & n15368;
  assign n15370 = po11  & n15367;
  assign n15371 = ~n14801 & ~n15370;
  assign n15372 = ~n15369 & ~n15371;
  assign n15373 = ~po58  & ~n15356;
  assign n15374 = ~n15364 & n15373;
  assign n15375 = ~n15372 & ~n15374;
  assign n15376 = ~n15366 & ~n15375;
  assign n15377 = po59  & ~n15376;
  assign n15378 = ~n14805 & ~n14813;
  assign n15379 = n14811 & n15378;
  assign n15380 = po11  & n15379;
  assign n15381 = po11  & n15378;
  assign n15382 = ~n14811 & ~n15381;
  assign n15383 = ~n15380 & ~n15382;
  assign n15384 = ~po59  & n15376;
  assign n15385 = ~n15383 & ~n15384;
  assign n15386 = ~n15377 & ~n15385;
  assign n15387 = po60  & ~n15386;
  assign n15388 = ~n14816 & ~n14823;
  assign n15389 = n14822 & n15388;
  assign n15390 = po11  & n15389;
  assign n15391 = po11  & n15388;
  assign n15392 = ~n14822 & ~n15391;
  assign n15393 = ~n15390 & ~n15392;
  assign n15394 = ~po60  & ~n15377;
  assign n15395 = ~n15385 & n15394;
  assign n15396 = ~n15393 & ~n15395;
  assign n15397 = ~n15387 & ~n15396;
  assign n15398 = po61  & ~n15397;
  assign n15399 = ~n14826 & ~n14834;
  assign n15400 = n14832 & n15399;
  assign n15401 = po11  & n15400;
  assign n15402 = po11  & n15399;
  assign n15403 = ~n14832 & ~n15402;
  assign n15404 = ~n15401 & ~n15403;
  assign n15405 = ~po61  & n15397;
  assign n15406 = ~n15404 & ~n15405;
  assign n15407 = ~n15398 & ~n15406;
  assign n15408 = po62  & ~n15407;
  assign n15409 = ~n14837 & ~n14844;
  assign n15410 = n14843 & n15409;
  assign n15411 = po11  & n15410;
  assign n15412 = po11  & n15409;
  assign n15413 = ~n14843 & ~n15412;
  assign n15414 = ~n15411 & ~n15413;
  assign n15415 = ~po62  & ~n15398;
  assign n15416 = ~n15406 & n15415;
  assign n15417 = ~n15414 & ~n15416;
  assign n15418 = ~n15408 & ~n15417;
  assign n15419 = ~n14847 & ~n14855;
  assign n15420 = po11  & n15419;
  assign n15421 = ~n14853 & ~n15420;
  assign n15422 = n14853 & n15420;
  assign n15423 = ~n15421 & ~n15422;
  assign n15424 = ~n14857 & ~n14862;
  assign n15425 = po11  & n15424;
  assign n15426 = ~n14875 & ~n15425;
  assign n15427 = ~n15423 & n15426;
  assign n15428 = ~n15418 & n15427;
  assign n15429 = ~po63  & ~n15428;
  assign n15430 = ~n14862 & po11 ;
  assign n15431 = n14857 & ~n15430;
  assign n15432 = po63  & ~n15424;
  assign n15433 = ~n15431 & n15432;
  assign n15434 = n14862 & ~po11 ;
  assign n15435 = ~n15433 & ~n15434;
  assign n15436 = n15418 & n15423;
  assign n15437 = n15435 & ~n15436;
  assign po10  = n15429 | ~n15437;
  assign n15439 = pi20  & po10 ;
  assign n15440 = ~pi18  & ~pi19 ;
  assign n15441 = ~pi20  & n15440;
  assign n15442 = ~n15439 & ~n15441;
  assign n15443 = po11  & ~n15442;
  assign n15444 = n14874 & ~n15441;
  assign n15445 = ~n14875 & n15444;
  assign n15446 = ~n14868 & n15445;
  assign n15447 = ~n15439 & n15446;
  assign n15448 = ~pi20  & po10 ;
  assign n15449 = pi21  & ~n15448;
  assign n15450 = n14879 & po10 ;
  assign n15451 = ~n15449 & ~n15450;
  assign n15452 = ~n15447 & n15451;
  assign n15453 = ~n15443 & ~n15452;
  assign n15454 = po12  & ~n15453;
  assign n15455 = ~po12  & ~n15443;
  assign n15456 = ~n15452 & n15455;
  assign n15457 = po11  & n15435;
  assign n15458 = ~n15436 & n15457;
  assign n15459 = ~n15429 & n15458;
  assign n15460 = ~n15450 & ~n15459;
  assign n15461 = pi22  & ~n15460;
  assign n15462 = ~pi22  & n15460;
  assign n15463 = ~n15461 & ~n15462;
  assign n15464 = ~n15456 & ~n15463;
  assign n15465 = ~n15454 & ~n15464;
  assign n15466 = po13  & ~n15465;
  assign n15467 = ~n14882 & ~n14886;
  assign n15468 = ~n14890 & n15467;
  assign n15469 = po10  & n15468;
  assign n15470 = po10  & n15467;
  assign n15471 = n14890 & ~n15470;
  assign n15472 = ~n15469 & ~n15471;
  assign n15473 = ~po13  & n15465;
  assign n15474 = ~n15472 & ~n15473;
  assign n15475 = ~n15466 & ~n15474;
  assign n15476 = po14  & ~n15475;
  assign n15477 = ~n14893 & ~n14901;
  assign n15478 = n14900 & n15477;
  assign n15479 = po10  & n15478;
  assign n15480 = po10  & n15477;
  assign n15481 = ~n14900 & ~n15480;
  assign n15482 = ~n15479 & ~n15481;
  assign n15483 = ~po14  & ~n15466;
  assign n15484 = ~n15474 & n15483;
  assign n15485 = ~n15482 & ~n15484;
  assign n15486 = ~n15476 & ~n15485;
  assign n15487 = po15  & ~n15486;
  assign n15488 = ~n14904 & ~n14912;
  assign n15489 = n14910 & n15488;
  assign n15490 = po10  & n15489;
  assign n15491 = po10  & n15488;
  assign n15492 = ~n14910 & ~n15491;
  assign n15493 = ~n15490 & ~n15492;
  assign n15494 = ~po15  & n15486;
  assign n15495 = ~n15493 & ~n15494;
  assign n15496 = ~n15487 & ~n15495;
  assign n15497 = po16  & ~n15496;
  assign n15498 = ~n14915 & ~n14922;
  assign n15499 = n14921 & n15498;
  assign n15500 = po10  & n15499;
  assign n15501 = po10  & n15498;
  assign n15502 = ~n14921 & ~n15501;
  assign n15503 = ~n15500 & ~n15502;
  assign n15504 = ~po16  & ~n15487;
  assign n15505 = ~n15495 & n15504;
  assign n15506 = ~n15503 & ~n15505;
  assign n15507 = ~n15497 & ~n15506;
  assign n15508 = po17  & ~n15507;
  assign n15509 = ~n14925 & ~n14933;
  assign n15510 = n14931 & n15509;
  assign n15511 = po10  & n15510;
  assign n15512 = po10  & n15509;
  assign n15513 = ~n14931 & ~n15512;
  assign n15514 = ~n15511 & ~n15513;
  assign n15515 = ~po17  & n15507;
  assign n15516 = ~n15514 & ~n15515;
  assign n15517 = ~n15508 & ~n15516;
  assign n15518 = po18  & ~n15517;
  assign n15519 = ~n14936 & ~n14943;
  assign n15520 = n14942 & n15519;
  assign n15521 = po10  & n15520;
  assign n15522 = po10  & n15519;
  assign n15523 = ~n14942 & ~n15522;
  assign n15524 = ~n15521 & ~n15523;
  assign n15525 = ~po18  & ~n15508;
  assign n15526 = ~n15516 & n15525;
  assign n15527 = ~n15524 & ~n15526;
  assign n15528 = ~n15518 & ~n15527;
  assign n15529 = po19  & ~n15528;
  assign n15530 = ~n14946 & ~n14954;
  assign n15531 = n14952 & n15530;
  assign n15532 = po10  & n15531;
  assign n15533 = po10  & n15530;
  assign n15534 = ~n14952 & ~n15533;
  assign n15535 = ~n15532 & ~n15534;
  assign n15536 = ~po19  & n15528;
  assign n15537 = ~n15535 & ~n15536;
  assign n15538 = ~n15529 & ~n15537;
  assign n15539 = po20  & ~n15538;
  assign n15540 = ~n14957 & ~n14964;
  assign n15541 = n14963 & n15540;
  assign n15542 = po10  & n15541;
  assign n15543 = po10  & n15540;
  assign n15544 = ~n14963 & ~n15543;
  assign n15545 = ~n15542 & ~n15544;
  assign n15546 = ~po20  & ~n15529;
  assign n15547 = ~n15537 & n15546;
  assign n15548 = ~n15545 & ~n15547;
  assign n15549 = ~n15539 & ~n15548;
  assign n15550 = po21  & ~n15549;
  assign n15551 = ~n14967 & ~n14975;
  assign n15552 = n14973 & n15551;
  assign n15553 = po10  & n15552;
  assign n15554 = po10  & n15551;
  assign n15555 = ~n14973 & ~n15554;
  assign n15556 = ~n15553 & ~n15555;
  assign n15557 = ~po21  & n15549;
  assign n15558 = ~n15556 & ~n15557;
  assign n15559 = ~n15550 & ~n15558;
  assign n15560 = po22  & ~n15559;
  assign n15561 = ~n14978 & ~n14985;
  assign n15562 = n14984 & n15561;
  assign n15563 = po10  & n15562;
  assign n15564 = po10  & n15561;
  assign n15565 = ~n14984 & ~n15564;
  assign n15566 = ~n15563 & ~n15565;
  assign n15567 = ~po22  & ~n15550;
  assign n15568 = ~n15558 & n15567;
  assign n15569 = ~n15566 & ~n15568;
  assign n15570 = ~n15560 & ~n15569;
  assign n15571 = po23  & ~n15570;
  assign n15572 = ~n14988 & ~n14996;
  assign n15573 = n14994 & n15572;
  assign n15574 = po10  & n15573;
  assign n15575 = po10  & n15572;
  assign n15576 = ~n14994 & ~n15575;
  assign n15577 = ~n15574 & ~n15576;
  assign n15578 = ~po23  & n15570;
  assign n15579 = ~n15577 & ~n15578;
  assign n15580 = ~n15571 & ~n15579;
  assign n15581 = po24  & ~n15580;
  assign n15582 = ~n14999 & ~n15006;
  assign n15583 = n15005 & n15582;
  assign n15584 = po10  & n15583;
  assign n15585 = po10  & n15582;
  assign n15586 = ~n15005 & ~n15585;
  assign n15587 = ~n15584 & ~n15586;
  assign n15588 = ~po24  & ~n15571;
  assign n15589 = ~n15579 & n15588;
  assign n15590 = ~n15587 & ~n15589;
  assign n15591 = ~n15581 & ~n15590;
  assign n15592 = po25  & ~n15591;
  assign n15593 = ~n15009 & ~n15017;
  assign n15594 = n15015 & n15593;
  assign n15595 = po10  & n15594;
  assign n15596 = po10  & n15593;
  assign n15597 = ~n15015 & ~n15596;
  assign n15598 = ~n15595 & ~n15597;
  assign n15599 = ~po25  & n15591;
  assign n15600 = ~n15598 & ~n15599;
  assign n15601 = ~n15592 & ~n15600;
  assign n15602 = po26  & ~n15601;
  assign n15603 = ~n15020 & ~n15027;
  assign n15604 = n15026 & n15603;
  assign n15605 = po10  & n15604;
  assign n15606 = po10  & n15603;
  assign n15607 = ~n15026 & ~n15606;
  assign n15608 = ~n15605 & ~n15607;
  assign n15609 = ~po26  & ~n15592;
  assign n15610 = ~n15600 & n15609;
  assign n15611 = ~n15608 & ~n15610;
  assign n15612 = ~n15602 & ~n15611;
  assign n15613 = po27  & ~n15612;
  assign n15614 = ~n15030 & ~n15038;
  assign n15615 = n15036 & n15614;
  assign n15616 = po10  & n15615;
  assign n15617 = po10  & n15614;
  assign n15618 = ~n15036 & ~n15617;
  assign n15619 = ~n15616 & ~n15618;
  assign n15620 = ~po27  & n15612;
  assign n15621 = ~n15619 & ~n15620;
  assign n15622 = ~n15613 & ~n15621;
  assign n15623 = po28  & ~n15622;
  assign n15624 = ~n15041 & ~n15048;
  assign n15625 = n15047 & n15624;
  assign n15626 = po10  & n15625;
  assign n15627 = po10  & n15624;
  assign n15628 = ~n15047 & ~n15627;
  assign n15629 = ~n15626 & ~n15628;
  assign n15630 = ~po28  & ~n15613;
  assign n15631 = ~n15621 & n15630;
  assign n15632 = ~n15629 & ~n15631;
  assign n15633 = ~n15623 & ~n15632;
  assign n15634 = po29  & ~n15633;
  assign n15635 = ~n15051 & ~n15059;
  assign n15636 = n15057 & n15635;
  assign n15637 = po10  & n15636;
  assign n15638 = po10  & n15635;
  assign n15639 = ~n15057 & ~n15638;
  assign n15640 = ~n15637 & ~n15639;
  assign n15641 = ~po29  & n15633;
  assign n15642 = ~n15640 & ~n15641;
  assign n15643 = ~n15634 & ~n15642;
  assign n15644 = po30  & ~n15643;
  assign n15645 = ~n15062 & ~n15069;
  assign n15646 = n15068 & n15645;
  assign n15647 = po10  & n15646;
  assign n15648 = po10  & n15645;
  assign n15649 = ~n15068 & ~n15648;
  assign n15650 = ~n15647 & ~n15649;
  assign n15651 = ~po30  & ~n15634;
  assign n15652 = ~n15642 & n15651;
  assign n15653 = ~n15650 & ~n15652;
  assign n15654 = ~n15644 & ~n15653;
  assign n15655 = po31  & ~n15654;
  assign n15656 = ~n15072 & ~n15080;
  assign n15657 = n15078 & n15656;
  assign n15658 = po10  & n15657;
  assign n15659 = po10  & n15656;
  assign n15660 = ~n15078 & ~n15659;
  assign n15661 = ~n15658 & ~n15660;
  assign n15662 = ~po31  & n15654;
  assign n15663 = ~n15661 & ~n15662;
  assign n15664 = ~n15655 & ~n15663;
  assign n15665 = po32  & ~n15664;
  assign n15666 = ~n15083 & ~n15090;
  assign n15667 = n15089 & n15666;
  assign n15668 = po10  & n15667;
  assign n15669 = po10  & n15666;
  assign n15670 = ~n15089 & ~n15669;
  assign n15671 = ~n15668 & ~n15670;
  assign n15672 = ~po32  & ~n15655;
  assign n15673 = ~n15663 & n15672;
  assign n15674 = ~n15671 & ~n15673;
  assign n15675 = ~n15665 & ~n15674;
  assign n15676 = po33  & ~n15675;
  assign n15677 = ~n15093 & ~n15101;
  assign n15678 = n15099 & n15677;
  assign n15679 = po10  & n15678;
  assign n15680 = po10  & n15677;
  assign n15681 = ~n15099 & ~n15680;
  assign n15682 = ~n15679 & ~n15681;
  assign n15683 = ~po33  & n15675;
  assign n15684 = ~n15682 & ~n15683;
  assign n15685 = ~n15676 & ~n15684;
  assign n15686 = po34  & ~n15685;
  assign n15687 = ~n15104 & ~n15111;
  assign n15688 = n15110 & n15687;
  assign n15689 = po10  & n15688;
  assign n15690 = po10  & n15687;
  assign n15691 = ~n15110 & ~n15690;
  assign n15692 = ~n15689 & ~n15691;
  assign n15693 = ~po34  & ~n15676;
  assign n15694 = ~n15684 & n15693;
  assign n15695 = ~n15692 & ~n15694;
  assign n15696 = ~n15686 & ~n15695;
  assign n15697 = po35  & ~n15696;
  assign n15698 = ~n15114 & ~n15122;
  assign n15699 = n15120 & n15698;
  assign n15700 = po10  & n15699;
  assign n15701 = po10  & n15698;
  assign n15702 = ~n15120 & ~n15701;
  assign n15703 = ~n15700 & ~n15702;
  assign n15704 = ~po35  & n15696;
  assign n15705 = ~n15703 & ~n15704;
  assign n15706 = ~n15697 & ~n15705;
  assign n15707 = po36  & ~n15706;
  assign n15708 = ~n15125 & ~n15132;
  assign n15709 = n15131 & n15708;
  assign n15710 = po10  & n15709;
  assign n15711 = po10  & n15708;
  assign n15712 = ~n15131 & ~n15711;
  assign n15713 = ~n15710 & ~n15712;
  assign n15714 = ~po36  & ~n15697;
  assign n15715 = ~n15705 & n15714;
  assign n15716 = ~n15713 & ~n15715;
  assign n15717 = ~n15707 & ~n15716;
  assign n15718 = po37  & ~n15717;
  assign n15719 = ~n15135 & ~n15143;
  assign n15720 = n15141 & n15719;
  assign n15721 = po10  & n15720;
  assign n15722 = po10  & n15719;
  assign n15723 = ~n15141 & ~n15722;
  assign n15724 = ~n15721 & ~n15723;
  assign n15725 = ~po37  & n15717;
  assign n15726 = ~n15724 & ~n15725;
  assign n15727 = ~n15718 & ~n15726;
  assign n15728 = po38  & ~n15727;
  assign n15729 = ~n15146 & ~n15153;
  assign n15730 = n15152 & n15729;
  assign n15731 = po10  & n15730;
  assign n15732 = po10  & n15729;
  assign n15733 = ~n15152 & ~n15732;
  assign n15734 = ~n15731 & ~n15733;
  assign n15735 = ~po38  & ~n15718;
  assign n15736 = ~n15726 & n15735;
  assign n15737 = ~n15734 & ~n15736;
  assign n15738 = ~n15728 & ~n15737;
  assign n15739 = po39  & ~n15738;
  assign n15740 = ~n15156 & ~n15164;
  assign n15741 = n15162 & n15740;
  assign n15742 = po10  & n15741;
  assign n15743 = po10  & n15740;
  assign n15744 = ~n15162 & ~n15743;
  assign n15745 = ~n15742 & ~n15744;
  assign n15746 = ~po39  & n15738;
  assign n15747 = ~n15745 & ~n15746;
  assign n15748 = ~n15739 & ~n15747;
  assign n15749 = po40  & ~n15748;
  assign n15750 = ~n15167 & ~n15174;
  assign n15751 = n15173 & n15750;
  assign n15752 = po10  & n15751;
  assign n15753 = po10  & n15750;
  assign n15754 = ~n15173 & ~n15753;
  assign n15755 = ~n15752 & ~n15754;
  assign n15756 = ~po40  & ~n15739;
  assign n15757 = ~n15747 & n15756;
  assign n15758 = ~n15755 & ~n15757;
  assign n15759 = ~n15749 & ~n15758;
  assign n15760 = po41  & ~n15759;
  assign n15761 = ~n15177 & ~n15185;
  assign n15762 = n15183 & n15761;
  assign n15763 = po10  & n15762;
  assign n15764 = po10  & n15761;
  assign n15765 = ~n15183 & ~n15764;
  assign n15766 = ~n15763 & ~n15765;
  assign n15767 = ~po41  & n15759;
  assign n15768 = ~n15766 & ~n15767;
  assign n15769 = ~n15760 & ~n15768;
  assign n15770 = po42  & ~n15769;
  assign n15771 = ~n15188 & ~n15195;
  assign n15772 = n15194 & n15771;
  assign n15773 = po10  & n15772;
  assign n15774 = po10  & n15771;
  assign n15775 = ~n15194 & ~n15774;
  assign n15776 = ~n15773 & ~n15775;
  assign n15777 = ~po42  & ~n15760;
  assign n15778 = ~n15768 & n15777;
  assign n15779 = ~n15776 & ~n15778;
  assign n15780 = ~n15770 & ~n15779;
  assign n15781 = po43  & ~n15780;
  assign n15782 = ~n15198 & ~n15206;
  assign n15783 = n15204 & n15782;
  assign n15784 = po10  & n15783;
  assign n15785 = po10  & n15782;
  assign n15786 = ~n15204 & ~n15785;
  assign n15787 = ~n15784 & ~n15786;
  assign n15788 = ~po43  & n15780;
  assign n15789 = ~n15787 & ~n15788;
  assign n15790 = ~n15781 & ~n15789;
  assign n15791 = po44  & ~n15790;
  assign n15792 = ~n15209 & ~n15216;
  assign n15793 = n15215 & n15792;
  assign n15794 = po10  & n15793;
  assign n15795 = po10  & n15792;
  assign n15796 = ~n15215 & ~n15795;
  assign n15797 = ~n15794 & ~n15796;
  assign n15798 = ~po44  & ~n15781;
  assign n15799 = ~n15789 & n15798;
  assign n15800 = ~n15797 & ~n15799;
  assign n15801 = ~n15791 & ~n15800;
  assign n15802 = po45  & ~n15801;
  assign n15803 = ~n15219 & ~n15227;
  assign n15804 = n15225 & n15803;
  assign n15805 = po10  & n15804;
  assign n15806 = po10  & n15803;
  assign n15807 = ~n15225 & ~n15806;
  assign n15808 = ~n15805 & ~n15807;
  assign n15809 = ~po45  & n15801;
  assign n15810 = ~n15808 & ~n15809;
  assign n15811 = ~n15802 & ~n15810;
  assign n15812 = po46  & ~n15811;
  assign n15813 = ~n15230 & ~n15237;
  assign n15814 = n15236 & n15813;
  assign n15815 = po10  & n15814;
  assign n15816 = po10  & n15813;
  assign n15817 = ~n15236 & ~n15816;
  assign n15818 = ~n15815 & ~n15817;
  assign n15819 = ~po46  & ~n15802;
  assign n15820 = ~n15810 & n15819;
  assign n15821 = ~n15818 & ~n15820;
  assign n15822 = ~n15812 & ~n15821;
  assign n15823 = po47  & ~n15822;
  assign n15824 = ~n15240 & ~n15248;
  assign n15825 = n15246 & n15824;
  assign n15826 = po10  & n15825;
  assign n15827 = po10  & n15824;
  assign n15828 = ~n15246 & ~n15827;
  assign n15829 = ~n15826 & ~n15828;
  assign n15830 = ~po47  & n15822;
  assign n15831 = ~n15829 & ~n15830;
  assign n15832 = ~n15823 & ~n15831;
  assign n15833 = po48  & ~n15832;
  assign n15834 = ~n15251 & ~n15258;
  assign n15835 = n15257 & n15834;
  assign n15836 = po10  & n15835;
  assign n15837 = po10  & n15834;
  assign n15838 = ~n15257 & ~n15837;
  assign n15839 = ~n15836 & ~n15838;
  assign n15840 = ~po48  & ~n15823;
  assign n15841 = ~n15831 & n15840;
  assign n15842 = ~n15839 & ~n15841;
  assign n15843 = ~n15833 & ~n15842;
  assign n15844 = po49  & ~n15843;
  assign n15845 = ~n15261 & ~n15269;
  assign n15846 = n15267 & n15845;
  assign n15847 = po10  & n15846;
  assign n15848 = po10  & n15845;
  assign n15849 = ~n15267 & ~n15848;
  assign n15850 = ~n15847 & ~n15849;
  assign n15851 = ~po49  & n15843;
  assign n15852 = ~n15850 & ~n15851;
  assign n15853 = ~n15844 & ~n15852;
  assign n15854 = po50  & ~n15853;
  assign n15855 = ~n15272 & ~n15279;
  assign n15856 = n15278 & n15855;
  assign n15857 = po10  & n15856;
  assign n15858 = po10  & n15855;
  assign n15859 = ~n15278 & ~n15858;
  assign n15860 = ~n15857 & ~n15859;
  assign n15861 = ~po50  & ~n15844;
  assign n15862 = ~n15852 & n15861;
  assign n15863 = ~n15860 & ~n15862;
  assign n15864 = ~n15854 & ~n15863;
  assign n15865 = po51  & ~n15864;
  assign n15866 = ~n15282 & ~n15290;
  assign n15867 = n15288 & n15866;
  assign n15868 = po10  & n15867;
  assign n15869 = po10  & n15866;
  assign n15870 = ~n15288 & ~n15869;
  assign n15871 = ~n15868 & ~n15870;
  assign n15872 = ~po51  & n15864;
  assign n15873 = ~n15871 & ~n15872;
  assign n15874 = ~n15865 & ~n15873;
  assign n15875 = po52  & ~n15874;
  assign n15876 = ~n15293 & ~n15300;
  assign n15877 = n15299 & n15876;
  assign n15878 = po10  & n15877;
  assign n15879 = po10  & n15876;
  assign n15880 = ~n15299 & ~n15879;
  assign n15881 = ~n15878 & ~n15880;
  assign n15882 = ~po52  & ~n15865;
  assign n15883 = ~n15873 & n15882;
  assign n15884 = ~n15881 & ~n15883;
  assign n15885 = ~n15875 & ~n15884;
  assign n15886 = po53  & ~n15885;
  assign n15887 = ~n15303 & ~n15311;
  assign n15888 = n15309 & n15887;
  assign n15889 = po10  & n15888;
  assign n15890 = po10  & n15887;
  assign n15891 = ~n15309 & ~n15890;
  assign n15892 = ~n15889 & ~n15891;
  assign n15893 = ~po53  & n15885;
  assign n15894 = ~n15892 & ~n15893;
  assign n15895 = ~n15886 & ~n15894;
  assign n15896 = po54  & ~n15895;
  assign n15897 = ~n15314 & ~n15321;
  assign n15898 = n15320 & n15897;
  assign n15899 = po10  & n15898;
  assign n15900 = po10  & n15897;
  assign n15901 = ~n15320 & ~n15900;
  assign n15902 = ~n15899 & ~n15901;
  assign n15903 = ~po54  & ~n15886;
  assign n15904 = ~n15894 & n15903;
  assign n15905 = ~n15902 & ~n15904;
  assign n15906 = ~n15896 & ~n15905;
  assign n15907 = po55  & ~n15906;
  assign n15908 = ~n15324 & ~n15326;
  assign n15909 = n15332 & n15908;
  assign n15910 = po10  & n15909;
  assign n15911 = po10  & n15908;
  assign n15912 = ~n15332 & ~n15911;
  assign n15913 = ~n15910 & ~n15912;
  assign n15914 = ~po55  & n15906;
  assign n15915 = ~n15913 & ~n15914;
  assign n15916 = ~n15907 & ~n15915;
  assign n15917 = po56  & ~n15916;
  assign n15918 = ~n15335 & ~n15342;
  assign n15919 = n15341 & n15918;
  assign n15920 = po10  & n15919;
  assign n15921 = po10  & n15918;
  assign n15922 = ~n15341 & ~n15921;
  assign n15923 = ~n15920 & ~n15922;
  assign n15924 = ~po56  & ~n15907;
  assign n15925 = ~n15915 & n15924;
  assign n15926 = ~n15923 & ~n15925;
  assign n15927 = ~n15917 & ~n15926;
  assign n15928 = po57  & ~n15927;
  assign n15929 = ~n15345 & ~n15353;
  assign n15930 = n15351 & n15929;
  assign n15931 = po10  & n15930;
  assign n15932 = po10  & n15929;
  assign n15933 = ~n15351 & ~n15932;
  assign n15934 = ~n15931 & ~n15933;
  assign n15935 = ~po57  & n15927;
  assign n15936 = ~n15934 & ~n15935;
  assign n15937 = ~n15928 & ~n15936;
  assign n15938 = po58  & ~n15937;
  assign n15939 = ~n15356 & ~n15363;
  assign n15940 = n15362 & n15939;
  assign n15941 = po10  & n15940;
  assign n15942 = po10  & n15939;
  assign n15943 = ~n15362 & ~n15942;
  assign n15944 = ~n15941 & ~n15943;
  assign n15945 = ~po58  & ~n15928;
  assign n15946 = ~n15936 & n15945;
  assign n15947 = ~n15944 & ~n15946;
  assign n15948 = ~n15938 & ~n15947;
  assign n15949 = po59  & ~n15948;
  assign n15950 = ~n15366 & ~n15374;
  assign n15951 = n15372 & n15950;
  assign n15952 = po10  & n15951;
  assign n15953 = po10  & n15950;
  assign n15954 = ~n15372 & ~n15953;
  assign n15955 = ~n15952 & ~n15954;
  assign n15956 = ~po59  & n15948;
  assign n15957 = ~n15955 & ~n15956;
  assign n15958 = ~n15949 & ~n15957;
  assign n15959 = po60  & ~n15958;
  assign n15960 = ~n15377 & ~n15384;
  assign n15961 = n15383 & n15960;
  assign n15962 = po10  & n15961;
  assign n15963 = po10  & n15960;
  assign n15964 = ~n15383 & ~n15963;
  assign n15965 = ~n15962 & ~n15964;
  assign n15966 = ~po60  & ~n15949;
  assign n15967 = ~n15957 & n15966;
  assign n15968 = ~n15965 & ~n15967;
  assign n15969 = ~n15959 & ~n15968;
  assign n15970 = po61  & ~n15969;
  assign n15971 = ~n15387 & ~n15395;
  assign n15972 = n15393 & n15971;
  assign n15973 = po10  & n15972;
  assign n15974 = po10  & n15971;
  assign n15975 = ~n15393 & ~n15974;
  assign n15976 = ~n15973 & ~n15975;
  assign n15977 = ~po61  & n15969;
  assign n15978 = ~n15976 & ~n15977;
  assign n15979 = ~n15970 & ~n15978;
  assign n15980 = po62  & ~n15979;
  assign n15981 = ~n15398 & ~n15405;
  assign n15982 = n15404 & n15981;
  assign n15983 = po10  & n15982;
  assign n15984 = po10  & n15981;
  assign n15985 = ~n15404 & ~n15984;
  assign n15986 = ~n15983 & ~n15985;
  assign n15987 = ~po62  & ~n15970;
  assign n15988 = ~n15978 & n15987;
  assign n15989 = ~n15986 & ~n15988;
  assign n15990 = ~n15980 & ~n15989;
  assign n15991 = ~n15408 & ~n15416;
  assign n15992 = po10  & n15991;
  assign n15993 = ~n15414 & ~n15992;
  assign n15994 = n15414 & n15992;
  assign n15995 = ~n15993 & ~n15994;
  assign n15996 = ~n15418 & ~n15423;
  assign n15997 = po10  & n15996;
  assign n15998 = ~n15436 & ~n15997;
  assign n15999 = ~n15995 & n15998;
  assign n16000 = ~n15990 & n15999;
  assign n16001 = ~po63  & ~n16000;
  assign n16002 = ~n15423 & po10 ;
  assign n16003 = n15418 & ~n16002;
  assign n16004 = po63  & ~n15996;
  assign n16005 = ~n16003 & n16004;
  assign n16006 = n15423 & ~po10 ;
  assign n16007 = ~n16005 & ~n16006;
  assign n16008 = n15990 & n15995;
  assign n16009 = n16007 & ~n16008;
  assign po9  = n16001 | ~n16009;
  assign n16011 = pi18  & po9 ;
  assign n16012 = ~pi16  & ~pi17 ;
  assign n16013 = ~pi18  & n16012;
  assign n16014 = ~n16011 & ~n16013;
  assign n16015 = po10  & ~n16014;
  assign n16016 = n15435 & ~n16013;
  assign n16017 = ~n15436 & n16016;
  assign n16018 = ~n15429 & n16017;
  assign n16019 = ~n16011 & n16018;
  assign n16020 = ~pi18  & po9 ;
  assign n16021 = pi19  & ~n16020;
  assign n16022 = n15440 & po9 ;
  assign n16023 = ~n16021 & ~n16022;
  assign n16024 = ~n16019 & n16023;
  assign n16025 = ~n16015 & ~n16024;
  assign n16026 = po11  & ~n16025;
  assign n16027 = po10  & n16007;
  assign n16028 = ~n16008 & n16027;
  assign n16029 = ~n16001 & n16028;
  assign n16030 = ~n16022 & ~n16029;
  assign n16031 = pi20  & ~n16030;
  assign n16032 = ~pi20  & n16030;
  assign n16033 = ~n16031 & ~n16032;
  assign n16034 = ~po11  & n16025;
  assign n16035 = ~n16033 & ~n16034;
  assign n16036 = ~n16026 & ~n16035;
  assign n16037 = po12  & ~n16036;
  assign n16038 = ~n15443 & ~n15447;
  assign n16039 = ~n15451 & n16038;
  assign n16040 = po9  & n16039;
  assign n16041 = po9  & n16038;
  assign n16042 = n15451 & ~n16041;
  assign n16043 = ~n16040 & ~n16042;
  assign n16044 = ~po12  & ~n16026;
  assign n16045 = ~n16035 & n16044;
  assign n16046 = ~n16043 & ~n16045;
  assign n16047 = ~n16037 & ~n16046;
  assign n16048 = po13  & ~n16047;
  assign n16049 = ~n15454 & ~n15456;
  assign n16050 = n15463 & n16049;
  assign n16051 = po9  & n16050;
  assign n16052 = po9  & n16049;
  assign n16053 = ~n15463 & ~n16052;
  assign n16054 = ~n16051 & ~n16053;
  assign n16055 = ~po13  & n16047;
  assign n16056 = ~n16054 & ~n16055;
  assign n16057 = ~n16048 & ~n16056;
  assign n16058 = po14  & ~n16057;
  assign n16059 = ~n15466 & ~n15473;
  assign n16060 = n15472 & n16059;
  assign n16061 = po9  & n16060;
  assign n16062 = po9  & n16059;
  assign n16063 = ~n15472 & ~n16062;
  assign n16064 = ~n16061 & ~n16063;
  assign n16065 = ~po14  & ~n16048;
  assign n16066 = ~n16056 & n16065;
  assign n16067 = ~n16064 & ~n16066;
  assign n16068 = ~n16058 & ~n16067;
  assign n16069 = po15  & ~n16068;
  assign n16070 = ~n15476 & ~n15484;
  assign n16071 = n15482 & n16070;
  assign n16072 = po9  & n16071;
  assign n16073 = po9  & n16070;
  assign n16074 = ~n15482 & ~n16073;
  assign n16075 = ~n16072 & ~n16074;
  assign n16076 = ~po15  & n16068;
  assign n16077 = ~n16075 & ~n16076;
  assign n16078 = ~n16069 & ~n16077;
  assign n16079 = po16  & ~n16078;
  assign n16080 = ~n15487 & ~n15494;
  assign n16081 = n15493 & n16080;
  assign n16082 = po9  & n16081;
  assign n16083 = po9  & n16080;
  assign n16084 = ~n15493 & ~n16083;
  assign n16085 = ~n16082 & ~n16084;
  assign n16086 = ~po16  & ~n16069;
  assign n16087 = ~n16077 & n16086;
  assign n16088 = ~n16085 & ~n16087;
  assign n16089 = ~n16079 & ~n16088;
  assign n16090 = po17  & ~n16089;
  assign n16091 = ~n15497 & ~n15505;
  assign n16092 = n15503 & n16091;
  assign n16093 = po9  & n16092;
  assign n16094 = po9  & n16091;
  assign n16095 = ~n15503 & ~n16094;
  assign n16096 = ~n16093 & ~n16095;
  assign n16097 = ~po17  & n16089;
  assign n16098 = ~n16096 & ~n16097;
  assign n16099 = ~n16090 & ~n16098;
  assign n16100 = po18  & ~n16099;
  assign n16101 = ~n15508 & ~n15515;
  assign n16102 = n15514 & n16101;
  assign n16103 = po9  & n16102;
  assign n16104 = po9  & n16101;
  assign n16105 = ~n15514 & ~n16104;
  assign n16106 = ~n16103 & ~n16105;
  assign n16107 = ~po18  & ~n16090;
  assign n16108 = ~n16098 & n16107;
  assign n16109 = ~n16106 & ~n16108;
  assign n16110 = ~n16100 & ~n16109;
  assign n16111 = po19  & ~n16110;
  assign n16112 = ~n15518 & ~n15526;
  assign n16113 = n15524 & n16112;
  assign n16114 = po9  & n16113;
  assign n16115 = po9  & n16112;
  assign n16116 = ~n15524 & ~n16115;
  assign n16117 = ~n16114 & ~n16116;
  assign n16118 = ~po19  & n16110;
  assign n16119 = ~n16117 & ~n16118;
  assign n16120 = ~n16111 & ~n16119;
  assign n16121 = po20  & ~n16120;
  assign n16122 = ~n15529 & ~n15536;
  assign n16123 = n15535 & n16122;
  assign n16124 = po9  & n16123;
  assign n16125 = po9  & n16122;
  assign n16126 = ~n15535 & ~n16125;
  assign n16127 = ~n16124 & ~n16126;
  assign n16128 = ~po20  & ~n16111;
  assign n16129 = ~n16119 & n16128;
  assign n16130 = ~n16127 & ~n16129;
  assign n16131 = ~n16121 & ~n16130;
  assign n16132 = po21  & ~n16131;
  assign n16133 = ~n15539 & ~n15547;
  assign n16134 = n15545 & n16133;
  assign n16135 = po9  & n16134;
  assign n16136 = po9  & n16133;
  assign n16137 = ~n15545 & ~n16136;
  assign n16138 = ~n16135 & ~n16137;
  assign n16139 = ~po21  & n16131;
  assign n16140 = ~n16138 & ~n16139;
  assign n16141 = ~n16132 & ~n16140;
  assign n16142 = po22  & ~n16141;
  assign n16143 = ~n15550 & ~n15557;
  assign n16144 = n15556 & n16143;
  assign n16145 = po9  & n16144;
  assign n16146 = po9  & n16143;
  assign n16147 = ~n15556 & ~n16146;
  assign n16148 = ~n16145 & ~n16147;
  assign n16149 = ~po22  & ~n16132;
  assign n16150 = ~n16140 & n16149;
  assign n16151 = ~n16148 & ~n16150;
  assign n16152 = ~n16142 & ~n16151;
  assign n16153 = po23  & ~n16152;
  assign n16154 = ~n15560 & ~n15568;
  assign n16155 = n15566 & n16154;
  assign n16156 = po9  & n16155;
  assign n16157 = po9  & n16154;
  assign n16158 = ~n15566 & ~n16157;
  assign n16159 = ~n16156 & ~n16158;
  assign n16160 = ~po23  & n16152;
  assign n16161 = ~n16159 & ~n16160;
  assign n16162 = ~n16153 & ~n16161;
  assign n16163 = po24  & ~n16162;
  assign n16164 = ~n15571 & ~n15578;
  assign n16165 = n15577 & n16164;
  assign n16166 = po9  & n16165;
  assign n16167 = po9  & n16164;
  assign n16168 = ~n15577 & ~n16167;
  assign n16169 = ~n16166 & ~n16168;
  assign n16170 = ~po24  & ~n16153;
  assign n16171 = ~n16161 & n16170;
  assign n16172 = ~n16169 & ~n16171;
  assign n16173 = ~n16163 & ~n16172;
  assign n16174 = po25  & ~n16173;
  assign n16175 = ~n15581 & ~n15589;
  assign n16176 = n15587 & n16175;
  assign n16177 = po9  & n16176;
  assign n16178 = po9  & n16175;
  assign n16179 = ~n15587 & ~n16178;
  assign n16180 = ~n16177 & ~n16179;
  assign n16181 = ~po25  & n16173;
  assign n16182 = ~n16180 & ~n16181;
  assign n16183 = ~n16174 & ~n16182;
  assign n16184 = po26  & ~n16183;
  assign n16185 = ~n15592 & ~n15599;
  assign n16186 = n15598 & n16185;
  assign n16187 = po9  & n16186;
  assign n16188 = po9  & n16185;
  assign n16189 = ~n15598 & ~n16188;
  assign n16190 = ~n16187 & ~n16189;
  assign n16191 = ~po26  & ~n16174;
  assign n16192 = ~n16182 & n16191;
  assign n16193 = ~n16190 & ~n16192;
  assign n16194 = ~n16184 & ~n16193;
  assign n16195 = po27  & ~n16194;
  assign n16196 = ~n15602 & ~n15610;
  assign n16197 = n15608 & n16196;
  assign n16198 = po9  & n16197;
  assign n16199 = po9  & n16196;
  assign n16200 = ~n15608 & ~n16199;
  assign n16201 = ~n16198 & ~n16200;
  assign n16202 = ~po27  & n16194;
  assign n16203 = ~n16201 & ~n16202;
  assign n16204 = ~n16195 & ~n16203;
  assign n16205 = po28  & ~n16204;
  assign n16206 = ~n15613 & ~n15620;
  assign n16207 = n15619 & n16206;
  assign n16208 = po9  & n16207;
  assign n16209 = po9  & n16206;
  assign n16210 = ~n15619 & ~n16209;
  assign n16211 = ~n16208 & ~n16210;
  assign n16212 = ~po28  & ~n16195;
  assign n16213 = ~n16203 & n16212;
  assign n16214 = ~n16211 & ~n16213;
  assign n16215 = ~n16205 & ~n16214;
  assign n16216 = po29  & ~n16215;
  assign n16217 = ~n15623 & ~n15631;
  assign n16218 = n15629 & n16217;
  assign n16219 = po9  & n16218;
  assign n16220 = po9  & n16217;
  assign n16221 = ~n15629 & ~n16220;
  assign n16222 = ~n16219 & ~n16221;
  assign n16223 = ~po29  & n16215;
  assign n16224 = ~n16222 & ~n16223;
  assign n16225 = ~n16216 & ~n16224;
  assign n16226 = po30  & ~n16225;
  assign n16227 = ~n15634 & ~n15641;
  assign n16228 = n15640 & n16227;
  assign n16229 = po9  & n16228;
  assign n16230 = po9  & n16227;
  assign n16231 = ~n15640 & ~n16230;
  assign n16232 = ~n16229 & ~n16231;
  assign n16233 = ~po30  & ~n16216;
  assign n16234 = ~n16224 & n16233;
  assign n16235 = ~n16232 & ~n16234;
  assign n16236 = ~n16226 & ~n16235;
  assign n16237 = po31  & ~n16236;
  assign n16238 = ~n15644 & ~n15652;
  assign n16239 = n15650 & n16238;
  assign n16240 = po9  & n16239;
  assign n16241 = po9  & n16238;
  assign n16242 = ~n15650 & ~n16241;
  assign n16243 = ~n16240 & ~n16242;
  assign n16244 = ~po31  & n16236;
  assign n16245 = ~n16243 & ~n16244;
  assign n16246 = ~n16237 & ~n16245;
  assign n16247 = po32  & ~n16246;
  assign n16248 = ~n15655 & ~n15662;
  assign n16249 = n15661 & n16248;
  assign n16250 = po9  & n16249;
  assign n16251 = po9  & n16248;
  assign n16252 = ~n15661 & ~n16251;
  assign n16253 = ~n16250 & ~n16252;
  assign n16254 = ~po32  & ~n16237;
  assign n16255 = ~n16245 & n16254;
  assign n16256 = ~n16253 & ~n16255;
  assign n16257 = ~n16247 & ~n16256;
  assign n16258 = po33  & ~n16257;
  assign n16259 = ~n15665 & ~n15673;
  assign n16260 = n15671 & n16259;
  assign n16261 = po9  & n16260;
  assign n16262 = po9  & n16259;
  assign n16263 = ~n15671 & ~n16262;
  assign n16264 = ~n16261 & ~n16263;
  assign n16265 = ~po33  & n16257;
  assign n16266 = ~n16264 & ~n16265;
  assign n16267 = ~n16258 & ~n16266;
  assign n16268 = po34  & ~n16267;
  assign n16269 = ~n15676 & ~n15683;
  assign n16270 = n15682 & n16269;
  assign n16271 = po9  & n16270;
  assign n16272 = po9  & n16269;
  assign n16273 = ~n15682 & ~n16272;
  assign n16274 = ~n16271 & ~n16273;
  assign n16275 = ~po34  & ~n16258;
  assign n16276 = ~n16266 & n16275;
  assign n16277 = ~n16274 & ~n16276;
  assign n16278 = ~n16268 & ~n16277;
  assign n16279 = po35  & ~n16278;
  assign n16280 = ~n15686 & ~n15694;
  assign n16281 = n15692 & n16280;
  assign n16282 = po9  & n16281;
  assign n16283 = po9  & n16280;
  assign n16284 = ~n15692 & ~n16283;
  assign n16285 = ~n16282 & ~n16284;
  assign n16286 = ~po35  & n16278;
  assign n16287 = ~n16285 & ~n16286;
  assign n16288 = ~n16279 & ~n16287;
  assign n16289 = po36  & ~n16288;
  assign n16290 = ~n15697 & ~n15704;
  assign n16291 = n15703 & n16290;
  assign n16292 = po9  & n16291;
  assign n16293 = po9  & n16290;
  assign n16294 = ~n15703 & ~n16293;
  assign n16295 = ~n16292 & ~n16294;
  assign n16296 = ~po36  & ~n16279;
  assign n16297 = ~n16287 & n16296;
  assign n16298 = ~n16295 & ~n16297;
  assign n16299 = ~n16289 & ~n16298;
  assign n16300 = po37  & ~n16299;
  assign n16301 = ~n15707 & ~n15715;
  assign n16302 = n15713 & n16301;
  assign n16303 = po9  & n16302;
  assign n16304 = po9  & n16301;
  assign n16305 = ~n15713 & ~n16304;
  assign n16306 = ~n16303 & ~n16305;
  assign n16307 = ~po37  & n16299;
  assign n16308 = ~n16306 & ~n16307;
  assign n16309 = ~n16300 & ~n16308;
  assign n16310 = po38  & ~n16309;
  assign n16311 = ~n15718 & ~n15725;
  assign n16312 = n15724 & n16311;
  assign n16313 = po9  & n16312;
  assign n16314 = po9  & n16311;
  assign n16315 = ~n15724 & ~n16314;
  assign n16316 = ~n16313 & ~n16315;
  assign n16317 = ~po38  & ~n16300;
  assign n16318 = ~n16308 & n16317;
  assign n16319 = ~n16316 & ~n16318;
  assign n16320 = ~n16310 & ~n16319;
  assign n16321 = po39  & ~n16320;
  assign n16322 = ~n15728 & ~n15736;
  assign n16323 = n15734 & n16322;
  assign n16324 = po9  & n16323;
  assign n16325 = po9  & n16322;
  assign n16326 = ~n15734 & ~n16325;
  assign n16327 = ~n16324 & ~n16326;
  assign n16328 = ~po39  & n16320;
  assign n16329 = ~n16327 & ~n16328;
  assign n16330 = ~n16321 & ~n16329;
  assign n16331 = po40  & ~n16330;
  assign n16332 = ~n15739 & ~n15746;
  assign n16333 = n15745 & n16332;
  assign n16334 = po9  & n16333;
  assign n16335 = po9  & n16332;
  assign n16336 = ~n15745 & ~n16335;
  assign n16337 = ~n16334 & ~n16336;
  assign n16338 = ~po40  & ~n16321;
  assign n16339 = ~n16329 & n16338;
  assign n16340 = ~n16337 & ~n16339;
  assign n16341 = ~n16331 & ~n16340;
  assign n16342 = po41  & ~n16341;
  assign n16343 = ~n15749 & ~n15757;
  assign n16344 = n15755 & n16343;
  assign n16345 = po9  & n16344;
  assign n16346 = po9  & n16343;
  assign n16347 = ~n15755 & ~n16346;
  assign n16348 = ~n16345 & ~n16347;
  assign n16349 = ~po41  & n16341;
  assign n16350 = ~n16348 & ~n16349;
  assign n16351 = ~n16342 & ~n16350;
  assign n16352 = po42  & ~n16351;
  assign n16353 = ~n15760 & ~n15767;
  assign n16354 = n15766 & n16353;
  assign n16355 = po9  & n16354;
  assign n16356 = po9  & n16353;
  assign n16357 = ~n15766 & ~n16356;
  assign n16358 = ~n16355 & ~n16357;
  assign n16359 = ~po42  & ~n16342;
  assign n16360 = ~n16350 & n16359;
  assign n16361 = ~n16358 & ~n16360;
  assign n16362 = ~n16352 & ~n16361;
  assign n16363 = po43  & ~n16362;
  assign n16364 = ~n15770 & ~n15778;
  assign n16365 = n15776 & n16364;
  assign n16366 = po9  & n16365;
  assign n16367 = po9  & n16364;
  assign n16368 = ~n15776 & ~n16367;
  assign n16369 = ~n16366 & ~n16368;
  assign n16370 = ~po43  & n16362;
  assign n16371 = ~n16369 & ~n16370;
  assign n16372 = ~n16363 & ~n16371;
  assign n16373 = po44  & ~n16372;
  assign n16374 = ~n15781 & ~n15788;
  assign n16375 = n15787 & n16374;
  assign n16376 = po9  & n16375;
  assign n16377 = po9  & n16374;
  assign n16378 = ~n15787 & ~n16377;
  assign n16379 = ~n16376 & ~n16378;
  assign n16380 = ~po44  & ~n16363;
  assign n16381 = ~n16371 & n16380;
  assign n16382 = ~n16379 & ~n16381;
  assign n16383 = ~n16373 & ~n16382;
  assign n16384 = po45  & ~n16383;
  assign n16385 = ~n15791 & ~n15799;
  assign n16386 = n15797 & n16385;
  assign n16387 = po9  & n16386;
  assign n16388 = po9  & n16385;
  assign n16389 = ~n15797 & ~n16388;
  assign n16390 = ~n16387 & ~n16389;
  assign n16391 = ~po45  & n16383;
  assign n16392 = ~n16390 & ~n16391;
  assign n16393 = ~n16384 & ~n16392;
  assign n16394 = po46  & ~n16393;
  assign n16395 = ~n15802 & ~n15809;
  assign n16396 = n15808 & n16395;
  assign n16397 = po9  & n16396;
  assign n16398 = po9  & n16395;
  assign n16399 = ~n15808 & ~n16398;
  assign n16400 = ~n16397 & ~n16399;
  assign n16401 = ~po46  & ~n16384;
  assign n16402 = ~n16392 & n16401;
  assign n16403 = ~n16400 & ~n16402;
  assign n16404 = ~n16394 & ~n16403;
  assign n16405 = po47  & ~n16404;
  assign n16406 = ~n15812 & ~n15820;
  assign n16407 = n15818 & n16406;
  assign n16408 = po9  & n16407;
  assign n16409 = po9  & n16406;
  assign n16410 = ~n15818 & ~n16409;
  assign n16411 = ~n16408 & ~n16410;
  assign n16412 = ~po47  & n16404;
  assign n16413 = ~n16411 & ~n16412;
  assign n16414 = ~n16405 & ~n16413;
  assign n16415 = po48  & ~n16414;
  assign n16416 = ~n15823 & ~n15830;
  assign n16417 = n15829 & n16416;
  assign n16418 = po9  & n16417;
  assign n16419 = po9  & n16416;
  assign n16420 = ~n15829 & ~n16419;
  assign n16421 = ~n16418 & ~n16420;
  assign n16422 = ~po48  & ~n16405;
  assign n16423 = ~n16413 & n16422;
  assign n16424 = ~n16421 & ~n16423;
  assign n16425 = ~n16415 & ~n16424;
  assign n16426 = po49  & ~n16425;
  assign n16427 = ~n15833 & ~n15841;
  assign n16428 = n15839 & n16427;
  assign n16429 = po9  & n16428;
  assign n16430 = po9  & n16427;
  assign n16431 = ~n15839 & ~n16430;
  assign n16432 = ~n16429 & ~n16431;
  assign n16433 = ~po49  & n16425;
  assign n16434 = ~n16432 & ~n16433;
  assign n16435 = ~n16426 & ~n16434;
  assign n16436 = po50  & ~n16435;
  assign n16437 = ~n15844 & ~n15851;
  assign n16438 = n15850 & n16437;
  assign n16439 = po9  & n16438;
  assign n16440 = po9  & n16437;
  assign n16441 = ~n15850 & ~n16440;
  assign n16442 = ~n16439 & ~n16441;
  assign n16443 = ~po50  & ~n16426;
  assign n16444 = ~n16434 & n16443;
  assign n16445 = ~n16442 & ~n16444;
  assign n16446 = ~n16436 & ~n16445;
  assign n16447 = po51  & ~n16446;
  assign n16448 = ~n15854 & ~n15862;
  assign n16449 = n15860 & n16448;
  assign n16450 = po9  & n16449;
  assign n16451 = po9  & n16448;
  assign n16452 = ~n15860 & ~n16451;
  assign n16453 = ~n16450 & ~n16452;
  assign n16454 = ~po51  & n16446;
  assign n16455 = ~n16453 & ~n16454;
  assign n16456 = ~n16447 & ~n16455;
  assign n16457 = po52  & ~n16456;
  assign n16458 = ~n15865 & ~n15872;
  assign n16459 = n15871 & n16458;
  assign n16460 = po9  & n16459;
  assign n16461 = po9  & n16458;
  assign n16462 = ~n15871 & ~n16461;
  assign n16463 = ~n16460 & ~n16462;
  assign n16464 = ~po52  & ~n16447;
  assign n16465 = ~n16455 & n16464;
  assign n16466 = ~n16463 & ~n16465;
  assign n16467 = ~n16457 & ~n16466;
  assign n16468 = po53  & ~n16467;
  assign n16469 = ~n15875 & ~n15883;
  assign n16470 = n15881 & n16469;
  assign n16471 = po9  & n16470;
  assign n16472 = po9  & n16469;
  assign n16473 = ~n15881 & ~n16472;
  assign n16474 = ~n16471 & ~n16473;
  assign n16475 = ~po53  & n16467;
  assign n16476 = ~n16474 & ~n16475;
  assign n16477 = ~n16468 & ~n16476;
  assign n16478 = po54  & ~n16477;
  assign n16479 = ~n15886 & ~n15893;
  assign n16480 = n15892 & n16479;
  assign n16481 = po9  & n16480;
  assign n16482 = po9  & n16479;
  assign n16483 = ~n15892 & ~n16482;
  assign n16484 = ~n16481 & ~n16483;
  assign n16485 = ~po54  & ~n16468;
  assign n16486 = ~n16476 & n16485;
  assign n16487 = ~n16484 & ~n16486;
  assign n16488 = ~n16478 & ~n16487;
  assign n16489 = po55  & ~n16488;
  assign n16490 = ~n15896 & ~n15904;
  assign n16491 = n15902 & n16490;
  assign n16492 = po9  & n16491;
  assign n16493 = po9  & n16490;
  assign n16494 = ~n15902 & ~n16493;
  assign n16495 = ~n16492 & ~n16494;
  assign n16496 = ~po55  & n16488;
  assign n16497 = ~n16495 & ~n16496;
  assign n16498 = ~n16489 & ~n16497;
  assign n16499 = po56  & ~n16498;
  assign n16500 = ~po56  & ~n16489;
  assign n16501 = ~n16497 & n16500;
  assign n16502 = ~n15907 & ~n15914;
  assign n16503 = n15913 & n16502;
  assign n16504 = po9  & n16503;
  assign n16505 = po9  & n16502;
  assign n16506 = ~n15913 & ~n16505;
  assign n16507 = ~n16504 & ~n16506;
  assign n16508 = ~n16501 & ~n16507;
  assign n16509 = ~n16499 & ~n16508;
  assign n16510 = po57  & ~n16509;
  assign n16511 = ~n15917 & ~n15925;
  assign n16512 = n15923 & n16511;
  assign n16513 = po9  & n16512;
  assign n16514 = po9  & n16511;
  assign n16515 = ~n15923 & ~n16514;
  assign n16516 = ~n16513 & ~n16515;
  assign n16517 = ~po57  & n16509;
  assign n16518 = ~n16516 & ~n16517;
  assign n16519 = ~n16510 & ~n16518;
  assign n16520 = po58  & ~n16519;
  assign n16521 = ~n15928 & ~n15935;
  assign n16522 = n15934 & n16521;
  assign n16523 = po9  & n16522;
  assign n16524 = po9  & n16521;
  assign n16525 = ~n15934 & ~n16524;
  assign n16526 = ~n16523 & ~n16525;
  assign n16527 = ~po58  & ~n16510;
  assign n16528 = ~n16518 & n16527;
  assign n16529 = ~n16526 & ~n16528;
  assign n16530 = ~n16520 & ~n16529;
  assign n16531 = po59  & ~n16530;
  assign n16532 = ~n15938 & ~n15946;
  assign n16533 = n15944 & n16532;
  assign n16534 = po9  & n16533;
  assign n16535 = po9  & n16532;
  assign n16536 = ~n15944 & ~n16535;
  assign n16537 = ~n16534 & ~n16536;
  assign n16538 = ~po59  & n16530;
  assign n16539 = ~n16537 & ~n16538;
  assign n16540 = ~n16531 & ~n16539;
  assign n16541 = po60  & ~n16540;
  assign n16542 = ~n15949 & ~n15956;
  assign n16543 = n15955 & n16542;
  assign n16544 = po9  & n16543;
  assign n16545 = po9  & n16542;
  assign n16546 = ~n15955 & ~n16545;
  assign n16547 = ~n16544 & ~n16546;
  assign n16548 = ~po60  & ~n16531;
  assign n16549 = ~n16539 & n16548;
  assign n16550 = ~n16547 & ~n16549;
  assign n16551 = ~n16541 & ~n16550;
  assign n16552 = po61  & ~n16551;
  assign n16553 = ~n15959 & ~n15967;
  assign n16554 = n15965 & n16553;
  assign n16555 = po9  & n16554;
  assign n16556 = po9  & n16553;
  assign n16557 = ~n15965 & ~n16556;
  assign n16558 = ~n16555 & ~n16557;
  assign n16559 = ~po61  & n16551;
  assign n16560 = ~n16558 & ~n16559;
  assign n16561 = ~n16552 & ~n16560;
  assign n16562 = po62  & ~n16561;
  assign n16563 = ~n15970 & ~n15977;
  assign n16564 = n15976 & n16563;
  assign n16565 = po9  & n16564;
  assign n16566 = po9  & n16563;
  assign n16567 = ~n15976 & ~n16566;
  assign n16568 = ~n16565 & ~n16567;
  assign n16569 = ~po62  & ~n16552;
  assign n16570 = ~n16560 & n16569;
  assign n16571 = ~n16568 & ~n16570;
  assign n16572 = ~n16562 & ~n16571;
  assign n16573 = ~n15980 & ~n15988;
  assign n16574 = po9  & n16573;
  assign n16575 = ~n15986 & ~n16574;
  assign n16576 = n15986 & n16574;
  assign n16577 = ~n16575 & ~n16576;
  assign n16578 = ~n15990 & ~n15995;
  assign n16579 = po9  & n16578;
  assign n16580 = ~n16008 & ~n16579;
  assign n16581 = ~n16577 & n16580;
  assign n16582 = ~n16572 & n16581;
  assign n16583 = ~po63  & ~n16582;
  assign n16584 = ~n15995 & po9 ;
  assign n16585 = n15990 & ~n16584;
  assign n16586 = po63  & ~n16578;
  assign n16587 = ~n16585 & n16586;
  assign n16588 = n15995 & ~po9 ;
  assign n16589 = ~n16587 & ~n16588;
  assign n16590 = n16572 & n16577;
  assign n16591 = n16589 & ~n16590;
  assign po8  = n16583 | ~n16591;
  assign n16593 = pi16  & po8 ;
  assign n16594 = ~pi14  & ~pi15 ;
  assign n16595 = ~pi16  & n16594;
  assign n16596 = ~n16593 & ~n16595;
  assign n16597 = po9  & ~n16596;
  assign n16598 = n16007 & ~n16595;
  assign n16599 = ~n16008 & n16598;
  assign n16600 = ~n16001 & n16599;
  assign n16601 = ~n16593 & n16600;
  assign n16602 = ~pi16  & po8 ;
  assign n16603 = pi17  & ~n16602;
  assign n16604 = n16012 & po8 ;
  assign n16605 = ~n16603 & ~n16604;
  assign n16606 = ~n16601 & n16605;
  assign n16607 = ~n16597 & ~n16606;
  assign n16608 = po10  & ~n16607;
  assign n16609 = ~po10  & ~n16597;
  assign n16610 = ~n16606 & n16609;
  assign n16611 = po9  & n16589;
  assign n16612 = ~n16590 & n16611;
  assign n16613 = ~n16583 & n16612;
  assign n16614 = ~n16604 & ~n16613;
  assign n16615 = pi18  & ~n16614;
  assign n16616 = ~pi18  & n16614;
  assign n16617 = ~n16615 & ~n16616;
  assign n16618 = ~n16610 & ~n16617;
  assign n16619 = ~n16608 & ~n16618;
  assign n16620 = po11  & ~n16619;
  assign n16621 = ~n16015 & ~n16019;
  assign n16622 = ~n16023 & n16621;
  assign n16623 = po8  & n16622;
  assign n16624 = po8  & n16621;
  assign n16625 = n16023 & ~n16624;
  assign n16626 = ~n16623 & ~n16625;
  assign n16627 = ~po11  & n16619;
  assign n16628 = ~n16626 & ~n16627;
  assign n16629 = ~n16620 & ~n16628;
  assign n16630 = po12  & ~n16629;
  assign n16631 = ~n16026 & ~n16034;
  assign n16632 = n16033 & n16631;
  assign n16633 = po8  & n16632;
  assign n16634 = po8  & n16631;
  assign n16635 = ~n16033 & ~n16634;
  assign n16636 = ~n16633 & ~n16635;
  assign n16637 = ~po12  & ~n16620;
  assign n16638 = ~n16628 & n16637;
  assign n16639 = ~n16636 & ~n16638;
  assign n16640 = ~n16630 & ~n16639;
  assign n16641 = po13  & ~n16640;
  assign n16642 = ~n16037 & ~n16045;
  assign n16643 = n16043 & n16642;
  assign n16644 = po8  & n16643;
  assign n16645 = po8  & n16642;
  assign n16646 = ~n16043 & ~n16645;
  assign n16647 = ~n16644 & ~n16646;
  assign n16648 = ~po13  & n16640;
  assign n16649 = ~n16647 & ~n16648;
  assign n16650 = ~n16641 & ~n16649;
  assign n16651 = po14  & ~n16650;
  assign n16652 = ~n16048 & ~n16055;
  assign n16653 = n16054 & n16652;
  assign n16654 = po8  & n16653;
  assign n16655 = po8  & n16652;
  assign n16656 = ~n16054 & ~n16655;
  assign n16657 = ~n16654 & ~n16656;
  assign n16658 = ~po14  & ~n16641;
  assign n16659 = ~n16649 & n16658;
  assign n16660 = ~n16657 & ~n16659;
  assign n16661 = ~n16651 & ~n16660;
  assign n16662 = po15  & ~n16661;
  assign n16663 = ~n16058 & ~n16066;
  assign n16664 = n16064 & n16663;
  assign n16665 = po8  & n16664;
  assign n16666 = po8  & n16663;
  assign n16667 = ~n16064 & ~n16666;
  assign n16668 = ~n16665 & ~n16667;
  assign n16669 = ~po15  & n16661;
  assign n16670 = ~n16668 & ~n16669;
  assign n16671 = ~n16662 & ~n16670;
  assign n16672 = po16  & ~n16671;
  assign n16673 = ~n16069 & ~n16076;
  assign n16674 = n16075 & n16673;
  assign n16675 = po8  & n16674;
  assign n16676 = po8  & n16673;
  assign n16677 = ~n16075 & ~n16676;
  assign n16678 = ~n16675 & ~n16677;
  assign n16679 = ~po16  & ~n16662;
  assign n16680 = ~n16670 & n16679;
  assign n16681 = ~n16678 & ~n16680;
  assign n16682 = ~n16672 & ~n16681;
  assign n16683 = po17  & ~n16682;
  assign n16684 = ~n16079 & ~n16087;
  assign n16685 = n16085 & n16684;
  assign n16686 = po8  & n16685;
  assign n16687 = po8  & n16684;
  assign n16688 = ~n16085 & ~n16687;
  assign n16689 = ~n16686 & ~n16688;
  assign n16690 = ~po17  & n16682;
  assign n16691 = ~n16689 & ~n16690;
  assign n16692 = ~n16683 & ~n16691;
  assign n16693 = po18  & ~n16692;
  assign n16694 = ~n16090 & ~n16097;
  assign n16695 = n16096 & n16694;
  assign n16696 = po8  & n16695;
  assign n16697 = po8  & n16694;
  assign n16698 = ~n16096 & ~n16697;
  assign n16699 = ~n16696 & ~n16698;
  assign n16700 = ~po18  & ~n16683;
  assign n16701 = ~n16691 & n16700;
  assign n16702 = ~n16699 & ~n16701;
  assign n16703 = ~n16693 & ~n16702;
  assign n16704 = po19  & ~n16703;
  assign n16705 = ~n16100 & ~n16108;
  assign n16706 = n16106 & n16705;
  assign n16707 = po8  & n16706;
  assign n16708 = po8  & n16705;
  assign n16709 = ~n16106 & ~n16708;
  assign n16710 = ~n16707 & ~n16709;
  assign n16711 = ~po19  & n16703;
  assign n16712 = ~n16710 & ~n16711;
  assign n16713 = ~n16704 & ~n16712;
  assign n16714 = po20  & ~n16713;
  assign n16715 = ~n16111 & ~n16118;
  assign n16716 = n16117 & n16715;
  assign n16717 = po8  & n16716;
  assign n16718 = po8  & n16715;
  assign n16719 = ~n16117 & ~n16718;
  assign n16720 = ~n16717 & ~n16719;
  assign n16721 = ~po20  & ~n16704;
  assign n16722 = ~n16712 & n16721;
  assign n16723 = ~n16720 & ~n16722;
  assign n16724 = ~n16714 & ~n16723;
  assign n16725 = po21  & ~n16724;
  assign n16726 = ~n16121 & ~n16129;
  assign n16727 = n16127 & n16726;
  assign n16728 = po8  & n16727;
  assign n16729 = po8  & n16726;
  assign n16730 = ~n16127 & ~n16729;
  assign n16731 = ~n16728 & ~n16730;
  assign n16732 = ~po21  & n16724;
  assign n16733 = ~n16731 & ~n16732;
  assign n16734 = ~n16725 & ~n16733;
  assign n16735 = po22  & ~n16734;
  assign n16736 = ~n16132 & ~n16139;
  assign n16737 = n16138 & n16736;
  assign n16738 = po8  & n16737;
  assign n16739 = po8  & n16736;
  assign n16740 = ~n16138 & ~n16739;
  assign n16741 = ~n16738 & ~n16740;
  assign n16742 = ~po22  & ~n16725;
  assign n16743 = ~n16733 & n16742;
  assign n16744 = ~n16741 & ~n16743;
  assign n16745 = ~n16735 & ~n16744;
  assign n16746 = po23  & ~n16745;
  assign n16747 = ~n16142 & ~n16150;
  assign n16748 = n16148 & n16747;
  assign n16749 = po8  & n16748;
  assign n16750 = po8  & n16747;
  assign n16751 = ~n16148 & ~n16750;
  assign n16752 = ~n16749 & ~n16751;
  assign n16753 = ~po23  & n16745;
  assign n16754 = ~n16752 & ~n16753;
  assign n16755 = ~n16746 & ~n16754;
  assign n16756 = po24  & ~n16755;
  assign n16757 = ~n16153 & ~n16160;
  assign n16758 = n16159 & n16757;
  assign n16759 = po8  & n16758;
  assign n16760 = po8  & n16757;
  assign n16761 = ~n16159 & ~n16760;
  assign n16762 = ~n16759 & ~n16761;
  assign n16763 = ~po24  & ~n16746;
  assign n16764 = ~n16754 & n16763;
  assign n16765 = ~n16762 & ~n16764;
  assign n16766 = ~n16756 & ~n16765;
  assign n16767 = po25  & ~n16766;
  assign n16768 = ~n16163 & ~n16171;
  assign n16769 = n16169 & n16768;
  assign n16770 = po8  & n16769;
  assign n16771 = po8  & n16768;
  assign n16772 = ~n16169 & ~n16771;
  assign n16773 = ~n16770 & ~n16772;
  assign n16774 = ~po25  & n16766;
  assign n16775 = ~n16773 & ~n16774;
  assign n16776 = ~n16767 & ~n16775;
  assign n16777 = po26  & ~n16776;
  assign n16778 = ~n16174 & ~n16181;
  assign n16779 = n16180 & n16778;
  assign n16780 = po8  & n16779;
  assign n16781 = po8  & n16778;
  assign n16782 = ~n16180 & ~n16781;
  assign n16783 = ~n16780 & ~n16782;
  assign n16784 = ~po26  & ~n16767;
  assign n16785 = ~n16775 & n16784;
  assign n16786 = ~n16783 & ~n16785;
  assign n16787 = ~n16777 & ~n16786;
  assign n16788 = po27  & ~n16787;
  assign n16789 = ~n16184 & ~n16192;
  assign n16790 = n16190 & n16789;
  assign n16791 = po8  & n16790;
  assign n16792 = po8  & n16789;
  assign n16793 = ~n16190 & ~n16792;
  assign n16794 = ~n16791 & ~n16793;
  assign n16795 = ~po27  & n16787;
  assign n16796 = ~n16794 & ~n16795;
  assign n16797 = ~n16788 & ~n16796;
  assign n16798 = po28  & ~n16797;
  assign n16799 = ~n16195 & ~n16202;
  assign n16800 = n16201 & n16799;
  assign n16801 = po8  & n16800;
  assign n16802 = po8  & n16799;
  assign n16803 = ~n16201 & ~n16802;
  assign n16804 = ~n16801 & ~n16803;
  assign n16805 = ~po28  & ~n16788;
  assign n16806 = ~n16796 & n16805;
  assign n16807 = ~n16804 & ~n16806;
  assign n16808 = ~n16798 & ~n16807;
  assign n16809 = po29  & ~n16808;
  assign n16810 = ~n16205 & ~n16213;
  assign n16811 = n16211 & n16810;
  assign n16812 = po8  & n16811;
  assign n16813 = po8  & n16810;
  assign n16814 = ~n16211 & ~n16813;
  assign n16815 = ~n16812 & ~n16814;
  assign n16816 = ~po29  & n16808;
  assign n16817 = ~n16815 & ~n16816;
  assign n16818 = ~n16809 & ~n16817;
  assign n16819 = po30  & ~n16818;
  assign n16820 = ~n16216 & ~n16223;
  assign n16821 = n16222 & n16820;
  assign n16822 = po8  & n16821;
  assign n16823 = po8  & n16820;
  assign n16824 = ~n16222 & ~n16823;
  assign n16825 = ~n16822 & ~n16824;
  assign n16826 = ~po30  & ~n16809;
  assign n16827 = ~n16817 & n16826;
  assign n16828 = ~n16825 & ~n16827;
  assign n16829 = ~n16819 & ~n16828;
  assign n16830 = po31  & ~n16829;
  assign n16831 = ~n16226 & ~n16234;
  assign n16832 = n16232 & n16831;
  assign n16833 = po8  & n16832;
  assign n16834 = po8  & n16831;
  assign n16835 = ~n16232 & ~n16834;
  assign n16836 = ~n16833 & ~n16835;
  assign n16837 = ~po31  & n16829;
  assign n16838 = ~n16836 & ~n16837;
  assign n16839 = ~n16830 & ~n16838;
  assign n16840 = po32  & ~n16839;
  assign n16841 = ~n16237 & ~n16244;
  assign n16842 = n16243 & n16841;
  assign n16843 = po8  & n16842;
  assign n16844 = po8  & n16841;
  assign n16845 = ~n16243 & ~n16844;
  assign n16846 = ~n16843 & ~n16845;
  assign n16847 = ~po32  & ~n16830;
  assign n16848 = ~n16838 & n16847;
  assign n16849 = ~n16846 & ~n16848;
  assign n16850 = ~n16840 & ~n16849;
  assign n16851 = po33  & ~n16850;
  assign n16852 = ~n16247 & ~n16255;
  assign n16853 = n16253 & n16852;
  assign n16854 = po8  & n16853;
  assign n16855 = po8  & n16852;
  assign n16856 = ~n16253 & ~n16855;
  assign n16857 = ~n16854 & ~n16856;
  assign n16858 = ~po33  & n16850;
  assign n16859 = ~n16857 & ~n16858;
  assign n16860 = ~n16851 & ~n16859;
  assign n16861 = po34  & ~n16860;
  assign n16862 = ~n16258 & ~n16265;
  assign n16863 = n16264 & n16862;
  assign n16864 = po8  & n16863;
  assign n16865 = po8  & n16862;
  assign n16866 = ~n16264 & ~n16865;
  assign n16867 = ~n16864 & ~n16866;
  assign n16868 = ~po34  & ~n16851;
  assign n16869 = ~n16859 & n16868;
  assign n16870 = ~n16867 & ~n16869;
  assign n16871 = ~n16861 & ~n16870;
  assign n16872 = po35  & ~n16871;
  assign n16873 = ~n16268 & ~n16276;
  assign n16874 = n16274 & n16873;
  assign n16875 = po8  & n16874;
  assign n16876 = po8  & n16873;
  assign n16877 = ~n16274 & ~n16876;
  assign n16878 = ~n16875 & ~n16877;
  assign n16879 = ~po35  & n16871;
  assign n16880 = ~n16878 & ~n16879;
  assign n16881 = ~n16872 & ~n16880;
  assign n16882 = po36  & ~n16881;
  assign n16883 = ~n16279 & ~n16286;
  assign n16884 = n16285 & n16883;
  assign n16885 = po8  & n16884;
  assign n16886 = po8  & n16883;
  assign n16887 = ~n16285 & ~n16886;
  assign n16888 = ~n16885 & ~n16887;
  assign n16889 = ~po36  & ~n16872;
  assign n16890 = ~n16880 & n16889;
  assign n16891 = ~n16888 & ~n16890;
  assign n16892 = ~n16882 & ~n16891;
  assign n16893 = po37  & ~n16892;
  assign n16894 = ~n16289 & ~n16297;
  assign n16895 = n16295 & n16894;
  assign n16896 = po8  & n16895;
  assign n16897 = po8  & n16894;
  assign n16898 = ~n16295 & ~n16897;
  assign n16899 = ~n16896 & ~n16898;
  assign n16900 = ~po37  & n16892;
  assign n16901 = ~n16899 & ~n16900;
  assign n16902 = ~n16893 & ~n16901;
  assign n16903 = po38  & ~n16902;
  assign n16904 = ~n16300 & ~n16307;
  assign n16905 = n16306 & n16904;
  assign n16906 = po8  & n16905;
  assign n16907 = po8  & n16904;
  assign n16908 = ~n16306 & ~n16907;
  assign n16909 = ~n16906 & ~n16908;
  assign n16910 = ~po38  & ~n16893;
  assign n16911 = ~n16901 & n16910;
  assign n16912 = ~n16909 & ~n16911;
  assign n16913 = ~n16903 & ~n16912;
  assign n16914 = po39  & ~n16913;
  assign n16915 = ~n16310 & ~n16318;
  assign n16916 = n16316 & n16915;
  assign n16917 = po8  & n16916;
  assign n16918 = po8  & n16915;
  assign n16919 = ~n16316 & ~n16918;
  assign n16920 = ~n16917 & ~n16919;
  assign n16921 = ~po39  & n16913;
  assign n16922 = ~n16920 & ~n16921;
  assign n16923 = ~n16914 & ~n16922;
  assign n16924 = po40  & ~n16923;
  assign n16925 = ~n16321 & ~n16328;
  assign n16926 = n16327 & n16925;
  assign n16927 = po8  & n16926;
  assign n16928 = po8  & n16925;
  assign n16929 = ~n16327 & ~n16928;
  assign n16930 = ~n16927 & ~n16929;
  assign n16931 = ~po40  & ~n16914;
  assign n16932 = ~n16922 & n16931;
  assign n16933 = ~n16930 & ~n16932;
  assign n16934 = ~n16924 & ~n16933;
  assign n16935 = po41  & ~n16934;
  assign n16936 = ~n16331 & ~n16339;
  assign n16937 = n16337 & n16936;
  assign n16938 = po8  & n16937;
  assign n16939 = po8  & n16936;
  assign n16940 = ~n16337 & ~n16939;
  assign n16941 = ~n16938 & ~n16940;
  assign n16942 = ~po41  & n16934;
  assign n16943 = ~n16941 & ~n16942;
  assign n16944 = ~n16935 & ~n16943;
  assign n16945 = po42  & ~n16944;
  assign n16946 = ~n16342 & ~n16349;
  assign n16947 = n16348 & n16946;
  assign n16948 = po8  & n16947;
  assign n16949 = po8  & n16946;
  assign n16950 = ~n16348 & ~n16949;
  assign n16951 = ~n16948 & ~n16950;
  assign n16952 = ~po42  & ~n16935;
  assign n16953 = ~n16943 & n16952;
  assign n16954 = ~n16951 & ~n16953;
  assign n16955 = ~n16945 & ~n16954;
  assign n16956 = po43  & ~n16955;
  assign n16957 = ~n16352 & ~n16360;
  assign n16958 = n16358 & n16957;
  assign n16959 = po8  & n16958;
  assign n16960 = po8  & n16957;
  assign n16961 = ~n16358 & ~n16960;
  assign n16962 = ~n16959 & ~n16961;
  assign n16963 = ~po43  & n16955;
  assign n16964 = ~n16962 & ~n16963;
  assign n16965 = ~n16956 & ~n16964;
  assign n16966 = po44  & ~n16965;
  assign n16967 = ~n16363 & ~n16370;
  assign n16968 = n16369 & n16967;
  assign n16969 = po8  & n16968;
  assign n16970 = po8  & n16967;
  assign n16971 = ~n16369 & ~n16970;
  assign n16972 = ~n16969 & ~n16971;
  assign n16973 = ~po44  & ~n16956;
  assign n16974 = ~n16964 & n16973;
  assign n16975 = ~n16972 & ~n16974;
  assign n16976 = ~n16966 & ~n16975;
  assign n16977 = po45  & ~n16976;
  assign n16978 = ~n16373 & ~n16381;
  assign n16979 = n16379 & n16978;
  assign n16980 = po8  & n16979;
  assign n16981 = po8  & n16978;
  assign n16982 = ~n16379 & ~n16981;
  assign n16983 = ~n16980 & ~n16982;
  assign n16984 = ~po45  & n16976;
  assign n16985 = ~n16983 & ~n16984;
  assign n16986 = ~n16977 & ~n16985;
  assign n16987 = po46  & ~n16986;
  assign n16988 = ~n16384 & ~n16391;
  assign n16989 = n16390 & n16988;
  assign n16990 = po8  & n16989;
  assign n16991 = po8  & n16988;
  assign n16992 = ~n16390 & ~n16991;
  assign n16993 = ~n16990 & ~n16992;
  assign n16994 = ~po46  & ~n16977;
  assign n16995 = ~n16985 & n16994;
  assign n16996 = ~n16993 & ~n16995;
  assign n16997 = ~n16987 & ~n16996;
  assign n16998 = po47  & ~n16997;
  assign n16999 = ~n16394 & ~n16402;
  assign n17000 = n16400 & n16999;
  assign n17001 = po8  & n17000;
  assign n17002 = po8  & n16999;
  assign n17003 = ~n16400 & ~n17002;
  assign n17004 = ~n17001 & ~n17003;
  assign n17005 = ~po47  & n16997;
  assign n17006 = ~n17004 & ~n17005;
  assign n17007 = ~n16998 & ~n17006;
  assign n17008 = po48  & ~n17007;
  assign n17009 = ~n16405 & ~n16412;
  assign n17010 = n16411 & n17009;
  assign n17011 = po8  & n17010;
  assign n17012 = po8  & n17009;
  assign n17013 = ~n16411 & ~n17012;
  assign n17014 = ~n17011 & ~n17013;
  assign n17015 = ~po48  & ~n16998;
  assign n17016 = ~n17006 & n17015;
  assign n17017 = ~n17014 & ~n17016;
  assign n17018 = ~n17008 & ~n17017;
  assign n17019 = po49  & ~n17018;
  assign n17020 = ~n16415 & ~n16423;
  assign n17021 = n16421 & n17020;
  assign n17022 = po8  & n17021;
  assign n17023 = po8  & n17020;
  assign n17024 = ~n16421 & ~n17023;
  assign n17025 = ~n17022 & ~n17024;
  assign n17026 = ~po49  & n17018;
  assign n17027 = ~n17025 & ~n17026;
  assign n17028 = ~n17019 & ~n17027;
  assign n17029 = po50  & ~n17028;
  assign n17030 = ~n16426 & ~n16433;
  assign n17031 = n16432 & n17030;
  assign n17032 = po8  & n17031;
  assign n17033 = po8  & n17030;
  assign n17034 = ~n16432 & ~n17033;
  assign n17035 = ~n17032 & ~n17034;
  assign n17036 = ~po50  & ~n17019;
  assign n17037 = ~n17027 & n17036;
  assign n17038 = ~n17035 & ~n17037;
  assign n17039 = ~n17029 & ~n17038;
  assign n17040 = po51  & ~n17039;
  assign n17041 = ~n16436 & ~n16444;
  assign n17042 = n16442 & n17041;
  assign n17043 = po8  & n17042;
  assign n17044 = po8  & n17041;
  assign n17045 = ~n16442 & ~n17044;
  assign n17046 = ~n17043 & ~n17045;
  assign n17047 = ~po51  & n17039;
  assign n17048 = ~n17046 & ~n17047;
  assign n17049 = ~n17040 & ~n17048;
  assign n17050 = po52  & ~n17049;
  assign n17051 = ~n16447 & ~n16454;
  assign n17052 = n16453 & n17051;
  assign n17053 = po8  & n17052;
  assign n17054 = po8  & n17051;
  assign n17055 = ~n16453 & ~n17054;
  assign n17056 = ~n17053 & ~n17055;
  assign n17057 = ~po52  & ~n17040;
  assign n17058 = ~n17048 & n17057;
  assign n17059 = ~n17056 & ~n17058;
  assign n17060 = ~n17050 & ~n17059;
  assign n17061 = po53  & ~n17060;
  assign n17062 = ~n16457 & ~n16465;
  assign n17063 = n16463 & n17062;
  assign n17064 = po8  & n17063;
  assign n17065 = po8  & n17062;
  assign n17066 = ~n16463 & ~n17065;
  assign n17067 = ~n17064 & ~n17066;
  assign n17068 = ~po53  & n17060;
  assign n17069 = ~n17067 & ~n17068;
  assign n17070 = ~n17061 & ~n17069;
  assign n17071 = po54  & ~n17070;
  assign n17072 = ~n16468 & ~n16475;
  assign n17073 = n16474 & n17072;
  assign n17074 = po8  & n17073;
  assign n17075 = po8  & n17072;
  assign n17076 = ~n16474 & ~n17075;
  assign n17077 = ~n17074 & ~n17076;
  assign n17078 = ~po54  & ~n17061;
  assign n17079 = ~n17069 & n17078;
  assign n17080 = ~n17077 & ~n17079;
  assign n17081 = ~n17071 & ~n17080;
  assign n17082 = po55  & ~n17081;
  assign n17083 = ~n16478 & ~n16486;
  assign n17084 = n16484 & n17083;
  assign n17085 = po8  & n17084;
  assign n17086 = po8  & n17083;
  assign n17087 = ~n16484 & ~n17086;
  assign n17088 = ~n17085 & ~n17087;
  assign n17089 = ~po55  & n17081;
  assign n17090 = ~n17088 & ~n17089;
  assign n17091 = ~n17082 & ~n17090;
  assign n17092 = po56  & ~n17091;
  assign n17093 = ~n16489 & ~n16496;
  assign n17094 = n16495 & n17093;
  assign n17095 = po8  & n17094;
  assign n17096 = po8  & n17093;
  assign n17097 = ~n16495 & ~n17096;
  assign n17098 = ~n17095 & ~n17097;
  assign n17099 = ~po56  & ~n17082;
  assign n17100 = ~n17090 & n17099;
  assign n17101 = ~n17098 & ~n17100;
  assign n17102 = ~n17092 & ~n17101;
  assign n17103 = po57  & ~n17102;
  assign n17104 = ~n16499 & ~n16501;
  assign n17105 = n16507 & n17104;
  assign n17106 = po8  & n17105;
  assign n17107 = po8  & n17104;
  assign n17108 = ~n16507 & ~n17107;
  assign n17109 = ~n17106 & ~n17108;
  assign n17110 = ~po57  & n17102;
  assign n17111 = ~n17109 & ~n17110;
  assign n17112 = ~n17103 & ~n17111;
  assign n17113 = po58  & ~n17112;
  assign n17114 = ~n16510 & ~n16517;
  assign n17115 = n16516 & n17114;
  assign n17116 = po8  & n17115;
  assign n17117 = po8  & n17114;
  assign n17118 = ~n16516 & ~n17117;
  assign n17119 = ~n17116 & ~n17118;
  assign n17120 = ~po58  & ~n17103;
  assign n17121 = ~n17111 & n17120;
  assign n17122 = ~n17119 & ~n17121;
  assign n17123 = ~n17113 & ~n17122;
  assign n17124 = po59  & ~n17123;
  assign n17125 = ~n16520 & ~n16528;
  assign n17126 = n16526 & n17125;
  assign n17127 = po8  & n17126;
  assign n17128 = po8  & n17125;
  assign n17129 = ~n16526 & ~n17128;
  assign n17130 = ~n17127 & ~n17129;
  assign n17131 = ~po59  & n17123;
  assign n17132 = ~n17130 & ~n17131;
  assign n17133 = ~n17124 & ~n17132;
  assign n17134 = po60  & ~n17133;
  assign n17135 = ~n16531 & ~n16538;
  assign n17136 = n16537 & n17135;
  assign n17137 = po8  & n17136;
  assign n17138 = po8  & n17135;
  assign n17139 = ~n16537 & ~n17138;
  assign n17140 = ~n17137 & ~n17139;
  assign n17141 = ~po60  & ~n17124;
  assign n17142 = ~n17132 & n17141;
  assign n17143 = ~n17140 & ~n17142;
  assign n17144 = ~n17134 & ~n17143;
  assign n17145 = po61  & ~n17144;
  assign n17146 = ~n16541 & ~n16549;
  assign n17147 = n16547 & n17146;
  assign n17148 = po8  & n17147;
  assign n17149 = po8  & n17146;
  assign n17150 = ~n16547 & ~n17149;
  assign n17151 = ~n17148 & ~n17150;
  assign n17152 = ~po61  & n17144;
  assign n17153 = ~n17151 & ~n17152;
  assign n17154 = ~n17145 & ~n17153;
  assign n17155 = po62  & ~n17154;
  assign n17156 = ~n16552 & ~n16559;
  assign n17157 = n16558 & n17156;
  assign n17158 = po8  & n17157;
  assign n17159 = po8  & n17156;
  assign n17160 = ~n16558 & ~n17159;
  assign n17161 = ~n17158 & ~n17160;
  assign n17162 = ~po62  & ~n17145;
  assign n17163 = ~n17153 & n17162;
  assign n17164 = ~n17161 & ~n17163;
  assign n17165 = ~n17155 & ~n17164;
  assign n17166 = ~n16562 & ~n16570;
  assign n17167 = po8  & n17166;
  assign n17168 = ~n16568 & ~n17167;
  assign n17169 = n16568 & n17167;
  assign n17170 = ~n17168 & ~n17169;
  assign n17171 = ~n16572 & ~n16577;
  assign n17172 = po8  & n17171;
  assign n17173 = ~n16590 & ~n17172;
  assign n17174 = ~n17170 & n17173;
  assign n17175 = ~n17165 & n17174;
  assign n17176 = ~po63  & ~n17175;
  assign n17177 = ~n16577 & po8 ;
  assign n17178 = n16572 & ~n17177;
  assign n17179 = po63  & ~n17171;
  assign n17180 = ~n17178 & n17179;
  assign n17181 = n16577 & ~po8 ;
  assign n17182 = ~n17180 & ~n17181;
  assign n17183 = n17165 & n17170;
  assign n17184 = n17182 & ~n17183;
  assign po7  = n17176 | ~n17184;
  assign n17186 = pi14  & po7 ;
  assign n17187 = ~pi12  & ~pi13 ;
  assign n17188 = ~pi14  & n17187;
  assign n17189 = ~n17186 & ~n17188;
  assign n17190 = po8  & ~n17189;
  assign n17191 = n16589 & ~n17188;
  assign n17192 = ~n16590 & n17191;
  assign n17193 = ~n16583 & n17192;
  assign n17194 = ~n17186 & n17193;
  assign n17195 = ~pi14  & po7 ;
  assign n17196 = pi15  & ~n17195;
  assign n17197 = n16594 & po7 ;
  assign n17198 = ~n17196 & ~n17197;
  assign n17199 = ~n17194 & n17198;
  assign n17200 = ~n17190 & ~n17199;
  assign n17201 = po9  & ~n17200;
  assign n17202 = po8  & n17182;
  assign n17203 = ~n17183 & n17202;
  assign n17204 = ~n17176 & n17203;
  assign n17205 = ~n17197 & ~n17204;
  assign n17206 = pi16  & ~n17205;
  assign n17207 = ~pi16  & n17205;
  assign n17208 = ~n17206 & ~n17207;
  assign n17209 = ~po9  & n17200;
  assign n17210 = ~n17208 & ~n17209;
  assign n17211 = ~n17201 & ~n17210;
  assign n17212 = po10  & ~n17211;
  assign n17213 = ~n16597 & ~n16601;
  assign n17214 = ~n16605 & n17213;
  assign n17215 = po7  & n17214;
  assign n17216 = po7  & n17213;
  assign n17217 = n16605 & ~n17216;
  assign n17218 = ~n17215 & ~n17217;
  assign n17219 = ~po10  & ~n17201;
  assign n17220 = ~n17210 & n17219;
  assign n17221 = ~n17218 & ~n17220;
  assign n17222 = ~n17212 & ~n17221;
  assign n17223 = po11  & ~n17222;
  assign n17224 = ~n16608 & ~n16610;
  assign n17225 = n16617 & n17224;
  assign n17226 = po7  & n17225;
  assign n17227 = po7  & n17224;
  assign n17228 = ~n16617 & ~n17227;
  assign n17229 = ~n17226 & ~n17228;
  assign n17230 = ~po11  & n17222;
  assign n17231 = ~n17229 & ~n17230;
  assign n17232 = ~n17223 & ~n17231;
  assign n17233 = po12  & ~n17232;
  assign n17234 = ~n16620 & ~n16627;
  assign n17235 = n16626 & n17234;
  assign n17236 = po7  & n17235;
  assign n17237 = po7  & n17234;
  assign n17238 = ~n16626 & ~n17237;
  assign n17239 = ~n17236 & ~n17238;
  assign n17240 = ~po12  & ~n17223;
  assign n17241 = ~n17231 & n17240;
  assign n17242 = ~n17239 & ~n17241;
  assign n17243 = ~n17233 & ~n17242;
  assign n17244 = po13  & ~n17243;
  assign n17245 = ~n16630 & ~n16638;
  assign n17246 = n16636 & n17245;
  assign n17247 = po7  & n17246;
  assign n17248 = po7  & n17245;
  assign n17249 = ~n16636 & ~n17248;
  assign n17250 = ~n17247 & ~n17249;
  assign n17251 = ~po13  & n17243;
  assign n17252 = ~n17250 & ~n17251;
  assign n17253 = ~n17244 & ~n17252;
  assign n17254 = po14  & ~n17253;
  assign n17255 = ~n16641 & ~n16648;
  assign n17256 = n16647 & n17255;
  assign n17257 = po7  & n17256;
  assign n17258 = po7  & n17255;
  assign n17259 = ~n16647 & ~n17258;
  assign n17260 = ~n17257 & ~n17259;
  assign n17261 = ~po14  & ~n17244;
  assign n17262 = ~n17252 & n17261;
  assign n17263 = ~n17260 & ~n17262;
  assign n17264 = ~n17254 & ~n17263;
  assign n17265 = po15  & ~n17264;
  assign n17266 = ~n16651 & ~n16659;
  assign n17267 = n16657 & n17266;
  assign n17268 = po7  & n17267;
  assign n17269 = po7  & n17266;
  assign n17270 = ~n16657 & ~n17269;
  assign n17271 = ~n17268 & ~n17270;
  assign n17272 = ~po15  & n17264;
  assign n17273 = ~n17271 & ~n17272;
  assign n17274 = ~n17265 & ~n17273;
  assign n17275 = po16  & ~n17274;
  assign n17276 = ~n16662 & ~n16669;
  assign n17277 = n16668 & n17276;
  assign n17278 = po7  & n17277;
  assign n17279 = po7  & n17276;
  assign n17280 = ~n16668 & ~n17279;
  assign n17281 = ~n17278 & ~n17280;
  assign n17282 = ~po16  & ~n17265;
  assign n17283 = ~n17273 & n17282;
  assign n17284 = ~n17281 & ~n17283;
  assign n17285 = ~n17275 & ~n17284;
  assign n17286 = po17  & ~n17285;
  assign n17287 = ~n16672 & ~n16680;
  assign n17288 = n16678 & n17287;
  assign n17289 = po7  & n17288;
  assign n17290 = po7  & n17287;
  assign n17291 = ~n16678 & ~n17290;
  assign n17292 = ~n17289 & ~n17291;
  assign n17293 = ~po17  & n17285;
  assign n17294 = ~n17292 & ~n17293;
  assign n17295 = ~n17286 & ~n17294;
  assign n17296 = po18  & ~n17295;
  assign n17297 = ~n16683 & ~n16690;
  assign n17298 = n16689 & n17297;
  assign n17299 = po7  & n17298;
  assign n17300 = po7  & n17297;
  assign n17301 = ~n16689 & ~n17300;
  assign n17302 = ~n17299 & ~n17301;
  assign n17303 = ~po18  & ~n17286;
  assign n17304 = ~n17294 & n17303;
  assign n17305 = ~n17302 & ~n17304;
  assign n17306 = ~n17296 & ~n17305;
  assign n17307 = po19  & ~n17306;
  assign n17308 = ~n16693 & ~n16701;
  assign n17309 = n16699 & n17308;
  assign n17310 = po7  & n17309;
  assign n17311 = po7  & n17308;
  assign n17312 = ~n16699 & ~n17311;
  assign n17313 = ~n17310 & ~n17312;
  assign n17314 = ~po19  & n17306;
  assign n17315 = ~n17313 & ~n17314;
  assign n17316 = ~n17307 & ~n17315;
  assign n17317 = po20  & ~n17316;
  assign n17318 = ~n16704 & ~n16711;
  assign n17319 = n16710 & n17318;
  assign n17320 = po7  & n17319;
  assign n17321 = po7  & n17318;
  assign n17322 = ~n16710 & ~n17321;
  assign n17323 = ~n17320 & ~n17322;
  assign n17324 = ~po20  & ~n17307;
  assign n17325 = ~n17315 & n17324;
  assign n17326 = ~n17323 & ~n17325;
  assign n17327 = ~n17317 & ~n17326;
  assign n17328 = po21  & ~n17327;
  assign n17329 = ~n16714 & ~n16722;
  assign n17330 = n16720 & n17329;
  assign n17331 = po7  & n17330;
  assign n17332 = po7  & n17329;
  assign n17333 = ~n16720 & ~n17332;
  assign n17334 = ~n17331 & ~n17333;
  assign n17335 = ~po21  & n17327;
  assign n17336 = ~n17334 & ~n17335;
  assign n17337 = ~n17328 & ~n17336;
  assign n17338 = po22  & ~n17337;
  assign n17339 = ~n16725 & ~n16732;
  assign n17340 = n16731 & n17339;
  assign n17341 = po7  & n17340;
  assign n17342 = po7  & n17339;
  assign n17343 = ~n16731 & ~n17342;
  assign n17344 = ~n17341 & ~n17343;
  assign n17345 = ~po22  & ~n17328;
  assign n17346 = ~n17336 & n17345;
  assign n17347 = ~n17344 & ~n17346;
  assign n17348 = ~n17338 & ~n17347;
  assign n17349 = po23  & ~n17348;
  assign n17350 = ~n16735 & ~n16743;
  assign n17351 = n16741 & n17350;
  assign n17352 = po7  & n17351;
  assign n17353 = po7  & n17350;
  assign n17354 = ~n16741 & ~n17353;
  assign n17355 = ~n17352 & ~n17354;
  assign n17356 = ~po23  & n17348;
  assign n17357 = ~n17355 & ~n17356;
  assign n17358 = ~n17349 & ~n17357;
  assign n17359 = po24  & ~n17358;
  assign n17360 = ~n16746 & ~n16753;
  assign n17361 = n16752 & n17360;
  assign n17362 = po7  & n17361;
  assign n17363 = po7  & n17360;
  assign n17364 = ~n16752 & ~n17363;
  assign n17365 = ~n17362 & ~n17364;
  assign n17366 = ~po24  & ~n17349;
  assign n17367 = ~n17357 & n17366;
  assign n17368 = ~n17365 & ~n17367;
  assign n17369 = ~n17359 & ~n17368;
  assign n17370 = po25  & ~n17369;
  assign n17371 = ~n16756 & ~n16764;
  assign n17372 = n16762 & n17371;
  assign n17373 = po7  & n17372;
  assign n17374 = po7  & n17371;
  assign n17375 = ~n16762 & ~n17374;
  assign n17376 = ~n17373 & ~n17375;
  assign n17377 = ~po25  & n17369;
  assign n17378 = ~n17376 & ~n17377;
  assign n17379 = ~n17370 & ~n17378;
  assign n17380 = po26  & ~n17379;
  assign n17381 = ~n16767 & ~n16774;
  assign n17382 = n16773 & n17381;
  assign n17383 = po7  & n17382;
  assign n17384 = po7  & n17381;
  assign n17385 = ~n16773 & ~n17384;
  assign n17386 = ~n17383 & ~n17385;
  assign n17387 = ~po26  & ~n17370;
  assign n17388 = ~n17378 & n17387;
  assign n17389 = ~n17386 & ~n17388;
  assign n17390 = ~n17380 & ~n17389;
  assign n17391 = po27  & ~n17390;
  assign n17392 = ~n16777 & ~n16785;
  assign n17393 = n16783 & n17392;
  assign n17394 = po7  & n17393;
  assign n17395 = po7  & n17392;
  assign n17396 = ~n16783 & ~n17395;
  assign n17397 = ~n17394 & ~n17396;
  assign n17398 = ~po27  & n17390;
  assign n17399 = ~n17397 & ~n17398;
  assign n17400 = ~n17391 & ~n17399;
  assign n17401 = po28  & ~n17400;
  assign n17402 = ~n16788 & ~n16795;
  assign n17403 = n16794 & n17402;
  assign n17404 = po7  & n17403;
  assign n17405 = po7  & n17402;
  assign n17406 = ~n16794 & ~n17405;
  assign n17407 = ~n17404 & ~n17406;
  assign n17408 = ~po28  & ~n17391;
  assign n17409 = ~n17399 & n17408;
  assign n17410 = ~n17407 & ~n17409;
  assign n17411 = ~n17401 & ~n17410;
  assign n17412 = po29  & ~n17411;
  assign n17413 = ~n16798 & ~n16806;
  assign n17414 = n16804 & n17413;
  assign n17415 = po7  & n17414;
  assign n17416 = po7  & n17413;
  assign n17417 = ~n16804 & ~n17416;
  assign n17418 = ~n17415 & ~n17417;
  assign n17419 = ~po29  & n17411;
  assign n17420 = ~n17418 & ~n17419;
  assign n17421 = ~n17412 & ~n17420;
  assign n17422 = po30  & ~n17421;
  assign n17423 = ~n16809 & ~n16816;
  assign n17424 = n16815 & n17423;
  assign n17425 = po7  & n17424;
  assign n17426 = po7  & n17423;
  assign n17427 = ~n16815 & ~n17426;
  assign n17428 = ~n17425 & ~n17427;
  assign n17429 = ~po30  & ~n17412;
  assign n17430 = ~n17420 & n17429;
  assign n17431 = ~n17428 & ~n17430;
  assign n17432 = ~n17422 & ~n17431;
  assign n17433 = po31  & ~n17432;
  assign n17434 = ~n16819 & ~n16827;
  assign n17435 = n16825 & n17434;
  assign n17436 = po7  & n17435;
  assign n17437 = po7  & n17434;
  assign n17438 = ~n16825 & ~n17437;
  assign n17439 = ~n17436 & ~n17438;
  assign n17440 = ~po31  & n17432;
  assign n17441 = ~n17439 & ~n17440;
  assign n17442 = ~n17433 & ~n17441;
  assign n17443 = po32  & ~n17442;
  assign n17444 = ~n16830 & ~n16837;
  assign n17445 = n16836 & n17444;
  assign n17446 = po7  & n17445;
  assign n17447 = po7  & n17444;
  assign n17448 = ~n16836 & ~n17447;
  assign n17449 = ~n17446 & ~n17448;
  assign n17450 = ~po32  & ~n17433;
  assign n17451 = ~n17441 & n17450;
  assign n17452 = ~n17449 & ~n17451;
  assign n17453 = ~n17443 & ~n17452;
  assign n17454 = po33  & ~n17453;
  assign n17455 = ~n16840 & ~n16848;
  assign n17456 = n16846 & n17455;
  assign n17457 = po7  & n17456;
  assign n17458 = po7  & n17455;
  assign n17459 = ~n16846 & ~n17458;
  assign n17460 = ~n17457 & ~n17459;
  assign n17461 = ~po33  & n17453;
  assign n17462 = ~n17460 & ~n17461;
  assign n17463 = ~n17454 & ~n17462;
  assign n17464 = po34  & ~n17463;
  assign n17465 = ~n16851 & ~n16858;
  assign n17466 = n16857 & n17465;
  assign n17467 = po7  & n17466;
  assign n17468 = po7  & n17465;
  assign n17469 = ~n16857 & ~n17468;
  assign n17470 = ~n17467 & ~n17469;
  assign n17471 = ~po34  & ~n17454;
  assign n17472 = ~n17462 & n17471;
  assign n17473 = ~n17470 & ~n17472;
  assign n17474 = ~n17464 & ~n17473;
  assign n17475 = po35  & ~n17474;
  assign n17476 = ~n16861 & ~n16869;
  assign n17477 = n16867 & n17476;
  assign n17478 = po7  & n17477;
  assign n17479 = po7  & n17476;
  assign n17480 = ~n16867 & ~n17479;
  assign n17481 = ~n17478 & ~n17480;
  assign n17482 = ~po35  & n17474;
  assign n17483 = ~n17481 & ~n17482;
  assign n17484 = ~n17475 & ~n17483;
  assign n17485 = po36  & ~n17484;
  assign n17486 = ~n16872 & ~n16879;
  assign n17487 = n16878 & n17486;
  assign n17488 = po7  & n17487;
  assign n17489 = po7  & n17486;
  assign n17490 = ~n16878 & ~n17489;
  assign n17491 = ~n17488 & ~n17490;
  assign n17492 = ~po36  & ~n17475;
  assign n17493 = ~n17483 & n17492;
  assign n17494 = ~n17491 & ~n17493;
  assign n17495 = ~n17485 & ~n17494;
  assign n17496 = po37  & ~n17495;
  assign n17497 = ~n16882 & ~n16890;
  assign n17498 = n16888 & n17497;
  assign n17499 = po7  & n17498;
  assign n17500 = po7  & n17497;
  assign n17501 = ~n16888 & ~n17500;
  assign n17502 = ~n17499 & ~n17501;
  assign n17503 = ~po37  & n17495;
  assign n17504 = ~n17502 & ~n17503;
  assign n17505 = ~n17496 & ~n17504;
  assign n17506 = po38  & ~n17505;
  assign n17507 = ~n16893 & ~n16900;
  assign n17508 = n16899 & n17507;
  assign n17509 = po7  & n17508;
  assign n17510 = po7  & n17507;
  assign n17511 = ~n16899 & ~n17510;
  assign n17512 = ~n17509 & ~n17511;
  assign n17513 = ~po38  & ~n17496;
  assign n17514 = ~n17504 & n17513;
  assign n17515 = ~n17512 & ~n17514;
  assign n17516 = ~n17506 & ~n17515;
  assign n17517 = po39  & ~n17516;
  assign n17518 = ~n16903 & ~n16911;
  assign n17519 = n16909 & n17518;
  assign n17520 = po7  & n17519;
  assign n17521 = po7  & n17518;
  assign n17522 = ~n16909 & ~n17521;
  assign n17523 = ~n17520 & ~n17522;
  assign n17524 = ~po39  & n17516;
  assign n17525 = ~n17523 & ~n17524;
  assign n17526 = ~n17517 & ~n17525;
  assign n17527 = po40  & ~n17526;
  assign n17528 = ~n16914 & ~n16921;
  assign n17529 = n16920 & n17528;
  assign n17530 = po7  & n17529;
  assign n17531 = po7  & n17528;
  assign n17532 = ~n16920 & ~n17531;
  assign n17533 = ~n17530 & ~n17532;
  assign n17534 = ~po40  & ~n17517;
  assign n17535 = ~n17525 & n17534;
  assign n17536 = ~n17533 & ~n17535;
  assign n17537 = ~n17527 & ~n17536;
  assign n17538 = po41  & ~n17537;
  assign n17539 = ~n16924 & ~n16932;
  assign n17540 = n16930 & n17539;
  assign n17541 = po7  & n17540;
  assign n17542 = po7  & n17539;
  assign n17543 = ~n16930 & ~n17542;
  assign n17544 = ~n17541 & ~n17543;
  assign n17545 = ~po41  & n17537;
  assign n17546 = ~n17544 & ~n17545;
  assign n17547 = ~n17538 & ~n17546;
  assign n17548 = po42  & ~n17547;
  assign n17549 = ~n16935 & ~n16942;
  assign n17550 = n16941 & n17549;
  assign n17551 = po7  & n17550;
  assign n17552 = po7  & n17549;
  assign n17553 = ~n16941 & ~n17552;
  assign n17554 = ~n17551 & ~n17553;
  assign n17555 = ~po42  & ~n17538;
  assign n17556 = ~n17546 & n17555;
  assign n17557 = ~n17554 & ~n17556;
  assign n17558 = ~n17548 & ~n17557;
  assign n17559 = po43  & ~n17558;
  assign n17560 = ~n16945 & ~n16953;
  assign n17561 = n16951 & n17560;
  assign n17562 = po7  & n17561;
  assign n17563 = po7  & n17560;
  assign n17564 = ~n16951 & ~n17563;
  assign n17565 = ~n17562 & ~n17564;
  assign n17566 = ~po43  & n17558;
  assign n17567 = ~n17565 & ~n17566;
  assign n17568 = ~n17559 & ~n17567;
  assign n17569 = po44  & ~n17568;
  assign n17570 = ~n16956 & ~n16963;
  assign n17571 = n16962 & n17570;
  assign n17572 = po7  & n17571;
  assign n17573 = po7  & n17570;
  assign n17574 = ~n16962 & ~n17573;
  assign n17575 = ~n17572 & ~n17574;
  assign n17576 = ~po44  & ~n17559;
  assign n17577 = ~n17567 & n17576;
  assign n17578 = ~n17575 & ~n17577;
  assign n17579 = ~n17569 & ~n17578;
  assign n17580 = po45  & ~n17579;
  assign n17581 = ~n16966 & ~n16974;
  assign n17582 = n16972 & n17581;
  assign n17583 = po7  & n17582;
  assign n17584 = po7  & n17581;
  assign n17585 = ~n16972 & ~n17584;
  assign n17586 = ~n17583 & ~n17585;
  assign n17587 = ~po45  & n17579;
  assign n17588 = ~n17586 & ~n17587;
  assign n17589 = ~n17580 & ~n17588;
  assign n17590 = po46  & ~n17589;
  assign n17591 = ~n16977 & ~n16984;
  assign n17592 = n16983 & n17591;
  assign n17593 = po7  & n17592;
  assign n17594 = po7  & n17591;
  assign n17595 = ~n16983 & ~n17594;
  assign n17596 = ~n17593 & ~n17595;
  assign n17597 = ~po46  & ~n17580;
  assign n17598 = ~n17588 & n17597;
  assign n17599 = ~n17596 & ~n17598;
  assign n17600 = ~n17590 & ~n17599;
  assign n17601 = po47  & ~n17600;
  assign n17602 = ~n16987 & ~n16995;
  assign n17603 = n16993 & n17602;
  assign n17604 = po7  & n17603;
  assign n17605 = po7  & n17602;
  assign n17606 = ~n16993 & ~n17605;
  assign n17607 = ~n17604 & ~n17606;
  assign n17608 = ~po47  & n17600;
  assign n17609 = ~n17607 & ~n17608;
  assign n17610 = ~n17601 & ~n17609;
  assign n17611 = po48  & ~n17610;
  assign n17612 = ~n16998 & ~n17005;
  assign n17613 = n17004 & n17612;
  assign n17614 = po7  & n17613;
  assign n17615 = po7  & n17612;
  assign n17616 = ~n17004 & ~n17615;
  assign n17617 = ~n17614 & ~n17616;
  assign n17618 = ~po48  & ~n17601;
  assign n17619 = ~n17609 & n17618;
  assign n17620 = ~n17617 & ~n17619;
  assign n17621 = ~n17611 & ~n17620;
  assign n17622 = po49  & ~n17621;
  assign n17623 = ~n17008 & ~n17016;
  assign n17624 = n17014 & n17623;
  assign n17625 = po7  & n17624;
  assign n17626 = po7  & n17623;
  assign n17627 = ~n17014 & ~n17626;
  assign n17628 = ~n17625 & ~n17627;
  assign n17629 = ~po49  & n17621;
  assign n17630 = ~n17628 & ~n17629;
  assign n17631 = ~n17622 & ~n17630;
  assign n17632 = po50  & ~n17631;
  assign n17633 = ~n17019 & ~n17026;
  assign n17634 = n17025 & n17633;
  assign n17635 = po7  & n17634;
  assign n17636 = po7  & n17633;
  assign n17637 = ~n17025 & ~n17636;
  assign n17638 = ~n17635 & ~n17637;
  assign n17639 = ~po50  & ~n17622;
  assign n17640 = ~n17630 & n17639;
  assign n17641 = ~n17638 & ~n17640;
  assign n17642 = ~n17632 & ~n17641;
  assign n17643 = po51  & ~n17642;
  assign n17644 = ~n17029 & ~n17037;
  assign n17645 = n17035 & n17644;
  assign n17646 = po7  & n17645;
  assign n17647 = po7  & n17644;
  assign n17648 = ~n17035 & ~n17647;
  assign n17649 = ~n17646 & ~n17648;
  assign n17650 = ~po51  & n17642;
  assign n17651 = ~n17649 & ~n17650;
  assign n17652 = ~n17643 & ~n17651;
  assign n17653 = po52  & ~n17652;
  assign n17654 = ~n17040 & ~n17047;
  assign n17655 = n17046 & n17654;
  assign n17656 = po7  & n17655;
  assign n17657 = po7  & n17654;
  assign n17658 = ~n17046 & ~n17657;
  assign n17659 = ~n17656 & ~n17658;
  assign n17660 = ~po52  & ~n17643;
  assign n17661 = ~n17651 & n17660;
  assign n17662 = ~n17659 & ~n17661;
  assign n17663 = ~n17653 & ~n17662;
  assign n17664 = po53  & ~n17663;
  assign n17665 = ~n17050 & ~n17058;
  assign n17666 = n17056 & n17665;
  assign n17667 = po7  & n17666;
  assign n17668 = po7  & n17665;
  assign n17669 = ~n17056 & ~n17668;
  assign n17670 = ~n17667 & ~n17669;
  assign n17671 = ~po53  & n17663;
  assign n17672 = ~n17670 & ~n17671;
  assign n17673 = ~n17664 & ~n17672;
  assign n17674 = po54  & ~n17673;
  assign n17675 = ~n17061 & ~n17068;
  assign n17676 = n17067 & n17675;
  assign n17677 = po7  & n17676;
  assign n17678 = po7  & n17675;
  assign n17679 = ~n17067 & ~n17678;
  assign n17680 = ~n17677 & ~n17679;
  assign n17681 = ~po54  & ~n17664;
  assign n17682 = ~n17672 & n17681;
  assign n17683 = ~n17680 & ~n17682;
  assign n17684 = ~n17674 & ~n17683;
  assign n17685 = po55  & ~n17684;
  assign n17686 = ~n17071 & ~n17079;
  assign n17687 = n17077 & n17686;
  assign n17688 = po7  & n17687;
  assign n17689 = po7  & n17686;
  assign n17690 = ~n17077 & ~n17689;
  assign n17691 = ~n17688 & ~n17690;
  assign n17692 = ~po55  & n17684;
  assign n17693 = ~n17691 & ~n17692;
  assign n17694 = ~n17685 & ~n17693;
  assign n17695 = po56  & ~n17694;
  assign n17696 = ~n17082 & ~n17089;
  assign n17697 = n17088 & n17696;
  assign n17698 = po7  & n17697;
  assign n17699 = po7  & n17696;
  assign n17700 = ~n17088 & ~n17699;
  assign n17701 = ~n17698 & ~n17700;
  assign n17702 = ~po56  & ~n17685;
  assign n17703 = ~n17693 & n17702;
  assign n17704 = ~n17701 & ~n17703;
  assign n17705 = ~n17695 & ~n17704;
  assign n17706 = po57  & ~n17705;
  assign n17707 = ~n17092 & ~n17100;
  assign n17708 = n17098 & n17707;
  assign n17709 = po7  & n17708;
  assign n17710 = po7  & n17707;
  assign n17711 = ~n17098 & ~n17710;
  assign n17712 = ~n17709 & ~n17711;
  assign n17713 = ~po57  & n17705;
  assign n17714 = ~n17712 & ~n17713;
  assign n17715 = ~n17706 & ~n17714;
  assign n17716 = po58  & ~n17715;
  assign n17717 = ~po58  & ~n17706;
  assign n17718 = ~n17714 & n17717;
  assign n17719 = ~n17103 & ~n17110;
  assign n17720 = n17109 & n17719;
  assign n17721 = po7  & n17720;
  assign n17722 = po7  & n17719;
  assign n17723 = ~n17109 & ~n17722;
  assign n17724 = ~n17721 & ~n17723;
  assign n17725 = ~n17718 & ~n17724;
  assign n17726 = ~n17716 & ~n17725;
  assign n17727 = po59  & ~n17726;
  assign n17728 = ~n17113 & ~n17121;
  assign n17729 = n17119 & n17728;
  assign n17730 = po7  & n17729;
  assign n17731 = po7  & n17728;
  assign n17732 = ~n17119 & ~n17731;
  assign n17733 = ~n17730 & ~n17732;
  assign n17734 = ~po59  & n17726;
  assign n17735 = ~n17733 & ~n17734;
  assign n17736 = ~n17727 & ~n17735;
  assign n17737 = po60  & ~n17736;
  assign n17738 = ~n17124 & ~n17131;
  assign n17739 = n17130 & n17738;
  assign n17740 = po7  & n17739;
  assign n17741 = po7  & n17738;
  assign n17742 = ~n17130 & ~n17741;
  assign n17743 = ~n17740 & ~n17742;
  assign n17744 = ~po60  & ~n17727;
  assign n17745 = ~n17735 & n17744;
  assign n17746 = ~n17743 & ~n17745;
  assign n17747 = ~n17737 & ~n17746;
  assign n17748 = po61  & ~n17747;
  assign n17749 = ~n17134 & ~n17142;
  assign n17750 = n17140 & n17749;
  assign n17751 = po7  & n17750;
  assign n17752 = po7  & n17749;
  assign n17753 = ~n17140 & ~n17752;
  assign n17754 = ~n17751 & ~n17753;
  assign n17755 = ~po61  & n17747;
  assign n17756 = ~n17754 & ~n17755;
  assign n17757 = ~n17748 & ~n17756;
  assign n17758 = po62  & ~n17757;
  assign n17759 = ~n17145 & ~n17152;
  assign n17760 = n17151 & n17759;
  assign n17761 = po7  & n17760;
  assign n17762 = po7  & n17759;
  assign n17763 = ~n17151 & ~n17762;
  assign n17764 = ~n17761 & ~n17763;
  assign n17765 = ~po62  & ~n17748;
  assign n17766 = ~n17756 & n17765;
  assign n17767 = ~n17764 & ~n17766;
  assign n17768 = ~n17758 & ~n17767;
  assign n17769 = ~n17155 & ~n17163;
  assign n17770 = po7  & n17769;
  assign n17771 = ~n17161 & ~n17770;
  assign n17772 = n17161 & n17770;
  assign n17773 = ~n17771 & ~n17772;
  assign n17774 = ~n17165 & ~n17170;
  assign n17775 = po7  & n17774;
  assign n17776 = ~n17183 & ~n17775;
  assign n17777 = ~n17773 & n17776;
  assign n17778 = ~n17768 & n17777;
  assign n17779 = ~po63  & ~n17778;
  assign n17780 = ~n17170 & po7 ;
  assign n17781 = n17165 & ~n17780;
  assign n17782 = po63  & ~n17774;
  assign n17783 = ~n17781 & n17782;
  assign n17784 = n17170 & ~po7 ;
  assign n17785 = ~n17783 & ~n17784;
  assign n17786 = n17768 & n17773;
  assign n17787 = n17785 & ~n17786;
  assign po6  = n17779 | ~n17787;
  assign n17789 = pi12  & po6 ;
  assign n17790 = ~pi10  & ~pi11 ;
  assign n17791 = ~pi12  & n17790;
  assign n17792 = ~n17789 & ~n17791;
  assign n17793 = po7  & ~n17792;
  assign n17794 = n17182 & ~n17791;
  assign n17795 = ~n17183 & n17794;
  assign n17796 = ~n17176 & n17795;
  assign n17797 = ~n17789 & n17796;
  assign n17798 = ~pi12  & po6 ;
  assign n17799 = pi13  & ~n17798;
  assign n17800 = n17187 & po6 ;
  assign n17801 = ~n17799 & ~n17800;
  assign n17802 = ~n17797 & n17801;
  assign n17803 = ~n17793 & ~n17802;
  assign n17804 = po8  & ~n17803;
  assign n17805 = ~po8  & ~n17793;
  assign n17806 = ~n17802 & n17805;
  assign n17807 = po7  & n17785;
  assign n17808 = ~n17786 & n17807;
  assign n17809 = ~n17779 & n17808;
  assign n17810 = ~n17800 & ~n17809;
  assign n17811 = pi14  & ~n17810;
  assign n17812 = ~pi14  & n17810;
  assign n17813 = ~n17811 & ~n17812;
  assign n17814 = ~n17806 & ~n17813;
  assign n17815 = ~n17804 & ~n17814;
  assign n17816 = po9  & ~n17815;
  assign n17817 = ~n17190 & ~n17194;
  assign n17818 = ~n17198 & n17817;
  assign n17819 = po6  & n17818;
  assign n17820 = po6  & n17817;
  assign n17821 = n17198 & ~n17820;
  assign n17822 = ~n17819 & ~n17821;
  assign n17823 = ~po9  & n17815;
  assign n17824 = ~n17822 & ~n17823;
  assign n17825 = ~n17816 & ~n17824;
  assign n17826 = po10  & ~n17825;
  assign n17827 = ~n17201 & ~n17209;
  assign n17828 = n17208 & n17827;
  assign n17829 = po6  & n17828;
  assign n17830 = po6  & n17827;
  assign n17831 = ~n17208 & ~n17830;
  assign n17832 = ~n17829 & ~n17831;
  assign n17833 = ~po10  & ~n17816;
  assign n17834 = ~n17824 & n17833;
  assign n17835 = ~n17832 & ~n17834;
  assign n17836 = ~n17826 & ~n17835;
  assign n17837 = po11  & ~n17836;
  assign n17838 = ~n17212 & ~n17220;
  assign n17839 = n17218 & n17838;
  assign n17840 = po6  & n17839;
  assign n17841 = po6  & n17838;
  assign n17842 = ~n17218 & ~n17841;
  assign n17843 = ~n17840 & ~n17842;
  assign n17844 = ~po11  & n17836;
  assign n17845 = ~n17843 & ~n17844;
  assign n17846 = ~n17837 & ~n17845;
  assign n17847 = po12  & ~n17846;
  assign n17848 = ~n17223 & ~n17230;
  assign n17849 = n17229 & n17848;
  assign n17850 = po6  & n17849;
  assign n17851 = po6  & n17848;
  assign n17852 = ~n17229 & ~n17851;
  assign n17853 = ~n17850 & ~n17852;
  assign n17854 = ~po12  & ~n17837;
  assign n17855 = ~n17845 & n17854;
  assign n17856 = ~n17853 & ~n17855;
  assign n17857 = ~n17847 & ~n17856;
  assign n17858 = po13  & ~n17857;
  assign n17859 = ~n17233 & ~n17241;
  assign n17860 = n17239 & n17859;
  assign n17861 = po6  & n17860;
  assign n17862 = po6  & n17859;
  assign n17863 = ~n17239 & ~n17862;
  assign n17864 = ~n17861 & ~n17863;
  assign n17865 = ~po13  & n17857;
  assign n17866 = ~n17864 & ~n17865;
  assign n17867 = ~n17858 & ~n17866;
  assign n17868 = po14  & ~n17867;
  assign n17869 = ~n17244 & ~n17251;
  assign n17870 = n17250 & n17869;
  assign n17871 = po6  & n17870;
  assign n17872 = po6  & n17869;
  assign n17873 = ~n17250 & ~n17872;
  assign n17874 = ~n17871 & ~n17873;
  assign n17875 = ~po14  & ~n17858;
  assign n17876 = ~n17866 & n17875;
  assign n17877 = ~n17874 & ~n17876;
  assign n17878 = ~n17868 & ~n17877;
  assign n17879 = po15  & ~n17878;
  assign n17880 = ~n17254 & ~n17262;
  assign n17881 = n17260 & n17880;
  assign n17882 = po6  & n17881;
  assign n17883 = po6  & n17880;
  assign n17884 = ~n17260 & ~n17883;
  assign n17885 = ~n17882 & ~n17884;
  assign n17886 = ~po15  & n17878;
  assign n17887 = ~n17885 & ~n17886;
  assign n17888 = ~n17879 & ~n17887;
  assign n17889 = po16  & ~n17888;
  assign n17890 = ~n17265 & ~n17272;
  assign n17891 = n17271 & n17890;
  assign n17892 = po6  & n17891;
  assign n17893 = po6  & n17890;
  assign n17894 = ~n17271 & ~n17893;
  assign n17895 = ~n17892 & ~n17894;
  assign n17896 = ~po16  & ~n17879;
  assign n17897 = ~n17887 & n17896;
  assign n17898 = ~n17895 & ~n17897;
  assign n17899 = ~n17889 & ~n17898;
  assign n17900 = po17  & ~n17899;
  assign n17901 = ~n17275 & ~n17283;
  assign n17902 = n17281 & n17901;
  assign n17903 = po6  & n17902;
  assign n17904 = po6  & n17901;
  assign n17905 = ~n17281 & ~n17904;
  assign n17906 = ~n17903 & ~n17905;
  assign n17907 = ~po17  & n17899;
  assign n17908 = ~n17906 & ~n17907;
  assign n17909 = ~n17900 & ~n17908;
  assign n17910 = po18  & ~n17909;
  assign n17911 = ~n17286 & ~n17293;
  assign n17912 = n17292 & n17911;
  assign n17913 = po6  & n17912;
  assign n17914 = po6  & n17911;
  assign n17915 = ~n17292 & ~n17914;
  assign n17916 = ~n17913 & ~n17915;
  assign n17917 = ~po18  & ~n17900;
  assign n17918 = ~n17908 & n17917;
  assign n17919 = ~n17916 & ~n17918;
  assign n17920 = ~n17910 & ~n17919;
  assign n17921 = po19  & ~n17920;
  assign n17922 = ~n17296 & ~n17304;
  assign n17923 = n17302 & n17922;
  assign n17924 = po6  & n17923;
  assign n17925 = po6  & n17922;
  assign n17926 = ~n17302 & ~n17925;
  assign n17927 = ~n17924 & ~n17926;
  assign n17928 = ~po19  & n17920;
  assign n17929 = ~n17927 & ~n17928;
  assign n17930 = ~n17921 & ~n17929;
  assign n17931 = po20  & ~n17930;
  assign n17932 = ~n17307 & ~n17314;
  assign n17933 = n17313 & n17932;
  assign n17934 = po6  & n17933;
  assign n17935 = po6  & n17932;
  assign n17936 = ~n17313 & ~n17935;
  assign n17937 = ~n17934 & ~n17936;
  assign n17938 = ~po20  & ~n17921;
  assign n17939 = ~n17929 & n17938;
  assign n17940 = ~n17937 & ~n17939;
  assign n17941 = ~n17931 & ~n17940;
  assign n17942 = po21  & ~n17941;
  assign n17943 = ~n17317 & ~n17325;
  assign n17944 = n17323 & n17943;
  assign n17945 = po6  & n17944;
  assign n17946 = po6  & n17943;
  assign n17947 = ~n17323 & ~n17946;
  assign n17948 = ~n17945 & ~n17947;
  assign n17949 = ~po21  & n17941;
  assign n17950 = ~n17948 & ~n17949;
  assign n17951 = ~n17942 & ~n17950;
  assign n17952 = po22  & ~n17951;
  assign n17953 = ~n17328 & ~n17335;
  assign n17954 = n17334 & n17953;
  assign n17955 = po6  & n17954;
  assign n17956 = po6  & n17953;
  assign n17957 = ~n17334 & ~n17956;
  assign n17958 = ~n17955 & ~n17957;
  assign n17959 = ~po22  & ~n17942;
  assign n17960 = ~n17950 & n17959;
  assign n17961 = ~n17958 & ~n17960;
  assign n17962 = ~n17952 & ~n17961;
  assign n17963 = po23  & ~n17962;
  assign n17964 = ~n17338 & ~n17346;
  assign n17965 = n17344 & n17964;
  assign n17966 = po6  & n17965;
  assign n17967 = po6  & n17964;
  assign n17968 = ~n17344 & ~n17967;
  assign n17969 = ~n17966 & ~n17968;
  assign n17970 = ~po23  & n17962;
  assign n17971 = ~n17969 & ~n17970;
  assign n17972 = ~n17963 & ~n17971;
  assign n17973 = po24  & ~n17972;
  assign n17974 = ~n17349 & ~n17356;
  assign n17975 = n17355 & n17974;
  assign n17976 = po6  & n17975;
  assign n17977 = po6  & n17974;
  assign n17978 = ~n17355 & ~n17977;
  assign n17979 = ~n17976 & ~n17978;
  assign n17980 = ~po24  & ~n17963;
  assign n17981 = ~n17971 & n17980;
  assign n17982 = ~n17979 & ~n17981;
  assign n17983 = ~n17973 & ~n17982;
  assign n17984 = po25  & ~n17983;
  assign n17985 = ~n17359 & ~n17367;
  assign n17986 = n17365 & n17985;
  assign n17987 = po6  & n17986;
  assign n17988 = po6  & n17985;
  assign n17989 = ~n17365 & ~n17988;
  assign n17990 = ~n17987 & ~n17989;
  assign n17991 = ~po25  & n17983;
  assign n17992 = ~n17990 & ~n17991;
  assign n17993 = ~n17984 & ~n17992;
  assign n17994 = po26  & ~n17993;
  assign n17995 = ~n17370 & ~n17377;
  assign n17996 = n17376 & n17995;
  assign n17997 = po6  & n17996;
  assign n17998 = po6  & n17995;
  assign n17999 = ~n17376 & ~n17998;
  assign n18000 = ~n17997 & ~n17999;
  assign n18001 = ~po26  & ~n17984;
  assign n18002 = ~n17992 & n18001;
  assign n18003 = ~n18000 & ~n18002;
  assign n18004 = ~n17994 & ~n18003;
  assign n18005 = po27  & ~n18004;
  assign n18006 = ~n17380 & ~n17388;
  assign n18007 = n17386 & n18006;
  assign n18008 = po6  & n18007;
  assign n18009 = po6  & n18006;
  assign n18010 = ~n17386 & ~n18009;
  assign n18011 = ~n18008 & ~n18010;
  assign n18012 = ~po27  & n18004;
  assign n18013 = ~n18011 & ~n18012;
  assign n18014 = ~n18005 & ~n18013;
  assign n18015 = po28  & ~n18014;
  assign n18016 = ~n17391 & ~n17398;
  assign n18017 = n17397 & n18016;
  assign n18018 = po6  & n18017;
  assign n18019 = po6  & n18016;
  assign n18020 = ~n17397 & ~n18019;
  assign n18021 = ~n18018 & ~n18020;
  assign n18022 = ~po28  & ~n18005;
  assign n18023 = ~n18013 & n18022;
  assign n18024 = ~n18021 & ~n18023;
  assign n18025 = ~n18015 & ~n18024;
  assign n18026 = po29  & ~n18025;
  assign n18027 = ~n17401 & ~n17409;
  assign n18028 = n17407 & n18027;
  assign n18029 = po6  & n18028;
  assign n18030 = po6  & n18027;
  assign n18031 = ~n17407 & ~n18030;
  assign n18032 = ~n18029 & ~n18031;
  assign n18033 = ~po29  & n18025;
  assign n18034 = ~n18032 & ~n18033;
  assign n18035 = ~n18026 & ~n18034;
  assign n18036 = po30  & ~n18035;
  assign n18037 = ~n17412 & ~n17419;
  assign n18038 = n17418 & n18037;
  assign n18039 = po6  & n18038;
  assign n18040 = po6  & n18037;
  assign n18041 = ~n17418 & ~n18040;
  assign n18042 = ~n18039 & ~n18041;
  assign n18043 = ~po30  & ~n18026;
  assign n18044 = ~n18034 & n18043;
  assign n18045 = ~n18042 & ~n18044;
  assign n18046 = ~n18036 & ~n18045;
  assign n18047 = po31  & ~n18046;
  assign n18048 = ~n17422 & ~n17430;
  assign n18049 = n17428 & n18048;
  assign n18050 = po6  & n18049;
  assign n18051 = po6  & n18048;
  assign n18052 = ~n17428 & ~n18051;
  assign n18053 = ~n18050 & ~n18052;
  assign n18054 = ~po31  & n18046;
  assign n18055 = ~n18053 & ~n18054;
  assign n18056 = ~n18047 & ~n18055;
  assign n18057 = po32  & ~n18056;
  assign n18058 = ~n17433 & ~n17440;
  assign n18059 = n17439 & n18058;
  assign n18060 = po6  & n18059;
  assign n18061 = po6  & n18058;
  assign n18062 = ~n17439 & ~n18061;
  assign n18063 = ~n18060 & ~n18062;
  assign n18064 = ~po32  & ~n18047;
  assign n18065 = ~n18055 & n18064;
  assign n18066 = ~n18063 & ~n18065;
  assign n18067 = ~n18057 & ~n18066;
  assign n18068 = po33  & ~n18067;
  assign n18069 = ~n17443 & ~n17451;
  assign n18070 = n17449 & n18069;
  assign n18071 = po6  & n18070;
  assign n18072 = po6  & n18069;
  assign n18073 = ~n17449 & ~n18072;
  assign n18074 = ~n18071 & ~n18073;
  assign n18075 = ~po33  & n18067;
  assign n18076 = ~n18074 & ~n18075;
  assign n18077 = ~n18068 & ~n18076;
  assign n18078 = po34  & ~n18077;
  assign n18079 = ~n17454 & ~n17461;
  assign n18080 = n17460 & n18079;
  assign n18081 = po6  & n18080;
  assign n18082 = po6  & n18079;
  assign n18083 = ~n17460 & ~n18082;
  assign n18084 = ~n18081 & ~n18083;
  assign n18085 = ~po34  & ~n18068;
  assign n18086 = ~n18076 & n18085;
  assign n18087 = ~n18084 & ~n18086;
  assign n18088 = ~n18078 & ~n18087;
  assign n18089 = po35  & ~n18088;
  assign n18090 = ~n17464 & ~n17472;
  assign n18091 = n17470 & n18090;
  assign n18092 = po6  & n18091;
  assign n18093 = po6  & n18090;
  assign n18094 = ~n17470 & ~n18093;
  assign n18095 = ~n18092 & ~n18094;
  assign n18096 = ~po35  & n18088;
  assign n18097 = ~n18095 & ~n18096;
  assign n18098 = ~n18089 & ~n18097;
  assign n18099 = po36  & ~n18098;
  assign n18100 = ~n17475 & ~n17482;
  assign n18101 = n17481 & n18100;
  assign n18102 = po6  & n18101;
  assign n18103 = po6  & n18100;
  assign n18104 = ~n17481 & ~n18103;
  assign n18105 = ~n18102 & ~n18104;
  assign n18106 = ~po36  & ~n18089;
  assign n18107 = ~n18097 & n18106;
  assign n18108 = ~n18105 & ~n18107;
  assign n18109 = ~n18099 & ~n18108;
  assign n18110 = po37  & ~n18109;
  assign n18111 = ~n17485 & ~n17493;
  assign n18112 = n17491 & n18111;
  assign n18113 = po6  & n18112;
  assign n18114 = po6  & n18111;
  assign n18115 = ~n17491 & ~n18114;
  assign n18116 = ~n18113 & ~n18115;
  assign n18117 = ~po37  & n18109;
  assign n18118 = ~n18116 & ~n18117;
  assign n18119 = ~n18110 & ~n18118;
  assign n18120 = po38  & ~n18119;
  assign n18121 = ~n17496 & ~n17503;
  assign n18122 = n17502 & n18121;
  assign n18123 = po6  & n18122;
  assign n18124 = po6  & n18121;
  assign n18125 = ~n17502 & ~n18124;
  assign n18126 = ~n18123 & ~n18125;
  assign n18127 = ~po38  & ~n18110;
  assign n18128 = ~n18118 & n18127;
  assign n18129 = ~n18126 & ~n18128;
  assign n18130 = ~n18120 & ~n18129;
  assign n18131 = po39  & ~n18130;
  assign n18132 = ~n17506 & ~n17514;
  assign n18133 = n17512 & n18132;
  assign n18134 = po6  & n18133;
  assign n18135 = po6  & n18132;
  assign n18136 = ~n17512 & ~n18135;
  assign n18137 = ~n18134 & ~n18136;
  assign n18138 = ~po39  & n18130;
  assign n18139 = ~n18137 & ~n18138;
  assign n18140 = ~n18131 & ~n18139;
  assign n18141 = po40  & ~n18140;
  assign n18142 = ~n17517 & ~n17524;
  assign n18143 = n17523 & n18142;
  assign n18144 = po6  & n18143;
  assign n18145 = po6  & n18142;
  assign n18146 = ~n17523 & ~n18145;
  assign n18147 = ~n18144 & ~n18146;
  assign n18148 = ~po40  & ~n18131;
  assign n18149 = ~n18139 & n18148;
  assign n18150 = ~n18147 & ~n18149;
  assign n18151 = ~n18141 & ~n18150;
  assign n18152 = po41  & ~n18151;
  assign n18153 = ~n17527 & ~n17535;
  assign n18154 = n17533 & n18153;
  assign n18155 = po6  & n18154;
  assign n18156 = po6  & n18153;
  assign n18157 = ~n17533 & ~n18156;
  assign n18158 = ~n18155 & ~n18157;
  assign n18159 = ~po41  & n18151;
  assign n18160 = ~n18158 & ~n18159;
  assign n18161 = ~n18152 & ~n18160;
  assign n18162 = po42  & ~n18161;
  assign n18163 = ~n17538 & ~n17545;
  assign n18164 = n17544 & n18163;
  assign n18165 = po6  & n18164;
  assign n18166 = po6  & n18163;
  assign n18167 = ~n17544 & ~n18166;
  assign n18168 = ~n18165 & ~n18167;
  assign n18169 = ~po42  & ~n18152;
  assign n18170 = ~n18160 & n18169;
  assign n18171 = ~n18168 & ~n18170;
  assign n18172 = ~n18162 & ~n18171;
  assign n18173 = po43  & ~n18172;
  assign n18174 = ~n17548 & ~n17556;
  assign n18175 = n17554 & n18174;
  assign n18176 = po6  & n18175;
  assign n18177 = po6  & n18174;
  assign n18178 = ~n17554 & ~n18177;
  assign n18179 = ~n18176 & ~n18178;
  assign n18180 = ~po43  & n18172;
  assign n18181 = ~n18179 & ~n18180;
  assign n18182 = ~n18173 & ~n18181;
  assign n18183 = po44  & ~n18182;
  assign n18184 = ~n17559 & ~n17566;
  assign n18185 = n17565 & n18184;
  assign n18186 = po6  & n18185;
  assign n18187 = po6  & n18184;
  assign n18188 = ~n17565 & ~n18187;
  assign n18189 = ~n18186 & ~n18188;
  assign n18190 = ~po44  & ~n18173;
  assign n18191 = ~n18181 & n18190;
  assign n18192 = ~n18189 & ~n18191;
  assign n18193 = ~n18183 & ~n18192;
  assign n18194 = po45  & ~n18193;
  assign n18195 = ~n17569 & ~n17577;
  assign n18196 = n17575 & n18195;
  assign n18197 = po6  & n18196;
  assign n18198 = po6  & n18195;
  assign n18199 = ~n17575 & ~n18198;
  assign n18200 = ~n18197 & ~n18199;
  assign n18201 = ~po45  & n18193;
  assign n18202 = ~n18200 & ~n18201;
  assign n18203 = ~n18194 & ~n18202;
  assign n18204 = po46  & ~n18203;
  assign n18205 = ~n17580 & ~n17587;
  assign n18206 = n17586 & n18205;
  assign n18207 = po6  & n18206;
  assign n18208 = po6  & n18205;
  assign n18209 = ~n17586 & ~n18208;
  assign n18210 = ~n18207 & ~n18209;
  assign n18211 = ~po46  & ~n18194;
  assign n18212 = ~n18202 & n18211;
  assign n18213 = ~n18210 & ~n18212;
  assign n18214 = ~n18204 & ~n18213;
  assign n18215 = po47  & ~n18214;
  assign n18216 = ~n17590 & ~n17598;
  assign n18217 = n17596 & n18216;
  assign n18218 = po6  & n18217;
  assign n18219 = po6  & n18216;
  assign n18220 = ~n17596 & ~n18219;
  assign n18221 = ~n18218 & ~n18220;
  assign n18222 = ~po47  & n18214;
  assign n18223 = ~n18221 & ~n18222;
  assign n18224 = ~n18215 & ~n18223;
  assign n18225 = po48  & ~n18224;
  assign n18226 = ~n17601 & ~n17608;
  assign n18227 = n17607 & n18226;
  assign n18228 = po6  & n18227;
  assign n18229 = po6  & n18226;
  assign n18230 = ~n17607 & ~n18229;
  assign n18231 = ~n18228 & ~n18230;
  assign n18232 = ~po48  & ~n18215;
  assign n18233 = ~n18223 & n18232;
  assign n18234 = ~n18231 & ~n18233;
  assign n18235 = ~n18225 & ~n18234;
  assign n18236 = po49  & ~n18235;
  assign n18237 = ~n17611 & ~n17619;
  assign n18238 = n17617 & n18237;
  assign n18239 = po6  & n18238;
  assign n18240 = po6  & n18237;
  assign n18241 = ~n17617 & ~n18240;
  assign n18242 = ~n18239 & ~n18241;
  assign n18243 = ~po49  & n18235;
  assign n18244 = ~n18242 & ~n18243;
  assign n18245 = ~n18236 & ~n18244;
  assign n18246 = po50  & ~n18245;
  assign n18247 = ~n17622 & ~n17629;
  assign n18248 = n17628 & n18247;
  assign n18249 = po6  & n18248;
  assign n18250 = po6  & n18247;
  assign n18251 = ~n17628 & ~n18250;
  assign n18252 = ~n18249 & ~n18251;
  assign n18253 = ~po50  & ~n18236;
  assign n18254 = ~n18244 & n18253;
  assign n18255 = ~n18252 & ~n18254;
  assign n18256 = ~n18246 & ~n18255;
  assign n18257 = po51  & ~n18256;
  assign n18258 = ~n17632 & ~n17640;
  assign n18259 = n17638 & n18258;
  assign n18260 = po6  & n18259;
  assign n18261 = po6  & n18258;
  assign n18262 = ~n17638 & ~n18261;
  assign n18263 = ~n18260 & ~n18262;
  assign n18264 = ~po51  & n18256;
  assign n18265 = ~n18263 & ~n18264;
  assign n18266 = ~n18257 & ~n18265;
  assign n18267 = po52  & ~n18266;
  assign n18268 = ~n17643 & ~n17650;
  assign n18269 = n17649 & n18268;
  assign n18270 = po6  & n18269;
  assign n18271 = po6  & n18268;
  assign n18272 = ~n17649 & ~n18271;
  assign n18273 = ~n18270 & ~n18272;
  assign n18274 = ~po52  & ~n18257;
  assign n18275 = ~n18265 & n18274;
  assign n18276 = ~n18273 & ~n18275;
  assign n18277 = ~n18267 & ~n18276;
  assign n18278 = po53  & ~n18277;
  assign n18279 = ~n17653 & ~n17661;
  assign n18280 = n17659 & n18279;
  assign n18281 = po6  & n18280;
  assign n18282 = po6  & n18279;
  assign n18283 = ~n17659 & ~n18282;
  assign n18284 = ~n18281 & ~n18283;
  assign n18285 = ~po53  & n18277;
  assign n18286 = ~n18284 & ~n18285;
  assign n18287 = ~n18278 & ~n18286;
  assign n18288 = po54  & ~n18287;
  assign n18289 = ~n17664 & ~n17671;
  assign n18290 = n17670 & n18289;
  assign n18291 = po6  & n18290;
  assign n18292 = po6  & n18289;
  assign n18293 = ~n17670 & ~n18292;
  assign n18294 = ~n18291 & ~n18293;
  assign n18295 = ~po54  & ~n18278;
  assign n18296 = ~n18286 & n18295;
  assign n18297 = ~n18294 & ~n18296;
  assign n18298 = ~n18288 & ~n18297;
  assign n18299 = po55  & ~n18298;
  assign n18300 = ~n17674 & ~n17682;
  assign n18301 = n17680 & n18300;
  assign n18302 = po6  & n18301;
  assign n18303 = po6  & n18300;
  assign n18304 = ~n17680 & ~n18303;
  assign n18305 = ~n18302 & ~n18304;
  assign n18306 = ~po55  & n18298;
  assign n18307 = ~n18305 & ~n18306;
  assign n18308 = ~n18299 & ~n18307;
  assign n18309 = po56  & ~n18308;
  assign n18310 = ~n17685 & ~n17692;
  assign n18311 = n17691 & n18310;
  assign n18312 = po6  & n18311;
  assign n18313 = po6  & n18310;
  assign n18314 = ~n17691 & ~n18313;
  assign n18315 = ~n18312 & ~n18314;
  assign n18316 = ~po56  & ~n18299;
  assign n18317 = ~n18307 & n18316;
  assign n18318 = ~n18315 & ~n18317;
  assign n18319 = ~n18309 & ~n18318;
  assign n18320 = po57  & ~n18319;
  assign n18321 = ~n17695 & ~n17703;
  assign n18322 = n17701 & n18321;
  assign n18323 = po6  & n18322;
  assign n18324 = po6  & n18321;
  assign n18325 = ~n17701 & ~n18324;
  assign n18326 = ~n18323 & ~n18325;
  assign n18327 = ~po57  & n18319;
  assign n18328 = ~n18326 & ~n18327;
  assign n18329 = ~n18320 & ~n18328;
  assign n18330 = po58  & ~n18329;
  assign n18331 = ~n17706 & ~n17713;
  assign n18332 = n17712 & n18331;
  assign n18333 = po6  & n18332;
  assign n18334 = po6  & n18331;
  assign n18335 = ~n17712 & ~n18334;
  assign n18336 = ~n18333 & ~n18335;
  assign n18337 = ~po58  & ~n18320;
  assign n18338 = ~n18328 & n18337;
  assign n18339 = ~n18336 & ~n18338;
  assign n18340 = ~n18330 & ~n18339;
  assign n18341 = po59  & ~n18340;
  assign n18342 = ~n17716 & ~n17718;
  assign n18343 = n17724 & n18342;
  assign n18344 = po6  & n18343;
  assign n18345 = po6  & n18342;
  assign n18346 = ~n17724 & ~n18345;
  assign n18347 = ~n18344 & ~n18346;
  assign n18348 = ~po59  & n18340;
  assign n18349 = ~n18347 & ~n18348;
  assign n18350 = ~n18341 & ~n18349;
  assign n18351 = po60  & ~n18350;
  assign n18352 = ~n17727 & ~n17734;
  assign n18353 = n17733 & n18352;
  assign n18354 = po6  & n18353;
  assign n18355 = po6  & n18352;
  assign n18356 = ~n17733 & ~n18355;
  assign n18357 = ~n18354 & ~n18356;
  assign n18358 = ~po60  & ~n18341;
  assign n18359 = ~n18349 & n18358;
  assign n18360 = ~n18357 & ~n18359;
  assign n18361 = ~n18351 & ~n18360;
  assign n18362 = po61  & ~n18361;
  assign n18363 = ~n17737 & ~n17745;
  assign n18364 = n17743 & n18363;
  assign n18365 = po6  & n18364;
  assign n18366 = po6  & n18363;
  assign n18367 = ~n17743 & ~n18366;
  assign n18368 = ~n18365 & ~n18367;
  assign n18369 = ~po61  & n18361;
  assign n18370 = ~n18368 & ~n18369;
  assign n18371 = ~n18362 & ~n18370;
  assign n18372 = po62  & ~n18371;
  assign n18373 = ~n17748 & ~n17755;
  assign n18374 = n17754 & n18373;
  assign n18375 = po6  & n18374;
  assign n18376 = po6  & n18373;
  assign n18377 = ~n17754 & ~n18376;
  assign n18378 = ~n18375 & ~n18377;
  assign n18379 = ~po62  & ~n18362;
  assign n18380 = ~n18370 & n18379;
  assign n18381 = ~n18378 & ~n18380;
  assign n18382 = ~n18372 & ~n18381;
  assign n18383 = ~n17758 & ~n17766;
  assign n18384 = po6  & n18383;
  assign n18385 = ~n17764 & ~n18384;
  assign n18386 = n17764 & n18384;
  assign n18387 = ~n18385 & ~n18386;
  assign n18388 = ~n17768 & ~n17773;
  assign n18389 = po6  & n18388;
  assign n18390 = ~n17786 & ~n18389;
  assign n18391 = ~n18387 & n18390;
  assign n18392 = ~n18382 & n18391;
  assign n18393 = ~po63  & ~n18392;
  assign n18394 = ~n17773 & po6 ;
  assign n18395 = n17768 & ~n18394;
  assign n18396 = po63  & ~n18388;
  assign n18397 = ~n18395 & n18396;
  assign n18398 = n18382 & n18387;
  assign n18399 = ~n18397 & ~n18398;
  assign po5  = n18393 | ~n18399;
  assign n18401 = pi10  & po5 ;
  assign n18402 = ~pi8  & ~pi9 ;
  assign n18403 = ~pi10  & n18402;
  assign n18404 = ~n18401 & ~n18403;
  assign n18405 = po6  & ~n18404;
  assign n18406 = n17785 & ~n18403;
  assign n18407 = ~n17786 & n18406;
  assign n18408 = ~n17779 & n18407;
  assign n18409 = ~n18401 & n18408;
  assign n18410 = ~pi10  & po5 ;
  assign n18411 = pi11  & ~n18410;
  assign n18412 = n17790 & po5 ;
  assign n18413 = ~n18411 & ~n18412;
  assign n18414 = ~n18409 & n18413;
  assign n18415 = ~n18405 & ~n18414;
  assign n18416 = po7  & ~n18415;
  assign n18417 = po6  & ~n18397;
  assign n18418 = ~n18398 & n18417;
  assign n18419 = ~n18393 & n18418;
  assign n18420 = ~n18412 & ~n18419;
  assign n18421 = pi12  & ~n18420;
  assign n18422 = ~pi12  & n18420;
  assign n18423 = ~n18421 & ~n18422;
  assign n18424 = ~po7  & n18415;
  assign n18425 = ~n18423 & ~n18424;
  assign n18426 = ~n18416 & ~n18425;
  assign n18427 = po8  & ~n18426;
  assign n18428 = ~n17793 & ~n17797;
  assign n18429 = ~n17801 & n18428;
  assign n18430 = po5  & n18429;
  assign n18431 = po5  & n18428;
  assign n18432 = n17801 & ~n18431;
  assign n18433 = ~n18430 & ~n18432;
  assign n18434 = ~po8  & ~n18416;
  assign n18435 = ~n18425 & n18434;
  assign n18436 = ~n18433 & ~n18435;
  assign n18437 = ~n18427 & ~n18436;
  assign n18438 = po9  & ~n18437;
  assign n18439 = ~n17804 & ~n17806;
  assign n18440 = n17813 & n18439;
  assign n18441 = po5  & n18440;
  assign n18442 = po5  & n18439;
  assign n18443 = ~n17813 & ~n18442;
  assign n18444 = ~n18441 & ~n18443;
  assign n18445 = ~po9  & n18437;
  assign n18446 = ~n18444 & ~n18445;
  assign n18447 = ~n18438 & ~n18446;
  assign n18448 = po10  & ~n18447;
  assign n18449 = ~n17816 & ~n17823;
  assign n18450 = n17822 & n18449;
  assign n18451 = po5  & n18450;
  assign n18452 = po5  & n18449;
  assign n18453 = ~n17822 & ~n18452;
  assign n18454 = ~n18451 & ~n18453;
  assign n18455 = ~po10  & ~n18438;
  assign n18456 = ~n18446 & n18455;
  assign n18457 = ~n18454 & ~n18456;
  assign n18458 = ~n18448 & ~n18457;
  assign n18459 = po11  & ~n18458;
  assign n18460 = ~n17826 & ~n17834;
  assign n18461 = n17832 & n18460;
  assign n18462 = po5  & n18461;
  assign n18463 = po5  & n18460;
  assign n18464 = ~n17832 & ~n18463;
  assign n18465 = ~n18462 & ~n18464;
  assign n18466 = ~po11  & n18458;
  assign n18467 = ~n18465 & ~n18466;
  assign n18468 = ~n18459 & ~n18467;
  assign n18469 = po12  & ~n18468;
  assign n18470 = ~n17837 & ~n17844;
  assign n18471 = n17843 & n18470;
  assign n18472 = po5  & n18471;
  assign n18473 = po5  & n18470;
  assign n18474 = ~n17843 & ~n18473;
  assign n18475 = ~n18472 & ~n18474;
  assign n18476 = ~po12  & ~n18459;
  assign n18477 = ~n18467 & n18476;
  assign n18478 = ~n18475 & ~n18477;
  assign n18479 = ~n18469 & ~n18478;
  assign n18480 = po13  & ~n18479;
  assign n18481 = ~n17847 & ~n17855;
  assign n18482 = n17853 & n18481;
  assign n18483 = po5  & n18482;
  assign n18484 = po5  & n18481;
  assign n18485 = ~n17853 & ~n18484;
  assign n18486 = ~n18483 & ~n18485;
  assign n18487 = ~po13  & n18479;
  assign n18488 = ~n18486 & ~n18487;
  assign n18489 = ~n18480 & ~n18488;
  assign n18490 = po14  & ~n18489;
  assign n18491 = ~n17858 & ~n17865;
  assign n18492 = n17864 & n18491;
  assign n18493 = po5  & n18492;
  assign n18494 = po5  & n18491;
  assign n18495 = ~n17864 & ~n18494;
  assign n18496 = ~n18493 & ~n18495;
  assign n18497 = ~po14  & ~n18480;
  assign n18498 = ~n18488 & n18497;
  assign n18499 = ~n18496 & ~n18498;
  assign n18500 = ~n18490 & ~n18499;
  assign n18501 = po15  & ~n18500;
  assign n18502 = ~n17868 & ~n17876;
  assign n18503 = n17874 & n18502;
  assign n18504 = po5  & n18503;
  assign n18505 = po5  & n18502;
  assign n18506 = ~n17874 & ~n18505;
  assign n18507 = ~n18504 & ~n18506;
  assign n18508 = ~po15  & n18500;
  assign n18509 = ~n18507 & ~n18508;
  assign n18510 = ~n18501 & ~n18509;
  assign n18511 = po16  & ~n18510;
  assign n18512 = ~n17879 & ~n17886;
  assign n18513 = n17885 & n18512;
  assign n18514 = po5  & n18513;
  assign n18515 = po5  & n18512;
  assign n18516 = ~n17885 & ~n18515;
  assign n18517 = ~n18514 & ~n18516;
  assign n18518 = ~po16  & ~n18501;
  assign n18519 = ~n18509 & n18518;
  assign n18520 = ~n18517 & ~n18519;
  assign n18521 = ~n18511 & ~n18520;
  assign n18522 = po17  & ~n18521;
  assign n18523 = ~n17889 & ~n17897;
  assign n18524 = n17895 & n18523;
  assign n18525 = po5  & n18524;
  assign n18526 = po5  & n18523;
  assign n18527 = ~n17895 & ~n18526;
  assign n18528 = ~n18525 & ~n18527;
  assign n18529 = ~po17  & n18521;
  assign n18530 = ~n18528 & ~n18529;
  assign n18531 = ~n18522 & ~n18530;
  assign n18532 = po18  & ~n18531;
  assign n18533 = ~n17900 & ~n17907;
  assign n18534 = n17906 & n18533;
  assign n18535 = po5  & n18534;
  assign n18536 = po5  & n18533;
  assign n18537 = ~n17906 & ~n18536;
  assign n18538 = ~n18535 & ~n18537;
  assign n18539 = ~po18  & ~n18522;
  assign n18540 = ~n18530 & n18539;
  assign n18541 = ~n18538 & ~n18540;
  assign n18542 = ~n18532 & ~n18541;
  assign n18543 = po19  & ~n18542;
  assign n18544 = ~n17910 & ~n17918;
  assign n18545 = n17916 & n18544;
  assign n18546 = po5  & n18545;
  assign n18547 = po5  & n18544;
  assign n18548 = ~n17916 & ~n18547;
  assign n18549 = ~n18546 & ~n18548;
  assign n18550 = ~po19  & n18542;
  assign n18551 = ~n18549 & ~n18550;
  assign n18552 = ~n18543 & ~n18551;
  assign n18553 = po20  & ~n18552;
  assign n18554 = ~n17921 & ~n17928;
  assign n18555 = n17927 & n18554;
  assign n18556 = po5  & n18555;
  assign n18557 = po5  & n18554;
  assign n18558 = ~n17927 & ~n18557;
  assign n18559 = ~n18556 & ~n18558;
  assign n18560 = ~po20  & ~n18543;
  assign n18561 = ~n18551 & n18560;
  assign n18562 = ~n18559 & ~n18561;
  assign n18563 = ~n18553 & ~n18562;
  assign n18564 = po21  & ~n18563;
  assign n18565 = ~n17931 & ~n17939;
  assign n18566 = n17937 & n18565;
  assign n18567 = po5  & n18566;
  assign n18568 = po5  & n18565;
  assign n18569 = ~n17937 & ~n18568;
  assign n18570 = ~n18567 & ~n18569;
  assign n18571 = ~po21  & n18563;
  assign n18572 = ~n18570 & ~n18571;
  assign n18573 = ~n18564 & ~n18572;
  assign n18574 = po22  & ~n18573;
  assign n18575 = ~n17942 & ~n17949;
  assign n18576 = n17948 & n18575;
  assign n18577 = po5  & n18576;
  assign n18578 = po5  & n18575;
  assign n18579 = ~n17948 & ~n18578;
  assign n18580 = ~n18577 & ~n18579;
  assign n18581 = ~po22  & ~n18564;
  assign n18582 = ~n18572 & n18581;
  assign n18583 = ~n18580 & ~n18582;
  assign n18584 = ~n18574 & ~n18583;
  assign n18585 = po23  & ~n18584;
  assign n18586 = ~n17952 & ~n17960;
  assign n18587 = n17958 & n18586;
  assign n18588 = po5  & n18587;
  assign n18589 = po5  & n18586;
  assign n18590 = ~n17958 & ~n18589;
  assign n18591 = ~n18588 & ~n18590;
  assign n18592 = ~po23  & n18584;
  assign n18593 = ~n18591 & ~n18592;
  assign n18594 = ~n18585 & ~n18593;
  assign n18595 = po24  & ~n18594;
  assign n18596 = ~n17963 & ~n17970;
  assign n18597 = n17969 & n18596;
  assign n18598 = po5  & n18597;
  assign n18599 = po5  & n18596;
  assign n18600 = ~n17969 & ~n18599;
  assign n18601 = ~n18598 & ~n18600;
  assign n18602 = ~po24  & ~n18585;
  assign n18603 = ~n18593 & n18602;
  assign n18604 = ~n18601 & ~n18603;
  assign n18605 = ~n18595 & ~n18604;
  assign n18606 = po25  & ~n18605;
  assign n18607 = ~n17973 & ~n17981;
  assign n18608 = n17979 & n18607;
  assign n18609 = po5  & n18608;
  assign n18610 = po5  & n18607;
  assign n18611 = ~n17979 & ~n18610;
  assign n18612 = ~n18609 & ~n18611;
  assign n18613 = ~po25  & n18605;
  assign n18614 = ~n18612 & ~n18613;
  assign n18615 = ~n18606 & ~n18614;
  assign n18616 = po26  & ~n18615;
  assign n18617 = ~n17984 & ~n17991;
  assign n18618 = n17990 & n18617;
  assign n18619 = po5  & n18618;
  assign n18620 = po5  & n18617;
  assign n18621 = ~n17990 & ~n18620;
  assign n18622 = ~n18619 & ~n18621;
  assign n18623 = ~po26  & ~n18606;
  assign n18624 = ~n18614 & n18623;
  assign n18625 = ~n18622 & ~n18624;
  assign n18626 = ~n18616 & ~n18625;
  assign n18627 = po27  & ~n18626;
  assign n18628 = ~n17994 & ~n18002;
  assign n18629 = n18000 & n18628;
  assign n18630 = po5  & n18629;
  assign n18631 = po5  & n18628;
  assign n18632 = ~n18000 & ~n18631;
  assign n18633 = ~n18630 & ~n18632;
  assign n18634 = ~po27  & n18626;
  assign n18635 = ~n18633 & ~n18634;
  assign n18636 = ~n18627 & ~n18635;
  assign n18637 = po28  & ~n18636;
  assign n18638 = ~n18005 & ~n18012;
  assign n18639 = n18011 & n18638;
  assign n18640 = po5  & n18639;
  assign n18641 = po5  & n18638;
  assign n18642 = ~n18011 & ~n18641;
  assign n18643 = ~n18640 & ~n18642;
  assign n18644 = ~po28  & ~n18627;
  assign n18645 = ~n18635 & n18644;
  assign n18646 = ~n18643 & ~n18645;
  assign n18647 = ~n18637 & ~n18646;
  assign n18648 = po29  & ~n18647;
  assign n18649 = ~n18015 & ~n18023;
  assign n18650 = n18021 & n18649;
  assign n18651 = po5  & n18650;
  assign n18652 = po5  & n18649;
  assign n18653 = ~n18021 & ~n18652;
  assign n18654 = ~n18651 & ~n18653;
  assign n18655 = ~po29  & n18647;
  assign n18656 = ~n18654 & ~n18655;
  assign n18657 = ~n18648 & ~n18656;
  assign n18658 = po30  & ~n18657;
  assign n18659 = ~n18026 & ~n18033;
  assign n18660 = n18032 & n18659;
  assign n18661 = po5  & n18660;
  assign n18662 = po5  & n18659;
  assign n18663 = ~n18032 & ~n18662;
  assign n18664 = ~n18661 & ~n18663;
  assign n18665 = ~po30  & ~n18648;
  assign n18666 = ~n18656 & n18665;
  assign n18667 = ~n18664 & ~n18666;
  assign n18668 = ~n18658 & ~n18667;
  assign n18669 = po31  & ~n18668;
  assign n18670 = ~n18036 & ~n18044;
  assign n18671 = n18042 & n18670;
  assign n18672 = po5  & n18671;
  assign n18673 = po5  & n18670;
  assign n18674 = ~n18042 & ~n18673;
  assign n18675 = ~n18672 & ~n18674;
  assign n18676 = ~po31  & n18668;
  assign n18677 = ~n18675 & ~n18676;
  assign n18678 = ~n18669 & ~n18677;
  assign n18679 = po32  & ~n18678;
  assign n18680 = ~n18047 & ~n18054;
  assign n18681 = n18053 & n18680;
  assign n18682 = po5  & n18681;
  assign n18683 = po5  & n18680;
  assign n18684 = ~n18053 & ~n18683;
  assign n18685 = ~n18682 & ~n18684;
  assign n18686 = ~po32  & ~n18669;
  assign n18687 = ~n18677 & n18686;
  assign n18688 = ~n18685 & ~n18687;
  assign n18689 = ~n18679 & ~n18688;
  assign n18690 = po33  & ~n18689;
  assign n18691 = ~n18057 & ~n18065;
  assign n18692 = n18063 & n18691;
  assign n18693 = po5  & n18692;
  assign n18694 = po5  & n18691;
  assign n18695 = ~n18063 & ~n18694;
  assign n18696 = ~n18693 & ~n18695;
  assign n18697 = ~po33  & n18689;
  assign n18698 = ~n18696 & ~n18697;
  assign n18699 = ~n18690 & ~n18698;
  assign n18700 = po34  & ~n18699;
  assign n18701 = ~n18068 & ~n18075;
  assign n18702 = n18074 & n18701;
  assign n18703 = po5  & n18702;
  assign n18704 = po5  & n18701;
  assign n18705 = ~n18074 & ~n18704;
  assign n18706 = ~n18703 & ~n18705;
  assign n18707 = ~po34  & ~n18690;
  assign n18708 = ~n18698 & n18707;
  assign n18709 = ~n18706 & ~n18708;
  assign n18710 = ~n18700 & ~n18709;
  assign n18711 = po35  & ~n18710;
  assign n18712 = ~n18078 & ~n18086;
  assign n18713 = n18084 & n18712;
  assign n18714 = po5  & n18713;
  assign n18715 = po5  & n18712;
  assign n18716 = ~n18084 & ~n18715;
  assign n18717 = ~n18714 & ~n18716;
  assign n18718 = ~po35  & n18710;
  assign n18719 = ~n18717 & ~n18718;
  assign n18720 = ~n18711 & ~n18719;
  assign n18721 = po36  & ~n18720;
  assign n18722 = ~n18089 & ~n18096;
  assign n18723 = n18095 & n18722;
  assign n18724 = po5  & n18723;
  assign n18725 = po5  & n18722;
  assign n18726 = ~n18095 & ~n18725;
  assign n18727 = ~n18724 & ~n18726;
  assign n18728 = ~po36  & ~n18711;
  assign n18729 = ~n18719 & n18728;
  assign n18730 = ~n18727 & ~n18729;
  assign n18731 = ~n18721 & ~n18730;
  assign n18732 = po37  & ~n18731;
  assign n18733 = ~n18099 & ~n18107;
  assign n18734 = n18105 & n18733;
  assign n18735 = po5  & n18734;
  assign n18736 = po5  & n18733;
  assign n18737 = ~n18105 & ~n18736;
  assign n18738 = ~n18735 & ~n18737;
  assign n18739 = ~po37  & n18731;
  assign n18740 = ~n18738 & ~n18739;
  assign n18741 = ~n18732 & ~n18740;
  assign n18742 = po38  & ~n18741;
  assign n18743 = ~n18110 & ~n18117;
  assign n18744 = n18116 & n18743;
  assign n18745 = po5  & n18744;
  assign n18746 = po5  & n18743;
  assign n18747 = ~n18116 & ~n18746;
  assign n18748 = ~n18745 & ~n18747;
  assign n18749 = ~po38  & ~n18732;
  assign n18750 = ~n18740 & n18749;
  assign n18751 = ~n18748 & ~n18750;
  assign n18752 = ~n18742 & ~n18751;
  assign n18753 = po39  & ~n18752;
  assign n18754 = ~n18120 & ~n18128;
  assign n18755 = n18126 & n18754;
  assign n18756 = po5  & n18755;
  assign n18757 = po5  & n18754;
  assign n18758 = ~n18126 & ~n18757;
  assign n18759 = ~n18756 & ~n18758;
  assign n18760 = ~po39  & n18752;
  assign n18761 = ~n18759 & ~n18760;
  assign n18762 = ~n18753 & ~n18761;
  assign n18763 = po40  & ~n18762;
  assign n18764 = ~n18131 & ~n18138;
  assign n18765 = n18137 & n18764;
  assign n18766 = po5  & n18765;
  assign n18767 = po5  & n18764;
  assign n18768 = ~n18137 & ~n18767;
  assign n18769 = ~n18766 & ~n18768;
  assign n18770 = ~po40  & ~n18753;
  assign n18771 = ~n18761 & n18770;
  assign n18772 = ~n18769 & ~n18771;
  assign n18773 = ~n18763 & ~n18772;
  assign n18774 = po41  & ~n18773;
  assign n18775 = ~n18141 & ~n18149;
  assign n18776 = n18147 & n18775;
  assign n18777 = po5  & n18776;
  assign n18778 = po5  & n18775;
  assign n18779 = ~n18147 & ~n18778;
  assign n18780 = ~n18777 & ~n18779;
  assign n18781 = ~po41  & n18773;
  assign n18782 = ~n18780 & ~n18781;
  assign n18783 = ~n18774 & ~n18782;
  assign n18784 = po42  & ~n18783;
  assign n18785 = ~n18152 & ~n18159;
  assign n18786 = n18158 & n18785;
  assign n18787 = po5  & n18786;
  assign n18788 = po5  & n18785;
  assign n18789 = ~n18158 & ~n18788;
  assign n18790 = ~n18787 & ~n18789;
  assign n18791 = ~po42  & ~n18774;
  assign n18792 = ~n18782 & n18791;
  assign n18793 = ~n18790 & ~n18792;
  assign n18794 = ~n18784 & ~n18793;
  assign n18795 = po43  & ~n18794;
  assign n18796 = ~n18162 & ~n18170;
  assign n18797 = n18168 & n18796;
  assign n18798 = po5  & n18797;
  assign n18799 = po5  & n18796;
  assign n18800 = ~n18168 & ~n18799;
  assign n18801 = ~n18798 & ~n18800;
  assign n18802 = ~po43  & n18794;
  assign n18803 = ~n18801 & ~n18802;
  assign n18804 = ~n18795 & ~n18803;
  assign n18805 = po44  & ~n18804;
  assign n18806 = ~n18173 & ~n18180;
  assign n18807 = n18179 & n18806;
  assign n18808 = po5  & n18807;
  assign n18809 = po5  & n18806;
  assign n18810 = ~n18179 & ~n18809;
  assign n18811 = ~n18808 & ~n18810;
  assign n18812 = ~po44  & ~n18795;
  assign n18813 = ~n18803 & n18812;
  assign n18814 = ~n18811 & ~n18813;
  assign n18815 = ~n18805 & ~n18814;
  assign n18816 = po45  & ~n18815;
  assign n18817 = ~n18183 & ~n18191;
  assign n18818 = n18189 & n18817;
  assign n18819 = po5  & n18818;
  assign n18820 = po5  & n18817;
  assign n18821 = ~n18189 & ~n18820;
  assign n18822 = ~n18819 & ~n18821;
  assign n18823 = ~po45  & n18815;
  assign n18824 = ~n18822 & ~n18823;
  assign n18825 = ~n18816 & ~n18824;
  assign n18826 = po46  & ~n18825;
  assign n18827 = ~n18194 & ~n18201;
  assign n18828 = n18200 & n18827;
  assign n18829 = po5  & n18828;
  assign n18830 = po5  & n18827;
  assign n18831 = ~n18200 & ~n18830;
  assign n18832 = ~n18829 & ~n18831;
  assign n18833 = ~po46  & ~n18816;
  assign n18834 = ~n18824 & n18833;
  assign n18835 = ~n18832 & ~n18834;
  assign n18836 = ~n18826 & ~n18835;
  assign n18837 = po47  & ~n18836;
  assign n18838 = ~n18204 & ~n18212;
  assign n18839 = n18210 & n18838;
  assign n18840 = po5  & n18839;
  assign n18841 = po5  & n18838;
  assign n18842 = ~n18210 & ~n18841;
  assign n18843 = ~n18840 & ~n18842;
  assign n18844 = ~po47  & n18836;
  assign n18845 = ~n18843 & ~n18844;
  assign n18846 = ~n18837 & ~n18845;
  assign n18847 = po48  & ~n18846;
  assign n18848 = ~n18215 & ~n18222;
  assign n18849 = n18221 & n18848;
  assign n18850 = po5  & n18849;
  assign n18851 = po5  & n18848;
  assign n18852 = ~n18221 & ~n18851;
  assign n18853 = ~n18850 & ~n18852;
  assign n18854 = ~po48  & ~n18837;
  assign n18855 = ~n18845 & n18854;
  assign n18856 = ~n18853 & ~n18855;
  assign n18857 = ~n18847 & ~n18856;
  assign n18858 = po49  & ~n18857;
  assign n18859 = ~n18225 & ~n18233;
  assign n18860 = n18231 & n18859;
  assign n18861 = po5  & n18860;
  assign n18862 = po5  & n18859;
  assign n18863 = ~n18231 & ~n18862;
  assign n18864 = ~n18861 & ~n18863;
  assign n18865 = ~po49  & n18857;
  assign n18866 = ~n18864 & ~n18865;
  assign n18867 = ~n18858 & ~n18866;
  assign n18868 = po50  & ~n18867;
  assign n18869 = ~n18236 & ~n18243;
  assign n18870 = n18242 & n18869;
  assign n18871 = po5  & n18870;
  assign n18872 = po5  & n18869;
  assign n18873 = ~n18242 & ~n18872;
  assign n18874 = ~n18871 & ~n18873;
  assign n18875 = ~po50  & ~n18858;
  assign n18876 = ~n18866 & n18875;
  assign n18877 = ~n18874 & ~n18876;
  assign n18878 = ~n18868 & ~n18877;
  assign n18879 = po51  & ~n18878;
  assign n18880 = ~n18246 & ~n18254;
  assign n18881 = n18252 & n18880;
  assign n18882 = po5  & n18881;
  assign n18883 = po5  & n18880;
  assign n18884 = ~n18252 & ~n18883;
  assign n18885 = ~n18882 & ~n18884;
  assign n18886 = ~po51  & n18878;
  assign n18887 = ~n18885 & ~n18886;
  assign n18888 = ~n18879 & ~n18887;
  assign n18889 = po52  & ~n18888;
  assign n18890 = ~n18257 & ~n18264;
  assign n18891 = n18263 & n18890;
  assign n18892 = po5  & n18891;
  assign n18893 = po5  & n18890;
  assign n18894 = ~n18263 & ~n18893;
  assign n18895 = ~n18892 & ~n18894;
  assign n18896 = ~po52  & ~n18879;
  assign n18897 = ~n18887 & n18896;
  assign n18898 = ~n18895 & ~n18897;
  assign n18899 = ~n18889 & ~n18898;
  assign n18900 = po53  & ~n18899;
  assign n18901 = ~n18267 & ~n18275;
  assign n18902 = n18273 & n18901;
  assign n18903 = po5  & n18902;
  assign n18904 = po5  & n18901;
  assign n18905 = ~n18273 & ~n18904;
  assign n18906 = ~n18903 & ~n18905;
  assign n18907 = ~po53  & n18899;
  assign n18908 = ~n18906 & ~n18907;
  assign n18909 = ~n18900 & ~n18908;
  assign n18910 = po54  & ~n18909;
  assign n18911 = ~n18278 & ~n18285;
  assign n18912 = n18284 & n18911;
  assign n18913 = po5  & n18912;
  assign n18914 = po5  & n18911;
  assign n18915 = ~n18284 & ~n18914;
  assign n18916 = ~n18913 & ~n18915;
  assign n18917 = ~po54  & ~n18900;
  assign n18918 = ~n18908 & n18917;
  assign n18919 = ~n18916 & ~n18918;
  assign n18920 = ~n18910 & ~n18919;
  assign n18921 = po55  & ~n18920;
  assign n18922 = ~n18288 & ~n18296;
  assign n18923 = n18294 & n18922;
  assign n18924 = po5  & n18923;
  assign n18925 = po5  & n18922;
  assign n18926 = ~n18294 & ~n18925;
  assign n18927 = ~n18924 & ~n18926;
  assign n18928 = ~po55  & n18920;
  assign n18929 = ~n18927 & ~n18928;
  assign n18930 = ~n18921 & ~n18929;
  assign n18931 = po56  & ~n18930;
  assign n18932 = ~n18299 & ~n18306;
  assign n18933 = n18305 & n18932;
  assign n18934 = po5  & n18933;
  assign n18935 = po5  & n18932;
  assign n18936 = ~n18305 & ~n18935;
  assign n18937 = ~n18934 & ~n18936;
  assign n18938 = ~po56  & ~n18921;
  assign n18939 = ~n18929 & n18938;
  assign n18940 = ~n18937 & ~n18939;
  assign n18941 = ~n18931 & ~n18940;
  assign n18942 = po57  & ~n18941;
  assign n18943 = ~n18309 & ~n18317;
  assign n18944 = n18315 & n18943;
  assign n18945 = po5  & n18944;
  assign n18946 = po5  & n18943;
  assign n18947 = ~n18315 & ~n18946;
  assign n18948 = ~n18945 & ~n18947;
  assign n18949 = ~po57  & n18941;
  assign n18950 = ~n18948 & ~n18949;
  assign n18951 = ~n18942 & ~n18950;
  assign n18952 = po58  & ~n18951;
  assign n18953 = ~n18320 & ~n18327;
  assign n18954 = n18326 & n18953;
  assign n18955 = po5  & n18954;
  assign n18956 = po5  & n18953;
  assign n18957 = ~n18326 & ~n18956;
  assign n18958 = ~n18955 & ~n18957;
  assign n18959 = ~po58  & ~n18942;
  assign n18960 = ~n18950 & n18959;
  assign n18961 = ~n18958 & ~n18960;
  assign n18962 = ~n18952 & ~n18961;
  assign n18963 = po59  & ~n18962;
  assign n18964 = ~n18330 & ~n18338;
  assign n18965 = n18336 & n18964;
  assign n18966 = po5  & n18965;
  assign n18967 = po5  & n18964;
  assign n18968 = ~n18336 & ~n18967;
  assign n18969 = ~n18966 & ~n18968;
  assign n18970 = ~po59  & n18962;
  assign n18971 = ~n18969 & ~n18970;
  assign n18972 = ~n18963 & ~n18971;
  assign n18973 = po60  & ~n18972;
  assign n18974 = ~po60  & ~n18963;
  assign n18975 = ~n18971 & n18974;
  assign n18976 = ~n18341 & ~n18348;
  assign n18977 = n18347 & n18976;
  assign n18978 = po5  & n18977;
  assign n18979 = po5  & n18976;
  assign n18980 = ~n18347 & ~n18979;
  assign n18981 = ~n18978 & ~n18980;
  assign n18982 = ~n18975 & ~n18981;
  assign n18983 = ~n18973 & ~n18982;
  assign n18984 = po61  & ~n18983;
  assign n18985 = ~n18351 & ~n18359;
  assign n18986 = n18357 & n18985;
  assign n18987 = po5  & n18986;
  assign n18988 = po5  & n18985;
  assign n18989 = ~n18357 & ~n18988;
  assign n18990 = ~n18987 & ~n18989;
  assign n18991 = ~po61  & n18983;
  assign n18992 = ~n18990 & ~n18991;
  assign n18993 = ~n18984 & ~n18992;
  assign n18994 = po62  & ~n18993;
  assign n18995 = ~n18362 & ~n18369;
  assign n18996 = n18368 & n18995;
  assign n18997 = po5  & n18996;
  assign n18998 = po5  & n18995;
  assign n18999 = ~n18368 & ~n18998;
  assign n19000 = ~n18997 & ~n18999;
  assign n19001 = ~po62  & ~n18984;
  assign n19002 = ~n18992 & n19001;
  assign n19003 = ~n19000 & ~n19002;
  assign n19004 = ~n18994 & ~n19003;
  assign n19005 = ~n18372 & ~n18380;
  assign n19006 = po5  & n19005;
  assign n19007 = ~n18378 & ~n19006;
  assign n19008 = n18378 & n19006;
  assign n19009 = ~n19007 & ~n19008;
  assign n19010 = ~n18382 & ~n18387;
  assign n19011 = po5  & n19010;
  assign n19012 = ~n18398 & ~n19011;
  assign n19013 = ~n19009 & n19012;
  assign n19014 = ~n19004 & n19013;
  assign n19015 = ~po63  & ~n19014;
  assign n19016 = ~n18387 & po5 ;
  assign n19017 = n18382 & ~n19016;
  assign n19018 = po63  & ~n19010;
  assign n19019 = ~n19017 & n19018;
  assign n19020 = n19004 & n19009;
  assign n19021 = ~n19019 & ~n19020;
  assign po4  = n19015 | ~n19021;
  assign n19023 = pi8  & po4 ;
  assign n19024 = ~pi6  & ~pi7 ;
  assign n19025 = ~pi8  & n19024;
  assign n19026 = ~n19023 & ~n19025;
  assign n19027 = po5  & ~n19026;
  assign n19028 = ~n18397 & ~n19025;
  assign n19029 = ~n18398 & n19028;
  assign n19030 = ~n18393 & n19029;
  assign n19031 = ~n19023 & n19030;
  assign n19032 = ~pi8  & po4 ;
  assign n19033 = pi9  & ~n19032;
  assign n19034 = n18402 & po4 ;
  assign n19035 = ~n19033 & ~n19034;
  assign n19036 = ~n19031 & n19035;
  assign n19037 = ~n19027 & ~n19036;
  assign n19038 = po6  & ~n19037;
  assign n19039 = ~po6  & ~n19027;
  assign n19040 = ~n19036 & n19039;
  assign n19041 = po5  & ~n19019;
  assign n19042 = ~n19020 & n19041;
  assign n19043 = ~n19015 & n19042;
  assign n19044 = ~n19034 & ~n19043;
  assign n19045 = pi10  & ~n19044;
  assign n19046 = ~pi10  & n19044;
  assign n19047 = ~n19045 & ~n19046;
  assign n19048 = ~n19040 & ~n19047;
  assign n19049 = ~n19038 & ~n19048;
  assign n19050 = po7  & ~n19049;
  assign n19051 = ~n18405 & ~n18409;
  assign n19052 = ~n18413 & n19051;
  assign n19053 = po4  & n19052;
  assign n19054 = po4  & n19051;
  assign n19055 = n18413 & ~n19054;
  assign n19056 = ~n19053 & ~n19055;
  assign n19057 = ~po7  & n19049;
  assign n19058 = ~n19056 & ~n19057;
  assign n19059 = ~n19050 & ~n19058;
  assign n19060 = po8  & ~n19059;
  assign n19061 = ~n18416 & ~n18424;
  assign n19062 = ~n18425 & n19061;
  assign n19063 = po4  & n19062;
  assign n19064 = po4  & n19061;
  assign n19065 = ~n18423 & ~n19064;
  assign n19066 = ~n19063 & ~n19065;
  assign n19067 = ~po8  & ~n19050;
  assign n19068 = ~n19058 & n19067;
  assign n19069 = ~n19066 & ~n19068;
  assign n19070 = ~n19060 & ~n19069;
  assign n19071 = po9  & ~n19070;
  assign n19072 = ~n18427 & ~n18435;
  assign n19073 = n18433 & n19072;
  assign n19074 = po4  & n19073;
  assign n19075 = po4  & n19072;
  assign n19076 = ~n18433 & ~n19075;
  assign n19077 = ~n19074 & ~n19076;
  assign n19078 = ~po9  & n19070;
  assign n19079 = ~n19077 & ~n19078;
  assign n19080 = ~n19071 & ~n19079;
  assign n19081 = po10  & ~n19080;
  assign n19082 = ~n18438 & ~n18445;
  assign n19083 = n18444 & n19082;
  assign n19084 = po4  & n19083;
  assign n19085 = po4  & n19082;
  assign n19086 = ~n18444 & ~n19085;
  assign n19087 = ~n19084 & ~n19086;
  assign n19088 = ~po10  & ~n19071;
  assign n19089 = ~n19079 & n19088;
  assign n19090 = ~n19087 & ~n19089;
  assign n19091 = ~n19081 & ~n19090;
  assign n19092 = po11  & ~n19091;
  assign n19093 = ~n18448 & ~n18456;
  assign n19094 = n18454 & n19093;
  assign n19095 = po4  & n19094;
  assign n19096 = po4  & n19093;
  assign n19097 = ~n18454 & ~n19096;
  assign n19098 = ~n19095 & ~n19097;
  assign n19099 = ~po11  & n19091;
  assign n19100 = ~n19098 & ~n19099;
  assign n19101 = ~n19092 & ~n19100;
  assign n19102 = po12  & ~n19101;
  assign n19103 = ~n18459 & ~n18466;
  assign n19104 = n18465 & n19103;
  assign n19105 = po4  & n19104;
  assign n19106 = po4  & n19103;
  assign n19107 = ~n18465 & ~n19106;
  assign n19108 = ~n19105 & ~n19107;
  assign n19109 = ~po12  & ~n19092;
  assign n19110 = ~n19100 & n19109;
  assign n19111 = ~n19108 & ~n19110;
  assign n19112 = ~n19102 & ~n19111;
  assign n19113 = po13  & ~n19112;
  assign n19114 = ~n18469 & ~n18477;
  assign n19115 = n18475 & n19114;
  assign n19116 = po4  & n19115;
  assign n19117 = po4  & n19114;
  assign n19118 = ~n18475 & ~n19117;
  assign n19119 = ~n19116 & ~n19118;
  assign n19120 = ~po13  & n19112;
  assign n19121 = ~n19119 & ~n19120;
  assign n19122 = ~n19113 & ~n19121;
  assign n19123 = po14  & ~n19122;
  assign n19124 = ~n18480 & ~n18487;
  assign n19125 = n18486 & n19124;
  assign n19126 = po4  & n19125;
  assign n19127 = po4  & n19124;
  assign n19128 = ~n18486 & ~n19127;
  assign n19129 = ~n19126 & ~n19128;
  assign n19130 = ~po14  & ~n19113;
  assign n19131 = ~n19121 & n19130;
  assign n19132 = ~n19129 & ~n19131;
  assign n19133 = ~n19123 & ~n19132;
  assign n19134 = po15  & ~n19133;
  assign n19135 = ~n18490 & ~n18498;
  assign n19136 = n18496 & n19135;
  assign n19137 = po4  & n19136;
  assign n19138 = po4  & n19135;
  assign n19139 = ~n18496 & ~n19138;
  assign n19140 = ~n19137 & ~n19139;
  assign n19141 = ~po15  & n19133;
  assign n19142 = ~n19140 & ~n19141;
  assign n19143 = ~n19134 & ~n19142;
  assign n19144 = po16  & ~n19143;
  assign n19145 = ~n18501 & ~n18508;
  assign n19146 = n18507 & n19145;
  assign n19147 = po4  & n19146;
  assign n19148 = po4  & n19145;
  assign n19149 = ~n18507 & ~n19148;
  assign n19150 = ~n19147 & ~n19149;
  assign n19151 = ~po16  & ~n19134;
  assign n19152 = ~n19142 & n19151;
  assign n19153 = ~n19150 & ~n19152;
  assign n19154 = ~n19144 & ~n19153;
  assign n19155 = po17  & ~n19154;
  assign n19156 = ~n18511 & ~n18519;
  assign n19157 = n18517 & n19156;
  assign n19158 = po4  & n19157;
  assign n19159 = po4  & n19156;
  assign n19160 = ~n18517 & ~n19159;
  assign n19161 = ~n19158 & ~n19160;
  assign n19162 = ~po17  & n19154;
  assign n19163 = ~n19161 & ~n19162;
  assign n19164 = ~n19155 & ~n19163;
  assign n19165 = po18  & ~n19164;
  assign n19166 = ~n18522 & ~n18529;
  assign n19167 = n18528 & n19166;
  assign n19168 = po4  & n19167;
  assign n19169 = po4  & n19166;
  assign n19170 = ~n18528 & ~n19169;
  assign n19171 = ~n19168 & ~n19170;
  assign n19172 = ~po18  & ~n19155;
  assign n19173 = ~n19163 & n19172;
  assign n19174 = ~n19171 & ~n19173;
  assign n19175 = ~n19165 & ~n19174;
  assign n19176 = po19  & ~n19175;
  assign n19177 = ~n18532 & ~n18540;
  assign n19178 = n18538 & n19177;
  assign n19179 = po4  & n19178;
  assign n19180 = po4  & n19177;
  assign n19181 = ~n18538 & ~n19180;
  assign n19182 = ~n19179 & ~n19181;
  assign n19183 = ~po19  & n19175;
  assign n19184 = ~n19182 & ~n19183;
  assign n19185 = ~n19176 & ~n19184;
  assign n19186 = po20  & ~n19185;
  assign n19187 = ~n18543 & ~n18550;
  assign n19188 = n18549 & n19187;
  assign n19189 = po4  & n19188;
  assign n19190 = po4  & n19187;
  assign n19191 = ~n18549 & ~n19190;
  assign n19192 = ~n19189 & ~n19191;
  assign n19193 = ~po20  & ~n19176;
  assign n19194 = ~n19184 & n19193;
  assign n19195 = ~n19192 & ~n19194;
  assign n19196 = ~n19186 & ~n19195;
  assign n19197 = po21  & ~n19196;
  assign n19198 = ~n18553 & ~n18561;
  assign n19199 = n18559 & n19198;
  assign n19200 = po4  & n19199;
  assign n19201 = po4  & n19198;
  assign n19202 = ~n18559 & ~n19201;
  assign n19203 = ~n19200 & ~n19202;
  assign n19204 = ~po21  & n19196;
  assign n19205 = ~n19203 & ~n19204;
  assign n19206 = ~n19197 & ~n19205;
  assign n19207 = po22  & ~n19206;
  assign n19208 = ~n18564 & ~n18571;
  assign n19209 = n18570 & n19208;
  assign n19210 = po4  & n19209;
  assign n19211 = po4  & n19208;
  assign n19212 = ~n18570 & ~n19211;
  assign n19213 = ~n19210 & ~n19212;
  assign n19214 = ~po22  & ~n19197;
  assign n19215 = ~n19205 & n19214;
  assign n19216 = ~n19213 & ~n19215;
  assign n19217 = ~n19207 & ~n19216;
  assign n19218 = po23  & ~n19217;
  assign n19219 = ~n18574 & ~n18582;
  assign n19220 = n18580 & n19219;
  assign n19221 = po4  & n19220;
  assign n19222 = po4  & n19219;
  assign n19223 = ~n18580 & ~n19222;
  assign n19224 = ~n19221 & ~n19223;
  assign n19225 = ~po23  & n19217;
  assign n19226 = ~n19224 & ~n19225;
  assign n19227 = ~n19218 & ~n19226;
  assign n19228 = po24  & ~n19227;
  assign n19229 = ~n18585 & ~n18592;
  assign n19230 = n18591 & n19229;
  assign n19231 = po4  & n19230;
  assign n19232 = po4  & n19229;
  assign n19233 = ~n18591 & ~n19232;
  assign n19234 = ~n19231 & ~n19233;
  assign n19235 = ~po24  & ~n19218;
  assign n19236 = ~n19226 & n19235;
  assign n19237 = ~n19234 & ~n19236;
  assign n19238 = ~n19228 & ~n19237;
  assign n19239 = po25  & ~n19238;
  assign n19240 = ~n18595 & ~n18603;
  assign n19241 = n18601 & n19240;
  assign n19242 = po4  & n19241;
  assign n19243 = po4  & n19240;
  assign n19244 = ~n18601 & ~n19243;
  assign n19245 = ~n19242 & ~n19244;
  assign n19246 = ~po25  & n19238;
  assign n19247 = ~n19245 & ~n19246;
  assign n19248 = ~n19239 & ~n19247;
  assign n19249 = po26  & ~n19248;
  assign n19250 = ~n18606 & ~n18613;
  assign n19251 = n18612 & n19250;
  assign n19252 = po4  & n19251;
  assign n19253 = po4  & n19250;
  assign n19254 = ~n18612 & ~n19253;
  assign n19255 = ~n19252 & ~n19254;
  assign n19256 = ~po26  & ~n19239;
  assign n19257 = ~n19247 & n19256;
  assign n19258 = ~n19255 & ~n19257;
  assign n19259 = ~n19249 & ~n19258;
  assign n19260 = po27  & ~n19259;
  assign n19261 = ~n18616 & ~n18624;
  assign n19262 = n18622 & n19261;
  assign n19263 = po4  & n19262;
  assign n19264 = po4  & n19261;
  assign n19265 = ~n18622 & ~n19264;
  assign n19266 = ~n19263 & ~n19265;
  assign n19267 = ~po27  & n19259;
  assign n19268 = ~n19266 & ~n19267;
  assign n19269 = ~n19260 & ~n19268;
  assign n19270 = po28  & ~n19269;
  assign n19271 = ~n18627 & ~n18634;
  assign n19272 = n18633 & n19271;
  assign n19273 = po4  & n19272;
  assign n19274 = po4  & n19271;
  assign n19275 = ~n18633 & ~n19274;
  assign n19276 = ~n19273 & ~n19275;
  assign n19277 = ~po28  & ~n19260;
  assign n19278 = ~n19268 & n19277;
  assign n19279 = ~n19276 & ~n19278;
  assign n19280 = ~n19270 & ~n19279;
  assign n19281 = po29  & ~n19280;
  assign n19282 = ~n18637 & ~n18645;
  assign n19283 = n18643 & n19282;
  assign n19284 = po4  & n19283;
  assign n19285 = po4  & n19282;
  assign n19286 = ~n18643 & ~n19285;
  assign n19287 = ~n19284 & ~n19286;
  assign n19288 = ~po29  & n19280;
  assign n19289 = ~n19287 & ~n19288;
  assign n19290 = ~n19281 & ~n19289;
  assign n19291 = po30  & ~n19290;
  assign n19292 = ~n18648 & ~n18655;
  assign n19293 = n18654 & n19292;
  assign n19294 = po4  & n19293;
  assign n19295 = po4  & n19292;
  assign n19296 = ~n18654 & ~n19295;
  assign n19297 = ~n19294 & ~n19296;
  assign n19298 = ~po30  & ~n19281;
  assign n19299 = ~n19289 & n19298;
  assign n19300 = ~n19297 & ~n19299;
  assign n19301 = ~n19291 & ~n19300;
  assign n19302 = po31  & ~n19301;
  assign n19303 = ~n18658 & ~n18666;
  assign n19304 = n18664 & n19303;
  assign n19305 = po4  & n19304;
  assign n19306 = po4  & n19303;
  assign n19307 = ~n18664 & ~n19306;
  assign n19308 = ~n19305 & ~n19307;
  assign n19309 = ~po31  & n19301;
  assign n19310 = ~n19308 & ~n19309;
  assign n19311 = ~n19302 & ~n19310;
  assign n19312 = po32  & ~n19311;
  assign n19313 = ~n18669 & ~n18676;
  assign n19314 = n18675 & n19313;
  assign n19315 = po4  & n19314;
  assign n19316 = po4  & n19313;
  assign n19317 = ~n18675 & ~n19316;
  assign n19318 = ~n19315 & ~n19317;
  assign n19319 = ~po32  & ~n19302;
  assign n19320 = ~n19310 & n19319;
  assign n19321 = ~n19318 & ~n19320;
  assign n19322 = ~n19312 & ~n19321;
  assign n19323 = po33  & ~n19322;
  assign n19324 = ~n18679 & ~n18687;
  assign n19325 = n18685 & n19324;
  assign n19326 = po4  & n19325;
  assign n19327 = po4  & n19324;
  assign n19328 = ~n18685 & ~n19327;
  assign n19329 = ~n19326 & ~n19328;
  assign n19330 = ~po33  & n19322;
  assign n19331 = ~n19329 & ~n19330;
  assign n19332 = ~n19323 & ~n19331;
  assign n19333 = po34  & ~n19332;
  assign n19334 = ~n18690 & ~n18697;
  assign n19335 = n18696 & n19334;
  assign n19336 = po4  & n19335;
  assign n19337 = po4  & n19334;
  assign n19338 = ~n18696 & ~n19337;
  assign n19339 = ~n19336 & ~n19338;
  assign n19340 = ~po34  & ~n19323;
  assign n19341 = ~n19331 & n19340;
  assign n19342 = ~n19339 & ~n19341;
  assign n19343 = ~n19333 & ~n19342;
  assign n19344 = po35  & ~n19343;
  assign n19345 = ~n18700 & ~n18708;
  assign n19346 = n18706 & n19345;
  assign n19347 = po4  & n19346;
  assign n19348 = po4  & n19345;
  assign n19349 = ~n18706 & ~n19348;
  assign n19350 = ~n19347 & ~n19349;
  assign n19351 = ~po35  & n19343;
  assign n19352 = ~n19350 & ~n19351;
  assign n19353 = ~n19344 & ~n19352;
  assign n19354 = po36  & ~n19353;
  assign n19355 = ~n18711 & ~n18718;
  assign n19356 = n18717 & n19355;
  assign n19357 = po4  & n19356;
  assign n19358 = po4  & n19355;
  assign n19359 = ~n18717 & ~n19358;
  assign n19360 = ~n19357 & ~n19359;
  assign n19361 = ~po36  & ~n19344;
  assign n19362 = ~n19352 & n19361;
  assign n19363 = ~n19360 & ~n19362;
  assign n19364 = ~n19354 & ~n19363;
  assign n19365 = po37  & ~n19364;
  assign n19366 = ~n18721 & ~n18729;
  assign n19367 = n18727 & n19366;
  assign n19368 = po4  & n19367;
  assign n19369 = po4  & n19366;
  assign n19370 = ~n18727 & ~n19369;
  assign n19371 = ~n19368 & ~n19370;
  assign n19372 = ~po37  & n19364;
  assign n19373 = ~n19371 & ~n19372;
  assign n19374 = ~n19365 & ~n19373;
  assign n19375 = po38  & ~n19374;
  assign n19376 = ~n18732 & ~n18739;
  assign n19377 = n18738 & n19376;
  assign n19378 = po4  & n19377;
  assign n19379 = po4  & n19376;
  assign n19380 = ~n18738 & ~n19379;
  assign n19381 = ~n19378 & ~n19380;
  assign n19382 = ~po38  & ~n19365;
  assign n19383 = ~n19373 & n19382;
  assign n19384 = ~n19381 & ~n19383;
  assign n19385 = ~n19375 & ~n19384;
  assign n19386 = po39  & ~n19385;
  assign n19387 = ~n18742 & ~n18750;
  assign n19388 = n18748 & n19387;
  assign n19389 = po4  & n19388;
  assign n19390 = po4  & n19387;
  assign n19391 = ~n18748 & ~n19390;
  assign n19392 = ~n19389 & ~n19391;
  assign n19393 = ~po39  & n19385;
  assign n19394 = ~n19392 & ~n19393;
  assign n19395 = ~n19386 & ~n19394;
  assign n19396 = po40  & ~n19395;
  assign n19397 = ~n18753 & ~n18760;
  assign n19398 = n18759 & n19397;
  assign n19399 = po4  & n19398;
  assign n19400 = po4  & n19397;
  assign n19401 = ~n18759 & ~n19400;
  assign n19402 = ~n19399 & ~n19401;
  assign n19403 = ~po40  & ~n19386;
  assign n19404 = ~n19394 & n19403;
  assign n19405 = ~n19402 & ~n19404;
  assign n19406 = ~n19396 & ~n19405;
  assign n19407 = po41  & ~n19406;
  assign n19408 = ~n18763 & ~n18771;
  assign n19409 = n18769 & n19408;
  assign n19410 = po4  & n19409;
  assign n19411 = po4  & n19408;
  assign n19412 = ~n18769 & ~n19411;
  assign n19413 = ~n19410 & ~n19412;
  assign n19414 = ~po41  & n19406;
  assign n19415 = ~n19413 & ~n19414;
  assign n19416 = ~n19407 & ~n19415;
  assign n19417 = po42  & ~n19416;
  assign n19418 = ~n18774 & ~n18781;
  assign n19419 = n18780 & n19418;
  assign n19420 = po4  & n19419;
  assign n19421 = po4  & n19418;
  assign n19422 = ~n18780 & ~n19421;
  assign n19423 = ~n19420 & ~n19422;
  assign n19424 = ~po42  & ~n19407;
  assign n19425 = ~n19415 & n19424;
  assign n19426 = ~n19423 & ~n19425;
  assign n19427 = ~n19417 & ~n19426;
  assign n19428 = po43  & ~n19427;
  assign n19429 = ~n18784 & ~n18792;
  assign n19430 = n18790 & n19429;
  assign n19431 = po4  & n19430;
  assign n19432 = po4  & n19429;
  assign n19433 = ~n18790 & ~n19432;
  assign n19434 = ~n19431 & ~n19433;
  assign n19435 = ~po43  & n19427;
  assign n19436 = ~n19434 & ~n19435;
  assign n19437 = ~n19428 & ~n19436;
  assign n19438 = po44  & ~n19437;
  assign n19439 = ~n18795 & ~n18802;
  assign n19440 = n18801 & n19439;
  assign n19441 = po4  & n19440;
  assign n19442 = po4  & n19439;
  assign n19443 = ~n18801 & ~n19442;
  assign n19444 = ~n19441 & ~n19443;
  assign n19445 = ~po44  & ~n19428;
  assign n19446 = ~n19436 & n19445;
  assign n19447 = ~n19444 & ~n19446;
  assign n19448 = ~n19438 & ~n19447;
  assign n19449 = po45  & ~n19448;
  assign n19450 = ~n18805 & ~n18813;
  assign n19451 = n18811 & n19450;
  assign n19452 = po4  & n19451;
  assign n19453 = po4  & n19450;
  assign n19454 = ~n18811 & ~n19453;
  assign n19455 = ~n19452 & ~n19454;
  assign n19456 = ~po45  & n19448;
  assign n19457 = ~n19455 & ~n19456;
  assign n19458 = ~n19449 & ~n19457;
  assign n19459 = po46  & ~n19458;
  assign n19460 = ~n18816 & ~n18823;
  assign n19461 = n18822 & n19460;
  assign n19462 = po4  & n19461;
  assign n19463 = po4  & n19460;
  assign n19464 = ~n18822 & ~n19463;
  assign n19465 = ~n19462 & ~n19464;
  assign n19466 = ~po46  & ~n19449;
  assign n19467 = ~n19457 & n19466;
  assign n19468 = ~n19465 & ~n19467;
  assign n19469 = ~n19459 & ~n19468;
  assign n19470 = po47  & ~n19469;
  assign n19471 = ~n18826 & ~n18834;
  assign n19472 = n18832 & n19471;
  assign n19473 = po4  & n19472;
  assign n19474 = po4  & n19471;
  assign n19475 = ~n18832 & ~n19474;
  assign n19476 = ~n19473 & ~n19475;
  assign n19477 = ~po47  & n19469;
  assign n19478 = ~n19476 & ~n19477;
  assign n19479 = ~n19470 & ~n19478;
  assign n19480 = po48  & ~n19479;
  assign n19481 = ~n18837 & ~n18844;
  assign n19482 = n18843 & n19481;
  assign n19483 = po4  & n19482;
  assign n19484 = po4  & n19481;
  assign n19485 = ~n18843 & ~n19484;
  assign n19486 = ~n19483 & ~n19485;
  assign n19487 = ~po48  & ~n19470;
  assign n19488 = ~n19478 & n19487;
  assign n19489 = ~n19486 & ~n19488;
  assign n19490 = ~n19480 & ~n19489;
  assign n19491 = po49  & ~n19490;
  assign n19492 = ~n18847 & ~n18855;
  assign n19493 = n18853 & n19492;
  assign n19494 = po4  & n19493;
  assign n19495 = po4  & n19492;
  assign n19496 = ~n18853 & ~n19495;
  assign n19497 = ~n19494 & ~n19496;
  assign n19498 = ~po49  & n19490;
  assign n19499 = ~n19497 & ~n19498;
  assign n19500 = ~n19491 & ~n19499;
  assign n19501 = po50  & ~n19500;
  assign n19502 = ~n18858 & ~n18865;
  assign n19503 = n18864 & n19502;
  assign n19504 = po4  & n19503;
  assign n19505 = po4  & n19502;
  assign n19506 = ~n18864 & ~n19505;
  assign n19507 = ~n19504 & ~n19506;
  assign n19508 = ~po50  & ~n19491;
  assign n19509 = ~n19499 & n19508;
  assign n19510 = ~n19507 & ~n19509;
  assign n19511 = ~n19501 & ~n19510;
  assign n19512 = po51  & ~n19511;
  assign n19513 = ~n18868 & ~n18876;
  assign n19514 = n18874 & n19513;
  assign n19515 = po4  & n19514;
  assign n19516 = po4  & n19513;
  assign n19517 = ~n18874 & ~n19516;
  assign n19518 = ~n19515 & ~n19517;
  assign n19519 = ~po51  & n19511;
  assign n19520 = ~n19518 & ~n19519;
  assign n19521 = ~n19512 & ~n19520;
  assign n19522 = po52  & ~n19521;
  assign n19523 = ~n18879 & ~n18886;
  assign n19524 = n18885 & n19523;
  assign n19525 = po4  & n19524;
  assign n19526 = po4  & n19523;
  assign n19527 = ~n18885 & ~n19526;
  assign n19528 = ~n19525 & ~n19527;
  assign n19529 = ~po52  & ~n19512;
  assign n19530 = ~n19520 & n19529;
  assign n19531 = ~n19528 & ~n19530;
  assign n19532 = ~n19522 & ~n19531;
  assign n19533 = po53  & ~n19532;
  assign n19534 = ~n18889 & ~n18897;
  assign n19535 = n18895 & n19534;
  assign n19536 = po4  & n19535;
  assign n19537 = po4  & n19534;
  assign n19538 = ~n18895 & ~n19537;
  assign n19539 = ~n19536 & ~n19538;
  assign n19540 = ~po53  & n19532;
  assign n19541 = ~n19539 & ~n19540;
  assign n19542 = ~n19533 & ~n19541;
  assign n19543 = po54  & ~n19542;
  assign n19544 = ~n18900 & ~n18907;
  assign n19545 = n18906 & n19544;
  assign n19546 = po4  & n19545;
  assign n19547 = po4  & n19544;
  assign n19548 = ~n18906 & ~n19547;
  assign n19549 = ~n19546 & ~n19548;
  assign n19550 = ~po54  & ~n19533;
  assign n19551 = ~n19541 & n19550;
  assign n19552 = ~n19549 & ~n19551;
  assign n19553 = ~n19543 & ~n19552;
  assign n19554 = po55  & ~n19553;
  assign n19555 = ~n18910 & ~n18918;
  assign n19556 = n18916 & n19555;
  assign n19557 = po4  & n19556;
  assign n19558 = po4  & n19555;
  assign n19559 = ~n18916 & ~n19558;
  assign n19560 = ~n19557 & ~n19559;
  assign n19561 = ~po55  & n19553;
  assign n19562 = ~n19560 & ~n19561;
  assign n19563 = ~n19554 & ~n19562;
  assign n19564 = po56  & ~n19563;
  assign n19565 = ~n18921 & ~n18928;
  assign n19566 = n18927 & n19565;
  assign n19567 = po4  & n19566;
  assign n19568 = po4  & n19565;
  assign n19569 = ~n18927 & ~n19568;
  assign n19570 = ~n19567 & ~n19569;
  assign n19571 = ~po56  & ~n19554;
  assign n19572 = ~n19562 & n19571;
  assign n19573 = ~n19570 & ~n19572;
  assign n19574 = ~n19564 & ~n19573;
  assign n19575 = po57  & ~n19574;
  assign n19576 = ~n18931 & ~n18939;
  assign n19577 = n18937 & n19576;
  assign n19578 = po4  & n19577;
  assign n19579 = po4  & n19576;
  assign n19580 = ~n18937 & ~n19579;
  assign n19581 = ~n19578 & ~n19580;
  assign n19582 = ~po57  & n19574;
  assign n19583 = ~n19581 & ~n19582;
  assign n19584 = ~n19575 & ~n19583;
  assign n19585 = po58  & ~n19584;
  assign n19586 = ~n18942 & ~n18949;
  assign n19587 = n18948 & n19586;
  assign n19588 = po4  & n19587;
  assign n19589 = po4  & n19586;
  assign n19590 = ~n18948 & ~n19589;
  assign n19591 = ~n19588 & ~n19590;
  assign n19592 = ~po58  & ~n19575;
  assign n19593 = ~n19583 & n19592;
  assign n19594 = ~n19591 & ~n19593;
  assign n19595 = ~n19585 & ~n19594;
  assign n19596 = po59  & ~n19595;
  assign n19597 = ~n18952 & ~n18960;
  assign n19598 = n18958 & n19597;
  assign n19599 = po4  & n19598;
  assign n19600 = po4  & n19597;
  assign n19601 = ~n18958 & ~n19600;
  assign n19602 = ~n19599 & ~n19601;
  assign n19603 = ~po59  & n19595;
  assign n19604 = ~n19602 & ~n19603;
  assign n19605 = ~n19596 & ~n19604;
  assign n19606 = po60  & ~n19605;
  assign n19607 = ~n18963 & ~n18970;
  assign n19608 = n18969 & n19607;
  assign n19609 = po4  & n19608;
  assign n19610 = po4  & n19607;
  assign n19611 = ~n18969 & ~n19610;
  assign n19612 = ~n19609 & ~n19611;
  assign n19613 = ~po60  & ~n19596;
  assign n19614 = ~n19604 & n19613;
  assign n19615 = ~n19612 & ~n19614;
  assign n19616 = ~n19606 & ~n19615;
  assign n19617 = po61  & ~n19616;
  assign n19618 = ~n18973 & ~n18975;
  assign n19619 = n18981 & n19618;
  assign n19620 = po4  & n19619;
  assign n19621 = po4  & n19618;
  assign n19622 = ~n18981 & ~n19621;
  assign n19623 = ~n19620 & ~n19622;
  assign n19624 = ~po61  & n19616;
  assign n19625 = ~n19623 & ~n19624;
  assign n19626 = ~n19617 & ~n19625;
  assign n19627 = po62  & ~n19626;
  assign n19628 = ~n18984 & ~n18991;
  assign n19629 = n18990 & n19628;
  assign n19630 = po4  & n19629;
  assign n19631 = po4  & n19628;
  assign n19632 = ~n18990 & ~n19631;
  assign n19633 = ~n19630 & ~n19632;
  assign n19634 = ~po62  & ~n19617;
  assign n19635 = ~n19625 & n19634;
  assign n19636 = ~n19633 & ~n19635;
  assign n19637 = ~n19627 & ~n19636;
  assign n19638 = ~n18994 & ~n19002;
  assign n19639 = po4  & n19638;
  assign n19640 = ~n19000 & ~n19639;
  assign n19641 = n19000 & n19639;
  assign n19642 = ~n19640 & ~n19641;
  assign n19643 = ~n19004 & ~n19009;
  assign n19644 = po4  & n19643;
  assign n19645 = ~n19020 & ~n19644;
  assign n19646 = ~n19642 & n19645;
  assign n19647 = ~n19637 & n19646;
  assign n19648 = ~po63  & ~n19647;
  assign n19649 = ~n19009 & po4 ;
  assign n19650 = n19004 & ~n19649;
  assign n19651 = po63  & ~n19643;
  assign n19652 = ~n19650 & n19651;
  assign n19653 = n19637 & n19642;
  assign n19654 = ~n19652 & ~n19653;
  assign po3  = n19648 | ~n19654;
  assign n19656 = pi6  & po3 ;
  assign n19657 = ~pi4  & ~pi5 ;
  assign n19658 = ~pi6  & n19657;
  assign n19659 = ~n19656 & ~n19658;
  assign n19660 = po4  & ~n19659;
  assign n19661 = ~n19019 & ~n19658;
  assign n19662 = ~n19020 & n19661;
  assign n19663 = ~n19015 & n19662;
  assign n19664 = ~n19656 & n19663;
  assign n19665 = ~pi6  & po3 ;
  assign n19666 = pi7  & ~n19665;
  assign n19667 = n19024 & po3 ;
  assign n19668 = ~n19666 & ~n19667;
  assign n19669 = ~n19664 & n19668;
  assign n19670 = ~n19660 & ~n19669;
  assign n19671 = po5  & ~n19670;
  assign n19672 = po4  & ~n19652;
  assign n19673 = ~n19653 & n19672;
  assign n19674 = ~n19648 & n19673;
  assign n19675 = ~n19667 & ~n19674;
  assign n19676 = pi8  & ~n19675;
  assign n19677 = ~pi8  & n19675;
  assign n19678 = ~n19676 & ~n19677;
  assign n19679 = ~po5  & n19670;
  assign n19680 = ~n19678 & ~n19679;
  assign n19681 = ~n19671 & ~n19680;
  assign n19682 = po6  & ~n19681;
  assign n19683 = ~n19027 & ~n19031;
  assign n19684 = ~n19035 & n19683;
  assign n19685 = po3  & n19684;
  assign n19686 = po3  & n19683;
  assign n19687 = n19035 & ~n19686;
  assign n19688 = ~n19685 & ~n19687;
  assign n19689 = ~po6  & ~n19671;
  assign n19690 = ~n19680 & n19689;
  assign n19691 = ~n19688 & ~n19690;
  assign n19692 = ~n19682 & ~n19691;
  assign n19693 = po7  & ~n19692;
  assign n19694 = ~n19038 & ~n19040;
  assign n19695 = ~n19048 & n19694;
  assign n19696 = po3  & n19695;
  assign n19697 = po3  & n19694;
  assign n19698 = ~n19047 & ~n19697;
  assign n19699 = ~n19696 & ~n19698;
  assign n19700 = ~po7  & n19692;
  assign n19701 = ~n19699 & ~n19700;
  assign n19702 = ~n19693 & ~n19701;
  assign n19703 = po8  & ~n19702;
  assign n19704 = ~n19050 & ~n19057;
  assign n19705 = n19056 & n19704;
  assign n19706 = po3  & n19705;
  assign n19707 = po3  & n19704;
  assign n19708 = ~n19056 & ~n19707;
  assign n19709 = ~n19706 & ~n19708;
  assign n19710 = ~po8  & ~n19693;
  assign n19711 = ~n19701 & n19710;
  assign n19712 = ~n19709 & ~n19711;
  assign n19713 = ~n19703 & ~n19712;
  assign n19714 = po9  & ~n19713;
  assign n19715 = ~n19060 & ~n19068;
  assign n19716 = n19066 & n19715;
  assign n19717 = po3  & n19716;
  assign n19718 = po3  & n19715;
  assign n19719 = ~n19066 & ~n19718;
  assign n19720 = ~n19717 & ~n19719;
  assign n19721 = ~po9  & n19713;
  assign n19722 = ~n19720 & ~n19721;
  assign n19723 = ~n19714 & ~n19722;
  assign n19724 = po10  & ~n19723;
  assign n19725 = ~n19071 & ~n19078;
  assign n19726 = n19077 & n19725;
  assign n19727 = po3  & n19726;
  assign n19728 = po3  & n19725;
  assign n19729 = ~n19077 & ~n19728;
  assign n19730 = ~n19727 & ~n19729;
  assign n19731 = ~po10  & ~n19714;
  assign n19732 = ~n19722 & n19731;
  assign n19733 = ~n19730 & ~n19732;
  assign n19734 = ~n19724 & ~n19733;
  assign n19735 = po11  & ~n19734;
  assign n19736 = ~n19081 & ~n19089;
  assign n19737 = n19087 & n19736;
  assign n19738 = po3  & n19737;
  assign n19739 = po3  & n19736;
  assign n19740 = ~n19087 & ~n19739;
  assign n19741 = ~n19738 & ~n19740;
  assign n19742 = ~po11  & n19734;
  assign n19743 = ~n19741 & ~n19742;
  assign n19744 = ~n19735 & ~n19743;
  assign n19745 = po12  & ~n19744;
  assign n19746 = ~n19092 & ~n19099;
  assign n19747 = n19098 & n19746;
  assign n19748 = po3  & n19747;
  assign n19749 = po3  & n19746;
  assign n19750 = ~n19098 & ~n19749;
  assign n19751 = ~n19748 & ~n19750;
  assign n19752 = ~po12  & ~n19735;
  assign n19753 = ~n19743 & n19752;
  assign n19754 = ~n19751 & ~n19753;
  assign n19755 = ~n19745 & ~n19754;
  assign n19756 = po13  & ~n19755;
  assign n19757 = ~n19102 & ~n19110;
  assign n19758 = n19108 & n19757;
  assign n19759 = po3  & n19758;
  assign n19760 = po3  & n19757;
  assign n19761 = ~n19108 & ~n19760;
  assign n19762 = ~n19759 & ~n19761;
  assign n19763 = ~po13  & n19755;
  assign n19764 = ~n19762 & ~n19763;
  assign n19765 = ~n19756 & ~n19764;
  assign n19766 = po14  & ~n19765;
  assign n19767 = ~n19113 & ~n19120;
  assign n19768 = n19119 & n19767;
  assign n19769 = po3  & n19768;
  assign n19770 = po3  & n19767;
  assign n19771 = ~n19119 & ~n19770;
  assign n19772 = ~n19769 & ~n19771;
  assign n19773 = ~po14  & ~n19756;
  assign n19774 = ~n19764 & n19773;
  assign n19775 = ~n19772 & ~n19774;
  assign n19776 = ~n19766 & ~n19775;
  assign n19777 = po15  & ~n19776;
  assign n19778 = ~n19123 & ~n19131;
  assign n19779 = n19129 & n19778;
  assign n19780 = po3  & n19779;
  assign n19781 = po3  & n19778;
  assign n19782 = ~n19129 & ~n19781;
  assign n19783 = ~n19780 & ~n19782;
  assign n19784 = ~po15  & n19776;
  assign n19785 = ~n19783 & ~n19784;
  assign n19786 = ~n19777 & ~n19785;
  assign n19787 = po16  & ~n19786;
  assign n19788 = ~n19134 & ~n19141;
  assign n19789 = n19140 & n19788;
  assign n19790 = po3  & n19789;
  assign n19791 = po3  & n19788;
  assign n19792 = ~n19140 & ~n19791;
  assign n19793 = ~n19790 & ~n19792;
  assign n19794 = ~po16  & ~n19777;
  assign n19795 = ~n19785 & n19794;
  assign n19796 = ~n19793 & ~n19795;
  assign n19797 = ~n19787 & ~n19796;
  assign n19798 = po17  & ~n19797;
  assign n19799 = ~n19144 & ~n19152;
  assign n19800 = n19150 & n19799;
  assign n19801 = po3  & n19800;
  assign n19802 = po3  & n19799;
  assign n19803 = ~n19150 & ~n19802;
  assign n19804 = ~n19801 & ~n19803;
  assign n19805 = ~po17  & n19797;
  assign n19806 = ~n19804 & ~n19805;
  assign n19807 = ~n19798 & ~n19806;
  assign n19808 = po18  & ~n19807;
  assign n19809 = ~n19155 & ~n19162;
  assign n19810 = n19161 & n19809;
  assign n19811 = po3  & n19810;
  assign n19812 = po3  & n19809;
  assign n19813 = ~n19161 & ~n19812;
  assign n19814 = ~n19811 & ~n19813;
  assign n19815 = ~po18  & ~n19798;
  assign n19816 = ~n19806 & n19815;
  assign n19817 = ~n19814 & ~n19816;
  assign n19818 = ~n19808 & ~n19817;
  assign n19819 = po19  & ~n19818;
  assign n19820 = ~n19165 & ~n19173;
  assign n19821 = n19171 & n19820;
  assign n19822 = po3  & n19821;
  assign n19823 = po3  & n19820;
  assign n19824 = ~n19171 & ~n19823;
  assign n19825 = ~n19822 & ~n19824;
  assign n19826 = ~po19  & n19818;
  assign n19827 = ~n19825 & ~n19826;
  assign n19828 = ~n19819 & ~n19827;
  assign n19829 = po20  & ~n19828;
  assign n19830 = ~n19176 & ~n19183;
  assign n19831 = n19182 & n19830;
  assign n19832 = po3  & n19831;
  assign n19833 = po3  & n19830;
  assign n19834 = ~n19182 & ~n19833;
  assign n19835 = ~n19832 & ~n19834;
  assign n19836 = ~po20  & ~n19819;
  assign n19837 = ~n19827 & n19836;
  assign n19838 = ~n19835 & ~n19837;
  assign n19839 = ~n19829 & ~n19838;
  assign n19840 = po21  & ~n19839;
  assign n19841 = ~n19186 & ~n19194;
  assign n19842 = n19192 & n19841;
  assign n19843 = po3  & n19842;
  assign n19844 = po3  & n19841;
  assign n19845 = ~n19192 & ~n19844;
  assign n19846 = ~n19843 & ~n19845;
  assign n19847 = ~po21  & n19839;
  assign n19848 = ~n19846 & ~n19847;
  assign n19849 = ~n19840 & ~n19848;
  assign n19850 = po22  & ~n19849;
  assign n19851 = ~n19197 & ~n19204;
  assign n19852 = n19203 & n19851;
  assign n19853 = po3  & n19852;
  assign n19854 = po3  & n19851;
  assign n19855 = ~n19203 & ~n19854;
  assign n19856 = ~n19853 & ~n19855;
  assign n19857 = ~po22  & ~n19840;
  assign n19858 = ~n19848 & n19857;
  assign n19859 = ~n19856 & ~n19858;
  assign n19860 = ~n19850 & ~n19859;
  assign n19861 = po23  & ~n19860;
  assign n19862 = ~n19207 & ~n19215;
  assign n19863 = n19213 & n19862;
  assign n19864 = po3  & n19863;
  assign n19865 = po3  & n19862;
  assign n19866 = ~n19213 & ~n19865;
  assign n19867 = ~n19864 & ~n19866;
  assign n19868 = ~po23  & n19860;
  assign n19869 = ~n19867 & ~n19868;
  assign n19870 = ~n19861 & ~n19869;
  assign n19871 = po24  & ~n19870;
  assign n19872 = ~n19218 & ~n19225;
  assign n19873 = n19224 & n19872;
  assign n19874 = po3  & n19873;
  assign n19875 = po3  & n19872;
  assign n19876 = ~n19224 & ~n19875;
  assign n19877 = ~n19874 & ~n19876;
  assign n19878 = ~po24  & ~n19861;
  assign n19879 = ~n19869 & n19878;
  assign n19880 = ~n19877 & ~n19879;
  assign n19881 = ~n19871 & ~n19880;
  assign n19882 = po25  & ~n19881;
  assign n19883 = ~n19228 & ~n19236;
  assign n19884 = n19234 & n19883;
  assign n19885 = po3  & n19884;
  assign n19886 = po3  & n19883;
  assign n19887 = ~n19234 & ~n19886;
  assign n19888 = ~n19885 & ~n19887;
  assign n19889 = ~po25  & n19881;
  assign n19890 = ~n19888 & ~n19889;
  assign n19891 = ~n19882 & ~n19890;
  assign n19892 = po26  & ~n19891;
  assign n19893 = ~n19239 & ~n19246;
  assign n19894 = n19245 & n19893;
  assign n19895 = po3  & n19894;
  assign n19896 = po3  & n19893;
  assign n19897 = ~n19245 & ~n19896;
  assign n19898 = ~n19895 & ~n19897;
  assign n19899 = ~po26  & ~n19882;
  assign n19900 = ~n19890 & n19899;
  assign n19901 = ~n19898 & ~n19900;
  assign n19902 = ~n19892 & ~n19901;
  assign n19903 = po27  & ~n19902;
  assign n19904 = ~n19249 & ~n19257;
  assign n19905 = n19255 & n19904;
  assign n19906 = po3  & n19905;
  assign n19907 = po3  & n19904;
  assign n19908 = ~n19255 & ~n19907;
  assign n19909 = ~n19906 & ~n19908;
  assign n19910 = ~po27  & n19902;
  assign n19911 = ~n19909 & ~n19910;
  assign n19912 = ~n19903 & ~n19911;
  assign n19913 = po28  & ~n19912;
  assign n19914 = ~n19260 & ~n19267;
  assign n19915 = n19266 & n19914;
  assign n19916 = po3  & n19915;
  assign n19917 = po3  & n19914;
  assign n19918 = ~n19266 & ~n19917;
  assign n19919 = ~n19916 & ~n19918;
  assign n19920 = ~po28  & ~n19903;
  assign n19921 = ~n19911 & n19920;
  assign n19922 = ~n19919 & ~n19921;
  assign n19923 = ~n19913 & ~n19922;
  assign n19924 = po29  & ~n19923;
  assign n19925 = ~n19270 & ~n19278;
  assign n19926 = n19276 & n19925;
  assign n19927 = po3  & n19926;
  assign n19928 = po3  & n19925;
  assign n19929 = ~n19276 & ~n19928;
  assign n19930 = ~n19927 & ~n19929;
  assign n19931 = ~po29  & n19923;
  assign n19932 = ~n19930 & ~n19931;
  assign n19933 = ~n19924 & ~n19932;
  assign n19934 = po30  & ~n19933;
  assign n19935 = ~n19281 & ~n19288;
  assign n19936 = n19287 & n19935;
  assign n19937 = po3  & n19936;
  assign n19938 = po3  & n19935;
  assign n19939 = ~n19287 & ~n19938;
  assign n19940 = ~n19937 & ~n19939;
  assign n19941 = ~po30  & ~n19924;
  assign n19942 = ~n19932 & n19941;
  assign n19943 = ~n19940 & ~n19942;
  assign n19944 = ~n19934 & ~n19943;
  assign n19945 = po31  & ~n19944;
  assign n19946 = ~n19291 & ~n19299;
  assign n19947 = n19297 & n19946;
  assign n19948 = po3  & n19947;
  assign n19949 = po3  & n19946;
  assign n19950 = ~n19297 & ~n19949;
  assign n19951 = ~n19948 & ~n19950;
  assign n19952 = ~po31  & n19944;
  assign n19953 = ~n19951 & ~n19952;
  assign n19954 = ~n19945 & ~n19953;
  assign n19955 = po32  & ~n19954;
  assign n19956 = ~n19302 & ~n19309;
  assign n19957 = n19308 & n19956;
  assign n19958 = po3  & n19957;
  assign n19959 = po3  & n19956;
  assign n19960 = ~n19308 & ~n19959;
  assign n19961 = ~n19958 & ~n19960;
  assign n19962 = ~po32  & ~n19945;
  assign n19963 = ~n19953 & n19962;
  assign n19964 = ~n19961 & ~n19963;
  assign n19965 = ~n19955 & ~n19964;
  assign n19966 = po33  & ~n19965;
  assign n19967 = ~n19312 & ~n19320;
  assign n19968 = n19318 & n19967;
  assign n19969 = po3  & n19968;
  assign n19970 = po3  & n19967;
  assign n19971 = ~n19318 & ~n19970;
  assign n19972 = ~n19969 & ~n19971;
  assign n19973 = ~po33  & n19965;
  assign n19974 = ~n19972 & ~n19973;
  assign n19975 = ~n19966 & ~n19974;
  assign n19976 = po34  & ~n19975;
  assign n19977 = ~n19323 & ~n19330;
  assign n19978 = n19329 & n19977;
  assign n19979 = po3  & n19978;
  assign n19980 = po3  & n19977;
  assign n19981 = ~n19329 & ~n19980;
  assign n19982 = ~n19979 & ~n19981;
  assign n19983 = ~po34  & ~n19966;
  assign n19984 = ~n19974 & n19983;
  assign n19985 = ~n19982 & ~n19984;
  assign n19986 = ~n19976 & ~n19985;
  assign n19987 = po35  & ~n19986;
  assign n19988 = ~n19333 & ~n19341;
  assign n19989 = n19339 & n19988;
  assign n19990 = po3  & n19989;
  assign n19991 = po3  & n19988;
  assign n19992 = ~n19339 & ~n19991;
  assign n19993 = ~n19990 & ~n19992;
  assign n19994 = ~po35  & n19986;
  assign n19995 = ~n19993 & ~n19994;
  assign n19996 = ~n19987 & ~n19995;
  assign n19997 = po36  & ~n19996;
  assign n19998 = ~n19344 & ~n19351;
  assign n19999 = n19350 & n19998;
  assign n20000 = po3  & n19999;
  assign n20001 = po3  & n19998;
  assign n20002 = ~n19350 & ~n20001;
  assign n20003 = ~n20000 & ~n20002;
  assign n20004 = ~po36  & ~n19987;
  assign n20005 = ~n19995 & n20004;
  assign n20006 = ~n20003 & ~n20005;
  assign n20007 = ~n19997 & ~n20006;
  assign n20008 = po37  & ~n20007;
  assign n20009 = ~n19354 & ~n19362;
  assign n20010 = n19360 & n20009;
  assign n20011 = po3  & n20010;
  assign n20012 = po3  & n20009;
  assign n20013 = ~n19360 & ~n20012;
  assign n20014 = ~n20011 & ~n20013;
  assign n20015 = ~po37  & n20007;
  assign n20016 = ~n20014 & ~n20015;
  assign n20017 = ~n20008 & ~n20016;
  assign n20018 = po38  & ~n20017;
  assign n20019 = ~n19365 & ~n19372;
  assign n20020 = n19371 & n20019;
  assign n20021 = po3  & n20020;
  assign n20022 = po3  & n20019;
  assign n20023 = ~n19371 & ~n20022;
  assign n20024 = ~n20021 & ~n20023;
  assign n20025 = ~po38  & ~n20008;
  assign n20026 = ~n20016 & n20025;
  assign n20027 = ~n20024 & ~n20026;
  assign n20028 = ~n20018 & ~n20027;
  assign n20029 = po39  & ~n20028;
  assign n20030 = ~n19375 & ~n19383;
  assign n20031 = n19381 & n20030;
  assign n20032 = po3  & n20031;
  assign n20033 = po3  & n20030;
  assign n20034 = ~n19381 & ~n20033;
  assign n20035 = ~n20032 & ~n20034;
  assign n20036 = ~po39  & n20028;
  assign n20037 = ~n20035 & ~n20036;
  assign n20038 = ~n20029 & ~n20037;
  assign n20039 = po40  & ~n20038;
  assign n20040 = ~n19386 & ~n19393;
  assign n20041 = n19392 & n20040;
  assign n20042 = po3  & n20041;
  assign n20043 = po3  & n20040;
  assign n20044 = ~n19392 & ~n20043;
  assign n20045 = ~n20042 & ~n20044;
  assign n20046 = ~po40  & ~n20029;
  assign n20047 = ~n20037 & n20046;
  assign n20048 = ~n20045 & ~n20047;
  assign n20049 = ~n20039 & ~n20048;
  assign n20050 = po41  & ~n20049;
  assign n20051 = ~n19396 & ~n19404;
  assign n20052 = n19402 & n20051;
  assign n20053 = po3  & n20052;
  assign n20054 = po3  & n20051;
  assign n20055 = ~n19402 & ~n20054;
  assign n20056 = ~n20053 & ~n20055;
  assign n20057 = ~po41  & n20049;
  assign n20058 = ~n20056 & ~n20057;
  assign n20059 = ~n20050 & ~n20058;
  assign n20060 = po42  & ~n20059;
  assign n20061 = ~n19407 & ~n19414;
  assign n20062 = n19413 & n20061;
  assign n20063 = po3  & n20062;
  assign n20064 = po3  & n20061;
  assign n20065 = ~n19413 & ~n20064;
  assign n20066 = ~n20063 & ~n20065;
  assign n20067 = ~po42  & ~n20050;
  assign n20068 = ~n20058 & n20067;
  assign n20069 = ~n20066 & ~n20068;
  assign n20070 = ~n20060 & ~n20069;
  assign n20071 = po43  & ~n20070;
  assign n20072 = ~n19417 & ~n19425;
  assign n20073 = n19423 & n20072;
  assign n20074 = po3  & n20073;
  assign n20075 = po3  & n20072;
  assign n20076 = ~n19423 & ~n20075;
  assign n20077 = ~n20074 & ~n20076;
  assign n20078 = ~po43  & n20070;
  assign n20079 = ~n20077 & ~n20078;
  assign n20080 = ~n20071 & ~n20079;
  assign n20081 = po44  & ~n20080;
  assign n20082 = ~n19428 & ~n19435;
  assign n20083 = n19434 & n20082;
  assign n20084 = po3  & n20083;
  assign n20085 = po3  & n20082;
  assign n20086 = ~n19434 & ~n20085;
  assign n20087 = ~n20084 & ~n20086;
  assign n20088 = ~po44  & ~n20071;
  assign n20089 = ~n20079 & n20088;
  assign n20090 = ~n20087 & ~n20089;
  assign n20091 = ~n20081 & ~n20090;
  assign n20092 = po45  & ~n20091;
  assign n20093 = ~n19438 & ~n19446;
  assign n20094 = n19444 & n20093;
  assign n20095 = po3  & n20094;
  assign n20096 = po3  & n20093;
  assign n20097 = ~n19444 & ~n20096;
  assign n20098 = ~n20095 & ~n20097;
  assign n20099 = ~po45  & n20091;
  assign n20100 = ~n20098 & ~n20099;
  assign n20101 = ~n20092 & ~n20100;
  assign n20102 = po46  & ~n20101;
  assign n20103 = ~n19449 & ~n19456;
  assign n20104 = n19455 & n20103;
  assign n20105 = po3  & n20104;
  assign n20106 = po3  & n20103;
  assign n20107 = ~n19455 & ~n20106;
  assign n20108 = ~n20105 & ~n20107;
  assign n20109 = ~po46  & ~n20092;
  assign n20110 = ~n20100 & n20109;
  assign n20111 = ~n20108 & ~n20110;
  assign n20112 = ~n20102 & ~n20111;
  assign n20113 = po47  & ~n20112;
  assign n20114 = ~n19459 & ~n19467;
  assign n20115 = n19465 & n20114;
  assign n20116 = po3  & n20115;
  assign n20117 = po3  & n20114;
  assign n20118 = ~n19465 & ~n20117;
  assign n20119 = ~n20116 & ~n20118;
  assign n20120 = ~po47  & n20112;
  assign n20121 = ~n20119 & ~n20120;
  assign n20122 = ~n20113 & ~n20121;
  assign n20123 = po48  & ~n20122;
  assign n20124 = ~n19470 & ~n19477;
  assign n20125 = n19476 & n20124;
  assign n20126 = po3  & n20125;
  assign n20127 = po3  & n20124;
  assign n20128 = ~n19476 & ~n20127;
  assign n20129 = ~n20126 & ~n20128;
  assign n20130 = ~po48  & ~n20113;
  assign n20131 = ~n20121 & n20130;
  assign n20132 = ~n20129 & ~n20131;
  assign n20133 = ~n20123 & ~n20132;
  assign n20134 = po49  & ~n20133;
  assign n20135 = ~n19480 & ~n19488;
  assign n20136 = n19486 & n20135;
  assign n20137 = po3  & n20136;
  assign n20138 = po3  & n20135;
  assign n20139 = ~n19486 & ~n20138;
  assign n20140 = ~n20137 & ~n20139;
  assign n20141 = ~po49  & n20133;
  assign n20142 = ~n20140 & ~n20141;
  assign n20143 = ~n20134 & ~n20142;
  assign n20144 = po50  & ~n20143;
  assign n20145 = ~n19491 & ~n19498;
  assign n20146 = n19497 & n20145;
  assign n20147 = po3  & n20146;
  assign n20148 = po3  & n20145;
  assign n20149 = ~n19497 & ~n20148;
  assign n20150 = ~n20147 & ~n20149;
  assign n20151 = ~po50  & ~n20134;
  assign n20152 = ~n20142 & n20151;
  assign n20153 = ~n20150 & ~n20152;
  assign n20154 = ~n20144 & ~n20153;
  assign n20155 = po51  & ~n20154;
  assign n20156 = ~n19501 & ~n19509;
  assign n20157 = n19507 & n20156;
  assign n20158 = po3  & n20157;
  assign n20159 = po3  & n20156;
  assign n20160 = ~n19507 & ~n20159;
  assign n20161 = ~n20158 & ~n20160;
  assign n20162 = ~po51  & n20154;
  assign n20163 = ~n20161 & ~n20162;
  assign n20164 = ~n20155 & ~n20163;
  assign n20165 = po52  & ~n20164;
  assign n20166 = ~n19512 & ~n19519;
  assign n20167 = n19518 & n20166;
  assign n20168 = po3  & n20167;
  assign n20169 = po3  & n20166;
  assign n20170 = ~n19518 & ~n20169;
  assign n20171 = ~n20168 & ~n20170;
  assign n20172 = ~po52  & ~n20155;
  assign n20173 = ~n20163 & n20172;
  assign n20174 = ~n20171 & ~n20173;
  assign n20175 = ~n20165 & ~n20174;
  assign n20176 = po53  & ~n20175;
  assign n20177 = ~n19522 & ~n19530;
  assign n20178 = n19528 & n20177;
  assign n20179 = po3  & n20178;
  assign n20180 = po3  & n20177;
  assign n20181 = ~n19528 & ~n20180;
  assign n20182 = ~n20179 & ~n20181;
  assign n20183 = ~po53  & n20175;
  assign n20184 = ~n20182 & ~n20183;
  assign n20185 = ~n20176 & ~n20184;
  assign n20186 = po54  & ~n20185;
  assign n20187 = ~n19533 & ~n19540;
  assign n20188 = n19539 & n20187;
  assign n20189 = po3  & n20188;
  assign n20190 = po3  & n20187;
  assign n20191 = ~n19539 & ~n20190;
  assign n20192 = ~n20189 & ~n20191;
  assign n20193 = ~po54  & ~n20176;
  assign n20194 = ~n20184 & n20193;
  assign n20195 = ~n20192 & ~n20194;
  assign n20196 = ~n20186 & ~n20195;
  assign n20197 = po55  & ~n20196;
  assign n20198 = ~n19543 & ~n19551;
  assign n20199 = n19549 & n20198;
  assign n20200 = po3  & n20199;
  assign n20201 = po3  & n20198;
  assign n20202 = ~n19549 & ~n20201;
  assign n20203 = ~n20200 & ~n20202;
  assign n20204 = ~po55  & n20196;
  assign n20205 = ~n20203 & ~n20204;
  assign n20206 = ~n20197 & ~n20205;
  assign n20207 = po56  & ~n20206;
  assign n20208 = ~n19554 & ~n19561;
  assign n20209 = n19560 & n20208;
  assign n20210 = po3  & n20209;
  assign n20211 = po3  & n20208;
  assign n20212 = ~n19560 & ~n20211;
  assign n20213 = ~n20210 & ~n20212;
  assign n20214 = ~po56  & ~n20197;
  assign n20215 = ~n20205 & n20214;
  assign n20216 = ~n20213 & ~n20215;
  assign n20217 = ~n20207 & ~n20216;
  assign n20218 = po57  & ~n20217;
  assign n20219 = ~n19564 & ~n19572;
  assign n20220 = n19570 & n20219;
  assign n20221 = po3  & n20220;
  assign n20222 = po3  & n20219;
  assign n20223 = ~n19570 & ~n20222;
  assign n20224 = ~n20221 & ~n20223;
  assign n20225 = ~po57  & n20217;
  assign n20226 = ~n20224 & ~n20225;
  assign n20227 = ~n20218 & ~n20226;
  assign n20228 = po58  & ~n20227;
  assign n20229 = ~n19575 & ~n19582;
  assign n20230 = n19581 & n20229;
  assign n20231 = po3  & n20230;
  assign n20232 = po3  & n20229;
  assign n20233 = ~n19581 & ~n20232;
  assign n20234 = ~n20231 & ~n20233;
  assign n20235 = ~po58  & ~n20218;
  assign n20236 = ~n20226 & n20235;
  assign n20237 = ~n20234 & ~n20236;
  assign n20238 = ~n20228 & ~n20237;
  assign n20239 = po59  & ~n20238;
  assign n20240 = ~n19585 & ~n19593;
  assign n20241 = n19591 & n20240;
  assign n20242 = po3  & n20241;
  assign n20243 = po3  & n20240;
  assign n20244 = ~n19591 & ~n20243;
  assign n20245 = ~n20242 & ~n20244;
  assign n20246 = ~po59  & n20238;
  assign n20247 = ~n20245 & ~n20246;
  assign n20248 = ~n20239 & ~n20247;
  assign n20249 = po60  & ~n20248;
  assign n20250 = ~n19596 & ~n19603;
  assign n20251 = n19602 & n20250;
  assign n20252 = po3  & n20251;
  assign n20253 = po3  & n20250;
  assign n20254 = ~n19602 & ~n20253;
  assign n20255 = ~n20252 & ~n20254;
  assign n20256 = ~po60  & ~n20239;
  assign n20257 = ~n20247 & n20256;
  assign n20258 = ~n20255 & ~n20257;
  assign n20259 = ~n20249 & ~n20258;
  assign n20260 = po61  & ~n20259;
  assign n20261 = ~n19606 & ~n19614;
  assign n20262 = n19612 & n20261;
  assign n20263 = po3  & n20262;
  assign n20264 = po3  & n20261;
  assign n20265 = ~n19612 & ~n20264;
  assign n20266 = ~n20263 & ~n20265;
  assign n20267 = ~po61  & n20259;
  assign n20268 = ~n20266 & ~n20267;
  assign n20269 = ~n20260 & ~n20268;
  assign n20270 = po62  & ~n20269;
  assign n20271 = ~po62  & ~n20260;
  assign n20272 = ~n20268 & n20271;
  assign n20273 = ~n19617 & ~n19624;
  assign n20274 = n19623 & n20273;
  assign n20275 = po3  & n20274;
  assign n20276 = po3  & n20273;
  assign n20277 = ~n19623 & ~n20276;
  assign n20278 = ~n20275 & ~n20277;
  assign n20279 = ~n20272 & ~n20278;
  assign n20280 = ~n20270 & ~n20279;
  assign n20281 = ~n19627 & ~n19635;
  assign n20282 = po3  & n20281;
  assign n20283 = ~n19633 & ~n20282;
  assign n20284 = n19633 & n20282;
  assign n20285 = ~n20283 & ~n20284;
  assign n20286 = ~n19637 & ~n19642;
  assign n20287 = po3  & n20286;
  assign n20288 = ~n19653 & ~n20287;
  assign n20289 = ~n20285 & n20288;
  assign n20290 = ~n20280 & n20289;
  assign n20291 = ~po63  & ~n20290;
  assign n20292 = ~n19642 & po3 ;
  assign n20293 = n19637 & ~n20292;
  assign n20294 = po63  & ~n20286;
  assign n20295 = ~n20293 & n20294;
  assign n20296 = n20280 & n20285;
  assign n20297 = ~n20295 & ~n20296;
  assign po2  = n20291 | ~n20297;
  assign n20299 = ~n20249 & ~n20257;
  assign n20300 = n20255 & n20299;
  assign n20301 = po2  & n20300;
  assign n20302 = po2  & n20299;
  assign n20303 = ~n20255 & ~n20302;
  assign n20304 = ~n20301 & ~n20303;
  assign n20305 = pi4  & po2 ;
  assign n20306 = ~pi2  & ~pi3 ;
  assign n20307 = ~pi4  & n20306;
  assign n20308 = ~n20305 & ~n20307;
  assign n20309 = po3  & ~n20308;
  assign n20310 = ~n19652 & ~n20307;
  assign n20311 = ~n19653 & n20310;
  assign n20312 = ~n19648 & n20311;
  assign n20313 = ~n20305 & n20312;
  assign n20314 = ~pi4  & po2 ;
  assign n20315 = pi5  & ~n20314;
  assign n20316 = n19657 & po2 ;
  assign n20317 = ~n20315 & ~n20316;
  assign n20318 = ~n20313 & n20317;
  assign n20319 = ~n20309 & ~n20318;
  assign n20320 = po4  & ~n20319;
  assign n20321 = ~po4  & ~n20309;
  assign n20322 = ~n20318 & n20321;
  assign n20323 = po3  & ~n20295;
  assign n20324 = ~n20296 & n20323;
  assign n20325 = ~n20291 & n20324;
  assign n20326 = ~n20316 & ~n20325;
  assign n20327 = pi6  & ~n20326;
  assign n20328 = ~pi6  & n20326;
  assign n20329 = ~n20327 & ~n20328;
  assign n20330 = ~n20322 & ~n20329;
  assign n20331 = ~n20320 & ~n20330;
  assign n20332 = po5  & ~n20331;
  assign n20333 = ~n19660 & ~n19664;
  assign n20334 = ~n19668 & n20333;
  assign n20335 = po2  & n20334;
  assign n20336 = po2  & n20333;
  assign n20337 = n19668 & ~n20336;
  assign n20338 = ~n20335 & ~n20337;
  assign n20339 = ~po5  & n20331;
  assign n20340 = ~n20338 & ~n20339;
  assign n20341 = ~n20332 & ~n20340;
  assign n20342 = po6  & ~n20341;
  assign n20343 = ~n19671 & ~n19679;
  assign n20344 = ~n19680 & n20343;
  assign n20345 = po2  & n20344;
  assign n20346 = po2  & n20343;
  assign n20347 = ~n19678 & ~n20346;
  assign n20348 = ~n20345 & ~n20347;
  assign n20349 = ~po6  & ~n20332;
  assign n20350 = ~n20340 & n20349;
  assign n20351 = ~n20348 & ~n20350;
  assign n20352 = ~n20342 & ~n20351;
  assign n20353 = po7  & ~n20352;
  assign n20354 = ~n19682 & ~n19690;
  assign n20355 = n19688 & n20354;
  assign n20356 = po2  & n20355;
  assign n20357 = po2  & n20354;
  assign n20358 = ~n19688 & ~n20357;
  assign n20359 = ~n20356 & ~n20358;
  assign n20360 = ~po7  & n20352;
  assign n20361 = ~n20359 & ~n20360;
  assign n20362 = ~n20353 & ~n20361;
  assign n20363 = po8  & ~n20362;
  assign n20364 = ~n19693 & ~n19700;
  assign n20365 = n19699 & n20364;
  assign n20366 = po2  & n20365;
  assign n20367 = po2  & n20364;
  assign n20368 = ~n19699 & ~n20367;
  assign n20369 = ~n20366 & ~n20368;
  assign n20370 = ~po8  & ~n20353;
  assign n20371 = ~n20361 & n20370;
  assign n20372 = ~n20369 & ~n20371;
  assign n20373 = ~n20363 & ~n20372;
  assign n20374 = po9  & ~n20373;
  assign n20375 = ~n19703 & ~n19711;
  assign n20376 = n19709 & n20375;
  assign n20377 = po2  & n20376;
  assign n20378 = po2  & n20375;
  assign n20379 = ~n19709 & ~n20378;
  assign n20380 = ~n20377 & ~n20379;
  assign n20381 = ~po9  & n20373;
  assign n20382 = ~n20380 & ~n20381;
  assign n20383 = ~n20374 & ~n20382;
  assign n20384 = po10  & ~n20383;
  assign n20385 = ~n19714 & ~n19721;
  assign n20386 = n19720 & n20385;
  assign n20387 = po2  & n20386;
  assign n20388 = po2  & n20385;
  assign n20389 = ~n19720 & ~n20388;
  assign n20390 = ~n20387 & ~n20389;
  assign n20391 = ~po10  & ~n20374;
  assign n20392 = ~n20382 & n20391;
  assign n20393 = ~n20390 & ~n20392;
  assign n20394 = ~n20384 & ~n20393;
  assign n20395 = po11  & ~n20394;
  assign n20396 = ~n19724 & ~n19732;
  assign n20397 = n19730 & n20396;
  assign n20398 = po2  & n20397;
  assign n20399 = po2  & n20396;
  assign n20400 = ~n19730 & ~n20399;
  assign n20401 = ~n20398 & ~n20400;
  assign n20402 = ~po11  & n20394;
  assign n20403 = ~n20401 & ~n20402;
  assign n20404 = ~n20395 & ~n20403;
  assign n20405 = po12  & ~n20404;
  assign n20406 = ~n19735 & ~n19742;
  assign n20407 = n19741 & n20406;
  assign n20408 = po2  & n20407;
  assign n20409 = po2  & n20406;
  assign n20410 = ~n19741 & ~n20409;
  assign n20411 = ~n20408 & ~n20410;
  assign n20412 = ~po12  & ~n20395;
  assign n20413 = ~n20403 & n20412;
  assign n20414 = ~n20411 & ~n20413;
  assign n20415 = ~n20405 & ~n20414;
  assign n20416 = po13  & ~n20415;
  assign n20417 = ~n19745 & ~n19753;
  assign n20418 = n19751 & n20417;
  assign n20419 = po2  & n20418;
  assign n20420 = po2  & n20417;
  assign n20421 = ~n19751 & ~n20420;
  assign n20422 = ~n20419 & ~n20421;
  assign n20423 = ~po13  & n20415;
  assign n20424 = ~n20422 & ~n20423;
  assign n20425 = ~n20416 & ~n20424;
  assign n20426 = po14  & ~n20425;
  assign n20427 = ~n19756 & ~n19763;
  assign n20428 = n19762 & n20427;
  assign n20429 = po2  & n20428;
  assign n20430 = po2  & n20427;
  assign n20431 = ~n19762 & ~n20430;
  assign n20432 = ~n20429 & ~n20431;
  assign n20433 = ~po14  & ~n20416;
  assign n20434 = ~n20424 & n20433;
  assign n20435 = ~n20432 & ~n20434;
  assign n20436 = ~n20426 & ~n20435;
  assign n20437 = po15  & ~n20436;
  assign n20438 = ~n19766 & ~n19774;
  assign n20439 = n19772 & n20438;
  assign n20440 = po2  & n20439;
  assign n20441 = po2  & n20438;
  assign n20442 = ~n19772 & ~n20441;
  assign n20443 = ~n20440 & ~n20442;
  assign n20444 = ~po15  & n20436;
  assign n20445 = ~n20443 & ~n20444;
  assign n20446 = ~n20437 & ~n20445;
  assign n20447 = po16  & ~n20446;
  assign n20448 = ~n19777 & ~n19784;
  assign n20449 = n19783 & n20448;
  assign n20450 = po2  & n20449;
  assign n20451 = po2  & n20448;
  assign n20452 = ~n19783 & ~n20451;
  assign n20453 = ~n20450 & ~n20452;
  assign n20454 = ~po16  & ~n20437;
  assign n20455 = ~n20445 & n20454;
  assign n20456 = ~n20453 & ~n20455;
  assign n20457 = ~n20447 & ~n20456;
  assign n20458 = po17  & ~n20457;
  assign n20459 = ~n19787 & ~n19795;
  assign n20460 = n19793 & n20459;
  assign n20461 = po2  & n20460;
  assign n20462 = po2  & n20459;
  assign n20463 = ~n19793 & ~n20462;
  assign n20464 = ~n20461 & ~n20463;
  assign n20465 = ~po17  & n20457;
  assign n20466 = ~n20464 & ~n20465;
  assign n20467 = ~n20458 & ~n20466;
  assign n20468 = po18  & ~n20467;
  assign n20469 = ~n19798 & ~n19805;
  assign n20470 = n19804 & n20469;
  assign n20471 = po2  & n20470;
  assign n20472 = po2  & n20469;
  assign n20473 = ~n19804 & ~n20472;
  assign n20474 = ~n20471 & ~n20473;
  assign n20475 = ~po18  & ~n20458;
  assign n20476 = ~n20466 & n20475;
  assign n20477 = ~n20474 & ~n20476;
  assign n20478 = ~n20468 & ~n20477;
  assign n20479 = po19  & ~n20478;
  assign n20480 = ~n19808 & ~n19816;
  assign n20481 = n19814 & n20480;
  assign n20482 = po2  & n20481;
  assign n20483 = po2  & n20480;
  assign n20484 = ~n19814 & ~n20483;
  assign n20485 = ~n20482 & ~n20484;
  assign n20486 = ~po19  & n20478;
  assign n20487 = ~n20485 & ~n20486;
  assign n20488 = ~n20479 & ~n20487;
  assign n20489 = po20  & ~n20488;
  assign n20490 = ~n19819 & ~n19826;
  assign n20491 = n19825 & n20490;
  assign n20492 = po2  & n20491;
  assign n20493 = po2  & n20490;
  assign n20494 = ~n19825 & ~n20493;
  assign n20495 = ~n20492 & ~n20494;
  assign n20496 = ~po20  & ~n20479;
  assign n20497 = ~n20487 & n20496;
  assign n20498 = ~n20495 & ~n20497;
  assign n20499 = ~n20489 & ~n20498;
  assign n20500 = po21  & ~n20499;
  assign n20501 = ~n19829 & ~n19837;
  assign n20502 = n19835 & n20501;
  assign n20503 = po2  & n20502;
  assign n20504 = po2  & n20501;
  assign n20505 = ~n19835 & ~n20504;
  assign n20506 = ~n20503 & ~n20505;
  assign n20507 = ~po21  & n20499;
  assign n20508 = ~n20506 & ~n20507;
  assign n20509 = ~n20500 & ~n20508;
  assign n20510 = po22  & ~n20509;
  assign n20511 = ~n19840 & ~n19847;
  assign n20512 = n19846 & n20511;
  assign n20513 = po2  & n20512;
  assign n20514 = po2  & n20511;
  assign n20515 = ~n19846 & ~n20514;
  assign n20516 = ~n20513 & ~n20515;
  assign n20517 = ~po22  & ~n20500;
  assign n20518 = ~n20508 & n20517;
  assign n20519 = ~n20516 & ~n20518;
  assign n20520 = ~n20510 & ~n20519;
  assign n20521 = po23  & ~n20520;
  assign n20522 = ~n19850 & ~n19858;
  assign n20523 = n19856 & n20522;
  assign n20524 = po2  & n20523;
  assign n20525 = po2  & n20522;
  assign n20526 = ~n19856 & ~n20525;
  assign n20527 = ~n20524 & ~n20526;
  assign n20528 = ~po23  & n20520;
  assign n20529 = ~n20527 & ~n20528;
  assign n20530 = ~n20521 & ~n20529;
  assign n20531 = po24  & ~n20530;
  assign n20532 = ~n19861 & ~n19868;
  assign n20533 = n19867 & n20532;
  assign n20534 = po2  & n20533;
  assign n20535 = po2  & n20532;
  assign n20536 = ~n19867 & ~n20535;
  assign n20537 = ~n20534 & ~n20536;
  assign n20538 = ~po24  & ~n20521;
  assign n20539 = ~n20529 & n20538;
  assign n20540 = ~n20537 & ~n20539;
  assign n20541 = ~n20531 & ~n20540;
  assign n20542 = po25  & ~n20541;
  assign n20543 = ~n19871 & ~n19879;
  assign n20544 = n19877 & n20543;
  assign n20545 = po2  & n20544;
  assign n20546 = po2  & n20543;
  assign n20547 = ~n19877 & ~n20546;
  assign n20548 = ~n20545 & ~n20547;
  assign n20549 = ~po25  & n20541;
  assign n20550 = ~n20548 & ~n20549;
  assign n20551 = ~n20542 & ~n20550;
  assign n20552 = po26  & ~n20551;
  assign n20553 = ~n19882 & ~n19889;
  assign n20554 = n19888 & n20553;
  assign n20555 = po2  & n20554;
  assign n20556 = po2  & n20553;
  assign n20557 = ~n19888 & ~n20556;
  assign n20558 = ~n20555 & ~n20557;
  assign n20559 = ~po26  & ~n20542;
  assign n20560 = ~n20550 & n20559;
  assign n20561 = ~n20558 & ~n20560;
  assign n20562 = ~n20552 & ~n20561;
  assign n20563 = po27  & ~n20562;
  assign n20564 = ~n19892 & ~n19900;
  assign n20565 = n19898 & n20564;
  assign n20566 = po2  & n20565;
  assign n20567 = po2  & n20564;
  assign n20568 = ~n19898 & ~n20567;
  assign n20569 = ~n20566 & ~n20568;
  assign n20570 = ~po27  & n20562;
  assign n20571 = ~n20569 & ~n20570;
  assign n20572 = ~n20563 & ~n20571;
  assign n20573 = po28  & ~n20572;
  assign n20574 = ~n19903 & ~n19910;
  assign n20575 = n19909 & n20574;
  assign n20576 = po2  & n20575;
  assign n20577 = po2  & n20574;
  assign n20578 = ~n19909 & ~n20577;
  assign n20579 = ~n20576 & ~n20578;
  assign n20580 = ~po28  & ~n20563;
  assign n20581 = ~n20571 & n20580;
  assign n20582 = ~n20579 & ~n20581;
  assign n20583 = ~n20573 & ~n20582;
  assign n20584 = po29  & ~n20583;
  assign n20585 = ~n19913 & ~n19921;
  assign n20586 = n19919 & n20585;
  assign n20587 = po2  & n20586;
  assign n20588 = po2  & n20585;
  assign n20589 = ~n19919 & ~n20588;
  assign n20590 = ~n20587 & ~n20589;
  assign n20591 = ~po29  & n20583;
  assign n20592 = ~n20590 & ~n20591;
  assign n20593 = ~n20584 & ~n20592;
  assign n20594 = po30  & ~n20593;
  assign n20595 = ~n19924 & ~n19931;
  assign n20596 = n19930 & n20595;
  assign n20597 = po2  & n20596;
  assign n20598 = po2  & n20595;
  assign n20599 = ~n19930 & ~n20598;
  assign n20600 = ~n20597 & ~n20599;
  assign n20601 = ~po30  & ~n20584;
  assign n20602 = ~n20592 & n20601;
  assign n20603 = ~n20600 & ~n20602;
  assign n20604 = ~n20594 & ~n20603;
  assign n20605 = po31  & ~n20604;
  assign n20606 = ~n19934 & ~n19942;
  assign n20607 = n19940 & n20606;
  assign n20608 = po2  & n20607;
  assign n20609 = po2  & n20606;
  assign n20610 = ~n19940 & ~n20609;
  assign n20611 = ~n20608 & ~n20610;
  assign n20612 = ~po31  & n20604;
  assign n20613 = ~n20611 & ~n20612;
  assign n20614 = ~n20605 & ~n20613;
  assign n20615 = po32  & ~n20614;
  assign n20616 = ~n19945 & ~n19952;
  assign n20617 = n19951 & n20616;
  assign n20618 = po2  & n20617;
  assign n20619 = po2  & n20616;
  assign n20620 = ~n19951 & ~n20619;
  assign n20621 = ~n20618 & ~n20620;
  assign n20622 = ~po32  & ~n20605;
  assign n20623 = ~n20613 & n20622;
  assign n20624 = ~n20621 & ~n20623;
  assign n20625 = ~n20615 & ~n20624;
  assign n20626 = po33  & ~n20625;
  assign n20627 = ~n19955 & ~n19963;
  assign n20628 = n19961 & n20627;
  assign n20629 = po2  & n20628;
  assign n20630 = po2  & n20627;
  assign n20631 = ~n19961 & ~n20630;
  assign n20632 = ~n20629 & ~n20631;
  assign n20633 = ~po33  & n20625;
  assign n20634 = ~n20632 & ~n20633;
  assign n20635 = ~n20626 & ~n20634;
  assign n20636 = po34  & ~n20635;
  assign n20637 = ~n19966 & ~n19973;
  assign n20638 = n19972 & n20637;
  assign n20639 = po2  & n20638;
  assign n20640 = po2  & n20637;
  assign n20641 = ~n19972 & ~n20640;
  assign n20642 = ~n20639 & ~n20641;
  assign n20643 = ~po34  & ~n20626;
  assign n20644 = ~n20634 & n20643;
  assign n20645 = ~n20642 & ~n20644;
  assign n20646 = ~n20636 & ~n20645;
  assign n20647 = po35  & ~n20646;
  assign n20648 = ~n19976 & ~n19984;
  assign n20649 = n19982 & n20648;
  assign n20650 = po2  & n20649;
  assign n20651 = po2  & n20648;
  assign n20652 = ~n19982 & ~n20651;
  assign n20653 = ~n20650 & ~n20652;
  assign n20654 = ~po35  & n20646;
  assign n20655 = ~n20653 & ~n20654;
  assign n20656 = ~n20647 & ~n20655;
  assign n20657 = po36  & ~n20656;
  assign n20658 = ~n19987 & ~n19994;
  assign n20659 = n19993 & n20658;
  assign n20660 = po2  & n20659;
  assign n20661 = po2  & n20658;
  assign n20662 = ~n19993 & ~n20661;
  assign n20663 = ~n20660 & ~n20662;
  assign n20664 = ~po36  & ~n20647;
  assign n20665 = ~n20655 & n20664;
  assign n20666 = ~n20663 & ~n20665;
  assign n20667 = ~n20657 & ~n20666;
  assign n20668 = po37  & ~n20667;
  assign n20669 = ~n19997 & ~n20005;
  assign n20670 = n20003 & n20669;
  assign n20671 = po2  & n20670;
  assign n20672 = po2  & n20669;
  assign n20673 = ~n20003 & ~n20672;
  assign n20674 = ~n20671 & ~n20673;
  assign n20675 = ~po37  & n20667;
  assign n20676 = ~n20674 & ~n20675;
  assign n20677 = ~n20668 & ~n20676;
  assign n20678 = po38  & ~n20677;
  assign n20679 = ~n20008 & ~n20015;
  assign n20680 = n20014 & n20679;
  assign n20681 = po2  & n20680;
  assign n20682 = po2  & n20679;
  assign n20683 = ~n20014 & ~n20682;
  assign n20684 = ~n20681 & ~n20683;
  assign n20685 = ~po38  & ~n20668;
  assign n20686 = ~n20676 & n20685;
  assign n20687 = ~n20684 & ~n20686;
  assign n20688 = ~n20678 & ~n20687;
  assign n20689 = po39  & ~n20688;
  assign n20690 = ~n20018 & ~n20026;
  assign n20691 = n20024 & n20690;
  assign n20692 = po2  & n20691;
  assign n20693 = po2  & n20690;
  assign n20694 = ~n20024 & ~n20693;
  assign n20695 = ~n20692 & ~n20694;
  assign n20696 = ~po39  & n20688;
  assign n20697 = ~n20695 & ~n20696;
  assign n20698 = ~n20689 & ~n20697;
  assign n20699 = po40  & ~n20698;
  assign n20700 = ~n20029 & ~n20036;
  assign n20701 = n20035 & n20700;
  assign n20702 = po2  & n20701;
  assign n20703 = po2  & n20700;
  assign n20704 = ~n20035 & ~n20703;
  assign n20705 = ~n20702 & ~n20704;
  assign n20706 = ~po40  & ~n20689;
  assign n20707 = ~n20697 & n20706;
  assign n20708 = ~n20705 & ~n20707;
  assign n20709 = ~n20699 & ~n20708;
  assign n20710 = po41  & ~n20709;
  assign n20711 = ~n20039 & ~n20047;
  assign n20712 = n20045 & n20711;
  assign n20713 = po2  & n20712;
  assign n20714 = po2  & n20711;
  assign n20715 = ~n20045 & ~n20714;
  assign n20716 = ~n20713 & ~n20715;
  assign n20717 = ~po41  & n20709;
  assign n20718 = ~n20716 & ~n20717;
  assign n20719 = ~n20710 & ~n20718;
  assign n20720 = po42  & ~n20719;
  assign n20721 = ~n20050 & ~n20057;
  assign n20722 = n20056 & n20721;
  assign n20723 = po2  & n20722;
  assign n20724 = po2  & n20721;
  assign n20725 = ~n20056 & ~n20724;
  assign n20726 = ~n20723 & ~n20725;
  assign n20727 = ~po42  & ~n20710;
  assign n20728 = ~n20718 & n20727;
  assign n20729 = ~n20726 & ~n20728;
  assign n20730 = ~n20720 & ~n20729;
  assign n20731 = po43  & ~n20730;
  assign n20732 = ~n20060 & ~n20068;
  assign n20733 = n20066 & n20732;
  assign n20734 = po2  & n20733;
  assign n20735 = po2  & n20732;
  assign n20736 = ~n20066 & ~n20735;
  assign n20737 = ~n20734 & ~n20736;
  assign n20738 = ~po43  & n20730;
  assign n20739 = ~n20737 & ~n20738;
  assign n20740 = ~n20731 & ~n20739;
  assign n20741 = po44  & ~n20740;
  assign n20742 = ~n20071 & ~n20078;
  assign n20743 = n20077 & n20742;
  assign n20744 = po2  & n20743;
  assign n20745 = po2  & n20742;
  assign n20746 = ~n20077 & ~n20745;
  assign n20747 = ~n20744 & ~n20746;
  assign n20748 = ~po44  & ~n20731;
  assign n20749 = ~n20739 & n20748;
  assign n20750 = ~n20747 & ~n20749;
  assign n20751 = ~n20741 & ~n20750;
  assign n20752 = po45  & ~n20751;
  assign n20753 = ~n20081 & ~n20089;
  assign n20754 = n20087 & n20753;
  assign n20755 = po2  & n20754;
  assign n20756 = po2  & n20753;
  assign n20757 = ~n20087 & ~n20756;
  assign n20758 = ~n20755 & ~n20757;
  assign n20759 = ~po45  & n20751;
  assign n20760 = ~n20758 & ~n20759;
  assign n20761 = ~n20752 & ~n20760;
  assign n20762 = po46  & ~n20761;
  assign n20763 = ~n20092 & ~n20099;
  assign n20764 = n20098 & n20763;
  assign n20765 = po2  & n20764;
  assign n20766 = po2  & n20763;
  assign n20767 = ~n20098 & ~n20766;
  assign n20768 = ~n20765 & ~n20767;
  assign n20769 = ~po46  & ~n20752;
  assign n20770 = ~n20760 & n20769;
  assign n20771 = ~n20768 & ~n20770;
  assign n20772 = ~n20762 & ~n20771;
  assign n20773 = po47  & ~n20772;
  assign n20774 = ~n20102 & ~n20110;
  assign n20775 = n20108 & n20774;
  assign n20776 = po2  & n20775;
  assign n20777 = po2  & n20774;
  assign n20778 = ~n20108 & ~n20777;
  assign n20779 = ~n20776 & ~n20778;
  assign n20780 = ~po47  & n20772;
  assign n20781 = ~n20779 & ~n20780;
  assign n20782 = ~n20773 & ~n20781;
  assign n20783 = po48  & ~n20782;
  assign n20784 = ~n20113 & ~n20120;
  assign n20785 = n20119 & n20784;
  assign n20786 = po2  & n20785;
  assign n20787 = po2  & n20784;
  assign n20788 = ~n20119 & ~n20787;
  assign n20789 = ~n20786 & ~n20788;
  assign n20790 = ~po48  & ~n20773;
  assign n20791 = ~n20781 & n20790;
  assign n20792 = ~n20789 & ~n20791;
  assign n20793 = ~n20783 & ~n20792;
  assign n20794 = po49  & ~n20793;
  assign n20795 = ~n20123 & ~n20131;
  assign n20796 = n20129 & n20795;
  assign n20797 = po2  & n20796;
  assign n20798 = po2  & n20795;
  assign n20799 = ~n20129 & ~n20798;
  assign n20800 = ~n20797 & ~n20799;
  assign n20801 = ~po49  & n20793;
  assign n20802 = ~n20800 & ~n20801;
  assign n20803 = ~n20794 & ~n20802;
  assign n20804 = po50  & ~n20803;
  assign n20805 = ~n20134 & ~n20141;
  assign n20806 = n20140 & n20805;
  assign n20807 = po2  & n20806;
  assign n20808 = po2  & n20805;
  assign n20809 = ~n20140 & ~n20808;
  assign n20810 = ~n20807 & ~n20809;
  assign n20811 = ~po50  & ~n20794;
  assign n20812 = ~n20802 & n20811;
  assign n20813 = ~n20810 & ~n20812;
  assign n20814 = ~n20804 & ~n20813;
  assign n20815 = po51  & ~n20814;
  assign n20816 = ~n20144 & ~n20152;
  assign n20817 = n20150 & n20816;
  assign n20818 = po2  & n20817;
  assign n20819 = po2  & n20816;
  assign n20820 = ~n20150 & ~n20819;
  assign n20821 = ~n20818 & ~n20820;
  assign n20822 = ~po51  & n20814;
  assign n20823 = ~n20821 & ~n20822;
  assign n20824 = ~n20815 & ~n20823;
  assign n20825 = po52  & ~n20824;
  assign n20826 = ~n20155 & ~n20162;
  assign n20827 = n20161 & n20826;
  assign n20828 = po2  & n20827;
  assign n20829 = po2  & n20826;
  assign n20830 = ~n20161 & ~n20829;
  assign n20831 = ~n20828 & ~n20830;
  assign n20832 = ~po52  & ~n20815;
  assign n20833 = ~n20823 & n20832;
  assign n20834 = ~n20831 & ~n20833;
  assign n20835 = ~n20825 & ~n20834;
  assign n20836 = po53  & ~n20835;
  assign n20837 = ~n20165 & ~n20173;
  assign n20838 = n20171 & n20837;
  assign n20839 = po2  & n20838;
  assign n20840 = po2  & n20837;
  assign n20841 = ~n20171 & ~n20840;
  assign n20842 = ~n20839 & ~n20841;
  assign n20843 = ~po53  & n20835;
  assign n20844 = ~n20842 & ~n20843;
  assign n20845 = ~n20836 & ~n20844;
  assign n20846 = po54  & ~n20845;
  assign n20847 = ~n20176 & ~n20183;
  assign n20848 = n20182 & n20847;
  assign n20849 = po2  & n20848;
  assign n20850 = po2  & n20847;
  assign n20851 = ~n20182 & ~n20850;
  assign n20852 = ~n20849 & ~n20851;
  assign n20853 = ~po54  & ~n20836;
  assign n20854 = ~n20844 & n20853;
  assign n20855 = ~n20852 & ~n20854;
  assign n20856 = ~n20846 & ~n20855;
  assign n20857 = po55  & ~n20856;
  assign n20858 = ~n20186 & ~n20194;
  assign n20859 = n20192 & n20858;
  assign n20860 = po2  & n20859;
  assign n20861 = po2  & n20858;
  assign n20862 = ~n20192 & ~n20861;
  assign n20863 = ~n20860 & ~n20862;
  assign n20864 = ~po55  & n20856;
  assign n20865 = ~n20863 & ~n20864;
  assign n20866 = ~n20857 & ~n20865;
  assign n20867 = po56  & ~n20866;
  assign n20868 = ~n20197 & ~n20204;
  assign n20869 = n20203 & n20868;
  assign n20870 = po2  & n20869;
  assign n20871 = po2  & n20868;
  assign n20872 = ~n20203 & ~n20871;
  assign n20873 = ~n20870 & ~n20872;
  assign n20874 = ~po56  & ~n20857;
  assign n20875 = ~n20865 & n20874;
  assign n20876 = ~n20873 & ~n20875;
  assign n20877 = ~n20867 & ~n20876;
  assign n20878 = po57  & ~n20877;
  assign n20879 = ~n20207 & ~n20215;
  assign n20880 = n20213 & n20879;
  assign n20881 = po2  & n20880;
  assign n20882 = po2  & n20879;
  assign n20883 = ~n20213 & ~n20882;
  assign n20884 = ~n20881 & ~n20883;
  assign n20885 = ~po57  & n20877;
  assign n20886 = ~n20884 & ~n20885;
  assign n20887 = ~n20878 & ~n20886;
  assign n20888 = po58  & ~n20887;
  assign n20889 = ~n20218 & ~n20225;
  assign n20890 = n20224 & n20889;
  assign n20891 = po2  & n20890;
  assign n20892 = po2  & n20889;
  assign n20893 = ~n20224 & ~n20892;
  assign n20894 = ~n20891 & ~n20893;
  assign n20895 = ~po58  & ~n20878;
  assign n20896 = ~n20886 & n20895;
  assign n20897 = ~n20894 & ~n20896;
  assign n20898 = ~n20888 & ~n20897;
  assign n20899 = po59  & ~n20898;
  assign n20900 = ~n20228 & ~n20236;
  assign n20901 = n20234 & n20900;
  assign n20902 = po2  & n20901;
  assign n20903 = po2  & n20900;
  assign n20904 = ~n20234 & ~n20903;
  assign n20905 = ~n20902 & ~n20904;
  assign n20906 = ~po59  & n20898;
  assign n20907 = ~n20905 & ~n20906;
  assign n20908 = ~n20899 & ~n20907;
  assign n20909 = po60  & ~n20908;
  assign n20910 = ~n20239 & ~n20246;
  assign n20911 = n20245 & n20910;
  assign n20912 = po2  & n20911;
  assign n20913 = po2  & n20910;
  assign n20914 = ~n20245 & ~n20913;
  assign n20915 = ~n20912 & ~n20914;
  assign n20916 = ~po60  & ~n20899;
  assign n20917 = ~n20907 & n20916;
  assign n20918 = ~n20915 & ~n20917;
  assign n20919 = ~n20909 & ~n20918;
  assign n20920 = po61  & ~n20919;
  assign n20921 = ~po61  & n20919;
  assign n20922 = ~n20304 & ~n20921;
  assign n20923 = ~n20920 & ~n20922;
  assign n20924 = po62  & ~n20923;
  assign n20925 = ~n20260 & ~n20267;
  assign n20926 = n20266 & n20925;
  assign n20927 = po2  & n20926;
  assign n20928 = po2  & n20925;
  assign n20929 = ~n20266 & ~n20928;
  assign n20930 = ~n20927 & ~n20929;
  assign n20931 = ~po62  & ~n20920;
  assign n20932 = ~n20922 & n20931;
  assign n20933 = ~n20930 & ~n20932;
  assign n20934 = ~n20924 & ~n20933;
  assign n20935 = ~n20270 & ~n20272;
  assign n20936 = po2  & n20935;
  assign n20937 = ~n20278 & ~n20936;
  assign n20938 = n20278 & n20936;
  assign n20939 = ~n20937 & ~n20938;
  assign n20940 = ~n20280 & ~n20285;
  assign n20941 = po2  & n20940;
  assign n20942 = ~n20296 & ~n20941;
  assign n20943 = ~n20939 & n20942;
  assign n20944 = ~n20934 & n20943;
  assign n20945 = ~po63  & ~n20944;
  assign n20946 = ~n20285 & po2 ;
  assign n20947 = n20280 & ~n20946;
  assign n20948 = po63  & ~n20940;
  assign n20949 = ~n20947 & n20948;
  assign n20950 = n20934 & n20939;
  assign n20951 = ~n20949 & ~n20950;
  assign po1  = n20945 | ~n20951;
  assign n20953 = ~n20920 & ~n20921;
  assign n20954 = po1  & n20953;
  assign n20955 = ~n20304 & ~n20954;
  assign n20956 = n20304 & n20953;
  assign n20957 = po1  & n20956;
  assign n20958 = ~n20955 & ~n20957;
  assign n20959 = ~n20909 & ~n20917;
  assign n20960 = po1  & n20959;
  assign n20961 = ~n20915 & ~n20960;
  assign n20962 = n20915 & n20959;
  assign n20963 = po1  & n20962;
  assign n20964 = ~n20961 & ~n20963;
  assign n20965 = ~n20899 & ~n20906;
  assign n20966 = po1  & n20965;
  assign n20967 = ~n20905 & ~n20966;
  assign n20968 = n20905 & n20965;
  assign n20969 = po1  & n20968;
  assign n20970 = ~n20967 & ~n20969;
  assign n20971 = ~n20888 & ~n20896;
  assign n20972 = po1  & n20971;
  assign n20973 = ~n20894 & ~n20972;
  assign n20974 = n20894 & n20971;
  assign n20975 = po1  & n20974;
  assign n20976 = ~n20973 & ~n20975;
  assign n20977 = ~n20878 & ~n20885;
  assign n20978 = po1  & n20977;
  assign n20979 = ~n20884 & ~n20978;
  assign n20980 = n20884 & n20977;
  assign n20981 = po1  & n20980;
  assign n20982 = ~n20979 & ~n20981;
  assign n20983 = ~n20867 & ~n20875;
  assign n20984 = po1  & n20983;
  assign n20985 = ~n20873 & ~n20984;
  assign n20986 = n20873 & n20983;
  assign n20987 = po1  & n20986;
  assign n20988 = ~n20985 & ~n20987;
  assign n20989 = ~n20857 & ~n20864;
  assign n20990 = po1  & n20989;
  assign n20991 = ~n20863 & ~n20990;
  assign n20992 = n20863 & n20989;
  assign n20993 = po1  & n20992;
  assign n20994 = ~n20991 & ~n20993;
  assign n20995 = ~n20846 & ~n20854;
  assign n20996 = po1  & n20995;
  assign n20997 = ~n20852 & ~n20996;
  assign n20998 = n20852 & n20995;
  assign n20999 = po1  & n20998;
  assign n21000 = ~n20997 & ~n20999;
  assign n21001 = ~n20836 & ~n20843;
  assign n21002 = po1  & n21001;
  assign n21003 = ~n20842 & ~n21002;
  assign n21004 = n20842 & n21001;
  assign n21005 = po1  & n21004;
  assign n21006 = ~n21003 & ~n21005;
  assign n21007 = ~n20825 & ~n20833;
  assign n21008 = po1  & n21007;
  assign n21009 = ~n20831 & ~n21008;
  assign n21010 = n20831 & n21007;
  assign n21011 = po1  & n21010;
  assign n21012 = ~n21009 & ~n21011;
  assign n21013 = ~n20815 & ~n20822;
  assign n21014 = po1  & n21013;
  assign n21015 = ~n20821 & ~n21014;
  assign n21016 = n20821 & n21013;
  assign n21017 = po1  & n21016;
  assign n21018 = ~n21015 & ~n21017;
  assign n21019 = ~n20804 & ~n20812;
  assign n21020 = po1  & n21019;
  assign n21021 = ~n20810 & ~n21020;
  assign n21022 = n20810 & n21019;
  assign n21023 = po1  & n21022;
  assign n21024 = ~n21021 & ~n21023;
  assign n21025 = ~n20794 & ~n20801;
  assign n21026 = po1  & n21025;
  assign n21027 = ~n20800 & ~n21026;
  assign n21028 = n20800 & n21025;
  assign n21029 = po1  & n21028;
  assign n21030 = ~n21027 & ~n21029;
  assign n21031 = ~n20783 & ~n20791;
  assign n21032 = po1  & n21031;
  assign n21033 = ~n20789 & ~n21032;
  assign n21034 = n20789 & n21031;
  assign n21035 = po1  & n21034;
  assign n21036 = ~n21033 & ~n21035;
  assign n21037 = ~n20773 & ~n20780;
  assign n21038 = po1  & n21037;
  assign n21039 = ~n20779 & ~n21038;
  assign n21040 = n20779 & n21037;
  assign n21041 = po1  & n21040;
  assign n21042 = ~n21039 & ~n21041;
  assign n21043 = ~n20762 & ~n20770;
  assign n21044 = po1  & n21043;
  assign n21045 = ~n20768 & ~n21044;
  assign n21046 = n20768 & n21043;
  assign n21047 = po1  & n21046;
  assign n21048 = ~n21045 & ~n21047;
  assign n21049 = ~n20752 & ~n20759;
  assign n21050 = po1  & n21049;
  assign n21051 = ~n20758 & ~n21050;
  assign n21052 = n20758 & n21049;
  assign n21053 = po1  & n21052;
  assign n21054 = ~n21051 & ~n21053;
  assign n21055 = ~n20741 & ~n20749;
  assign n21056 = po1  & n21055;
  assign n21057 = ~n20747 & ~n21056;
  assign n21058 = n20747 & n21055;
  assign n21059 = po1  & n21058;
  assign n21060 = ~n21057 & ~n21059;
  assign n21061 = ~n20731 & ~n20738;
  assign n21062 = po1  & n21061;
  assign n21063 = ~n20737 & ~n21062;
  assign n21064 = n20737 & n21061;
  assign n21065 = po1  & n21064;
  assign n21066 = ~n21063 & ~n21065;
  assign n21067 = ~n20720 & ~n20728;
  assign n21068 = po1  & n21067;
  assign n21069 = ~n20726 & ~n21068;
  assign n21070 = n20726 & n21067;
  assign n21071 = po1  & n21070;
  assign n21072 = ~n21069 & ~n21071;
  assign n21073 = ~n20710 & ~n20717;
  assign n21074 = po1  & n21073;
  assign n21075 = ~n20716 & ~n21074;
  assign n21076 = n20716 & n21073;
  assign n21077 = po1  & n21076;
  assign n21078 = ~n21075 & ~n21077;
  assign n21079 = ~n20699 & ~n20707;
  assign n21080 = po1  & n21079;
  assign n21081 = ~n20705 & ~n21080;
  assign n21082 = n20705 & n21079;
  assign n21083 = po1  & n21082;
  assign n21084 = ~n21081 & ~n21083;
  assign n21085 = ~n20689 & ~n20696;
  assign n21086 = po1  & n21085;
  assign n21087 = ~n20695 & ~n21086;
  assign n21088 = n20695 & n21085;
  assign n21089 = po1  & n21088;
  assign n21090 = ~n21087 & ~n21089;
  assign n21091 = ~n20678 & ~n20686;
  assign n21092 = po1  & n21091;
  assign n21093 = ~n20684 & ~n21092;
  assign n21094 = n20684 & n21091;
  assign n21095 = po1  & n21094;
  assign n21096 = ~n21093 & ~n21095;
  assign n21097 = ~n20668 & ~n20675;
  assign n21098 = po1  & n21097;
  assign n21099 = ~n20674 & ~n21098;
  assign n21100 = n20674 & n21097;
  assign n21101 = po1  & n21100;
  assign n21102 = ~n21099 & ~n21101;
  assign n21103 = ~n20657 & ~n20665;
  assign n21104 = po1  & n21103;
  assign n21105 = ~n20663 & ~n21104;
  assign n21106 = n20663 & n21103;
  assign n21107 = po1  & n21106;
  assign n21108 = ~n21105 & ~n21107;
  assign n21109 = ~n20647 & ~n20654;
  assign n21110 = po1  & n21109;
  assign n21111 = ~n20653 & ~n21110;
  assign n21112 = n20653 & n21109;
  assign n21113 = po1  & n21112;
  assign n21114 = ~n21111 & ~n21113;
  assign n21115 = ~n20636 & ~n20644;
  assign n21116 = po1  & n21115;
  assign n21117 = ~n20642 & ~n21116;
  assign n21118 = n20642 & n21115;
  assign n21119 = po1  & n21118;
  assign n21120 = ~n21117 & ~n21119;
  assign n21121 = ~n20626 & ~n20633;
  assign n21122 = po1  & n21121;
  assign n21123 = ~n20632 & ~n21122;
  assign n21124 = n20632 & n21121;
  assign n21125 = po1  & n21124;
  assign n21126 = ~n21123 & ~n21125;
  assign n21127 = ~n20615 & ~n20623;
  assign n21128 = po1  & n21127;
  assign n21129 = ~n20621 & ~n21128;
  assign n21130 = n20621 & n21127;
  assign n21131 = po1  & n21130;
  assign n21132 = ~n21129 & ~n21131;
  assign n21133 = ~n20605 & ~n20612;
  assign n21134 = po1  & n21133;
  assign n21135 = ~n20611 & ~n21134;
  assign n21136 = n20611 & n21133;
  assign n21137 = po1  & n21136;
  assign n21138 = ~n21135 & ~n21137;
  assign n21139 = ~n20594 & ~n20602;
  assign n21140 = po1  & n21139;
  assign n21141 = ~n20600 & ~n21140;
  assign n21142 = n20600 & n21139;
  assign n21143 = po1  & n21142;
  assign n21144 = ~n21141 & ~n21143;
  assign n21145 = ~n20584 & ~n20591;
  assign n21146 = po1  & n21145;
  assign n21147 = ~n20590 & ~n21146;
  assign n21148 = n20590 & n21145;
  assign n21149 = po1  & n21148;
  assign n21150 = ~n21147 & ~n21149;
  assign n21151 = ~n20573 & ~n20581;
  assign n21152 = po1  & n21151;
  assign n21153 = ~n20579 & ~n21152;
  assign n21154 = n20579 & n21151;
  assign n21155 = po1  & n21154;
  assign n21156 = ~n21153 & ~n21155;
  assign n21157 = ~n20563 & ~n20570;
  assign n21158 = po1  & n21157;
  assign n21159 = ~n20569 & ~n21158;
  assign n21160 = n20569 & n21157;
  assign n21161 = po1  & n21160;
  assign n21162 = ~n21159 & ~n21161;
  assign n21163 = ~n20552 & ~n20560;
  assign n21164 = po1  & n21163;
  assign n21165 = ~n20558 & ~n21164;
  assign n21166 = n20558 & n21163;
  assign n21167 = po1  & n21166;
  assign n21168 = ~n21165 & ~n21167;
  assign n21169 = ~n20542 & ~n20549;
  assign n21170 = po1  & n21169;
  assign n21171 = ~n20548 & ~n21170;
  assign n21172 = n20548 & n21169;
  assign n21173 = po1  & n21172;
  assign n21174 = ~n21171 & ~n21173;
  assign n21175 = ~n20531 & ~n20539;
  assign n21176 = po1  & n21175;
  assign n21177 = ~n20537 & ~n21176;
  assign n21178 = n20537 & n21175;
  assign n21179 = po1  & n21178;
  assign n21180 = ~n21177 & ~n21179;
  assign n21181 = ~n20521 & ~n20528;
  assign n21182 = po1  & n21181;
  assign n21183 = ~n20527 & ~n21182;
  assign n21184 = n20527 & n21181;
  assign n21185 = po1  & n21184;
  assign n21186 = ~n21183 & ~n21185;
  assign n21187 = ~n20510 & ~n20518;
  assign n21188 = po1  & n21187;
  assign n21189 = ~n20516 & ~n21188;
  assign n21190 = n20516 & n21187;
  assign n21191 = po1  & n21190;
  assign n21192 = ~n21189 & ~n21191;
  assign n21193 = ~n20500 & ~n20507;
  assign n21194 = po1  & n21193;
  assign n21195 = ~n20506 & ~n21194;
  assign n21196 = n20506 & n21193;
  assign n21197 = po1  & n21196;
  assign n21198 = ~n21195 & ~n21197;
  assign n21199 = ~n20489 & ~n20497;
  assign n21200 = po1  & n21199;
  assign n21201 = ~n20495 & ~n21200;
  assign n21202 = n20495 & n21199;
  assign n21203 = po1  & n21202;
  assign n21204 = ~n21201 & ~n21203;
  assign n21205 = ~n20479 & ~n20486;
  assign n21206 = po1  & n21205;
  assign n21207 = ~n20485 & ~n21206;
  assign n21208 = n20485 & n21205;
  assign n21209 = po1  & n21208;
  assign n21210 = ~n21207 & ~n21209;
  assign n21211 = ~n20468 & ~n20476;
  assign n21212 = po1  & n21211;
  assign n21213 = ~n20474 & ~n21212;
  assign n21214 = n20474 & n21211;
  assign n21215 = po1  & n21214;
  assign n21216 = ~n21213 & ~n21215;
  assign n21217 = ~n20458 & ~n20465;
  assign n21218 = po1  & n21217;
  assign n21219 = ~n20464 & ~n21218;
  assign n21220 = n20464 & n21217;
  assign n21221 = po1  & n21220;
  assign n21222 = ~n21219 & ~n21221;
  assign n21223 = ~n20447 & ~n20455;
  assign n21224 = po1  & n21223;
  assign n21225 = ~n20453 & ~n21224;
  assign n21226 = n20453 & n21223;
  assign n21227 = po1  & n21226;
  assign n21228 = ~n21225 & ~n21227;
  assign n21229 = ~n20437 & ~n20444;
  assign n21230 = po1  & n21229;
  assign n21231 = ~n20443 & ~n21230;
  assign n21232 = n20443 & n21229;
  assign n21233 = po1  & n21232;
  assign n21234 = ~n21231 & ~n21233;
  assign n21235 = ~n20426 & ~n20434;
  assign n21236 = po1  & n21235;
  assign n21237 = ~n20432 & ~n21236;
  assign n21238 = n20432 & n21235;
  assign n21239 = po1  & n21238;
  assign n21240 = ~n21237 & ~n21239;
  assign n21241 = ~n20416 & ~n20423;
  assign n21242 = po1  & n21241;
  assign n21243 = ~n20422 & ~n21242;
  assign n21244 = n20422 & n21241;
  assign n21245 = po1  & n21244;
  assign n21246 = ~n21243 & ~n21245;
  assign n21247 = ~n20405 & ~n20413;
  assign n21248 = po1  & n21247;
  assign n21249 = ~n20411 & ~n21248;
  assign n21250 = n20411 & n21247;
  assign n21251 = po1  & n21250;
  assign n21252 = ~n21249 & ~n21251;
  assign n21253 = ~n20395 & ~n20402;
  assign n21254 = po1  & n21253;
  assign n21255 = ~n20401 & ~n21254;
  assign n21256 = n20401 & n21253;
  assign n21257 = po1  & n21256;
  assign n21258 = ~n21255 & ~n21257;
  assign n21259 = ~n20384 & ~n20392;
  assign n21260 = po1  & n21259;
  assign n21261 = ~n20390 & ~n21260;
  assign n21262 = n20390 & n21259;
  assign n21263 = po1  & n21262;
  assign n21264 = ~n21261 & ~n21263;
  assign n21265 = ~n20374 & ~n20381;
  assign n21266 = po1  & n21265;
  assign n21267 = ~n20380 & ~n21266;
  assign n21268 = n20380 & n21265;
  assign n21269 = po1  & n21268;
  assign n21270 = ~n21267 & ~n21269;
  assign n21271 = ~n20363 & ~n20371;
  assign n21272 = po1  & n21271;
  assign n21273 = ~n20369 & ~n21272;
  assign n21274 = n20369 & n21271;
  assign n21275 = po1  & n21274;
  assign n21276 = ~n21273 & ~n21275;
  assign n21277 = ~n20353 & ~n20360;
  assign n21278 = po1  & n21277;
  assign n21279 = ~n20359 & ~n21278;
  assign n21280 = n20359 & n21277;
  assign n21281 = po1  & n21280;
  assign n21282 = ~n21279 & ~n21281;
  assign n21283 = ~n20342 & ~n20350;
  assign n21284 = po1  & n21283;
  assign n21285 = ~n20348 & ~n21284;
  assign n21286 = n20348 & n21283;
  assign n21287 = po1  & n21286;
  assign n21288 = ~n21285 & ~n21287;
  assign n21289 = ~n20332 & ~n20339;
  assign n21290 = n20338 & n21289;
  assign n21291 = po1  & n21290;
  assign n21292 = po1  & n21289;
  assign n21293 = ~n20338 & ~n21292;
  assign n21294 = ~n21291 & ~n21293;
  assign n21295 = ~n20320 & ~n20322;
  assign n21296 = po1  & n21295;
  assign n21297 = ~n20329 & ~n21296;
  assign n21298 = ~n20330 & n21295;
  assign n21299 = po1  & n21298;
  assign n21300 = ~n21297 & ~n21299;
  assign n21301 = ~n20309 & ~n20313;
  assign n21302 = ~n20317 & n21301;
  assign n21303 = po1  & n21302;
  assign n21304 = po1  & n21301;
  assign n21305 = n20317 & ~n21304;
  assign n21306 = ~n21303 & ~n21305;
  assign n21307 = n20306 & po1 ;
  assign n21308 = po2  & ~n20949;
  assign n21309 = ~n20950 & n21308;
  assign n21310 = ~n20945 & n21309;
  assign n21311 = ~n21307 & ~n21310;
  assign n21312 = pi4  & ~n21311;
  assign n21313 = ~pi4  & n21311;
  assign n21314 = ~n21312 & ~n21313;
  assign n21315 = ~pi2  & po1 ;
  assign n21316 = pi3  & ~n21315;
  assign n21317 = ~pi0  & ~pi1 ;
  assign n21318 = ~pi2  & ~n21317;
  assign n21319 = pi2  & ~n20949;
  assign n21320 = ~n20950 & n21319;
  assign n21321 = ~n20945 & n21320;
  assign n21322 = ~n21318 & ~n21321;
  assign n21323 = ~n21307 & n21322;
  assign n21324 = ~n21316 & n21323;
  assign n21325 = ~po2  & ~n21324;
  assign n21326 = ~n21307 & ~n21316;
  assign n21327 = ~n21322 & ~n21326;
  assign n21328 = ~n21325 & ~n21327;
  assign n21329 = ~n21314 & n21328;
  assign n21330 = ~po3  & ~n21329;
  assign n21331 = n21314 & ~n21328;
  assign n21332 = ~n21330 & ~n21331;
  assign n21333 = n21306 & ~n21332;
  assign n21334 = ~n21306 & ~n21331;
  assign n21335 = ~n21330 & n21334;
  assign n21336 = ~po4  & ~n21335;
  assign n21337 = ~n21333 & ~n21336;
  assign n21338 = ~n21300 & n21337;
  assign n21339 = ~po5  & ~n21338;
  assign n21340 = n21300 & ~n21337;
  assign n21341 = ~n21339 & ~n21340;
  assign n21342 = n21294 & ~n21341;
  assign n21343 = ~n21294 & ~n21340;
  assign n21344 = ~n21339 & n21343;
  assign n21345 = ~po6  & ~n21344;
  assign n21346 = ~n21342 & ~n21345;
  assign n21347 = ~n21288 & n21346;
  assign n21348 = ~po7  & ~n21347;
  assign n21349 = n21288 & ~n21346;
  assign n21350 = ~n21348 & ~n21349;
  assign n21351 = n21282 & ~n21350;
  assign n21352 = ~n21282 & ~n21349;
  assign n21353 = ~n21348 & n21352;
  assign n21354 = ~po8  & ~n21353;
  assign n21355 = ~n21351 & ~n21354;
  assign n21356 = ~n21276 & n21355;
  assign n21357 = ~po9  & ~n21356;
  assign n21358 = n21276 & ~n21355;
  assign n21359 = ~n21357 & ~n21358;
  assign n21360 = n21270 & ~n21359;
  assign n21361 = ~n21270 & ~n21358;
  assign n21362 = ~n21357 & n21361;
  assign n21363 = ~po10  & ~n21362;
  assign n21364 = ~n21360 & ~n21363;
  assign n21365 = ~n21264 & n21364;
  assign n21366 = ~po11  & ~n21365;
  assign n21367 = n21264 & ~n21364;
  assign n21368 = ~n21366 & ~n21367;
  assign n21369 = n21258 & ~n21368;
  assign n21370 = ~n21258 & ~n21367;
  assign n21371 = ~n21366 & n21370;
  assign n21372 = ~po12  & ~n21371;
  assign n21373 = ~n21369 & ~n21372;
  assign n21374 = ~n21252 & n21373;
  assign n21375 = ~po13  & ~n21374;
  assign n21376 = n21252 & ~n21373;
  assign n21377 = ~n21375 & ~n21376;
  assign n21378 = n21246 & ~n21377;
  assign n21379 = ~n21246 & ~n21376;
  assign n21380 = ~n21375 & n21379;
  assign n21381 = ~po14  & ~n21380;
  assign n21382 = ~n21378 & ~n21381;
  assign n21383 = ~n21240 & n21382;
  assign n21384 = ~po15  & ~n21383;
  assign n21385 = n21240 & ~n21382;
  assign n21386 = ~n21384 & ~n21385;
  assign n21387 = n21234 & ~n21386;
  assign n21388 = ~n21234 & ~n21385;
  assign n21389 = ~n21384 & n21388;
  assign n21390 = ~po16  & ~n21389;
  assign n21391 = ~n21387 & ~n21390;
  assign n21392 = ~n21228 & n21391;
  assign n21393 = ~po17  & ~n21392;
  assign n21394 = n21228 & ~n21391;
  assign n21395 = ~n21393 & ~n21394;
  assign n21396 = n21222 & ~n21395;
  assign n21397 = ~n21222 & ~n21394;
  assign n21398 = ~n21393 & n21397;
  assign n21399 = ~po18  & ~n21398;
  assign n21400 = ~n21396 & ~n21399;
  assign n21401 = ~n21216 & n21400;
  assign n21402 = ~po19  & ~n21401;
  assign n21403 = n21216 & ~n21400;
  assign n21404 = ~n21402 & ~n21403;
  assign n21405 = n21210 & ~n21404;
  assign n21406 = ~n21210 & ~n21403;
  assign n21407 = ~n21402 & n21406;
  assign n21408 = ~po20  & ~n21407;
  assign n21409 = ~n21405 & ~n21408;
  assign n21410 = ~n21204 & n21409;
  assign n21411 = ~po21  & ~n21410;
  assign n21412 = n21204 & ~n21409;
  assign n21413 = ~n21411 & ~n21412;
  assign n21414 = n21198 & ~n21413;
  assign n21415 = ~n21198 & ~n21412;
  assign n21416 = ~n21411 & n21415;
  assign n21417 = ~po22  & ~n21416;
  assign n21418 = ~n21414 & ~n21417;
  assign n21419 = ~n21192 & n21418;
  assign n21420 = ~po23  & ~n21419;
  assign n21421 = n21192 & ~n21418;
  assign n21422 = ~n21420 & ~n21421;
  assign n21423 = n21186 & ~n21422;
  assign n21424 = ~n21186 & ~n21421;
  assign n21425 = ~n21420 & n21424;
  assign n21426 = ~po24  & ~n21425;
  assign n21427 = ~n21423 & ~n21426;
  assign n21428 = ~n21180 & n21427;
  assign n21429 = ~po25  & ~n21428;
  assign n21430 = n21180 & ~n21427;
  assign n21431 = ~n21429 & ~n21430;
  assign n21432 = n21174 & ~n21431;
  assign n21433 = ~n21174 & ~n21430;
  assign n21434 = ~n21429 & n21433;
  assign n21435 = ~po26  & ~n21434;
  assign n21436 = ~n21432 & ~n21435;
  assign n21437 = ~n21168 & n21436;
  assign n21438 = ~po27  & ~n21437;
  assign n21439 = n21168 & ~n21436;
  assign n21440 = ~n21438 & ~n21439;
  assign n21441 = n21162 & ~n21440;
  assign n21442 = ~n21162 & ~n21439;
  assign n21443 = ~n21438 & n21442;
  assign n21444 = ~po28  & ~n21443;
  assign n21445 = ~n21441 & ~n21444;
  assign n21446 = ~n21156 & n21445;
  assign n21447 = ~po29  & ~n21446;
  assign n21448 = n21156 & ~n21445;
  assign n21449 = ~n21447 & ~n21448;
  assign n21450 = n21150 & ~n21449;
  assign n21451 = ~n21150 & ~n21448;
  assign n21452 = ~n21447 & n21451;
  assign n21453 = ~po30  & ~n21452;
  assign n21454 = ~n21450 & ~n21453;
  assign n21455 = ~n21144 & n21454;
  assign n21456 = ~po31  & ~n21455;
  assign n21457 = n21144 & ~n21454;
  assign n21458 = ~n21456 & ~n21457;
  assign n21459 = n21138 & ~n21458;
  assign n21460 = ~n21138 & ~n21457;
  assign n21461 = ~n21456 & n21460;
  assign n21462 = ~po32  & ~n21461;
  assign n21463 = ~n21459 & ~n21462;
  assign n21464 = ~n21132 & n21463;
  assign n21465 = ~po33  & ~n21464;
  assign n21466 = n21132 & ~n21463;
  assign n21467 = ~n21465 & ~n21466;
  assign n21468 = n21126 & ~n21467;
  assign n21469 = ~n21126 & ~n21466;
  assign n21470 = ~n21465 & n21469;
  assign n21471 = ~po34  & ~n21470;
  assign n21472 = ~n21468 & ~n21471;
  assign n21473 = ~n21120 & n21472;
  assign n21474 = ~po35  & ~n21473;
  assign n21475 = n21120 & ~n21472;
  assign n21476 = ~n21474 & ~n21475;
  assign n21477 = n21114 & ~n21476;
  assign n21478 = ~n21114 & ~n21475;
  assign n21479 = ~n21474 & n21478;
  assign n21480 = ~po36  & ~n21479;
  assign n21481 = ~n21477 & ~n21480;
  assign n21482 = ~n21108 & n21481;
  assign n21483 = ~po37  & ~n21482;
  assign n21484 = n21108 & ~n21481;
  assign n21485 = ~n21483 & ~n21484;
  assign n21486 = n21102 & ~n21485;
  assign n21487 = ~n21102 & ~n21484;
  assign n21488 = ~n21483 & n21487;
  assign n21489 = ~po38  & ~n21488;
  assign n21490 = ~n21486 & ~n21489;
  assign n21491 = ~n21096 & n21490;
  assign n21492 = ~po39  & ~n21491;
  assign n21493 = n21096 & ~n21490;
  assign n21494 = ~n21492 & ~n21493;
  assign n21495 = n21090 & ~n21494;
  assign n21496 = ~n21090 & ~n21493;
  assign n21497 = ~n21492 & n21496;
  assign n21498 = ~po40  & ~n21497;
  assign n21499 = ~n21495 & ~n21498;
  assign n21500 = ~n21084 & n21499;
  assign n21501 = ~po41  & ~n21500;
  assign n21502 = n21084 & ~n21499;
  assign n21503 = ~n21501 & ~n21502;
  assign n21504 = n21078 & ~n21503;
  assign n21505 = ~n21078 & ~n21502;
  assign n21506 = ~n21501 & n21505;
  assign n21507 = ~po42  & ~n21506;
  assign n21508 = ~n21504 & ~n21507;
  assign n21509 = ~n21072 & n21508;
  assign n21510 = ~po43  & ~n21509;
  assign n21511 = n21072 & ~n21508;
  assign n21512 = ~n21510 & ~n21511;
  assign n21513 = n21066 & ~n21512;
  assign n21514 = ~n21066 & ~n21511;
  assign n21515 = ~n21510 & n21514;
  assign n21516 = ~po44  & ~n21515;
  assign n21517 = ~n21513 & ~n21516;
  assign n21518 = ~n21060 & n21517;
  assign n21519 = ~po45  & ~n21518;
  assign n21520 = n21060 & ~n21517;
  assign n21521 = ~n21519 & ~n21520;
  assign n21522 = n21054 & ~n21521;
  assign n21523 = ~n21054 & ~n21520;
  assign n21524 = ~n21519 & n21523;
  assign n21525 = ~po46  & ~n21524;
  assign n21526 = ~n21522 & ~n21525;
  assign n21527 = ~n21048 & n21526;
  assign n21528 = ~po47  & ~n21527;
  assign n21529 = n21048 & ~n21526;
  assign n21530 = ~n21528 & ~n21529;
  assign n21531 = n21042 & ~n21530;
  assign n21532 = ~n21042 & ~n21529;
  assign n21533 = ~n21528 & n21532;
  assign n21534 = ~po48  & ~n21533;
  assign n21535 = ~n21531 & ~n21534;
  assign n21536 = ~n21036 & n21535;
  assign n21537 = ~po49  & ~n21536;
  assign n21538 = n21036 & ~n21535;
  assign n21539 = ~n21537 & ~n21538;
  assign n21540 = n21030 & ~n21539;
  assign n21541 = ~n21030 & ~n21538;
  assign n21542 = ~n21537 & n21541;
  assign n21543 = ~po50  & ~n21542;
  assign n21544 = ~n21540 & ~n21543;
  assign n21545 = ~n21024 & n21544;
  assign n21546 = ~po51  & ~n21545;
  assign n21547 = n21024 & ~n21544;
  assign n21548 = ~n21546 & ~n21547;
  assign n21549 = n21018 & ~n21548;
  assign n21550 = ~n21018 & ~n21547;
  assign n21551 = ~n21546 & n21550;
  assign n21552 = ~po52  & ~n21551;
  assign n21553 = ~n21549 & ~n21552;
  assign n21554 = ~n21012 & n21553;
  assign n21555 = ~po53  & ~n21554;
  assign n21556 = n21012 & ~n21553;
  assign n21557 = ~n21555 & ~n21556;
  assign n21558 = n21006 & ~n21557;
  assign n21559 = ~n21006 & ~n21556;
  assign n21560 = ~n21555 & n21559;
  assign n21561 = ~po54  & ~n21560;
  assign n21562 = ~n21558 & ~n21561;
  assign n21563 = ~n21000 & n21562;
  assign n21564 = ~po55  & ~n21563;
  assign n21565 = n21000 & ~n21562;
  assign n21566 = ~n21564 & ~n21565;
  assign n21567 = n20994 & ~n21566;
  assign n21568 = ~n20994 & ~n21565;
  assign n21569 = ~n21564 & n21568;
  assign n21570 = ~po56  & ~n21569;
  assign n21571 = ~n21567 & ~n21570;
  assign n21572 = ~n20988 & n21571;
  assign n21573 = ~po57  & ~n21572;
  assign n21574 = n20988 & ~n21571;
  assign n21575 = ~n21573 & ~n21574;
  assign n21576 = n20982 & ~n21575;
  assign n21577 = ~n20982 & ~n21574;
  assign n21578 = ~n21573 & n21577;
  assign n21579 = ~po58  & ~n21578;
  assign n21580 = ~n21576 & ~n21579;
  assign n21581 = ~n20976 & n21580;
  assign n21582 = ~po59  & ~n21581;
  assign n21583 = n20976 & ~n21580;
  assign n21584 = ~n21582 & ~n21583;
  assign n21585 = n20970 & ~n21584;
  assign n21586 = ~n20970 & ~n21583;
  assign n21587 = ~n21582 & n21586;
  assign n21588 = ~po60  & ~n21587;
  assign n21589 = ~n21585 & ~n21588;
  assign n21590 = ~n20964 & n21589;
  assign n21591 = ~po61  & ~n21590;
  assign n21592 = n20964 & ~n21589;
  assign n21593 = ~n21591 & ~n21592;
  assign n21594 = n20958 & ~n21593;
  assign n21595 = ~n20958 & ~n21592;
  assign n21596 = ~n21591 & n21595;
  assign n21597 = ~po62  & ~n21596;
  assign n21598 = ~n21594 & ~n21597;
  assign n21599 = ~n20924 & ~n20932;
  assign n21600 = po1  & n21599;
  assign n21601 = ~n20930 & ~n21600;
  assign n21602 = n20930 & n21600;
  assign n21603 = ~n21601 & ~n21602;
  assign n21604 = ~n20934 & ~n20939;
  assign n21605 = po1  & n21604;
  assign n21606 = ~n20950 & ~n21605;
  assign n21607 = ~n21603 & n21606;
  assign n21608 = n21598 & n21607;
  assign n21609 = ~po63  & ~n21608;
  assign n21610 = ~n21598 & n21603;
  assign n21611 = ~n20939 & po1 ;
  assign n21612 = n20934 & ~n21611;
  assign n21613 = po63  & ~n21604;
  assign n21614 = ~n21612 & n21613;
  assign n21615 = ~n21610 & ~n21614;
  assign po0  = n21609 | ~n21615;
endmodule
