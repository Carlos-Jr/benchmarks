module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n208, n209, n210,
    n211, n212, n213, n214, n215, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n345,
    n346, n347;
  assign n92 = ~pi9  & ~pi10 ;
  assign n93 = pi11  & ~n92;
  assign n94 = ~pi12  & ~n93;
  assign n95 = ~pi13  & n94;
  assign n96 = pi14  & ~n95;
  assign n97 = pi15  & n96;
  assign n98 = ~pi16  & ~n97;
  assign n99 = pi17  & ~n98;
  assign n100 = ~pi18  & ~n99;
  assign n101 = pi19  & ~n100;
  assign n102 = pi20  & n101;
  assign n103 = ~pi21  & ~n102;
  assign n104 = ~pi22  & n103;
  assign n105 = pi23  & ~n104;
  assign n106 = pi24  & n105;
  assign n107 = pi25  & n106;
  assign n108 = ~pi26  & ~n107;
  assign n109 = pi27  & ~n108;
  assign n110 = pi28  & n109;
  assign n111 = ~pi29  & n110;
  assign n112 = pi29  & ~n110;
  assign n113 = ~n111 & ~n112;
  assign n114 = pi28  & ~n109;
  assign n115 = ~pi28  & n109;
  assign n116 = ~n114 & ~n115;
  assign n117 = ~pi27  & n108;
  assign n118 = ~n109 & ~n117;
  assign n119 = pi26  & n107;
  assign n120 = ~n108 & ~n119;
  assign n121 = pi25  & ~n106;
  assign n122 = ~pi25  & n106;
  assign n123 = ~n121 & ~n122;
  assign n124 = pi24  & ~n105;
  assign n125 = ~pi24  & n105;
  assign n126 = ~n124 & ~n125;
  assign n127 = ~pi23  & n104;
  assign n128 = ~n105 & ~n127;
  assign n129 = pi22  & ~n103;
  assign n130 = ~n104 & ~n129;
  assign n131 = pi21  & n102;
  assign n132 = ~n103 & ~n131;
  assign n133 = pi20  & ~n101;
  assign n134 = ~pi20  & n101;
  assign n135 = ~n133 & ~n134;
  assign n136 = ~pi19  & n100;
  assign n137 = ~n101 & ~n136;
  assign n138 = pi18  & n99;
  assign n139 = ~n100 & ~n138;
  assign n140 = ~pi17  & n98;
  assign n141 = ~n99 & ~n140;
  assign n142 = pi16  & n97;
  assign n143 = ~n98 & ~n142;
  assign n144 = pi15  & ~n96;
  assign n145 = ~pi15  & n96;
  assign n146 = ~n144 & ~n145;
  assign n147 = ~pi14  & n95;
  assign n148 = ~n96 & ~n147;
  assign n149 = pi13  & ~n94;
  assign n150 = ~n95 & ~n149;
  assign n151 = pi12  & n93;
  assign n152 = ~n94 & ~n151;
  assign n153 = ~pi11  & n92;
  assign n154 = ~n93 & ~n153;
  assign n155 = pi9  & pi10 ;
  assign n156 = ~n92 & ~n155;
  assign n157 = pi0  & pi1 ;
  assign n158 = pi2  & pi3 ;
  assign n159 = pi4  & pi5 ;
  assign n160 = pi6  & pi7 ;
  assign n161 = pi8  & ~pi9 ;
  assign n162 = n160 & n161;
  assign n163 = n158 & n159;
  assign n164 = n157 & n163;
  assign n165 = ~n156 & n162;
  assign n166 = n164 & n165;
  assign n167 = n154 & n166;
  assign n168 = ~n152 & n167;
  assign n169 = ~n150 & n168;
  assign n170 = n148 & n169;
  assign n171 = ~n146 & n170;
  assign n172 = ~n143 & n171;
  assign n173 = n141 & n172;
  assign n174 = ~n139 & n173;
  assign n175 = n137 & n174;
  assign n176 = ~n135 & n175;
  assign n177 = ~n132 & n176;
  assign n178 = ~n130 & n177;
  assign n179 = n128 & n178;
  assign n180 = ~n126 & n179;
  assign n181 = ~n123 & n180;
  assign n182 = ~n120 & n181;
  assign n183 = n118 & n182;
  assign n184 = ~n116 & n183;
  assign n185 = ~n113 & n184;
  assign n186 = pi29  & n110;
  assign n187 = ~n185 & ~n186;
  assign n188 = ~pi1  & ~pi2 ;
  assign n189 = ~pi3  & ~pi4 ;
  assign n190 = ~pi5  & ~pi6 ;
  assign n191 = ~pi7  & ~pi8 ;
  assign n192 = pi9  & n191;
  assign n193 = n189 & n190;
  assign n194 = n188 & n193;
  assign n195 = n156 & n192;
  assign n196 = n194 & n195;
  assign n197 = ~n154 & n196;
  assign n198 = n152 & n197;
  assign n199 = n150 & n198;
  assign n200 = ~n148 & n199;
  assign n201 = n146 & n200;
  assign n202 = n143 & n201;
  assign n203 = ~n141 & n202;
  assign n204 = n139 & n203;
  assign n205 = ~n137 & n204;
  assign n206 = n135 & n205;
  assign n207 = n132 & n206;
  assign n208 = n130 & n207;
  assign n209 = ~n128 & n208;
  assign n210 = n126 & n209;
  assign n211 = n123 & n210;
  assign n212 = n120 & n211;
  assign n213 = ~n118 & n212;
  assign n214 = n116 & n213;
  assign n215 = n186 & ~n214;
  assign po0  = n187 | n215;
  assign n217 = ~pi39  & ~pi40 ;
  assign n218 = pi41  & ~n217;
  assign n219 = ~pi42  & ~n218;
  assign n220 = ~pi43  & n219;
  assign n221 = pi44  & ~n220;
  assign n222 = pi45  & n221;
  assign n223 = ~pi46  & ~n222;
  assign n224 = pi47  & ~n223;
  assign n225 = ~pi48  & ~n224;
  assign n226 = pi49  & ~n225;
  assign n227 = pi50  & n226;
  assign n228 = ~pi51  & ~n227;
  assign n229 = ~pi52  & n228;
  assign n230 = pi53  & ~n229;
  assign n231 = pi54  & n230;
  assign n232 = pi55  & n231;
  assign n233 = ~pi56  & ~n232;
  assign n234 = pi57  & ~n233;
  assign n235 = pi58  & pi59 ;
  assign n236 = n234 & n235;
  assign n237 = pi58  & ~n234;
  assign n238 = ~pi58  & n234;
  assign n239 = ~n237 & ~n238;
  assign n240 = ~pi57  & n233;
  assign n241 = ~n234 & ~n240;
  assign n242 = pi56  & n232;
  assign n243 = ~n233 & ~n242;
  assign n244 = pi55  & ~n231;
  assign n245 = ~pi55  & n231;
  assign n246 = ~n244 & ~n245;
  assign n247 = pi54  & ~n230;
  assign n248 = ~pi54  & n230;
  assign n249 = ~n247 & ~n248;
  assign n250 = ~pi53  & n229;
  assign n251 = ~n230 & ~n250;
  assign n252 = pi52  & ~n228;
  assign n253 = ~n229 & ~n252;
  assign n254 = pi51  & n227;
  assign n255 = ~n228 & ~n254;
  assign n256 = pi50  & ~n226;
  assign n257 = ~pi50  & n226;
  assign n258 = ~n256 & ~n257;
  assign n259 = ~pi49  & n225;
  assign n260 = ~n226 & ~n259;
  assign n261 = pi48  & n224;
  assign n262 = ~n225 & ~n261;
  assign n263 = ~pi47  & n223;
  assign n264 = ~n224 & ~n263;
  assign n265 = pi46  & n222;
  assign n266 = ~n223 & ~n265;
  assign n267 = pi45  & ~n221;
  assign n268 = ~pi45  & n221;
  assign n269 = ~n267 & ~n268;
  assign n270 = ~pi44  & n220;
  assign n271 = ~n221 & ~n270;
  assign n272 = pi43  & ~n219;
  assign n273 = ~n220 & ~n272;
  assign n274 = pi42  & n218;
  assign n275 = ~n219 & ~n274;
  assign n276 = ~pi41  & n217;
  assign n277 = ~n218 & ~n276;
  assign n278 = pi39  & pi40 ;
  assign n279 = ~n217 & ~n278;
  assign n280 = ~pi31  & ~pi32 ;
  assign n281 = ~pi33  & ~pi34 ;
  assign n282 = ~pi35  & ~pi36 ;
  assign n283 = ~pi37  & ~pi38 ;
  assign n284 = pi39  & n283;
  assign n285 = n281 & n282;
  assign n286 = n280 & n285;
  assign n287 = n279 & n284;
  assign n288 = n286 & n287;
  assign n289 = ~n277 & n288;
  assign n290 = n275 & n289;
  assign n291 = n273 & n290;
  assign n292 = ~n271 & n291;
  assign n293 = n269 & n292;
  assign n294 = n266 & n293;
  assign n295 = ~n264 & n294;
  assign n296 = n262 & n295;
  assign n297 = ~n260 & n296;
  assign n298 = n258 & n297;
  assign n299 = n255 & n298;
  assign n300 = n253 & n299;
  assign n301 = ~n251 & n300;
  assign n302 = n249 & n301;
  assign n303 = n246 & n302;
  assign n304 = n243 & n303;
  assign n305 = ~n241 & n304;
  assign n306 = n239 & n305;
  assign n307 = n236 & ~n306;
  assign n308 = ~pi0  & ~pi30 ;
  assign n309 = n236 & ~n308;
  assign n310 = pi30  & pi31 ;
  assign n311 = pi32  & pi33 ;
  assign n312 = pi34  & pi35 ;
  assign n313 = pi36  & pi37 ;
  assign n314 = pi38  & ~pi39 ;
  assign n315 = pi59  & n314;
  assign n316 = n312 & n313;
  assign n317 = n310 & n311;
  assign n318 = n316 & n317;
  assign n319 = ~n279 & n315;
  assign n320 = n318 & n319;
  assign n321 = n277 & n320;
  assign n322 = ~n275 & n321;
  assign n323 = ~n273 & n322;
  assign n324 = n271 & n323;
  assign n325 = ~n269 & n324;
  assign n326 = ~n266 & n325;
  assign n327 = n264 & n326;
  assign n328 = ~n262 & n327;
  assign n329 = n260 & n328;
  assign n330 = ~n258 & n329;
  assign n331 = ~n255 & n330;
  assign n332 = ~n253 & n331;
  assign n333 = n251 & n332;
  assign n334 = ~n249 & n333;
  assign n335 = ~n246 & n334;
  assign n336 = ~n243 & n335;
  assign n337 = n241 & n336;
  assign n338 = ~n239 & n337;
  assign n339 = ~n309 & ~n338;
  assign n340 = ~n307 & n339;
  assign n341 = pi0  & ~n236;
  assign n342 = ~n187 & ~n341;
  assign n343 = ~n340 & n342;
  assign po1  = ~n215 & ~n343;
  assign n345 = pi0  & pi30 ;
  assign n346 = n236 & n345;
  assign n347 = ~n307 & ~n346;
  assign po2  = ~po0  & ~n347;
  assign po3  = 1'b0;
  assign po4  = 1'b0;
  assign po5  = 1'b0;
  assign po6  = 1'b0;
  assign po7  = 1'b0;
  assign po8  = 1'b0;
  assign po9  = 1'b0;
  assign po10  = 1'b0;
  assign po11  = 1'b0;
  assign po12  = 1'b0;
  assign po13  = 1'b0;
  assign po14  = 1'b0;
  assign po15  = 1'b0;
  assign po16  = 1'b0;
  assign po17  = 1'b0;
  assign po18  = 1'b0;
  assign po19  = 1'b0;
  assign po20  = 1'b0;
  assign po21  = 1'b0;
  assign po22  = 1'b0;
  assign po23  = 1'b0;
  assign po24  = 1'b0;
  assign po25  = 1'b0;
  assign po26  = 1'b0;
  assign po27  = 1'b0;
  assign po28  = 1'b0;
  assign po29  = 1'b0;
endmodule
