module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n329, n330, n331;
  assign n92 = ~pi9  & ~pi10 ;
  assign n93 = pi11  & ~n92;
  assign n94 = ~pi12  & ~n93;
  assign n95 = ~pi13  & n94;
  assign n96 = pi14  & ~n95;
  assign n97 = pi15  & n96;
  assign n98 = ~pi16  & ~n97;
  assign n99 = pi17  & ~n98;
  assign n100 = ~pi18  & ~n99;
  assign n101 = pi19  & ~n100;
  assign n102 = pi20  & n101;
  assign n103 = ~pi21  & ~n102;
  assign n104 = ~pi22  & n103;
  assign n105 = pi23  & ~n104;
  assign n106 = pi24  & n105;
  assign n107 = pi25  & n106;
  assign n108 = ~pi26  & ~n107;
  assign n109 = pi27  & ~n108;
  assign n110 = pi28  & n109;
  assign n111 = pi29  & n110;
  assign n112 = ~pi28  & ~n109;
  assign n113 = pi26  & n107;
  assign n114 = ~n108 & ~n113;
  assign n115 = pi25  & ~n106;
  assign n116 = ~pi25  & n106;
  assign n117 = ~n115 & ~n116;
  assign n118 = pi22  & ~n103;
  assign n119 = ~n104 & ~n118;
  assign n120 = pi21  & n102;
  assign n121 = ~n103 & ~n120;
  assign n122 = ~pi19  & n100;
  assign n123 = ~n101 & ~n122;
  assign n124 = pi18  & n99;
  assign n125 = ~n100 & ~n124;
  assign n126 = pi20  & ~n101;
  assign n127 = ~pi20  & n101;
  assign n128 = ~n126 & ~n127;
  assign n129 = ~pi17  & n98;
  assign n130 = ~n99 & ~n129;
  assign n131 = pi16  & n97;
  assign n132 = ~n98 & ~n131;
  assign n133 = ~pi11  & n92;
  assign n134 = ~n93 & ~n133;
  assign n135 = pi15  & ~n96;
  assign n136 = ~pi15  & n96;
  assign n137 = ~n135 & ~n136;
  assign n138 = ~pi14  & n95;
  assign n139 = ~n96 & ~n138;
  assign n140 = pi13  & ~n94;
  assign n141 = ~n95 & ~n140;
  assign n142 = pi12  & n93;
  assign n143 = ~n94 & ~n142;
  assign n144 = ~pi27  & n108;
  assign n145 = ~n109 & ~n144;
  assign n146 = pi24  & ~n105;
  assign n147 = ~pi24  & n105;
  assign n148 = ~n146 & ~n147;
  assign n149 = ~pi23  & n104;
  assign n150 = ~n105 & ~n149;
  assign n151 = pi0  & pi1 ;
  assign n152 = pi2  & pi3 ;
  assign n153 = pi4  & pi5 ;
  assign n154 = pi6  & pi7 ;
  assign n155 = pi8  & pi29 ;
  assign n156 = n154 & n155;
  assign n157 = n152 & n153;
  assign n158 = n92 & n151;
  assign n159 = n157 & n158;
  assign n160 = n156 & n159;
  assign n161 = n134 & n160;
  assign n162 = ~n143 & n161;
  assign n163 = ~n141 & n162;
  assign n164 = n139 & n163;
  assign n165 = ~n137 & n164;
  assign n166 = ~n132 & n165;
  assign n167 = n130 & n166;
  assign n168 = ~n125 & n167;
  assign n169 = n123 & n168;
  assign n170 = ~n128 & n169;
  assign n171 = ~n121 & n170;
  assign n172 = ~n119 & n171;
  assign n173 = n150 & n172;
  assign n174 = ~n148 & n173;
  assign n175 = ~n117 & n174;
  assign n176 = ~n114 & n175;
  assign n177 = ~n110 & ~n112;
  assign n178 = n145 & n177;
  assign n179 = n176 & n178;
  assign n180 = ~n111 & ~n179;
  assign n181 = ~pi1  & ~pi2 ;
  assign n182 = ~pi3  & ~pi4 ;
  assign n183 = ~pi5  & ~pi6 ;
  assign n184 = ~pi7  & ~pi8 ;
  assign n185 = pi9  & ~pi10 ;
  assign n186 = n184 & n185;
  assign n187 = n182 & n183;
  assign n188 = n181 & n187;
  assign n189 = n186 & n188;
  assign n190 = ~n134 & n189;
  assign n191 = n143 & n190;
  assign n192 = n141 & n191;
  assign n193 = ~n139 & n192;
  assign n194 = n137 & n193;
  assign n195 = n132 & n194;
  assign n196 = ~n130 & n195;
  assign n197 = n125 & n196;
  assign n198 = ~n123 & n197;
  assign n199 = n128 & n198;
  assign n200 = n121 & n199;
  assign n201 = n119 & n200;
  assign n202 = ~n150 & n201;
  assign n203 = n148 & n202;
  assign n204 = n117 & n203;
  assign n205 = n114 & n204;
  assign n206 = ~n145 & n205;
  assign n207 = n111 & ~n206;
  assign po0  = n180 | n207;
  assign n209 = ~pi39  & ~pi40 ;
  assign n210 = pi41  & ~n209;
  assign n211 = ~pi42  & ~n210;
  assign n212 = ~pi43  & n211;
  assign n213 = pi44  & ~n212;
  assign n214 = pi45  & n213;
  assign n215 = ~pi46  & ~n214;
  assign n216 = pi47  & ~n215;
  assign n217 = ~pi48  & ~n216;
  assign n218 = pi49  & ~n217;
  assign n219 = pi50  & n218;
  assign n220 = ~pi51  & ~n219;
  assign n221 = ~pi52  & n220;
  assign n222 = pi53  & ~n221;
  assign n223 = pi54  & n222;
  assign n224 = pi55  & ~n223;
  assign n225 = ~pi55  & n223;
  assign n226 = ~n224 & ~n225;
  assign n227 = pi52  & ~n220;
  assign n228 = ~n221 & ~n227;
  assign n229 = pi51  & n219;
  assign n230 = ~n220 & ~n229;
  assign n231 = ~pi49  & n217;
  assign n232 = ~n218 & ~n231;
  assign n233 = pi48  & n216;
  assign n234 = ~n217 & ~n233;
  assign n235 = pi50  & ~n218;
  assign n236 = ~pi50  & n218;
  assign n237 = ~n235 & ~n236;
  assign n238 = ~pi47  & n215;
  assign n239 = ~n216 & ~n238;
  assign n240 = pi46  & n214;
  assign n241 = ~n215 & ~n240;
  assign n242 = ~pi44  & n212;
  assign n243 = ~n213 & ~n242;
  assign n244 = ~pi41  & n209;
  assign n245 = ~n210 & ~n244;
  assign n246 = pi45  & ~n213;
  assign n247 = ~pi45  & n213;
  assign n248 = ~n246 & ~n247;
  assign n249 = pi43  & ~n211;
  assign n250 = ~n212 & ~n249;
  assign n251 = pi42  & n210;
  assign n252 = ~n211 & ~n251;
  assign n253 = pi55  & n223;
  assign n254 = ~pi56  & ~n253;
  assign n255 = pi56  & n253;
  assign n256 = ~n254 & ~n255;
  assign n257 = pi54  & ~n222;
  assign n258 = ~pi54  & n222;
  assign n259 = ~n257 & ~n258;
  assign n260 = ~pi53  & n221;
  assign n261 = ~n222 & ~n260;
  assign n262 = pi57  & ~n254;
  assign n263 = ~pi57  & n254;
  assign n264 = ~n262 & ~n263;
  assign n265 = pi30  & pi31 ;
  assign n266 = pi32  & pi33 ;
  assign n267 = pi34  & pi35 ;
  assign n268 = pi36  & pi37 ;
  assign n269 = pi38  & pi58 ;
  assign n270 = pi59  & n269;
  assign n271 = n267 & n268;
  assign n272 = n265 & n266;
  assign n273 = n209 & n272;
  assign n274 = n270 & n271;
  assign n275 = n273 & n274;
  assign n276 = n245 & n275;
  assign n277 = ~n252 & n276;
  assign n278 = ~n250 & n277;
  assign n279 = n243 & n278;
  assign n280 = ~n248 & n279;
  assign n281 = ~n241 & n280;
  assign n282 = n239 & n281;
  assign n283 = ~n234 & n282;
  assign n284 = n232 & n283;
  assign n285 = ~n237 & n284;
  assign n286 = ~n230 & n285;
  assign n287 = ~n228 & n286;
  assign n288 = n261 & n287;
  assign n289 = ~n259 & n288;
  assign n290 = ~n226 & n289;
  assign n291 = ~n256 & n290;
  assign n292 = n264 & n291;
  assign n293 = pi58  & pi59 ;
  assign n294 = n262 & n293;
  assign n295 = ~pi31  & ~pi32 ;
  assign n296 = ~pi33  & ~pi34 ;
  assign n297 = ~pi35  & ~pi36 ;
  assign n298 = ~pi37  & ~pi38 ;
  assign n299 = pi39  & ~pi40 ;
  assign n300 = n298 & n299;
  assign n301 = n296 & n297;
  assign n302 = n295 & n301;
  assign n303 = n300 & n302;
  assign n304 = ~n245 & n303;
  assign n305 = n252 & n304;
  assign n306 = n250 & n305;
  assign n307 = ~n243 & n306;
  assign n308 = n248 & n307;
  assign n309 = n241 & n308;
  assign n310 = ~n239 & n309;
  assign n311 = n234 & n310;
  assign n312 = ~n232 & n311;
  assign n313 = n237 & n312;
  assign n314 = n230 & n313;
  assign n315 = n228 & n314;
  assign n316 = ~n261 & n315;
  assign n317 = n259 & n316;
  assign n318 = n226 & n317;
  assign n319 = n256 & n318;
  assign n320 = ~n264 & n319;
  assign n321 = ~pi0  & ~pi30 ;
  assign n322 = n320 & n321;
  assign n323 = n294 & ~n322;
  assign n324 = ~n292 & ~n323;
  assign n325 = pi0  & ~n294;
  assign n326 = ~n180 & ~n325;
  assign n327 = ~n324 & n326;
  assign po1  = ~n207 & ~n327;
  assign n329 = pi0  & pi30 ;
  assign n330 = n320 & ~n329;
  assign n331 = n294 & ~n330;
  assign po2  = ~po0  & n331;
  assign po3  = 1'b0;
  assign po4  = 1'b0;
  assign po5  = 1'b0;
  assign po6  = 1'b0;
  assign po7  = 1'b0;
  assign po8  = 1'b0;
  assign po9  = 1'b0;
  assign po10  = 1'b0;
  assign po11  = 1'b0;
  assign po12  = 1'b0;
  assign po13  = 1'b0;
  assign po14  = 1'b0;
  assign po15  = 1'b0;
  assign po16  = 1'b0;
  assign po17  = 1'b0;
  assign po18  = 1'b0;
  assign po19  = 1'b0;
  assign po20  = 1'b0;
  assign po21  = 1'b0;
  assign po22  = 1'b0;
  assign po23  = 1'b0;
  assign po24  = 1'b0;
  assign po25  = 1'b0;
  assign po26  = 1'b0;
  assign po27  = 1'b0;
  assign po28  = 1'b0;
  assign po29  = 1'b0;
endmodule
