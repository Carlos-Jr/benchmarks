module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24 ;
  wire n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n100, n101, n102, n103,
    n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061,
    n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331,
    n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231,
    n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3296, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321,
    n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561,
    n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591,
    n3592, n3593, n3594, n3595, n3596, n3597,
    n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621,
    n3622, n3623, n3624, n3625, n3626, n3627,
    n3629, n3630, n3631, n3632, n3633, n3634,
    n3635, n3636, n3637, n3638, n3639, n3640,
    n3641, n3642, n3643, n3644, n3645, n3646,
    n3647, n3648, n3649, n3650, n3651, n3652,
    n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664,
    n3665, n3666, n3667, n3668, n3669, n3670,
    n3671, n3672, n3673, n3674, n3675, n3676,
    n3677, n3678, n3679, n3680, n3681, n3682,
    n3683, n3684, n3685, n3686, n3687, n3688,
    n3689, n3690, n3691, n3692, n3693, n3694,
    n3695, n3696, n3697, n3698, n3699, n3700,
    n3701, n3702, n3703, n3704, n3705, n3706,
    n3707, n3708, n3709, n3710, n3711, n3712,
    n3713, n3714, n3715, n3716, n3717, n3718,
    n3719, n3720, n3721, n3722, n3723, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730,
    n3731, n3732, n3733, n3734, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742,
    n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3770, n3771, n3772, n3773,
    n3774, n3775, n3776, n3777, n3778, n3779,
    n3780, n3781, n3782, n3783, n3784, n3785,
    n3786, n3787, n3788, n3789, n3790, n3791,
    n3792, n3793, n3794, n3795, n3796, n3797,
    n3798, n3799, n3800, n3801, n3802, n3803,
    n3804, n3805, n3806, n3807, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815,
    n3816, n3817, n3818, n3819, n3820, n3821,
    n3822, n3823, n3824, n3825, n3826, n3827,
    n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3842, n3843, n3844, n3845,
    n3846, n3847, n3848, n3849, n3850, n3851,
    n3852, n3853, n3854, n3855, n3856, n3857,
    n3858, n3859, n3860, n3861, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881,
    n3882, n3883, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894,
    n3895, n3896, n3897, n3898, n3899, n3900,
    n3901, n3902, n3903, n3904, n3905, n3906,
    n3907, n3908, n3909, n3910, n3911, n3912,
    n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924,
    n3925, n3926, n3927, n3928, n3929, n3930,
    n3931, n3932, n3933, n3934, n3935, n3936,
    n3937, n3938, n3939, n3940, n3941, n3942,
    n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954,
    n3955, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966,
    n3967, n3968, n3969, n3970, n3971, n3972,
    n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990,
    n3991, n3992, n3993, n3995, n3996, n3997,
    n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027,
    n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057,
    n4058, n4059, n4060, n4061, n4062, n4063,
    n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4083, n4084, n4085, n4086, n4087,
    n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4095, n4096, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227,
    n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4249, n4250, n4251,
    n4252, n4253, n4254, n4255, n4256, n4257,
    n4258, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4303, n4304, n4305, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312,
    n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324,
    n4325, n4326, n4327, n4328, n4329, n4330,
    n4331, n4332, n4333, n4334, n4335, n4336,
    n4337, n4338, n4339, n4340, n4341, n4342,
    n4343, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354,
    n4355, n4356, n4357, n4358, n4359, n4360,
    n4361, n4362, n4363, n4364, n4365, n4366,
    n4367, n4368, n4369, n4370, n4371, n4372,
    n4373, n4374, n4375, n4376, n4377, n4378,
    n4379, n4380, n4381, n4382, n4383, n4384,
    n4385, n4386, n4387, n4388, n4389, n4390,
    n4391, n4392, n4394, n4395, n4396, n4397,
    n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415,
    n4416, n4417, n4418, n4419, n4420, n4421,
    n4422, n4423, n4424, n4425, n4426, n4427,
    n4428, n4429, n4430, n4431, n4432, n4433,
    n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445,
    n4446, n4447, n4448, n4449, n4450, n4451,
    n4452, n4453, n4454, n4455, n4456, n4457,
    n4458, n4459, n4460, n4461, n4462, n4463,
    n4464, n4465, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481,
    n4482, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560,
    n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682,
    n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700,
    n4702, n4703, n4704, n4705, n4706, n4707,
    n4708, n4709, n4710, n4711, n4712, n4713,
    n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737,
    n4738, n4739, n4740, n4741, n4742, n4743,
    n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761,
    n4762, n4764, n4765, n4766, n4767, n4768,
    n4769, n4770, n4771, n4772, n4773, n4774,
    n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786,
    n4787, n4788, n4789, n4790, n4791, n4792,
    n4793, n4794, n4795, n4796, n4797, n4798,
    n4799, n4800, n4801, n4802, n4803, n4804,
    n4805, n4806, n4807, n4808, n4809, n4810,
    n4811, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822,
    n4823, n4824, n4825, n4826, n4827, n4829,
    n4830, n4831, n4832, n4833, n4834, n4835,
    n4836, n4837, n4838, n4839, n4840, n4841,
    n4842, n4843, n4844, n4845, n4846, n4847,
    n4848, n4849, n4850, n4851, n4852, n4853,
    n4854, n4855, n4856, n4857, n4858, n4859,
    n4860, n4861, n4862, n4863, n4864, n4865,
    n4866, n4867, n4868, n4869, n4870, n4871,
    n4872, n4873, n4874, n4875, n4876, n4877,
    n4878, n4879, n4881, n4882, n4883, n4884,
    n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914,
    n4915, n4916, n4917, n4918, n4919, n4920,
    n4921, n4922, n4923, n4924, n4925, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963,
    n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4989,
    n4990, n4991, n4992, n4993, n4994, n4995,
    n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5003, n5004, n5005, n5006, n5007,
    n5009, n5010, n5011, n5012, n5013, n5014,
    n5015, n5016, n5017, n5018, n5019, n5020,
    n5021, n5022, n5023, n5024, n5025, n5026,
    n5027, n5028, n5029, n5030, n5031, n5033,
    n5034, n5035, n5036, n5037, n5038, n5039,
    n5040, n5041, n5042, n5043, n5044, n5045,
    n5046, n5047, n5048, n5050, n5051, n5052,
    n5053, n5054, n5055, n5056, n5057, n5058,
    n5059, n5060, n5061, n5062, n5063, n5064,
    n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5085,
    n5086, n5087, n5088, n5089;
  assign n50 = ~pi0  & ~pi1 ;
  assign n51 = ~pi2  & n50;
  assign n52 = ~pi3  & n51;
  assign n53 = ~pi4  & n52;
  assign n54 = ~pi22  & ~n53;
  assign n55 = ~pi5  & ~n54;
  assign n56 = pi5  & n54;
  assign n57 = ~n55 & ~n56;
  assign n58 = pi18  & pi22 ;
  assign n59 = ~pi5  & n53;
  assign n60 = ~pi6  & n59;
  assign n61 = ~pi7  & n60;
  assign n62 = ~pi8  & n61;
  assign n63 = ~pi9  & n62;
  assign n64 = ~pi10  & n63;
  assign n65 = ~pi11  & n64;
  assign n66 = ~pi12  & n65;
  assign n67 = ~pi13  & n66;
  assign n68 = ~pi14  & n67;
  assign n69 = ~pi15  & n68;
  assign n70 = ~pi16  & n69;
  assign n71 = ~pi17  & n70;
  assign n72 = ~pi18  & n71;
  assign n73 = ~pi22  & ~n72;
  assign n74 = pi18  & ~n71;
  assign n75 = n73 & ~n74;
  assign n76 = ~n58 & ~n75;
  assign n77 = ~pi19  & ~n73;
  assign n78 = pi19  & n73;
  assign n79 = ~n77 & ~n78;
  assign n80 = ~n76 & n79;
  assign n81 = ~pi22  & ~n70;
  assign n82 = pi17  & ~n81;
  assign n83 = ~pi17  & n81;
  assign n84 = ~n82 & ~n83;
  assign n85 = ~pi22  & ~n69;
  assign n86 = pi16  & ~n85;
  assign n87 = ~pi16  & n85;
  assign n88 = ~n86 & ~n87;
  assign n89 = ~n84 & ~n88;
  assign n90 = n80 & n89;
  assign n91 = ~pi22  & ~n68;
  assign n92 = pi15  & ~n91;
  assign n93 = ~pi15  & n91;
  assign n94 = ~n92 & ~n93;
  assign n95 = pi20  & pi22 ;
  assign n96 = ~pi19  & n72;
  assign n97 = pi20  & ~n96;
  assign n98 = ~pi20  & n96;
  assign n99 = ~pi22  & ~n98;
  assign n100 = ~n97 & n99;
  assign n101 = ~n95 & ~n100;
  assign n102 = pi21  & ~n99;
  assign n103 = ~pi21  & ~pi22 ;
  assign n104 = ~n98 & n103;
  assign n105 = ~n102 & ~n104;
  assign n106 = ~n101 & n105;
  assign n107 = ~n94 & n106;
  assign n108 = n90 & n107;
  assign n109 = n84 & ~n88;
  assign n110 = n80 & n109;
  assign n111 = n101 & n105;
  assign n112 = n94 & n111;
  assign n113 = n110 & n112;
  assign n114 = ~n108 & ~n113;
  assign n115 = ~n101 & ~n105;
  assign n116 = n94 & n115;
  assign n117 = n76 & ~n79;
  assign n118 = n89 & n117;
  assign n119 = n116 & n118;
  assign n120 = n101 & ~n105;
  assign n121 = n94 & n120;
  assign n122 = n84 & n88;
  assign n123 = n76 & n79;
  assign n124 = n122 & n123;
  assign n125 = n121 & n124;
  assign n126 = ~n84 & n88;
  assign n127 = n80 & n126;
  assign n128 = n94 & n106;
  assign n129 = n127 & n128;
  assign n130 = ~n76 & ~n79;
  assign n131 = n89 & n130;
  assign n132 = n112 & n131;
  assign n133 = n109 & n123;
  assign n134 = n112 & n133;
  assign n135 = n109 & n130;
  assign n136 = ~n94 & n111;
  assign n137 = n135 & n136;
  assign n138 = n122 & n130;
  assign n139 = n121 & n138;
  assign n140 = n136 & n138;
  assign n141 = ~n139 & ~n140;
  assign n142 = ~n137 & n141;
  assign n143 = n126 & n130;
  assign n144 = n136 & n143;
  assign n145 = n107 & n124;
  assign n146 = ~n144 & ~n145;
  assign n147 = n80 & n122;
  assign n148 = n121 & n147;
  assign n149 = n128 & n135;
  assign n150 = n123 & n126;
  assign n151 = n120 & n150;
  assign n152 = n94 & n151;
  assign n153 = n121 & n143;
  assign n154 = n116 & n131;
  assign n155 = ~n94 & n115;
  assign n156 = n124 & n155;
  assign n157 = ~n154 & ~n156;
  assign n158 = ~n148 & ~n149;
  assign n159 = ~n152 & ~n153;
  assign n160 = n158 & n159;
  assign n161 = n157 & n160;
  assign n162 = ~n119 & ~n125;
  assign n163 = ~n129 & ~n132;
  assign n164 = ~n134 & n163;
  assign n165 = n114 & n162;
  assign n166 = n146 & n165;
  assign n167 = n142 & n164;
  assign n168 = n166 & n167;
  assign n169 = n161 & n168;
  assign n170 = n110 & n120;
  assign n171 = ~n94 & n170;
  assign n172 = ~n94 & n120;
  assign n173 = n117 & n126;
  assign n174 = n172 & n173;
  assign n175 = n109 & n117;
  assign n176 = n121 & n175;
  assign n177 = ~n171 & ~n174;
  assign n178 = ~n176 & n177;
  assign n179 = n117 & n122;
  assign n180 = n107 & n179;
  assign n181 = n138 & n172;
  assign n182 = n135 & n172;
  assign n183 = ~n181 & ~n182;
  assign n184 = ~n180 & n183;
  assign n185 = n136 & n173;
  assign n186 = n112 & n127;
  assign n187 = ~n185 & ~n186;
  assign n188 = n136 & n175;
  assign n189 = n128 & n150;
  assign n190 = n133 & n172;
  assign n191 = n89 & n123;
  assign n192 = n172 & n191;
  assign n193 = ~n188 & ~n189;
  assign n194 = ~n190 & ~n192;
  assign n195 = n193 & n194;
  assign n196 = n107 & n175;
  assign n197 = n112 & n124;
  assign n198 = n128 & n143;
  assign n199 = n127 & n136;
  assign n200 = n116 & n124;
  assign n201 = n128 & n133;
  assign n202 = ~n196 & ~n197;
  assign n203 = ~n198 & ~n199;
  assign n204 = ~n200 & ~n201;
  assign n205 = n203 & n204;
  assign n206 = n202 & n205;
  assign n207 = n107 & n131;
  assign n208 = n116 & n133;
  assign n209 = n107 & n173;
  assign n210 = n107 & n147;
  assign n211 = ~n209 & ~n210;
  assign n212 = ~n207 & ~n208;
  assign n213 = n187 & n212;
  assign n214 = n211 & n213;
  assign n215 = n184 & n195;
  assign n216 = n214 & n215;
  assign n217 = n206 & n216;
  assign n218 = n116 & n179;
  assign n219 = n116 & n175;
  assign n220 = n136 & n179;
  assign n221 = ~n219 & ~n220;
  assign n222 = n118 & n155;
  assign n223 = n112 & n150;
  assign n224 = n128 & n138;
  assign n225 = n110 & n128;
  assign n226 = n112 & n147;
  assign n227 = ~n218 & ~n222;
  assign n228 = ~n223 & ~n224;
  assign n229 = ~n225 & ~n226;
  assign n230 = n228 & n229;
  assign n231 = n221 & n227;
  assign n232 = n230 & n231;
  assign n233 = n131 & n172;
  assign n234 = n90 & n111;
  assign n235 = ~n94 & n234;
  assign n236 = n106 & n191;
  assign n237 = ~n94 & n236;
  assign n238 = n118 & n128;
  assign n239 = n131 & n155;
  assign n240 = n112 & n191;
  assign n241 = ~n239 & ~n240;
  assign n242 = ~n233 & ~n235;
  assign n243 = ~n237 & ~n238;
  assign n244 = n242 & n243;
  assign n245 = n241 & n244;
  assign n246 = n120 & n127;
  assign n247 = n116 & n138;
  assign n248 = n118 & n136;
  assign n249 = n155 & n179;
  assign n250 = n138 & n155;
  assign n251 = n107 & n143;
  assign n252 = ~n249 & ~n250;
  assign n253 = ~n251 & n252;
  assign n254 = ~n246 & ~n247;
  assign n255 = ~n248 & n254;
  assign n256 = n178 & n255;
  assign n257 = n253 & n256;
  assign n258 = n232 & n245;
  assign n259 = n257 & n258;
  assign n260 = n169 & n259;
  assign n261 = n217 & n260;
  assign n262 = n116 & n173;
  assign n263 = n150 & n155;
  assign n264 = n121 & n173;
  assign n265 = ~n263 & ~n264;
  assign n266 = ~n262 & n265;
  assign n267 = n128 & n147;
  assign n268 = n110 & n155;
  assign n269 = ~n226 & ~n267;
  assign n270 = ~n268 & n269;
  assign n271 = n107 & n133;
  assign n272 = n133 & n136;
  assign n273 = n147 & n172;
  assign n274 = n90 & n128;
  assign n275 = ~n271 & ~n272;
  assign n276 = ~n273 & ~n274;
  assign n277 = n275 & n276;
  assign n278 = ~n152 & ~n238;
  assign n279 = n94 & n170;
  assign n280 = ~n94 & n246;
  assign n281 = ~n186 & ~n280;
  assign n282 = n133 & n155;
  assign n283 = n115 & n147;
  assign n284 = n94 & n283;
  assign n285 = ~n108 & ~n282;
  assign n286 = ~n284 & n285;
  assign n287 = ~n222 & ~n279;
  assign n288 = n278 & n287;
  assign n289 = n281 & n288;
  assign n290 = n266 & n270;
  assign n291 = n277 & n286;
  assign n292 = n290 & n291;
  assign n293 = n289 & n292;
  assign n294 = n128 & n173;
  assign n295 = n136 & n191;
  assign n296 = n121 & n133;
  assign n297 = ~n171 & ~n296;
  assign n298 = n110 & n136;
  assign n299 = n94 & n246;
  assign n300 = ~n225 & ~n299;
  assign n301 = ~n248 & ~n298;
  assign n302 = n300 & n301;
  assign n303 = n124 & n172;
  assign n304 = n110 & n116;
  assign n305 = ~n303 & ~n304;
  assign n306 = n90 & n155;
  assign n307 = n116 & n127;
  assign n308 = ~n119 & ~n307;
  assign n309 = n128 & n131;
  assign n310 = n112 & n135;
  assign n311 = n128 & n179;
  assign n312 = ~n199 & ~n311;
  assign n313 = n115 & n191;
  assign n314 = ~n94 & n313;
  assign n315 = n155 & n173;
  assign n316 = ~n250 & ~n315;
  assign n317 = n131 & n136;
  assign n318 = n121 & n135;
  assign n319 = ~n153 & ~n318;
  assign n320 = ~n314 & ~n317;
  assign n321 = n312 & n320;
  assign n322 = n316 & n319;
  assign n323 = n321 & n322;
  assign n324 = n127 & n155;
  assign n325 = n155 & n175;
  assign n326 = ~n324 & ~n325;
  assign n327 = n94 & n313;
  assign n328 = n326 & ~n327;
  assign n329 = n116 & n150;
  assign n330 = ~n189 & ~n207;
  assign n331 = ~n182 & ~n247;
  assign n332 = ~n309 & ~n310;
  assign n333 = ~n329 & n332;
  assign n334 = n308 & n331;
  assign n335 = n330 & n334;
  assign n336 = n328 & n333;
  assign n337 = n335 & n336;
  assign n338 = n323 & n337;
  assign n339 = ~n197 & ~n306;
  assign n340 = n338 & n339;
  assign n341 = n112 & n175;
  assign n342 = n112 & n118;
  assign n343 = n172 & n175;
  assign n344 = ~n342 & ~n343;
  assign n345 = n107 & n127;
  assign n346 = ~n149 & ~n345;
  assign n347 = ~n137 & ~n174;
  assign n348 = ~n223 & ~n341;
  assign n349 = n344 & n348;
  assign n350 = n346 & n347;
  assign n351 = n349 & n350;
  assign n352 = n211 & n351;
  assign n353 = ~n94 & n283;
  assign n354 = ~n190 & ~n353;
  assign n355 = n90 & n116;
  assign n356 = n107 & n138;
  assign n357 = ~n355 & ~n356;
  assign n358 = ~n180 & ~n188;
  assign n359 = ~n294 & ~n295;
  assign n360 = n358 & n359;
  assign n361 = n297 & n305;
  assign n362 = n354 & n357;
  assign n363 = n361 & n362;
  assign n364 = n302 & n360;
  assign n365 = n363 & n364;
  assign n366 = n352 & n365;
  assign n367 = n293 & n366;
  assign n368 = n340 & n367;
  assign n369 = ~n261 & ~n368;
  assign n370 = n112 & n173;
  assign n371 = ~n170 & ~n295;
  assign n372 = n107 & n118;
  assign n373 = ~n235 & ~n248;
  assign n374 = ~n372 & n373;
  assign n375 = ~n263 & ~n306;
  assign n376 = ~n314 & n375;
  assign n377 = n115 & n135;
  assign n378 = n112 & n143;
  assign n379 = ~n185 & ~n378;
  assign n380 = n94 & n234;
  assign n381 = n379 & ~n380;
  assign n382 = ~n377 & n381;
  assign n383 = ~n240 & ~n271;
  assign n384 = n121 & n191;
  assign n385 = ~n180 & ~n268;
  assign n386 = ~n139 & ~n284;
  assign n387 = ~n353 & ~n384;
  assign n388 = n383 & n387;
  assign n389 = n385 & n386;
  assign n390 = n388 & n389;
  assign n391 = ~n153 & ~n307;
  assign n392 = ~n370 & n391;
  assign n393 = n371 & n392;
  assign n394 = n374 & n376;
  assign n395 = n393 & n394;
  assign n396 = n382 & n390;
  assign n397 = n395 & n396;
  assign n398 = ~n182 & ~n189;
  assign n399 = ~n94 & n151;
  assign n400 = ~n197 & ~n299;
  assign n401 = ~n399 & n400;
  assign n402 = n398 & n401;
  assign n403 = n136 & n150;
  assign n404 = n124 & n128;
  assign n405 = ~n201 & ~n403;
  assign n406 = ~n404 & n405;
  assign n407 = n357 & n406;
  assign n408 = ~n327 & ~n329;
  assign n409 = ~n317 & ~n324;
  assign n410 = n346 & n408;
  assign n411 = n409 & n410;
  assign n412 = n116 & n143;
  assign n413 = ~n208 & ~n412;
  assign n414 = ~n129 & ~n304;
  assign n415 = ~n144 & ~n154;
  assign n416 = ~n239 & ~n280;
  assign n417 = ~n282 & n416;
  assign n418 = n413 & n415;
  assign n419 = n414 & n418;
  assign n420 = n417 & n419;
  assign n421 = n411 & n420;
  assign n422 = ~n156 & ~n224;
  assign n423 = n421 & n422;
  assign n424 = ~n145 & ~n274;
  assign n425 = ~n311 & n424;
  assign n426 = ~n273 & ~n342;
  assign n427 = n118 & n120;
  assign n428 = n94 & n427;
  assign n429 = n107 & n110;
  assign n430 = ~n148 & ~n318;
  assign n431 = ~n428 & ~n429;
  assign n432 = n430 & n431;
  assign n433 = n143 & n155;
  assign n434 = ~n181 & ~n192;
  assign n435 = ~n433 & n434;
  assign n436 = ~n94 & n427;
  assign n437 = ~n108 & ~n200;
  assign n438 = ~n226 & ~n436;
  assign n439 = n437 & n438;
  assign n440 = n435 & n439;
  assign n441 = ~n132 & n426;
  assign n442 = n425 & n441;
  assign n443 = n432 & n442;
  assign n444 = n402 & n407;
  assign n445 = n440 & n444;
  assign n446 = n443 & n445;
  assign n447 = n397 & n446;
  assign n448 = n423 & n447;
  assign n449 = ~n369 & ~n448;
  assign n450 = ~pi22  & ~n62;
  assign n451 = ~pi9  & ~n450;
  assign n452 = pi9  & n450;
  assign n453 = ~n451 & ~n452;
  assign n454 = ~n94 & n377;
  assign n455 = ~n233 & ~n454;
  assign n456 = ~n200 & ~n384;
  assign n457 = n143 & n172;
  assign n458 = n121 & n131;
  assign n459 = ~n457 & ~n458;
  assign n460 = ~n412 & n459;
  assign n461 = n94 & n377;
  assign n462 = ~n151 & ~n156;
  assign n463 = ~n192 & ~n208;
  assign n464 = ~n461 & n463;
  assign n465 = n455 & n462;
  assign n466 = n456 & n465;
  assign n467 = n460 & n464;
  assign n468 = n466 & n467;
  assign n469 = n90 & n121;
  assign n470 = ~n314 & ~n469;
  assign n471 = ~n246 & ~n283;
  assign n472 = n470 & n471;
  assign n473 = ~n154 & ~n247;
  assign n474 = ~n296 & ~n433;
  assign n475 = n473 & n474;
  assign n476 = ~n125 & ~n239;
  assign n477 = ~n303 & n476;
  assign n478 = ~n190 & ~n250;
  assign n479 = n475 & n478;
  assign n480 = n477 & n479;
  assign n481 = n90 & n172;
  assign n482 = ~n218 & ~n481;
  assign n483 = ~n119 & ~n273;
  assign n484 = ~n222 & ~n327;
  assign n485 = ~n171 & ~n263;
  assign n486 = ~n329 & n485;
  assign n487 = n483 & n484;
  assign n488 = n486 & n487;
  assign n489 = ~n148 & ~n279;
  assign n490 = n488 & n489;
  assign n491 = ~n249 & ~n268;
  assign n492 = ~n219 & ~n282;
  assign n493 = ~n304 & ~n307;
  assign n494 = n492 & n493;
  assign n495 = n482 & n491;
  assign n496 = n494 & n495;
  assign n497 = n480 & n496;
  assign n498 = n490 & n497;
  assign n499 = ~n90 & ~n173;
  assign n500 = n115 & ~n499;
  assign n501 = n326 & ~n500;
  assign n502 = n472 & n501;
  assign n503 = n468 & n502;
  assign n504 = n498 & n503;
  assign n505 = n453 & ~n504;
  assign n506 = ~n449 & n505;
  assign n507 = pi10  & pi22 ;
  assign n508 = ~pi22  & ~n64;
  assign n509 = pi10  & ~n63;
  assign n510 = n508 & ~n509;
  assign n511 = ~n507 & ~n510;
  assign n512 = ~n504 & ~n511;
  assign n513 = n449 & ~n505;
  assign n514 = ~n506 & ~n513;
  assign n515 = n512 & n514;
  assign n516 = ~n506 & ~n515;
  assign n517 = ~pi11  & ~n508;
  assign n518 = pi11  & n508;
  assign n519 = ~n517 & ~n518;
  assign n520 = n128 & n175;
  assign n521 = ~n356 & ~n520;
  assign n522 = ~n196 & ~n238;
  assign n523 = ~n294 & n522;
  assign n524 = n521 & n523;
  assign n525 = ~n209 & ~n224;
  assign n526 = ~n372 & n525;
  assign n527 = n524 & n526;
  assign n528 = ~n149 & n527;
  assign n529 = ~n271 & ~n404;
  assign n530 = n107 & n135;
  assign n531 = ~n198 & ~n309;
  assign n532 = ~n530 & n531;
  assign n533 = ~n145 & ~n201;
  assign n534 = ~n251 & n533;
  assign n535 = n330 & n529;
  assign n536 = n534 & n535;
  assign n537 = n532 & n536;
  assign n538 = ~n139 & ~n318;
  assign n539 = ~n210 & ~n429;
  assign n540 = ~n225 & n539;
  assign n541 = ~n236 & ~n345;
  assign n542 = n540 & n541;
  assign n543 = n107 & n150;
  assign n544 = ~n108 & ~n129;
  assign n545 = ~n176 & ~n428;
  assign n546 = ~n543 & n545;
  assign n547 = n544 & n546;
  assign n548 = n121 & n179;
  assign n549 = ~n153 & ~n274;
  assign n550 = ~n264 & ~n436;
  assign n551 = ~n174 & ~n343;
  assign n552 = n172 & n179;
  assign n553 = ~n267 & ~n552;
  assign n554 = ~n548 & n549;
  assign n555 = n550 & n551;
  assign n556 = n553 & n555;
  assign n557 = n554 & n556;
  assign n558 = n542 & n547;
  assign n559 = n557 & n558;
  assign n560 = n183 & n538;
  assign n561 = n537 & n560;
  assign n562 = n559 & n561;
  assign n563 = n528 & n562;
  assign n564 = n136 & n147;
  assign n565 = ~n298 & ~n564;
  assign n566 = ~n113 & ~n234;
  assign n567 = ~n186 & n566;
  assign n568 = n312 & n538;
  assign n569 = n565 & n568;
  assign n570 = n184 & n567;
  assign n571 = n569 & n570;
  assign n572 = ~n226 & ~n240;
  assign n573 = ~n295 & ~n403;
  assign n574 = n572 & n573;
  assign n575 = n571 & n574;
  assign n576 = n124 & n136;
  assign n577 = ~n134 & ~n576;
  assign n578 = ~n223 & ~n272;
  assign n579 = n577 & n578;
  assign n580 = n559 & n579;
  assign n581 = n575 & n580;
  assign n582 = n563 & n581;
  assign n583 = ~n563 & ~n581;
  assign n584 = ~n582 & ~n583;
  assign n585 = n504 & ~n563;
  assign n586 = ~n584 & ~n585;
  assign n587 = n519 & n586;
  assign n588 = ~n504 & ~n583;
  assign n589 = ~n584 & ~n588;
  assign n590 = ~n519 & n589;
  assign n591 = pi12  & pi22 ;
  assign n592 = ~pi22  & ~n66;
  assign n593 = pi12  & ~n65;
  assign n594 = n592 & ~n593;
  assign n595 = ~n591 & ~n594;
  assign n596 = ~n504 & ~n595;
  assign n597 = n504 & n595;
  assign n598 = ~n596 & ~n597;
  assign n599 = n584 & ~n598;
  assign n600 = ~n587 & ~n599;
  assign n601 = ~n590 & n600;
  assign n602 = pi14  & pi22 ;
  assign n603 = pi14  & ~n67;
  assign n604 = n91 & ~n603;
  assign n605 = ~n602 & ~n604;
  assign n606 = ~n176 & ~n481;
  assign n607 = ~n144 & ~n235;
  assign n608 = ~n304 & ~n454;
  assign n609 = n607 & n608;
  assign n610 = n606 & n609;
  assign n611 = n266 & n610;
  assign n612 = ~n222 & ~n343;
  assign n613 = n611 & n612;
  assign n614 = ~n218 & ~n469;
  assign n615 = ~n201 & ~n268;
  assign n616 = ~n174 & ~n251;
  assign n617 = ~n353 & ~n355;
  assign n618 = n616 & n617;
  assign n619 = n614 & n615;
  assign n620 = n618 & n619;
  assign n621 = ~n145 & ~n198;
  assign n622 = ~n140 & ~n186;
  assign n623 = ~n180 & ~n282;
  assign n624 = ~n378 & ~n433;
  assign n625 = n623 & n624;
  assign n626 = n413 & n621;
  assign n627 = n622 & n626;
  assign n628 = n625 & n627;
  assign n629 = ~n428 & ~n564;
  assign n630 = n112 & n138;
  assign n631 = ~n200 & ~n219;
  assign n632 = ~n404 & n631;
  assign n633 = ~n249 & ~n461;
  assign n634 = ~n239 & ~n271;
  assign n635 = n633 & n634;
  assign n636 = ~n137 & ~n181;
  assign n637 = ~n552 & ~n630;
  assign n638 = n636 & n637;
  assign n639 = n629 & n638;
  assign n640 = n632 & n635;
  assign n641 = n639 & n640;
  assign n642 = n628 & n641;
  assign n643 = n340 & n642;
  assign n644 = n157 & ~n298;
  assign n645 = ~n113 & ~n548;
  assign n646 = ~n436 & ~n530;
  assign n647 = ~n132 & ~n380;
  assign n648 = n386 & n647;
  assign n649 = n645 & n646;
  assign n650 = n648 & n649;
  assign n651 = n644 & n650;
  assign n652 = n620 & n651;
  assign n653 = n613 & n652;
  assign n654 = n643 & n653;
  assign n655 = n448 & n654;
  assign n656 = ~n448 & ~n654;
  assign n657 = ~n655 & ~n656;
  assign n658 = ~n581 & n657;
  assign n659 = ~n605 & n658;
  assign n660 = n581 & n657;
  assign n661 = n605 & n660;
  assign n662 = ~pi13  & ~n592;
  assign n663 = pi13  & n592;
  assign n664 = ~n662 & ~n663;
  assign n665 = ~n581 & ~n656;
  assign n666 = ~n657 & ~n665;
  assign n667 = ~n664 & n666;
  assign n668 = ~n448 & n581;
  assign n669 = ~n657 & ~n668;
  assign n670 = n664 & n669;
  assign n671 = ~n659 & ~n661;
  assign n672 = ~n667 & ~n670;
  assign n673 = n671 & n672;
  assign n674 = n601 & n673;
  assign n675 = n261 & n368;
  assign n676 = ~n369 & ~n675;
  assign n677 = ~n605 & ~n676;
  assign n678 = ~n449 & ~n677;
  assign n679 = ~n261 & n448;
  assign n680 = ~n676 & ~n679;
  assign n681 = ~n605 & n680;
  assign n682 = ~n678 & ~n681;
  assign n683 = ~n505 & n682;
  assign n684 = n505 & ~n682;
  assign n685 = ~n683 & ~n684;
  assign n686 = n658 & n664;
  assign n687 = n660 & ~n664;
  assign n688 = ~n595 & n669;
  assign n689 = n595 & n666;
  assign n690 = ~n686 & ~n687;
  assign n691 = ~n688 & ~n689;
  assign n692 = n690 & n691;
  assign n693 = n685 & n692;
  assign n694 = ~n683 & ~n693;
  assign n695 = ~n601 & ~n673;
  assign n696 = ~n674 & ~n695;
  assign n697 = ~n694 & n696;
  assign n698 = ~n674 & ~n697;
  assign n699 = ~n516 & ~n698;
  assign n700 = ~n504 & n519;
  assign n701 = ~n605 & ~n657;
  assign n702 = ~n665 & ~n701;
  assign n703 = ~n605 & n669;
  assign n704 = ~n702 & ~n703;
  assign n705 = ~n700 & n704;
  assign n706 = n700 & ~n704;
  assign n707 = ~n705 & ~n706;
  assign n708 = n586 & ~n595;
  assign n709 = n589 & n595;
  assign n710 = ~n504 & n664;
  assign n711 = n504 & ~n664;
  assign n712 = ~n710 & ~n711;
  assign n713 = n584 & ~n712;
  assign n714 = ~n708 & ~n713;
  assign n715 = ~n709 & n714;
  assign n716 = n707 & n715;
  assign n717 = ~n707 & ~n715;
  assign n718 = ~n716 & ~n717;
  assign n719 = n516 & n698;
  assign n720 = ~n699 & ~n719;
  assign n721 = n718 & n720;
  assign n722 = ~n699 & ~n721;
  assign n723 = ~n705 & ~n716;
  assign n724 = n586 & n664;
  assign n725 = n589 & ~n664;
  assign n726 = ~n504 & n605;
  assign n727 = n504 & ~n605;
  assign n728 = ~n726 & ~n727;
  assign n729 = n584 & n728;
  assign n730 = ~n724 & ~n729;
  assign n731 = ~n725 & n730;
  assign n732 = ~n723 & n731;
  assign n733 = n723 & ~n731;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~n665 & n700;
  assign n736 = n665 & ~n700;
  assign n737 = ~n735 & ~n736;
  assign n738 = n596 & n737;
  assign n739 = ~n596 & ~n737;
  assign n740 = ~n738 & ~n739;
  assign n741 = n734 & n740;
  assign n742 = ~n734 & ~n740;
  assign n743 = ~n741 & ~n742;
  assign n744 = ~n722 & n743;
  assign n745 = ~pi22  & ~n60;
  assign n746 = ~pi7  & ~n745;
  assign n747 = pi7  & n745;
  assign n748 = ~n746 & ~n747;
  assign n749 = ~n504 & n748;
  assign n750 = ~n264 & ~n274;
  assign n751 = n577 & n750;
  assign n752 = ~n208 & ~n458;
  assign n753 = ~n149 & ~n296;
  assign n754 = ~n189 & ~n263;
  assign n755 = ~n342 & ~n380;
  assign n756 = n754 & n755;
  assign n757 = n477 & n756;
  assign n758 = ~n222 & n615;
  assign n759 = n752 & n753;
  assign n760 = n758 & n759;
  assign n761 = n374 & n751;
  assign n762 = n760 & n761;
  assign n763 = n757 & n762;
  assign n764 = n112 & n179;
  assign n765 = ~n190 & ~n764;
  assign n766 = ~n174 & ~n370;
  assign n767 = ~n225 & ~n552;
  assign n768 = ~n132 & ~n185;
  assign n769 = ~n295 & n768;
  assign n770 = n414 & n767;
  assign n771 = n769 & n770;
  assign n772 = ~n226 & ~n384;
  assign n773 = ~n152 & n221;
  assign n774 = n772 & n773;
  assign n775 = ~n108 & ~n454;
  assign n776 = ~n307 & ~n315;
  assign n777 = ~n457 & n776;
  assign n778 = ~n233 & ~n469;
  assign n779 = ~n238 & ~n404;
  assign n780 = n775 & n778;
  assign n781 = n779 & n780;
  assign n782 = n777 & n781;
  assign n783 = ~n251 & ~n267;
  assign n784 = ~n196 & ~n207;
  assign n785 = ~n273 & ~n317;
  assign n786 = ~n327 & ~n355;
  assign n787 = n785 & n786;
  assign n788 = n783 & n784;
  assign n789 = n787 & n788;
  assign n790 = n771 & n789;
  assign n791 = n774 & n790;
  assign n792 = n782 & n791;
  assign n793 = n94 & n236;
  assign n794 = ~n306 & ~n793;
  assign n795 = ~n199 & n794;
  assign n796 = ~n197 & ~n250;
  assign n797 = ~n324 & n796;
  assign n798 = ~n139 & ~n148;
  assign n799 = ~n188 & ~n249;
  assign n800 = ~n280 & ~n399;
  assign n801 = ~n564 & n800;
  assign n802 = n798 & n799;
  assign n803 = n801 & n802;
  assign n804 = ~n341 & ~n481;
  assign n805 = n521 & n804;
  assign n806 = n765 & n766;
  assign n807 = n805 & n806;
  assign n808 = n435 & n795;
  assign n809 = n797 & n808;
  assign n810 = n803 & n807;
  assign n811 = n809 & n810;
  assign n812 = n763 & n811;
  assign n813 = n792 & n812;
  assign n814 = ~n251 & ~n793;
  assign n815 = ~n384 & n814;
  assign n816 = ~n181 & ~n240;
  assign n817 = n815 & n816;
  assign n818 = ~n224 & ~n309;
  assign n819 = ~n237 & ~n271;
  assign n820 = ~n436 & n819;
  assign n821 = ~n148 & ~n152;
  assign n822 = ~n324 & ~n372;
  assign n823 = n821 & n822;
  assign n824 = n818 & n823;
  assign n825 = n820 & n824;
  assign n826 = ~n200 & ~n353;
  assign n827 = ~n219 & ~n247;
  assign n828 = ~n156 & ~n279;
  assign n829 = ~n306 & n828;
  assign n830 = n827 & n829;
  assign n831 = ~n284 & ~n307;
  assign n832 = ~n355 & ~n429;
  assign n833 = n831 & n832;
  assign n834 = ~n262 & ~n272;
  assign n835 = ~n433 & n834;
  assign n836 = n300 & n385;
  assign n837 = n606 & n836;
  assign n838 = n751 & n835;
  assign n839 = n833 & n838;
  assign n840 = n830 & n837;
  assign n841 = n839 & n840;
  assign n842 = ~n132 & ~n197;
  assign n843 = n826 & n842;
  assign n844 = n841 & n843;
  assign n845 = ~n235 & ~n403;
  assign n846 = ~n125 & ~n280;
  assign n847 = ~n223 & n846;
  assign n848 = ~n458 & ~n552;
  assign n849 = ~n238 & ~n304;
  assign n850 = n845 & n849;
  assign n851 = n848 & n850;
  assign n852 = n847 & n851;
  assign n853 = ~n201 & ~n296;
  assign n854 = ~n380 & n853;
  assign n855 = n413 & n854;
  assign n856 = n323 & n855;
  assign n857 = n817 & n856;
  assign n858 = n825 & n852;
  assign n859 = n857 & n858;
  assign n860 = n844 & n859;
  assign n861 = ~n813 & ~n860;
  assign n862 = ~n261 & ~n861;
  assign n863 = n749 & ~n862;
  assign n864 = ~n749 & n862;
  assign n865 = ~n863 & ~n864;
  assign n866 = pi8  & pi22 ;
  assign n867 = pi8  & ~n61;
  assign n868 = n450 & ~n867;
  assign n869 = ~n866 & ~n868;
  assign n870 = ~n504 & ~n869;
  assign n871 = n865 & n870;
  assign n872 = ~n863 & ~n871;
  assign n873 = ~n511 & n586;
  assign n874 = n511 & n589;
  assign n875 = n504 & ~n519;
  assign n876 = ~n700 & ~n875;
  assign n877 = n584 & ~n876;
  assign n878 = ~n873 & ~n877;
  assign n879 = ~n874 & n878;
  assign n880 = ~n872 & n879;
  assign n881 = ~n448 & n676;
  assign n882 = ~n605 & n881;
  assign n883 = n448 & n676;
  assign n884 = n605 & n883;
  assign n885 = ~n449 & ~n676;
  assign n886 = ~n664 & n885;
  assign n887 = n664 & n680;
  assign n888 = ~n882 & ~n884;
  assign n889 = ~n886 & ~n887;
  assign n890 = n888 & n889;
  assign n891 = ~n595 & n658;
  assign n892 = n595 & n660;
  assign n893 = ~n519 & n666;
  assign n894 = n519 & n669;
  assign n895 = ~n891 & ~n892;
  assign n896 = ~n893 & ~n894;
  assign n897 = n895 & n896;
  assign n898 = n890 & n897;
  assign n899 = ~n890 & ~n897;
  assign n900 = ~n898 & ~n899;
  assign n901 = n453 & n586;
  assign n902 = ~n453 & n589;
  assign n903 = n504 & n511;
  assign n904 = ~n512 & ~n903;
  assign n905 = n584 & ~n904;
  assign n906 = ~n901 & ~n905;
  assign n907 = ~n902 & n906;
  assign n908 = n900 & n907;
  assign n909 = ~n898 & ~n908;
  assign n910 = n872 & ~n879;
  assign n911 = ~n880 & ~n910;
  assign n912 = ~n909 & n911;
  assign n913 = ~n880 & ~n912;
  assign n914 = ~n512 & ~n514;
  assign n915 = ~n515 & ~n914;
  assign n916 = ~n913 & n915;
  assign n917 = n913 & ~n915;
  assign n918 = ~n916 & ~n917;
  assign n919 = n694 & ~n696;
  assign n920 = ~n697 & ~n919;
  assign n921 = n918 & n920;
  assign n922 = ~n916 & ~n921;
  assign n923 = ~n718 & ~n720;
  assign n924 = ~n721 & ~n923;
  assign n925 = ~n922 & n924;
  assign n926 = n586 & ~n869;
  assign n927 = n589 & n869;
  assign n928 = ~n453 & n504;
  assign n929 = ~n505 & ~n928;
  assign n930 = n584 & ~n929;
  assign n931 = ~n926 & ~n930;
  assign n932 = ~n927 & n931;
  assign n933 = n519 & n658;
  assign n934 = ~n519 & n660;
  assign n935 = ~n511 & n669;
  assign n936 = n511 & n666;
  assign n937 = ~n933 & ~n934;
  assign n938 = ~n935 & ~n936;
  assign n939 = n937 & n938;
  assign n940 = n932 & n939;
  assign n941 = ~n932 & ~n939;
  assign n942 = ~n940 & ~n941;
  assign n943 = ~n303 & ~n315;
  assign n944 = ~n145 & ~n181;
  assign n945 = ~n210 & ~n239;
  assign n946 = ~n295 & ~n296;
  assign n947 = n945 & n946;
  assign n948 = n347 & n944;
  assign n949 = n386 & n783;
  assign n950 = n948 & n949;
  assign n951 = n947 & n950;
  assign n952 = ~n148 & ~n207;
  assign n953 = ~n220 & ~n294;
  assign n954 = ~n576 & n953;
  assign n955 = n491 & n952;
  assign n956 = n550 & n955;
  assign n957 = n954 & n956;
  assign n958 = ~n272 & ~n630;
  assign n959 = ~n356 & ~n543;
  assign n960 = ~n151 & ~n199;
  assign n961 = ~n236 & n959;
  assign n962 = n960 & n961;
  assign n963 = ~n250 & ~n412;
  assign n964 = ~n299 & ~n370;
  assign n965 = ~n552 & n964;
  assign n966 = ~n153 & ~n196;
  assign n967 = ~n520 & n966;
  assign n968 = ~n113 & ~n201;
  assign n969 = ~n353 & ~n428;
  assign n970 = n968 & n969;
  assign n971 = ~n108 & ~n355;
  assign n972 = ~n403 & ~n458;
  assign n973 = n971 & n972;
  assign n974 = n346 & n973;
  assign n975 = n965 & n967;
  assign n976 = n970 & n975;
  assign n977 = n830 & n974;
  assign n978 = n976 & n977;
  assign n979 = ~n119 & ~n132;
  assign n980 = ~n209 & ~n225;
  assign n981 = ~n280 & n980;
  assign n982 = n765 & n979;
  assign n983 = n943 & n958;
  assign n984 = n963 & n983;
  assign n985 = n981 & n982;
  assign n986 = n984 & n985;
  assign n987 = n382 & n962;
  assign n988 = n986 & n987;
  assign n989 = n951 & n957;
  assign n990 = n988 & n989;
  assign n991 = n978 & n990;
  assign n992 = n813 & n991;
  assign n993 = ~n132 & ~n296;
  assign n994 = ~n153 & ~n188;
  assign n995 = ~n249 & ~n325;
  assign n996 = n994 & n995;
  assign n997 = n614 & n772;
  assign n998 = n993 & n997;
  assign n999 = n996 & n998;
  assign n1000 = ~n303 & n847;
  assign n1001 = ~n140 & ~n192;
  assign n1002 = ~n220 & ~n317;
  assign n1003 = ~n341 & ~n764;
  assign n1004 = n1002 & n1003;
  assign n1005 = n183 & n1001;
  assign n1006 = n371 & n1005;
  assign n1007 = n1004 & n1006;
  assign n1008 = n1000 & n1007;
  assign n1009 = n999 & n1008;
  assign n1010 = ~n129 & ~n247;
  assign n1011 = ~n267 & ~n461;
  assign n1012 = n1010 & n1011;
  assign n1013 = ~n271 & ~n355;
  assign n1014 = ~n306 & ~n433;
  assign n1015 = n354 & n1014;
  assign n1016 = n551 & n958;
  assign n1017 = n1015 & n1016;
  assign n1018 = ~n238 & ~n307;
  assign n1019 = ~n310 & ~n329;
  assign n1020 = ~n548 & n1019;
  assign n1021 = n455 & n1018;
  assign n1022 = n1013 & n1021;
  assign n1023 = n644 & n1020;
  assign n1024 = n797 & n1023;
  assign n1025 = n962 & n1022;
  assign n1026 = n1017 & n1025;
  assign n1027 = n1024 & n1026;
  assign n1028 = ~n294 & ~n311;
  assign n1029 = n646 & n1028;
  assign n1030 = n818 & n1029;
  assign n1031 = n114 & ~n520;
  assign n1032 = n330 & n413;
  assign n1033 = n484 & n1032;
  assign n1034 = n540 & n1031;
  assign n1035 = n1012 & n1034;
  assign n1036 = n1030 & n1033;
  assign n1037 = n1035 & n1036;
  assign n1038 = n1009 & n1037;
  assign n1039 = n1027 & n1038;
  assign n1040 = ~n991 & ~n1039;
  assign n1041 = ~n813 & ~n1040;
  assign n1042 = ~n991 & n1041;
  assign n1043 = pi6  & pi22 ;
  assign n1044 = pi6  & ~n59;
  assign n1045 = n745 & ~n1044;
  assign n1046 = ~n1043 & ~n1045;
  assign n1047 = ~n504 & ~n1046;
  assign n1048 = ~n1042 & n1047;
  assign n1049 = ~n992 & ~n1048;
  assign n1050 = n942 & ~n1049;
  assign n1051 = ~n940 & ~n1050;
  assign n1052 = n813 & n860;
  assign n1053 = ~n861 & ~n1052;
  assign n1054 = ~n605 & ~n1053;
  assign n1055 = ~n862 & ~n1054;
  assign n1056 = n261 & ~n1052;
  assign n1057 = n1054 & ~n1056;
  assign n1058 = ~n1055 & ~n1057;
  assign n1059 = ~n749 & n1058;
  assign n1060 = n749 & ~n1058;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = n664 & n881;
  assign n1063 = ~n664 & n883;
  assign n1064 = ~n595 & n680;
  assign n1065 = n595 & n885;
  assign n1066 = ~n1062 & ~n1063;
  assign n1067 = ~n1064 & ~n1065;
  assign n1068 = n1066 & n1067;
  assign n1069 = n1061 & n1068;
  assign n1070 = ~n1059 & ~n1069;
  assign n1071 = ~n1051 & ~n1070;
  assign n1072 = ~n865 & ~n870;
  assign n1073 = ~n871 & ~n1072;
  assign n1074 = n1051 & n1070;
  assign n1075 = ~n1071 & ~n1074;
  assign n1076 = n1073 & n1075;
  assign n1077 = ~n1071 & ~n1076;
  assign n1078 = ~n685 & ~n692;
  assign n1079 = ~n693 & ~n1078;
  assign n1080 = ~n1077 & n1079;
  assign n1081 = n1077 & ~n1079;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = n909 & ~n911;
  assign n1084 = ~n912 & ~n1083;
  assign n1085 = n1082 & n1084;
  assign n1086 = ~n1080 & ~n1085;
  assign n1087 = ~n918 & ~n920;
  assign n1088 = ~n921 & ~n1087;
  assign n1089 = ~n1086 & n1088;
  assign n1090 = n586 & n748;
  assign n1091 = n589 & ~n748;
  assign n1092 = n504 & n869;
  assign n1093 = ~n870 & ~n1092;
  assign n1094 = n584 & ~n1093;
  assign n1095 = ~n1090 & ~n1094;
  assign n1096 = ~n1091 & n1095;
  assign n1097 = ~n511 & n658;
  assign n1098 = n511 & n660;
  assign n1099 = ~n453 & n666;
  assign n1100 = n453 & n669;
  assign n1101 = ~n1097 & ~n1098;
  assign n1102 = ~n1099 & ~n1100;
  assign n1103 = n1101 & n1102;
  assign n1104 = n1096 & n1103;
  assign n1105 = ~n1096 & ~n1103;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = ~n862 & ~n1053;
  assign n1108 = ~n664 & ~n1107;
  assign n1109 = ~n1053 & ~n1056;
  assign n1110 = n664 & ~n1109;
  assign n1111 = ~n1108 & ~n1110;
  assign n1112 = n862 & ~n1052;
  assign n1113 = ~n605 & n1112;
  assign n1114 = ~n861 & n1056;
  assign n1115 = n605 & n1114;
  assign n1116 = ~n1113 & ~n1115;
  assign n1117 = ~n1111 & n1116;
  assign n1118 = n1106 & n1117;
  assign n1119 = ~n1104 & ~n1118;
  assign n1120 = ~n1061 & ~n1068;
  assign n1121 = ~n1069 & ~n1120;
  assign n1122 = ~n1119 & n1121;
  assign n1123 = ~n942 & n1049;
  assign n1124 = ~n1050 & ~n1123;
  assign n1125 = n1119 & ~n1121;
  assign n1126 = ~n1122 & ~n1125;
  assign n1127 = n1124 & n1126;
  assign n1128 = ~n1122 & ~n1127;
  assign n1129 = ~n900 & ~n907;
  assign n1130 = ~n908 & ~n1129;
  assign n1131 = ~n1128 & n1130;
  assign n1132 = n1128 & ~n1130;
  assign n1133 = ~n1131 & ~n1132;
  assign n1134 = ~n1073 & ~n1075;
  assign n1135 = ~n1076 & ~n1134;
  assign n1136 = n1133 & n1135;
  assign n1137 = ~n1131 & ~n1136;
  assign n1138 = ~n1082 & ~n1084;
  assign n1139 = ~n1085 & ~n1138;
  assign n1140 = ~n1137 & n1139;
  assign n1141 = ~n992 & ~n1042;
  assign n1142 = n1047 & ~n1141;
  assign n1143 = ~n1048 & n1141;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = ~n595 & n881;
  assign n1146 = n595 & n883;
  assign n1147 = ~n519 & n885;
  assign n1148 = n519 & n680;
  assign n1149 = ~n1145 & ~n1146;
  assign n1150 = ~n1147 & ~n1148;
  assign n1151 = n1149 & n1150;
  assign n1152 = ~n1144 & n1151;
  assign n1153 = n57 & ~n504;
  assign n1154 = ~n991 & n1153;
  assign n1155 = n991 & ~n1153;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = n991 & n1039;
  assign n1158 = ~n1040 & ~n1157;
  assign n1159 = ~n605 & ~n1158;
  assign n1160 = ~n1041 & ~n1159;
  assign n1161 = n813 & ~n1157;
  assign n1162 = n1159 & ~n1161;
  assign n1163 = ~n1160 & ~n1162;
  assign n1164 = n1156 & n1163;
  assign n1165 = ~n1154 & ~n1164;
  assign n1166 = n1144 & ~n1151;
  assign n1167 = ~n1152 & ~n1166;
  assign n1168 = ~n1165 & n1167;
  assign n1169 = ~n1152 & ~n1168;
  assign n1170 = n595 & ~n1107;
  assign n1171 = ~n595 & ~n1109;
  assign n1172 = ~n1170 & ~n1171;
  assign n1173 = ~n664 & n1114;
  assign n1174 = n664 & n1112;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = ~n1172 & n1175;
  assign n1177 = n519 & n881;
  assign n1178 = ~n519 & n883;
  assign n1179 = ~n511 & n680;
  assign n1180 = n511 & n885;
  assign n1181 = ~n1177 & ~n1178;
  assign n1182 = ~n1179 & ~n1180;
  assign n1183 = n1181 & n1182;
  assign n1184 = n1176 & n1183;
  assign n1185 = ~n1176 & ~n1183;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = n453 & n658;
  assign n1188 = ~n453 & n660;
  assign n1189 = n669 & ~n869;
  assign n1190 = n666 & n869;
  assign n1191 = ~n1187 & ~n1188;
  assign n1192 = ~n1189 & ~n1190;
  assign n1193 = n1191 & n1192;
  assign n1194 = n1186 & n1193;
  assign n1195 = ~n1184 & ~n1194;
  assign n1196 = ~n1106 & ~n1117;
  assign n1197 = ~n1118 & ~n1196;
  assign n1198 = ~n1195 & n1197;
  assign n1199 = pi4  & pi22 ;
  assign n1200 = pi4  & ~n52;
  assign n1201 = n54 & ~n1200;
  assign n1202 = ~n1199 & ~n1201;
  assign n1203 = ~n504 & ~n1202;
  assign n1204 = ~n991 & n1203;
  assign n1205 = n991 & ~n1203;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = ~n813 & n1040;
  assign n1208 = ~n1157 & ~n1207;
  assign n1209 = n664 & ~n1208;
  assign n1210 = ~n1041 & ~n1158;
  assign n1211 = ~n664 & n1210;
  assign n1212 = n1041 & ~n1157;
  assign n1213 = ~n605 & n1212;
  assign n1214 = ~n1040 & n1161;
  assign n1215 = n605 & n1214;
  assign n1216 = ~n1209 & ~n1211;
  assign n1217 = ~n1213 & ~n1215;
  assign n1218 = n1216 & n1217;
  assign n1219 = n1206 & n1218;
  assign n1220 = ~n1204 & ~n1219;
  assign n1221 = n586 & ~n1046;
  assign n1222 = n589 & n1046;
  assign n1223 = n504 & ~n748;
  assign n1224 = ~n749 & ~n1223;
  assign n1225 = n584 & ~n1224;
  assign n1226 = ~n1221 & ~n1225;
  assign n1227 = ~n1222 & n1226;
  assign n1228 = ~n1220 & n1227;
  assign n1229 = n1220 & ~n1227;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = ~n511 & n881;
  assign n1232 = n511 & n883;
  assign n1233 = ~n453 & n885;
  assign n1234 = n453 & n680;
  assign n1235 = ~n1231 & ~n1232;
  assign n1236 = ~n1233 & ~n1234;
  assign n1237 = n1235 & n1236;
  assign n1238 = ~n519 & ~n1107;
  assign n1239 = n519 & ~n1109;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = ~n595 & n1112;
  assign n1242 = n595 & n1114;
  assign n1243 = ~n1241 & ~n1242;
  assign n1244 = ~n1240 & n1243;
  assign n1245 = n1237 & n1244;
  assign n1246 = ~n1237 & ~n1244;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = n658 & ~n869;
  assign n1249 = n660 & n869;
  assign n1250 = n666 & ~n748;
  assign n1251 = n669 & n748;
  assign n1252 = ~n1248 & ~n1249;
  assign n1253 = ~n1250 & ~n1251;
  assign n1254 = n1252 & n1253;
  assign n1255 = n1247 & n1254;
  assign n1256 = ~n1245 & ~n1255;
  assign n1257 = n1230 & ~n1256;
  assign n1258 = ~n1228 & ~n1257;
  assign n1259 = n1195 & ~n1197;
  assign n1260 = ~n1198 & ~n1259;
  assign n1261 = ~n1258 & n1260;
  assign n1262 = ~n1198 & ~n1261;
  assign n1263 = ~n1169 & ~n1262;
  assign n1264 = ~n1124 & ~n1126;
  assign n1265 = ~n1127 & ~n1264;
  assign n1266 = n1169 & n1262;
  assign n1267 = ~n1263 & ~n1266;
  assign n1268 = n1265 & n1267;
  assign n1269 = ~n1263 & ~n1268;
  assign n1270 = ~n1133 & ~n1135;
  assign n1271 = ~n1136 & ~n1270;
  assign n1272 = ~n1269 & n1271;
  assign n1273 = ~n1156 & ~n1163;
  assign n1274 = ~n1164 & ~n1273;
  assign n1275 = ~n1186 & ~n1193;
  assign n1276 = ~n1194 & ~n1275;
  assign n1277 = n1274 & n1276;
  assign n1278 = ~pi22  & ~n51;
  assign n1279 = ~pi3  & ~n1278;
  assign n1280 = pi3  & n1278;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = ~n504 & n1281;
  assign n1283 = ~n132 & ~n190;
  assign n1284 = ~n274 & ~n384;
  assign n1285 = n1283 & n1284;
  assign n1286 = n344 & n766;
  assign n1287 = n775 & n1286;
  assign n1288 = n1285 & n1287;
  assign n1289 = ~n180 & ~n189;
  assign n1290 = ~n201 & ~n311;
  assign n1291 = ~n317 & ~n436;
  assign n1292 = ~n552 & ~n564;
  assign n1293 = ~n764 & n1292;
  assign n1294 = n1290 & n1291;
  assign n1295 = n1289 & n1294;
  assign n1296 = n1293 & n1295;
  assign n1297 = n278 & ~n433;
  assign n1298 = ~n200 & ~n249;
  assign n1299 = ~n279 & ~n372;
  assign n1300 = ~n380 & n1299;
  assign n1301 = n326 & n1298;
  assign n1302 = n645 & n846;
  assign n1303 = n1301 & n1302;
  assign n1304 = n432 & n1300;
  assign n1305 = n1297 & n1304;
  assign n1306 = n1303 & n1305;
  assign n1307 = ~n341 & ~n530;
  assign n1308 = ~n137 & ~n284;
  assign n1309 = ~n356 & ~n461;
  assign n1310 = ~n630 & n1309;
  assign n1311 = n622 & n1308;
  assign n1312 = n1307 & n1311;
  assign n1313 = n1310 & n1312;
  assign n1314 = n488 & n1313;
  assign n1315 = n1288 & n1296;
  assign n1316 = n1314 & n1315;
  assign n1317 = n1306 & n1316;
  assign n1318 = ~n991 & ~n1317;
  assign n1319 = n605 & ~n991;
  assign n1320 = ~n1318 & ~n1319;
  assign n1321 = n1282 & ~n1320;
  assign n1322 = ~n1282 & n1320;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = n595 & ~n1210;
  assign n1325 = ~n595 & n1208;
  assign n1326 = ~n1324 & ~n1325;
  assign n1327 = ~n664 & n1214;
  assign n1328 = n664 & n1212;
  assign n1329 = ~n1327 & ~n1328;
  assign n1330 = ~n1326 & n1329;
  assign n1331 = n1323 & n1330;
  assign n1332 = ~n1321 & ~n1331;
  assign n1333 = n57 & n586;
  assign n1334 = ~n57 & n589;
  assign n1335 = n504 & n1046;
  assign n1336 = ~n1047 & ~n1335;
  assign n1337 = n584 & ~n1336;
  assign n1338 = ~n1333 & ~n1337;
  assign n1339 = ~n1334 & n1338;
  assign n1340 = ~n1332 & n1339;
  assign n1341 = n1332 & ~n1339;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = n453 & n881;
  assign n1344 = ~n453 & n883;
  assign n1345 = n680 & ~n869;
  assign n1346 = n869 & n885;
  assign n1347 = ~n1343 & ~n1344;
  assign n1348 = ~n1345 & ~n1346;
  assign n1349 = n1347 & n1348;
  assign n1350 = n511 & ~n1107;
  assign n1351 = ~n511 & ~n1109;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = ~n519 & n1114;
  assign n1354 = n519 & n1112;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = ~n1352 & n1355;
  assign n1357 = n1349 & n1356;
  assign n1358 = ~n1349 & ~n1356;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = n658 & n748;
  assign n1361 = n660 & ~n748;
  assign n1362 = n669 & ~n1046;
  assign n1363 = n666 & n1046;
  assign n1364 = ~n1360 & ~n1361;
  assign n1365 = ~n1362 & ~n1363;
  assign n1366 = n1364 & n1365;
  assign n1367 = n1359 & n1366;
  assign n1368 = ~n1357 & ~n1367;
  assign n1369 = n1342 & ~n1368;
  assign n1370 = ~n1340 & ~n1369;
  assign n1371 = ~n1274 & ~n1276;
  assign n1372 = ~n1277 & ~n1371;
  assign n1373 = ~n1370 & n1372;
  assign n1374 = ~n1277 & ~n1373;
  assign n1375 = n1165 & ~n1167;
  assign n1376 = ~n1168 & ~n1375;
  assign n1377 = ~n1374 & n1376;
  assign n1378 = n1374 & ~n1376;
  assign n1379 = ~n1377 & ~n1378;
  assign n1380 = n1258 & ~n1260;
  assign n1381 = ~n1261 & ~n1380;
  assign n1382 = n1379 & n1381;
  assign n1383 = ~n1377 & ~n1382;
  assign n1384 = ~n1265 & ~n1267;
  assign n1385 = ~n1268 & ~n1384;
  assign n1386 = ~n1383 & n1385;
  assign n1387 = n584 & n1281;
  assign n1388 = n588 & ~n1387;
  assign n1389 = ~n605 & n1318;
  assign n1390 = ~n605 & ~n1317;
  assign n1391 = n991 & ~n1390;
  assign n1392 = n664 & n1317;
  assign n1393 = ~n1389 & ~n1392;
  assign n1394 = ~n1391 & n1393;
  assign n1395 = n1388 & n1394;
  assign n1396 = n586 & ~n1202;
  assign n1397 = n589 & n1202;
  assign n1398 = ~n57 & n504;
  assign n1399 = ~n1153 & ~n1398;
  assign n1400 = n584 & ~n1399;
  assign n1401 = ~n1396 & ~n1400;
  assign n1402 = ~n1397 & n1401;
  assign n1403 = n1395 & n1402;
  assign n1404 = ~n869 & n881;
  assign n1405 = n869 & n883;
  assign n1406 = ~n748 & n885;
  assign n1407 = n680 & n748;
  assign n1408 = ~n1404 & ~n1405;
  assign n1409 = ~n1406 & ~n1407;
  assign n1410 = n1408 & n1409;
  assign n1411 = n658 & ~n1046;
  assign n1412 = n660 & n1046;
  assign n1413 = ~n57 & n666;
  assign n1414 = n57 & n669;
  assign n1415 = ~n1411 & ~n1412;
  assign n1416 = ~n1413 & ~n1414;
  assign n1417 = n1415 & n1416;
  assign n1418 = n1410 & n1417;
  assign n1419 = ~n1410 & ~n1417;
  assign n1420 = ~n1418 & ~n1419;
  assign n1421 = ~n453 & ~n1107;
  assign n1422 = n453 & ~n1109;
  assign n1423 = ~n1421 & ~n1422;
  assign n1424 = ~n511 & n1112;
  assign n1425 = n511 & n1114;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = ~n1423 & n1426;
  assign n1428 = n1420 & n1427;
  assign n1429 = ~n1418 & ~n1428;
  assign n1430 = ~n1395 & ~n1402;
  assign n1431 = ~n1403 & ~n1430;
  assign n1432 = ~n1429 & n1431;
  assign n1433 = ~n1403 & ~n1432;
  assign n1434 = ~n1206 & ~n1218;
  assign n1435 = ~n1219 & ~n1434;
  assign n1436 = ~n1433 & n1435;
  assign n1437 = n1433 & ~n1435;
  assign n1438 = ~n1436 & ~n1437;
  assign n1439 = ~n1247 & ~n1254;
  assign n1440 = ~n1255 & ~n1439;
  assign n1441 = n1438 & n1440;
  assign n1442 = ~n1436 & ~n1441;
  assign n1443 = ~n1230 & n1256;
  assign n1444 = ~n1257 & ~n1443;
  assign n1445 = ~n1442 & n1444;
  assign n1446 = n1442 & ~n1444;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = n1370 & ~n1372;
  assign n1449 = ~n1373 & ~n1448;
  assign n1450 = n1447 & n1449;
  assign n1451 = ~n1445 & ~n1450;
  assign n1452 = ~n1379 & ~n1381;
  assign n1453 = ~n1382 & ~n1452;
  assign n1454 = ~n1451 & n1453;
  assign n1455 = n586 & n1281;
  assign n1456 = n589 & ~n1281;
  assign n1457 = n504 & n1202;
  assign n1458 = ~n1203 & ~n1457;
  assign n1459 = n584 & ~n1458;
  assign n1460 = ~n1455 & ~n1459;
  assign n1461 = ~n1456 & n1460;
  assign n1462 = n519 & ~n1208;
  assign n1463 = ~n519 & n1210;
  assign n1464 = ~n595 & n1212;
  assign n1465 = n595 & n1214;
  assign n1466 = ~n1462 & ~n1463;
  assign n1467 = ~n1464 & ~n1465;
  assign n1468 = n1466 & n1467;
  assign n1469 = n1461 & n1468;
  assign n1470 = ~n1388 & ~n1394;
  assign n1471 = ~n1395 & ~n1470;
  assign n1472 = ~n1461 & ~n1468;
  assign n1473 = ~n1469 & ~n1472;
  assign n1474 = n1471 & n1473;
  assign n1475 = ~n1469 & ~n1474;
  assign n1476 = ~n1323 & ~n1330;
  assign n1477 = ~n1331 & ~n1476;
  assign n1478 = ~n1475 & n1477;
  assign n1479 = n1475 & ~n1477;
  assign n1480 = ~n1478 & ~n1479;
  assign n1481 = ~n1359 & ~n1366;
  assign n1482 = ~n1367 & ~n1481;
  assign n1483 = n1480 & n1482;
  assign n1484 = ~n1478 & ~n1483;
  assign n1485 = ~n1342 & n1368;
  assign n1486 = ~n1369 & ~n1485;
  assign n1487 = ~n1484 & n1486;
  assign n1488 = n1484 & ~n1486;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = ~n1438 & ~n1440;
  assign n1491 = ~n1441 & ~n1490;
  assign n1492 = n1489 & n1491;
  assign n1493 = ~n1487 & ~n1492;
  assign n1494 = ~n1447 & ~n1449;
  assign n1495 = ~n1450 & ~n1494;
  assign n1496 = ~n1493 & n1495;
  assign n1497 = n869 & ~n1107;
  assign n1498 = ~n869 & ~n1109;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = ~n453 & n1114;
  assign n1501 = n453 & n1112;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = ~n1499 & n1502;
  assign n1504 = n748 & n881;
  assign n1505 = ~n748 & n883;
  assign n1506 = n680 & ~n1046;
  assign n1507 = n885 & n1046;
  assign n1508 = ~n1504 & ~n1505;
  assign n1509 = ~n1506 & ~n1507;
  assign n1510 = n1508 & n1509;
  assign n1511 = n1503 & n1510;
  assign n1512 = n657 & n1281;
  assign n1513 = n665 & ~n1512;
  assign n1514 = ~n595 & n1318;
  assign n1515 = ~n595 & ~n1317;
  assign n1516 = n991 & ~n1515;
  assign n1517 = n519 & n1317;
  assign n1518 = ~n1514 & ~n1517;
  assign n1519 = ~n1516 & n1518;
  assign n1520 = n1513 & n1519;
  assign n1521 = ~n1503 & ~n1510;
  assign n1522 = ~n1511 & ~n1521;
  assign n1523 = n1520 & n1522;
  assign n1524 = ~n1511 & ~n1523;
  assign n1525 = n664 & n1318;
  assign n1526 = n664 & ~n1317;
  assign n1527 = n991 & ~n1526;
  assign n1528 = ~n595 & n1317;
  assign n1529 = ~n1525 & ~n1528;
  assign n1530 = ~n1527 & n1529;
  assign n1531 = n511 & ~n1210;
  assign n1532 = ~n511 & n1208;
  assign n1533 = ~n1531 & ~n1532;
  assign n1534 = ~n519 & n1214;
  assign n1535 = n519 & n1212;
  assign n1536 = ~n1534 & ~n1535;
  assign n1537 = ~n1533 & n1536;
  assign n1538 = n1530 & n1537;
  assign n1539 = ~n1530 & ~n1537;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = n57 & n658;
  assign n1542 = ~n57 & n660;
  assign n1543 = n669 & ~n1202;
  assign n1544 = n666 & n1202;
  assign n1545 = ~n1541 & ~n1542;
  assign n1546 = ~n1543 & ~n1544;
  assign n1547 = n1545 & n1546;
  assign n1548 = n1540 & n1547;
  assign n1549 = ~n1538 & ~n1548;
  assign n1550 = ~n1524 & ~n1549;
  assign n1551 = n1524 & n1549;
  assign n1552 = ~n1550 & ~n1551;
  assign n1553 = ~n1420 & ~n1427;
  assign n1554 = ~n1428 & ~n1553;
  assign n1555 = n1552 & n1554;
  assign n1556 = ~n1550 & ~n1555;
  assign n1557 = n1429 & ~n1431;
  assign n1558 = ~n1432 & ~n1557;
  assign n1559 = ~n1556 & n1558;
  assign n1560 = n1556 & ~n1558;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = ~n1480 & ~n1482;
  assign n1563 = ~n1483 & ~n1562;
  assign n1564 = n1561 & n1563;
  assign n1565 = ~n1559 & ~n1564;
  assign n1566 = ~n1489 & ~n1491;
  assign n1567 = ~n1492 & ~n1566;
  assign n1568 = ~n1565 & n1567;
  assign n1569 = n453 & ~n1208;
  assign n1570 = ~n453 & n1210;
  assign n1571 = ~n511 & n1212;
  assign n1572 = n511 & n1214;
  assign n1573 = ~n1569 & ~n1570;
  assign n1574 = ~n1571 & ~n1572;
  assign n1575 = n1573 & n1574;
  assign n1576 = n881 & ~n1046;
  assign n1577 = n883 & n1046;
  assign n1578 = ~n57 & n885;
  assign n1579 = n57 & n680;
  assign n1580 = ~n1576 & ~n1577;
  assign n1581 = ~n1578 & ~n1579;
  assign n1582 = n1580 & n1581;
  assign n1583 = n1575 & n1582;
  assign n1584 = ~n1575 & ~n1582;
  assign n1585 = ~n1583 & ~n1584;
  assign n1586 = ~n748 & ~n1107;
  assign n1587 = n748 & ~n1109;
  assign n1588 = ~n1586 & ~n1587;
  assign n1589 = ~n869 & n1112;
  assign n1590 = n869 & n1114;
  assign n1591 = ~n1589 & ~n1590;
  assign n1592 = ~n1588 & n1591;
  assign n1593 = n1585 & n1592;
  assign n1594 = ~n1583 & ~n1593;
  assign n1595 = n1387 & ~n1594;
  assign n1596 = ~n1520 & ~n1522;
  assign n1597 = ~n1523 & ~n1596;
  assign n1598 = ~n1387 & n1594;
  assign n1599 = ~n1595 & ~n1598;
  assign n1600 = n1597 & n1599;
  assign n1601 = ~n1595 & ~n1600;
  assign n1602 = n1471 & ~n1473;
  assign n1603 = ~n1471 & n1473;
  assign n1604 = ~n1602 & ~n1603;
  assign n1605 = ~n1601 & ~n1604;
  assign n1606 = n1601 & n1604;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = ~n1552 & ~n1554;
  assign n1609 = ~n1555 & ~n1608;
  assign n1610 = n1607 & n1609;
  assign n1611 = ~n1605 & ~n1610;
  assign n1612 = ~n1561 & ~n1563;
  assign n1613 = ~n1564 & ~n1612;
  assign n1614 = ~n1611 & n1613;
  assign n1615 = n1611 & ~n1613;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = ~n1513 & ~n1519;
  assign n1618 = ~n1520 & ~n1617;
  assign n1619 = n658 & ~n1202;
  assign n1620 = n660 & n1202;
  assign n1621 = n666 & ~n1281;
  assign n1622 = n669 & n1281;
  assign n1623 = ~n1619 & ~n1620;
  assign n1624 = ~n1621 & ~n1622;
  assign n1625 = n1623 & n1624;
  assign n1626 = n1618 & n1625;
  assign n1627 = n519 & n1318;
  assign n1628 = n519 & ~n1317;
  assign n1629 = n991 & ~n1628;
  assign n1630 = ~n511 & n1317;
  assign n1631 = ~n1627 & ~n1630;
  assign n1632 = ~n1629 & n1631;
  assign n1633 = n869 & ~n1210;
  assign n1634 = ~n869 & n1208;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = ~n453 & n1214;
  assign n1637 = n453 & n1212;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = ~n1635 & n1638;
  assign n1640 = n1632 & n1639;
  assign n1641 = ~n1632 & ~n1639;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = n1046 & ~n1107;
  assign n1644 = ~n1046 & ~n1109;
  assign n1645 = ~n1643 & ~n1644;
  assign n1646 = ~n748 & n1114;
  assign n1647 = n748 & n1112;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = ~n1645 & n1648;
  assign n1650 = n1642 & n1649;
  assign n1651 = ~n1640 & ~n1650;
  assign n1652 = ~n1618 & ~n1625;
  assign n1653 = ~n1626 & ~n1652;
  assign n1654 = ~n1651 & n1653;
  assign n1655 = ~n1626 & ~n1654;
  assign n1656 = ~n1540 & ~n1547;
  assign n1657 = ~n1548 & ~n1656;
  assign n1658 = ~n1655 & n1657;
  assign n1659 = ~n1597 & ~n1599;
  assign n1660 = ~n1600 & ~n1659;
  assign n1661 = n1655 & ~n1657;
  assign n1662 = ~n1658 & ~n1661;
  assign n1663 = n1660 & n1662;
  assign n1664 = ~n1658 & ~n1663;
  assign n1665 = n676 & n1281;
  assign n1666 = n449 & ~n1665;
  assign n1667 = ~n511 & n1318;
  assign n1668 = ~n511 & ~n1317;
  assign n1669 = n991 & ~n1668;
  assign n1670 = n453 & n1317;
  assign n1671 = ~n1667 & ~n1670;
  assign n1672 = ~n1669 & n1671;
  assign n1673 = n1666 & n1672;
  assign n1674 = n57 & n881;
  assign n1675 = ~n57 & n883;
  assign n1676 = n680 & ~n1202;
  assign n1677 = n885 & n1202;
  assign n1678 = ~n1674 & ~n1675;
  assign n1679 = ~n1676 & ~n1677;
  assign n1680 = n1678 & n1679;
  assign n1681 = n1673 & n1680;
  assign n1682 = ~n1673 & ~n1680;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = n1512 & n1683;
  assign n1685 = ~n1681 & ~n1684;
  assign n1686 = ~n1585 & ~n1592;
  assign n1687 = ~n1593 & ~n1686;
  assign n1688 = ~n1685 & n1687;
  assign n1689 = n1685 & ~n1687;
  assign n1690 = ~n1688 & ~n1689;
  assign n1691 = n1651 & ~n1653;
  assign n1692 = ~n1654 & ~n1691;
  assign n1693 = n1690 & n1692;
  assign n1694 = ~n1688 & ~n1693;
  assign n1695 = n748 & ~n1208;
  assign n1696 = ~n748 & n1210;
  assign n1697 = ~n869 & n1212;
  assign n1698 = n869 & n1214;
  assign n1699 = ~n1695 & ~n1696;
  assign n1700 = ~n1697 & ~n1698;
  assign n1701 = n1699 & n1700;
  assign n1702 = ~n57 & ~n1107;
  assign n1703 = n57 & ~n1109;
  assign n1704 = ~n1702 & ~n1703;
  assign n1705 = ~n1046 & n1112;
  assign n1706 = n1046 & n1114;
  assign n1707 = ~n1705 & ~n1706;
  assign n1708 = ~n1704 & n1707;
  assign n1709 = n1701 & n1708;
  assign n1710 = ~n1701 & ~n1708;
  assign n1711 = ~n1709 & ~n1710;
  assign n1712 = n881 & ~n1202;
  assign n1713 = n883 & n1202;
  assign n1714 = n885 & ~n1281;
  assign n1715 = n680 & n1281;
  assign n1716 = ~n1712 & ~n1713;
  assign n1717 = ~n1714 & ~n1715;
  assign n1718 = n1716 & n1717;
  assign n1719 = n1711 & n1718;
  assign n1720 = ~n1709 & ~n1719;
  assign n1721 = ~n1642 & ~n1649;
  assign n1722 = ~n1650 & ~n1721;
  assign n1723 = ~n1720 & n1722;
  assign n1724 = ~n1512 & ~n1683;
  assign n1725 = ~n1684 & ~n1724;
  assign n1726 = n1720 & ~n1722;
  assign n1727 = ~n1723 & ~n1726;
  assign n1728 = n1725 & n1727;
  assign n1729 = ~n1723 & ~n1728;
  assign n1730 = ~n1666 & ~n1672;
  assign n1731 = ~n1673 & ~n1730;
  assign n1732 = n453 & n1318;
  assign n1733 = n453 & ~n1317;
  assign n1734 = n991 & ~n1733;
  assign n1735 = ~n869 & n1317;
  assign n1736 = ~n1732 & ~n1735;
  assign n1737 = ~n1734 & n1736;
  assign n1738 = n1046 & ~n1210;
  assign n1739 = ~n1046 & n1208;
  assign n1740 = ~n1738 & ~n1739;
  assign n1741 = ~n748 & n1214;
  assign n1742 = n748 & n1212;
  assign n1743 = ~n1741 & ~n1742;
  assign n1744 = ~n1740 & n1743;
  assign n1745 = n1737 & n1744;
  assign n1746 = ~n1737 & ~n1744;
  assign n1747 = ~n1745 & ~n1746;
  assign n1748 = ~n1107 & n1202;
  assign n1749 = ~n1109 & ~n1202;
  assign n1750 = ~n1748 & ~n1749;
  assign n1751 = ~n57 & n1114;
  assign n1752 = n57 & n1112;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = ~n1750 & n1753;
  assign n1755 = n1747 & n1754;
  assign n1756 = ~n1745 & ~n1755;
  assign n1757 = n1731 & ~n1756;
  assign n1758 = ~n1731 & n1756;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = ~n1711 & ~n1718;
  assign n1761 = ~n1719 & ~n1760;
  assign n1762 = n1759 & n1761;
  assign n1763 = ~n1757 & ~n1762;
  assign n1764 = n1053 & n1281;
  assign n1765 = n862 & ~n1764;
  assign n1766 = ~n869 & n1318;
  assign n1767 = ~n869 & ~n1317;
  assign n1768 = n991 & ~n1767;
  assign n1769 = n748 & n1317;
  assign n1770 = ~n1766 & ~n1769;
  assign n1771 = ~n1768 & n1770;
  assign n1772 = n1765 & n1771;
  assign n1773 = n1665 & n1772;
  assign n1774 = n57 & ~n1208;
  assign n1775 = ~n57 & n1210;
  assign n1776 = ~n1046 & n1212;
  assign n1777 = n1046 & n1214;
  assign n1778 = ~n1774 & ~n1775;
  assign n1779 = ~n1776 & ~n1777;
  assign n1780 = n1778 & n1779;
  assign n1781 = ~n1107 & ~n1281;
  assign n1782 = ~n1109 & n1281;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = n1112 & ~n1202;
  assign n1785 = n1114 & n1202;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = ~n1783 & n1786;
  assign n1788 = n1780 & n1787;
  assign n1789 = ~n1765 & ~n1771;
  assign n1790 = ~n1772 & ~n1789;
  assign n1791 = ~n1780 & ~n1787;
  assign n1792 = ~n1788 & ~n1791;
  assign n1793 = n1790 & n1792;
  assign n1794 = ~n1788 & ~n1793;
  assign n1795 = ~n1665 & ~n1772;
  assign n1796 = ~n1773 & ~n1795;
  assign n1797 = ~n1794 & n1796;
  assign n1798 = ~n1773 & ~n1797;
  assign n1799 = n1794 & ~n1796;
  assign n1800 = ~n1797 & ~n1799;
  assign n1801 = n748 & n1318;
  assign n1802 = n748 & ~n1317;
  assign n1803 = n991 & ~n1802;
  assign n1804 = ~n1046 & n1317;
  assign n1805 = ~n1801 & ~n1804;
  assign n1806 = ~n1803 & n1805;
  assign n1807 = n1202 & ~n1210;
  assign n1808 = ~n1202 & n1208;
  assign n1809 = ~n1807 & ~n1808;
  assign n1810 = ~n57 & n1214;
  assign n1811 = n57 & n1212;
  assign n1812 = ~n1810 & ~n1811;
  assign n1813 = ~n1809 & n1812;
  assign n1814 = n1806 & n1813;
  assign n1815 = ~n1157 & n1281;
  assign n1816 = n1041 & ~n1815;
  assign n1817 = ~n1046 & n1318;
  assign n1818 = ~n1046 & ~n1317;
  assign n1819 = n991 & ~n1818;
  assign n1820 = n57 & n1317;
  assign n1821 = ~n1817 & ~n1820;
  assign n1822 = ~n1819 & n1821;
  assign n1823 = n1816 & n1822;
  assign n1824 = ~n1806 & ~n1813;
  assign n1825 = ~n1814 & ~n1824;
  assign n1826 = n1823 & n1825;
  assign n1827 = ~n1814 & ~n1826;
  assign n1828 = ~n1790 & ~n1792;
  assign n1829 = ~n1793 & ~n1828;
  assign n1830 = n1827 & ~n1829;
  assign n1831 = ~n1827 & n1829;
  assign n1832 = ~n1202 & ~n1317;
  assign n1833 = ~n991 & ~n1281;
  assign n1834 = ~n1832 & n1833;
  assign n1835 = n57 & n1318;
  assign n1836 = n57 & ~n1317;
  assign n1837 = n991 & ~n1836;
  assign n1838 = ~n1202 & n1317;
  assign n1839 = ~n1835 & ~n1838;
  assign n1840 = ~n1837 & n1839;
  assign n1841 = n1158 & n1281;
  assign n1842 = n1840 & n1841;
  assign n1843 = ~n1834 & ~n1842;
  assign n1844 = ~n1840 & ~n1841;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = ~n1816 & ~n1822;
  assign n1847 = ~n1823 & ~n1846;
  assign n1848 = ~n1210 & ~n1281;
  assign n1849 = n1208 & n1281;
  assign n1850 = ~n1848 & ~n1849;
  assign n1851 = ~n1202 & n1212;
  assign n1852 = n1202 & n1214;
  assign n1853 = ~n1851 & ~n1852;
  assign n1854 = ~n1850 & n1853;
  assign n1855 = n1847 & n1854;
  assign n1856 = ~n1845 & ~n1855;
  assign n1857 = ~n1847 & ~n1854;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = ~n1823 & ~n1825;
  assign n1860 = ~n1826 & ~n1859;
  assign n1861 = n1764 & n1860;
  assign n1862 = ~n1858 & ~n1861;
  assign n1863 = ~n1764 & ~n1860;
  assign n1864 = ~n1862 & ~n1863;
  assign n1865 = ~n1831 & ~n1864;
  assign n1866 = ~n1830 & ~n1865;
  assign n1867 = n1800 & n1866;
  assign n1868 = ~n1800 & ~n1866;
  assign n1869 = ~n1747 & ~n1754;
  assign n1870 = ~n1755 & ~n1869;
  assign n1871 = ~n1868 & n1870;
  assign n1872 = ~n1867 & ~n1871;
  assign n1873 = ~n1798 & ~n1872;
  assign n1874 = n1798 & n1872;
  assign n1875 = ~n1759 & ~n1761;
  assign n1876 = ~n1762 & ~n1875;
  assign n1877 = ~n1874 & n1876;
  assign n1878 = ~n1873 & ~n1877;
  assign n1879 = ~n1763 & ~n1878;
  assign n1880 = n1763 & n1878;
  assign n1881 = ~n1725 & ~n1727;
  assign n1882 = ~n1728 & ~n1881;
  assign n1883 = ~n1880 & n1882;
  assign n1884 = ~n1879 & ~n1883;
  assign n1885 = ~n1729 & ~n1884;
  assign n1886 = n1729 & n1884;
  assign n1887 = ~n1690 & ~n1692;
  assign n1888 = ~n1693 & ~n1887;
  assign n1889 = ~n1886 & n1888;
  assign n1890 = ~n1885 & ~n1889;
  assign n1891 = ~n1694 & ~n1890;
  assign n1892 = n1694 & n1890;
  assign n1893 = ~n1660 & ~n1662;
  assign n1894 = ~n1663 & ~n1893;
  assign n1895 = ~n1892 & n1894;
  assign n1896 = ~n1891 & ~n1895;
  assign n1897 = ~n1664 & ~n1896;
  assign n1898 = n1664 & n1896;
  assign n1899 = ~n1607 & ~n1609;
  assign n1900 = ~n1610 & ~n1899;
  assign n1901 = ~n1898 & n1900;
  assign n1902 = ~n1897 & ~n1901;
  assign n1903 = n1616 & ~n1902;
  assign n1904 = ~n1614 & ~n1903;
  assign n1905 = n1565 & ~n1567;
  assign n1906 = ~n1568 & ~n1905;
  assign n1907 = ~n1904 & n1906;
  assign n1908 = ~n1568 & ~n1907;
  assign n1909 = n1493 & ~n1495;
  assign n1910 = ~n1496 & ~n1909;
  assign n1911 = ~n1908 & n1910;
  assign n1912 = ~n1496 & ~n1911;
  assign n1913 = n1451 & ~n1453;
  assign n1914 = ~n1454 & ~n1913;
  assign n1915 = ~n1912 & n1914;
  assign n1916 = ~n1454 & ~n1915;
  assign n1917 = n1383 & ~n1385;
  assign n1918 = ~n1386 & ~n1917;
  assign n1919 = ~n1916 & n1918;
  assign n1920 = ~n1386 & ~n1919;
  assign n1921 = n1269 & ~n1271;
  assign n1922 = ~n1272 & ~n1921;
  assign n1923 = ~n1920 & n1922;
  assign n1924 = ~n1272 & ~n1923;
  assign n1925 = n1137 & ~n1139;
  assign n1926 = ~n1140 & ~n1925;
  assign n1927 = ~n1924 & n1926;
  assign n1928 = ~n1140 & ~n1927;
  assign n1929 = n1086 & ~n1088;
  assign n1930 = ~n1089 & ~n1929;
  assign n1931 = ~n1928 & n1930;
  assign n1932 = ~n1089 & ~n1931;
  assign n1933 = n922 & ~n924;
  assign n1934 = ~n925 & ~n1933;
  assign n1935 = ~n1932 & n1934;
  assign n1936 = ~n925 & ~n1935;
  assign n1937 = n722 & ~n743;
  assign n1938 = ~n744 & ~n1937;
  assign n1939 = ~n1936 & n1938;
  assign n1940 = ~n744 & ~n1939;
  assign n1941 = ~n732 & ~n741;
  assign n1942 = ~n735 & ~n738;
  assign n1943 = n583 & n727;
  assign n1944 = ~n588 & ~n1943;
  assign n1945 = n582 & ~n605;
  assign n1946 = ~n1944 & ~n1945;
  assign n1947 = ~n710 & n1946;
  assign n1948 = n710 & ~n1946;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = ~n1942 & n1949;
  assign n1951 = n1942 & ~n1949;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = ~n1941 & n1952;
  assign n1954 = n1941 & ~n1952;
  assign n1955 = ~n1953 & ~n1954;
  assign n1956 = ~n1940 & n1955;
  assign n1957 = n1940 & ~n1955;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = ~n309 & ~n343;
  assign n1960 = ~n370 & ~n412;
  assign n1961 = n1959 & n1960;
  assign n1962 = n753 & n1961;
  assign n1963 = n277 & n1962;
  assign n1964 = ~n129 & ~n530;
  assign n1965 = n846 & n1964;
  assign n1966 = ~n210 & ~n218;
  assign n1967 = ~n311 & n1966;
  assign n1968 = n633 & n1967;
  assign n1969 = n146 & ~n317;
  assign n1970 = n379 & n1969;
  assign n1971 = n184 & n833;
  assign n1972 = n967 & n1965;
  assign n1973 = n1971 & n1972;
  assign n1974 = n1968 & n1970;
  assign n1975 = n1973 & n1974;
  assign n1976 = ~n176 & ~n294;
  assign n1977 = ~n310 & ~n318;
  assign n1978 = ~n564 & n1977;
  assign n1979 = n1976 & n1978;
  assign n1980 = ~n148 & ~n188;
  assign n1981 = ~n192 & ~n209;
  assign n1982 = ~n299 & ~n342;
  assign n1983 = ~n793 & n1982;
  assign n1984 = n1980 & n1981;
  assign n1985 = n114 & n1984;
  assign n1986 = n1983 & n1985;
  assign n1987 = n1979 & n1986;
  assign n1988 = ~n222 & ~n282;
  assign n1989 = ~n576 & n1988;
  assign n1990 = ~n156 & ~n207;
  assign n1991 = ~n262 & ~n380;
  assign n1992 = n1990 & n1991;
  assign n1993 = n141 & n305;
  assign n1994 = n408 & n459;
  assign n1995 = n1993 & n1994;
  assign n1996 = n1989 & n1992;
  assign n1997 = n1995 & n1996;
  assign n1998 = n245 & n1997;
  assign n1999 = n1963 & n1998;
  assign n2000 = n1975 & n1987;
  assign n2001 = n1999 & n2000;
  assign n2002 = ~n1958 & ~n2001;
  assign n2003 = n1936 & ~n1938;
  assign n2004 = ~n1939 & ~n2003;
  assign n2005 = ~n210 & ~n240;
  assign n2006 = ~n248 & ~n294;
  assign n2007 = ~n343 & n2006;
  assign n2008 = n312 & n2005;
  assign n2009 = n414 & n614;
  assign n2010 = n2008 & n2009;
  assign n2011 = n195 & n2007;
  assign n2012 = n270 & n777;
  assign n2013 = n2011 & n2012;
  assign n2014 = n2010 & n2013;
  assign n2015 = n628 & n825;
  assign n2016 = n2014 & n2015;
  assign n2017 = n978 & n2016;
  assign n2018 = ~n2004 & ~n2017;
  assign n2019 = n1932 & ~n1934;
  assign n2020 = ~n1935 & ~n2019;
  assign n2021 = ~n149 & ~n176;
  assign n2022 = ~n185 & ~n225;
  assign n2023 = ~n237 & n2022;
  assign n2024 = n553 & n2021;
  assign n2025 = n2023 & n2024;
  assign n2026 = ~n190 & ~n314;
  assign n2027 = ~n188 & ~n279;
  assign n2028 = n2026 & n2027;
  assign n2029 = n635 & n2028;
  assign n2030 = n407 & n2029;
  assign n2031 = n2025 & n2030;
  assign n2032 = ~n171 & ~n454;
  assign n2033 = ~n199 & ~n372;
  assign n2034 = ~n262 & ~n318;
  assign n2035 = ~n481 & n2034;
  assign n2036 = ~n209 & ~n306;
  assign n2037 = n347 & n2036;
  assign n2038 = n614 & n2032;
  assign n2039 = n2033 & n2038;
  assign n2040 = n1965 & n2037;
  assign n2041 = n1989 & n2035;
  assign n2042 = n2040 & n2041;
  assign n2043 = n402 & n2039;
  assign n2044 = n2042 & n2043;
  assign n2045 = ~n198 & ~n235;
  assign n2046 = ~n284 & n2045;
  assign n2047 = ~n134 & ~n233;
  assign n2048 = ~n251 & n2047;
  assign n2049 = ~n378 & n409;
  assign n2050 = n565 & n645;
  assign n2051 = n943 & n2050;
  assign n2052 = n2046 & n2049;
  assign n2053 = n2048 & n2052;
  assign n2054 = n440 & n2051;
  assign n2055 = n2053 & n2054;
  assign n2056 = n2031 & n2055;
  assign n2057 = n2044 & n2056;
  assign n2058 = ~n2020 & ~n2057;
  assign n2059 = n1928 & ~n1930;
  assign n2060 = ~n1931 & ~n2059;
  assign n2061 = ~n208 & ~n224;
  assign n2062 = ~n380 & ~n520;
  assign n2063 = ~n630 & n2062;
  assign n2064 = n308 & n2061;
  assign n2065 = n456 & n2064;
  assign n2066 = n540 & n2063;
  assign n2067 = n2046 & n2066;
  assign n2068 = n2065 & n2067;
  assign n2069 = ~n132 & ~n237;
  assign n2070 = ~n248 & n2069;
  assign n2071 = ~n140 & ~n295;
  assign n2072 = ~n327 & n2071;
  assign n2073 = n2044 & n2072;
  assign n2074 = ~n192 & ~n427;
  assign n2075 = ~n233 & ~n268;
  assign n2076 = n2074 & n2075;
  assign n2077 = n765 & n827;
  assign n2078 = n2076 & n2077;
  assign n2079 = n1297 & n2070;
  assign n2080 = n2078 & n2079;
  assign n2081 = n1963 & n2080;
  assign n2082 = n2068 & n2081;
  assign n2083 = n2073 & n2082;
  assign n2084 = ~n2060 & ~n2083;
  assign n2085 = n1924 & ~n1926;
  assign n2086 = ~n1927 & ~n2085;
  assign n2087 = ~n200 & ~n237;
  assign n2088 = ~n223 & ~n263;
  assign n2089 = ~n274 & ~n343;
  assign n2090 = n413 & n2089;
  assign n2091 = n645 & n958;
  assign n2092 = n2087 & n2088;
  assign n2093 = n2091 & n2092;
  assign n2094 = n2090 & n2093;
  assign n2095 = n803 & n2094;
  assign n2096 = ~n186 & ~n310;
  assign n2097 = n792 & n2096;
  assign n2098 = ~n189 & ~n372;
  assign n2099 = ~n154 & ~n180;
  assign n2100 = ~n240 & ~n309;
  assign n2101 = n2099 & n2100;
  assign n2102 = n2026 & n2098;
  assign n2103 = n2101 & n2102;
  assign n2104 = ~n137 & ~n156;
  assign n2105 = ~n182 & ~n345;
  assign n2106 = ~n403 & n2105;
  assign n2107 = n2104 & n2106;
  assign n2108 = ~n134 & ~n145;
  assign n2109 = ~n222 & ~n247;
  assign n2110 = ~n262 & ~n325;
  assign n2111 = n2109 & n2110;
  assign n2112 = n539 & n2108;
  assign n2113 = n2111 & n2112;
  assign n2114 = n2103 & n2113;
  assign n2115 = n2107 & n2114;
  assign n2116 = n2095 & n2115;
  assign n2117 = n2097 & n2116;
  assign n2118 = ~n2086 & ~n2117;
  assign n2119 = n1920 & ~n1922;
  assign n2120 = ~n1923 & ~n2119;
  assign n2121 = ~n188 & ~n220;
  assign n2122 = ~n548 & n2121;
  assign n2123 = n532 & n2122;
  assign n2124 = ~n154 & ~n345;
  assign n2125 = ~n153 & n187;
  assign n2126 = ~n182 & ~n196;
  assign n2127 = ~n310 & ~n403;
  assign n2128 = n529 & n752;
  assign n2129 = n783 & n2127;
  assign n2130 = n2128 & n2129;
  assign n2131 = n142 & n2130;
  assign n2132 = ~n356 & n455;
  assign n2133 = n629 & n960;
  assign n2134 = n2124 & n2126;
  assign n2135 = n2133 & n2134;
  assign n2136 = n328 & n2132;
  assign n2137 = n2125 & n2136;
  assign n2138 = n757 & n2135;
  assign n2139 = n2123 & n2138;
  assign n2140 = n2131 & n2137;
  assign n2141 = n2139 & n2140;
  assign n2142 = n841 & n2141;
  assign n2143 = ~n2120 & ~n2142;
  assign n2144 = n1916 & ~n1918;
  assign n2145 = ~n1919 & ~n2144;
  assign n2146 = ~n378 & ~n429;
  assign n2147 = ~n481 & n2146;
  assign n2148 = ~n248 & ~n325;
  assign n2149 = ~n119 & ~n181;
  assign n2150 = ~n201 & ~n458;
  assign n2151 = n2149 & n2150;
  assign n2152 = n319 & n2148;
  assign n2153 = n2151 & n2152;
  assign n2154 = n2147 & n2153;
  assign n2155 = n771 & n2154;
  assign n2156 = n90 & n115;
  assign n2157 = ~n264 & ~n380;
  assign n2158 = n2088 & n2157;
  assign n2159 = ~n272 & ~n280;
  assign n2160 = ~n345 & ~n384;
  assign n2161 = n2159 & n2160;
  assign n2162 = n622 & n2161;
  assign n2163 = n2158 & n2162;
  assign n2164 = n402 & n1030;
  assign n2165 = n2163 & n2164;
  assign n2166 = ~n152 & n409;
  assign n2167 = n2165 & n2166;
  assign n2168 = ~n199 & ~n279;
  assign n2169 = ~n370 & ~n543;
  assign n2170 = n2168 & n2169;
  assign n2171 = n413 & n778;
  assign n2172 = n2170 & n2171;
  assign n2173 = ~n236 & ~n2156;
  assign n2174 = ~n113 & n2173;
  assign n2175 = ~n192 & ~n274;
  assign n2176 = ~n454 & n2175;
  assign n2177 = n146 & n2174;
  assign n2178 = n2176 & n2177;
  assign n2179 = n2172 & n2178;
  assign n2180 = n2155 & n2179;
  assign n2181 = n2167 & n2180;
  assign n2182 = ~n2145 & ~n2181;
  assign n2183 = n1912 & ~n1914;
  assign n2184 = ~n1915 & ~n2183;
  assign n2185 = ~n156 & ~n299;
  assign n2186 = ~n272 & ~n310;
  assign n2187 = ~n404 & ~n436;
  assign n2188 = n2186 & n2187;
  assign n2189 = n767 & n2188;
  assign n2190 = n376 & n475;
  assign n2191 = n2048 & n2190;
  assign n2192 = n2189 & n2191;
  assign n2193 = ~n145 & ~n380;
  assign n2194 = n482 & n2193;
  assign n2195 = n538 & n959;
  assign n2196 = n2194 & n2195;
  assign n2197 = ~n222 & ~n295;
  assign n2198 = ~n303 & ~n341;
  assign n2199 = ~n372 & ~n378;
  assign n2200 = ~n564 & n2199;
  assign n2201 = n2197 & n2198;
  assign n2202 = n346 & n426;
  assign n2203 = n2185 & n2202;
  assign n2204 = n2200 & n2201;
  assign n2205 = n833 & n2204;
  assign n2206 = n2196 & n2203;
  assign n2207 = n2205 & n2206;
  assign n2208 = n217 & n2207;
  assign n2209 = n2192 & n2208;
  assign n2210 = ~n2184 & ~n2209;
  assign n2211 = n1908 & ~n1910;
  assign n2212 = ~n1911 & ~n2211;
  assign n2213 = ~n197 & ~n207;
  assign n2214 = ~n294 & n622;
  assign n2215 = ~n113 & ~n224;
  assign n2216 = ~n295 & ~n429;
  assign n2217 = ~n370 & ~n630;
  assign n2218 = ~n267 & ~n298;
  assign n2219 = ~n520 & n2218;
  assign n2220 = n2217 & n2219;
  assign n2221 = ~n272 & n845;
  assign n2222 = n2215 & n2216;
  assign n2223 = n2221 & n2222;
  assign n2224 = n751 & n2070;
  assign n2225 = n2214 & n2224;
  assign n2226 = n2123 & n2223;
  assign n2227 = n2220 & n2226;
  assign n2228 = n2225 & n2227;
  assign n2229 = ~n125 & ~n185;
  assign n2230 = ~n249 & ~n262;
  assign n2231 = ~n436 & n2230;
  assign n2232 = n297 & n2229;
  assign n2233 = n456 & n765;
  assign n2234 = n2213 & n2233;
  assign n2235 = n2231 & n2232;
  assign n2236 = n2234 & n2235;
  assign n2237 = n830 & n2196;
  assign n2238 = n2236 & n2237;
  assign n2239 = n782 & n2238;
  assign n2240 = n421 & n2239;
  assign n2241 = n2228 & n2240;
  assign n2242 = ~n2212 & ~n2241;
  assign n2243 = n1904 & ~n1906;
  assign n2244 = ~n1907 & ~n2243;
  assign n2245 = ~n282 & ~n461;
  assign n2246 = ~n303 & ~n412;
  assign n2247 = ~n274 & ~n313;
  assign n2248 = ~n378 & n2247;
  assign n2249 = n2246 & n2248;
  assign n2250 = n121 & ~n499;
  assign n2251 = ~n144 & ~n268;
  assign n2252 = ~n530 & ~n2250;
  assign n2253 = n2251 & n2252;
  assign n2254 = ~n132 & ~n224;
  assign n2255 = ~n317 & ~n343;
  assign n2256 = ~n428 & n2255;
  assign n2257 = n2254 & n2256;
  assign n2258 = n2253 & n2257;
  assign n2259 = n2249 & n2258;
  assign n2260 = ~n134 & ~n190;
  assign n2261 = ~n200 & ~n309;
  assign n2262 = ~n399 & ~n543;
  assign n2263 = n2261 & n2262;
  assign n2264 = n312 & n2260;
  assign n2265 = n606 & n2216;
  assign n2266 = n2245 & n2265;
  assign n2267 = n2263 & n2264;
  assign n2268 = n302 & n2267;
  assign n2269 = n2266 & n2268;
  assign n2270 = n2131 & n2269;
  assign n2271 = n2259 & n2270;
  assign n2272 = ~n2244 & ~n2271;
  assign n2273 = ~n1616 & n1902;
  assign n2274 = ~n1903 & ~n2273;
  assign n2275 = ~n399 & ~n793;
  assign n2276 = ~n279 & ~n630;
  assign n2277 = n2275 & n2276;
  assign n2278 = n178 & n2277;
  assign n2279 = n195 & n970;
  assign n2280 = n2214 & n2279;
  assign n2281 = n774 & n2278;
  assign n2282 = n2280 & n2281;
  assign n2283 = n1975 & n2282;
  assign n2284 = n2192 & n2283;
  assign n2285 = n2274 & n2284;
  assign n2286 = n2244 & n2271;
  assign n2287 = ~n2272 & ~n2286;
  assign n2288 = ~n2285 & n2287;
  assign n2289 = ~n2272 & ~n2288;
  assign n2290 = n2212 & n2241;
  assign n2291 = ~n2242 & ~n2290;
  assign n2292 = ~n2289 & n2291;
  assign n2293 = ~n2242 & ~n2292;
  assign n2294 = n2184 & n2209;
  assign n2295 = ~n2210 & ~n2294;
  assign n2296 = ~n2293 & n2295;
  assign n2297 = ~n2210 & ~n2296;
  assign n2298 = n2145 & n2181;
  assign n2299 = ~n2182 & ~n2298;
  assign n2300 = ~n2297 & n2299;
  assign n2301 = ~n2182 & ~n2300;
  assign n2302 = n2120 & n2142;
  assign n2303 = ~n2143 & ~n2302;
  assign n2304 = ~n2301 & n2303;
  assign n2305 = ~n2143 & ~n2304;
  assign n2306 = n2086 & n2117;
  assign n2307 = ~n2118 & ~n2306;
  assign n2308 = ~n2305 & n2307;
  assign n2309 = ~n2118 & ~n2308;
  assign n2310 = n2060 & n2083;
  assign n2311 = ~n2084 & ~n2310;
  assign n2312 = ~n2309 & n2311;
  assign n2313 = ~n2084 & ~n2312;
  assign n2314 = n2020 & n2057;
  assign n2315 = ~n2058 & ~n2314;
  assign n2316 = ~n2313 & n2315;
  assign n2317 = ~n2058 & ~n2316;
  assign n2318 = n2004 & n2017;
  assign n2319 = ~n2018 & ~n2318;
  assign n2320 = ~n2317 & n2319;
  assign n2321 = ~n2018 & ~n2320;
  assign n2322 = n1958 & n2001;
  assign n2323 = ~n2002 & ~n2322;
  assign n2324 = ~n2321 & n2323;
  assign n2325 = ~n2002 & ~n2324;
  assign n2326 = ~n125 & ~n341;
  assign n2327 = ~n220 & ~n329;
  assign n2328 = ~n240 & ~n310;
  assign n2329 = ~n458 & n2328;
  assign n2330 = n2035 & n2329;
  assign n2331 = ~n119 & ~n303;
  assign n2332 = ~n520 & n2331;
  assign n2333 = n826 & n2332;
  assign n2334 = n549 & n629;
  assign n2335 = n765 & n2245;
  assign n2336 = n2326 & n2327;
  assign n2337 = n2335 & n2336;
  assign n2338 = n2334 & n2337;
  assign n2339 = n2330 & n2333;
  assign n2340 = n2338 & n2339;
  assign n2341 = n782 & n951;
  assign n2342 = n2340 & n2341;
  assign n2343 = n2167 & n2342;
  assign n2344 = ~n605 & ~n664;
  assign n2345 = n605 & n664;
  assign n2346 = ~n2344 & ~n2345;
  assign n2347 = ~n583 & ~n2346;
  assign n2348 = n583 & n2346;
  assign n2349 = ~n504 & ~n2347;
  assign n2350 = ~n2348 & n2349;
  assign n2351 = ~n1953 & ~n1956;
  assign n2352 = ~n1947 & ~n1950;
  assign n2353 = n2351 & ~n2352;
  assign n2354 = ~n2351 & n2352;
  assign n2355 = ~n2353 & ~n2354;
  assign n2356 = n2350 & n2355;
  assign n2357 = ~n2350 & ~n2355;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = ~n2343 & ~n2358;
  assign n2360 = n2343 & n2358;
  assign n2361 = ~n2359 & ~n2360;
  assign n2362 = ~n2325 & n2361;
  assign n2363 = n2325 & ~n2361;
  assign n2364 = ~n2362 & ~n2363;
  assign n2365 = pi2  & pi22 ;
  assign n2366 = pi2  & ~n50;
  assign n2367 = n1278 & ~n2366;
  assign n2368 = ~n2365 & ~n2367;
  assign n2369 = ~n1281 & ~n2368;
  assign n2370 = n1281 & n2368;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = ~n57 & ~n1202;
  assign n2373 = n57 & n1202;
  assign n2374 = ~n2372 & ~n2373;
  assign n2375 = ~n2371 & n2374;
  assign n2376 = n2364 & n2375;
  assign n2377 = n2321 & ~n2323;
  assign n2378 = ~n2324 & ~n2377;
  assign n2379 = ~n1202 & ~n1281;
  assign n2380 = n1202 & n1281;
  assign n2381 = ~n2379 & ~n2380;
  assign n2382 = n2371 & ~n2381;
  assign n2383 = n2378 & n2382;
  assign n2384 = n2317 & ~n2319;
  assign n2385 = ~n2320 & ~n2384;
  assign n2386 = n2371 & ~n2374;
  assign n2387 = n2381 & n2386;
  assign n2388 = n2385 & n2387;
  assign n2389 = ~n2371 & ~n2374;
  assign n2390 = n2378 & n2385;
  assign n2391 = n2313 & ~n2315;
  assign n2392 = ~n2316 & ~n2391;
  assign n2393 = n2385 & n2392;
  assign n2394 = n2309 & ~n2311;
  assign n2395 = ~n2312 & ~n2394;
  assign n2396 = n2392 & n2395;
  assign n2397 = n2305 & ~n2307;
  assign n2398 = ~n2308 & ~n2397;
  assign n2399 = n2395 & n2398;
  assign n2400 = n2301 & ~n2303;
  assign n2401 = ~n2304 & ~n2400;
  assign n2402 = n2398 & n2401;
  assign n2403 = n2297 & ~n2299;
  assign n2404 = ~n2300 & ~n2403;
  assign n2405 = n2401 & n2404;
  assign n2406 = n2293 & ~n2295;
  assign n2407 = ~n2296 & ~n2406;
  assign n2408 = n2404 & n2407;
  assign n2409 = n2289 & ~n2291;
  assign n2410 = ~n2292 & ~n2409;
  assign n2411 = n2407 & n2410;
  assign n2412 = ~n2407 & ~n2410;
  assign n2413 = ~n2411 & ~n2412;
  assign n2414 = ~n2274 & ~n2284;
  assign n2415 = ~n2285 & ~n2414;
  assign n2416 = ~n2410 & n2415;
  assign n2417 = n2285 & ~n2287;
  assign n2418 = ~n2288 & ~n2417;
  assign n2419 = ~n2416 & n2418;
  assign n2420 = n2413 & n2419;
  assign n2421 = ~n2411 & ~n2420;
  assign n2422 = ~n2404 & ~n2407;
  assign n2423 = ~n2408 & ~n2422;
  assign n2424 = ~n2421 & n2423;
  assign n2425 = ~n2408 & ~n2424;
  assign n2426 = ~n2401 & ~n2404;
  assign n2427 = ~n2405 & ~n2426;
  assign n2428 = ~n2425 & n2427;
  assign n2429 = ~n2405 & ~n2428;
  assign n2430 = ~n2398 & ~n2401;
  assign n2431 = ~n2402 & ~n2430;
  assign n2432 = ~n2429 & n2431;
  assign n2433 = ~n2402 & ~n2432;
  assign n2434 = ~n2395 & ~n2398;
  assign n2435 = ~n2399 & ~n2434;
  assign n2436 = ~n2433 & n2435;
  assign n2437 = ~n2399 & ~n2436;
  assign n2438 = ~n2392 & ~n2395;
  assign n2439 = ~n2396 & ~n2438;
  assign n2440 = ~n2437 & n2439;
  assign n2441 = ~n2396 & ~n2440;
  assign n2442 = ~n2385 & ~n2392;
  assign n2443 = ~n2393 & ~n2442;
  assign n2444 = ~n2441 & n2443;
  assign n2445 = ~n2393 & ~n2444;
  assign n2446 = ~n2378 & ~n2385;
  assign n2447 = ~n2390 & ~n2446;
  assign n2448 = ~n2445 & n2447;
  assign n2449 = ~n2390 & ~n2448;
  assign n2450 = n2364 & n2378;
  assign n2451 = ~n2364 & ~n2378;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = ~n2449 & n2452;
  assign n2454 = n2449 & ~n2452;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = n2389 & n2455;
  assign n2457 = ~n2383 & ~n2388;
  assign n2458 = ~n2376 & n2457;
  assign n2459 = ~n2456 & n2458;
  assign n2460 = n57 & ~n2459;
  assign n2461 = ~n57 & n2459;
  assign n2462 = ~n2460 & ~n2461;
  assign n2463 = ~n57 & ~n1046;
  assign n2464 = n57 & n1046;
  assign n2465 = ~n2463 & ~n2464;
  assign n2466 = ~n748 & ~n869;
  assign n2467 = n748 & n869;
  assign n2468 = ~n2466 & ~n2467;
  assign n2469 = ~n2465 & n2468;
  assign n2470 = n2395 & n2469;
  assign n2471 = ~n748 & ~n1046;
  assign n2472 = n748 & n1046;
  assign n2473 = ~n2471 & ~n2472;
  assign n2474 = n2465 & ~n2473;
  assign n2475 = n2398 & n2474;
  assign n2476 = n2465 & n2473;
  assign n2477 = ~n2468 & n2476;
  assign n2478 = n2401 & n2477;
  assign n2479 = ~n2465 & ~n2468;
  assign n2480 = n2433 & ~n2435;
  assign n2481 = ~n2436 & ~n2480;
  assign n2482 = n2479 & n2481;
  assign n2483 = ~n2475 & ~n2478;
  assign n2484 = ~n2470 & n2483;
  assign n2485 = ~n2482 & n2484;
  assign n2486 = n869 & ~n2485;
  assign n2487 = ~n869 & n2485;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = ~n519 & ~n595;
  assign n2490 = n519 & n595;
  assign n2491 = ~n2489 & ~n2490;
  assign n2492 = ~n2415 & ~n2491;
  assign n2493 = ~n453 & ~n869;
  assign n2494 = n453 & n869;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = ~n2415 & ~n2495;
  assign n2497 = ~n2415 & ~n2418;
  assign n2498 = ~n2287 & n2415;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = ~n511 & ~n519;
  assign n2501 = n511 & n519;
  assign n2502 = ~n2500 & ~n2501;
  assign n2503 = ~n2495 & ~n2502;
  assign n2504 = ~n2499 & n2503;
  assign n2505 = ~n453 & ~n511;
  assign n2506 = n453 & n511;
  assign n2507 = ~n2505 & ~n2506;
  assign n2508 = n2495 & ~n2507;
  assign n2509 = ~n2415 & n2508;
  assign n2510 = ~n2495 & n2502;
  assign n2511 = n2418 & n2510;
  assign n2512 = ~n2509 & ~n2511;
  assign n2513 = ~n2504 & n2512;
  assign n2514 = n519 & ~n2496;
  assign n2515 = n2513 & n2514;
  assign n2516 = n2410 & n2510;
  assign n2517 = n2495 & ~n2502;
  assign n2518 = n2507 & n2517;
  assign n2519 = ~n2415 & n2518;
  assign n2520 = n2418 & n2508;
  assign n2521 = n2410 & ~n2498;
  assign n2522 = ~n2410 & n2498;
  assign n2523 = ~n2521 & ~n2522;
  assign n2524 = n2503 & ~n2523;
  assign n2525 = ~n2519 & ~n2520;
  assign n2526 = ~n2516 & n2525;
  assign n2527 = ~n2524 & n2526;
  assign n2528 = n2515 & n2527;
  assign n2529 = n2492 & n2528;
  assign n2530 = n2407 & n2510;
  assign n2531 = n2418 & n2518;
  assign n2532 = n2410 & n2508;
  assign n2533 = ~n2413 & ~n2419;
  assign n2534 = ~n2420 & ~n2533;
  assign n2535 = n2503 & n2534;
  assign n2536 = ~n2531 & ~n2532;
  assign n2537 = ~n2530 & n2536;
  assign n2538 = ~n2535 & n2537;
  assign n2539 = n519 & ~n2538;
  assign n2540 = ~n519 & n2538;
  assign n2541 = ~n2539 & ~n2540;
  assign n2542 = ~n2492 & ~n2528;
  assign n2543 = ~n2529 & ~n2542;
  assign n2544 = n2541 & n2543;
  assign n2545 = ~n2529 & ~n2544;
  assign n2546 = n2404 & n2510;
  assign n2547 = n2407 & n2508;
  assign n2548 = n2410 & n2518;
  assign n2549 = n2421 & ~n2423;
  assign n2550 = ~n2424 & ~n2549;
  assign n2551 = n2503 & n2550;
  assign n2552 = ~n2547 & ~n2548;
  assign n2553 = ~n2546 & n2552;
  assign n2554 = ~n2551 & n2553;
  assign n2555 = ~n519 & n2554;
  assign n2556 = n519 & ~n2554;
  assign n2557 = ~n2555 & ~n2556;
  assign n2558 = ~n2346 & ~n2491;
  assign n2559 = ~n2499 & n2558;
  assign n2560 = ~n595 & ~n664;
  assign n2561 = n595 & n664;
  assign n2562 = ~n2560 & ~n2561;
  assign n2563 = n2491 & ~n2562;
  assign n2564 = ~n2415 & n2563;
  assign n2565 = n2346 & ~n2491;
  assign n2566 = n2418 & n2565;
  assign n2567 = ~n2564 & ~n2566;
  assign n2568 = ~n2559 & n2567;
  assign n2569 = ~n605 & ~n2415;
  assign n2570 = ~n2491 & n2569;
  assign n2571 = ~n2568 & n2570;
  assign n2572 = n2568 & ~n2570;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = n2557 & n2573;
  assign n2575 = ~n2557 & ~n2573;
  assign n2576 = ~n2574 & ~n2575;
  assign n2577 = ~n2545 & n2576;
  assign n2578 = n2545 & ~n2576;
  assign n2579 = ~n2577 & ~n2578;
  assign n2580 = ~n2488 & n2579;
  assign n2581 = n2398 & n2469;
  assign n2582 = n2401 & n2474;
  assign n2583 = n2404 & n2477;
  assign n2584 = n2429 & ~n2431;
  assign n2585 = ~n2432 & ~n2584;
  assign n2586 = n2479 & n2585;
  assign n2587 = ~n2582 & ~n2583;
  assign n2588 = ~n2581 & n2587;
  assign n2589 = ~n2586 & n2588;
  assign n2590 = n869 & n2589;
  assign n2591 = ~n869 & ~n2589;
  assign n2592 = ~n2590 & ~n2591;
  assign n2593 = ~n2541 & ~n2543;
  assign n2594 = ~n2544 & ~n2593;
  assign n2595 = n2592 & n2594;
  assign n2596 = n2401 & n2469;
  assign n2597 = n2404 & n2474;
  assign n2598 = n2407 & n2477;
  assign n2599 = n2425 & ~n2427;
  assign n2600 = ~n2428 & ~n2599;
  assign n2601 = n2479 & n2600;
  assign n2602 = ~n2597 & ~n2598;
  assign n2603 = ~n2596 & n2602;
  assign n2604 = ~n2601 & n2603;
  assign n2605 = n869 & ~n2604;
  assign n2606 = ~n869 & n2604;
  assign n2607 = ~n2605 & ~n2606;
  assign n2608 = n519 & ~n2515;
  assign n2609 = ~n2527 & n2608;
  assign n2610 = n2527 & ~n2608;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = ~n2607 & n2611;
  assign n2613 = n2404 & n2469;
  assign n2614 = n2407 & n2474;
  assign n2615 = n2410 & n2477;
  assign n2616 = n2479 & n2550;
  assign n2617 = ~n2614 & ~n2615;
  assign n2618 = ~n2613 & n2617;
  assign n2619 = ~n2616 & n2618;
  assign n2620 = n869 & n2619;
  assign n2621 = ~n869 & ~n2619;
  assign n2622 = ~n2620 & ~n2621;
  assign n2623 = n519 & n2496;
  assign n2624 = ~n2513 & n2623;
  assign n2625 = n2513 & ~n2623;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = n2622 & n2626;
  assign n2628 = ~n2415 & ~n2465;
  assign n2629 = n2479 & ~n2499;
  assign n2630 = ~n2415 & n2474;
  assign n2631 = n2418 & n2469;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = ~n2629 & n2632;
  assign n2634 = ~n869 & ~n2628;
  assign n2635 = n2633 & n2634;
  assign n2636 = n2410 & n2469;
  assign n2637 = ~n2415 & n2477;
  assign n2638 = n2418 & n2474;
  assign n2639 = n2479 & ~n2523;
  assign n2640 = ~n2637 & ~n2638;
  assign n2641 = ~n2636 & n2640;
  assign n2642 = ~n2639 & n2641;
  assign n2643 = n2635 & n2642;
  assign n2644 = n2496 & n2643;
  assign n2645 = n2407 & n2469;
  assign n2646 = n2418 & n2477;
  assign n2647 = n2410 & n2474;
  assign n2648 = n2479 & n2534;
  assign n2649 = ~n2646 & ~n2647;
  assign n2650 = ~n2645 & n2649;
  assign n2651 = ~n2648 & n2650;
  assign n2652 = ~n869 & n2651;
  assign n2653 = n869 & ~n2651;
  assign n2654 = ~n2652 & ~n2653;
  assign n2655 = ~n2496 & ~n2643;
  assign n2656 = ~n2644 & ~n2655;
  assign n2657 = ~n2654 & n2656;
  assign n2658 = ~n2644 & ~n2657;
  assign n2659 = ~n2622 & ~n2626;
  assign n2660 = ~n2627 & ~n2659;
  assign n2661 = ~n2658 & n2660;
  assign n2662 = ~n2627 & ~n2661;
  assign n2663 = n2607 & ~n2611;
  assign n2664 = ~n2612 & ~n2663;
  assign n2665 = ~n2662 & n2664;
  assign n2666 = ~n2612 & ~n2665;
  assign n2667 = ~n2592 & ~n2594;
  assign n2668 = ~n2595 & ~n2667;
  assign n2669 = ~n2666 & n2668;
  assign n2670 = ~n2595 & ~n2669;
  assign n2671 = n2488 & ~n2579;
  assign n2672 = ~n2580 & ~n2671;
  assign n2673 = ~n2670 & n2672;
  assign n2674 = ~n2580 & ~n2673;
  assign n2675 = ~n2574 & ~n2577;
  assign n2676 = n2401 & n2510;
  assign n2677 = n2404 & n2508;
  assign n2678 = n2407 & n2518;
  assign n2679 = n2503 & n2600;
  assign n2680 = ~n2677 & ~n2678;
  assign n2681 = ~n2676 & n2680;
  assign n2682 = ~n2679 & n2681;
  assign n2683 = n519 & ~n2682;
  assign n2684 = ~n519 & n2682;
  assign n2685 = ~n2683 & ~n2684;
  assign n2686 = ~n605 & ~n2492;
  assign n2687 = n2568 & n2686;
  assign n2688 = ~n605 & ~n2687;
  assign n2689 = n2410 & n2565;
  assign n2690 = n2491 & n2562;
  assign n2691 = ~n2346 & n2690;
  assign n2692 = ~n2415 & n2691;
  assign n2693 = n2418 & n2563;
  assign n2694 = ~n2523 & n2558;
  assign n2695 = ~n2692 & ~n2693;
  assign n2696 = ~n2689 & n2695;
  assign n2697 = ~n2694 & n2696;
  assign n2698 = n2688 & ~n2697;
  assign n2699 = ~n2688 & n2697;
  assign n2700 = ~n2698 & ~n2699;
  assign n2701 = n2685 & n2700;
  assign n2702 = ~n2685 & ~n2700;
  assign n2703 = ~n2701 & ~n2702;
  assign n2704 = n2675 & ~n2703;
  assign n2705 = ~n2675 & n2703;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = n2392 & n2469;
  assign n2708 = n2398 & n2477;
  assign n2709 = n2395 & n2474;
  assign n2710 = n2437 & ~n2439;
  assign n2711 = ~n2440 & ~n2710;
  assign n2712 = n2479 & n2711;
  assign n2713 = ~n2708 & ~n2709;
  assign n2714 = ~n2707 & n2713;
  assign n2715 = ~n2712 & n2714;
  assign n2716 = n869 & n2715;
  assign n2717 = ~n869 & ~n2715;
  assign n2718 = ~n2716 & ~n2717;
  assign n2719 = n2706 & n2718;
  assign n2720 = ~n2706 & ~n2718;
  assign n2721 = ~n2719 & ~n2720;
  assign n2722 = ~n2674 & n2721;
  assign n2723 = n2674 & ~n2721;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = n2462 & n2724;
  assign n2726 = n2375 & n2378;
  assign n2727 = n2387 & n2392;
  assign n2728 = n2382 & n2385;
  assign n2729 = n2445 & ~n2447;
  assign n2730 = ~n2448 & ~n2729;
  assign n2731 = n2389 & n2730;
  assign n2732 = ~n2727 & ~n2728;
  assign n2733 = ~n2726 & n2732;
  assign n2734 = ~n2731 & n2733;
  assign n2735 = ~n57 & n2734;
  assign n2736 = n57 & ~n2734;
  assign n2737 = ~n2735 & ~n2736;
  assign n2738 = n2670 & ~n2672;
  assign n2739 = ~n2673 & ~n2738;
  assign n2740 = n2737 & n2739;
  assign n2741 = n2375 & n2385;
  assign n2742 = n2382 & n2392;
  assign n2743 = n2387 & n2395;
  assign n2744 = n2441 & ~n2443;
  assign n2745 = ~n2444 & ~n2744;
  assign n2746 = n2389 & n2745;
  assign n2747 = ~n2742 & ~n2743;
  assign n2748 = ~n2741 & n2747;
  assign n2749 = ~n2746 & n2748;
  assign n2750 = ~n57 & n2749;
  assign n2751 = n57 & ~n2749;
  assign n2752 = ~n2750 & ~n2751;
  assign n2753 = n2666 & ~n2668;
  assign n2754 = ~n2669 & ~n2753;
  assign n2755 = n2752 & n2754;
  assign n2756 = n2375 & n2392;
  assign n2757 = n2387 & n2398;
  assign n2758 = n2382 & n2395;
  assign n2759 = n2389 & n2711;
  assign n2760 = ~n2757 & ~n2758;
  assign n2761 = ~n2756 & n2760;
  assign n2762 = ~n2759 & n2761;
  assign n2763 = ~n57 & n2762;
  assign n2764 = n57 & ~n2762;
  assign n2765 = ~n2763 & ~n2764;
  assign n2766 = n2662 & ~n2664;
  assign n2767 = ~n2665 & ~n2766;
  assign n2768 = n2765 & n2767;
  assign n2769 = n2375 & n2395;
  assign n2770 = n2382 & n2398;
  assign n2771 = n2387 & n2401;
  assign n2772 = n2389 & n2481;
  assign n2773 = ~n2770 & ~n2771;
  assign n2774 = ~n2769 & n2773;
  assign n2775 = ~n2772 & n2774;
  assign n2776 = n57 & ~n2775;
  assign n2777 = ~n57 & n2775;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = n2658 & ~n2660;
  assign n2780 = ~n2661 & ~n2779;
  assign n2781 = n2778 & n2780;
  assign n2782 = n2375 & n2398;
  assign n2783 = n2382 & n2401;
  assign n2784 = n2387 & n2404;
  assign n2785 = n2389 & n2585;
  assign n2786 = ~n2783 & ~n2784;
  assign n2787 = ~n2782 & n2786;
  assign n2788 = ~n2785 & n2787;
  assign n2789 = ~n57 & n2788;
  assign n2790 = n57 & ~n2788;
  assign n2791 = ~n2789 & ~n2790;
  assign n2792 = n2654 & ~n2656;
  assign n2793 = ~n2657 & ~n2792;
  assign n2794 = n2791 & n2793;
  assign n2795 = n2375 & n2401;
  assign n2796 = n2382 & n2404;
  assign n2797 = n2387 & n2407;
  assign n2798 = n2389 & n2600;
  assign n2799 = ~n2796 & ~n2797;
  assign n2800 = ~n2795 & n2799;
  assign n2801 = ~n2798 & n2800;
  assign n2802 = n57 & ~n2801;
  assign n2803 = ~n57 & n2801;
  assign n2804 = ~n2802 & ~n2803;
  assign n2805 = ~n869 & ~n2635;
  assign n2806 = ~n2642 & n2805;
  assign n2807 = n2642 & ~n2805;
  assign n2808 = ~n2806 & ~n2807;
  assign n2809 = n2804 & n2808;
  assign n2810 = n2375 & n2404;
  assign n2811 = n2382 & n2407;
  assign n2812 = n2387 & n2410;
  assign n2813 = n2389 & n2550;
  assign n2814 = ~n2811 & ~n2812;
  assign n2815 = ~n2810 & n2814;
  assign n2816 = ~n2813 & n2815;
  assign n2817 = ~n57 & n2816;
  assign n2818 = n57 & ~n2816;
  assign n2819 = ~n2817 & ~n2818;
  assign n2820 = ~n869 & n2628;
  assign n2821 = ~n2633 & n2820;
  assign n2822 = n2633 & ~n2820;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = n2819 & n2823;
  assign n2825 = ~n2371 & ~n2415;
  assign n2826 = n2389 & ~n2499;
  assign n2827 = n2382 & ~n2415;
  assign n2828 = n2375 & n2418;
  assign n2829 = ~n2827 & ~n2828;
  assign n2830 = ~n2826 & n2829;
  assign n2831 = n57 & ~n2825;
  assign n2832 = n2830 & n2831;
  assign n2833 = n2375 & n2410;
  assign n2834 = n2387 & ~n2415;
  assign n2835 = n2382 & n2418;
  assign n2836 = n2389 & ~n2523;
  assign n2837 = ~n2834 & ~n2835;
  assign n2838 = ~n2833 & n2837;
  assign n2839 = ~n2836 & n2838;
  assign n2840 = n2832 & n2839;
  assign n2841 = n2628 & n2840;
  assign n2842 = n2375 & n2407;
  assign n2843 = n2387 & n2418;
  assign n2844 = n2382 & n2410;
  assign n2845 = n2389 & n2534;
  assign n2846 = ~n2843 & ~n2844;
  assign n2847 = ~n2842 & n2846;
  assign n2848 = ~n2845 & n2847;
  assign n2849 = n57 & ~n2848;
  assign n2850 = ~n57 & n2848;
  assign n2851 = ~n2849 & ~n2850;
  assign n2852 = ~n2628 & ~n2840;
  assign n2853 = ~n2841 & ~n2852;
  assign n2854 = n2851 & n2853;
  assign n2855 = ~n2841 & ~n2854;
  assign n2856 = ~n2819 & ~n2823;
  assign n2857 = ~n2824 & ~n2856;
  assign n2858 = ~n2855 & n2857;
  assign n2859 = ~n2824 & ~n2858;
  assign n2860 = ~n2804 & ~n2808;
  assign n2861 = ~n2809 & ~n2860;
  assign n2862 = ~n2859 & n2861;
  assign n2863 = ~n2809 & ~n2862;
  assign n2864 = ~n2791 & ~n2793;
  assign n2865 = ~n2794 & ~n2864;
  assign n2866 = ~n2863 & n2865;
  assign n2867 = ~n2794 & ~n2866;
  assign n2868 = ~n2778 & ~n2780;
  assign n2869 = ~n2781 & ~n2868;
  assign n2870 = ~n2867 & n2869;
  assign n2871 = ~n2781 & ~n2870;
  assign n2872 = ~n2765 & ~n2767;
  assign n2873 = ~n2768 & ~n2872;
  assign n2874 = ~n2871 & n2873;
  assign n2875 = ~n2768 & ~n2874;
  assign n2876 = ~n2752 & ~n2754;
  assign n2877 = ~n2755 & ~n2876;
  assign n2878 = ~n2875 & n2877;
  assign n2879 = ~n2755 & ~n2878;
  assign n2880 = ~n2737 & ~n2739;
  assign n2881 = ~n2740 & ~n2880;
  assign n2882 = ~n2879 & n2881;
  assign n2883 = ~n2740 & ~n2882;
  assign n2884 = ~n2462 & ~n2724;
  assign n2885 = ~n2725 & ~n2884;
  assign n2886 = ~n2883 & n2885;
  assign n2887 = ~n2725 & ~n2886;
  assign n2888 = ~n2359 & ~n2362;
  assign n2889 = ~n119 & ~n223;
  assign n2890 = ~n247 & ~n314;
  assign n2891 = ~n384 & n2890;
  assign n2892 = n2889 & n2891;
  assign n2893 = n286 & n2892;
  assign n2894 = ~n272 & ~n378;
  assign n2895 = n346 & n565;
  assign n2896 = n794 & n993;
  assign n2897 = n2894 & n2896;
  assign n2898 = n967 & n2895;
  assign n2899 = n2897 & n2898;
  assign n2900 = n611 & n2899;
  assign n2901 = n2131 & n2893;
  assign n2902 = n2900 & n2901;
  assign n2903 = n1306 & n2902;
  assign n2904 = n2888 & n2903;
  assign n2905 = ~n2888 & ~n2903;
  assign n2906 = ~n2904 & ~n2905;
  assign n2907 = n2375 & ~n2906;
  assign n2908 = n2378 & n2387;
  assign n2909 = n2364 & n2382;
  assign n2910 = ~n2450 & ~n2453;
  assign n2911 = n2364 & ~n2906;
  assign n2912 = ~n2364 & n2906;
  assign n2913 = ~n2911 & ~n2912;
  assign n2914 = ~n2910 & n2913;
  assign n2915 = n2910 & ~n2913;
  assign n2916 = ~n2914 & ~n2915;
  assign n2917 = n2389 & n2916;
  assign n2918 = ~n2908 & ~n2909;
  assign n2919 = ~n2907 & n2918;
  assign n2920 = ~n2917 & n2919;
  assign n2921 = n57 & ~n2920;
  assign n2922 = ~n57 & n2920;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = ~n2719 & ~n2722;
  assign n2925 = ~n2701 & ~n2705;
  assign n2926 = n2398 & n2510;
  assign n2927 = n2401 & n2508;
  assign n2928 = n2404 & n2518;
  assign n2929 = n2503 & n2585;
  assign n2930 = ~n2927 & ~n2928;
  assign n2931 = ~n2926 & n2930;
  assign n2932 = ~n2929 & n2931;
  assign n2933 = n519 & ~n2932;
  assign n2934 = ~n519 & n2932;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = n2407 & n2565;
  assign n2937 = n2418 & n2691;
  assign n2938 = n2410 & n2563;
  assign n2939 = n2534 & n2558;
  assign n2940 = ~n2937 & ~n2938;
  assign n2941 = ~n2936 & n2940;
  assign n2942 = ~n2939 & n2941;
  assign n2943 = n605 & ~n2942;
  assign n2944 = ~n605 & n2942;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = n2687 & n2697;
  assign n2947 = ~n2569 & ~n2946;
  assign n2948 = n2569 & n2946;
  assign n2949 = ~n2947 & ~n2948;
  assign n2950 = ~n2945 & n2949;
  assign n2951 = n2945 & ~n2949;
  assign n2952 = ~n2950 & ~n2951;
  assign n2953 = n2935 & n2952;
  assign n2954 = ~n2935 & ~n2952;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = n2925 & ~n2955;
  assign n2957 = ~n2925 & n2955;
  assign n2958 = ~n2956 & ~n2957;
  assign n2959 = n2385 & n2469;
  assign n2960 = n2392 & n2474;
  assign n2961 = n2395 & n2477;
  assign n2962 = n2479 & n2745;
  assign n2963 = ~n2960 & ~n2961;
  assign n2964 = ~n2959 & n2963;
  assign n2965 = ~n2962 & n2964;
  assign n2966 = n869 & n2965;
  assign n2967 = ~n869 & ~n2965;
  assign n2968 = ~n2966 & ~n2967;
  assign n2969 = n2958 & n2968;
  assign n2970 = ~n2958 & ~n2968;
  assign n2971 = ~n2969 & ~n2970;
  assign n2972 = ~n2924 & n2971;
  assign n2973 = n2924 & ~n2971;
  assign n2974 = ~n2972 & ~n2973;
  assign n2975 = n2923 & n2974;
  assign n2976 = ~n2923 & ~n2974;
  assign n2977 = ~n2975 & ~n2976;
  assign n2978 = n2887 & ~n2977;
  assign n2979 = ~n2887 & n2977;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = ~n209 & ~n457;
  assign n2982 = ~n461 & n2981;
  assign n2983 = ~n520 & ~n564;
  assign n2984 = ~n186 & ~n404;
  assign n2985 = ~n181 & ~n325;
  assign n2986 = ~n355 & n2985;
  assign n2987 = n2275 & n2986;
  assign n2988 = ~n174 & ~n310;
  assign n2989 = n305 & n2988;
  assign n2990 = ~n218 & ~n237;
  assign n2991 = ~n264 & ~n294;
  assign n2992 = ~n299 & ~n548;
  assign n2993 = n2991 & n2992;
  assign n2994 = n2983 & n2990;
  assign n2995 = n2984 & n2994;
  assign n2996 = n1989 & n2993;
  assign n2997 = n2989 & n2996;
  assign n2998 = n2987 & n2995;
  assign n2999 = n2997 & n2998;
  assign n3000 = ~n273 & ~n329;
  assign n3001 = ~n268 & ~n298;
  assign n3002 = ~n314 & ~n433;
  assign n3003 = ~n530 & ~n552;
  assign n3004 = n3002 & n3003;
  assign n3005 = n409 & n3001;
  assign n3006 = n3000 & n3005;
  assign n3007 = n2147 & n3004;
  assign n3008 = n2982 & n3007;
  assign n3009 = n206 & n3006;
  assign n3010 = n3008 & n3009;
  assign n3011 = n169 & n3010;
  assign n3012 = n2999 & n3011;
  assign n3013 = n2904 & n3012;
  assign n3014 = ~n108 & ~n207;
  assign n3015 = ~n210 & ~n248;
  assign n3016 = n1003 & n3015;
  assign n3017 = n344 & n3014;
  assign n3018 = n814 & n2217;
  assign n3019 = n3017 & n3018;
  assign n3020 = n3016 & n3019;
  assign n3021 = n2025 & n2123;
  assign n3022 = n3020 & n3021;
  assign n3023 = n571 & n3022;
  assign n3024 = n498 & n3023;
  assign n3025 = n3013 & n3024;
  assign n3026 = ~n250 & ~n282;
  assign n3027 = n455 & n549;
  assign n3028 = n3026 & n3027;
  assign n3029 = n460 & n472;
  assign n3030 = n1012 & n3029;
  assign n3031 = n542 & n3028;
  assign n3032 = n3030 & n3031;
  assign n3033 = n490 & n527;
  assign n3034 = n571 & n3033;
  assign n3035 = n3032 & n3034;
  assign n3036 = n3025 & n3035;
  assign n3037 = ~n3025 & ~n3035;
  assign n3038 = ~n3036 & ~n3037;
  assign n3039 = pi0  & ~pi22 ;
  assign n3040 = pi1  & ~n3039;
  assign n3041 = ~pi1  & n3039;
  assign n3042 = ~n3040 & ~n3041;
  assign n3043 = n2368 & n3042;
  assign n3044 = ~n2368 & ~n3042;
  assign n3045 = ~n3043 & ~n3044;
  assign n3046 = pi0  & ~n3045;
  assign n3047 = ~n3038 & n3046;
  assign n3048 = ~n3013 & ~n3024;
  assign n3049 = ~n3025 & ~n3048;
  assign n3050 = ~pi0  & ~n3042;
  assign n3051 = ~n3049 & n3050;
  assign n3052 = ~n2904 & ~n3012;
  assign n3053 = ~n3013 & ~n3052;
  assign n3054 = pi2  & n50;
  assign n3055 = ~n3053 & n3054;
  assign n3056 = pi0  & n3045;
  assign n3057 = ~n3049 & ~n3053;
  assign n3058 = ~n2906 & ~n3053;
  assign n3059 = ~n2911 & ~n2914;
  assign n3060 = n2906 & n3012;
  assign n3061 = ~n3058 & ~n3060;
  assign n3062 = ~n3059 & n3061;
  assign n3063 = ~n3058 & ~n3062;
  assign n3064 = n3024 & n3053;
  assign n3065 = ~n3057 & ~n3064;
  assign n3066 = ~n3063 & n3065;
  assign n3067 = ~n3057 & ~n3066;
  assign n3068 = ~n3038 & ~n3049;
  assign n3069 = n3035 & n3049;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = ~n3067 & n3070;
  assign n3072 = n3067 & ~n3070;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = n3056 & n3073;
  assign n3075 = ~n3051 & ~n3055;
  assign n3076 = ~n3047 & n3075;
  assign n3077 = ~n3074 & n3076;
  assign n3078 = n2368 & n3077;
  assign n3079 = ~n2368 & ~n3077;
  assign n3080 = ~n3078 & ~n3079;
  assign n3081 = n2980 & n3080;
  assign n3082 = n2883 & ~n2885;
  assign n3083 = ~n2886 & ~n3082;
  assign n3084 = n3046 & ~n3049;
  assign n3085 = n3050 & ~n3053;
  assign n3086 = ~n2906 & n3054;
  assign n3087 = n3063 & ~n3065;
  assign n3088 = ~n3066 & ~n3087;
  assign n3089 = n3056 & n3088;
  assign n3090 = ~n3085 & ~n3086;
  assign n3091 = ~n3084 & n3090;
  assign n3092 = ~n3089 & n3091;
  assign n3093 = n2368 & n3092;
  assign n3094 = ~n2368 & ~n3092;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = n3083 & n3095;
  assign n3097 = ~n3083 & ~n3095;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = n2879 & ~n2881;
  assign n3100 = ~n2882 & ~n3099;
  assign n3101 = n2875 & ~n2877;
  assign n3102 = ~n2878 & ~n3101;
  assign n3103 = n2871 & ~n2873;
  assign n3104 = ~n2874 & ~n3103;
  assign n3105 = n2867 & ~n2869;
  assign n3106 = ~n2870 & ~n3105;
  assign n3107 = n2863 & ~n2865;
  assign n3108 = ~n2866 & ~n3107;
  assign n3109 = n2859 & ~n2861;
  assign n3110 = ~n2862 & ~n3109;
  assign n3111 = n2855 & ~n2857;
  assign n3112 = ~n2858 & ~n3111;
  assign n3113 = n2398 & n3046;
  assign n3114 = n2401 & n3050;
  assign n3115 = n2404 & n3054;
  assign n3116 = n2585 & n3056;
  assign n3117 = ~n3114 & ~n3115;
  assign n3118 = ~n3113 & n3117;
  assign n3119 = ~n3116 & n3118;
  assign n3120 = n2368 & ~n3119;
  assign n3121 = ~n2368 & n3119;
  assign n3122 = ~n3120 & ~n3121;
  assign n3123 = n57 & ~n2832;
  assign n3124 = ~n2839 & n3123;
  assign n3125 = n2839 & ~n3123;
  assign n3126 = ~n3124 & ~n3125;
  assign n3127 = n57 & n2825;
  assign n3128 = ~n2830 & n3127;
  assign n3129 = n2830 & ~n3127;
  assign n3130 = ~n3128 & ~n3129;
  assign n3131 = n2418 & n3050;
  assign n3132 = ~n2410 & n2499;
  assign n3133 = n3056 & ~n3132;
  assign n3134 = ~n2410 & ~n2418;
  assign n3135 = n3046 & ~n3134;
  assign n3136 = ~n51 & ~n2415;
  assign n3137 = ~n2368 & ~n3136;
  assign n3138 = ~n3131 & n3137;
  assign n3139 = ~n3133 & n3138;
  assign n3140 = ~n3135 & n3139;
  assign n3141 = n2825 & n3140;
  assign n3142 = ~n2825 & ~n3140;
  assign n3143 = n2407 & n3046;
  assign n3144 = n2410 & n3050;
  assign n3145 = n2534 & n3056;
  assign n3146 = ~n3143 & ~n3144;
  assign n3147 = ~n3145 & n3146;
  assign n3148 = n2368 & ~n3147;
  assign n3149 = n2418 & n3054;
  assign n3150 = ~n2368 & ~n3149;
  assign n3151 = n3147 & n3150;
  assign n3152 = ~n3148 & ~n3151;
  assign n3153 = ~n3142 & ~n3152;
  assign n3154 = ~n3141 & ~n3153;
  assign n3155 = n3130 & ~n3154;
  assign n3156 = ~n3130 & n3154;
  assign n3157 = n2404 & n3046;
  assign n3158 = n2407 & n3050;
  assign n3159 = n2410 & n3054;
  assign n3160 = n2550 & n3056;
  assign n3161 = ~n3158 & ~n3159;
  assign n3162 = ~n3157 & n3161;
  assign n3163 = ~n3160 & n3162;
  assign n3164 = ~n2368 & ~n3163;
  assign n3165 = n2368 & n3163;
  assign n3166 = ~n3164 & ~n3165;
  assign n3167 = ~n3156 & n3166;
  assign n3168 = ~n3155 & ~n3167;
  assign n3169 = ~n3126 & n3168;
  assign n3170 = n3126 & ~n3168;
  assign n3171 = n2401 & n3046;
  assign n3172 = n2404 & n3050;
  assign n3173 = n2407 & n3054;
  assign n3174 = n2600 & n3056;
  assign n3175 = ~n3172 & ~n3173;
  assign n3176 = ~n3171 & n3175;
  assign n3177 = ~n3174 & n3176;
  assign n3178 = n2368 & ~n3177;
  assign n3179 = ~n2368 & n3177;
  assign n3180 = ~n3178 & ~n3179;
  assign n3181 = ~n3170 & n3180;
  assign n3182 = ~n3169 & ~n3181;
  assign n3183 = ~n3122 & n3182;
  assign n3184 = n3122 & ~n3182;
  assign n3185 = ~n2851 & ~n2853;
  assign n3186 = ~n2854 & ~n3185;
  assign n3187 = ~n3184 & n3186;
  assign n3188 = ~n3183 & ~n3187;
  assign n3189 = ~n3112 & n3188;
  assign n3190 = n3112 & ~n3188;
  assign n3191 = n2395 & n3046;
  assign n3192 = n2398 & n3050;
  assign n3193 = n2401 & n3054;
  assign n3194 = n2481 & n3056;
  assign n3195 = ~n3192 & ~n3193;
  assign n3196 = ~n3191 & n3195;
  assign n3197 = ~n3194 & n3196;
  assign n3198 = n2368 & ~n3197;
  assign n3199 = ~n2368 & n3197;
  assign n3200 = ~n3198 & ~n3199;
  assign n3201 = ~n3190 & n3200;
  assign n3202 = ~n3189 & ~n3201;
  assign n3203 = n3110 & n3202;
  assign n3204 = ~n3110 & ~n3202;
  assign n3205 = n2392 & n3046;
  assign n3206 = n2395 & n3050;
  assign n3207 = n2711 & n3056;
  assign n3208 = ~n3205 & ~n3206;
  assign n3209 = ~n3207 & n3208;
  assign n3210 = n2368 & ~n3209;
  assign n3211 = n50 & n2398;
  assign n3212 = ~n2368 & ~n3211;
  assign n3213 = n3209 & n3212;
  assign n3214 = ~n3210 & ~n3213;
  assign n3215 = ~n3204 & ~n3214;
  assign n3216 = ~n3203 & ~n3215;
  assign n3217 = n3108 & ~n3216;
  assign n3218 = ~n3108 & n3216;
  assign n3219 = n2385 & n3046;
  assign n3220 = n2392 & n3050;
  assign n3221 = n2395 & n3054;
  assign n3222 = n2745 & n3056;
  assign n3223 = ~n3220 & ~n3221;
  assign n3224 = ~n3219 & n3223;
  assign n3225 = ~n3222 & n3224;
  assign n3226 = ~n2368 & ~n3225;
  assign n3227 = n2368 & n3225;
  assign n3228 = ~n3226 & ~n3227;
  assign n3229 = ~n3218 & n3228;
  assign n3230 = ~n3217 & ~n3229;
  assign n3231 = n3106 & ~n3230;
  assign n3232 = ~n3106 & n3230;
  assign n3233 = n2378 & n3046;
  assign n3234 = n2385 & n3050;
  assign n3235 = n2730 & n3056;
  assign n3236 = ~n3233 & ~n3234;
  assign n3237 = ~n3235 & n3236;
  assign n3238 = n2368 & ~n3237;
  assign n3239 = n50 & n2392;
  assign n3240 = ~n2368 & ~n3239;
  assign n3241 = n3237 & n3240;
  assign n3242 = ~n3238 & ~n3241;
  assign n3243 = ~n3232 & ~n3242;
  assign n3244 = ~n3231 & ~n3243;
  assign n3245 = ~n3104 & n3244;
  assign n3246 = n3104 & ~n3244;
  assign n3247 = n2364 & n3046;
  assign n3248 = n2378 & n3050;
  assign n3249 = n2385 & n3054;
  assign n3250 = n2455 & n3056;
  assign n3251 = ~n3248 & ~n3249;
  assign n3252 = ~n3247 & n3251;
  assign n3253 = ~n3250 & n3252;
  assign n3254 = n2368 & ~n3253;
  assign n3255 = ~n2368 & n3253;
  assign n3256 = ~n3254 & ~n3255;
  assign n3257 = ~n3246 & n3256;
  assign n3258 = ~n3245 & ~n3257;
  assign n3259 = n3102 & n3258;
  assign n3260 = ~n3102 & ~n3258;
  assign n3261 = ~n2906 & n3046;
  assign n3262 = n2364 & n3050;
  assign n3263 = n2916 & n3056;
  assign n3264 = ~n3261 & ~n3262;
  assign n3265 = ~n3263 & n3264;
  assign n3266 = n2368 & ~n3265;
  assign n3267 = n50 & n2378;
  assign n3268 = ~n2368 & ~n3267;
  assign n3269 = n3265 & n3268;
  assign n3270 = ~n3266 & ~n3269;
  assign n3271 = ~n3260 & ~n3270;
  assign n3272 = ~n3259 & ~n3271;
  assign n3273 = ~n3100 & n3272;
  assign n3274 = n3100 & ~n3272;
  assign n3275 = n3046 & ~n3053;
  assign n3276 = ~n2906 & n3050;
  assign n3277 = n2364 & n3054;
  assign n3278 = n3059 & ~n3061;
  assign n3279 = ~n3062 & ~n3278;
  assign n3280 = n3056 & n3279;
  assign n3281 = ~n3276 & ~n3277;
  assign n3282 = ~n3275 & n3281;
  assign n3283 = ~n3280 & n3282;
  assign n3284 = n2368 & ~n3283;
  assign n3285 = ~n2368 & n3283;
  assign n3286 = ~n3284 & ~n3285;
  assign n3287 = ~n3274 & n3286;
  assign n3288 = ~n3273 & ~n3287;
  assign n3289 = n3098 & n3288;
  assign n3290 = ~n3096 & ~n3289;
  assign n3291 = ~n2980 & ~n3080;
  assign n3292 = ~n3081 & ~n3291;
  assign n3293 = ~n3290 & n3292;
  assign n3294 = ~n3081 & ~n3293;
  assign n3295 = ~n2975 & ~n2979;
  assign n3296 = n2375 & ~n3053;
  assign n3297 = n2382 & ~n2906;
  assign n3298 = n2364 & n2387;
  assign n3299 = n2389 & n3279;
  assign n3300 = ~n3297 & ~n3298;
  assign n3301 = ~n3296 & n3300;
  assign n3302 = ~n3299 & n3301;
  assign n3303 = n57 & ~n3302;
  assign n3304 = ~n57 & n3302;
  assign n3305 = ~n3303 & ~n3304;
  assign n3306 = ~n2969 & ~n2972;
  assign n3307 = n2378 & n2469;
  assign n3308 = n2392 & n2477;
  assign n3309 = n2385 & n2474;
  assign n3310 = n2479 & n2730;
  assign n3311 = ~n3308 & ~n3309;
  assign n3312 = ~n3307 & n3311;
  assign n3313 = ~n3310 & n3312;
  assign n3314 = n869 & n3313;
  assign n3315 = ~n869 & ~n3313;
  assign n3316 = ~n3314 & ~n3315;
  assign n3317 = ~n2953 & ~n2957;
  assign n3318 = n2395 & n2510;
  assign n3319 = n2398 & n2508;
  assign n3320 = n2401 & n2518;
  assign n3321 = n2481 & n2503;
  assign n3322 = ~n3319 & ~n3320;
  assign n3323 = ~n3318 & n3322;
  assign n3324 = ~n3321 & n3323;
  assign n3325 = n519 & ~n3324;
  assign n3326 = ~n519 & n3324;
  assign n3327 = ~n3325 & ~n3326;
  assign n3328 = ~n2948 & ~n2950;
  assign n3329 = ~n605 & ~n2418;
  assign n3330 = n2404 & n2565;
  assign n3331 = n2407 & n2563;
  assign n3332 = n2410 & n2691;
  assign n3333 = n2550 & n2558;
  assign n3334 = ~n3331 & ~n3332;
  assign n3335 = ~n3330 & n3334;
  assign n3336 = ~n3333 & n3335;
  assign n3337 = n3329 & ~n3336;
  assign n3338 = ~n3329 & n3336;
  assign n3339 = ~n3337 & ~n3338;
  assign n3340 = ~n3328 & n3339;
  assign n3341 = n3328 & ~n3339;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = n3327 & n3342;
  assign n3344 = ~n3327 & ~n3342;
  assign n3345 = ~n3343 & ~n3344;
  assign n3346 = ~n3317 & n3345;
  assign n3347 = n3317 & ~n3345;
  assign n3348 = ~n3346 & ~n3347;
  assign n3349 = n3316 & n3348;
  assign n3350 = ~n3316 & ~n3348;
  assign n3351 = ~n3349 & ~n3350;
  assign n3352 = ~n3306 & n3351;
  assign n3353 = n3306 & ~n3351;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355 = n3305 & n3354;
  assign n3356 = ~n3305 & ~n3354;
  assign n3357 = ~n3355 & ~n3356;
  assign n3358 = ~n3295 & n3357;
  assign n3359 = n3295 & ~n3357;
  assign n3360 = ~n3358 & ~n3359;
  assign n3361 = ~n153 & n528;
  assign n3362 = n115 & n118;
  assign n3363 = ~n543 & ~n3362;
  assign n3364 = n468 & n3363;
  assign n3365 = n480 & n537;
  assign n3366 = n571 & n3365;
  assign n3367 = n3364 & n3366;
  assign n3368 = n3361 & n3367;
  assign n3369 = ~n3036 & ~n3368;
  assign n3370 = n3036 & n3368;
  assign n3371 = ~n3369 & ~n3370;
  assign n3372 = n3046 & ~n3371;
  assign n3373 = ~n3038 & n3050;
  assign n3374 = ~n3049 & n3054;
  assign n3375 = ~n3068 & ~n3071;
  assign n3376 = ~n3038 & ~n3371;
  assign n3377 = n3038 & n3368;
  assign n3378 = ~n3376 & ~n3377;
  assign n3379 = ~n3375 & n3378;
  assign n3380 = n3375 & ~n3378;
  assign n3381 = ~n3379 & ~n3380;
  assign n3382 = n3056 & n3381;
  assign n3383 = ~n3373 & ~n3374;
  assign n3384 = ~n3372 & n3383;
  assign n3385 = ~n3382 & n3384;
  assign n3386 = n2368 & n3385;
  assign n3387 = ~n2368 & ~n3385;
  assign n3388 = ~n3386 & ~n3387;
  assign n3389 = n3360 & n3388;
  assign n3390 = ~n3360 & ~n3388;
  assign n3391 = ~n3389 & ~n3390;
  assign n3392 = ~n3294 & n3391;
  assign n3393 = n3294 & ~n3391;
  assign n3394 = ~n3392 & ~n3393;
  assign n3395 = ~n192 & ~n225;
  assign n3396 = n483 & n3395;
  assign n3397 = n390 & n3396;
  assign n3398 = n2987 & n3397;
  assign n3399 = ~n108 & ~n548;
  assign n3400 = ~n185 & ~n248;
  assign n3401 = ~n171 & ~n272;
  assign n3402 = ~n314 & ~n543;
  assign n3403 = n3401 & n3402;
  assign n3404 = n2185 & n3403;
  assign n3405 = ~n140 & ~n148;
  assign n3406 = ~n219 & ~n222;
  assign n3407 = ~n433 & ~n454;
  assign n3408 = n3406 & n3407;
  assign n3409 = n398 & n3405;
  assign n3410 = n2033 & n3400;
  assign n3411 = n3409 & n3410;
  assign n3412 = n3408 & n3411;
  assign n3413 = n3404 & n3412;
  assign n3414 = ~n137 & ~n249;
  assign n3415 = n3399 & n3414;
  assign n3416 = n3413 & n3415;
  assign n3417 = ~n190 & ~n263;
  assign n3418 = ~n267 & ~n307;
  assign n3419 = ~n356 & n3418;
  assign n3420 = n606 & n3417;
  assign n3421 = n2326 & n2984;
  assign n3422 = n3420 & n3421;
  assign n3423 = n2982 & n3419;
  assign n3424 = n3422 & n3423;
  assign n3425 = n421 & n3424;
  assign n3426 = n3398 & n3425;
  assign n3427 = n3416 & n3426;
  assign n3428 = n3394 & ~n3427;
  assign n3429 = ~n3394 & n3427;
  assign n3430 = ~n3428 & ~n3429;
  assign n3431 = n3290 & ~n3292;
  assign n3432 = ~n3293 & ~n3431;
  assign n3433 = ~n188 & ~n198;
  assign n3434 = ~n295 & ~n317;
  assign n3435 = ~n404 & n3434;
  assign n3436 = n3433 & n3435;
  assign n3437 = ~n129 & ~n208;
  assign n3438 = ~n224 & ~n233;
  assign n3439 = n3437 & n3438;
  assign n3440 = n281 & n297;
  assign n3441 = n3000 & n3440;
  assign n3442 = n3439 & n3441;
  assign n3443 = n3436 & n3442;
  assign n3444 = ~n134 & ~n140;
  assign n3445 = ~n235 & ~n370;
  assign n3446 = ~n481 & n3445;
  assign n3447 = n330 & n3444;
  assign n3448 = n2126 & n3447;
  assign n3449 = n2158 & n3446;
  assign n3450 = n3448 & n3449;
  assign n3451 = n1017 & n3450;
  assign n3452 = ~n145 & ~n279;
  assign n3453 = n302 & n3452;
  assign n3454 = n3451 & n3453;
  assign n3455 = ~n176 & ~n210;
  assign n3456 = ~n226 & ~n239;
  assign n3457 = ~n345 & n3456;
  assign n3458 = n827 & n3455;
  assign n3459 = n848 & n2983;
  assign n3460 = n3458 & n3459;
  assign n3461 = n3457 & n3460;
  assign n3462 = n2249 & n3461;
  assign n3463 = n3443 & n3462;
  assign n3464 = n3454 & n3463;
  assign n3465 = ~n3432 & n3464;
  assign n3466 = n3432 & ~n3464;
  assign n3467 = ~n298 & ~n304;
  assign n3468 = n1290 & n3467;
  assign n3469 = n459 & n3468;
  assign n3470 = n2070 & n3469;
  assign n3471 = n2103 & n3470;
  assign n3472 = ~n239 & ~n324;
  assign n3473 = n351 & n3472;
  assign n3474 = n2333 & n3473;
  assign n3475 = ~n148 & ~n218;
  assign n3476 = ~n222 & ~n251;
  assign n3477 = ~n315 & ~n329;
  assign n3478 = ~n384 & n3477;
  assign n3479 = n3475 & n3476;
  assign n3480 = n550 & n629;
  assign n3481 = n2213 & n2216;
  assign n3482 = n3480 & n3481;
  assign n3483 = n3478 & n3479;
  assign n3484 = n3482 & n3483;
  assign n3485 = n2172 & n3484;
  assign n3486 = n3471 & n3485;
  assign n3487 = n3474 & n3486;
  assign n3488 = ~n3098 & ~n3288;
  assign n3489 = ~n3289 & ~n3487;
  assign n3490 = ~n3488 & n3489;
  assign n3491 = ~n3466 & ~n3490;
  assign n3492 = ~n3465 & ~n3491;
  assign n3493 = n3430 & n3492;
  assign n3494 = ~n3428 & ~n3493;
  assign n3495 = ~n3389 & ~n3392;
  assign n3496 = ~n152 & ~n190;
  assign n3497 = ~n403 & ~n457;
  assign n3498 = n3496 & n3497;
  assign n3499 = n426 & n2047;
  assign n3500 = n3400 & n3499;
  assign n3501 = n3498 & n3500;
  assign n3502 = ~n137 & ~n139;
  assign n3503 = ~n144 & ~n148;
  assign n3504 = ~n219 & ~n315;
  assign n3505 = ~n576 & n3504;
  assign n3506 = n3502 & n3503;
  assign n3507 = n2217 & n2894;
  assign n3508 = n3506 & n3507;
  assign n3509 = n401 & n3505;
  assign n3510 = n3508 & n3509;
  assign n3511 = n2330 & n3510;
  assign n3512 = n3501 & n3511;
  assign n3513 = n1009 & n3512;
  assign n3514 = n3370 & n3513;
  assign n3515 = ~n3370 & ~n3513;
  assign n3516 = ~n3514 & ~n3515;
  assign n3517 = n3046 & ~n3516;
  assign n3518 = n3050 & ~n3371;
  assign n3519 = ~n3038 & n3054;
  assign n3520 = ~n3376 & ~n3379;
  assign n3521 = ~n3371 & ~n3516;
  assign n3522 = n3371 & n3513;
  assign n3523 = ~n3521 & ~n3522;
  assign n3524 = ~n3520 & n3523;
  assign n3525 = n3520 & ~n3523;
  assign n3526 = ~n3524 & ~n3525;
  assign n3527 = n3056 & n3526;
  assign n3528 = ~n3518 & ~n3519;
  assign n3529 = ~n3517 & n3528;
  assign n3530 = ~n3527 & n3529;
  assign n3531 = n2368 & ~n3530;
  assign n3532 = ~n2368 & n3530;
  assign n3533 = ~n3531 & ~n3532;
  assign n3534 = ~n3355 & ~n3358;
  assign n3535 = ~n3349 & ~n3352;
  assign n3536 = n2364 & n2469;
  assign n3537 = n2378 & n2474;
  assign n3538 = n2385 & n2477;
  assign n3539 = n2455 & n2479;
  assign n3540 = ~n3537 & ~n3538;
  assign n3541 = ~n3536 & n3540;
  assign n3542 = ~n3539 & n3541;
  assign n3543 = n869 & ~n3542;
  assign n3544 = ~n869 & n3542;
  assign n3545 = ~n3543 & ~n3544;
  assign n3546 = ~n3343 & ~n3346;
  assign n3547 = ~n605 & ~n2410;
  assign n3548 = n2401 & n2565;
  assign n3549 = n2404 & n2563;
  assign n3550 = n2407 & n2691;
  assign n3551 = n2558 & n2600;
  assign n3552 = ~n3549 & ~n3550;
  assign n3553 = ~n3548 & n3552;
  assign n3554 = ~n3551 & n3553;
  assign n3555 = n3547 & ~n3554;
  assign n3556 = ~n3547 & n3554;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = ~n605 & n2418;
  assign n3559 = n3336 & n3558;
  assign n3560 = ~n3340 & ~n3559;
  assign n3561 = n3557 & ~n3560;
  assign n3562 = ~n3557 & n3560;
  assign n3563 = ~n3561 & ~n3562;
  assign n3564 = n2392 & n2510;
  assign n3565 = n2398 & n2518;
  assign n3566 = n2395 & n2508;
  assign n3567 = n2503 & n2711;
  assign n3568 = ~n3565 & ~n3566;
  assign n3569 = ~n3564 & n3568;
  assign n3570 = ~n3567 & n3569;
  assign n3571 = ~n519 & n3570;
  assign n3572 = n519 & ~n3570;
  assign n3573 = ~n3571 & ~n3572;
  assign n3574 = n3563 & n3573;
  assign n3575 = ~n3563 & ~n3573;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = ~n3546 & n3576;
  assign n3578 = n3546 & ~n3576;
  assign n3579 = ~n3577 & ~n3578;
  assign n3580 = ~n3545 & n3579;
  assign n3581 = n3545 & ~n3579;
  assign n3582 = ~n3580 & ~n3581;
  assign n3583 = n3535 & ~n3582;
  assign n3584 = ~n3535 & n3582;
  assign n3585 = ~n3583 & ~n3584;
  assign n3586 = n2375 & ~n3049;
  assign n3587 = n2382 & ~n3053;
  assign n3588 = n2387 & ~n2906;
  assign n3589 = n2389 & n3088;
  assign n3590 = ~n3587 & ~n3588;
  assign n3591 = ~n3586 & n3590;
  assign n3592 = ~n3589 & n3591;
  assign n3593 = ~n57 & n3592;
  assign n3594 = n57 & ~n3592;
  assign n3595 = ~n3593 & ~n3594;
  assign n3596 = n3585 & n3595;
  assign n3597 = ~n3585 & ~n3595;
  assign n3598 = ~n3596 & ~n3597;
  assign n3599 = ~n3534 & n3598;
  assign n3600 = n3534 & ~n3598;
  assign n3601 = ~n3599 & ~n3600;
  assign n3602 = ~n3533 & n3601;
  assign n3603 = n3533 & ~n3601;
  assign n3604 = ~n3602 & ~n3603;
  assign n3605 = n3495 & ~n3604;
  assign n3606 = ~n3495 & n3604;
  assign n3607 = ~n3605 & ~n3606;
  assign n3608 = ~n149 & ~n220;
  assign n3609 = ~n481 & n3608;
  assign n3610 = n297 & n3400;
  assign n3611 = n3609 & n3610;
  assign n3612 = n965 & n1297;
  assign n3613 = n2982 & n3612;
  assign n3614 = n620 & n3611;
  assign n3615 = n3613 & n3614;
  assign n3616 = n338 & n3615;
  assign n3617 = n2095 & n3616;
  assign n3618 = ~n3607 & n3617;
  assign n3619 = n3607 & ~n3617;
  assign n3620 = ~n3618 & ~n3619;
  assign n3621 = ~n3494 & n3620;
  assign n3622 = n3494 & ~n3620;
  assign n3623 = ~n3621 & ~n3622;
  assign n3624 = ~n3430 & ~n3492;
  assign n3625 = ~n3493 & ~n3624;
  assign n3626 = n3623 & n3625;
  assign n3627 = ~n3623 & ~n3625;
  assign po0  = ~n3626 & ~n3627;
  assign n3629 = ~n3619 & ~n3621;
  assign n3630 = ~n3602 & ~n3606;
  assign n3631 = ~n225 & ~n356;
  assign n3632 = n146 & n3631;
  assign n3633 = n383 & n2033;
  assign n3634 = n2213 & n3633;
  assign n3635 = n3632 & n3634;
  assign n3636 = n547 & n3635;
  assign n3637 = n779 & n814;
  assign n3638 = ~n196 & ~n226;
  assign n3639 = ~n310 & n3638;
  assign n3640 = n381 & n3639;
  assign n3641 = n3637 & n3640;
  assign n3642 = n352 & n3641;
  assign n3643 = n1296 & n3642;
  assign n3644 = n3636 & n3643;
  assign n3645 = n2228 & n3644;
  assign n3646 = n3514 & ~n3645;
  assign n3647 = ~n3514 & n3645;
  assign n3648 = ~n3646 & ~n3647;
  assign n3649 = n3046 & n3648;
  assign n3650 = n3050 & ~n3516;
  assign n3651 = n3054 & ~n3371;
  assign n3652 = ~n3521 & ~n3524;
  assign n3653 = ~n3516 & ~n3648;
  assign n3654 = n3516 & ~n3645;
  assign n3655 = ~n3653 & ~n3654;
  assign n3656 = ~n3652 & ~n3655;
  assign n3657 = n3652 & n3655;
  assign n3658 = ~n3656 & ~n3657;
  assign n3659 = n3056 & n3658;
  assign n3660 = ~n3650 & ~n3651;
  assign n3661 = ~n3649 & n3660;
  assign n3662 = ~n3659 & n3661;
  assign n3663 = n2368 & ~n3662;
  assign n3664 = ~n2368 & n3662;
  assign n3665 = ~n3663 & ~n3664;
  assign n3666 = ~n3596 & ~n3599;
  assign n3667 = ~n3580 & ~n3584;
  assign n3668 = n2469 & ~n2906;
  assign n3669 = n2378 & n2477;
  assign n3670 = n2364 & n2474;
  assign n3671 = n2479 & n2916;
  assign n3672 = ~n3669 & ~n3670;
  assign n3673 = ~n3668 & n3672;
  assign n3674 = ~n3671 & n3673;
  assign n3675 = n869 & ~n3674;
  assign n3676 = ~n869 & n3674;
  assign n3677 = ~n3675 & ~n3676;
  assign n3678 = ~n3574 & ~n3577;
  assign n3679 = n2385 & n2510;
  assign n3680 = n2392 & n2508;
  assign n3681 = n2395 & n2518;
  assign n3682 = n2503 & n2745;
  assign n3683 = ~n3680 & ~n3681;
  assign n3684 = ~n3679 & n3683;
  assign n3685 = ~n3682 & n3684;
  assign n3686 = ~n519 & n3685;
  assign n3687 = n519 & ~n3685;
  assign n3688 = ~n3686 & ~n3687;
  assign n3689 = ~n605 & ~n2407;
  assign n3690 = n2398 & n2565;
  assign n3691 = n2401 & n2563;
  assign n3692 = n2404 & n2691;
  assign n3693 = n2558 & n2585;
  assign n3694 = ~n3691 & ~n3692;
  assign n3695 = ~n3690 & n3694;
  assign n3696 = ~n3693 & n3695;
  assign n3697 = n3689 & ~n3696;
  assign n3698 = ~n3689 & n3696;
  assign n3699 = ~n3697 & ~n3698;
  assign n3700 = ~n605 & n2410;
  assign n3701 = n3554 & n3700;
  assign n3702 = ~n3561 & ~n3701;
  assign n3703 = n3699 & ~n3702;
  assign n3704 = ~n3699 & n3702;
  assign n3705 = ~n3703 & ~n3704;
  assign n3706 = n3688 & n3705;
  assign n3707 = ~n3688 & ~n3705;
  assign n3708 = ~n3706 & ~n3707;
  assign n3709 = ~n3678 & n3708;
  assign n3710 = n3678 & ~n3708;
  assign n3711 = ~n3709 & ~n3710;
  assign n3712 = ~n3677 & n3711;
  assign n3713 = n3677 & ~n3711;
  assign n3714 = ~n3712 & ~n3713;
  assign n3715 = n3667 & ~n3714;
  assign n3716 = ~n3667 & n3714;
  assign n3717 = ~n3715 & ~n3716;
  assign n3718 = n2375 & ~n3038;
  assign n3719 = n2382 & ~n3049;
  assign n3720 = n2387 & ~n3053;
  assign n3721 = n2389 & n3073;
  assign n3722 = ~n3719 & ~n3720;
  assign n3723 = ~n3718 & n3722;
  assign n3724 = ~n3721 & n3723;
  assign n3725 = ~n57 & n3724;
  assign n3726 = n57 & ~n3724;
  assign n3727 = ~n3725 & ~n3726;
  assign n3728 = n3717 & n3727;
  assign n3729 = ~n3717 & ~n3727;
  assign n3730 = ~n3728 & ~n3729;
  assign n3731 = ~n3666 & n3730;
  assign n3732 = n3666 & ~n3730;
  assign n3733 = ~n3731 & ~n3732;
  assign n3734 = ~n3665 & n3733;
  assign n3735 = n3665 & ~n3733;
  assign n3736 = ~n3734 & ~n3735;
  assign n3737 = n3630 & ~n3736;
  assign n3738 = ~n3630 & n3736;
  assign n3739 = ~n3737 & ~n3738;
  assign n3740 = n963 & n1307;
  assign n3741 = ~n134 & ~n181;
  assign n3742 = ~n324 & ~n353;
  assign n3743 = ~n356 & ~n458;
  assign n3744 = n3742 & n3743;
  assign n3745 = n146 & n3741;
  assign n3746 = n614 & n2124;
  assign n3747 = n3745 & n3746;
  assign n3748 = n2982 & n3744;
  assign n3749 = n2989 & n3740;
  assign n3750 = n3748 & n3749;
  assign n3751 = n3747 & n3750;
  assign n3752 = n2068 & n3751;
  assign n3753 = n3413 & n3752;
  assign n3754 = ~n3739 & n3753;
  assign n3755 = n3739 & ~n3753;
  assign n3756 = ~n3754 & ~n3755;
  assign n3757 = ~n3629 & n3756;
  assign n3758 = n3629 & ~n3756;
  assign n3759 = ~n3757 & ~n3758;
  assign n3760 = ~pi22  & ~pi23 ;
  assign n3761 = pi22  & pi23 ;
  assign n3762 = ~n3760 & ~n3761;
  assign n3763 = po0  & n3762;
  assign n3764 = ~n3759 & n3763;
  assign n3765 = n3626 & n3759;
  assign n3766 = ~n3626 & ~n3759;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = ~n3763 & n3767;
  assign po1  = n3764 | n3768;
  assign n3770 = ~n3755 & ~n3757;
  assign n3771 = ~n3734 & ~n3738;
  assign n3772 = ~n3728 & ~n3731;
  assign n3773 = ~n3712 & ~n3716;
  assign n3774 = n2469 & ~n3053;
  assign n3775 = n2474 & ~n2906;
  assign n3776 = n2364 & n2477;
  assign n3777 = n2479 & n3279;
  assign n3778 = ~n3775 & ~n3776;
  assign n3779 = ~n3774 & n3778;
  assign n3780 = ~n3777 & n3779;
  assign n3781 = n869 & ~n3780;
  assign n3782 = ~n869 & n3780;
  assign n3783 = ~n3781 & ~n3782;
  assign n3784 = ~n3706 & ~n3709;
  assign n3785 = n2378 & n2510;
  assign n3786 = n2392 & n2518;
  assign n3787 = n2385 & n2508;
  assign n3788 = n2503 & n2730;
  assign n3789 = ~n3786 & ~n3787;
  assign n3790 = ~n3785 & n3789;
  assign n3791 = ~n3788 & n3790;
  assign n3792 = ~n519 & n3791;
  assign n3793 = n519 & ~n3791;
  assign n3794 = ~n3792 & ~n3793;
  assign n3795 = ~n605 & ~n2404;
  assign n3796 = n2395 & n2565;
  assign n3797 = n2398 & n2563;
  assign n3798 = n2401 & n2691;
  assign n3799 = n2481 & n2558;
  assign n3800 = ~n3797 & ~n3798;
  assign n3801 = ~n3796 & n3800;
  assign n3802 = ~n3799 & n3801;
  assign n3803 = n3795 & ~n3802;
  assign n3804 = ~n3795 & n3802;
  assign n3805 = ~n3803 & ~n3804;
  assign n3806 = ~n605 & n2407;
  assign n3807 = n3696 & n3806;
  assign n3808 = ~n3703 & ~n3807;
  assign n3809 = n3805 & ~n3808;
  assign n3810 = ~n3805 & n3808;
  assign n3811 = ~n3809 & ~n3810;
  assign n3812 = n3794 & n3811;
  assign n3813 = ~n3794 & ~n3811;
  assign n3814 = ~n3812 & ~n3813;
  assign n3815 = ~n3784 & n3814;
  assign n3816 = n3784 & ~n3814;
  assign n3817 = ~n3815 & ~n3816;
  assign n3818 = ~n3783 & n3817;
  assign n3819 = n3783 & ~n3817;
  assign n3820 = ~n3818 & ~n3819;
  assign n3821 = n3773 & ~n3820;
  assign n3822 = ~n3773 & n3820;
  assign n3823 = ~n3821 & ~n3822;
  assign n3824 = n2375 & ~n3371;
  assign n3825 = n2382 & ~n3038;
  assign n3826 = n2387 & ~n3049;
  assign n3827 = n2389 & n3381;
  assign n3828 = ~n3825 & ~n3826;
  assign n3829 = ~n3824 & n3828;
  assign n3830 = ~n3827 & n3829;
  assign n3831 = ~n57 & n3830;
  assign n3832 = n57 & ~n3830;
  assign n3833 = ~n3831 & ~n3832;
  assign n3834 = n3823 & n3833;
  assign n3835 = ~n3823 & ~n3833;
  assign n3836 = ~n3834 & ~n3835;
  assign n3837 = ~n3772 & n3836;
  assign n3838 = n3772 & ~n3836;
  assign n3839 = ~n3837 & ~n3838;
  assign n3840 = n3050 & n3648;
  assign n3841 = ~n3648 & n3656;
  assign n3842 = n3654 & ~n3656;
  assign n3843 = ~n3841 & ~n3842;
  assign n3844 = n3056 & ~n3843;
  assign n3845 = ~n3840 & ~n3844;
  assign n3846 = n3054 & ~n3516;
  assign n3847 = ~n2368 & ~n3846;
  assign n3848 = n3845 & ~n3847;
  assign n3849 = ~n2368 & ~n3845;
  assign n3850 = ~n3848 & ~n3849;
  assign n3851 = n3839 & n3850;
  assign n3852 = ~n3839 & ~n3850;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = ~n3771 & n3853;
  assign n3855 = n3771 & ~n3853;
  assign n3856 = ~n3854 & ~n3855;
  assign n3857 = ~n144 & ~n156;
  assign n3858 = ~n307 & n3857;
  assign n3859 = n1010 & n2327;
  assign n3860 = n3858 & n3859;
  assign n3861 = ~n207 & ~n233;
  assign n3862 = ~n310 & ~n343;
  assign n3863 = ~n345 & n3862;
  assign n3864 = n482 & n3861;
  assign n3865 = n621 & n3864;
  assign n3866 = n632 & n3863;
  assign n3867 = n3865 & n3866;
  assign n3868 = n3860 & n3867;
  assign n3869 = n293 & n3868;
  assign n3870 = n3471 & n3869;
  assign n3871 = n3856 & ~n3870;
  assign n3872 = ~n3856 & n3870;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = ~n3770 & n3873;
  assign n3875 = n3770 & ~n3873;
  assign n3876 = ~n3874 & ~n3875;
  assign n3877 = ~n3765 & ~n3876;
  assign n3878 = n3765 & n3876;
  assign n3879 = ~n3877 & ~n3878;
  assign n3880 = ~po0  & ~n3767;
  assign n3881 = n3762 & ~n3880;
  assign n3882 = n3879 & ~n3881;
  assign n3883 = ~n3879 & n3881;
  assign po2  = n3882 | n3883;
  assign n3885 = ~n3879 & n3880;
  assign n3886 = n3762 & ~n3885;
  assign n3887 = ~n3871 & ~n3874;
  assign n3888 = ~n3851 & ~n3854;
  assign n3889 = ~n3834 & ~n3837;
  assign n3890 = n3516 & ~n3656;
  assign n3891 = n3056 & ~n3890;
  assign n3892 = ~n3054 & ~n3891;
  assign n3893 = n3648 & ~n3892;
  assign n3894 = n2368 & n3893;
  assign n3895 = ~n2368 & ~n3893;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = ~n3818 & ~n3822;
  assign n3898 = n2469 & ~n3049;
  assign n3899 = n2474 & ~n3053;
  assign n3900 = n2477 & ~n2906;
  assign n3901 = n2479 & n3088;
  assign n3902 = ~n3899 & ~n3900;
  assign n3903 = ~n3898 & n3902;
  assign n3904 = ~n3901 & n3903;
  assign n3905 = n869 & ~n3904;
  assign n3906 = ~n869 & n3904;
  assign n3907 = ~n3905 & ~n3906;
  assign n3908 = ~n3812 & ~n3815;
  assign n3909 = n2364 & n2510;
  assign n3910 = n2378 & n2508;
  assign n3911 = n2385 & n2518;
  assign n3912 = n2455 & n2503;
  assign n3913 = ~n3910 & ~n3911;
  assign n3914 = ~n3909 & n3913;
  assign n3915 = ~n3912 & n3914;
  assign n3916 = ~n519 & n3915;
  assign n3917 = n519 & ~n3915;
  assign n3918 = ~n3916 & ~n3917;
  assign n3919 = ~n605 & ~n2401;
  assign n3920 = n2392 & n2565;
  assign n3921 = n2398 & n2691;
  assign n3922 = n2395 & n2563;
  assign n3923 = n2558 & n2711;
  assign n3924 = ~n3921 & ~n3922;
  assign n3925 = ~n3920 & n3924;
  assign n3926 = ~n3923 & n3925;
  assign n3927 = n3919 & ~n3926;
  assign n3928 = ~n3919 & n3926;
  assign n3929 = ~n3927 & ~n3928;
  assign n3930 = ~n605 & n2404;
  assign n3931 = n3802 & n3930;
  assign n3932 = ~n3809 & ~n3931;
  assign n3933 = n3929 & ~n3932;
  assign n3934 = ~n3929 & n3932;
  assign n3935 = ~n3933 & ~n3934;
  assign n3936 = n3918 & n3935;
  assign n3937 = ~n3918 & ~n3935;
  assign n3938 = ~n3936 & ~n3937;
  assign n3939 = ~n3908 & n3938;
  assign n3940 = n3908 & ~n3938;
  assign n3941 = ~n3939 & ~n3940;
  assign n3942 = ~n3907 & n3941;
  assign n3943 = n3907 & ~n3941;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = n3897 & ~n3944;
  assign n3946 = ~n3897 & n3944;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = n2375 & ~n3516;
  assign n3949 = n2382 & ~n3371;
  assign n3950 = n2387 & ~n3038;
  assign n3951 = n2389 & n3526;
  assign n3952 = ~n3949 & ~n3950;
  assign n3953 = ~n3948 & n3952;
  assign n3954 = ~n3951 & n3953;
  assign n3955 = ~n57 & n3954;
  assign n3956 = n57 & ~n3954;
  assign n3957 = ~n3955 & ~n3956;
  assign n3958 = n3947 & n3957;
  assign n3959 = ~n3947 & ~n3957;
  assign n3960 = ~n3958 & ~n3959;
  assign n3961 = ~n3896 & n3960;
  assign n3962 = n3896 & ~n3960;
  assign n3963 = ~n3961 & ~n3962;
  assign n3964 = ~n3889 & n3963;
  assign n3965 = n3889 & ~n3963;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = ~n3888 & n3966;
  assign n3968 = n3888 & ~n3966;
  assign n3969 = ~n3967 & ~n3968;
  assign n3970 = ~n185 & ~n264;
  assign n3971 = ~n267 & ~n315;
  assign n3972 = ~n341 & ~n353;
  assign n3973 = n3971 & n3972;
  assign n3974 = n459 & n3970;
  assign n3975 = n2124 & n3974;
  assign n3976 = n795 & n3973;
  assign n3977 = n3975 & n3976;
  assign n3978 = n232 & n402;
  assign n3979 = n3436 & n3978;
  assign n3980 = n1963 & n3977;
  assign n3981 = n3979 & n3980;
  assign n3982 = n1306 & n3981;
  assign n3983 = n3969 & ~n3982;
  assign n3984 = ~n3969 & n3982;
  assign n3985 = ~n3983 & ~n3984;
  assign n3986 = ~n3887 & n3985;
  assign n3987 = n3887 & ~n3985;
  assign n3988 = ~n3986 & ~n3987;
  assign n3989 = n3878 & n3988;
  assign n3990 = ~n3878 & ~n3988;
  assign n3991 = ~n3989 & ~n3990;
  assign n3992 = n3886 & n3991;
  assign n3993 = ~n3886 & ~n3991;
  assign po3  = ~n3992 & ~n3993;
  assign n3995 = ~n3983 & ~n3986;
  assign n3996 = ~n3964 & ~n3967;
  assign n3997 = ~n3958 & ~n3961;
  assign n3998 = ~n3942 & ~n3946;
  assign n3999 = n2469 & ~n3038;
  assign n4000 = n2474 & ~n3049;
  assign n4001 = n2477 & ~n3053;
  assign n4002 = n2479 & n3073;
  assign n4003 = ~n4000 & ~n4001;
  assign n4004 = ~n3999 & n4003;
  assign n4005 = ~n4002 & n4004;
  assign n4006 = ~n869 & n4005;
  assign n4007 = n869 & ~n4005;
  assign n4008 = ~n4006 & ~n4007;
  assign n4009 = ~n3936 & ~n3939;
  assign n4010 = n2385 & n2565;
  assign n4011 = n2392 & n2563;
  assign n4012 = n2395 & n2691;
  assign n4013 = n2558 & n2745;
  assign n4014 = ~n4011 & ~n4012;
  assign n4015 = ~n4010 & n4014;
  assign n4016 = ~n4013 & n4015;
  assign n4017 = n605 & ~n4016;
  assign n4018 = ~n605 & n4016;
  assign n4019 = ~n4017 & ~n4018;
  assign n4020 = ~n605 & n2398;
  assign n4021 = ~n2368 & n4020;
  assign n4022 = n2368 & ~n4020;
  assign n4023 = ~n4021 & ~n4022;
  assign n4024 = ~n4019 & n4023;
  assign n4025 = n4019 & ~n4023;
  assign n4026 = ~n4024 & ~n4025;
  assign n4027 = ~n605 & n2401;
  assign n4028 = n3926 & n4027;
  assign n4029 = ~n3933 & ~n4028;
  assign n4030 = n4026 & ~n4029;
  assign n4031 = ~n4026 & n4029;
  assign n4032 = ~n4030 & ~n4031;
  assign n4033 = n2510 & ~n2906;
  assign n4034 = n2378 & n2518;
  assign n4035 = n2364 & n2508;
  assign n4036 = n2503 & n2916;
  assign n4037 = ~n4034 & ~n4035;
  assign n4038 = ~n4033 & n4037;
  assign n4039 = ~n4036 & n4038;
  assign n4040 = n519 & ~n4039;
  assign n4041 = ~n519 & n4039;
  assign n4042 = ~n4040 & ~n4041;
  assign n4043 = n4032 & n4042;
  assign n4044 = ~n4032 & ~n4042;
  assign n4045 = ~n4043 & ~n4044;
  assign n4046 = ~n4009 & n4045;
  assign n4047 = n4009 & ~n4045;
  assign n4048 = ~n4046 & ~n4047;
  assign n4049 = ~n4008 & n4048;
  assign n4050 = n4008 & ~n4048;
  assign n4051 = ~n4049 & ~n4050;
  assign n4052 = ~n3998 & n4051;
  assign n4053 = n3998 & ~n4051;
  assign n4054 = ~n4052 & ~n4053;
  assign n4055 = n2375 & n3648;
  assign n4056 = n2382 & ~n3516;
  assign n4057 = n2387 & ~n3371;
  assign n4058 = n2389 & n3658;
  assign n4059 = ~n4056 & ~n4057;
  assign n4060 = ~n4055 & n4059;
  assign n4061 = ~n4058 & n4060;
  assign n4062 = n57 & ~n4061;
  assign n4063 = ~n57 & n4061;
  assign n4064 = ~n4062 & ~n4063;
  assign n4065 = n4054 & n4064;
  assign n4066 = ~n4054 & ~n4064;
  assign n4067 = ~n4065 & ~n4066;
  assign n4068 = ~n3997 & n4067;
  assign n4069 = n3997 & ~n4067;
  assign n4070 = ~n4068 & ~n4069;
  assign n4071 = n3996 & ~n4070;
  assign n4072 = ~n3996 & n4070;
  assign n4073 = ~n4071 & ~n4072;
  assign n4074 = ~n284 & ~n325;
  assign n4075 = ~n342 & n4074;
  assign n4076 = n347 & n521;
  assign n4077 = n645 & n2217;
  assign n4078 = n2327 & n4077;
  assign n4079 = n4075 & n4076;
  assign n4080 = n4078 & n4079;
  assign n4081 = n852 & n4080;
  assign n4082 = n217 & n4081;
  assign n4083 = n2259 & n4082;
  assign n4084 = ~n4073 & n4083;
  assign n4085 = n4073 & ~n4083;
  assign n4086 = ~n4084 & ~n4085;
  assign n4087 = ~n3995 & n4086;
  assign n4088 = n3995 & ~n4086;
  assign n4089 = ~n4087 & ~n4088;
  assign n4090 = ~n3989 & ~n4089;
  assign n4091 = n3989 & n4089;
  assign n4092 = ~n4090 & ~n4091;
  assign n4093 = n3885 & ~n3991;
  assign n4094 = n3762 & ~n4093;
  assign n4095 = n4092 & ~n4094;
  assign n4096 = ~n4092 & n4094;
  assign po4  = n4095 | n4096;
  assign n4098 = ~n4085 & ~n4087;
  assign n4099 = ~n4068 & ~n4072;
  assign n4100 = ~n4052 & ~n4065;
  assign n4101 = n2389 & ~n3843;
  assign n4102 = n2387 & ~n3516;
  assign n4103 = n2382 & n3648;
  assign n4104 = ~n4102 & ~n4103;
  assign n4105 = ~n4101 & n4104;
  assign n4106 = n57 & ~n4105;
  assign n4107 = ~n57 & n4105;
  assign n4108 = ~n4106 & ~n4107;
  assign n4109 = ~n4046 & ~n4049;
  assign n4110 = n2469 & ~n3371;
  assign n4111 = n2474 & ~n3038;
  assign n4112 = n2477 & ~n3049;
  assign n4113 = n2479 & n3381;
  assign n4114 = ~n4111 & ~n4112;
  assign n4115 = ~n4110 & n4114;
  assign n4116 = ~n4113 & n4115;
  assign n4117 = n869 & ~n4116;
  assign n4118 = ~n869 & n4116;
  assign n4119 = ~n4117 & ~n4118;
  assign n4120 = ~n4030 & ~n4043;
  assign n4121 = n2510 & ~n3053;
  assign n4122 = n2508 & ~n2906;
  assign n4123 = n2364 & n2518;
  assign n4124 = n2503 & n3279;
  assign n4125 = ~n4122 & ~n4123;
  assign n4126 = ~n4121 & n4125;
  assign n4127 = ~n4124 & n4126;
  assign n4128 = n519 & ~n4127;
  assign n4129 = ~n519 & n4127;
  assign n4130 = ~n4128 & ~n4129;
  assign n4131 = n2378 & n2565;
  assign n4132 = n2392 & n2691;
  assign n4133 = n2385 & n2563;
  assign n4134 = n2558 & n2730;
  assign n4135 = ~n4132 & ~n4133;
  assign n4136 = ~n4131 & n4135;
  assign n4137 = ~n4134 & n4136;
  assign n4138 = n605 & n4137;
  assign n4139 = ~n605 & ~n4137;
  assign n4140 = ~n4138 & ~n4139;
  assign n4141 = ~n4021 & ~n4024;
  assign n4142 = ~n605 & n2395;
  assign n4143 = ~n2368 & n4142;
  assign n4144 = n2368 & ~n4142;
  assign n4145 = ~n4143 & ~n4144;
  assign n4146 = ~n4141 & n4145;
  assign n4147 = n4141 & ~n4145;
  assign n4148 = ~n4146 & ~n4147;
  assign n4149 = n4140 & n4148;
  assign n4150 = ~n4140 & ~n4148;
  assign n4151 = ~n4149 & ~n4150;
  assign n4152 = n4130 & n4151;
  assign n4153 = ~n4130 & ~n4151;
  assign n4154 = ~n4152 & ~n4153;
  assign n4155 = ~n4120 & n4154;
  assign n4156 = n4120 & ~n4154;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = ~n4119 & n4157;
  assign n4159 = n4119 & ~n4157;
  assign n4160 = ~n4158 & ~n4159;
  assign n4161 = ~n4109 & n4160;
  assign n4162 = n4109 & ~n4160;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = n4108 & n4163;
  assign n4165 = ~n4108 & ~n4163;
  assign n4166 = ~n4164 & ~n4165;
  assign n4167 = ~n4100 & n4166;
  assign n4168 = n4100 & ~n4166;
  assign n4169 = ~n4167 & ~n4168;
  assign n4170 = ~n4099 & n4169;
  assign n4171 = n4099 & ~n4169;
  assign n4172 = ~n4170 & ~n4171;
  assign n4173 = ~n315 & n2215;
  assign n4174 = n483 & n2088;
  assign n4175 = ~n248 & ~n279;
  assign n4176 = ~n284 & ~n296;
  assign n4177 = n4175 & n4176;
  assign n4178 = n354 & n455;
  assign n4179 = n4177 & n4178;
  assign n4180 = n3740 & n4173;
  assign n4181 = n4174 & n4180;
  assign n4182 = n2107 & n4179;
  assign n4183 = n4181 & n4182;
  assign n4184 = n2999 & n4183;
  assign n4185 = n3636 & n4184;
  assign n4186 = ~n4172 & n4185;
  assign n4187 = n4172 & ~n4185;
  assign n4188 = ~n4186 & ~n4187;
  assign n4189 = ~n4098 & n4188;
  assign n4190 = n4098 & ~n4188;
  assign n4191 = ~n4189 & ~n4190;
  assign n4192 = ~n4091 & ~n4191;
  assign n4193 = n4091 & n4191;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = ~n4092 & n4093;
  assign n4196 = n3762 & ~n4195;
  assign n4197 = n4194 & ~n4196;
  assign n4198 = ~n4194 & n4196;
  assign po5  = n4197 | n4198;
  assign n4200 = ~n4187 & ~n4189;
  assign n4201 = ~n4167 & ~n4170;
  assign n4202 = ~n4161 & ~n4164;
  assign n4203 = ~n4155 & ~n4158;
  assign n4204 = n2389 & ~n3890;
  assign n4205 = ~n2387 & ~n4204;
  assign n4206 = n3648 & ~n4205;
  assign n4207 = ~n57 & n4206;
  assign n4208 = n57 & ~n4206;
  assign n4209 = ~n4207 & ~n4208;
  assign n4210 = ~n4203 & ~n4209;
  assign n4211 = n4203 & n4209;
  assign n4212 = ~n4210 & ~n4211;
  assign n4213 = n2469 & ~n3516;
  assign n4214 = n2474 & ~n3371;
  assign n4215 = n2477 & ~n3038;
  assign n4216 = n2479 & n3526;
  assign n4217 = ~n4214 & ~n4215;
  assign n4218 = ~n4213 & n4217;
  assign n4219 = ~n4216 & n4218;
  assign n4220 = n869 & ~n4219;
  assign n4221 = ~n869 & n4219;
  assign n4222 = ~n4220 & ~n4221;
  assign n4223 = ~n4149 & ~n4152;
  assign n4224 = n2510 & ~n3049;
  assign n4225 = n2508 & ~n3053;
  assign n4226 = n2518 & ~n2906;
  assign n4227 = n2503 & n3088;
  assign n4228 = ~n4225 & ~n4226;
  assign n4229 = ~n4224 & n4228;
  assign n4230 = ~n4227 & n4229;
  assign n4231 = n519 & ~n4230;
  assign n4232 = ~n519 & n4230;
  assign n4233 = ~n4231 & ~n4232;
  assign n4234 = n2364 & n2565;
  assign n4235 = n2378 & n2563;
  assign n4236 = n2385 & n2691;
  assign n4237 = n2455 & n2558;
  assign n4238 = ~n4235 & ~n4236;
  assign n4239 = ~n4234 & n4238;
  assign n4240 = ~n4237 & n4239;
  assign n4241 = n605 & n4240;
  assign n4242 = ~n605 & ~n4240;
  assign n4243 = ~n4241 & ~n4242;
  assign n4244 = ~n4143 & ~n4146;
  assign n4245 = ~n605 & n2392;
  assign n4246 = ~n2368 & n4245;
  assign n4247 = n2368 & ~n4245;
  assign n4248 = ~n4246 & ~n4247;
  assign n4249 = ~n4244 & n4248;
  assign n4250 = n4244 & ~n4248;
  assign n4251 = ~n4249 & ~n4250;
  assign n4252 = n4243 & n4251;
  assign n4253 = ~n4243 & ~n4251;
  assign n4254 = ~n4252 & ~n4253;
  assign n4255 = n4233 & n4254;
  assign n4256 = ~n4233 & ~n4254;
  assign n4257 = ~n4255 & ~n4256;
  assign n4258 = ~n4223 & n4257;
  assign n4259 = n4223 & ~n4257;
  assign n4260 = ~n4258 & ~n4259;
  assign n4261 = ~n4222 & n4260;
  assign n4262 = n4222 & ~n4260;
  assign n4263 = ~n4261 & ~n4262;
  assign n4264 = n4212 & n4263;
  assign n4265 = ~n4212 & ~n4263;
  assign n4266 = ~n4264 & ~n4265;
  assign n4267 = ~n4202 & n4266;
  assign n4268 = n4202 & ~n4266;
  assign n4269 = ~n4267 & ~n4268;
  assign n4270 = ~n4201 & n4269;
  assign n4271 = n4201 & ~n4269;
  assign n4272 = ~n4270 & ~n4271;
  assign n4273 = ~n309 & n409;
  assign n4274 = n2088 & n2124;
  assign n4275 = n2246 & n4274;
  assign n4276 = n425 & n4273;
  assign n4277 = n3637 & n4276;
  assign n4278 = n2220 & n4275;
  assign n4279 = n4277 & n4278;
  assign n4280 = ~n149 & ~n180;
  assign n4281 = ~n271 & ~n329;
  assign n4282 = n4280 & n4281;
  assign n4283 = n845 & n2087;
  assign n4284 = n3026 & n4283;
  assign n4285 = n2253 & n4282;
  assign n4286 = n4284 & n4285;
  assign n4287 = n4279 & n4286;
  assign n4288 = n3416 & n4287;
  assign n4289 = ~n4272 & n4288;
  assign n4290 = n4272 & ~n4288;
  assign n4291 = ~n4289 & ~n4290;
  assign n4292 = ~n4200 & n4291;
  assign n4293 = n4200 & ~n4291;
  assign n4294 = ~n4292 & ~n4293;
  assign n4295 = ~n4193 & ~n4294;
  assign n4296 = n4193 & n4294;
  assign n4297 = ~n4295 & ~n4296;
  assign n4298 = ~n4194 & n4195;
  assign n4299 = n3762 & ~n4298;
  assign n4300 = n4297 & ~n4299;
  assign n4301 = ~n4297 & n4299;
  assign po6  = n4300 | n4301;
  assign n4303 = ~n4290 & ~n4292;
  assign n4304 = ~n4267 & ~n4270;
  assign n4305 = ~n4210 & ~n4264;
  assign n4306 = ~n4258 & ~n4261;
  assign n4307 = n2469 & n3648;
  assign n4308 = n2474 & ~n3516;
  assign n4309 = n2477 & ~n3371;
  assign n4310 = n2479 & n3658;
  assign n4311 = ~n4308 & ~n4309;
  assign n4312 = ~n4307 & n4311;
  assign n4313 = ~n4310 & n4312;
  assign n4314 = n869 & n4313;
  assign n4315 = ~n869 & ~n4313;
  assign n4316 = ~n4314 & ~n4315;
  assign n4317 = ~n4306 & n4316;
  assign n4318 = n4306 & ~n4316;
  assign n4319 = ~n4317 & ~n4318;
  assign n4320 = ~n4252 & ~n4255;
  assign n4321 = ~n4246 & ~n4249;
  assign n4322 = n2565 & ~n2906;
  assign n4323 = n2378 & n2691;
  assign n4324 = n2364 & n2563;
  assign n4325 = n2558 & n2916;
  assign n4326 = ~n4323 & ~n4324;
  assign n4327 = ~n4322 & n4326;
  assign n4328 = ~n4325 & n4327;
  assign n4329 = n605 & ~n4328;
  assign n4330 = ~n605 & n4328;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = ~n605 & n2385;
  assign n4333 = ~n57 & n2368;
  assign n4334 = n57 & ~n2368;
  assign n4335 = ~n4333 & ~n4334;
  assign n4336 = n4332 & n4335;
  assign n4337 = ~n4332 & ~n4335;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = ~n4331 & n4338;
  assign n4340 = n4331 & ~n4338;
  assign n4341 = ~n4339 & ~n4340;
  assign n4342 = ~n4321 & n4341;
  assign n4343 = n4321 & ~n4341;
  assign n4344 = ~n4342 & ~n4343;
  assign n4345 = n2510 & ~n3038;
  assign n4346 = n2508 & ~n3049;
  assign n4347 = n2518 & ~n3053;
  assign n4348 = n2503 & n3073;
  assign n4349 = ~n4346 & ~n4347;
  assign n4350 = ~n4345 & n4349;
  assign n4351 = ~n4348 & n4350;
  assign n4352 = ~n519 & n4351;
  assign n4353 = n519 & ~n4351;
  assign n4354 = ~n4352 & ~n4353;
  assign n4355 = n4344 & n4354;
  assign n4356 = ~n4344 & ~n4354;
  assign n4357 = ~n4355 & ~n4356;
  assign n4358 = ~n4320 & n4357;
  assign n4359 = n4320 & ~n4357;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = n4319 & n4360;
  assign n4362 = ~n4319 & ~n4360;
  assign n4363 = ~n4361 & ~n4362;
  assign n4364 = ~n4305 & n4363;
  assign n4365 = n4305 & ~n4363;
  assign n4366 = ~n4364 & ~n4365;
  assign n4367 = n4304 & ~n4366;
  assign n4368 = ~n4304 & n4366;
  assign n4369 = ~n4367 & ~n4368;
  assign n4370 = ~n148 & ~n325;
  assign n4371 = ~n134 & ~n307;
  assign n4372 = n241 & n4371;
  assign n4373 = n344 & n752;
  assign n4374 = n966 & n4370;
  assign n4375 = n4373 & n4374;
  assign n4376 = n4173 & n4372;
  assign n4377 = n4375 & n4376;
  assign n4378 = n4279 & n4377;
  assign n4379 = n2073 & n4378;
  assign n4380 = n4369 & ~n4379;
  assign n4381 = ~n4369 & n4379;
  assign n4382 = ~n4380 & ~n4381;
  assign n4383 = ~n4303 & n4382;
  assign n4384 = n4303 & ~n4382;
  assign n4385 = ~n4383 & ~n4384;
  assign n4386 = n4296 & n4385;
  assign n4387 = ~n4296 & ~n4385;
  assign n4388 = ~n4386 & ~n4387;
  assign n4389 = ~n4297 & n4298;
  assign n4390 = n3762 & ~n4389;
  assign n4391 = n4388 & ~n4390;
  assign n4392 = ~n4388 & n4390;
  assign po7  = n4391 | n4392;
  assign n4394 = ~n4380 & ~n4383;
  assign n4395 = ~n4364 & ~n4368;
  assign n4396 = ~n4317 & ~n4361;
  assign n4397 = n2479 & ~n3843;
  assign n4398 = n2477 & ~n3516;
  assign n4399 = n2474 & n3648;
  assign n4400 = ~n4398 & ~n4399;
  assign n4401 = ~n4397 & n4400;
  assign n4402 = n869 & ~n4401;
  assign n4403 = ~n869 & n4401;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = ~n4355 & ~n4358;
  assign n4406 = n2510 & ~n3371;
  assign n4407 = n2508 & ~n3038;
  assign n4408 = n2518 & ~n3049;
  assign n4409 = n2503 & n3381;
  assign n4410 = ~n4407 & ~n4408;
  assign n4411 = ~n4406 & n4410;
  assign n4412 = ~n4409 & n4411;
  assign n4413 = n519 & ~n4412;
  assign n4414 = ~n519 & n4412;
  assign n4415 = ~n4413 & ~n4414;
  assign n4416 = ~n4339 & ~n4342;
  assign n4417 = n2565 & ~n3053;
  assign n4418 = n2563 & ~n2906;
  assign n4419 = n2364 & n2691;
  assign n4420 = n2558 & n3279;
  assign n4421 = ~n4418 & ~n4419;
  assign n4422 = ~n4417 & n4421;
  assign n4423 = ~n4420 & n4422;
  assign n4424 = n605 & n4423;
  assign n4425 = ~n605 & ~n4423;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = ~n605 & n2378;
  assign n4428 = ~n4333 & ~n4336;
  assign n4429 = ~n4427 & ~n4428;
  assign n4430 = n4427 & n4428;
  assign n4431 = ~n4429 & ~n4430;
  assign n4432 = n4426 & n4431;
  assign n4433 = ~n4426 & ~n4431;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = ~n4416 & n4434;
  assign n4436 = n4416 & ~n4434;
  assign n4437 = ~n4435 & ~n4436;
  assign n4438 = n4415 & n4437;
  assign n4439 = ~n4415 & ~n4437;
  assign n4440 = ~n4438 & ~n4439;
  assign n4441 = ~n4405 & n4440;
  assign n4442 = n4405 & ~n4440;
  assign n4443 = ~n4441 & ~n4442;
  assign n4444 = ~n4404 & n4443;
  assign n4445 = n4404 & ~n4443;
  assign n4446 = ~n4444 & ~n4445;
  assign n4447 = ~n4396 & n4446;
  assign n4448 = n4396 & ~n4446;
  assign n4449 = ~n4447 & ~n4448;
  assign n4450 = ~n4395 & n4449;
  assign n4451 = n4395 & ~n4449;
  assign n4452 = ~n4450 & ~n4451;
  assign n4453 = ~n137 & ~n192;
  assign n4454 = ~n222 & n4453;
  assign n4455 = n316 & n553;
  assign n4456 = n2032 & n4455;
  assign n4457 = n4454 & n4456;
  assign n4458 = n1968 & n4457;
  assign n4459 = n421 & n4458;
  assign n4460 = ~n125 & ~n247;
  assign n4461 = ~n457 & ~n530;
  assign n4462 = ~n543 & n4461;
  assign n4463 = n2127 & n4460;
  assign n4464 = n4462 & n4463;
  assign n4465 = n820 & n2125;
  assign n4466 = n4464 & n4465;
  assign n4467 = n817 & n4466;
  assign n4468 = n3454 & n4467;
  assign n4469 = n4459 & n4468;
  assign n4470 = ~n4452 & n4469;
  assign n4471 = n4452 & ~n4469;
  assign n4472 = ~n4470 & ~n4471;
  assign n4473 = ~n4394 & n4472;
  assign n4474 = n4394 & ~n4472;
  assign n4475 = ~n4473 & ~n4474;
  assign n4476 = ~n4386 & ~n4475;
  assign n4477 = n4386 & n4475;
  assign n4478 = ~n4476 & ~n4477;
  assign n4479 = ~n4388 & n4389;
  assign n4480 = n3762 & ~n4479;
  assign n4481 = n4478 & ~n4480;
  assign n4482 = ~n4478 & n4480;
  assign po8  = n4481 | n4482;
  assign n4484 = ~n4471 & ~n4473;
  assign n4485 = ~n4447 & ~n4450;
  assign n4486 = ~n4441 & ~n4444;
  assign n4487 = ~n4435 & ~n4438;
  assign n4488 = n2479 & ~n3890;
  assign n4489 = ~n2477 & ~n4488;
  assign n4490 = n3648 & ~n4489;
  assign n4491 = ~n869 & ~n4490;
  assign n4492 = n869 & n4490;
  assign n4493 = ~n4491 & ~n4492;
  assign n4494 = ~n4487 & ~n4493;
  assign n4495 = n4487 & n4493;
  assign n4496 = ~n4494 & ~n4495;
  assign n4497 = ~n4429 & ~n4432;
  assign n4498 = n2565 & ~n3049;
  assign n4499 = n2563 & ~n3053;
  assign n4500 = n2691 & ~n2906;
  assign n4501 = n2558 & n3088;
  assign n4502 = ~n4499 & ~n4500;
  assign n4503 = ~n4498 & n4502;
  assign n4504 = ~n4501 & n4503;
  assign n4505 = n605 & ~n4504;
  assign n4506 = ~n605 & n4504;
  assign n4507 = ~n4505 & ~n4506;
  assign n4508 = ~n605 & n2452;
  assign n4509 = ~n4507 & ~n4508;
  assign n4510 = n4507 & n4508;
  assign n4511 = ~n4509 & ~n4510;
  assign n4512 = ~n4497 & n4511;
  assign n4513 = n4497 & ~n4511;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = n2510 & ~n3516;
  assign n4516 = n2508 & ~n3371;
  assign n4517 = n2518 & ~n3038;
  assign n4518 = n2503 & n3526;
  assign n4519 = ~n4516 & ~n4517;
  assign n4520 = ~n4515 & n4519;
  assign n4521 = ~n4518 & n4520;
  assign n4522 = n519 & ~n4521;
  assign n4523 = ~n519 & n4521;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = n4514 & n4524;
  assign n4526 = ~n4514 & ~n4524;
  assign n4527 = ~n4525 & ~n4526;
  assign n4528 = n4496 & n4527;
  assign n4529 = ~n4496 & ~n4527;
  assign n4530 = ~n4528 & ~n4529;
  assign n4531 = ~n4486 & n4530;
  assign n4532 = n4486 & ~n4530;
  assign n4533 = ~n4531 & ~n4532;
  assign n4534 = n4485 & ~n4533;
  assign n4535 = ~n4485 & n4533;
  assign n4536 = ~n4534 & ~n4535;
  assign n4537 = ~n171 & ~n200;
  assign n4538 = ~n280 & ~n311;
  assign n4539 = ~n458 & n4538;
  assign n4540 = n344 & n4537;
  assign n4541 = n2098 & n3026;
  assign n4542 = n4540 & n4541;
  assign n4543 = n2989 & n4539;
  assign n4544 = n4542 & n4543;
  assign n4545 = n161 & n4544;
  assign n4546 = n3398 & n4545;
  assign n4547 = n2228 & n4546;
  assign n4548 = ~n4536 & n4547;
  assign n4549 = n4536 & ~n4547;
  assign n4550 = ~n4548 & ~n4549;
  assign n4551 = ~n4484 & n4550;
  assign n4552 = n4484 & ~n4550;
  assign n4553 = ~n4551 & ~n4552;
  assign n4554 = ~n4477 & ~n4553;
  assign n4555 = n4477 & n4553;
  assign n4556 = ~n4554 & ~n4555;
  assign n4557 = ~n4478 & n4479;
  assign n4558 = n3762 & ~n4557;
  assign n4559 = n4556 & ~n4558;
  assign n4560 = ~n4556 & n4558;
  assign po9  = n4559 | n4560;
  assign n4562 = ~n4549 & ~n4551;
  assign n4563 = ~n4531 & ~n4535;
  assign n4564 = ~n4494 & ~n4528;
  assign n4565 = ~n4512 & ~n4525;
  assign n4566 = n2510 & n3648;
  assign n4567 = n2508 & ~n3516;
  assign n4568 = n2518 & ~n3371;
  assign n4569 = n2503 & n3658;
  assign n4570 = ~n4567 & ~n4568;
  assign n4571 = ~n4566 & n4570;
  assign n4572 = ~n4569 & n4571;
  assign n4573 = ~n519 & n4572;
  assign n4574 = n519 & ~n4572;
  assign n4575 = ~n4573 & ~n4574;
  assign n4576 = ~n4565 & n4575;
  assign n4577 = n4565 & ~n4575;
  assign n4578 = ~n4576 & ~n4577;
  assign n4579 = n2565 & ~n3038;
  assign n4580 = n2563 & ~n3049;
  assign n4581 = n2691 & ~n3053;
  assign n4582 = n2558 & n3073;
  assign n4583 = ~n4580 & ~n4581;
  assign n4584 = ~n4579 & n4583;
  assign n4585 = ~n4582 & n4584;
  assign n4586 = ~n605 & n4585;
  assign n4587 = n605 & ~n4585;
  assign n4588 = ~n4586 & ~n4587;
  assign n4589 = ~n605 & ~n2906;
  assign n4590 = ~n869 & ~n4589;
  assign n4591 = n869 & n4589;
  assign n4592 = ~n4590 & ~n4591;
  assign n4593 = n4427 & ~n4592;
  assign n4594 = ~n4427 & n4592;
  assign n4595 = ~n4593 & ~n4594;
  assign n4596 = ~n605 & ~n2378;
  assign n4597 = n2364 & n4596;
  assign n4598 = ~n4509 & ~n4597;
  assign n4599 = ~n4595 & ~n4598;
  assign n4600 = n4595 & n4598;
  assign n4601 = ~n4599 & ~n4600;
  assign n4602 = n4588 & ~n4601;
  assign n4603 = ~n4588 & n4601;
  assign n4604 = ~n4602 & ~n4603;
  assign n4605 = n4578 & n4604;
  assign n4606 = ~n4578 & ~n4604;
  assign n4607 = ~n4605 & ~n4606;
  assign n4608 = ~n4564 & n4607;
  assign n4609 = n4564 & ~n4607;
  assign n4610 = ~n4608 & ~n4609;
  assign n4611 = ~n4563 & n4610;
  assign n4612 = n4563 & ~n4610;
  assign n4613 = ~n4611 & ~n4612;
  assign n4614 = ~n238 & ~n399;
  assign n4615 = ~n469 & n4614;
  assign n4616 = n330 & n2326;
  assign n4617 = n3026 & n4616;
  assign n4618 = n184 & n4615;
  assign n4619 = n815 & n2982;
  assign n4620 = n4618 & n4619;
  assign n4621 = n4617 & n4620;
  assign n4622 = n613 & n4621;
  assign n4623 = n978 & n3443;
  assign n4624 = n4622 & n4623;
  assign n4625 = ~n4613 & n4624;
  assign n4626 = n4613 & ~n4624;
  assign n4627 = ~n4625 & ~n4626;
  assign n4628 = ~n4562 & n4627;
  assign n4629 = n4562 & ~n4627;
  assign n4630 = ~n4628 & ~n4629;
  assign n4631 = ~n4555 & ~n4630;
  assign n4632 = n4555 & n4630;
  assign n4633 = ~n4631 & ~n4632;
  assign n4634 = ~n4556 & n4557;
  assign n4635 = n3762 & ~n4634;
  assign n4636 = n4633 & ~n4635;
  assign n4637 = ~n4633 & n4635;
  assign po10  = n4636 | n4637;
  assign n4639 = ~n4626 & ~n4628;
  assign n4640 = ~n4608 & ~n4611;
  assign n4641 = ~n4576 & ~n4605;
  assign n4642 = n2503 & ~n3843;
  assign n4643 = n2518 & ~n3516;
  assign n4644 = n2508 & n3648;
  assign n4645 = ~n4643 & ~n4644;
  assign n4646 = ~n4642 & n4645;
  assign n4647 = n519 & ~n4646;
  assign n4648 = ~n519 & n4646;
  assign n4649 = ~n4647 & ~n4648;
  assign n4650 = n2565 & ~n3371;
  assign n4651 = n2563 & ~n3038;
  assign n4652 = n2691 & ~n3049;
  assign n4653 = n2558 & n3381;
  assign n4654 = ~n4651 & ~n4652;
  assign n4655 = ~n4650 & n4654;
  assign n4656 = ~n4653 & n4655;
  assign n4657 = n605 & n4656;
  assign n4658 = ~n605 & ~n4656;
  assign n4659 = ~n4657 & ~n4658;
  assign n4660 = ~n605 & ~n3053;
  assign n4661 = ~n4427 & ~n4591;
  assign n4662 = ~n4590 & ~n4661;
  assign n4663 = ~n4660 & n4662;
  assign n4664 = n4660 & ~n4662;
  assign n4665 = ~n4663 & ~n4664;
  assign n4666 = n4659 & n4665;
  assign n4667 = ~n4659 & ~n4665;
  assign n4668 = ~n4666 & ~n4667;
  assign n4669 = n4588 & ~n4599;
  assign n4670 = ~n4600 & ~n4669;
  assign n4671 = n4668 & n4670;
  assign n4672 = ~n4668 & ~n4670;
  assign n4673 = ~n4671 & ~n4672;
  assign n4674 = n4649 & n4673;
  assign n4675 = ~n4649 & ~n4673;
  assign n4676 = ~n4674 & ~n4675;
  assign n4677 = ~n4641 & n4676;
  assign n4678 = n4641 & ~n4676;
  assign n4679 = ~n4677 & ~n4678;
  assign n4680 = ~n4640 & n4679;
  assign n4681 = n4640 & ~n4679;
  assign n4682 = ~n4680 & ~n4681;
  assign n4683 = n524 & n772;
  assign n4684 = n542 & n1000;
  assign n4685 = n4683 & n4684;
  assign n4686 = n3501 & n4685;
  assign n4687 = n643 & n4686;
  assign n4688 = ~n4682 & n4687;
  assign n4689 = n4682 & ~n4687;
  assign n4690 = ~n4688 & ~n4689;
  assign n4691 = ~n4639 & n4690;
  assign n4692 = n4639 & ~n4690;
  assign n4693 = ~n4691 & ~n4692;
  assign n4694 = ~n4632 & ~n4693;
  assign n4695 = n4632 & n4693;
  assign n4696 = ~n4694 & ~n4695;
  assign n4697 = ~n4633 & n4634;
  assign n4698 = n3762 & ~n4697;
  assign n4699 = n4696 & ~n4698;
  assign n4700 = ~n4696 & n4698;
  assign po11  = n4699 | n4700;
  assign n4702 = ~n4689 & ~n4691;
  assign n4703 = ~n4677 & ~n4680;
  assign n4704 = ~n4671 & ~n4674;
  assign n4705 = ~n4663 & ~n4666;
  assign n4706 = ~n605 & n3065;
  assign n4707 = ~n4705 & ~n4706;
  assign n4708 = n4705 & n4706;
  assign n4709 = ~n4707 & ~n4708;
  assign n4710 = n2565 & ~n3516;
  assign n4711 = n2563 & ~n3371;
  assign n4712 = n2691 & ~n3038;
  assign n4713 = n2558 & n3526;
  assign n4714 = ~n4711 & ~n4712;
  assign n4715 = ~n4710 & n4714;
  assign n4716 = ~n4713 & n4715;
  assign n4717 = ~n605 & n4716;
  assign n4718 = n605 & ~n4716;
  assign n4719 = ~n4717 & ~n4718;
  assign n4720 = n2503 & ~n3890;
  assign n4721 = ~n2518 & ~n4720;
  assign n4722 = n3648 & ~n4721;
  assign n4723 = ~n519 & n4722;
  assign n4724 = n519 & ~n4722;
  assign n4725 = ~n4723 & ~n4724;
  assign n4726 = ~n4719 & ~n4725;
  assign n4727 = n4719 & n4725;
  assign n4728 = ~n4726 & ~n4727;
  assign n4729 = n4709 & n4728;
  assign n4730 = ~n4709 & ~n4728;
  assign n4731 = ~n4729 & ~n4730;
  assign n4732 = ~n4704 & n4731;
  assign n4733 = n4704 & ~n4731;
  assign n4734 = ~n4732 & ~n4733;
  assign n4735 = ~n4703 & n4734;
  assign n4736 = n4703 & ~n4734;
  assign n4737 = ~n4735 & ~n4736;
  assign n4738 = n115 & n133;
  assign n4739 = ~n139 & ~n273;
  assign n4740 = ~n372 & ~n457;
  assign n4741 = ~n520 & n4740;
  assign n4742 = n4739 & n4741;
  assign n4743 = ~n137 & ~n4738;
  assign n4744 = n2148 & n4743;
  assign n4745 = n795 & n4744;
  assign n4746 = n3860 & n4745;
  assign n4747 = n4742 & n4746;
  assign n4748 = n2031 & n4747;
  assign n4749 = n2165 & n4748;
  assign n4750 = ~n4737 & n4749;
  assign n4751 = n4737 & ~n4749;
  assign n4752 = ~n4750 & ~n4751;
  assign n4753 = ~n4702 & n4752;
  assign n4754 = n4702 & ~n4752;
  assign n4755 = ~n4753 & ~n4754;
  assign n4756 = ~n4695 & ~n4755;
  assign n4757 = n4695 & n4755;
  assign n4758 = ~n4756 & ~n4757;
  assign n4759 = ~n4696 & n4697;
  assign n4760 = n3762 & ~n4759;
  assign n4761 = n4758 & ~n4760;
  assign n4762 = ~n4758 & n4760;
  assign po12  = n4761 | n4762;
  assign n4764 = ~n4751 & ~n4753;
  assign n4765 = ~n4732 & ~n4735;
  assign n4766 = ~n4726 & ~n4729;
  assign n4767 = n3049 & n4660;
  assign n4768 = ~n4707 & ~n4767;
  assign n4769 = n2565 & n3648;
  assign n4770 = n2563 & ~n3516;
  assign n4771 = n2691 & ~n3371;
  assign n4772 = n2558 & n3658;
  assign n4773 = ~n4770 & ~n4771;
  assign n4774 = ~n4769 & n4773;
  assign n4775 = ~n4772 & n4774;
  assign n4776 = n605 & ~n4775;
  assign n4777 = ~n605 & n4775;
  assign n4778 = ~n4776 & ~n4777;
  assign n4779 = ~n605 & ~n3049;
  assign n4780 = ~n519 & n4779;
  assign n4781 = n519 & ~n4779;
  assign n4782 = ~n4780 & ~n4781;
  assign n4783 = ~n605 & ~n3038;
  assign n4784 = n4782 & n4783;
  assign n4785 = ~n4782 & ~n4783;
  assign n4786 = ~n4784 & ~n4785;
  assign n4787 = ~n4778 & n4786;
  assign n4788 = n4778 & ~n4786;
  assign n4789 = ~n4787 & ~n4788;
  assign n4790 = ~n4768 & n4789;
  assign n4791 = n4768 & ~n4789;
  assign n4792 = ~n4790 & ~n4791;
  assign n4793 = ~n4766 & n4792;
  assign n4794 = n4766 & ~n4792;
  assign n4795 = ~n4793 & ~n4794;
  assign n4796 = ~n4765 & n4795;
  assign n4797 = n4765 & ~n4795;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = ~n306 & ~n325;
  assign n4800 = ~n356 & ~n436;
  assign n4801 = ~n481 & n4800;
  assign n4802 = n4799 & n4801;
  assign n4803 = ~n125 & ~n129;
  assign n4804 = ~n197 & ~n226;
  assign n4805 = ~n428 & n4804;
  assign n4806 = n409 & n4803;
  assign n4807 = n827 & n1013;
  assign n4808 = n4806 & n4807;
  assign n4809 = n3740 & n4805;
  assign n4810 = n4808 & n4809;
  assign n4811 = n4802 & n4810;
  assign n4812 = n951 & n4811;
  assign n4813 = n1987 & n3471;
  assign n4814 = n4812 & n4813;
  assign n4815 = n4798 & ~n4814;
  assign n4816 = ~n4798 & n4814;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = ~n4764 & n4817;
  assign n4819 = n4764 & ~n4817;
  assign n4820 = ~n4818 & ~n4819;
  assign n4821 = ~n4757 & ~n4820;
  assign n4822 = n4757 & n4820;
  assign n4823 = ~n4821 & ~n4822;
  assign n4824 = ~n4758 & n4759;
  assign n4825 = n3762 & ~n4824;
  assign n4826 = n4823 & ~n4825;
  assign n4827 = ~n4823 & n4825;
  assign po13  = n4826 | n4827;
  assign n4829 = ~n4815 & ~n4818;
  assign n4830 = ~n4793 & ~n4796;
  assign n4831 = ~n4787 & ~n4790;
  assign n4832 = n2558 & ~n3843;
  assign n4833 = n2691 & ~n3516;
  assign n4834 = n2563 & n3648;
  assign n4835 = ~n4833 & ~n4834;
  assign n4836 = ~n4832 & n4835;
  assign n4837 = n605 & n4836;
  assign n4838 = ~n605 & ~n4836;
  assign n4839 = ~n4837 & ~n4838;
  assign n4840 = ~n605 & ~n3371;
  assign n4841 = ~n4780 & ~n4784;
  assign n4842 = ~n4840 & ~n4841;
  assign n4843 = n4840 & n4841;
  assign n4844 = ~n4842 & ~n4843;
  assign n4845 = n4839 & n4844;
  assign n4846 = ~n4839 & ~n4844;
  assign n4847 = ~n4845 & ~n4846;
  assign n4848 = ~n4831 & n4847;
  assign n4849 = n4831 & ~n4847;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n4830 & n4850;
  assign n4852 = n4830 & ~n4850;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = ~n154 & ~n198;
  assign n4855 = ~n268 & ~n303;
  assign n4856 = ~n428 & n4855;
  assign n4857 = n265 & n4854;
  assign n4858 = n538 & n2148;
  assign n4859 = n2213 & n3026;
  assign n4860 = n4858 & n4859;
  assign n4861 = n4856 & n4857;
  assign n4862 = n4860 & n4861;
  assign n4863 = n830 & n4862;
  assign n4864 = n825 & n1288;
  assign n4865 = n4863 & n4864;
  assign n4866 = n1975 & n4865;
  assign n4867 = ~n4853 & n4866;
  assign n4868 = n4853 & ~n4866;
  assign n4869 = ~n4867 & ~n4868;
  assign n4870 = ~n4829 & n4869;
  assign n4871 = n4829 & ~n4869;
  assign n4872 = ~n4870 & ~n4871;
  assign n4873 = ~n4822 & ~n4872;
  assign n4874 = n4822 & n4872;
  assign n4875 = ~n4873 & ~n4874;
  assign n4876 = ~n4823 & n4824;
  assign n4877 = n3762 & ~n4876;
  assign n4878 = n4875 & ~n4877;
  assign n4879 = ~n4875 & n4877;
  assign po14  = n4878 | n4879;
  assign n4881 = ~n4868 & ~n4870;
  assign n4882 = ~n4842 & ~n4845;
  assign n4883 = n2558 & ~n3890;
  assign n4884 = ~n2691 & ~n4883;
  assign n4885 = n3648 & ~n4884;
  assign n4886 = n605 & n4885;
  assign n4887 = ~n605 & ~n4885;
  assign n4888 = ~n4886 & ~n4887;
  assign n4889 = ~n605 & n3523;
  assign n4890 = ~n4888 & ~n4889;
  assign n4891 = n4885 & n4889;
  assign n4892 = ~n4890 & ~n4891;
  assign n4893 = n4882 & ~n4892;
  assign n4894 = ~n4882 & n4892;
  assign n4895 = ~n4893 & ~n4894;
  assign n4896 = ~n4848 & ~n4851;
  assign n4897 = ~n4895 & n4896;
  assign n4898 = n4895 & ~n4896;
  assign n4899 = ~n4897 & ~n4898;
  assign n4900 = ~n176 & ~n200;
  assign n4901 = ~n262 & n4900;
  assign n4902 = n1027 & n4901;
  assign n4903 = ~n182 & ~n263;
  assign n4904 = ~n299 & ~n311;
  assign n4905 = n4903 & n4904;
  assign n4906 = n629 & n845;
  assign n4907 = n3433 & n4906;
  assign n4908 = n4905 & n4907;
  assign n4909 = n4742 & n4908;
  assign n4910 = n957 & n4909;
  assign n4911 = n2155 & n4910;
  assign n4912 = n4902 & n4911;
  assign n4913 = n4899 & ~n4912;
  assign n4914 = ~n4899 & n4912;
  assign n4915 = ~n4913 & ~n4914;
  assign n4916 = ~n4881 & n4915;
  assign n4917 = n4881 & ~n4915;
  assign n4918 = ~n4916 & ~n4917;
  assign n4919 = ~n4874 & ~n4918;
  assign n4920 = n4874 & n4918;
  assign n4921 = ~n4919 & ~n4920;
  assign n4922 = ~n4875 & n4876;
  assign n4923 = n3762 & ~n4922;
  assign n4924 = n4921 & ~n4923;
  assign n4925 = ~n4921 & n4923;
  assign po15  = n4924 | n4925;
  assign n4927 = ~n4913 & ~n4916;
  assign n4928 = ~n237 & ~n298;
  assign n4929 = ~n461 & n4928;
  assign n4930 = n183 & n615;
  assign n4931 = n4929 & n4930;
  assign n4932 = n2046 & n4931;
  assign n4933 = n3404 & n4802;
  assign n4934 = n4932 & n4933;
  assign n4935 = n3474 & n4934;
  assign n4936 = n2097 & n4935;
  assign n4937 = ~n605 & ~n3513;
  assign n4938 = n3371 & n4937;
  assign n4939 = ~n4890 & ~n4938;
  assign n4940 = ~n4894 & ~n4898;
  assign n4941 = ~n3371 & ~n3648;
  assign n4942 = n3371 & ~n3645;
  assign n4943 = ~n605 & ~n4942;
  assign n4944 = ~n4941 & n4943;
  assign n4945 = n4940 & ~n4944;
  assign n4946 = ~n4940 & n4944;
  assign n4947 = ~n4945 & ~n4946;
  assign n4948 = n4939 & n4947;
  assign n4949 = ~n4939 & ~n4947;
  assign n4950 = ~n4948 & ~n4949;
  assign n4951 = ~n4936 & n4950;
  assign n4952 = n4936 & ~n4950;
  assign n4953 = ~n4951 & ~n4952;
  assign n4954 = n4927 & n4953;
  assign n4955 = ~n4927 & ~n4953;
  assign n4956 = ~n4954 & ~n4955;
  assign n4957 = ~n4920 & n4956;
  assign n4958 = n4920 & ~n4956;
  assign n4959 = ~n4957 & ~n4958;
  assign n4960 = ~n4921 & n4922;
  assign n4961 = n3762 & ~n4960;
  assign n4962 = n4959 & ~n4961;
  assign n4963 = ~n4959 & n4961;
  assign po16  = n4962 | n4963;
  assign n4965 = ~n4959 & n4960;
  assign n4966 = n3762 & ~n4965;
  assign n4967 = n4927 & ~n4951;
  assign n4968 = ~n4952 & ~n4967;
  assign n4969 = ~n140 & ~n208;
  assign n4970 = ~n210 & ~n223;
  assign n4971 = ~n457 & n4970;
  assign n4972 = n767 & n4969;
  assign n4973 = n827 & n2326;
  assign n4974 = n4972 & n4973;
  assign n4975 = n253 & n4971;
  assign n4976 = n4974 & n4975;
  assign n4977 = n411 & n4976;
  assign n4978 = n397 & n4977;
  assign n4979 = n2999 & n4978;
  assign n4980 = n4968 & ~n4979;
  assign n4981 = ~n4968 & n4979;
  assign n4982 = ~n4980 & ~n4981;
  assign n4983 = n4958 & n4982;
  assign n4984 = ~n4958 & ~n4982;
  assign n4985 = ~n4983 & ~n4984;
  assign n4986 = n4966 & n4985;
  assign n4987 = ~n4966 & ~n4985;
  assign po17  = ~n4986 & ~n4987;
  assign n4989 = n4965 & ~n4985;
  assign n4990 = n3762 & ~n4989;
  assign n4991 = ~n4980 & ~n4983;
  assign n4992 = ~n185 & ~n268;
  assign n4993 = ~n309 & ~n314;
  assign n4994 = ~n457 & n4993;
  assign n4995 = n4992 & n4994;
  assign n4996 = n632 & n833;
  assign n4997 = n4995 & n4996;
  assign n4998 = n962 & n1979;
  assign n4999 = n4997 & n4998;
  assign n5000 = n999 & n4999;
  assign n5001 = n3451 & n5000;
  assign n5002 = n423 & n5001;
  assign n5003 = ~n4991 & n5002;
  assign n5004 = n4991 & ~n5002;
  assign n5005 = ~n5003 & ~n5004;
  assign n5006 = n4990 & n5005;
  assign n5007 = ~n4990 & ~n5005;
  assign po18  = n5006 | n5007;
  assign n5009 = n4980 & ~n5002;
  assign n5010 = ~n145 & ~n209;
  assign n5011 = ~n304 & ~n327;
  assign n5012 = ~n412 & ~n461;
  assign n5013 = ~n552 & n5012;
  assign n5014 = n5010 & n5011;
  assign n5015 = n622 & n5014;
  assign n5016 = n4173 & n5013;
  assign n5017 = n5015 & n5016;
  assign n5018 = n2893 & n5017;
  assign n5019 = n763 & n5018;
  assign n5020 = n4902 & n5019;
  assign n5021 = ~n5009 & n5020;
  assign n5022 = n5009 & ~n5020;
  assign n5023 = ~n5021 & ~n5022;
  assign n5024 = n4983 & ~n5002;
  assign n5025 = ~n5023 & ~n5024;
  assign n5026 = n5023 & n5024;
  assign n5027 = ~n5025 & ~n5026;
  assign n5028 = n4989 & n5005;
  assign n5029 = n3762 & ~n5028;
  assign n5030 = n5027 & ~n5029;
  assign n5031 = ~n5027 & n5029;
  assign po19  = n5030 | n5031;
  assign n5033 = ~n5027 & n5028;
  assign n5034 = n3762 & ~n5033;
  assign n5035 = ~n5022 & ~n5026;
  assign n5036 = ~n378 & n470;
  assign n5037 = n551 & n3399;
  assign n5038 = n4370 & n5037;
  assign n5039 = n4174 & n5036;
  assign n5040 = n5038 & n5039;
  assign n5041 = n527 & n5040;
  assign n5042 = n844 & n5041;
  assign n5043 = n4459 & n5042;
  assign n5044 = ~n5035 & n5043;
  assign n5045 = n5035 & ~n5043;
  assign n5046 = ~n5044 & ~n5045;
  assign n5047 = n5034 & n5046;
  assign n5048 = ~n5034 & ~n5046;
  assign po20  = n5047 | n5048;
  assign n5050 = n5022 & ~n5043;
  assign n5051 = ~n427 & n575;
  assign n5052 = n3361 & n5051;
  assign n5053 = n504 & n5052;
  assign n5054 = ~n5050 & n5053;
  assign n5055 = n5050 & ~n5053;
  assign n5056 = ~n5054 & ~n5055;
  assign n5057 = n5026 & ~n5043;
  assign n5058 = ~n5056 & ~n5057;
  assign n5059 = n5056 & n5057;
  assign n5060 = ~n5058 & ~n5059;
  assign n5061 = n5033 & n5046;
  assign n5062 = n3762 & ~n5061;
  assign n5063 = n5060 & ~n5062;
  assign n5064 = ~n5060 & n5062;
  assign po21  = n5063 | n5064;
  assign n5066 = ~n5060 & n5061;
  assign n5067 = n3762 & ~n5066;
  assign n5068 = n504 & n562;
  assign n5069 = ~n5055 & ~n5059;
  assign n5070 = ~n5068 & ~n5069;
  assign n5071 = n5068 & n5069;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = ~n5067 & n5072;
  assign n5074 = n5067 & ~n5072;
  assign po22  = n5073 | n5074;
  assign n5076 = n5066 & ~n5072;
  assign n5077 = n3762 & ~n5076;
  assign n5078 = n5055 & n5059;
  assign n5079 = n5070 & ~n5078;
  assign n5080 = ~n5077 & n5079;
  assign n5081 = n98 & n103;
  assign n5082 = n5077 & ~n5079;
  assign n5083 = ~n5080 & ~n5081;
  assign po23  = n5082 | ~n5083;
  assign n5085 = ~n5068 & n5078;
  assign n5086 = ~n5076 & ~n5085;
  assign n5087 = n5066 & n5070;
  assign n5088 = ~n5081 & ~n5087;
  assign n5089 = ~n5086 & n5088;
  assign po24  = n3762 & ~n5089;
endmodule
