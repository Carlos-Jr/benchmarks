module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 , pi132 ,
    pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 , pi140 ,
    pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 , pi148 ,
    pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 , pi156 ,
    pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 , pi164 ,
    pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 , pi172 ,
    pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 , pi180 ,
    pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 , pi188 ,
    pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 , pi196 ,
    pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 , pi204 ,
    pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 , pi212 ,
    pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 , pi220 ,
    pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 ,
    po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 ,
    po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 , po30 , po31 , po32 ,
    po33 , po34 , po35 , po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 , po46 , po47 , po48 ,
    po49 , po50 , po51 , po52 , po53 , po54 , po55 , po56 ,
    po57 , po58 , po59 , po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 , po70 , po71 , po72 ,
    po73 , po74 , po75 , po76 , po77 , po78 , po79 , po80 ,
    po81 , po82 , po83 , po84 , po85 , po86 , po87 , po88 ,
    po89 , po90 , po91 , po92 , po93 , po94 , po95 , po96 ,
    po97 , po98 , po99 , po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 , po108 , po109 , po110 ,
    po111 , po112 , po113 , po114 , po115 , po116 , po117 ,
    po118 , po119 , po120 , po121 , po122 , po123 , po124 ,
    po125 , po126 , po127 , po128  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 ,
    pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 ,
    pi140 , pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 ,
    pi148 , pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 ,
    pi156 , pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 ,
    pi164 , pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 ,
    pi172 , pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 ,
    pi180 , pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 ,
    pi188 , pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 ,
    pi196 , pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 ,
    pi204 , pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 ,
    pi212 , pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 ,
    pi220 , pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 , po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 , po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 , po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 , po100 , po101 , po102 ,
    po103 , po104 , po105 , po106 , po107 , po108 , po109 ,
    po110 , po111 , po112 , po113 , po114 , po115 , po116 ,
    po117 , po118 , po119 , po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 , po128;
  wire n386, n387, n389, n390, n391, n392, n393,
    n394, n396, n397, n398, n399, n400, n401,
    n402, n403, n405, n406, n407, n408, n409,
    n410, n411, n413, n414, n415, n416, n417,
    n418, n419, n421, n422, n423, n424, n425,
    n426, n427, n429, n430, n431, n432, n433,
    n434, n435, n437, n438, n439, n440, n441,
    n442, n443, n445, n446, n447, n448, n449,
    n450, n451, n453, n454, n455, n456, n457,
    n458, n459, n461, n462, n463, n464, n465,
    n466, n467, n469, n470, n471, n472, n473,
    n474, n475, n477, n478, n479, n480, n481,
    n482, n483, n485, n486, n487, n488, n489,
    n490, n491, n493, n494, n495, n496, n497,
    n498, n499, n501, n502, n503, n504, n505,
    n506, n507, n509, n510, n511, n512, n513,
    n514, n515, n517, n518, n519, n520, n521,
    n522, n523, n525, n526, n527, n528, n529,
    n530, n531, n533, n534, n535, n536, n537,
    n538, n539, n541, n542, n543, n544, n545,
    n546, n547, n549, n550, n551, n552, n553,
    n554, n555, n557, n558, n559, n560, n561,
    n562, n563, n565, n566, n567, n568, n569,
    n570, n571, n573, n574, n575, n576, n577,
    n578, n579, n581, n582, n583, n584, n585,
    n586, n587, n589, n590, n591, n592, n593,
    n594, n595, n597, n598, n599, n600, n601,
    n602, n603, n605, n606, n607, n608, n609,
    n610, n611, n613, n614, n615, n616, n617,
    n618, n619, n621, n622, n623, n624, n625,
    n626, n627, n629, n630, n631, n632, n633,
    n634, n635, n637, n638, n639, n640, n641,
    n642, n643, n645, n646, n647, n648, n649,
    n650, n651, n653, n654, n655, n656, n657,
    n658, n659, n661, n662, n663, n664, n665,
    n666, n667, n669, n670, n671, n672, n673,
    n674, n675, n677, n678, n679, n680, n681,
    n682, n683, n685, n686, n687, n688, n689,
    n690, n691, n693, n694, n695, n696, n697,
    n698, n699, n701, n702, n703, n704, n705,
    n706, n707, n709, n710, n711, n712, n713,
    n714, n715, n717, n718, n719, n720, n721,
    n722, n723, n725, n726, n727, n728, n729,
    n730, n731, n733, n734, n735, n736, n737,
    n738, n739, n741, n742, n743, n744, n745,
    n746, n747, n749, n750, n751, n752, n753,
    n754, n755, n757, n758, n759, n760, n761,
    n762, n763, n765, n766, n767, n768, n769,
    n770, n771, n773, n774, n775, n776, n777,
    n778, n779, n781, n782, n783, n784, n785,
    n786, n787, n789, n790, n791, n792, n793,
    n794, n795, n797, n798, n799, n800, n801,
    n802, n803, n805, n806, n807, n808, n809,
    n810, n811, n813, n814, n815, n816, n817,
    n818, n819, n821, n822, n823, n824, n825,
    n826, n827, n829, n830, n831, n832, n833,
    n834, n835, n837, n838, n839, n840, n841,
    n842, n843, n845, n846, n847, n848, n849,
    n850, n851, n853, n854, n855, n856, n857,
    n858, n859, n861, n862, n863, n864, n865,
    n866, n867, n869, n870, n871, n872, n873,
    n874, n875, n877, n878, n879, n880, n881,
    n882, n883, n885, n886, n887, n888, n889,
    n890, n891, n893, n894, n895, n896, n897,
    n898, n899, n901, n902, n903, n904, n905,
    n906, n907, n909, n910, n911, n912, n913,
    n914, n915, n917, n918, n919, n920, n921,
    n922, n923, n925, n926, n927, n928, n929,
    n930, n931, n933, n934, n935, n936, n937,
    n938, n939, n941, n942, n943, n944, n945,
    n946, n947, n949, n950, n951, n952, n953,
    n954, n955, n957, n958, n959, n960, n961,
    n962, n963, n965, n966, n967, n968, n969,
    n970, n971, n973, n974, n975, n976, n977,
    n978, n979, n981, n982, n983, n984, n985,
    n986, n987, n989, n990, n991, n992, n993,
    n994, n995, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227,
    n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1237, n1238, n1239, n1240, n1241,
    n1242, n1243, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275,
    n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1349, n1350, n1351,
    n1352, n1353, n1354, n1355, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1397, n1398, n1399,
    n1400, n1401, n1402, n1404;
  assign n386 = pi0  & ~pi128 ;
  assign n387 = ~pi0  & pi128 ;
  assign po0  = n386 | n387;
  assign n389 = pi0  & pi128 ;
  assign n390 = ~pi1  & ~pi129 ;
  assign n391 = pi1  & pi129 ;
  assign n392 = ~n390 & ~n391;
  assign n393 = n389 & ~n392;
  assign n394 = ~n389 & n392;
  assign po1  = n393 | n394;
  assign n396 = ~pi2  & ~pi130 ;
  assign n397 = pi2  & pi130 ;
  assign n398 = ~n396 & ~n397;
  assign n399 = ~n389 & ~n391;
  assign n400 = ~n390 & ~n399;
  assign n401 = ~n398 & n400;
  assign n402 = ~n397 & ~n400;
  assign n403 = ~n396 & n402;
  assign po2  = n401 | n403;
  assign n405 = ~pi3  & ~pi131 ;
  assign n406 = pi3  & pi131 ;
  assign n407 = ~n405 & ~n406;
  assign n408 = ~n396 & ~n402;
  assign n409 = ~n407 & n408;
  assign n410 = ~n406 & ~n408;
  assign n411 = ~n405 & n410;
  assign po3  = n409 | n411;
  assign n413 = ~pi4  & ~pi132 ;
  assign n414 = pi4  & pi132 ;
  assign n415 = ~n413 & ~n414;
  assign n416 = ~n405 & ~n410;
  assign n417 = ~n415 & n416;
  assign n418 = ~n414 & ~n416;
  assign n419 = ~n413 & n418;
  assign po4  = n417 | n419;
  assign n421 = ~pi5  & ~pi133 ;
  assign n422 = pi5  & pi133 ;
  assign n423 = ~n421 & ~n422;
  assign n424 = ~n413 & ~n418;
  assign n425 = ~n423 & n424;
  assign n426 = ~n422 & ~n424;
  assign n427 = ~n421 & n426;
  assign po5  = n425 | n427;
  assign n429 = ~pi6  & ~pi134 ;
  assign n430 = pi6  & pi134 ;
  assign n431 = ~n429 & ~n430;
  assign n432 = ~n421 & ~n426;
  assign n433 = ~n431 & n432;
  assign n434 = ~n430 & ~n432;
  assign n435 = ~n429 & n434;
  assign po6  = n433 | n435;
  assign n437 = ~pi7  & ~pi135 ;
  assign n438 = pi7  & pi135 ;
  assign n439 = ~n437 & ~n438;
  assign n440 = ~n429 & ~n434;
  assign n441 = ~n439 & n440;
  assign n442 = ~n438 & ~n440;
  assign n443 = ~n437 & n442;
  assign po7  = n441 | n443;
  assign n445 = ~pi8  & ~pi136 ;
  assign n446 = pi8  & pi136 ;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~n437 & ~n442;
  assign n449 = ~n447 & n448;
  assign n450 = ~n446 & ~n448;
  assign n451 = ~n445 & n450;
  assign po8  = n449 | n451;
  assign n453 = ~pi9  & ~pi137 ;
  assign n454 = pi9  & pi137 ;
  assign n455 = ~n453 & ~n454;
  assign n456 = ~n445 & ~n450;
  assign n457 = ~n455 & n456;
  assign n458 = ~n454 & ~n456;
  assign n459 = ~n453 & n458;
  assign po9  = n457 | n459;
  assign n461 = ~pi10  & ~pi138 ;
  assign n462 = pi10  & pi138 ;
  assign n463 = ~n461 & ~n462;
  assign n464 = ~n453 & ~n458;
  assign n465 = ~n463 & n464;
  assign n466 = ~n462 & ~n464;
  assign n467 = ~n461 & n466;
  assign po10  = n465 | n467;
  assign n469 = ~pi11  & ~pi139 ;
  assign n470 = pi11  & pi139 ;
  assign n471 = ~n469 & ~n470;
  assign n472 = ~n461 & ~n466;
  assign n473 = ~n471 & n472;
  assign n474 = ~n470 & ~n472;
  assign n475 = ~n469 & n474;
  assign po11  = n473 | n475;
  assign n477 = ~pi12  & ~pi140 ;
  assign n478 = pi12  & pi140 ;
  assign n479 = ~n477 & ~n478;
  assign n480 = ~n469 & ~n474;
  assign n481 = ~n479 & n480;
  assign n482 = ~n478 & ~n480;
  assign n483 = ~n477 & n482;
  assign po12  = n481 | n483;
  assign n485 = ~pi13  & ~pi141 ;
  assign n486 = pi13  & pi141 ;
  assign n487 = ~n485 & ~n486;
  assign n488 = ~n477 & ~n482;
  assign n489 = ~n487 & n488;
  assign n490 = ~n486 & ~n488;
  assign n491 = ~n485 & n490;
  assign po13  = n489 | n491;
  assign n493 = ~pi14  & ~pi142 ;
  assign n494 = pi14  & pi142 ;
  assign n495 = ~n493 & ~n494;
  assign n496 = ~n485 & ~n490;
  assign n497 = ~n495 & n496;
  assign n498 = ~n494 & ~n496;
  assign n499 = ~n493 & n498;
  assign po14  = n497 | n499;
  assign n501 = ~pi15  & ~pi143 ;
  assign n502 = pi15  & pi143 ;
  assign n503 = ~n501 & ~n502;
  assign n504 = ~n493 & ~n498;
  assign n505 = ~n503 & n504;
  assign n506 = ~n502 & ~n504;
  assign n507 = ~n501 & n506;
  assign po15  = n505 | n507;
  assign n509 = ~pi16  & ~pi144 ;
  assign n510 = pi16  & pi144 ;
  assign n511 = ~n509 & ~n510;
  assign n512 = ~n501 & ~n506;
  assign n513 = ~n511 & n512;
  assign n514 = ~n510 & ~n512;
  assign n515 = ~n509 & n514;
  assign po16  = n513 | n515;
  assign n517 = ~pi17  & ~pi145 ;
  assign n518 = pi17  & pi145 ;
  assign n519 = ~n517 & ~n518;
  assign n520 = ~n509 & ~n514;
  assign n521 = ~n519 & n520;
  assign n522 = ~n518 & ~n520;
  assign n523 = ~n517 & n522;
  assign po17  = n521 | n523;
  assign n525 = ~pi18  & ~pi146 ;
  assign n526 = pi18  & pi146 ;
  assign n527 = ~n525 & ~n526;
  assign n528 = ~n517 & ~n522;
  assign n529 = ~n527 & n528;
  assign n530 = ~n526 & ~n528;
  assign n531 = ~n525 & n530;
  assign po18  = n529 | n531;
  assign n533 = ~pi19  & ~pi147 ;
  assign n534 = pi19  & pi147 ;
  assign n535 = ~n533 & ~n534;
  assign n536 = ~n525 & ~n530;
  assign n537 = ~n535 & n536;
  assign n538 = ~n534 & ~n536;
  assign n539 = ~n533 & n538;
  assign po19  = n537 | n539;
  assign n541 = ~pi20  & ~pi148 ;
  assign n542 = pi20  & pi148 ;
  assign n543 = ~n541 & ~n542;
  assign n544 = ~n533 & ~n538;
  assign n545 = ~n543 & n544;
  assign n546 = ~n542 & ~n544;
  assign n547 = ~n541 & n546;
  assign po20  = n545 | n547;
  assign n549 = ~pi21  & ~pi149 ;
  assign n550 = pi21  & pi149 ;
  assign n551 = ~n549 & ~n550;
  assign n552 = ~n541 & ~n546;
  assign n553 = ~n551 & n552;
  assign n554 = ~n550 & ~n552;
  assign n555 = ~n549 & n554;
  assign po21  = n553 | n555;
  assign n557 = ~pi22  & ~pi150 ;
  assign n558 = pi22  & pi150 ;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~n549 & ~n554;
  assign n561 = ~n559 & n560;
  assign n562 = ~n558 & ~n560;
  assign n563 = ~n557 & n562;
  assign po22  = n561 | n563;
  assign n565 = ~pi23  & ~pi151 ;
  assign n566 = pi23  & pi151 ;
  assign n567 = ~n565 & ~n566;
  assign n568 = ~n557 & ~n562;
  assign n569 = ~n567 & n568;
  assign n570 = ~n566 & ~n568;
  assign n571 = ~n565 & n570;
  assign po23  = n569 | n571;
  assign n573 = ~pi24  & ~pi152 ;
  assign n574 = pi24  & pi152 ;
  assign n575 = ~n573 & ~n574;
  assign n576 = ~n565 & ~n570;
  assign n577 = ~n575 & n576;
  assign n578 = ~n574 & ~n576;
  assign n579 = ~n573 & n578;
  assign po24  = n577 | n579;
  assign n581 = ~pi25  & ~pi153 ;
  assign n582 = pi25  & pi153 ;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~n573 & ~n578;
  assign n585 = ~n583 & n584;
  assign n586 = ~n582 & ~n584;
  assign n587 = ~n581 & n586;
  assign po25  = n585 | n587;
  assign n589 = ~pi26  & ~pi154 ;
  assign n590 = pi26  & pi154 ;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~n581 & ~n586;
  assign n593 = ~n591 & n592;
  assign n594 = ~n590 & ~n592;
  assign n595 = ~n589 & n594;
  assign po26  = n593 | n595;
  assign n597 = ~pi27  & ~pi155 ;
  assign n598 = pi27  & pi155 ;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~n589 & ~n594;
  assign n601 = ~n599 & n600;
  assign n602 = ~n598 & ~n600;
  assign n603 = ~n597 & n602;
  assign po27  = n601 | n603;
  assign n605 = ~pi28  & ~pi156 ;
  assign n606 = pi28  & pi156 ;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~n597 & ~n602;
  assign n609 = ~n607 & n608;
  assign n610 = ~n606 & ~n608;
  assign n611 = ~n605 & n610;
  assign po28  = n609 | n611;
  assign n613 = ~pi29  & ~pi157 ;
  assign n614 = pi29  & pi157 ;
  assign n615 = ~n613 & ~n614;
  assign n616 = ~n605 & ~n610;
  assign n617 = ~n615 & n616;
  assign n618 = ~n614 & ~n616;
  assign n619 = ~n613 & n618;
  assign po29  = n617 | n619;
  assign n621 = ~pi30  & ~pi158 ;
  assign n622 = pi30  & pi158 ;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~n613 & ~n618;
  assign n625 = ~n623 & n624;
  assign n626 = ~n622 & ~n624;
  assign n627 = ~n621 & n626;
  assign po30  = n625 | n627;
  assign n629 = ~pi31  & ~pi159 ;
  assign n630 = pi31  & pi159 ;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~n621 & ~n626;
  assign n633 = ~n631 & n632;
  assign n634 = ~n630 & ~n632;
  assign n635 = ~n629 & n634;
  assign po31  = n633 | n635;
  assign n637 = ~pi32  & ~pi160 ;
  assign n638 = pi32  & pi160 ;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~n629 & ~n634;
  assign n641 = ~n639 & n640;
  assign n642 = ~n638 & ~n640;
  assign n643 = ~n637 & n642;
  assign po32  = n641 | n643;
  assign n645 = ~pi33  & ~pi161 ;
  assign n646 = pi33  & pi161 ;
  assign n647 = ~n645 & ~n646;
  assign n648 = ~n637 & ~n642;
  assign n649 = ~n647 & n648;
  assign n650 = ~n646 & ~n648;
  assign n651 = ~n645 & n650;
  assign po33  = n649 | n651;
  assign n653 = ~pi34  & ~pi162 ;
  assign n654 = pi34  & pi162 ;
  assign n655 = ~n653 & ~n654;
  assign n656 = ~n645 & ~n650;
  assign n657 = ~n655 & n656;
  assign n658 = ~n654 & ~n656;
  assign n659 = ~n653 & n658;
  assign po34  = n657 | n659;
  assign n661 = ~pi35  & ~pi163 ;
  assign n662 = pi35  & pi163 ;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~n653 & ~n658;
  assign n665 = ~n663 & n664;
  assign n666 = ~n662 & ~n664;
  assign n667 = ~n661 & n666;
  assign po35  = n665 | n667;
  assign n669 = ~pi36  & ~pi164 ;
  assign n670 = pi36  & pi164 ;
  assign n671 = ~n669 & ~n670;
  assign n672 = ~n661 & ~n666;
  assign n673 = ~n671 & n672;
  assign n674 = ~n670 & ~n672;
  assign n675 = ~n669 & n674;
  assign po36  = n673 | n675;
  assign n677 = ~pi37  & ~pi165 ;
  assign n678 = pi37  & pi165 ;
  assign n679 = ~n677 & ~n678;
  assign n680 = ~n669 & ~n674;
  assign n681 = ~n679 & n680;
  assign n682 = ~n678 & ~n680;
  assign n683 = ~n677 & n682;
  assign po37  = n681 | n683;
  assign n685 = ~pi38  & ~pi166 ;
  assign n686 = pi38  & pi166 ;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~n677 & ~n682;
  assign n689 = ~n687 & n688;
  assign n690 = ~n686 & ~n688;
  assign n691 = ~n685 & n690;
  assign po38  = n689 | n691;
  assign n693 = ~pi39  & ~pi167 ;
  assign n694 = pi39  & pi167 ;
  assign n695 = ~n693 & ~n694;
  assign n696 = ~n685 & ~n690;
  assign n697 = ~n695 & n696;
  assign n698 = ~n694 & ~n696;
  assign n699 = ~n693 & n698;
  assign po39  = n697 | n699;
  assign n701 = ~pi40  & ~pi168 ;
  assign n702 = pi40  & pi168 ;
  assign n703 = ~n701 & ~n702;
  assign n704 = ~n693 & ~n698;
  assign n705 = ~n703 & n704;
  assign n706 = ~n702 & ~n704;
  assign n707 = ~n701 & n706;
  assign po40  = n705 | n707;
  assign n709 = ~pi41  & ~pi169 ;
  assign n710 = pi41  & pi169 ;
  assign n711 = ~n709 & ~n710;
  assign n712 = ~n701 & ~n706;
  assign n713 = ~n711 & n712;
  assign n714 = ~n710 & ~n712;
  assign n715 = ~n709 & n714;
  assign po41  = n713 | n715;
  assign n717 = ~pi42  & ~pi170 ;
  assign n718 = pi42  & pi170 ;
  assign n719 = ~n717 & ~n718;
  assign n720 = ~n709 & ~n714;
  assign n721 = ~n719 & n720;
  assign n722 = ~n718 & ~n720;
  assign n723 = ~n717 & n722;
  assign po42  = n721 | n723;
  assign n725 = ~pi43  & ~pi171 ;
  assign n726 = pi43  & pi171 ;
  assign n727 = ~n725 & ~n726;
  assign n728 = ~n717 & ~n722;
  assign n729 = ~n727 & n728;
  assign n730 = ~n726 & ~n728;
  assign n731 = ~n725 & n730;
  assign po43  = n729 | n731;
  assign n733 = ~pi44  & ~pi172 ;
  assign n734 = pi44  & pi172 ;
  assign n735 = ~n733 & ~n734;
  assign n736 = ~n725 & ~n730;
  assign n737 = ~n735 & n736;
  assign n738 = ~n734 & ~n736;
  assign n739 = ~n733 & n738;
  assign po44  = n737 | n739;
  assign n741 = ~pi45  & ~pi173 ;
  assign n742 = pi45  & pi173 ;
  assign n743 = ~n741 & ~n742;
  assign n744 = ~n733 & ~n738;
  assign n745 = ~n743 & n744;
  assign n746 = ~n742 & ~n744;
  assign n747 = ~n741 & n746;
  assign po45  = n745 | n747;
  assign n749 = ~pi46  & ~pi174 ;
  assign n750 = pi46  & pi174 ;
  assign n751 = ~n749 & ~n750;
  assign n752 = ~n741 & ~n746;
  assign n753 = ~n751 & n752;
  assign n754 = ~n750 & ~n752;
  assign n755 = ~n749 & n754;
  assign po46  = n753 | n755;
  assign n757 = ~pi47  & ~pi175 ;
  assign n758 = pi47  & pi175 ;
  assign n759 = ~n757 & ~n758;
  assign n760 = ~n749 & ~n754;
  assign n761 = ~n759 & n760;
  assign n762 = ~n758 & ~n760;
  assign n763 = ~n757 & n762;
  assign po47  = n761 | n763;
  assign n765 = ~pi48  & ~pi176 ;
  assign n766 = pi48  & pi176 ;
  assign n767 = ~n765 & ~n766;
  assign n768 = ~n757 & ~n762;
  assign n769 = ~n767 & n768;
  assign n770 = ~n766 & ~n768;
  assign n771 = ~n765 & n770;
  assign po48  = n769 | n771;
  assign n773 = ~pi49  & ~pi177 ;
  assign n774 = pi49  & pi177 ;
  assign n775 = ~n773 & ~n774;
  assign n776 = ~n765 & ~n770;
  assign n777 = ~n775 & n776;
  assign n778 = ~n774 & ~n776;
  assign n779 = ~n773 & n778;
  assign po49  = n777 | n779;
  assign n781 = ~pi50  & ~pi178 ;
  assign n782 = pi50  & pi178 ;
  assign n783 = ~n781 & ~n782;
  assign n784 = ~n773 & ~n778;
  assign n785 = ~n783 & n784;
  assign n786 = ~n782 & ~n784;
  assign n787 = ~n781 & n786;
  assign po50  = n785 | n787;
  assign n789 = ~pi51  & ~pi179 ;
  assign n790 = pi51  & pi179 ;
  assign n791 = ~n789 & ~n790;
  assign n792 = ~n781 & ~n786;
  assign n793 = ~n791 & n792;
  assign n794 = ~n790 & ~n792;
  assign n795 = ~n789 & n794;
  assign po51  = n793 | n795;
  assign n797 = ~pi52  & ~pi180 ;
  assign n798 = pi52  & pi180 ;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~n789 & ~n794;
  assign n801 = ~n799 & n800;
  assign n802 = ~n798 & ~n800;
  assign n803 = ~n797 & n802;
  assign po52  = n801 | n803;
  assign n805 = ~pi53  & ~pi181 ;
  assign n806 = pi53  & pi181 ;
  assign n807 = ~n805 & ~n806;
  assign n808 = ~n797 & ~n802;
  assign n809 = ~n807 & n808;
  assign n810 = ~n806 & ~n808;
  assign n811 = ~n805 & n810;
  assign po53  = n809 | n811;
  assign n813 = ~pi54  & ~pi182 ;
  assign n814 = pi54  & pi182 ;
  assign n815 = ~n813 & ~n814;
  assign n816 = ~n805 & ~n810;
  assign n817 = ~n815 & n816;
  assign n818 = ~n814 & ~n816;
  assign n819 = ~n813 & n818;
  assign po54  = n817 | n819;
  assign n821 = ~pi55  & ~pi183 ;
  assign n822 = pi55  & pi183 ;
  assign n823 = ~n821 & ~n822;
  assign n824 = ~n813 & ~n818;
  assign n825 = ~n823 & n824;
  assign n826 = ~n822 & ~n824;
  assign n827 = ~n821 & n826;
  assign po55  = n825 | n827;
  assign n829 = ~pi56  & ~pi184 ;
  assign n830 = pi56  & pi184 ;
  assign n831 = ~n829 & ~n830;
  assign n832 = ~n821 & ~n826;
  assign n833 = ~n831 & n832;
  assign n834 = ~n830 & ~n832;
  assign n835 = ~n829 & n834;
  assign po56  = n833 | n835;
  assign n837 = ~pi57  & ~pi185 ;
  assign n838 = pi57  & pi185 ;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~n829 & ~n834;
  assign n841 = ~n839 & n840;
  assign n842 = ~n838 & ~n840;
  assign n843 = ~n837 & n842;
  assign po57  = n841 | n843;
  assign n845 = ~pi58  & ~pi186 ;
  assign n846 = pi58  & pi186 ;
  assign n847 = ~n845 & ~n846;
  assign n848 = ~n837 & ~n842;
  assign n849 = ~n847 & n848;
  assign n850 = ~n846 & ~n848;
  assign n851 = ~n845 & n850;
  assign po58  = n849 | n851;
  assign n853 = ~pi59  & ~pi187 ;
  assign n854 = pi59  & pi187 ;
  assign n855 = ~n853 & ~n854;
  assign n856 = ~n845 & ~n850;
  assign n857 = ~n855 & n856;
  assign n858 = ~n854 & ~n856;
  assign n859 = ~n853 & n858;
  assign po59  = n857 | n859;
  assign n861 = ~pi60  & ~pi188 ;
  assign n862 = pi60  & pi188 ;
  assign n863 = ~n861 & ~n862;
  assign n864 = ~n853 & ~n858;
  assign n865 = ~n863 & n864;
  assign n866 = ~n862 & ~n864;
  assign n867 = ~n861 & n866;
  assign po60  = n865 | n867;
  assign n869 = ~pi61  & ~pi189 ;
  assign n870 = pi61  & pi189 ;
  assign n871 = ~n869 & ~n870;
  assign n872 = ~n861 & ~n866;
  assign n873 = ~n871 & n872;
  assign n874 = ~n870 & ~n872;
  assign n875 = ~n869 & n874;
  assign po61  = n873 | n875;
  assign n877 = ~pi62  & ~pi190 ;
  assign n878 = pi62  & pi190 ;
  assign n879 = ~n877 & ~n878;
  assign n880 = ~n869 & ~n874;
  assign n881 = ~n879 & n880;
  assign n882 = ~n878 & ~n880;
  assign n883 = ~n877 & n882;
  assign po62  = n881 | n883;
  assign n885 = ~pi63  & ~pi191 ;
  assign n886 = pi63  & pi191 ;
  assign n887 = ~n885 & ~n886;
  assign n888 = ~n877 & ~n882;
  assign n889 = ~n887 & n888;
  assign n890 = ~n886 & ~n888;
  assign n891 = ~n885 & n890;
  assign po63  = n889 | n891;
  assign n893 = ~pi64  & ~pi192 ;
  assign n894 = pi64  & pi192 ;
  assign n895 = ~n893 & ~n894;
  assign n896 = ~n885 & ~n890;
  assign n897 = ~n895 & n896;
  assign n898 = ~n894 & ~n896;
  assign n899 = ~n893 & n898;
  assign po64  = n897 | n899;
  assign n901 = ~pi65  & ~pi193 ;
  assign n902 = pi65  & pi193 ;
  assign n903 = ~n901 & ~n902;
  assign n904 = ~n893 & ~n898;
  assign n905 = ~n903 & n904;
  assign n906 = ~n902 & ~n904;
  assign n907 = ~n901 & n906;
  assign po65  = n905 | n907;
  assign n909 = ~pi66  & ~pi194 ;
  assign n910 = pi66  & pi194 ;
  assign n911 = ~n909 & ~n910;
  assign n912 = ~n901 & ~n906;
  assign n913 = ~n911 & n912;
  assign n914 = ~n910 & ~n912;
  assign n915 = ~n909 & n914;
  assign po66  = n913 | n915;
  assign n917 = ~pi67  & ~pi195 ;
  assign n918 = pi67  & pi195 ;
  assign n919 = ~n917 & ~n918;
  assign n920 = ~n909 & ~n914;
  assign n921 = ~n919 & n920;
  assign n922 = ~n918 & ~n920;
  assign n923 = ~n917 & n922;
  assign po67  = n921 | n923;
  assign n925 = ~pi68  & ~pi196 ;
  assign n926 = pi68  & pi196 ;
  assign n927 = ~n925 & ~n926;
  assign n928 = ~n917 & ~n922;
  assign n929 = ~n927 & n928;
  assign n930 = ~n926 & ~n928;
  assign n931 = ~n925 & n930;
  assign po68  = n929 | n931;
  assign n933 = ~pi69  & ~pi197 ;
  assign n934 = pi69  & pi197 ;
  assign n935 = ~n933 & ~n934;
  assign n936 = ~n925 & ~n930;
  assign n937 = ~n935 & n936;
  assign n938 = ~n934 & ~n936;
  assign n939 = ~n933 & n938;
  assign po69  = n937 | n939;
  assign n941 = ~pi70  & ~pi198 ;
  assign n942 = pi70  & pi198 ;
  assign n943 = ~n941 & ~n942;
  assign n944 = ~n933 & ~n938;
  assign n945 = ~n943 & n944;
  assign n946 = ~n942 & ~n944;
  assign n947 = ~n941 & n946;
  assign po70  = n945 | n947;
  assign n949 = ~pi71  & ~pi199 ;
  assign n950 = pi71  & pi199 ;
  assign n951 = ~n949 & ~n950;
  assign n952 = ~n941 & ~n946;
  assign n953 = ~n951 & n952;
  assign n954 = ~n950 & ~n952;
  assign n955 = ~n949 & n954;
  assign po71  = n953 | n955;
  assign n957 = ~pi72  & ~pi200 ;
  assign n958 = pi72  & pi200 ;
  assign n959 = ~n957 & ~n958;
  assign n960 = ~n949 & ~n954;
  assign n961 = ~n959 & n960;
  assign n962 = ~n958 & ~n960;
  assign n963 = ~n957 & n962;
  assign po72  = n961 | n963;
  assign n965 = ~pi73  & ~pi201 ;
  assign n966 = pi73  & pi201 ;
  assign n967 = ~n965 & ~n966;
  assign n968 = ~n957 & ~n962;
  assign n969 = ~n967 & n968;
  assign n970 = ~n966 & ~n968;
  assign n971 = ~n965 & n970;
  assign po73  = n969 | n971;
  assign n973 = ~pi74  & ~pi202 ;
  assign n974 = pi74  & pi202 ;
  assign n975 = ~n973 & ~n974;
  assign n976 = ~n965 & ~n970;
  assign n977 = ~n975 & n976;
  assign n978 = ~n974 & ~n976;
  assign n979 = ~n973 & n978;
  assign po74  = n977 | n979;
  assign n981 = ~pi75  & ~pi203 ;
  assign n982 = pi75  & pi203 ;
  assign n983 = ~n981 & ~n982;
  assign n984 = ~n973 & ~n978;
  assign n985 = ~n983 & n984;
  assign n986 = ~n982 & ~n984;
  assign n987 = ~n981 & n986;
  assign po75  = n985 | n987;
  assign n989 = ~pi76  & ~pi204 ;
  assign n990 = pi76  & pi204 ;
  assign n991 = ~n989 & ~n990;
  assign n992 = ~n981 & ~n986;
  assign n993 = ~n991 & n992;
  assign n994 = ~n990 & ~n992;
  assign n995 = ~n989 & n994;
  assign po76  = n993 | n995;
  assign n997 = ~pi77  & ~pi205 ;
  assign n998 = pi77  & pi205 ;
  assign n999 = ~n997 & ~n998;
  assign n1000 = ~n989 & ~n994;
  assign n1001 = ~n999 & n1000;
  assign n1002 = ~n998 & ~n1000;
  assign n1003 = ~n997 & n1002;
  assign po77  = n1001 | n1003;
  assign n1005 = ~pi78  & ~pi206 ;
  assign n1006 = pi78  & pi206 ;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = ~n997 & ~n1002;
  assign n1009 = ~n1007 & n1008;
  assign n1010 = ~n1006 & ~n1008;
  assign n1011 = ~n1005 & n1010;
  assign po78  = n1009 | n1011;
  assign n1013 = ~pi79  & ~pi207 ;
  assign n1014 = pi79  & pi207 ;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = ~n1005 & ~n1010;
  assign n1017 = ~n1015 & n1016;
  assign n1018 = ~n1014 & ~n1016;
  assign n1019 = ~n1013 & n1018;
  assign po79  = n1017 | n1019;
  assign n1021 = ~pi80  & ~pi208 ;
  assign n1022 = pi80  & pi208 ;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = ~n1013 & ~n1018;
  assign n1025 = ~n1023 & n1024;
  assign n1026 = ~n1022 & ~n1024;
  assign n1027 = ~n1021 & n1026;
  assign po80  = n1025 | n1027;
  assign n1029 = ~pi81  & ~pi209 ;
  assign n1030 = pi81  & pi209 ;
  assign n1031 = ~n1029 & ~n1030;
  assign n1032 = ~n1021 & ~n1026;
  assign n1033 = ~n1031 & n1032;
  assign n1034 = ~n1030 & ~n1032;
  assign n1035 = ~n1029 & n1034;
  assign po81  = n1033 | n1035;
  assign n1037 = ~pi82  & ~pi210 ;
  assign n1038 = pi82  & pi210 ;
  assign n1039 = ~n1037 & ~n1038;
  assign n1040 = ~n1029 & ~n1034;
  assign n1041 = ~n1039 & n1040;
  assign n1042 = ~n1038 & ~n1040;
  assign n1043 = ~n1037 & n1042;
  assign po82  = n1041 | n1043;
  assign n1045 = ~pi83  & ~pi211 ;
  assign n1046 = pi83  & pi211 ;
  assign n1047 = ~n1045 & ~n1046;
  assign n1048 = ~n1037 & ~n1042;
  assign n1049 = ~n1047 & n1048;
  assign n1050 = ~n1046 & ~n1048;
  assign n1051 = ~n1045 & n1050;
  assign po83  = n1049 | n1051;
  assign n1053 = ~pi84  & ~pi212 ;
  assign n1054 = pi84  & pi212 ;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = ~n1045 & ~n1050;
  assign n1057 = ~n1055 & n1056;
  assign n1058 = ~n1054 & ~n1056;
  assign n1059 = ~n1053 & n1058;
  assign po84  = n1057 | n1059;
  assign n1061 = ~pi85  & ~pi213 ;
  assign n1062 = pi85  & pi213 ;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = ~n1053 & ~n1058;
  assign n1065 = ~n1063 & n1064;
  assign n1066 = ~n1062 & ~n1064;
  assign n1067 = ~n1061 & n1066;
  assign po85  = n1065 | n1067;
  assign n1069 = ~pi86  & ~pi214 ;
  assign n1070 = pi86  & pi214 ;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = ~n1061 & ~n1066;
  assign n1073 = ~n1071 & n1072;
  assign n1074 = ~n1070 & ~n1072;
  assign n1075 = ~n1069 & n1074;
  assign po86  = n1073 | n1075;
  assign n1077 = ~pi87  & ~pi215 ;
  assign n1078 = pi87  & pi215 ;
  assign n1079 = ~n1077 & ~n1078;
  assign n1080 = ~n1069 & ~n1074;
  assign n1081 = ~n1079 & n1080;
  assign n1082 = ~n1078 & ~n1080;
  assign n1083 = ~n1077 & n1082;
  assign po87  = n1081 | n1083;
  assign n1085 = ~pi88  & ~pi216 ;
  assign n1086 = pi88  & pi216 ;
  assign n1087 = ~n1085 & ~n1086;
  assign n1088 = ~n1077 & ~n1082;
  assign n1089 = ~n1087 & n1088;
  assign n1090 = ~n1086 & ~n1088;
  assign n1091 = ~n1085 & n1090;
  assign po88  = n1089 | n1091;
  assign n1093 = ~pi89  & ~pi217 ;
  assign n1094 = pi89  & pi217 ;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = ~n1085 & ~n1090;
  assign n1097 = ~n1095 & n1096;
  assign n1098 = ~n1094 & ~n1096;
  assign n1099 = ~n1093 & n1098;
  assign po89  = n1097 | n1099;
  assign n1101 = ~pi90  & ~pi218 ;
  assign n1102 = pi90  & pi218 ;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = ~n1093 & ~n1098;
  assign n1105 = ~n1103 & n1104;
  assign n1106 = ~n1102 & ~n1104;
  assign n1107 = ~n1101 & n1106;
  assign po90  = n1105 | n1107;
  assign n1109 = ~pi91  & ~pi219 ;
  assign n1110 = pi91  & pi219 ;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = ~n1101 & ~n1106;
  assign n1113 = ~n1111 & n1112;
  assign n1114 = ~n1110 & ~n1112;
  assign n1115 = ~n1109 & n1114;
  assign po91  = n1113 | n1115;
  assign n1117 = ~pi92  & ~pi220 ;
  assign n1118 = pi92  & pi220 ;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = ~n1109 & ~n1114;
  assign n1121 = ~n1119 & n1120;
  assign n1122 = ~n1118 & ~n1120;
  assign n1123 = ~n1117 & n1122;
  assign po92  = n1121 | n1123;
  assign n1125 = ~pi93  & ~pi221 ;
  assign n1126 = pi93  & pi221 ;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = ~n1117 & ~n1122;
  assign n1129 = ~n1127 & n1128;
  assign n1130 = ~n1126 & ~n1128;
  assign n1131 = ~n1125 & n1130;
  assign po93  = n1129 | n1131;
  assign n1133 = ~pi94  & ~pi222 ;
  assign n1134 = pi94  & pi222 ;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = ~n1125 & ~n1130;
  assign n1137 = ~n1135 & n1136;
  assign n1138 = ~n1134 & ~n1136;
  assign n1139 = ~n1133 & n1138;
  assign po94  = n1137 | n1139;
  assign n1141 = ~pi95  & ~pi223 ;
  assign n1142 = pi95  & pi223 ;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n1133 & ~n1138;
  assign n1145 = ~n1143 & n1144;
  assign n1146 = ~n1142 & ~n1144;
  assign n1147 = ~n1141 & n1146;
  assign po95  = n1145 | n1147;
  assign n1149 = ~pi96  & ~pi224 ;
  assign n1150 = pi96  & pi224 ;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = ~n1141 & ~n1146;
  assign n1153 = ~n1151 & n1152;
  assign n1154 = ~n1150 & ~n1152;
  assign n1155 = ~n1149 & n1154;
  assign po96  = n1153 | n1155;
  assign n1157 = ~pi97  & ~pi225 ;
  assign n1158 = pi97  & pi225 ;
  assign n1159 = ~n1157 & ~n1158;
  assign n1160 = ~n1149 & ~n1154;
  assign n1161 = ~n1159 & n1160;
  assign n1162 = ~n1158 & ~n1160;
  assign n1163 = ~n1157 & n1162;
  assign po97  = n1161 | n1163;
  assign n1165 = ~pi98  & ~pi226 ;
  assign n1166 = pi98  & pi226 ;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = ~n1157 & ~n1162;
  assign n1169 = ~n1167 & n1168;
  assign n1170 = ~n1166 & ~n1168;
  assign n1171 = ~n1165 & n1170;
  assign po98  = n1169 | n1171;
  assign n1173 = ~pi99  & ~pi227 ;
  assign n1174 = pi99  & pi227 ;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = ~n1165 & ~n1170;
  assign n1177 = ~n1175 & n1176;
  assign n1178 = ~n1174 & ~n1176;
  assign n1179 = ~n1173 & n1178;
  assign po99  = n1177 | n1179;
  assign n1181 = ~pi100  & ~pi228 ;
  assign n1182 = pi100  & pi228 ;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = ~n1173 & ~n1178;
  assign n1185 = ~n1183 & n1184;
  assign n1186 = ~n1182 & ~n1184;
  assign n1187 = ~n1181 & n1186;
  assign po100  = n1185 | n1187;
  assign n1189 = ~pi101  & ~pi229 ;
  assign n1190 = pi101  & pi229 ;
  assign n1191 = ~n1189 & ~n1190;
  assign n1192 = ~n1181 & ~n1186;
  assign n1193 = ~n1191 & n1192;
  assign n1194 = ~n1190 & ~n1192;
  assign n1195 = ~n1189 & n1194;
  assign po101  = n1193 | n1195;
  assign n1197 = ~pi102  & ~pi230 ;
  assign n1198 = pi102  & pi230 ;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = ~n1189 & ~n1194;
  assign n1201 = ~n1199 & n1200;
  assign n1202 = ~n1198 & ~n1200;
  assign n1203 = ~n1197 & n1202;
  assign po102  = n1201 | n1203;
  assign n1205 = ~pi103  & ~pi231 ;
  assign n1206 = pi103  & pi231 ;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = ~n1197 & ~n1202;
  assign n1209 = ~n1207 & n1208;
  assign n1210 = ~n1206 & ~n1208;
  assign n1211 = ~n1205 & n1210;
  assign po103  = n1209 | n1211;
  assign n1213 = ~pi104  & ~pi232 ;
  assign n1214 = pi104  & pi232 ;
  assign n1215 = ~n1213 & ~n1214;
  assign n1216 = ~n1205 & ~n1210;
  assign n1217 = ~n1215 & n1216;
  assign n1218 = ~n1214 & ~n1216;
  assign n1219 = ~n1213 & n1218;
  assign po104  = n1217 | n1219;
  assign n1221 = ~pi105  & ~pi233 ;
  assign n1222 = pi105  & pi233 ;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = ~n1213 & ~n1218;
  assign n1225 = ~n1223 & n1224;
  assign n1226 = ~n1222 & ~n1224;
  assign n1227 = ~n1221 & n1226;
  assign po105  = n1225 | n1227;
  assign n1229 = ~pi106  & ~pi234 ;
  assign n1230 = pi106  & pi234 ;
  assign n1231 = ~n1229 & ~n1230;
  assign n1232 = ~n1221 & ~n1226;
  assign n1233 = ~n1231 & n1232;
  assign n1234 = ~n1230 & ~n1232;
  assign n1235 = ~n1229 & n1234;
  assign po106  = n1233 | n1235;
  assign n1237 = ~pi107  & ~pi235 ;
  assign n1238 = pi107  & pi235 ;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = ~n1229 & ~n1234;
  assign n1241 = ~n1239 & n1240;
  assign n1242 = ~n1238 & ~n1240;
  assign n1243 = ~n1237 & n1242;
  assign po107  = n1241 | n1243;
  assign n1245 = ~pi108  & ~pi236 ;
  assign n1246 = pi108  & pi236 ;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = ~n1237 & ~n1242;
  assign n1249 = ~n1247 & n1248;
  assign n1250 = ~n1246 & ~n1248;
  assign n1251 = ~n1245 & n1250;
  assign po108  = n1249 | n1251;
  assign n1253 = ~pi109  & ~pi237 ;
  assign n1254 = pi109  & pi237 ;
  assign n1255 = ~n1253 & ~n1254;
  assign n1256 = ~n1245 & ~n1250;
  assign n1257 = ~n1255 & n1256;
  assign n1258 = ~n1254 & ~n1256;
  assign n1259 = ~n1253 & n1258;
  assign po109  = n1257 | n1259;
  assign n1261 = ~pi110  & ~pi238 ;
  assign n1262 = pi110  & pi238 ;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = ~n1253 & ~n1258;
  assign n1265 = ~n1263 & n1264;
  assign n1266 = ~n1262 & ~n1264;
  assign n1267 = ~n1261 & n1266;
  assign po110  = n1265 | n1267;
  assign n1269 = ~pi111  & ~pi239 ;
  assign n1270 = pi111  & pi239 ;
  assign n1271 = ~n1269 & ~n1270;
  assign n1272 = ~n1261 & ~n1266;
  assign n1273 = ~n1271 & n1272;
  assign n1274 = ~n1270 & ~n1272;
  assign n1275 = ~n1269 & n1274;
  assign po111  = n1273 | n1275;
  assign n1277 = ~pi112  & ~pi240 ;
  assign n1278 = pi112  & pi240 ;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = ~n1269 & ~n1274;
  assign n1281 = ~n1279 & n1280;
  assign n1282 = ~n1278 & ~n1280;
  assign n1283 = ~n1277 & n1282;
  assign po112  = n1281 | n1283;
  assign n1285 = ~pi113  & ~pi241 ;
  assign n1286 = pi113  & pi241 ;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = ~n1277 & ~n1282;
  assign n1289 = ~n1287 & n1288;
  assign n1290 = ~n1286 & ~n1288;
  assign n1291 = ~n1285 & n1290;
  assign po113  = n1289 | n1291;
  assign n1293 = ~pi114  & ~pi242 ;
  assign n1294 = pi114  & pi242 ;
  assign n1295 = ~n1293 & ~n1294;
  assign n1296 = ~n1285 & ~n1290;
  assign n1297 = ~n1295 & n1296;
  assign n1298 = ~n1294 & ~n1296;
  assign n1299 = ~n1293 & n1298;
  assign po114  = n1297 | n1299;
  assign n1301 = ~pi115  & ~pi243 ;
  assign n1302 = pi115  & pi243 ;
  assign n1303 = ~n1301 & ~n1302;
  assign n1304 = ~n1293 & ~n1298;
  assign n1305 = ~n1303 & n1304;
  assign n1306 = ~n1302 & ~n1304;
  assign n1307 = ~n1301 & n1306;
  assign po115  = n1305 | n1307;
  assign n1309 = ~pi116  & ~pi244 ;
  assign n1310 = pi116  & pi244 ;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = ~n1301 & ~n1306;
  assign n1313 = ~n1311 & n1312;
  assign n1314 = ~n1310 & ~n1312;
  assign n1315 = ~n1309 & n1314;
  assign po116  = n1313 | n1315;
  assign n1317 = ~pi117  & ~pi245 ;
  assign n1318 = pi117  & pi245 ;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = ~n1309 & ~n1314;
  assign n1321 = ~n1319 & n1320;
  assign n1322 = ~n1318 & ~n1320;
  assign n1323 = ~n1317 & n1322;
  assign po117  = n1321 | n1323;
  assign n1325 = ~pi118  & ~pi246 ;
  assign n1326 = pi118  & pi246 ;
  assign n1327 = ~n1325 & ~n1326;
  assign n1328 = ~n1317 & ~n1322;
  assign n1329 = ~n1327 & n1328;
  assign n1330 = ~n1326 & ~n1328;
  assign n1331 = ~n1325 & n1330;
  assign po118  = n1329 | n1331;
  assign n1333 = ~pi119  & ~pi247 ;
  assign n1334 = pi119  & pi247 ;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = ~n1325 & ~n1330;
  assign n1337 = ~n1335 & n1336;
  assign n1338 = ~n1334 & ~n1336;
  assign n1339 = ~n1333 & n1338;
  assign po119  = n1337 | n1339;
  assign n1341 = ~pi120  & ~pi248 ;
  assign n1342 = pi120  & pi248 ;
  assign n1343 = ~n1341 & ~n1342;
  assign n1344 = ~n1333 & ~n1338;
  assign n1345 = ~n1343 & n1344;
  assign n1346 = ~n1342 & ~n1344;
  assign n1347 = ~n1341 & n1346;
  assign po120  = n1345 | n1347;
  assign n1349 = ~pi121  & ~pi249 ;
  assign n1350 = pi121  & pi249 ;
  assign n1351 = ~n1349 & ~n1350;
  assign n1352 = ~n1341 & ~n1346;
  assign n1353 = ~n1351 & n1352;
  assign n1354 = ~n1350 & ~n1352;
  assign n1355 = ~n1349 & n1354;
  assign po121  = n1353 | n1355;
  assign n1357 = ~pi122  & ~pi250 ;
  assign n1358 = pi122  & pi250 ;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = ~n1349 & ~n1354;
  assign n1361 = ~n1359 & n1360;
  assign n1362 = ~n1358 & ~n1360;
  assign n1363 = ~n1357 & n1362;
  assign po122  = n1361 | n1363;
  assign n1365 = ~pi123  & ~pi251 ;
  assign n1366 = pi123  & pi251 ;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = ~n1357 & ~n1362;
  assign n1369 = ~n1367 & n1368;
  assign n1370 = ~n1366 & ~n1368;
  assign n1371 = ~n1365 & n1370;
  assign po123  = n1369 | n1371;
  assign n1373 = ~pi124  & ~pi252 ;
  assign n1374 = pi124  & pi252 ;
  assign n1375 = ~n1373 & ~n1374;
  assign n1376 = ~n1365 & ~n1370;
  assign n1377 = ~n1375 & n1376;
  assign n1378 = ~n1374 & ~n1376;
  assign n1379 = ~n1373 & n1378;
  assign po124  = n1377 | n1379;
  assign n1381 = ~pi125  & ~pi253 ;
  assign n1382 = pi125  & pi253 ;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = ~n1373 & ~n1378;
  assign n1385 = ~n1383 & n1384;
  assign n1386 = ~n1382 & ~n1384;
  assign n1387 = ~n1381 & n1386;
  assign po125  = n1385 | n1387;
  assign n1389 = ~pi126  & ~pi254 ;
  assign n1390 = pi126  & pi254 ;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = ~n1381 & ~n1386;
  assign n1393 = ~n1391 & n1392;
  assign n1394 = ~n1390 & ~n1392;
  assign n1395 = ~n1389 & n1394;
  assign po126  = n1393 | n1395;
  assign n1397 = ~pi127  & ~pi255 ;
  assign n1398 = pi127  & pi255 ;
  assign n1399 = ~n1397 & ~n1398;
  assign n1400 = ~n1389 & ~n1394;
  assign n1401 = n1399 & ~n1400;
  assign n1402 = ~n1399 & n1400;
  assign po127  = n1401 | n1402;
  assign n1404 = ~n1398 & ~n1400;
  assign po128 = ~n1397 & ~n1404;
endmodule
