module dec ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 ,
    pi6 , pi7 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 ,
    po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 ,
    po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 ,
    po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 ,
    po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 ,
    po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 ,
    po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 ,
    po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 ,
    po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 ,
    po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ,
    po128 , po129 , po130 , po131 ,
    po132 , po133 , po134 , po135 ,
    po136 , po137 , po138 , po139 ,
    po140 , po141 , po142 , po143 ,
    po144 , po145 , po146 , po147 ,
    po148 , po149 , po150 , po151 ,
    po152 , po153 , po154 , po155 ,
    po156 , po157 , po158 , po159 ,
    po160 , po161 , po162 , po163 ,
    po164 , po165 , po166 , po167 ,
    po168 , po169 , po170 , po171 ,
    po172 , po173 , po174 , po175 ,
    po176 , po177 , po178 , po179 ,
    po180 , po181 , po182 , po183 ,
    po184 , po185 , po186 , po187 ,
    po188 , po189 , po190 , po191 ,
    po192 , po193 , po194 , po195 ,
    po196 , po197 , po198 , po199 ,
    po200 , po201 , po202 , po203 ,
    po204 , po205 , po206 , po207 ,
    po208 , po209 , po210 , po211 ,
    po212 , po213 , po214 , po215 ,
    po216 , po217 , po218 , po219 ,
    po220 , po221 , po222 , po223 ,
    po224 , po225 , po226 , po227 ,
    po228 , po229 , po230 , po231 ,
    po232 , po233 , po234 , po235 ,
    po236 , po237 , po238 , po239 ,
    po240 , po241 , po242 , po243 ,
    po244 , po245 , po246 , po247 ,
    po248 , po249 , po250 , po251 ,
    po252 , po253 , po254 , po255   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 ;
  output po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 ,
    po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 ,
    po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 ,
    po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 ,
    po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 ,
    po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 ,
    po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 ,
    po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 ,
    po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 ,
    po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ,
    po128 , po129 , po130 , po131 ,
    po132 , po133 , po134 , po135 ,
    po136 , po137 , po138 , po139 ,
    po140 , po141 , po142 , po143 ,
    po144 , po145 , po146 , po147 ,
    po148 , po149 , po150 , po151 ,
    po152 , po153 , po154 , po155 ,
    po156 , po157 , po158 , po159 ,
    po160 , po161 , po162 , po163 ,
    po164 , po165 , po166 , po167 ,
    po168 , po169 , po170 , po171 ,
    po172 , po173 , po174 , po175 ,
    po176 , po177 , po178 , po179 ,
    po180 , po181 , po182 , po183 ,
    po184 , po185 , po186 , po187 ,
    po188 , po189 , po190 , po191 ,
    po192 , po193 , po194 , po195 ,
    po196 , po197 , po198 , po199 ,
    po200 , po201 , po202 , po203 ,
    po204 , po205 , po206 , po207 ,
    po208 , po209 , po210 , po211 ,
    po212 , po213 , po214 , po215 ,
    po216 , po217 , po218 , po219 ,
    po220 , po221 , po222 , po223 ,
    po224 , po225 , po226 , po227 ,
    po228 , po229 , po230 , po231 ,
    po232 , po233 , po234 , po235 ,
    po236 , po237 , po238 , po239 ,
    po240 , po241 , po242 , po243 ,
    po244 , po245 , po246 , po247 ,
    po248 , po249 , po250 , po251 ,
    po252 , po253 , po254 , po255 ;
  wire n265, n266, n267, n268, n269, n270, n272,
    n273, n275, n276, n278, n280, n281, n283,
    n284, n286, n288, n290, n291, n293, n295,
    n296, n298, n300, n302, n304, n306, n308,
    n309, n326, n327, n344, n345, n362, n363,
    n380, n397, n414, n431, n432, n449, n466,
    n483, n500, n501, n518, n535, n552;
  assign n265 = ~pi4  & ~pi5 ;
  assign n266 = ~pi6  & pi7 ;
  assign n267 = n265 & n266;
  assign n268 = ~pi0  & ~pi2 ;
  assign n269 = ~pi1  & ~pi3 ;
  assign n270 = n268 & n269;
  assign po0  = n267 & n270;
  assign n272 = pi0  & ~pi2 ;
  assign n273 = n269 & n272;
  assign po1  = n267 & n273;
  assign n275 = pi1  & ~pi3 ;
  assign n276 = n268 & n275;
  assign po2  = n267 & n276;
  assign n278 = n272 & n275;
  assign po3  = n267 & n278;
  assign n280 = ~pi0  & pi2 ;
  assign n281 = n269 & n280;
  assign po4  = n267 & n281;
  assign n283 = pi0  & pi2 ;
  assign n284 = n269 & n283;
  assign po5  = n267 & n284;
  assign n286 = n275 & n280;
  assign po6  = n267 & n286;
  assign n288 = n275 & n283;
  assign po7  = n267 & n288;
  assign n290 = ~pi1  & pi3 ;
  assign n291 = n268 & n290;
  assign po8  = n267 & n291;
  assign n293 = n272 & n290;
  assign po9  = n267 & n293;
  assign n295 = pi1  & pi3 ;
  assign n296 = n268 & n295;
  assign po10  = n267 & n296;
  assign n298 = n272 & n295;
  assign po11  = n267 & n298;
  assign n300 = n280 & n290;
  assign po12  = n267 & n300;
  assign n302 = n283 & n290;
  assign po13  = n267 & n302;
  assign n304 = n280 & n295;
  assign po14  = n267 & n304;
  assign n306 = n283 & n295;
  assign po15  = n267 & n306;
  assign n308 = pi4  & ~pi5 ;
  assign n309 = n266 & n308;
  assign po16  = n270 & n309;
  assign po17  = n273 & n309;
  assign po18  = n276 & n309;
  assign po19  = n278 & n309;
  assign po20  = n281 & n309;
  assign po21  = n284 & n309;
  assign po22  = n286 & n309;
  assign po23  = n288 & n309;
  assign po24  = n291 & n309;
  assign po25  = n293 & n309;
  assign po26  = n296 & n309;
  assign po27  = n298 & n309;
  assign po28  = n300 & n309;
  assign po29  = n302 & n309;
  assign po30  = n304 & n309;
  assign po31  = n306 & n309;
  assign n326 = ~pi4  & pi5 ;
  assign n327 = n266 & n326;
  assign po32  = n270 & n327;
  assign po33  = n273 & n327;
  assign po34  = n276 & n327;
  assign po35  = n278 & n327;
  assign po36  = n281 & n327;
  assign po37  = n284 & n327;
  assign po38  = n286 & n327;
  assign po39  = n288 & n327;
  assign po40  = n291 & n327;
  assign po41  = n293 & n327;
  assign po42  = n296 & n327;
  assign po43  = n298 & n327;
  assign po44  = n300 & n327;
  assign po45  = n302 & n327;
  assign po46  = n304 & n327;
  assign po47  = n306 & n327;
  assign n344 = pi4  & pi5 ;
  assign n345 = n266 & n344;
  assign po48  = n270 & n345;
  assign po49  = n273 & n345;
  assign po50  = n276 & n345;
  assign po51  = n278 & n345;
  assign po52  = n281 & n345;
  assign po53  = n284 & n345;
  assign po54  = n286 & n345;
  assign po55  = n288 & n345;
  assign po56  = n291 & n345;
  assign po57  = n293 & n345;
  assign po58  = n296 & n345;
  assign po59  = n298 & n345;
  assign po60  = n300 & n345;
  assign po61  = n302 & n345;
  assign po62  = n304 & n345;
  assign po63  = n306 & n345;
  assign n362 = pi6  & pi7 ;
  assign n363 = n265 & n362;
  assign po64  = n270 & n363;
  assign po65  = n273 & n363;
  assign po66  = n276 & n363;
  assign po67  = n278 & n363;
  assign po68  = n281 & n363;
  assign po69  = n284 & n363;
  assign po70  = n286 & n363;
  assign po71  = n288 & n363;
  assign po72  = n291 & n363;
  assign po73  = n293 & n363;
  assign po74  = n296 & n363;
  assign po75  = n298 & n363;
  assign po76  = n300 & n363;
  assign po77  = n302 & n363;
  assign po78  = n304 & n363;
  assign po79  = n306 & n363;
  assign n380 = n308 & n362;
  assign po80  = n270 & n380;
  assign po81  = n273 & n380;
  assign po82  = n276 & n380;
  assign po83  = n278 & n380;
  assign po84  = n281 & n380;
  assign po85  = n284 & n380;
  assign po86  = n286 & n380;
  assign po87  = n288 & n380;
  assign po88  = n291 & n380;
  assign po89  = n293 & n380;
  assign po90  = n296 & n380;
  assign po91  = n298 & n380;
  assign po92  = n300 & n380;
  assign po93  = n302 & n380;
  assign po94  = n304 & n380;
  assign po95  = n306 & n380;
  assign n397 = n326 & n362;
  assign po96  = n270 & n397;
  assign po97  = n273 & n397;
  assign po98  = n276 & n397;
  assign po99  = n278 & n397;
  assign po100  = n281 & n397;
  assign po101  = n284 & n397;
  assign po102  = n286 & n397;
  assign po103  = n288 & n397;
  assign po104  = n291 & n397;
  assign po105  = n293 & n397;
  assign po106  = n296 & n397;
  assign po107  = n298 & n397;
  assign po108  = n300 & n397;
  assign po109  = n302 & n397;
  assign po110  = n304 & n397;
  assign po111  = n306 & n397;
  assign n414 = n344 & n362;
  assign po112  = n270 & n414;
  assign po113  = n273 & n414;
  assign po114  = n276 & n414;
  assign po115  = n278 & n414;
  assign po116  = n281 & n414;
  assign po117  = n284 & n414;
  assign po118  = n286 & n414;
  assign po119  = n288 & n414;
  assign po120  = n291 & n414;
  assign po121  = n293 & n414;
  assign po122  = n296 & n414;
  assign po123  = n298 & n414;
  assign po124  = n300 & n414;
  assign po125  = n302 & n414;
  assign po126  = n304 & n414;
  assign po127  = n306 & n414;
  assign n431 = ~pi6  & ~pi7 ;
  assign n432 = n265 & n431;
  assign po128  = n270 & n432;
  assign po129  = n273 & n432;
  assign po130  = n276 & n432;
  assign po131  = n278 & n432;
  assign po132  = n281 & n432;
  assign po133  = n284 & n432;
  assign po134  = n286 & n432;
  assign po135  = n288 & n432;
  assign po136  = n291 & n432;
  assign po137  = n293 & n432;
  assign po138  = n296 & n432;
  assign po139  = n298 & n432;
  assign po140  = n300 & n432;
  assign po141  = n302 & n432;
  assign po142  = n304 & n432;
  assign po143  = n306 & n432;
  assign n449 = n308 & n431;
  assign po144  = n270 & n449;
  assign po145  = n273 & n449;
  assign po146  = n276 & n449;
  assign po147  = n278 & n449;
  assign po148  = n281 & n449;
  assign po149  = n284 & n449;
  assign po150  = n286 & n449;
  assign po151  = n288 & n449;
  assign po152  = n291 & n449;
  assign po153  = n293 & n449;
  assign po154  = n296 & n449;
  assign po155  = n298 & n449;
  assign po156  = n300 & n449;
  assign po157  = n302 & n449;
  assign po158  = n304 & n449;
  assign po159  = n306 & n449;
  assign n466 = n326 & n431;
  assign po160  = n270 & n466;
  assign po161  = n273 & n466;
  assign po162  = n276 & n466;
  assign po163  = n278 & n466;
  assign po164  = n281 & n466;
  assign po165  = n284 & n466;
  assign po166  = n286 & n466;
  assign po167  = n288 & n466;
  assign po168  = n291 & n466;
  assign po169  = n293 & n466;
  assign po170  = n296 & n466;
  assign po171  = n298 & n466;
  assign po172  = n300 & n466;
  assign po173  = n302 & n466;
  assign po174  = n304 & n466;
  assign po175  = n306 & n466;
  assign n483 = n344 & n431;
  assign po176  = n270 & n483;
  assign po177  = n273 & n483;
  assign po178  = n276 & n483;
  assign po179  = n278 & n483;
  assign po180  = n281 & n483;
  assign po181  = n284 & n483;
  assign po182  = n286 & n483;
  assign po183  = n288 & n483;
  assign po184  = n291 & n483;
  assign po185  = n293 & n483;
  assign po186  = n296 & n483;
  assign po187  = n298 & n483;
  assign po188  = n300 & n483;
  assign po189  = n302 & n483;
  assign po190  = n304 & n483;
  assign po191  = n306 & n483;
  assign n500 = pi6  & ~pi7 ;
  assign n501 = n265 & n500;
  assign po192  = n270 & n501;
  assign po193  = n273 & n501;
  assign po194  = n276 & n501;
  assign po195  = n278 & n501;
  assign po196  = n281 & n501;
  assign po197  = n284 & n501;
  assign po198  = n286 & n501;
  assign po199  = n288 & n501;
  assign po200  = n291 & n501;
  assign po201  = n293 & n501;
  assign po202  = n296 & n501;
  assign po203  = n298 & n501;
  assign po204  = n300 & n501;
  assign po205  = n302 & n501;
  assign po206  = n304 & n501;
  assign po207  = n306 & n501;
  assign n518 = n308 & n500;
  assign po208  = n270 & n518;
  assign po209  = n273 & n518;
  assign po210  = n276 & n518;
  assign po211  = n278 & n518;
  assign po212  = n281 & n518;
  assign po213  = n284 & n518;
  assign po214  = n286 & n518;
  assign po215  = n288 & n518;
  assign po216  = n291 & n518;
  assign po217  = n293 & n518;
  assign po218  = n296 & n518;
  assign po219  = n298 & n518;
  assign po220  = n300 & n518;
  assign po221  = n302 & n518;
  assign po222  = n304 & n518;
  assign po223  = n306 & n518;
  assign n535 = n326 & n500;
  assign po224  = n270 & n535;
  assign po225  = n273 & n535;
  assign po226  = n276 & n535;
  assign po227  = n278 & n535;
  assign po228  = n281 & n535;
  assign po229  = n284 & n535;
  assign po230  = n286 & n535;
  assign po231  = n288 & n535;
  assign po232  = n291 & n535;
  assign po233  = n293 & n535;
  assign po234  = n296 & n535;
  assign po235  = n298 & n535;
  assign po236  = n300 & n535;
  assign po237  = n302 & n535;
  assign po238  = n304 & n535;
  assign po239  = n306 & n535;
  assign n552 = n344 & n500;
  assign po240  = n270 & n552;
  assign po241  = n273 & n552;
  assign po242  = n276 & n552;
  assign po243  = n278 & n552;
  assign po244  = n281 & n552;
  assign po245  = n284 & n552;
  assign po246  = n286 & n552;
  assign po247  = n288 & n552;
  assign po248  = n291 & n552;
  assign po249  = n293 & n552;
  assign po250  = n296 & n552;
  assign po251  = n298 & n552;
  assign po252  = n300 & n552;
  assign po253  = n302 & n552;
  assign po254  = n304 & n552;
  assign po255  = n306 & n552;
endmodule
