module alu4_cl ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    po0, po1, po2, po3, po4, po5  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9;
  output po0, po1, po2, po3, po4, po5;
  wire n17, n18, n20, n21, n22, n23, n24,
    n25, n26, n27, n28, n29, n30, n31, n32,
    n33, n34, n35, n36, n37, n38, n39, n40,
    n41, n42, n43, n44, n45, n46, n47, n48,
    n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n100, n101, n102, n103,
    n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n630,
    n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715,
    n716, n717, n718, n719, n720, n721, n722,
    n723, n724;
  assign n17 = pi6 & ~pi7;
  assign n18 = ~pi0 & pi2;
  assign po3 = pi1 & pi3;
  assign n20 = n18 & po3;
  assign n21 = ~pi1 & pi3;
  assign n22 = pi5 & ~n18;
  assign n23 = pi5 & n21;
  assign n24 = ~n18 & n23;
  assign n25 = n21 & n22;
  assign n26 = ~n20 & ~n630;
  assign n27 = n17 & ~n26;
  assign n28 = ~pi1 & ~pi3;
  assign n29 = n18 & ~n28;
  assign n30 = pi1 & ~pi3;
  assign n31 = ~n18 & ~n30;
  assign n32 = pi5 & ~n31;
  assign n33 = n18 & n28;
  assign n34 = ~n18 & n30;
  assign n35 = ~n33 & ~n34;
  assign n36 = pi5 & ~n35;
  assign n37 = ~n29 & n32;
  assign n38 = ~n27 & ~n631;
  assign n39 = pi9 & ~n38;
  assign n40 = ~pi6 & ~pi9;
  assign n41 = pi5 & pi7;
  assign n42 = ~pi6 & ~n41;
  assign n43 = ~pi9 & n42;
  assign n44 = n40 & ~n41;
  assign n45 = ~pi1 & n632;
  assign n46 = ~n39 & ~n45;
  assign n47 = ~pi4 & ~n46;
  assign n48 = ~pi5 & pi6;
  assign n49 = pi4 & ~pi9;
  assign n50 = pi7 & n49;
  assign n51 = pi7 & n48;
  assign n52 = n49 & n51;
  assign n53 = n48 & n50;
  assign n54 = pi4 & pi5;
  assign n55 = pi6 & n54;
  assign n56 = ~pi7 & n55;
  assign n57 = n17 & n54;
  assign n58 = ~pi4 & pi5;
  assign n59 = pi9 & n58;
  assign n60 = pi5 & pi9;
  assign n61 = ~n17 & n60;
  assign n62 = ~pi4 & n61;
  assign n63 = ~n17 & n59;
  assign n64 = ~n634 & ~n635;
  assign n65 = ~n633 & ~n635;
  assign n66 = ~n634 & n65;
  assign n67 = ~n633 & n64;
  assign n68 = ~pi3 & ~n636;
  assign n69 = ~pi4 & ~pi5;
  assign n70 = ~n54 & ~n69;
  assign n71 = ~pi6 & pi9;
  assign n72 = po3 & n71;
  assign n73 = ~pi6 & po3;
  assign n74 = pi9 & n69;
  assign n75 = pi4 & n60;
  assign n76 = ~n74 & ~n75;
  assign n77 = pi9 & ~n70;
  assign n78 = n73 & ~n637;
  assign n79 = ~n70 & n72;
  assign n80 = pi0 & pi6;
  assign n81 = ~pi4 & pi9;
  assign n82 = ~pi5 & n80;
  assign n83 = n81 & n82;
  assign n84 = n74 & n80;
  assign n85 = ~n638 & ~n639;
  assign n86 = pi7 & ~n85;
  assign n87 = ~pi7 & n48;
  assign n88 = ~pi5 & n17;
  assign n89 = po3 & ~n49;
  assign n90 = ~pi5 & po3;
  assign n91 = n17 & n90;
  assign n92 = ~n49 & n91;
  assign n93 = n640 & n89;
  assign n94 = pi6 & pi9;
  assign n95 = ~pi7 & ~pi9;
  assign n96 = ~pi6 & n95;
  assign n97 = ~pi7 & n40;
  assign n98 = ~n94 & ~n642;
  assign n99 = pi4 & ~pi5;
  assign n100 = ~n28 & n99;
  assign n101 = ~n98 & n100;
  assign n102 = ~n641 & ~n101;
  assign n103 = ~n86 & n102;
  assign n104 = ~n68 & n103;
  assign n105 = ~n68 & ~n101;
  assign n106 = ~n47 & n105;
  assign n107 = ~n86 & n106;
  assign n108 = ~n641 & n107;
  assign n109 = ~n47 & n104;
  assign n110 = pi6 & ~n643;
  assign n111 = pi4 & ~pi6;
  assign n112 = n21 & n111;
  assign n113 = pi1 & ~pi4;
  assign n114 = ~n30 & ~n113;
  assign n115 = ~n112 & n114;
  assign n116 = ~n30 & ~n110;
  assign n117 = ~n112 & ~n113;
  assign n118 = n116 & n117;
  assign n119 = ~n110 & n115;
  assign n120 = pi7 & ~n644;
  assign n121 = ~pi4 & pi6;
  assign n122 = ~pi7 & ~n643;
  assign n123 = n121 & ~n122;
  assign n124 = ~pi6 & ~n643;
  assign n125 = pi4 & ~pi7;
  assign n126 = pi3 & pi6;
  assign n127 = n125 & ~n126;
  assign n128 = ~pi3 & pi6;
  assign n129 = ~pi6 & n643;
  assign n130 = ~n128 & ~n129;
  assign n131 = pi4 & ~n130;
  assign n132 = ~pi7 & n131;
  assign n133 = ~n124 & n127;
  assign n134 = ~pi4 & ~pi6;
  assign n135 = ~pi4 & n124;
  assign n136 = ~n643 & n134;
  assign n137 = ~n645 & ~n646;
  assign n138 = ~n123 & ~n646;
  assign n139 = ~n645 & n138;
  assign n140 = ~n123 & n137;
  assign n141 = ~n120 & ~n646;
  assign n142 = ~n123 & n141;
  assign n143 = ~n645 & n142;
  assign n144 = ~n120 & n647;
  assign n145 = ~pi5 & ~n648;
  assign n146 = pi4 & pi6;
  assign n147 = pi1 & ~n643;
  assign n148 = pi4 & n147;
  assign n149 = pi6 & n148;
  assign n150 = n146 & n147;
  assign n151 = po3 & n121;
  assign n152 = ~pi4 & n17;
  assign n153 = n17 & n28;
  assign n154 = ~pi4 & n153;
  assign n155 = n28 & n152;
  assign n156 = ~n151 & ~n650;
  assign n157 = ~n649 & n156;
  assign n158 = pi5 & ~n157;
  assign n159 = ~pi4 & pi7;
  assign n160 = pi5 & n159;
  assign n161 = pi7 & n58;
  assign n162 = ~n646 & ~n651;
  assign n163 = pi3 & ~n162;
  assign n164 = pi3 & pi5;
  assign n165 = ~pi6 & ~n164;
  assign n166 = pi1 & pi7;
  assign n167 = pi1 & pi6;
  assign n168 = pi5 & po3;
  assign n169 = ~n167 & ~n168;
  assign n170 = pi7 & ~n169;
  assign n171 = ~n165 & n166;
  assign n172 = ~n163 & ~n652;
  assign n173 = ~n158 & ~n163;
  assign n174 = ~n652 & n173;
  assign n175 = ~n158 & n172;
  assign n176 = ~n145 & n653;
  assign n177 = ~pi9 & ~n176;
  assign n178 = ~pi6 & n54;
  assign n179 = ~pi7 & n178;
  assign n180 = ~pi2 & ~n636;
  assign n181 = ~pi6 & pi7;
  assign n182 = pi9 & n181;
  assign n183 = pi7 & n71;
  assign n184 = ~n152 & ~n654;
  assign n185 = pi0 & pi2;
  assign n186 = ~n70 & n185;
  assign n187 = pi7 & ~n70;
  assign n188 = ~pi6 & n187;
  assign n189 = pi9 & n188;
  assign n190 = ~pi4 & n640;
  assign n191 = ~n189 & ~n190;
  assign n192 = n185 & ~n191;
  assign n193 = ~n184 & n186;
  assign n194 = ~pi0 & ~pi2;
  assign n195 = n99 & ~n194;
  assign n196 = ~n98 & n99;
  assign n197 = ~n194 & n196;
  assign n198 = ~n98 & n195;
  assign n199 = ~n655 & ~n656;
  assign n200 = ~n180 & n199;
  assign n201 = ~pi0 & n632;
  assign n202 = ~pi0 & ~n17;
  assign n203 = pi0 & ~pi2;
  assign n204 = ~n18 & ~n203;
  assign n205 = ~n185 & ~n194;
  assign n206 = n60 & ~n657;
  assign n207 = n17 & n18;
  assign n208 = ~n203 & ~n207;
  assign n209 = n60 & ~n208;
  assign n210 = ~n202 & n206;
  assign n211 = ~n201 & ~n658;
  assign n212 = ~pi4 & ~n211;
  assign n213 = ~n180 & ~n656;
  assign n214 = ~n212 & n213;
  assign n215 = ~n655 & n214;
  assign n216 = n200 & ~n212;
  assign n217 = n54 & n659;
  assign n218 = n54 & n200;
  assign n219 = ~pi6 & n660;
  assign n220 = ~pi6 & ~n69;
  assign n221 = ~pi0 & ~n220;
  assign n222 = ~n659 & n221;
  assign n223 = ~n219 & ~n222;
  assign n224 = pi7 & ~n223;
  assign n225 = ~pi0 & n659;
  assign n226 = pi9 & n651;
  assign n227 = n60 & n159;
  assign n228 = ~n225 & n661;
  assign n229 = pi9 & n17;
  assign n230 = pi0 & ~n659;
  assign n231 = n54 & n230;
  assign n232 = n99 & n185;
  assign n233 = n69 & n659;
  assign n234 = ~n232 & ~n233;
  assign n235 = ~n231 & n234;
  assign n236 = n229 & ~n235;
  assign n237 = ~n228 & ~n236;
  assign n238 = pi4 & n640;
  assign n239 = n48 & n125;
  assign n240 = pi9 & n662;
  assign n241 = n99 & n229;
  assign n242 = n237 & n663;
  assign n243 = pi0 & ~pi4;
  assign n244 = ~pi5 & ~pi6;
  assign n245 = ~pi6 & n243;
  assign n246 = ~pi5 & n245;
  assign n247 = n243 & n244;
  assign n248 = ~n242 & ~n664;
  assign n249 = n659 & ~n248;
  assign n250 = ~pi7 & n237;
  assign n251 = ~pi7 & ~n236;
  assign n252 = n237 & n243;
  assign n253 = ~pi7 & n252;
  assign n254 = n243 & n665;
  assign n255 = pi4 & ~n657;
  assign n256 = ~pi6 & n255;
  assign n257 = n111 & ~n657;
  assign n258 = ~n666 & ~n667;
  assign n259 = ~pi5 & ~n258;
  assign n260 = ~pi0 & pi7;
  assign n261 = ~n665 & ~n260;
  assign n262 = n55 & ~n261;
  assign n263 = pi6 & ~n659;
  assign n264 = pi0 & ~n54;
  assign n265 = ~n17 & ~n181;
  assign n266 = pi0 & ~n17;
  assign n267 = ~n54 & ~n181;
  assign n268 = n266 & n267;
  assign n269 = n264 & n265;
  assign n270 = n80 & n659;
  assign n271 = pi7 & n270;
  assign n272 = pi0 & ~pi7;
  assign n273 = ~pi6 & n272;
  assign n274 = ~n271 & ~n273;
  assign n275 = ~n54 & ~n274;
  assign n276 = ~n263 & n668;
  assign n277 = ~n262 & ~n669;
  assign n278 = ~n259 & n277;
  assign n279 = ~n249 & n278;
  assign n280 = ~pi6 & n659;
  assign n281 = ~pi6 & ~n659;
  assign n282 = pi6 & n659;
  assign n283 = ~n281 & ~n282;
  assign n284 = ~n263 & ~n280;
  assign n285 = n58 & ~n670;
  assign n286 = n181 & n185;
  assign n287 = ~pi6 & n185;
  assign n288 = n661 & n287;
  assign n289 = n59 & n286;
  assign n290 = ~n242 & ~n671;
  assign n291 = n99 & n263;
  assign n292 = n48 & ~n659;
  assign n293 = pi4 & n290;
  assign n294 = n292 & n293;
  assign n295 = n290 & n291;
  assign n296 = ~n285 & ~n672;
  assign n297 = ~pi7 & ~n296;
  assign n298 = ~pi6 & n651;
  assign n299 = n58 & n181;
  assign n300 = n58 & n290;
  assign n301 = n181 & n300;
  assign n302 = n290 & n673;
  assign n303 = ~pi0 & ~pi4;
  assign n304 = ~pi0 & ~pi7;
  assign n305 = ~pi4 & n48;
  assign n306 = n304 & n305;
  assign n307 = n640 & n303;
  assign n308 = ~n674 & ~n675;
  assign n309 = ~n237 & ~n308;
  assign n310 = ~n297 & ~n309;
  assign n311 = n278 & ~n309;
  assign n312 = ~n249 & ~n297;
  assign n313 = n311 & n312;
  assign n314 = n279 & n310;
  assign n315 = ~n259 & ~n297;
  assign n316 = ~n249 & n315;
  assign n317 = ~n224 & n316;
  assign n318 = ~n309 & n317;
  assign n319 = ~n262 & n318;
  assign n320 = ~n669 & n319;
  assign n321 = ~n224 & n676;
  assign n322 = pi9 & ~n677;
  assign n323 = ~pi8 & n322;
  assign n324 = n643 & n659;
  assign n325 = n54 & n324;
  assign n326 = ~pi1 & n643;
  assign n327 = n661 & ~n326;
  assign n328 = n54 & n147;
  assign n329 = n69 & n643;
  assign n330 = po3 & n99;
  assign n331 = ~n329 & ~n330;
  assign n332 = ~n328 & n331;
  assign n333 = n229 & ~n332;
  assign n334 = ~n327 & ~n333;
  assign n335 = n663 & n334;
  assign n336 = n73 & n661;
  assign n337 = n72 & n651;
  assign n338 = ~n335 & ~n678;
  assign n339 = n671 & ~n338;
  assign n340 = ~n671 & n338;
  assign n341 = n671 & n338;
  assign n342 = ~n671 & ~n338;
  assign n343 = ~n341 & ~n342;
  assign n344 = ~n339 & ~n340;
  assign n345 = ~n334 & ~n679;
  assign n346 = n334 & n679;
  assign n347 = n58 & ~n346;
  assign n348 = ~n334 & n679;
  assign n349 = n334 & ~n679;
  assign n350 = ~n348 & ~n349;
  assign n351 = n58 & ~n350;
  assign n352 = ~n345 & n347;
  assign n353 = ~n325 & ~n680;
  assign n354 = ~pi6 & ~n353;
  assign n355 = ~n48 & ~n69;
  assign n356 = ~n48 & ~n121;
  assign n357 = ~n69 & n356;
  assign n358 = ~n121 & n355;
  assign n359 = ~n643 & n230;
  assign n360 = n643 & ~n230;
  assign n361 = ~n359 & ~n360;
  assign n362 = ~n681 & n361;
  assign n363 = ~pi0 & n54;
  assign n364 = pi6 & n363;
  assign n365 = ~pi0 & n55;
  assign n366 = ~n362 & ~n682;
  assign n367 = ~pi1 & ~n366;
  assign n368 = pi1 & n80;
  assign n369 = ~n643 & n281;
  assign n370 = ~n368 & ~n369;
  assign n371 = n54 & ~n370;
  assign n372 = ~n367 & ~n371;
  assign n373 = ~n354 & ~n371;
  assign n374 = ~n367 & n373;
  assign n375 = ~n354 & n372;
  assign n376 = pi7 & ~n683;
  assign n377 = ~n659 & ~n290;
  assign n378 = n643 & ~n377;
  assign n379 = ~n643 & n377;
  assign n380 = ~n378 & ~n379;
  assign n381 = ~n338 & n380;
  assign n382 = n338 & ~n380;
  assign n383 = n99 & ~n382;
  assign n384 = n338 & ~n377;
  assign n385 = n338 & ~n379;
  assign n386 = ~n338 & n377;
  assign n387 = n338 & n377;
  assign n388 = ~n338 & ~n377;
  assign n389 = ~n387 & ~n388;
  assign n390 = ~n684 & ~n386;
  assign n391 = ~n643 & n685;
  assign n392 = n643 & ~n685;
  assign n393 = ~n391 & ~n392;
  assign n394 = n99 & ~n393;
  assign n395 = ~n381 & n383;
  assign n396 = pi0 & ~n237;
  assign n397 = n334 & ~n396;
  assign n398 = ~n334 & n396;
  assign n399 = ~n334 & ~n396;
  assign n400 = n334 & n396;
  assign n401 = ~n399 & ~n400;
  assign n402 = ~n397 & ~n398;
  assign n403 = ~pi1 & n69;
  assign n404 = ~n687 & n403;
  assign n405 = n54 & n237;
  assign n406 = n237 & n334;
  assign n407 = n54 & n406;
  assign n408 = n334 & n405;
  assign n409 = n54 & ~n237;
  assign n410 = ~n237 & ~n334;
  assign n411 = n54 & n410;
  assign n412 = ~n334 & n409;
  assign n413 = ~n688 & ~n689;
  assign n414 = ~n404 & n413;
  assign n415 = ~n686 & n414;
  assign n416 = pi6 & ~n415;
  assign n417 = pi1 & n69;
  assign n418 = ~pi5 & n687;
  assign n419 = n113 & n418;
  assign n420 = n687 & n417;
  assign n421 = pi6 & n324;
  assign n422 = ~n643 & ~n659;
  assign n423 = ~n421 & ~n422;
  assign n424 = n58 & ~n423;
  assign n425 = ~pi6 & ~n54;
  assign n426 = pi5 & ~n643;
  assign n427 = ~pi1 & ~n426;
  assign n428 = n58 & ~n643;
  assign n429 = pi1 & ~n54;
  assign n430 = ~n428 & ~n429;
  assign n431 = ~pi6 & ~n430;
  assign n432 = n425 & ~n427;
  assign n433 = ~n424 & ~n691;
  assign n434 = n69 & n687;
  assign n435 = ~n425 & ~n434;
  assign n436 = pi1 & ~n435;
  assign n437 = ~n124 & ~n422;
  assign n438 = ~n421 & n437;
  assign n439 = n58 & ~n438;
  assign n440 = ~n436 & ~n439;
  assign n441 = ~n690 & n433;
  assign n442 = ~n416 & ~n690;
  assign n443 = ~n424 & n442;
  assign n444 = ~n691 & n443;
  assign n445 = ~n416 & n692;
  assign n446 = ~pi7 & ~n693;
  assign n447 = n113 & n244;
  assign n448 = pi1 & ~n681;
  assign n449 = pi7 & n448;
  assign n450 = n166 & ~n681;
  assign n451 = ~n447 & ~n694;
  assign n452 = ~n361 & ~n451;
  assign n453 = ~pi5 & n111;
  assign n454 = pi4 & n244;
  assign n455 = pi7 & n28;
  assign n456 = ~po3 & ~n455;
  assign n457 = n185 & ~n456;
  assign n458 = ~n21 & ~n30;
  assign n459 = ~po3 & ~n28;
  assign n460 = ~n185 & ~po2;
  assign n461 = pi3 & ~pi7;
  assign n462 = ~n460 & ~n461;
  assign n463 = ~n457 & n462;
  assign n464 = n185 & n695;
  assign n465 = ~pi6 & n232;
  assign n466 = ~n456 & n697;
  assign n467 = n695 & ~n462;
  assign n468 = ~n466 & ~n467;
  assign n469 = n695 & ~n463;
  assign n470 = ~n452 & n698;
  assign n471 = ~n446 & n470;
  assign n472 = ~n376 & ~n446;
  assign n473 = ~n467 & n472;
  assign n474 = ~n452 & n473;
  assign n475 = ~n466 & n474;
  assign n476 = ~n376 & n471;
  assign n477 = pi9 & ~n699;
  assign n478 = n323 & n477;
  assign n479 = n323 & ~n699;
  assign n480 = ~n323 & n699;
  assign n481 = ~n700 & ~n480;
  assign n482 = ~n179 & ~n481;
  assign n483 = ~n323 & n477;
  assign n484 = n323 & ~n477;
  assign n485 = ~n179 & ~n484;
  assign n486 = ~n483 & n485;
  assign n487 = pi9 & ~n486;
  assign n488 = pi9 & ~n482;
  assign n489 = ~n177 & ~n701;
  assign n490 = pi5 & n121;
  assign n491 = ~pi7 & n490;
  assign n492 = n17 & n58;
  assign n493 = ~n178 & ~n702;
  assign n494 = n324 & ~n493;
  assign n495 = ~pi6 & n58;
  assign n496 = ~n340 & n495;
  assign n497 = ~n334 & n496;
  assign n498 = ~n334 & ~n340;
  assign n499 = ~n147 & ~n230;
  assign n500 = ~n326 & ~n681;
  assign n501 = n230 & ~n326;
  assign n502 = ~n147 & ~n501;
  assign n503 = ~n681 & ~n502;
  assign n504 = ~n499 & n500;
  assign n505 = ~n28 & n185;
  assign n506 = ~po3 & ~n505;
  assign n507 = po3 & n695;
  assign n508 = ~pi6 & n330;
  assign n509 = ~n28 & n697;
  assign n510 = ~n705 & ~n509;
  assign n511 = n695 & ~n506;
  assign n512 = ~pi0 & ~pi1;
  assign n513 = ~pi1 & n682;
  assign n514 = n55 & n512;
  assign n515 = pi7 & ~n707;
  assign n516 = n706 & n515;
  assign n517 = ~n704 & n516;
  assign n518 = ~n703 & n517;
  assign n519 = ~n338 & ~n378;
  assign n520 = pi4 & ~n379;
  assign n521 = ~n519 & n520;
  assign n522 = pi1 & ~n397;
  assign n523 = ~pi4 & ~n398;
  assign n524 = ~n522 & n523;
  assign n525 = n48 & ~n524;
  assign n526 = pi4 & ~n378;
  assign n527 = ~n379 & ~n519;
  assign n528 = ~n684 & n526;
  assign n529 = ~pi1 & ~n398;
  assign n530 = ~pi4 & ~n397;
  assign n531 = ~n529 & n530;
  assign n532 = ~pi1 & ~n396;
  assign n533 = ~pi4 & ~n532;
  assign n534 = ~n334 & n533;
  assign n535 = n113 & n396;
  assign n536 = n708 & ~n535;
  assign n537 = ~n534 & n536;
  assign n538 = n708 & ~n531;
  assign n539 = n48 & ~n709;
  assign n540 = ~n521 & n525;
  assign n541 = ~pi7 & ~n178;
  assign n542 = ~n688 & n541;
  assign n543 = ~n710 & n542;
  assign n544 = ~n518 & ~n543;
  assign n545 = ~n688 & ~n710;
  assign n546 = ~pi7 & ~n545;
  assign n547 = ~n705 & ~n707;
  assign n548 = ~n509 & n547;
  assign n549 = n706 & ~n707;
  assign n550 = ~n704 & n711;
  assign n551 = ~n703 & n550;
  assign n552 = pi7 & ~n551;
  assign n553 = ~n494 & ~n552;
  assign n554 = ~n546 & n553;
  assign n555 = ~n494 & ~n544;
  assign n556 = ~n700 & ~n552;
  assign n557 = ~n546 & n556;
  assign n558 = ~n494 & n557;
  assign n559 = ~n700 & n712;
  assign po4 = pi9 & ~n713;
  assign n561 = pi8 & ~n322;
  assign n562 = ~n323 & ~n561;
  assign n563 = pi8 & n322;
  assign n564 = ~pi8 & ~n322;
  assign n565 = ~n179 & ~n564;
  assign n566 = ~n563 & n565;
  assign n567 = ~n179 & ~n562;
  assign n568 = pi9 & ~n714;
  assign n569 = ~pi0 & ~n111;
  assign n570 = pi2 & ~n111;
  assign n571 = ~n657 & ~n570;
  assign n572 = ~n657 & ~n569;
  assign n573 = ~n121 & ~n243;
  assign n574 = ~n715 & n573;
  assign n575 = n18 & n111;
  assign n576 = ~n263 & ~n575;
  assign n577 = ~n203 & n573;
  assign n578 = n576 & n577;
  assign n579 = ~n263 & n574;
  assign n580 = ~pi5 & ~n716;
  assign n581 = pi5 & n185;
  assign n582 = ~n80 & ~n581;
  assign n583 = ~n580 & n582;
  assign n584 = pi7 & ~n583;
  assign n585 = ~pi4 & ~n670;
  assign n586 = pi2 & pi6;
  assign n587 = n125 & ~n586;
  assign n588 = ~pi2 & pi6;
  assign n589 = ~n280 & ~n588;
  assign n590 = pi4 & ~n589;
  assign n591 = ~pi7 & n590;
  assign n592 = ~n281 & n587;
  assign n593 = ~n585 & ~n717;
  assign n594 = ~pi5 & ~n593;
  assign n595 = pi6 & n230;
  assign n596 = pi4 & n595;
  assign n597 = n146 & n230;
  assign n598 = n121 & n185;
  assign n599 = n17 & n194;
  assign n600 = ~pi4 & n599;
  assign n601 = n152 & n194;
  assign n602 = ~n598 & ~n719;
  assign n603 = ~n718 & ~n598;
  assign n604 = ~n719 & n603;
  assign n605 = ~n718 & n602;
  assign n606 = pi5 & ~n720;
  assign n607 = ~n41 & ~n281;
  assign n608 = pi2 & ~pi4;
  assign n609 = ~pi4 & n281;
  assign n610 = ~n651 & ~n609;
  assign n611 = pi2 & ~n610;
  assign n612 = ~n607 & n608;
  assign n613 = ~n606 & ~n721;
  assign n614 = ~n594 & n613;
  assign n615 = pi7 & ~n716;
  assign n616 = ~n717 & ~n615;
  assign n617 = ~n585 & ~n615;
  assign n618 = ~n717 & n617;
  assign n619 = ~n585 & n616;
  assign n620 = ~pi5 & ~n722;
  assign n621 = pi7 & ~n582;
  assign n622 = ~n721 & ~n621;
  assign n623 = n613 & ~n621;
  assign n624 = ~n606 & n622;
  assign n625 = ~n620 & n723;
  assign n626 = ~n584 & n614;
  assign n627 = ~pi9 & ~n724;
  assign n628 = ~n568 & ~n627;
  assign po5 = n657 & po2;
  assign n630 = n24 | n25;
  assign n631 = n36 | n37;
  assign n632 = n43 | n44;
  assign n633 = n52 | n53;
  assign n634 = n56 | n57;
  assign n635 = n62 | n63;
  assign n636 = n66 | n67;
  assign n637 = n76 | ~n77;
  assign n638 = n78 | n79;
  assign n639 = n83 | n84;
  assign n640 = n87 | n88;
  assign n641 = n92 | n93;
  assign n642 = n96 | n97;
  assign n643 = n108 | n109;
  assign n644 = n118 | n119;
  assign n645 = n132 | n133;
  assign n646 = n135 | n136;
  assign n647 = n139 | n140;
  assign n648 = n143 | n144;
  assign n649 = n149 | n150;
  assign n650 = n154 | n155;
  assign n651 = n160 | n161;
  assign n652 = n170 | n171;
  assign n653 = n174 | n175;
  assign n654 = n182 | n183;
  assign n655 = n192 | n193;
  assign n656 = n197 | n198;
  assign n657 = n204 | ~n205;
  assign n658 = n209 | n210;
  assign n659 = n215 | n216;
  assign n660 = n217 | n218;
  assign n661 = n226 | n227;
  assign n662 = n238 | n239;
  assign n663 = n240 | n241;
  assign n664 = n246 | n247;
  assign n665 = n250 | n251;
  assign n666 = n253 | n254;
  assign n667 = n256 | n257;
  assign n668 = n268 | n269;
  assign n669 = n275 | n276;
  assign n670 = n283 | ~n284;
  assign n671 = n288 | n289;
  assign n672 = n294 | n295;
  assign n673 = n298 | n299;
  assign n674 = n301 | n302;
  assign n675 = n306 | n307;
  assign n676 = n313 | n314;
  assign n677 = n320 | n321;
  assign n678 = n336 | n337;
  assign n679 = n343 | ~n344;
  assign n680 = n351 | n352;
  assign n681 = n357 | n358;
  assign n682 = n364 | n365;
  assign n683 = n374 | n375;
  assign n684 = n384 | n385;
  assign n685 = n389 | ~n390;
  assign n686 = n394 | n395;
  assign n687 = n401 | ~n402;
  assign n688 = n407 | n408;
  assign n689 = n411 | n412;
  assign n690 = n419 | n420;
  assign n691 = n431 | n432;
  assign n692 = n440 | n441;
  assign n693 = n444 | n445;
  assign n694 = n449 | n450;
  assign n695 = n453 | n454;
  assign po2 = n458 | ~n459;
  assign n697 = n464 | n465;
  assign n698 = n468 | ~n469;
  assign n699 = n475 | n476;
  assign n700 = n478 | n479;
  assign n701 = n487 | n488;
  assign n702 = n491 | n492;
  assign n703 = n497 | n498;
  assign n704 = n503 | n504;
  assign n705 = n507 | n508;
  assign n706 = n510 | ~n511;
  assign n707 = n513 | n514;
  assign n708 = n527 | ~n528;
  assign n709 = n537 | n538;
  assign n710 = n539 | n540;
  assign n711 = n548 | n549;
  assign n712 = n554 | n555;
  assign n713 = n558 | n559;
  assign n714 = n566 | n567;
  assign n715 = n571 | n572;
  assign n716 = n578 | n579;
  assign n717 = n591 | n592;
  assign n718 = n596 | n597;
  assign n719 = n600 | n601;
  assign n720 = n604 | n605;
  assign n721 = n611 | n612;
  assign n722 = n618 | n619;
  assign n723 = n623 | n624;
  assign n724 = n625 | n626;
  assign po0 = ~n628;
  assign po1 = ~n489;
endmodule
