module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7;
  wire n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902,
    n903, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n924, n925,
    n926, n927, n928, n931, n932, n933, n934,
    n935, n936;
  assign n137 = ~pi123  & pi125 ;
  assign n138 = ~pi126  & n137;
  assign n139 = pi124  & ~pi125 ;
  assign n140 = ~pi126  & ~n139;
  assign n141 = pi123  & n140;
  assign n142 = ~pi127  & ~n138;
  assign n143 = ~n141 & n142;
  assign n144 = ~pi121  & ~n143;
  assign n145 = ~pi127  & ~n140;
  assign n146 = ~pi122  & ~n145;
  assign n147 = pi122  & ~n143;
  assign n148 = ~n146 & ~n147;
  assign n149 = pi121  & ~n148;
  assign n150 = ~n144 & ~n149;
  assign n151 = ~pi119  & ~n150;
  assign n152 = ~pi120  & ~n148;
  assign n153 = pi120  & ~n150;
  assign n154 = ~n152 & ~n153;
  assign n155 = pi119  & ~n154;
  assign n156 = ~n151 & ~n155;
  assign n157 = ~pi117  & ~n156;
  assign n158 = ~pi118  & ~n154;
  assign n159 = pi118  & ~n156;
  assign n160 = ~n158 & ~n159;
  assign n161 = pi117  & ~n160;
  assign n162 = ~n157 & ~n161;
  assign n163 = ~pi115  & ~n162;
  assign n164 = ~pi116  & ~n160;
  assign n165 = pi116  & ~n162;
  assign n166 = ~n164 & ~n165;
  assign n167 = pi115  & ~n166;
  assign n168 = ~n163 & ~n167;
  assign n169 = ~pi113  & ~n168;
  assign n170 = ~pi114  & ~n166;
  assign n171 = pi114  & ~n168;
  assign n172 = ~n170 & ~n171;
  assign n173 = pi113  & ~n172;
  assign n174 = ~n169 & ~n173;
  assign n175 = ~pi111  & ~n174;
  assign n176 = ~pi112  & ~n172;
  assign n177 = pi112  & ~n174;
  assign n178 = ~n176 & ~n177;
  assign n179 = pi111  & ~n178;
  assign n180 = ~n175 & ~n179;
  assign n181 = ~pi109  & ~n180;
  assign n182 = ~pi110  & ~n178;
  assign n183 = pi110  & ~n180;
  assign n184 = ~n182 & ~n183;
  assign n185 = pi109  & ~n184;
  assign n186 = ~n181 & ~n185;
  assign n187 = ~pi107  & ~n186;
  assign n188 = ~pi108  & ~n184;
  assign n189 = pi108  & ~n186;
  assign n190 = ~n188 & ~n189;
  assign n191 = pi107  & ~n190;
  assign n192 = ~n187 & ~n191;
  assign n193 = ~pi105  & ~n192;
  assign n194 = ~pi106  & ~n190;
  assign n195 = pi106  & ~n192;
  assign n196 = ~n194 & ~n195;
  assign n197 = pi105  & ~n196;
  assign n198 = ~n193 & ~n197;
  assign n199 = ~pi103  & ~n198;
  assign n200 = ~pi104  & ~n196;
  assign n201 = pi104  & ~n198;
  assign n202 = ~n200 & ~n201;
  assign n203 = pi103  & ~n202;
  assign n204 = ~n199 & ~n203;
  assign n205 = ~pi101  & ~n204;
  assign n206 = ~pi102  & ~n202;
  assign n207 = pi102  & ~n204;
  assign n208 = ~n206 & ~n207;
  assign n209 = pi101  & ~n208;
  assign n210 = ~n205 & ~n209;
  assign n211 = ~pi99  & ~n210;
  assign n212 = ~pi100  & ~n208;
  assign n213 = pi100  & ~n210;
  assign n214 = ~n212 & ~n213;
  assign n215 = pi99  & ~n214;
  assign n216 = ~n211 & ~n215;
  assign n217 = ~pi97  & ~n216;
  assign n218 = ~pi98  & ~n214;
  assign n219 = pi98  & ~n216;
  assign n220 = ~n218 & ~n219;
  assign n221 = pi97  & ~n220;
  assign n222 = ~n217 & ~n221;
  assign n223 = ~pi95  & ~n222;
  assign n224 = ~pi96  & ~n220;
  assign n225 = pi96  & ~n222;
  assign n226 = ~n224 & ~n225;
  assign n227 = pi95  & ~n226;
  assign n228 = ~n223 & ~n227;
  assign n229 = ~pi93  & ~n228;
  assign n230 = ~pi94  & ~n226;
  assign n231 = pi94  & ~n228;
  assign n232 = ~n230 & ~n231;
  assign n233 = pi93  & ~n232;
  assign n234 = ~n229 & ~n233;
  assign n235 = ~pi91  & ~n234;
  assign n236 = ~pi92  & ~n232;
  assign n237 = pi92  & ~n234;
  assign n238 = ~n236 & ~n237;
  assign n239 = pi91  & ~n238;
  assign n240 = ~n235 & ~n239;
  assign n241 = ~pi89  & ~n240;
  assign n242 = ~pi90  & ~n238;
  assign n243 = pi90  & ~n240;
  assign n244 = ~n242 & ~n243;
  assign n245 = pi89  & ~n244;
  assign n246 = ~n241 & ~n245;
  assign n247 = ~pi87  & ~n246;
  assign n248 = ~pi88  & ~n244;
  assign n249 = pi88  & ~n246;
  assign n250 = ~n248 & ~n249;
  assign n251 = pi87  & ~n250;
  assign n252 = ~n247 & ~n251;
  assign n253 = ~pi85  & ~n252;
  assign n254 = ~pi86  & ~n250;
  assign n255 = pi86  & ~n252;
  assign n256 = ~n254 & ~n255;
  assign n257 = pi85  & ~n256;
  assign n258 = ~n253 & ~n257;
  assign n259 = ~pi83  & ~n258;
  assign n260 = ~pi84  & ~n256;
  assign n261 = pi84  & ~n258;
  assign n262 = ~n260 & ~n261;
  assign n263 = pi83  & ~n262;
  assign n264 = ~n259 & ~n263;
  assign n265 = ~pi81  & ~n264;
  assign n266 = ~pi82  & ~n262;
  assign n267 = pi82  & ~n264;
  assign n268 = ~n266 & ~n267;
  assign n269 = pi81  & ~n268;
  assign n270 = ~n265 & ~n269;
  assign n271 = ~pi79  & ~n270;
  assign n272 = ~pi80  & ~n268;
  assign n273 = pi80  & ~n270;
  assign n274 = ~n272 & ~n273;
  assign n275 = pi79  & ~n274;
  assign n276 = ~n271 & ~n275;
  assign n277 = ~pi77  & ~n276;
  assign n278 = ~pi78  & ~n274;
  assign n279 = pi78  & ~n276;
  assign n280 = ~n278 & ~n279;
  assign n281 = pi77  & ~n280;
  assign n282 = ~n277 & ~n281;
  assign n283 = ~pi75  & ~n282;
  assign n284 = ~pi76  & ~n280;
  assign n285 = pi76  & ~n282;
  assign n286 = ~n284 & ~n285;
  assign n287 = pi75  & ~n286;
  assign n288 = ~n283 & ~n287;
  assign n289 = ~pi73  & ~n288;
  assign n290 = ~pi74  & ~n286;
  assign n291 = pi74  & ~n288;
  assign n292 = ~n290 & ~n291;
  assign n293 = pi73  & ~n292;
  assign n294 = ~n289 & ~n293;
  assign n295 = ~pi71  & ~n294;
  assign n296 = ~pi72  & ~n292;
  assign n297 = pi72  & ~n294;
  assign n298 = ~n296 & ~n297;
  assign n299 = pi71  & ~n298;
  assign n300 = ~n295 & ~n299;
  assign n301 = ~pi69  & ~n300;
  assign n302 = ~pi70  & ~n298;
  assign n303 = pi70  & ~n300;
  assign n304 = ~n302 & ~n303;
  assign n305 = pi69  & ~n304;
  assign n306 = ~n301 & ~n305;
  assign n307 = ~pi67  & ~n306;
  assign n308 = ~pi68  & ~n304;
  assign n309 = pi68  & ~n306;
  assign n310 = ~n308 & ~n309;
  assign n311 = pi67  & ~n310;
  assign n312 = ~n307 & ~n311;
  assign n313 = ~pi65  & ~n312;
  assign n314 = ~pi66  & ~n310;
  assign n315 = pi66  & ~n312;
  assign n316 = ~n314 & ~n315;
  assign n317 = pi65  & ~n316;
  assign n318 = ~n313 & ~n317;
  assign n319 = ~pi63  & ~n318;
  assign n320 = ~pi64  & ~n316;
  assign n321 = pi64  & ~n318;
  assign n322 = ~n320 & ~n321;
  assign n323 = pi63  & ~n322;
  assign n324 = ~n319 & ~n323;
  assign n325 = ~pi61  & ~n324;
  assign n326 = ~pi62  & ~n322;
  assign n327 = pi62  & ~n324;
  assign n328 = ~n326 & ~n327;
  assign n329 = pi61  & ~n328;
  assign n330 = ~n325 & ~n329;
  assign n331 = ~pi59  & ~n330;
  assign n332 = ~pi60  & ~n328;
  assign n333 = pi60  & ~n330;
  assign n334 = ~n332 & ~n333;
  assign n335 = pi59  & ~n334;
  assign n336 = ~n331 & ~n335;
  assign n337 = ~pi57  & ~n336;
  assign n338 = ~pi58  & ~n334;
  assign n339 = pi58  & ~n336;
  assign n340 = ~n338 & ~n339;
  assign n341 = pi57  & ~n340;
  assign n342 = ~n337 & ~n341;
  assign n343 = ~pi55  & ~n342;
  assign n344 = ~pi56  & ~n340;
  assign n345 = pi56  & ~n342;
  assign n346 = ~n344 & ~n345;
  assign n347 = pi55  & ~n346;
  assign n348 = ~n343 & ~n347;
  assign n349 = ~pi53  & ~n348;
  assign n350 = ~pi54  & ~n346;
  assign n351 = pi54  & ~n348;
  assign n352 = ~n350 & ~n351;
  assign n353 = pi53  & ~n352;
  assign n354 = ~n349 & ~n353;
  assign n355 = ~pi51  & ~n354;
  assign n356 = ~pi52  & ~n352;
  assign n357 = pi52  & ~n354;
  assign n358 = ~n356 & ~n357;
  assign n359 = pi51  & ~n358;
  assign n360 = ~n355 & ~n359;
  assign n361 = ~pi49  & ~n360;
  assign n362 = ~pi50  & ~n358;
  assign n363 = pi50  & ~n360;
  assign n364 = ~n362 & ~n363;
  assign n365 = pi49  & ~n364;
  assign n366 = ~n361 & ~n365;
  assign n367 = ~pi47  & ~n366;
  assign n368 = ~pi48  & ~n364;
  assign n369 = pi48  & ~n366;
  assign n370 = ~n368 & ~n369;
  assign n371 = pi47  & ~n370;
  assign n372 = ~n367 & ~n371;
  assign n373 = ~pi45  & ~n372;
  assign n374 = ~pi46  & ~n370;
  assign n375 = pi46  & ~n372;
  assign n376 = ~n374 & ~n375;
  assign n377 = pi45  & ~n376;
  assign n378 = ~n373 & ~n377;
  assign n379 = ~pi43  & ~n378;
  assign n380 = ~pi44  & ~n376;
  assign n381 = pi44  & ~n378;
  assign n382 = ~n380 & ~n381;
  assign n383 = pi43  & ~n382;
  assign n384 = ~n379 & ~n383;
  assign n385 = ~pi41  & ~n384;
  assign n386 = ~pi42  & ~n382;
  assign n387 = pi42  & ~n384;
  assign n388 = ~n386 & ~n387;
  assign n389 = pi41  & ~n388;
  assign n390 = ~n385 & ~n389;
  assign n391 = ~pi39  & ~n390;
  assign n392 = ~pi40  & ~n388;
  assign n393 = pi40  & ~n390;
  assign n394 = ~n392 & ~n393;
  assign n395 = pi39  & ~n394;
  assign n396 = ~n391 & ~n395;
  assign n397 = ~pi37  & ~n396;
  assign n398 = ~pi38  & ~n394;
  assign n399 = pi38  & ~n396;
  assign n400 = ~n398 & ~n399;
  assign n401 = pi37  & ~n400;
  assign n402 = ~n397 & ~n401;
  assign n403 = ~pi35  & ~n402;
  assign n404 = ~pi36  & ~n400;
  assign n405 = pi36  & ~n402;
  assign n406 = ~n404 & ~n405;
  assign n407 = pi35  & ~n406;
  assign n408 = ~n403 & ~n407;
  assign n409 = ~pi33  & ~n408;
  assign n410 = ~pi34  & ~n406;
  assign n411 = pi34  & ~n408;
  assign n412 = ~n410 & ~n411;
  assign n413 = pi33  & ~n412;
  assign n414 = ~n409 & ~n413;
  assign n415 = ~pi31  & ~n414;
  assign n416 = ~pi32  & ~n412;
  assign n417 = pi32  & ~n414;
  assign n418 = ~n416 & ~n417;
  assign n419 = pi31  & ~n418;
  assign n420 = ~n415 & ~n419;
  assign n421 = ~pi29  & ~n420;
  assign n422 = ~pi30  & ~n418;
  assign n423 = pi30  & ~n420;
  assign n424 = ~n422 & ~n423;
  assign n425 = pi29  & ~n424;
  assign n426 = ~n421 & ~n425;
  assign n427 = ~pi27  & ~n426;
  assign n428 = ~pi28  & ~n424;
  assign n429 = pi28  & ~n426;
  assign n430 = ~n428 & ~n429;
  assign n431 = pi27  & ~n430;
  assign n432 = ~n427 & ~n431;
  assign n433 = ~pi25  & ~n432;
  assign n434 = ~pi26  & ~n430;
  assign n435 = pi26  & ~n432;
  assign n436 = ~n434 & ~n435;
  assign n437 = pi25  & ~n436;
  assign n438 = ~n433 & ~n437;
  assign n439 = ~pi23  & ~n438;
  assign n440 = ~pi24  & ~n436;
  assign n441 = pi24  & ~n438;
  assign n442 = ~n440 & ~n441;
  assign n443 = pi23  & ~n442;
  assign n444 = ~n439 & ~n443;
  assign n445 = ~pi21  & ~n444;
  assign n446 = ~pi22  & ~n442;
  assign n447 = pi22  & ~n444;
  assign n448 = ~n446 & ~n447;
  assign n449 = pi21  & ~n448;
  assign n450 = ~n445 & ~n449;
  assign n451 = ~pi19  & ~n450;
  assign n452 = ~pi20  & ~n448;
  assign n453 = pi20  & ~n450;
  assign n454 = ~n452 & ~n453;
  assign n455 = pi19  & ~n454;
  assign n456 = ~n451 & ~n455;
  assign n457 = ~pi17  & ~n456;
  assign n458 = ~pi18  & ~n454;
  assign n459 = pi18  & ~n456;
  assign n460 = ~n458 & ~n459;
  assign n461 = pi17  & ~n460;
  assign n462 = ~n457 & ~n461;
  assign n463 = ~pi15  & ~n462;
  assign n464 = ~pi16  & ~n460;
  assign n465 = pi16  & ~n462;
  assign n466 = ~n464 & ~n465;
  assign n467 = pi15  & ~n466;
  assign n468 = ~n463 & ~n467;
  assign n469 = ~pi13  & ~n468;
  assign n470 = ~pi14  & ~n466;
  assign n471 = pi14  & ~n468;
  assign n472 = ~n470 & ~n471;
  assign n473 = pi13  & ~n472;
  assign n474 = ~n469 & ~n473;
  assign n475 = ~pi11  & ~n474;
  assign n476 = ~pi12  & ~n472;
  assign n477 = pi12  & ~n474;
  assign n478 = ~n476 & ~n477;
  assign n479 = pi11  & ~n478;
  assign n480 = ~n475 & ~n479;
  assign n481 = ~pi9  & ~n480;
  assign n482 = ~pi10  & ~n478;
  assign n483 = pi10  & ~n480;
  assign n484 = ~n482 & ~n483;
  assign n485 = pi9  & ~n484;
  assign n486 = ~n481 & ~n485;
  assign n487 = ~pi7  & ~n486;
  assign n488 = ~pi8  & ~n484;
  assign n489 = pi8  & ~n486;
  assign n490 = ~n488 & ~n489;
  assign n491 = pi7  & ~n490;
  assign n492 = pi1  & ~pi2 ;
  assign n493 = ~pi3  & ~n492;
  assign n494 = ~pi4  & ~n493;
  assign n495 = ~pi5  & ~n494;
  assign n496 = ~pi6  & ~n495;
  assign n497 = ~n487 & ~n496;
  assign n498 = ~n491 & n497;
  assign n499 = n490 & n496;
  assign po0  = ~n498 & ~n499;
  assign n501 = ~pi12  & ~pi13 ;
  assign n502 = ~pi14  & ~pi15 ;
  assign n503 = ~pi18  & ~pi19 ;
  assign n504 = ~pi22  & ~pi23 ;
  assign n505 = ~pi26  & ~pi27 ;
  assign n506 = ~pi30  & ~pi31 ;
  assign n507 = ~pi34  & ~pi35 ;
  assign n508 = ~pi38  & ~pi39 ;
  assign n509 = ~pi42  & ~pi43 ;
  assign n510 = ~pi46  & ~pi47 ;
  assign n511 = ~pi50  & ~pi51 ;
  assign n512 = ~pi54  & ~pi55 ;
  assign n513 = ~pi58  & ~pi59 ;
  assign n514 = ~pi62  & ~pi63 ;
  assign n515 = ~pi66  & ~pi67 ;
  assign n516 = ~pi70  & ~pi71 ;
  assign n517 = ~pi74  & ~pi75 ;
  assign n518 = ~pi78  & ~pi79 ;
  assign n519 = ~pi82  & ~pi83 ;
  assign n520 = ~pi86  & ~pi87 ;
  assign n521 = ~pi90  & ~pi91 ;
  assign n522 = ~pi94  & ~pi95 ;
  assign n523 = ~pi98  & ~pi99 ;
  assign n524 = ~pi102  & ~pi103 ;
  assign n525 = ~pi106  & ~pi107 ;
  assign n526 = ~pi110  & ~pi111 ;
  assign n527 = ~pi114  & ~pi115 ;
  assign n528 = ~pi116  & ~pi117 ;
  assign n529 = ~pi122  & ~pi123 ;
  assign n530 = pi121  & n529;
  assign n531 = ~pi124  & ~pi125 ;
  assign n532 = ~pi120  & n531;
  assign n533 = ~n530 & n532;
  assign n534 = ~pi126  & pi127 ;
  assign n535 = ~pi126  & ~n534;
  assign n536 = ~n529 & n531;
  assign n537 = pi120  & n536;
  assign n538 = ~n533 & n535;
  assign n539 = ~n537 & n538;
  assign n540 = n528 & ~n539;
  assign n541 = ~pi118  & ~pi119 ;
  assign n542 = n539 & ~n541;
  assign n543 = n535 & n541;
  assign n544 = ~n536 & n543;
  assign n545 = ~n542 & ~n544;
  assign n546 = ~n528 & n545;
  assign n547 = ~n540 & ~n546;
  assign n548 = ~n527 & ~n547;
  assign n549 = n527 & n545;
  assign n550 = ~n548 & ~n549;
  assign n551 = n526 & ~n550;
  assign n552 = ~pi112  & ~pi113 ;
  assign n553 = ~n550 & ~n552;
  assign n554 = ~n547 & n552;
  assign n555 = ~n553 & ~n554;
  assign n556 = ~n526 & ~n555;
  assign n557 = ~n551 & ~n556;
  assign n558 = n525 & ~n557;
  assign n559 = ~pi108  & ~pi109 ;
  assign n560 = ~n557 & ~n559;
  assign n561 = ~n555 & n559;
  assign n562 = ~n560 & ~n561;
  assign n563 = ~n525 & ~n562;
  assign n564 = ~n558 & ~n563;
  assign n565 = n524 & ~n564;
  assign n566 = ~pi104  & ~pi105 ;
  assign n567 = ~n564 & ~n566;
  assign n568 = ~n562 & n566;
  assign n569 = ~n567 & ~n568;
  assign n570 = ~n524 & ~n569;
  assign n571 = ~n565 & ~n570;
  assign n572 = n523 & ~n571;
  assign n573 = ~pi100  & ~pi101 ;
  assign n574 = ~n571 & ~n573;
  assign n575 = ~n569 & n573;
  assign n576 = ~n574 & ~n575;
  assign n577 = ~n523 & ~n576;
  assign n578 = ~n572 & ~n577;
  assign n579 = n522 & ~n578;
  assign n580 = ~pi96  & ~pi97 ;
  assign n581 = ~n578 & ~n580;
  assign n582 = ~n576 & n580;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~n522 & ~n583;
  assign n585 = ~n579 & ~n584;
  assign n586 = n521 & ~n585;
  assign n587 = ~pi92  & ~pi93 ;
  assign n588 = ~n585 & ~n587;
  assign n589 = ~n583 & n587;
  assign n590 = ~n588 & ~n589;
  assign n591 = ~n521 & ~n590;
  assign n592 = ~n586 & ~n591;
  assign n593 = n520 & ~n592;
  assign n594 = ~pi88  & ~pi89 ;
  assign n595 = ~n592 & ~n594;
  assign n596 = ~n590 & n594;
  assign n597 = ~n595 & ~n596;
  assign n598 = ~n520 & ~n597;
  assign n599 = ~n593 & ~n598;
  assign n600 = n519 & ~n599;
  assign n601 = ~pi84  & ~pi85 ;
  assign n602 = ~n599 & ~n601;
  assign n603 = ~n597 & n601;
  assign n604 = ~n602 & ~n603;
  assign n605 = ~n519 & ~n604;
  assign n606 = ~n600 & ~n605;
  assign n607 = n518 & ~n606;
  assign n608 = ~pi80  & ~pi81 ;
  assign n609 = ~n606 & ~n608;
  assign n610 = ~n604 & n608;
  assign n611 = ~n609 & ~n610;
  assign n612 = ~n518 & ~n611;
  assign n613 = ~n607 & ~n612;
  assign n614 = n517 & ~n613;
  assign n615 = ~pi76  & ~pi77 ;
  assign n616 = ~n613 & ~n615;
  assign n617 = ~n611 & n615;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~n517 & ~n618;
  assign n620 = ~n614 & ~n619;
  assign n621 = n516 & ~n620;
  assign n622 = ~pi72  & ~pi73 ;
  assign n623 = ~n620 & ~n622;
  assign n624 = ~n618 & n622;
  assign n625 = ~n623 & ~n624;
  assign n626 = ~n516 & ~n625;
  assign n627 = ~n621 & ~n626;
  assign n628 = n515 & ~n627;
  assign n629 = ~pi68  & ~pi69 ;
  assign n630 = ~n627 & ~n629;
  assign n631 = ~n625 & n629;
  assign n632 = ~n630 & ~n631;
  assign n633 = ~n515 & ~n632;
  assign n634 = ~n628 & ~n633;
  assign n635 = n514 & ~n634;
  assign n636 = ~pi64  & ~pi65 ;
  assign n637 = ~n634 & ~n636;
  assign n638 = ~n632 & n636;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~n514 & ~n639;
  assign n641 = ~n635 & ~n640;
  assign n642 = n513 & ~n641;
  assign n643 = ~pi60  & ~pi61 ;
  assign n644 = ~n641 & ~n643;
  assign n645 = ~n639 & n643;
  assign n646 = ~n644 & ~n645;
  assign n647 = ~n513 & ~n646;
  assign n648 = ~n642 & ~n647;
  assign n649 = n512 & ~n648;
  assign n650 = ~pi56  & ~pi57 ;
  assign n651 = ~n648 & ~n650;
  assign n652 = ~n646 & n650;
  assign n653 = ~n651 & ~n652;
  assign n654 = ~n512 & ~n653;
  assign n655 = ~n649 & ~n654;
  assign n656 = n511 & ~n655;
  assign n657 = ~pi52  & ~pi53 ;
  assign n658 = ~n655 & ~n657;
  assign n659 = ~n653 & n657;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n511 & ~n660;
  assign n662 = ~n656 & ~n661;
  assign n663 = n510 & ~n662;
  assign n664 = ~pi48  & ~pi49 ;
  assign n665 = ~n662 & ~n664;
  assign n666 = ~n660 & n664;
  assign n667 = ~n665 & ~n666;
  assign n668 = ~n510 & ~n667;
  assign n669 = ~n663 & ~n668;
  assign n670 = n509 & ~n669;
  assign n671 = ~pi44  & ~pi45 ;
  assign n672 = ~n669 & ~n671;
  assign n673 = ~n667 & n671;
  assign n674 = ~n672 & ~n673;
  assign n675 = ~n509 & ~n674;
  assign n676 = ~n670 & ~n675;
  assign n677 = n508 & ~n676;
  assign n678 = ~pi40  & ~pi41 ;
  assign n679 = ~n676 & ~n678;
  assign n680 = ~n674 & n678;
  assign n681 = ~n679 & ~n680;
  assign n682 = ~n508 & ~n681;
  assign n683 = ~n677 & ~n682;
  assign n684 = n507 & ~n683;
  assign n685 = ~pi36  & ~pi37 ;
  assign n686 = ~n683 & ~n685;
  assign n687 = ~n681 & n685;
  assign n688 = ~n686 & ~n687;
  assign n689 = ~n507 & ~n688;
  assign n690 = ~n684 & ~n689;
  assign n691 = n506 & ~n690;
  assign n692 = ~pi32  & ~pi33 ;
  assign n693 = ~n690 & ~n692;
  assign n694 = ~n688 & n692;
  assign n695 = ~n693 & ~n694;
  assign n696 = ~n506 & ~n695;
  assign n697 = ~n691 & ~n696;
  assign n698 = n505 & ~n697;
  assign n699 = ~pi28  & ~pi29 ;
  assign n700 = ~n697 & ~n699;
  assign n701 = ~n695 & n699;
  assign n702 = ~n700 & ~n701;
  assign n703 = ~n505 & ~n702;
  assign n704 = ~n698 & ~n703;
  assign n705 = n504 & ~n704;
  assign n706 = ~pi24  & ~pi25 ;
  assign n707 = ~n704 & ~n706;
  assign n708 = ~n702 & n706;
  assign n709 = ~n707 & ~n708;
  assign n710 = ~n504 & ~n709;
  assign n711 = ~n705 & ~n710;
  assign n712 = n503 & ~n711;
  assign n713 = ~pi20  & ~pi21 ;
  assign n714 = ~n711 & ~n713;
  assign n715 = ~n709 & n713;
  assign n716 = ~n714 & ~n715;
  assign n717 = ~n503 & ~n716;
  assign n718 = ~n712 & ~n717;
  assign n719 = n502 & ~n718;
  assign n720 = ~pi16  & ~pi17 ;
  assign n721 = ~n718 & ~n720;
  assign n722 = ~n716 & n720;
  assign n723 = ~n721 & ~n722;
  assign n724 = ~n502 & ~n723;
  assign n725 = ~n719 & ~n724;
  assign n726 = ~n501 & ~n725;
  assign n727 = n501 & ~n723;
  assign n728 = ~pi10  & ~pi11 ;
  assign n729 = ~pi8  & ~pi9 ;
  assign n730 = ~pi6  & ~pi7 ;
  assign n731 = ~pi4  & ~pi5 ;
  assign n732 = ~pi2  & ~pi3 ;
  assign n733 = n731 & ~n732;
  assign n734 = n730 & ~n733;
  assign n735 = n729 & ~n734;
  assign n736 = n728 & ~n735;
  assign n737 = ~n727 & ~n736;
  assign n738 = ~n726 & n737;
  assign n739 = n725 & n736;
  assign po1  = ~n738 & ~n739;
  assign n741 = n505 & n706;
  assign n742 = n507 & n692;
  assign n743 = n509 & n678;
  assign n744 = n511 & n664;
  assign n745 = n513 & n650;
  assign n746 = n515 & n636;
  assign n747 = n517 & n622;
  assign n748 = n519 & n608;
  assign n749 = n521 & n594;
  assign n750 = n523 & n580;
  assign n751 = n525 & n566;
  assign n752 = n531 & n535;
  assign n753 = n528 & n541;
  assign n754 = ~pi120  & ~pi121 ;
  assign n755 = n529 & n754;
  assign n756 = ~n753 & n755;
  assign n757 = n752 & ~n756;
  assign n758 = ~pi114  & n552;
  assign n759 = n757 & ~n758;
  assign n760 = pi115  & n753;
  assign n761 = n755 & ~n760;
  assign n762 = n752 & n758;
  assign n763 = ~n761 & n762;
  assign n764 = ~n759 & ~n763;
  assign n765 = n751 & ~n764;
  assign n766 = n526 & n559;
  assign n767 = ~n757 & n766;
  assign n768 = n764 & ~n766;
  assign n769 = ~n767 & ~n768;
  assign n770 = ~n751 & n769;
  assign n771 = ~n765 & ~n770;
  assign n772 = n750 & ~n771;
  assign n773 = n524 & n573;
  assign n774 = n771 & ~n773;
  assign n775 = ~n769 & n773;
  assign n776 = ~n774 & ~n775;
  assign n777 = ~n750 & n776;
  assign n778 = ~n772 & ~n777;
  assign n779 = n749 & ~n778;
  assign n780 = n522 & n587;
  assign n781 = ~n776 & n780;
  assign n782 = n778 & ~n780;
  assign n783 = ~n781 & ~n782;
  assign n784 = ~n749 & n783;
  assign n785 = ~n779 & ~n784;
  assign n786 = n748 & ~n785;
  assign n787 = n520 & n601;
  assign n788 = ~n783 & n787;
  assign n789 = n785 & ~n787;
  assign n790 = ~n788 & ~n789;
  assign n791 = ~n748 & n790;
  assign n792 = ~n786 & ~n791;
  assign n793 = n747 & ~n792;
  assign n794 = n518 & n615;
  assign n795 = n792 & ~n794;
  assign n796 = ~n790 & n794;
  assign n797 = ~n795 & ~n796;
  assign n798 = ~n747 & n797;
  assign n799 = ~n793 & ~n798;
  assign n800 = n746 & ~n799;
  assign n801 = n516 & n629;
  assign n802 = ~n797 & n801;
  assign n803 = n799 & ~n801;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~n746 & n804;
  assign n806 = ~n800 & ~n805;
  assign n807 = n745 & ~n806;
  assign n808 = n514 & n643;
  assign n809 = ~n804 & n808;
  assign n810 = n806 & ~n808;
  assign n811 = ~n809 & ~n810;
  assign n812 = ~n745 & n811;
  assign n813 = ~n807 & ~n812;
  assign n814 = n744 & ~n813;
  assign n815 = n512 & n657;
  assign n816 = ~n811 & n815;
  assign n817 = n813 & ~n815;
  assign n818 = ~n816 & ~n817;
  assign n819 = ~n744 & n818;
  assign n820 = ~n814 & ~n819;
  assign n821 = n743 & ~n820;
  assign n822 = n510 & n671;
  assign n823 = ~n818 & n822;
  assign n824 = n820 & ~n822;
  assign n825 = ~n823 & ~n824;
  assign n826 = ~n743 & n825;
  assign n827 = ~n821 & ~n826;
  assign n828 = n742 & ~n827;
  assign n829 = n508 & n685;
  assign n830 = ~n825 & n829;
  assign n831 = n827 & ~n829;
  assign n832 = ~n830 & ~n831;
  assign n833 = ~n742 & n832;
  assign n834 = ~n828 & ~n833;
  assign n835 = n741 & ~n834;
  assign n836 = n506 & n699;
  assign n837 = ~n832 & n836;
  assign n838 = n834 & ~n836;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~n741 & n839;
  assign n841 = n504 & n713;
  assign n842 = n503 & n720;
  assign n843 = n501 & n502;
  assign n844 = n728 & n729;
  assign n845 = n730 & n731;
  assign n846 = n844 & ~n845;
  assign n847 = n843 & ~n846;
  assign n848 = n842 & ~n847;
  assign n849 = n841 & ~n848;
  assign n850 = ~n835 & ~n849;
  assign n851 = ~n840 & n850;
  assign n852 = ~n839 & n849;
  assign po2  = n851 | n852;
  assign n854 = n744 & n815;
  assign n855 = n746 & n801;
  assign n856 = n748 & n787;
  assign n857 = n752 & n755;
  assign n858 = n751 & n766;
  assign n859 = ~pi115  & n753;
  assign n860 = n758 & n859;
  assign n861 = ~n858 & n860;
  assign n862 = n857 & ~n861;
  assign n863 = n573 & n750;
  assign n864 = ~pi102  & n863;
  assign n865 = n862 & ~n864;
  assign n866 = pi103  & n858;
  assign n867 = n860 & ~n866;
  assign n868 = n857 & n864;
  assign n869 = ~n867 & n868;
  assign n870 = ~n865 & ~n869;
  assign n871 = n856 & ~n870;
  assign n872 = n749 & n780;
  assign n873 = ~n862 & n872;
  assign n874 = n870 & ~n872;
  assign n875 = ~n873 & ~n874;
  assign n876 = ~n856 & n875;
  assign n877 = ~n871 & ~n876;
  assign n878 = n855 & ~n877;
  assign n879 = n615 & n747;
  assign n880 = n518 & n879;
  assign n881 = n877 & ~n880;
  assign n882 = ~n875 & n880;
  assign n883 = ~n881 & ~n882;
  assign n884 = ~n855 & n883;
  assign n885 = ~n878 & ~n884;
  assign n886 = n854 & ~n885;
  assign n887 = n745 & n808;
  assign n888 = ~n883 & n887;
  assign n889 = n885 & ~n887;
  assign n890 = ~n888 & ~n889;
  assign n891 = ~n854 & n890;
  assign n892 = n743 & n822;
  assign n893 = n742 & n829;
  assign n894 = n741 & n836;
  assign n895 = n841 & n842;
  assign n896 = n843 & n844;
  assign n897 = n895 & ~n896;
  assign n898 = n894 & ~n897;
  assign n899 = n893 & ~n898;
  assign n900 = n892 & ~n899;
  assign n901 = ~n886 & ~n900;
  assign n902 = ~n891 & n901;
  assign n903 = ~n890 & n900;
  assign po3  = n902 | n903;
  assign n905 = n857 & n860;
  assign n906 = n854 & n887;
  assign n907 = n892 & n893;
  assign n908 = n894 & n895;
  assign n909 = n907 & ~n908;
  assign n910 = n906 & ~n909;
  assign n911 = ~pi78  & n855;
  assign n912 = n879 & n911;
  assign n913 = ~n910 & n912;
  assign n914 = n856 & n872;
  assign n915 = pi79  & n914;
  assign n916 = n524 & n858;
  assign n917 = n863 & n916;
  assign n918 = ~n915 & n917;
  assign n919 = n913 & ~n918;
  assign n920 = ~n914 & n917;
  assign n921 = ~n913 & ~n920;
  assign n922 = ~n919 & ~n921;
  assign po4  = ~n905 | n922;
  assign n924 = n905 & n917;
  assign n925 = n906 & n907;
  assign n926 = ~pi79  & n914;
  assign n927 = n912 & n926;
  assign n928 = ~n925 & n927;
  assign po5  = ~n924 | n928;
  assign po6  = ~n924 | ~n927;
  assign n931 = ~pi0  & ~pi1 ;
  assign n932 = n732 & n931;
  assign n933 = n845 & n932;
  assign n934 = n896 & n933;
  assign n935 = n908 & n934;
  assign n936 = n925 & n935;
  assign po7 = po6  | ~n936;
endmodule
