module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24 ;
  wire n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n100, n101, n102, n103,
    n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061,
    n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331,
    n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231,
    n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3296, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321,
    n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561,
    n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591,
    n3592, n3593, n3594, n3595, n3596, n3597,
    n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621,
    n3622, n3623, n3624, n3625, n3627, n3628,
    n3629, n3630, n3631, n3632, n3633, n3634,
    n3635, n3636, n3637, n3638, n3639, n3640,
    n3641, n3642, n3643, n3644, n3645, n3646,
    n3647, n3648, n3649, n3650, n3651, n3652,
    n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664,
    n3665, n3666, n3667, n3668, n3669, n3670,
    n3671, n3672, n3673, n3674, n3675, n3676,
    n3677, n3678, n3679, n3680, n3681, n3682,
    n3683, n3684, n3685, n3686, n3687, n3688,
    n3689, n3690, n3691, n3692, n3693, n3694,
    n3695, n3696, n3697, n3698, n3699, n3700,
    n3701, n3702, n3703, n3704, n3705, n3706,
    n3707, n3708, n3709, n3710, n3711, n3712,
    n3713, n3714, n3715, n3716, n3717, n3718,
    n3719, n3720, n3721, n3722, n3723, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730,
    n3731, n3732, n3733, n3734, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742,
    n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3769, n3770, n3771, n3772, n3773,
    n3774, n3775, n3776, n3777, n3778, n3779,
    n3780, n3781, n3782, n3783, n3784, n3785,
    n3786, n3787, n3788, n3789, n3790, n3791,
    n3792, n3793, n3794, n3795, n3796, n3797,
    n3798, n3799, n3800, n3801, n3802, n3803,
    n3804, n3805, n3806, n3807, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815,
    n3816, n3817, n3818, n3819, n3820, n3821,
    n3822, n3823, n3824, n3825, n3826, n3827,
    n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3842, n3843, n3844, n3845,
    n3846, n3847, n3848, n3849, n3850, n3851,
    n3852, n3853, n3854, n3855, n3856, n3857,
    n3858, n3859, n3860, n3861, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881,
    n3882, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894,
    n3895, n3896, n3897, n3898, n3899, n3900,
    n3901, n3902, n3903, n3904, n3905, n3906,
    n3907, n3908, n3909, n3910, n3911, n3912,
    n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924,
    n3925, n3926, n3927, n3928, n3929, n3930,
    n3931, n3932, n3933, n3934, n3935, n3936,
    n3937, n3938, n3939, n3940, n3941, n3942,
    n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954,
    n3955, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966,
    n3967, n3968, n3969, n3970, n3971, n3972,
    n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990,
    n3991, n3993, n3994, n3995, n3996, n3997,
    n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027,
    n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057,
    n4058, n4059, n4060, n4061, n4062, n4063,
    n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4083, n4084, n4085, n4086, n4087,
    n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196,
    n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227,
    n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4249, n4250, n4251,
    n4252, n4253, n4254, n4255, n4256, n4257,
    n4258, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299,
    n4301, n4302, n4303, n4304, n4305, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312,
    n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324,
    n4325, n4326, n4327, n4328, n4329, n4330,
    n4331, n4332, n4333, n4334, n4335, n4336,
    n4337, n4338, n4339, n4340, n4341, n4342,
    n4343, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354,
    n4355, n4356, n4357, n4358, n4359, n4360,
    n4361, n4362, n4363, n4364, n4365, n4366,
    n4367, n4368, n4369, n4370, n4371, n4372,
    n4373, n4374, n4375, n4376, n4377, n4378,
    n4379, n4380, n4381, n4382, n4383, n4384,
    n4385, n4386, n4387, n4388, n4389, n4390,
    n4392, n4393, n4394, n4395, n4396, n4397,
    n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415,
    n4416, n4417, n4418, n4419, n4420, n4421,
    n4422, n4423, n4424, n4425, n4426, n4427,
    n4428, n4429, n4430, n4431, n4432, n4433,
    n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445,
    n4446, n4447, n4448, n4449, n4450, n4451,
    n4452, n4453, n4454, n4455, n4456, n4457,
    n4458, n4459, n4460, n4461, n4462, n4463,
    n4464, n4465, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682,
    n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707,
    n4708, n4709, n4710, n4711, n4712, n4713,
    n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737,
    n4738, n4739, n4740, n4741, n4742, n4743,
    n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761,
    n4763, n4764, n4765, n4766, n4767, n4768,
    n4769, n4770, n4771, n4772, n4773, n4774,
    n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786,
    n4787, n4788, n4789, n4790, n4791, n4792,
    n4793, n4794, n4795, n4796, n4797, n4798,
    n4799, n4800, n4801, n4802, n4803, n4804,
    n4805, n4806, n4807, n4808, n4809, n4810,
    n4811, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822,
    n4823, n4824, n4825, n4826, n4828, n4829,
    n4830, n4831, n4832, n4833, n4834, n4835,
    n4836, n4837, n4838, n4839, n4840, n4841,
    n4842, n4843, n4844, n4845, n4846, n4847,
    n4848, n4849, n4850, n4851, n4852, n4853,
    n4854, n4855, n4856, n4857, n4858, n4859,
    n4860, n4861, n4862, n4863, n4864, n4865,
    n4866, n4867, n4868, n4869, n4870, n4871,
    n4872, n4873, n4874, n4875, n4876, n4877,
    n4878, n4880, n4881, n4882, n4883, n4884,
    n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914,
    n4915, n4916, n4917, n4918, n4919, n4920,
    n4921, n4922, n4923, n4924, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4987, n4988, n4989,
    n4990, n4991, n4992, n4993, n4994, n4995,
    n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5003, n5004, n5005, n5007, n5008,
    n5009, n5010, n5011, n5012, n5013, n5014,
    n5015, n5016, n5017, n5018, n5019, n5020,
    n5021, n5022, n5023, n5024, n5025, n5026,
    n5027, n5028, n5029, n5031, n5032, n5033,
    n5034, n5035, n5036, n5037, n5038, n5039,
    n5040, n5041, n5042, n5043, n5044, n5045,
    n5046, n5048, n5049, n5050, n5051, n5052,
    n5053, n5054, n5055, n5056, n5057, n5058,
    n5059, n5060, n5061, n5062, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5083, n5084, n5085,
    n5086, n5087;
  assign n50 = ~pi0  & ~pi1 ;
  assign n51 = ~pi2  & n50;
  assign n52 = ~pi3  & n51;
  assign n53 = ~pi4  & n52;
  assign n54 = ~pi22  & ~n53;
  assign n55 = ~pi5  & ~n54;
  assign n56 = pi5  & n54;
  assign n57 = ~n55 & ~n56;
  assign n58 = pi18  & pi22 ;
  assign n59 = ~pi5  & n53;
  assign n60 = ~pi6  & n59;
  assign n61 = ~pi7  & n60;
  assign n62 = ~pi8  & n61;
  assign n63 = ~pi9  & n62;
  assign n64 = ~pi10  & n63;
  assign n65 = ~pi11  & n64;
  assign n66 = ~pi12  & n65;
  assign n67 = ~pi13  & n66;
  assign n68 = ~pi14  & n67;
  assign n69 = ~pi15  & n68;
  assign n70 = ~pi16  & n69;
  assign n71 = ~pi17  & n70;
  assign n72 = ~pi18  & n71;
  assign n73 = ~pi22  & ~n72;
  assign n74 = pi18  & ~n71;
  assign n75 = n73 & ~n74;
  assign n76 = ~n58 & ~n75;
  assign n77 = ~pi19  & ~n73;
  assign n78 = pi19  & n73;
  assign n79 = ~n77 & ~n78;
  assign n80 = ~n76 & n79;
  assign n81 = ~pi22  & ~n70;
  assign n82 = pi17  & ~n81;
  assign n83 = ~pi17  & n81;
  assign n84 = ~n82 & ~n83;
  assign n85 = ~pi22  & ~n69;
  assign n86 = pi16  & ~n85;
  assign n87 = ~pi16  & n85;
  assign n88 = ~n86 & ~n87;
  assign n89 = ~n84 & ~n88;
  assign n90 = n80 & n89;
  assign n91 = ~pi22  & ~n68;
  assign n92 = pi15  & ~n91;
  assign n93 = ~pi15  & n91;
  assign n94 = ~n92 & ~n93;
  assign n95 = pi20  & pi22 ;
  assign n96 = ~pi19  & n72;
  assign n97 = pi20  & ~n96;
  assign n98 = ~pi20  & n96;
  assign n99 = ~pi22  & ~n98;
  assign n100 = ~n97 & n99;
  assign n101 = ~n95 & ~n100;
  assign n102 = pi21  & ~n99;
  assign n103 = ~pi21  & ~pi22 ;
  assign n104 = ~n98 & n103;
  assign n105 = ~n102 & ~n104;
  assign n106 = ~n101 & n105;
  assign n107 = ~n94 & n106;
  assign n108 = n90 & n107;
  assign n109 = n84 & ~n88;
  assign n110 = n80 & n109;
  assign n111 = n101 & n105;
  assign n112 = n94 & n111;
  assign n113 = n110 & n112;
  assign n114 = ~n108 & ~n113;
  assign n115 = ~n101 & ~n105;
  assign n116 = n94 & n115;
  assign n117 = n76 & ~n79;
  assign n118 = n89 & n117;
  assign n119 = n116 & n118;
  assign n120 = n101 & ~n105;
  assign n121 = n94 & n120;
  assign n122 = n84 & n88;
  assign n123 = n76 & n79;
  assign n124 = n122 & n123;
  assign n125 = n121 & n124;
  assign n126 = n109 & n123;
  assign n127 = n112 & n126;
  assign n128 = ~n76 & ~n79;
  assign n129 = n109 & n128;
  assign n130 = ~n94 & n111;
  assign n131 = n129 & n130;
  assign n132 = n122 & n128;
  assign n133 = n121 & n132;
  assign n134 = n130 & n132;
  assign n135 = ~n133 & ~n134;
  assign n136 = ~n131 & n135;
  assign n137 = ~n84 & n88;
  assign n138 = n80 & n137;
  assign n139 = n94 & n106;
  assign n140 = n138 & n139;
  assign n141 = n89 & n128;
  assign n142 = n112 & n141;
  assign n143 = n128 & n137;
  assign n144 = n130 & n143;
  assign n145 = n107 & n124;
  assign n146 = ~n144 & ~n145;
  assign n147 = n116 & n141;
  assign n148 = ~n94 & n115;
  assign n149 = n124 & n148;
  assign n150 = ~n147 & ~n149;
  assign n151 = n80 & n122;
  assign n152 = n121 & n151;
  assign n153 = n123 & n137;
  assign n154 = n120 & n153;
  assign n155 = n94 & n154;
  assign n156 = ~n152 & ~n155;
  assign n157 = n129 & n139;
  assign n158 = n121 & n143;
  assign n159 = ~n157 & ~n158;
  assign n160 = n150 & n156;
  assign n161 = n159 & n160;
  assign n162 = ~n119 & ~n125;
  assign n163 = ~n127 & ~n140;
  assign n164 = ~n142 & n163;
  assign n165 = n114 & n162;
  assign n166 = n146 & n165;
  assign n167 = n136 & n164;
  assign n168 = n166 & n167;
  assign n169 = n161 & n168;
  assign n170 = n110 & n120;
  assign n171 = ~n94 & n170;
  assign n172 = ~n94 & n120;
  assign n173 = n117 & n137;
  assign n174 = n172 & n173;
  assign n175 = n109 & n117;
  assign n176 = n121 & n175;
  assign n177 = ~n171 & ~n174;
  assign n178 = ~n176 & n177;
  assign n179 = n117 & n122;
  assign n180 = n107 & n179;
  assign n181 = n132 & n172;
  assign n182 = n129 & n172;
  assign n183 = ~n181 & ~n182;
  assign n184 = ~n180 & n183;
  assign n185 = n130 & n173;
  assign n186 = n112 & n138;
  assign n187 = ~n185 & ~n186;
  assign n188 = n130 & n175;
  assign n189 = n139 & n153;
  assign n190 = n126 & n172;
  assign n191 = n89 & n123;
  assign n192 = n172 & n191;
  assign n193 = ~n188 & ~n189;
  assign n194 = ~n190 & ~n192;
  assign n195 = n193 & n194;
  assign n196 = n126 & n139;
  assign n197 = n130 & n138;
  assign n198 = n139 & n143;
  assign n199 = n112 & n124;
  assign n200 = n116 & n124;
  assign n201 = n107 & n175;
  assign n202 = ~n196 & ~n197;
  assign n203 = ~n198 & ~n199;
  assign n204 = ~n200 & ~n201;
  assign n205 = n203 & n204;
  assign n206 = n202 & n205;
  assign n207 = n107 & n141;
  assign n208 = n116 & n126;
  assign n209 = n107 & n173;
  assign n210 = n107 & n151;
  assign n211 = ~n209 & ~n210;
  assign n212 = ~n207 & ~n208;
  assign n213 = n187 & n212;
  assign n214 = n211 & n213;
  assign n215 = n184 & n195;
  assign n216 = n214 & n215;
  assign n217 = n206 & n216;
  assign n218 = n116 & n179;
  assign n219 = n116 & n175;
  assign n220 = n130 & n179;
  assign n221 = ~n219 & ~n220;
  assign n222 = n118 & n148;
  assign n223 = n112 & n153;
  assign n224 = n132 & n139;
  assign n225 = n110 & n139;
  assign n226 = n112 & n151;
  assign n227 = ~n218 & ~n222;
  assign n228 = ~n223 & ~n224;
  assign n229 = ~n225 & ~n226;
  assign n230 = n228 & n229;
  assign n231 = n221 & n227;
  assign n232 = n230 & n231;
  assign n233 = n141 & n172;
  assign n234 = n118 & n139;
  assign n235 = n90 & n111;
  assign n236 = ~n94 & n235;
  assign n237 = n141 & n148;
  assign n238 = n112 & n191;
  assign n239 = ~n237 & ~n238;
  assign n240 = n106 & n191;
  assign n241 = ~n94 & n240;
  assign n242 = ~n233 & ~n234;
  assign n243 = ~n236 & ~n241;
  assign n244 = n242 & n243;
  assign n245 = n239 & n244;
  assign n246 = n120 & n138;
  assign n247 = n116 & n132;
  assign n248 = n118 & n130;
  assign n249 = n148 & n179;
  assign n250 = n132 & n148;
  assign n251 = n107 & n143;
  assign n252 = ~n249 & ~n250;
  assign n253 = ~n251 & n252;
  assign n254 = ~n246 & ~n247;
  assign n255 = ~n248 & n254;
  assign n256 = n178 & n255;
  assign n257 = n253 & n256;
  assign n258 = n232 & n245;
  assign n259 = n257 & n258;
  assign n260 = n169 & n259;
  assign n261 = n217 & n260;
  assign n262 = n116 & n173;
  assign n263 = n148 & n153;
  assign n264 = n121 & n173;
  assign n265 = ~n263 & ~n264;
  assign n266 = ~n262 & n265;
  assign n267 = n139 & n151;
  assign n268 = n110 & n148;
  assign n269 = ~n226 & ~n267;
  assign n270 = ~n268 & n269;
  assign n271 = n107 & n126;
  assign n272 = n126 & n130;
  assign n273 = n151 & n172;
  assign n274 = n90 & n139;
  assign n275 = ~n271 & ~n272;
  assign n276 = ~n273 & ~n274;
  assign n277 = n275 & n276;
  assign n278 = ~n155 & ~n234;
  assign n279 = n94 & n170;
  assign n280 = ~n94 & n246;
  assign n281 = ~n186 & ~n280;
  assign n282 = n126 & n148;
  assign n283 = n115 & n151;
  assign n284 = n94 & n283;
  assign n285 = ~n108 & ~n282;
  assign n286 = ~n284 & n285;
  assign n287 = ~n222 & ~n279;
  assign n288 = n278 & n287;
  assign n289 = n281 & n288;
  assign n290 = n266 & n270;
  assign n291 = n277 & n286;
  assign n292 = n290 & n291;
  assign n293 = n289 & n292;
  assign n294 = n139 & n173;
  assign n295 = n121 & n126;
  assign n296 = ~n171 & ~n295;
  assign n297 = n130 & n191;
  assign n298 = n110 & n130;
  assign n299 = n94 & n246;
  assign n300 = ~n225 & ~n299;
  assign n301 = ~n248 & ~n298;
  assign n302 = n300 & n301;
  assign n303 = n124 & n172;
  assign n304 = n110 & n116;
  assign n305 = ~n303 & ~n304;
  assign n306 = n90 & n148;
  assign n307 = n116 & n138;
  assign n308 = ~n119 & ~n307;
  assign n309 = n139 & n141;
  assign n310 = n112 & n129;
  assign n311 = n139 & n179;
  assign n312 = ~n197 & ~n311;
  assign n313 = n115 & n191;
  assign n314 = ~n94 & n313;
  assign n315 = n148 & n173;
  assign n316 = ~n250 & ~n315;
  assign n317 = n130 & n141;
  assign n318 = n121 & n129;
  assign n319 = ~n158 & ~n318;
  assign n320 = ~n314 & ~n317;
  assign n321 = n312 & n320;
  assign n322 = n316 & n319;
  assign n323 = n321 & n322;
  assign n324 = n138 & n148;
  assign n325 = n148 & n175;
  assign n326 = ~n324 & ~n325;
  assign n327 = n94 & n313;
  assign n328 = n326 & ~n327;
  assign n329 = n116 & n153;
  assign n330 = ~n189 & ~n207;
  assign n331 = ~n182 & ~n247;
  assign n332 = ~n309 & ~n310;
  assign n333 = ~n329 & n332;
  assign n334 = n308 & n331;
  assign n335 = n330 & n334;
  assign n336 = n328 & n333;
  assign n337 = n335 & n336;
  assign n338 = n323 & n337;
  assign n339 = ~n199 & ~n306;
  assign n340 = n338 & n339;
  assign n341 = n112 & n175;
  assign n342 = n112 & n118;
  assign n343 = n172 & n175;
  assign n344 = ~n342 & ~n343;
  assign n345 = n107 & n138;
  assign n346 = ~n157 & ~n345;
  assign n347 = ~n131 & ~n174;
  assign n348 = ~n223 & ~n341;
  assign n349 = n344 & n348;
  assign n350 = n346 & n347;
  assign n351 = n349 & n350;
  assign n352 = n211 & n351;
  assign n353 = ~n94 & n283;
  assign n354 = ~n190 & ~n353;
  assign n355 = n90 & n116;
  assign n356 = n107 & n132;
  assign n357 = ~n355 & ~n356;
  assign n358 = ~n180 & ~n188;
  assign n359 = ~n294 & ~n297;
  assign n360 = n358 & n359;
  assign n361 = n296 & n305;
  assign n362 = n354 & n357;
  assign n363 = n361 & n362;
  assign n364 = n302 & n360;
  assign n365 = n363 & n364;
  assign n366 = n352 & n365;
  assign n367 = n293 & n366;
  assign n368 = n340 & n367;
  assign n369 = ~n261 & ~n368;
  assign n370 = n112 & n173;
  assign n371 = ~n170 & ~n297;
  assign n372 = n107 & n118;
  assign n373 = ~n236 & ~n248;
  assign n374 = ~n372 & n373;
  assign n375 = ~n263 & ~n306;
  assign n376 = ~n314 & n375;
  assign n377 = n94 & n235;
  assign n378 = n112 & n143;
  assign n379 = ~n185 & ~n378;
  assign n380 = n115 & n129;
  assign n381 = ~n377 & ~n380;
  assign n382 = n379 & n381;
  assign n383 = ~n238 & ~n271;
  assign n384 = n121 & n191;
  assign n385 = ~n180 & ~n268;
  assign n386 = ~n133 & ~n284;
  assign n387 = ~n353 & ~n384;
  assign n388 = n383 & n387;
  assign n389 = n385 & n386;
  assign n390 = n388 & n389;
  assign n391 = ~n158 & ~n307;
  assign n392 = ~n370 & n391;
  assign n393 = n371 & n392;
  assign n394 = n374 & n376;
  assign n395 = n382 & n394;
  assign n396 = n390 & n393;
  assign n397 = n395 & n396;
  assign n398 = ~n182 & ~n189;
  assign n399 = ~n94 & n154;
  assign n400 = ~n199 & ~n299;
  assign n401 = ~n399 & n400;
  assign n402 = n398 & n401;
  assign n403 = n124 & n139;
  assign n404 = ~n196 & ~n403;
  assign n405 = n130 & n153;
  assign n406 = n357 & ~n405;
  assign n407 = n404 & n406;
  assign n408 = ~n327 & ~n329;
  assign n409 = ~n317 & ~n324;
  assign n410 = n346 & n408;
  assign n411 = n409 & n410;
  assign n412 = n116 & n143;
  assign n413 = ~n208 & ~n412;
  assign n414 = ~n140 & ~n304;
  assign n415 = ~n144 & ~n147;
  assign n416 = ~n237 & ~n280;
  assign n417 = ~n282 & n416;
  assign n418 = n413 & n415;
  assign n419 = n414 & n418;
  assign n420 = n417 & n419;
  assign n421 = n411 & n420;
  assign n422 = ~n149 & ~n224;
  assign n423 = n421 & n422;
  assign n424 = ~n145 & ~n274;
  assign n425 = ~n311 & n424;
  assign n426 = ~n273 & ~n342;
  assign n427 = n118 & n120;
  assign n428 = n94 & n427;
  assign n429 = n107 & n110;
  assign n430 = ~n152 & ~n318;
  assign n431 = ~n428 & ~n429;
  assign n432 = n430 & n431;
  assign n433 = n143 & n148;
  assign n434 = ~n181 & ~n192;
  assign n435 = ~n433 & n434;
  assign n436 = ~n94 & n427;
  assign n437 = ~n108 & ~n200;
  assign n438 = ~n226 & ~n436;
  assign n439 = n437 & n438;
  assign n440 = n435 & n439;
  assign n441 = ~n142 & n426;
  assign n442 = n425 & n441;
  assign n443 = n432 & n442;
  assign n444 = n402 & n407;
  assign n445 = n440 & n444;
  assign n446 = n443 & n445;
  assign n447 = n397 & n446;
  assign n448 = n423 & n447;
  assign n449 = ~n369 & ~n448;
  assign n450 = ~pi22  & ~n62;
  assign n451 = ~pi9  & ~n450;
  assign n452 = pi9  & n450;
  assign n453 = ~n451 & ~n452;
  assign n454 = ~n94 & n380;
  assign n455 = ~n233 & ~n454;
  assign n456 = ~n200 & ~n384;
  assign n457 = n143 & n172;
  assign n458 = n121 & n141;
  assign n459 = ~n457 & ~n458;
  assign n460 = ~n412 & n459;
  assign n461 = n94 & n380;
  assign n462 = ~n149 & ~n154;
  assign n463 = ~n192 & ~n208;
  assign n464 = ~n461 & n463;
  assign n465 = n455 & n462;
  assign n466 = n456 & n465;
  assign n467 = n460 & n464;
  assign n468 = n466 & n467;
  assign n469 = n90 & n121;
  assign n470 = ~n314 & ~n469;
  assign n471 = ~n246 & ~n283;
  assign n472 = n470 & n471;
  assign n473 = ~n147 & ~n247;
  assign n474 = ~n295 & ~n433;
  assign n475 = n473 & n474;
  assign n476 = ~n125 & ~n237;
  assign n477 = ~n303 & n476;
  assign n478 = ~n190 & ~n250;
  assign n479 = n475 & n478;
  assign n480 = n477 & n479;
  assign n481 = n90 & n172;
  assign n482 = ~n218 & ~n481;
  assign n483 = ~n119 & ~n273;
  assign n484 = ~n222 & ~n327;
  assign n485 = ~n171 & ~n263;
  assign n486 = ~n329 & n485;
  assign n487 = n483 & n484;
  assign n488 = n486 & n487;
  assign n489 = ~n152 & ~n279;
  assign n490 = n488 & n489;
  assign n491 = ~n249 & ~n268;
  assign n492 = ~n219 & ~n282;
  assign n493 = ~n304 & ~n307;
  assign n494 = n492 & n493;
  assign n495 = n482 & n491;
  assign n496 = n494 & n495;
  assign n497 = n480 & n496;
  assign n498 = n490 & n497;
  assign n499 = ~n90 & ~n173;
  assign n500 = n115 & ~n499;
  assign n501 = n326 & ~n500;
  assign n502 = n472 & n501;
  assign n503 = n468 & n502;
  assign n504 = n498 & n503;
  assign n505 = n453 & ~n504;
  assign n506 = ~n449 & n505;
  assign n507 = pi10  & pi22 ;
  assign n508 = ~pi22  & ~n64;
  assign n509 = pi10  & ~n63;
  assign n510 = n508 & ~n509;
  assign n511 = ~n507 & ~n510;
  assign n512 = ~n504 & ~n511;
  assign n513 = n449 & ~n505;
  assign n514 = ~n506 & ~n513;
  assign n515 = n512 & n514;
  assign n516 = ~n506 & ~n515;
  assign n517 = ~pi11  & ~n508;
  assign n518 = pi11  & n508;
  assign n519 = ~n517 & ~n518;
  assign n520 = n130 & n151;
  assign n521 = ~n298 & ~n520;
  assign n522 = ~n133 & ~n318;
  assign n523 = ~n113 & ~n235;
  assign n524 = ~n186 & n523;
  assign n525 = n312 & n521;
  assign n526 = n522 & n525;
  assign n527 = n184 & n524;
  assign n528 = n526 & n527;
  assign n529 = ~n226 & ~n238;
  assign n530 = ~n297 & ~n405;
  assign n531 = n529 & n530;
  assign n532 = n528 & n531;
  assign n533 = ~n210 & ~n429;
  assign n534 = ~n225 & n533;
  assign n535 = ~n240 & ~n345;
  assign n536 = n534 & n535;
  assign n537 = n107 & n153;
  assign n538 = ~n108 & ~n140;
  assign n539 = ~n176 & ~n428;
  assign n540 = ~n537 & n539;
  assign n541 = n538 & n540;
  assign n542 = n121 & n179;
  assign n543 = ~n158 & ~n274;
  assign n544 = ~n264 & ~n436;
  assign n545 = ~n174 & ~n343;
  assign n546 = n172 & n179;
  assign n547 = ~n267 & ~n546;
  assign n548 = ~n542 & n543;
  assign n549 = n544 & n545;
  assign n550 = n547 & n549;
  assign n551 = n548 & n550;
  assign n552 = n536 & n541;
  assign n553 = n551 & n552;
  assign n554 = n124 & n130;
  assign n555 = ~n127 & ~n554;
  assign n556 = ~n223 & ~n272;
  assign n557 = n555 & n556;
  assign n558 = n532 & n557;
  assign n559 = n553 & n558;
  assign n560 = n107 & n129;
  assign n561 = ~n198 & ~n309;
  assign n562 = ~n560 & n561;
  assign n563 = ~n145 & ~n251;
  assign n564 = ~n271 & n563;
  assign n565 = n330 & n404;
  assign n566 = n564 & n565;
  assign n567 = n562 & n566;
  assign n568 = n183 & n522;
  assign n569 = n567 & n568;
  assign n570 = n553 & n569;
  assign n571 = n139 & n175;
  assign n572 = ~n356 & ~n571;
  assign n573 = ~n201 & ~n234;
  assign n574 = ~n294 & n573;
  assign n575 = n572 & n574;
  assign n576 = ~n209 & ~n224;
  assign n577 = ~n372 & n576;
  assign n578 = n575 & n577;
  assign n579 = ~n157 & n578;
  assign n580 = n570 & n579;
  assign n581 = n559 & n580;
  assign n582 = ~n559 & ~n580;
  assign n583 = ~n581 & ~n582;
  assign n584 = n504 & ~n559;
  assign n585 = ~n583 & ~n584;
  assign n586 = n519 & n585;
  assign n587 = ~n504 & ~n582;
  assign n588 = ~n583 & ~n587;
  assign n589 = ~n519 & n588;
  assign n590 = pi12  & pi22 ;
  assign n591 = ~pi22  & ~n66;
  assign n592 = pi12  & ~n65;
  assign n593 = n591 & ~n592;
  assign n594 = ~n590 & ~n593;
  assign n595 = ~n504 & ~n594;
  assign n596 = n504 & n594;
  assign n597 = ~n595 & ~n596;
  assign n598 = n583 & ~n597;
  assign n599 = ~n586 & ~n598;
  assign n600 = ~n589 & n599;
  assign n601 = pi14  & pi22 ;
  assign n602 = pi14  & ~n67;
  assign n603 = n91 & ~n602;
  assign n604 = ~n601 & ~n603;
  assign n605 = ~n176 & ~n481;
  assign n606 = ~n144 & ~n236;
  assign n607 = ~n304 & ~n454;
  assign n608 = n606 & n607;
  assign n609 = n605 & n608;
  assign n610 = n266 & n609;
  assign n611 = ~n222 & ~n343;
  assign n612 = n610 & n611;
  assign n613 = ~n436 & ~n560;
  assign n614 = ~n145 & ~n198;
  assign n615 = ~n134 & ~n186;
  assign n616 = ~n180 & ~n282;
  assign n617 = ~n378 & ~n433;
  assign n618 = n616 & n617;
  assign n619 = n413 & n614;
  assign n620 = n615 & n619;
  assign n621 = n618 & n620;
  assign n622 = ~n428 & ~n520;
  assign n623 = n112 & n132;
  assign n624 = ~n200 & ~n219;
  assign n625 = ~n403 & n624;
  assign n626 = ~n249 & ~n461;
  assign n627 = ~n237 & ~n271;
  assign n628 = n626 & n627;
  assign n629 = ~n131 & ~n181;
  assign n630 = ~n546 & ~n623;
  assign n631 = n629 & n630;
  assign n632 = n622 & n631;
  assign n633 = n625 & n628;
  assign n634 = n632 & n633;
  assign n635 = n621 & n634;
  assign n636 = n340 & n635;
  assign n637 = ~n113 & ~n542;
  assign n638 = n150 & ~n298;
  assign n639 = ~n218 & ~n469;
  assign n640 = ~n196 & ~n268;
  assign n641 = ~n174 & ~n251;
  assign n642 = ~n353 & ~n355;
  assign n643 = n641 & n642;
  assign n644 = n639 & n640;
  assign n645 = n643 & n644;
  assign n646 = ~n142 & ~n377;
  assign n647 = n386 & n646;
  assign n648 = n613 & n637;
  assign n649 = n647 & n648;
  assign n650 = n638 & n649;
  assign n651 = n645 & n650;
  assign n652 = n612 & n651;
  assign n653 = n636 & n652;
  assign n654 = n448 & n653;
  assign n655 = ~n448 & ~n653;
  assign n656 = ~n654 & ~n655;
  assign n657 = ~n559 & n656;
  assign n658 = ~n604 & n657;
  assign n659 = n559 & n656;
  assign n660 = n604 & n659;
  assign n661 = ~pi13  & ~n591;
  assign n662 = pi13  & n591;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~n559 & ~n655;
  assign n665 = ~n656 & ~n664;
  assign n666 = ~n663 & n665;
  assign n667 = ~n448 & n559;
  assign n668 = ~n656 & ~n667;
  assign n669 = n663 & n668;
  assign n670 = ~n658 & ~n660;
  assign n671 = ~n666 & ~n669;
  assign n672 = n670 & n671;
  assign n673 = n600 & n672;
  assign n674 = n261 & n368;
  assign n675 = ~n369 & ~n674;
  assign n676 = ~n604 & ~n675;
  assign n677 = ~n449 & ~n676;
  assign n678 = ~n261 & n448;
  assign n679 = ~n675 & ~n678;
  assign n680 = ~n604 & n679;
  assign n681 = ~n677 & ~n680;
  assign n682 = ~n505 & n681;
  assign n683 = n505 & ~n681;
  assign n684 = ~n682 & ~n683;
  assign n685 = n657 & n663;
  assign n686 = n659 & ~n663;
  assign n687 = ~n594 & n668;
  assign n688 = n594 & n665;
  assign n689 = ~n685 & ~n686;
  assign n690 = ~n687 & ~n688;
  assign n691 = n689 & n690;
  assign n692 = n684 & n691;
  assign n693 = ~n682 & ~n692;
  assign n694 = ~n600 & ~n672;
  assign n695 = ~n673 & ~n694;
  assign n696 = ~n693 & n695;
  assign n697 = ~n673 & ~n696;
  assign n698 = ~n516 & ~n697;
  assign n699 = ~n504 & n519;
  assign n700 = ~n604 & ~n656;
  assign n701 = ~n664 & ~n700;
  assign n702 = ~n604 & n668;
  assign n703 = ~n701 & ~n702;
  assign n704 = ~n699 & n703;
  assign n705 = n699 & ~n703;
  assign n706 = ~n704 & ~n705;
  assign n707 = n585 & ~n594;
  assign n708 = n588 & n594;
  assign n709 = ~n504 & n663;
  assign n710 = n504 & ~n663;
  assign n711 = ~n709 & ~n710;
  assign n712 = n583 & ~n711;
  assign n713 = ~n707 & ~n712;
  assign n714 = ~n708 & n713;
  assign n715 = n706 & n714;
  assign n716 = ~n706 & ~n714;
  assign n717 = ~n715 & ~n716;
  assign n718 = n516 & n697;
  assign n719 = ~n698 & ~n718;
  assign n720 = n717 & n719;
  assign n721 = ~n698 & ~n720;
  assign n722 = ~n704 & ~n715;
  assign n723 = n585 & n663;
  assign n724 = n588 & ~n663;
  assign n725 = ~n504 & n604;
  assign n726 = n504 & ~n604;
  assign n727 = ~n725 & ~n726;
  assign n728 = n583 & n727;
  assign n729 = ~n723 & ~n728;
  assign n730 = ~n724 & n729;
  assign n731 = ~n722 & n730;
  assign n732 = n722 & ~n730;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~n664 & n699;
  assign n735 = n664 & ~n699;
  assign n736 = ~n734 & ~n735;
  assign n737 = n595 & n736;
  assign n738 = ~n595 & ~n736;
  assign n739 = ~n737 & ~n738;
  assign n740 = n733 & n739;
  assign n741 = ~n733 & ~n739;
  assign n742 = ~n740 & ~n741;
  assign n743 = ~n721 & n742;
  assign n744 = ~pi22  & ~n60;
  assign n745 = ~pi7  & ~n744;
  assign n746 = pi7  & n744;
  assign n747 = ~n745 & ~n746;
  assign n748 = ~n504 & n747;
  assign n749 = ~n225 & ~n546;
  assign n750 = ~n142 & ~n185;
  assign n751 = ~n297 & n750;
  assign n752 = n414 & n749;
  assign n753 = n751 & n752;
  assign n754 = ~n226 & ~n384;
  assign n755 = ~n155 & n221;
  assign n756 = n754 & n755;
  assign n757 = ~n108 & ~n454;
  assign n758 = ~n307 & ~n315;
  assign n759 = ~n457 & n758;
  assign n760 = ~n233 & ~n469;
  assign n761 = ~n234 & ~n403;
  assign n762 = n757 & n760;
  assign n763 = n761 & n762;
  assign n764 = n759 & n763;
  assign n765 = ~n251 & ~n267;
  assign n766 = ~n201 & ~n207;
  assign n767 = ~n273 & ~n317;
  assign n768 = ~n327 & ~n355;
  assign n769 = n767 & n768;
  assign n770 = n765 & n766;
  assign n771 = n769 & n770;
  assign n772 = n753 & n771;
  assign n773 = n756 & n772;
  assign n774 = n764 & n773;
  assign n775 = n94 & n240;
  assign n776 = ~n306 & ~n775;
  assign n777 = ~n197 & n776;
  assign n778 = ~n199 & ~n250;
  assign n779 = ~n324 & n778;
  assign n780 = n112 & n179;
  assign n781 = ~n190 & ~n780;
  assign n782 = ~n174 & ~n370;
  assign n783 = ~n264 & ~n274;
  assign n784 = n555 & n783;
  assign n785 = ~n208 & ~n458;
  assign n786 = ~n157 & ~n295;
  assign n787 = ~n189 & ~n263;
  assign n788 = ~n342 & ~n377;
  assign n789 = n787 & n788;
  assign n790 = n477 & n789;
  assign n791 = ~n222 & n640;
  assign n792 = n785 & n786;
  assign n793 = n791 & n792;
  assign n794 = n374 & n784;
  assign n795 = n793 & n794;
  assign n796 = n790 & n795;
  assign n797 = ~n133 & ~n152;
  assign n798 = ~n188 & ~n249;
  assign n799 = ~n280 & ~n399;
  assign n800 = ~n520 & n799;
  assign n801 = n797 & n798;
  assign n802 = n800 & n801;
  assign n803 = ~n341 & ~n481;
  assign n804 = n572 & n803;
  assign n805 = n781 & n782;
  assign n806 = n804 & n805;
  assign n807 = n435 & n777;
  assign n808 = n779 & n807;
  assign n809 = n802 & n806;
  assign n810 = n808 & n809;
  assign n811 = n796 & n810;
  assign n812 = n774 & n811;
  assign n813 = ~n219 & ~n247;
  assign n814 = ~n149 & ~n279;
  assign n815 = ~n306 & n814;
  assign n816 = n813 & n815;
  assign n817 = ~n284 & ~n307;
  assign n818 = ~n355 & ~n429;
  assign n819 = n817 & n818;
  assign n820 = ~n262 & ~n272;
  assign n821 = ~n433 & n820;
  assign n822 = n300 & n385;
  assign n823 = n605 & n822;
  assign n824 = n784 & n821;
  assign n825 = n819 & n824;
  assign n826 = n816 & n823;
  assign n827 = n825 & n826;
  assign n828 = ~n200 & ~n353;
  assign n829 = ~n142 & ~n199;
  assign n830 = n828 & n829;
  assign n831 = n827 & n830;
  assign n832 = ~n324 & ~n372;
  assign n833 = ~n241 & ~n271;
  assign n834 = ~n436 & n833;
  assign n835 = ~n224 & ~n309;
  assign n836 = n156 & n832;
  assign n837 = n835 & n836;
  assign n838 = n834 & n837;
  assign n839 = ~n236 & ~n405;
  assign n840 = ~n125 & ~n280;
  assign n841 = ~n223 & n840;
  assign n842 = ~n458 & ~n546;
  assign n843 = ~n234 & ~n304;
  assign n844 = n839 & n843;
  assign n845 = n842 & n844;
  assign n846 = n841 & n845;
  assign n847 = ~n251 & ~n775;
  assign n848 = ~n384 & n847;
  assign n849 = ~n181 & ~n238;
  assign n850 = n848 & n849;
  assign n851 = ~n196 & ~n295;
  assign n852 = ~n377 & n851;
  assign n853 = n413 & n852;
  assign n854 = n323 & n853;
  assign n855 = n850 & n854;
  assign n856 = n838 & n846;
  assign n857 = n855 & n856;
  assign n858 = n831 & n857;
  assign n859 = ~n812 & ~n858;
  assign n860 = ~n261 & ~n859;
  assign n861 = n748 & ~n860;
  assign n862 = ~n748 & n860;
  assign n863 = ~n861 & ~n862;
  assign n864 = pi8  & pi22 ;
  assign n865 = pi8  & ~n61;
  assign n866 = n450 & ~n865;
  assign n867 = ~n864 & ~n866;
  assign n868 = ~n504 & ~n867;
  assign n869 = n863 & n868;
  assign n870 = ~n861 & ~n869;
  assign n871 = ~n511 & n585;
  assign n872 = n511 & n588;
  assign n873 = n504 & ~n519;
  assign n874 = ~n699 & ~n873;
  assign n875 = n583 & ~n874;
  assign n876 = ~n871 & ~n875;
  assign n877 = ~n872 & n876;
  assign n878 = ~n870 & n877;
  assign n879 = ~n448 & n675;
  assign n880 = ~n604 & n879;
  assign n881 = n448 & n675;
  assign n882 = n604 & n881;
  assign n883 = ~n449 & ~n675;
  assign n884 = ~n663 & n883;
  assign n885 = n663 & n679;
  assign n886 = ~n880 & ~n882;
  assign n887 = ~n884 & ~n885;
  assign n888 = n886 & n887;
  assign n889 = ~n594 & n657;
  assign n890 = n594 & n659;
  assign n891 = ~n519 & n665;
  assign n892 = n519 & n668;
  assign n893 = ~n889 & ~n890;
  assign n894 = ~n891 & ~n892;
  assign n895 = n893 & n894;
  assign n896 = n888 & n895;
  assign n897 = ~n888 & ~n895;
  assign n898 = ~n896 & ~n897;
  assign n899 = n453 & n585;
  assign n900 = ~n453 & n588;
  assign n901 = n504 & n511;
  assign n902 = ~n512 & ~n901;
  assign n903 = n583 & ~n902;
  assign n904 = ~n899 & ~n903;
  assign n905 = ~n900 & n904;
  assign n906 = n898 & n905;
  assign n907 = ~n896 & ~n906;
  assign n908 = n870 & ~n877;
  assign n909 = ~n878 & ~n908;
  assign n910 = ~n907 & n909;
  assign n911 = ~n878 & ~n910;
  assign n912 = ~n512 & ~n514;
  assign n913 = ~n515 & ~n912;
  assign n914 = ~n911 & n913;
  assign n915 = n911 & ~n913;
  assign n916 = ~n914 & ~n915;
  assign n917 = n693 & ~n695;
  assign n918 = ~n696 & ~n917;
  assign n919 = n916 & n918;
  assign n920 = ~n914 & ~n919;
  assign n921 = ~n717 & ~n719;
  assign n922 = ~n720 & ~n921;
  assign n923 = ~n920 & n922;
  assign n924 = n585 & ~n867;
  assign n925 = n588 & n867;
  assign n926 = ~n453 & n504;
  assign n927 = ~n505 & ~n926;
  assign n928 = n583 & ~n927;
  assign n929 = ~n924 & ~n928;
  assign n930 = ~n925 & n929;
  assign n931 = n519 & n657;
  assign n932 = ~n519 & n659;
  assign n933 = ~n511 & n668;
  assign n934 = n511 & n665;
  assign n935 = ~n931 & ~n932;
  assign n936 = ~n933 & ~n934;
  assign n937 = n935 & n936;
  assign n938 = n930 & n937;
  assign n939 = ~n930 & ~n937;
  assign n940 = ~n938 & ~n939;
  assign n941 = ~n113 & ~n196;
  assign n942 = ~n353 & ~n428;
  assign n943 = n941 & n942;
  assign n944 = ~n158 & ~n201;
  assign n945 = ~n571 & n944;
  assign n946 = ~n299 & ~n370;
  assign n947 = ~n546 & n946;
  assign n948 = ~n108 & ~n355;
  assign n949 = ~n405 & ~n458;
  assign n950 = n948 & n949;
  assign n951 = n346 & n950;
  assign n952 = n943 & n945;
  assign n953 = n947 & n952;
  assign n954 = n816 & n951;
  assign n955 = n953 & n954;
  assign n956 = ~n303 & ~n315;
  assign n957 = ~n272 & ~n623;
  assign n958 = ~n250 & ~n412;
  assign n959 = ~n152 & ~n207;
  assign n960 = ~n220 & ~n294;
  assign n961 = ~n554 & n960;
  assign n962 = n491 & n959;
  assign n963 = n544 & n962;
  assign n964 = n961 & n963;
  assign n965 = ~n145 & ~n181;
  assign n966 = ~n210 & ~n237;
  assign n967 = ~n295 & ~n297;
  assign n968 = n966 & n967;
  assign n969 = n347 & n965;
  assign n970 = n386 & n765;
  assign n971 = n969 & n970;
  assign n972 = n968 & n971;
  assign n973 = ~n356 & ~n537;
  assign n974 = ~n154 & ~n197;
  assign n975 = ~n240 & n973;
  assign n976 = n974 & n975;
  assign n977 = ~n119 & ~n142;
  assign n978 = ~n209 & ~n225;
  assign n979 = ~n280 & n978;
  assign n980 = n781 & n977;
  assign n981 = n956 & n957;
  assign n982 = n958 & n981;
  assign n983 = n979 & n980;
  assign n984 = n382 & n983;
  assign n985 = n976 & n982;
  assign n986 = n984 & n985;
  assign n987 = n964 & n972;
  assign n988 = n986 & n987;
  assign n989 = n955 & n988;
  assign n990 = n812 & n989;
  assign n991 = ~n271 & ~n355;
  assign n992 = ~n306 & ~n433;
  assign n993 = n354 & n992;
  assign n994 = n545 & n957;
  assign n995 = n993 & n994;
  assign n996 = ~n234 & ~n307;
  assign n997 = ~n310 & ~n329;
  assign n998 = ~n542 & n997;
  assign n999 = n455 & n996;
  assign n1000 = n991 & n999;
  assign n1001 = n638 & n998;
  assign n1002 = n779 & n1001;
  assign n1003 = n976 & n1000;
  assign n1004 = n995 & n1003;
  assign n1005 = n1002 & n1004;
  assign n1006 = ~n341 & ~n780;
  assign n1007 = ~n134 & ~n223;
  assign n1008 = ~n249 & ~n325;
  assign n1009 = ~n142 & ~n295;
  assign n1010 = ~n158 & ~n188;
  assign n1011 = n639 & n1010;
  assign n1012 = n754 & n1008;
  assign n1013 = n1009 & n1012;
  assign n1014 = n1011 & n1013;
  assign n1015 = ~n192 & ~n220;
  assign n1016 = ~n303 & ~n317;
  assign n1017 = n1015 & n1016;
  assign n1018 = n183 & n371;
  assign n1019 = n840 & n1006;
  assign n1020 = n1007 & n1019;
  assign n1021 = n1017 & n1018;
  assign n1022 = n1020 & n1021;
  assign n1023 = n1014 & n1022;
  assign n1024 = ~n140 & ~n247;
  assign n1025 = ~n267 & ~n461;
  assign n1026 = n1024 & n1025;
  assign n1027 = ~n294 & ~n311;
  assign n1028 = n613 & n1027;
  assign n1029 = n835 & n1028;
  assign n1030 = n114 & ~n571;
  assign n1031 = n330 & n413;
  assign n1032 = n484 & n1031;
  assign n1033 = n534 & n1030;
  assign n1034 = n1026 & n1033;
  assign n1035 = n1029 & n1032;
  assign n1036 = n1034 & n1035;
  assign n1037 = n1023 & n1036;
  assign n1038 = n1005 & n1037;
  assign n1039 = ~n989 & ~n1038;
  assign n1040 = ~n812 & ~n1039;
  assign n1041 = ~n989 & n1040;
  assign n1042 = pi6  & pi22 ;
  assign n1043 = pi6  & ~n59;
  assign n1044 = n744 & ~n1043;
  assign n1045 = ~n1042 & ~n1044;
  assign n1046 = ~n504 & ~n1045;
  assign n1047 = ~n1041 & n1046;
  assign n1048 = ~n990 & ~n1047;
  assign n1049 = n940 & ~n1048;
  assign n1050 = ~n938 & ~n1049;
  assign n1051 = n812 & n858;
  assign n1052 = ~n859 & ~n1051;
  assign n1053 = ~n604 & ~n1052;
  assign n1054 = ~n860 & ~n1053;
  assign n1055 = n261 & ~n1051;
  assign n1056 = n1053 & ~n1055;
  assign n1057 = ~n1054 & ~n1056;
  assign n1058 = ~n748 & n1057;
  assign n1059 = n748 & ~n1057;
  assign n1060 = ~n1058 & ~n1059;
  assign n1061 = n663 & n879;
  assign n1062 = ~n663 & n881;
  assign n1063 = ~n594 & n679;
  assign n1064 = n594 & n883;
  assign n1065 = ~n1061 & ~n1062;
  assign n1066 = ~n1063 & ~n1064;
  assign n1067 = n1065 & n1066;
  assign n1068 = n1060 & n1067;
  assign n1069 = ~n1058 & ~n1068;
  assign n1070 = ~n1050 & ~n1069;
  assign n1071 = ~n863 & ~n868;
  assign n1072 = ~n869 & ~n1071;
  assign n1073 = n1050 & n1069;
  assign n1074 = ~n1070 & ~n1073;
  assign n1075 = n1072 & n1074;
  assign n1076 = ~n1070 & ~n1075;
  assign n1077 = ~n684 & ~n691;
  assign n1078 = ~n692 & ~n1077;
  assign n1079 = ~n1076 & n1078;
  assign n1080 = n1076 & ~n1078;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = n907 & ~n909;
  assign n1083 = ~n910 & ~n1082;
  assign n1084 = n1081 & n1083;
  assign n1085 = ~n1079 & ~n1084;
  assign n1086 = ~n916 & ~n918;
  assign n1087 = ~n919 & ~n1086;
  assign n1088 = ~n1085 & n1087;
  assign n1089 = n585 & n747;
  assign n1090 = n588 & ~n747;
  assign n1091 = n504 & n867;
  assign n1092 = ~n868 & ~n1091;
  assign n1093 = n583 & ~n1092;
  assign n1094 = ~n1089 & ~n1093;
  assign n1095 = ~n1090 & n1094;
  assign n1096 = ~n511 & n657;
  assign n1097 = n511 & n659;
  assign n1098 = ~n453 & n665;
  assign n1099 = n453 & n668;
  assign n1100 = ~n1096 & ~n1097;
  assign n1101 = ~n1098 & ~n1099;
  assign n1102 = n1100 & n1101;
  assign n1103 = n1095 & n1102;
  assign n1104 = ~n1095 & ~n1102;
  assign n1105 = ~n1103 & ~n1104;
  assign n1106 = ~n860 & ~n1052;
  assign n1107 = ~n663 & ~n1106;
  assign n1108 = ~n1052 & ~n1055;
  assign n1109 = n663 & ~n1108;
  assign n1110 = ~n1107 & ~n1109;
  assign n1111 = n860 & ~n1051;
  assign n1112 = ~n604 & n1111;
  assign n1113 = ~n859 & n1055;
  assign n1114 = n604 & n1113;
  assign n1115 = ~n1112 & ~n1114;
  assign n1116 = ~n1110 & n1115;
  assign n1117 = n1105 & n1116;
  assign n1118 = ~n1103 & ~n1117;
  assign n1119 = ~n1060 & ~n1067;
  assign n1120 = ~n1068 & ~n1119;
  assign n1121 = ~n1118 & n1120;
  assign n1122 = ~n940 & n1048;
  assign n1123 = ~n1049 & ~n1122;
  assign n1124 = n1118 & ~n1120;
  assign n1125 = ~n1121 & ~n1124;
  assign n1126 = n1123 & n1125;
  assign n1127 = ~n1121 & ~n1126;
  assign n1128 = ~n898 & ~n905;
  assign n1129 = ~n906 & ~n1128;
  assign n1130 = ~n1127 & n1129;
  assign n1131 = n1127 & ~n1129;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = ~n1072 & ~n1074;
  assign n1134 = ~n1075 & ~n1133;
  assign n1135 = n1132 & n1134;
  assign n1136 = ~n1130 & ~n1135;
  assign n1137 = ~n1081 & ~n1083;
  assign n1138 = ~n1084 & ~n1137;
  assign n1139 = ~n1136 & n1138;
  assign n1140 = ~n990 & ~n1041;
  assign n1141 = n1046 & ~n1140;
  assign n1142 = ~n1047 & n1140;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n594 & n879;
  assign n1145 = n594 & n881;
  assign n1146 = ~n519 & n883;
  assign n1147 = n519 & n679;
  assign n1148 = ~n1144 & ~n1145;
  assign n1149 = ~n1146 & ~n1147;
  assign n1150 = n1148 & n1149;
  assign n1151 = ~n1143 & n1150;
  assign n1152 = n57 & ~n504;
  assign n1153 = ~n989 & n1152;
  assign n1154 = n989 & ~n1152;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156 = n989 & n1038;
  assign n1157 = ~n1039 & ~n1156;
  assign n1158 = ~n604 & ~n1157;
  assign n1159 = ~n1040 & ~n1158;
  assign n1160 = n812 & ~n1156;
  assign n1161 = n1158 & ~n1160;
  assign n1162 = ~n1159 & ~n1161;
  assign n1163 = n1155 & n1162;
  assign n1164 = ~n1153 & ~n1163;
  assign n1165 = n1143 & ~n1150;
  assign n1166 = ~n1151 & ~n1165;
  assign n1167 = ~n1164 & n1166;
  assign n1168 = ~n1151 & ~n1167;
  assign n1169 = n594 & ~n1106;
  assign n1170 = ~n594 & ~n1108;
  assign n1171 = ~n1169 & ~n1170;
  assign n1172 = ~n663 & n1113;
  assign n1173 = n663 & n1111;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = ~n1171 & n1174;
  assign n1176 = n519 & n879;
  assign n1177 = ~n519 & n881;
  assign n1178 = ~n511 & n679;
  assign n1179 = n511 & n883;
  assign n1180 = ~n1176 & ~n1177;
  assign n1181 = ~n1178 & ~n1179;
  assign n1182 = n1180 & n1181;
  assign n1183 = n1175 & n1182;
  assign n1184 = ~n1175 & ~n1182;
  assign n1185 = ~n1183 & ~n1184;
  assign n1186 = n453 & n657;
  assign n1187 = ~n453 & n659;
  assign n1188 = n668 & ~n867;
  assign n1189 = n665 & n867;
  assign n1190 = ~n1186 & ~n1187;
  assign n1191 = ~n1188 & ~n1189;
  assign n1192 = n1190 & n1191;
  assign n1193 = n1185 & n1192;
  assign n1194 = ~n1183 & ~n1193;
  assign n1195 = ~n1105 & ~n1116;
  assign n1196 = ~n1117 & ~n1195;
  assign n1197 = ~n1194 & n1196;
  assign n1198 = pi4  & pi22 ;
  assign n1199 = pi4  & ~n52;
  assign n1200 = n54 & ~n1199;
  assign n1201 = ~n1198 & ~n1200;
  assign n1202 = ~n504 & ~n1201;
  assign n1203 = ~n989 & n1202;
  assign n1204 = n989 & ~n1202;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = ~n812 & n1039;
  assign n1207 = ~n1156 & ~n1206;
  assign n1208 = n663 & ~n1207;
  assign n1209 = ~n1040 & ~n1157;
  assign n1210 = ~n663 & n1209;
  assign n1211 = n1040 & ~n1156;
  assign n1212 = ~n604 & n1211;
  assign n1213 = ~n1039 & n1160;
  assign n1214 = n604 & n1213;
  assign n1215 = ~n1208 & ~n1210;
  assign n1216 = ~n1212 & ~n1214;
  assign n1217 = n1215 & n1216;
  assign n1218 = n1205 & n1217;
  assign n1219 = ~n1203 & ~n1218;
  assign n1220 = n585 & ~n1045;
  assign n1221 = n588 & n1045;
  assign n1222 = n504 & ~n747;
  assign n1223 = ~n748 & ~n1222;
  assign n1224 = n583 & ~n1223;
  assign n1225 = ~n1220 & ~n1224;
  assign n1226 = ~n1221 & n1225;
  assign n1227 = ~n1219 & n1226;
  assign n1228 = n1219 & ~n1226;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~n511 & n879;
  assign n1231 = n511 & n881;
  assign n1232 = ~n453 & n883;
  assign n1233 = n453 & n679;
  assign n1234 = ~n1230 & ~n1231;
  assign n1235 = ~n1232 & ~n1233;
  assign n1236 = n1234 & n1235;
  assign n1237 = ~n519 & ~n1106;
  assign n1238 = n519 & ~n1108;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = ~n594 & n1111;
  assign n1241 = n594 & n1113;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = ~n1239 & n1242;
  assign n1244 = n1236 & n1243;
  assign n1245 = ~n1236 & ~n1243;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = n657 & ~n867;
  assign n1248 = n659 & n867;
  assign n1249 = n665 & ~n747;
  assign n1250 = n668 & n747;
  assign n1251 = ~n1247 & ~n1248;
  assign n1252 = ~n1249 & ~n1250;
  assign n1253 = n1251 & n1252;
  assign n1254 = n1246 & n1253;
  assign n1255 = ~n1244 & ~n1254;
  assign n1256 = n1229 & ~n1255;
  assign n1257 = ~n1227 & ~n1256;
  assign n1258 = n1194 & ~n1196;
  assign n1259 = ~n1197 & ~n1258;
  assign n1260 = ~n1257 & n1259;
  assign n1261 = ~n1197 & ~n1260;
  assign n1262 = ~n1168 & ~n1261;
  assign n1263 = ~n1123 & ~n1125;
  assign n1264 = ~n1126 & ~n1263;
  assign n1265 = n1168 & n1261;
  assign n1266 = ~n1262 & ~n1265;
  assign n1267 = n1264 & n1266;
  assign n1268 = ~n1262 & ~n1267;
  assign n1269 = ~n1132 & ~n1134;
  assign n1270 = ~n1135 & ~n1269;
  assign n1271 = ~n1268 & n1270;
  assign n1272 = ~n1155 & ~n1162;
  assign n1273 = ~n1163 & ~n1272;
  assign n1274 = ~n1185 & ~n1192;
  assign n1275 = ~n1193 & ~n1274;
  assign n1276 = n1273 & n1275;
  assign n1277 = ~pi22  & ~n51;
  assign n1278 = ~pi3  & ~n1277;
  assign n1279 = pi3  & n1277;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = ~n504 & n1280;
  assign n1282 = n278 & ~n433;
  assign n1283 = ~n200 & ~n279;
  assign n1284 = ~n377 & n1283;
  assign n1285 = n637 & n832;
  assign n1286 = n840 & n1008;
  assign n1287 = n1285 & n1286;
  assign n1288 = n432 & n1284;
  assign n1289 = n1282 & n1288;
  assign n1290 = n1287 & n1289;
  assign n1291 = ~n180 & ~n189;
  assign n1292 = ~n196 & ~n311;
  assign n1293 = ~n317 & ~n436;
  assign n1294 = ~n520 & ~n546;
  assign n1295 = ~n780 & n1294;
  assign n1296 = n1292 & n1293;
  assign n1297 = n1291 & n1296;
  assign n1298 = n1295 & n1297;
  assign n1299 = ~n341 & ~n560;
  assign n1300 = ~n356 & ~n461;
  assign n1301 = ~n142 & ~n190;
  assign n1302 = ~n274 & ~n384;
  assign n1303 = n1301 & n1302;
  assign n1304 = n344 & n757;
  assign n1305 = n782 & n1304;
  assign n1306 = n1303 & n1305;
  assign n1307 = ~n131 & ~n284;
  assign n1308 = ~n623 & n1307;
  assign n1309 = n615 & n1299;
  assign n1310 = n1300 & n1309;
  assign n1311 = n1308 & n1310;
  assign n1312 = n488 & n1311;
  assign n1313 = n1298 & n1306;
  assign n1314 = n1312 & n1313;
  assign n1315 = n1290 & n1314;
  assign n1316 = ~n989 & ~n1315;
  assign n1317 = n604 & ~n989;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = n1281 & ~n1318;
  assign n1320 = ~n1281 & n1318;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = n594 & ~n1209;
  assign n1323 = ~n594 & n1207;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = ~n663 & n1213;
  assign n1326 = n663 & n1211;
  assign n1327 = ~n1325 & ~n1326;
  assign n1328 = ~n1324 & n1327;
  assign n1329 = n1321 & n1328;
  assign n1330 = ~n1319 & ~n1329;
  assign n1331 = n57 & n585;
  assign n1332 = ~n57 & n588;
  assign n1333 = n504 & n1045;
  assign n1334 = ~n1046 & ~n1333;
  assign n1335 = n583 & ~n1334;
  assign n1336 = ~n1331 & ~n1335;
  assign n1337 = ~n1332 & n1336;
  assign n1338 = ~n1330 & n1337;
  assign n1339 = n1330 & ~n1337;
  assign n1340 = ~n1338 & ~n1339;
  assign n1341 = n453 & n879;
  assign n1342 = ~n453 & n881;
  assign n1343 = n679 & ~n867;
  assign n1344 = n867 & n883;
  assign n1345 = ~n1341 & ~n1342;
  assign n1346 = ~n1343 & ~n1344;
  assign n1347 = n1345 & n1346;
  assign n1348 = n511 & ~n1106;
  assign n1349 = ~n511 & ~n1108;
  assign n1350 = ~n1348 & ~n1349;
  assign n1351 = ~n519 & n1113;
  assign n1352 = n519 & n1111;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = ~n1350 & n1353;
  assign n1355 = n1347 & n1354;
  assign n1356 = ~n1347 & ~n1354;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = n657 & n747;
  assign n1359 = n659 & ~n747;
  assign n1360 = n668 & ~n1045;
  assign n1361 = n665 & n1045;
  assign n1362 = ~n1358 & ~n1359;
  assign n1363 = ~n1360 & ~n1361;
  assign n1364 = n1362 & n1363;
  assign n1365 = n1357 & n1364;
  assign n1366 = ~n1355 & ~n1365;
  assign n1367 = n1340 & ~n1366;
  assign n1368 = ~n1338 & ~n1367;
  assign n1369 = ~n1273 & ~n1275;
  assign n1370 = ~n1276 & ~n1369;
  assign n1371 = ~n1368 & n1370;
  assign n1372 = ~n1276 & ~n1371;
  assign n1373 = n1164 & ~n1166;
  assign n1374 = ~n1167 & ~n1373;
  assign n1375 = ~n1372 & n1374;
  assign n1376 = n1372 & ~n1374;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = n1257 & ~n1259;
  assign n1379 = ~n1260 & ~n1378;
  assign n1380 = n1377 & n1379;
  assign n1381 = ~n1375 & ~n1380;
  assign n1382 = ~n1264 & ~n1266;
  assign n1383 = ~n1267 & ~n1382;
  assign n1384 = ~n1381 & n1383;
  assign n1385 = n583 & n1280;
  assign n1386 = n587 & ~n1385;
  assign n1387 = ~n604 & n1316;
  assign n1388 = ~n604 & ~n1315;
  assign n1389 = n989 & ~n1388;
  assign n1390 = n663 & n1315;
  assign n1391 = ~n1387 & ~n1390;
  assign n1392 = ~n1389 & n1391;
  assign n1393 = n1386 & n1392;
  assign n1394 = n585 & ~n1201;
  assign n1395 = n588 & n1201;
  assign n1396 = ~n57 & n504;
  assign n1397 = ~n1152 & ~n1396;
  assign n1398 = n583 & ~n1397;
  assign n1399 = ~n1394 & ~n1398;
  assign n1400 = ~n1395 & n1399;
  assign n1401 = n1393 & n1400;
  assign n1402 = ~n867 & n879;
  assign n1403 = n867 & n881;
  assign n1404 = ~n747 & n883;
  assign n1405 = n679 & n747;
  assign n1406 = ~n1402 & ~n1403;
  assign n1407 = ~n1404 & ~n1405;
  assign n1408 = n1406 & n1407;
  assign n1409 = n657 & ~n1045;
  assign n1410 = n659 & n1045;
  assign n1411 = ~n57 & n665;
  assign n1412 = n57 & n668;
  assign n1413 = ~n1409 & ~n1410;
  assign n1414 = ~n1411 & ~n1412;
  assign n1415 = n1413 & n1414;
  assign n1416 = n1408 & n1415;
  assign n1417 = ~n1408 & ~n1415;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = ~n453 & ~n1106;
  assign n1420 = n453 & ~n1108;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = ~n511 & n1111;
  assign n1423 = n511 & n1113;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = ~n1421 & n1424;
  assign n1426 = n1418 & n1425;
  assign n1427 = ~n1416 & ~n1426;
  assign n1428 = ~n1393 & ~n1400;
  assign n1429 = ~n1401 & ~n1428;
  assign n1430 = ~n1427 & n1429;
  assign n1431 = ~n1401 & ~n1430;
  assign n1432 = ~n1205 & ~n1217;
  assign n1433 = ~n1218 & ~n1432;
  assign n1434 = ~n1431 & n1433;
  assign n1435 = n1431 & ~n1433;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = ~n1246 & ~n1253;
  assign n1438 = ~n1254 & ~n1437;
  assign n1439 = n1436 & n1438;
  assign n1440 = ~n1434 & ~n1439;
  assign n1441 = ~n1229 & n1255;
  assign n1442 = ~n1256 & ~n1441;
  assign n1443 = ~n1440 & n1442;
  assign n1444 = n1440 & ~n1442;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = n1368 & ~n1370;
  assign n1447 = ~n1371 & ~n1446;
  assign n1448 = n1445 & n1447;
  assign n1449 = ~n1443 & ~n1448;
  assign n1450 = ~n1377 & ~n1379;
  assign n1451 = ~n1380 & ~n1450;
  assign n1452 = ~n1449 & n1451;
  assign n1453 = n585 & n1280;
  assign n1454 = n588 & ~n1280;
  assign n1455 = n504 & n1201;
  assign n1456 = ~n1202 & ~n1455;
  assign n1457 = n583 & ~n1456;
  assign n1458 = ~n1453 & ~n1457;
  assign n1459 = ~n1454 & n1458;
  assign n1460 = n519 & ~n1207;
  assign n1461 = ~n519 & n1209;
  assign n1462 = ~n594 & n1211;
  assign n1463 = n594 & n1213;
  assign n1464 = ~n1460 & ~n1461;
  assign n1465 = ~n1462 & ~n1463;
  assign n1466 = n1464 & n1465;
  assign n1467 = n1459 & n1466;
  assign n1468 = ~n1386 & ~n1392;
  assign n1469 = ~n1393 & ~n1468;
  assign n1470 = ~n1459 & ~n1466;
  assign n1471 = ~n1467 & ~n1470;
  assign n1472 = n1469 & n1471;
  assign n1473 = ~n1467 & ~n1472;
  assign n1474 = ~n1321 & ~n1328;
  assign n1475 = ~n1329 & ~n1474;
  assign n1476 = ~n1473 & n1475;
  assign n1477 = n1473 & ~n1475;
  assign n1478 = ~n1476 & ~n1477;
  assign n1479 = ~n1357 & ~n1364;
  assign n1480 = ~n1365 & ~n1479;
  assign n1481 = n1478 & n1480;
  assign n1482 = ~n1476 & ~n1481;
  assign n1483 = ~n1340 & n1366;
  assign n1484 = ~n1367 & ~n1483;
  assign n1485 = ~n1482 & n1484;
  assign n1486 = n1482 & ~n1484;
  assign n1487 = ~n1485 & ~n1486;
  assign n1488 = ~n1436 & ~n1438;
  assign n1489 = ~n1439 & ~n1488;
  assign n1490 = n1487 & n1489;
  assign n1491 = ~n1485 & ~n1490;
  assign n1492 = ~n1445 & ~n1447;
  assign n1493 = ~n1448 & ~n1492;
  assign n1494 = ~n1491 & n1493;
  assign n1495 = n867 & ~n1106;
  assign n1496 = ~n867 & ~n1108;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = ~n453 & n1113;
  assign n1499 = n453 & n1111;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = ~n1497 & n1500;
  assign n1502 = n747 & n879;
  assign n1503 = ~n747 & n881;
  assign n1504 = n679 & ~n1045;
  assign n1505 = n883 & n1045;
  assign n1506 = ~n1502 & ~n1503;
  assign n1507 = ~n1504 & ~n1505;
  assign n1508 = n1506 & n1507;
  assign n1509 = n1501 & n1508;
  assign n1510 = n656 & n1280;
  assign n1511 = n664 & ~n1510;
  assign n1512 = ~n594 & n1316;
  assign n1513 = ~n594 & ~n1315;
  assign n1514 = n989 & ~n1513;
  assign n1515 = n519 & n1315;
  assign n1516 = ~n1512 & ~n1515;
  assign n1517 = ~n1514 & n1516;
  assign n1518 = n1511 & n1517;
  assign n1519 = ~n1501 & ~n1508;
  assign n1520 = ~n1509 & ~n1519;
  assign n1521 = n1518 & n1520;
  assign n1522 = ~n1509 & ~n1521;
  assign n1523 = n663 & n1316;
  assign n1524 = n663 & ~n1315;
  assign n1525 = n989 & ~n1524;
  assign n1526 = ~n594 & n1315;
  assign n1527 = ~n1523 & ~n1526;
  assign n1528 = ~n1525 & n1527;
  assign n1529 = n511 & ~n1209;
  assign n1530 = ~n511 & n1207;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = ~n519 & n1213;
  assign n1533 = n519 & n1211;
  assign n1534 = ~n1532 & ~n1533;
  assign n1535 = ~n1531 & n1534;
  assign n1536 = n1528 & n1535;
  assign n1537 = ~n1528 & ~n1535;
  assign n1538 = ~n1536 & ~n1537;
  assign n1539 = n57 & n657;
  assign n1540 = ~n57 & n659;
  assign n1541 = n668 & ~n1201;
  assign n1542 = n665 & n1201;
  assign n1543 = ~n1539 & ~n1540;
  assign n1544 = ~n1541 & ~n1542;
  assign n1545 = n1543 & n1544;
  assign n1546 = n1538 & n1545;
  assign n1547 = ~n1536 & ~n1546;
  assign n1548 = ~n1522 & ~n1547;
  assign n1549 = n1522 & n1547;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = ~n1418 & ~n1425;
  assign n1552 = ~n1426 & ~n1551;
  assign n1553 = n1550 & n1552;
  assign n1554 = ~n1548 & ~n1553;
  assign n1555 = n1427 & ~n1429;
  assign n1556 = ~n1430 & ~n1555;
  assign n1557 = ~n1554 & n1556;
  assign n1558 = n1554 & ~n1556;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = ~n1478 & ~n1480;
  assign n1561 = ~n1481 & ~n1560;
  assign n1562 = n1559 & n1561;
  assign n1563 = ~n1557 & ~n1562;
  assign n1564 = ~n1487 & ~n1489;
  assign n1565 = ~n1490 & ~n1564;
  assign n1566 = ~n1563 & n1565;
  assign n1567 = n453 & ~n1207;
  assign n1568 = ~n453 & n1209;
  assign n1569 = ~n511 & n1211;
  assign n1570 = n511 & n1213;
  assign n1571 = ~n1567 & ~n1568;
  assign n1572 = ~n1569 & ~n1570;
  assign n1573 = n1571 & n1572;
  assign n1574 = n879 & ~n1045;
  assign n1575 = n881 & n1045;
  assign n1576 = ~n57 & n883;
  assign n1577 = n57 & n679;
  assign n1578 = ~n1574 & ~n1575;
  assign n1579 = ~n1576 & ~n1577;
  assign n1580 = n1578 & n1579;
  assign n1581 = n1573 & n1580;
  assign n1582 = ~n1573 & ~n1580;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = ~n747 & ~n1106;
  assign n1585 = n747 & ~n1108;
  assign n1586 = ~n1584 & ~n1585;
  assign n1587 = ~n867 & n1111;
  assign n1588 = n867 & n1113;
  assign n1589 = ~n1587 & ~n1588;
  assign n1590 = ~n1586 & n1589;
  assign n1591 = n1583 & n1590;
  assign n1592 = ~n1581 & ~n1591;
  assign n1593 = n1385 & ~n1592;
  assign n1594 = ~n1518 & ~n1520;
  assign n1595 = ~n1521 & ~n1594;
  assign n1596 = ~n1385 & n1592;
  assign n1597 = ~n1593 & ~n1596;
  assign n1598 = n1595 & n1597;
  assign n1599 = ~n1593 & ~n1598;
  assign n1600 = n1469 & ~n1471;
  assign n1601 = ~n1469 & n1471;
  assign n1602 = ~n1600 & ~n1601;
  assign n1603 = ~n1599 & ~n1602;
  assign n1604 = n1599 & n1602;
  assign n1605 = ~n1603 & ~n1604;
  assign n1606 = ~n1550 & ~n1552;
  assign n1607 = ~n1553 & ~n1606;
  assign n1608 = n1605 & n1607;
  assign n1609 = ~n1603 & ~n1608;
  assign n1610 = ~n1559 & ~n1561;
  assign n1611 = ~n1562 & ~n1610;
  assign n1612 = ~n1609 & n1611;
  assign n1613 = n1609 & ~n1611;
  assign n1614 = ~n1612 & ~n1613;
  assign n1615 = ~n1511 & ~n1517;
  assign n1616 = ~n1518 & ~n1615;
  assign n1617 = n657 & ~n1201;
  assign n1618 = n659 & n1201;
  assign n1619 = n665 & ~n1280;
  assign n1620 = n668 & n1280;
  assign n1621 = ~n1617 & ~n1618;
  assign n1622 = ~n1619 & ~n1620;
  assign n1623 = n1621 & n1622;
  assign n1624 = n1616 & n1623;
  assign n1625 = n519 & n1316;
  assign n1626 = n519 & ~n1315;
  assign n1627 = n989 & ~n1626;
  assign n1628 = ~n511 & n1315;
  assign n1629 = ~n1625 & ~n1628;
  assign n1630 = ~n1627 & n1629;
  assign n1631 = n867 & ~n1209;
  assign n1632 = ~n867 & n1207;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = ~n453 & n1213;
  assign n1635 = n453 & n1211;
  assign n1636 = ~n1634 & ~n1635;
  assign n1637 = ~n1633 & n1636;
  assign n1638 = n1630 & n1637;
  assign n1639 = ~n1630 & ~n1637;
  assign n1640 = ~n1638 & ~n1639;
  assign n1641 = n1045 & ~n1106;
  assign n1642 = ~n1045 & ~n1108;
  assign n1643 = ~n1641 & ~n1642;
  assign n1644 = ~n747 & n1113;
  assign n1645 = n747 & n1111;
  assign n1646 = ~n1644 & ~n1645;
  assign n1647 = ~n1643 & n1646;
  assign n1648 = n1640 & n1647;
  assign n1649 = ~n1638 & ~n1648;
  assign n1650 = ~n1616 & ~n1623;
  assign n1651 = ~n1624 & ~n1650;
  assign n1652 = ~n1649 & n1651;
  assign n1653 = ~n1624 & ~n1652;
  assign n1654 = ~n1538 & ~n1545;
  assign n1655 = ~n1546 & ~n1654;
  assign n1656 = ~n1653 & n1655;
  assign n1657 = ~n1595 & ~n1597;
  assign n1658 = ~n1598 & ~n1657;
  assign n1659 = n1653 & ~n1655;
  assign n1660 = ~n1656 & ~n1659;
  assign n1661 = n1658 & n1660;
  assign n1662 = ~n1656 & ~n1661;
  assign n1663 = n675 & n1280;
  assign n1664 = n449 & ~n1663;
  assign n1665 = ~n511 & n1316;
  assign n1666 = ~n511 & ~n1315;
  assign n1667 = n989 & ~n1666;
  assign n1668 = n453 & n1315;
  assign n1669 = ~n1665 & ~n1668;
  assign n1670 = ~n1667 & n1669;
  assign n1671 = n1664 & n1670;
  assign n1672 = n57 & n879;
  assign n1673 = ~n57 & n881;
  assign n1674 = n679 & ~n1201;
  assign n1675 = n883 & n1201;
  assign n1676 = ~n1672 & ~n1673;
  assign n1677 = ~n1674 & ~n1675;
  assign n1678 = n1676 & n1677;
  assign n1679 = n1671 & n1678;
  assign n1680 = ~n1671 & ~n1678;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = n1510 & n1681;
  assign n1683 = ~n1679 & ~n1682;
  assign n1684 = ~n1583 & ~n1590;
  assign n1685 = ~n1591 & ~n1684;
  assign n1686 = ~n1683 & n1685;
  assign n1687 = n1683 & ~n1685;
  assign n1688 = ~n1686 & ~n1687;
  assign n1689 = n1649 & ~n1651;
  assign n1690 = ~n1652 & ~n1689;
  assign n1691 = n1688 & n1690;
  assign n1692 = ~n1686 & ~n1691;
  assign n1693 = n747 & ~n1207;
  assign n1694 = ~n747 & n1209;
  assign n1695 = ~n867 & n1211;
  assign n1696 = n867 & n1213;
  assign n1697 = ~n1693 & ~n1694;
  assign n1698 = ~n1695 & ~n1696;
  assign n1699 = n1697 & n1698;
  assign n1700 = ~n57 & ~n1106;
  assign n1701 = n57 & ~n1108;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n1045 & n1111;
  assign n1704 = n1045 & n1113;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = ~n1702 & n1705;
  assign n1707 = n1699 & n1706;
  assign n1708 = ~n1699 & ~n1706;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = n879 & ~n1201;
  assign n1711 = n881 & n1201;
  assign n1712 = n883 & ~n1280;
  assign n1713 = n679 & n1280;
  assign n1714 = ~n1710 & ~n1711;
  assign n1715 = ~n1712 & ~n1713;
  assign n1716 = n1714 & n1715;
  assign n1717 = n1709 & n1716;
  assign n1718 = ~n1707 & ~n1717;
  assign n1719 = ~n1640 & ~n1647;
  assign n1720 = ~n1648 & ~n1719;
  assign n1721 = ~n1718 & n1720;
  assign n1722 = ~n1510 & ~n1681;
  assign n1723 = ~n1682 & ~n1722;
  assign n1724 = n1718 & ~n1720;
  assign n1725 = ~n1721 & ~n1724;
  assign n1726 = n1723 & n1725;
  assign n1727 = ~n1721 & ~n1726;
  assign n1728 = ~n1664 & ~n1670;
  assign n1729 = ~n1671 & ~n1728;
  assign n1730 = n453 & n1316;
  assign n1731 = n453 & ~n1315;
  assign n1732 = n989 & ~n1731;
  assign n1733 = ~n867 & n1315;
  assign n1734 = ~n1730 & ~n1733;
  assign n1735 = ~n1732 & n1734;
  assign n1736 = n1045 & ~n1209;
  assign n1737 = ~n1045 & n1207;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = ~n747 & n1213;
  assign n1740 = n747 & n1211;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = ~n1738 & n1741;
  assign n1743 = n1735 & n1742;
  assign n1744 = ~n1735 & ~n1742;
  assign n1745 = ~n1743 & ~n1744;
  assign n1746 = ~n1106 & n1201;
  assign n1747 = ~n1108 & ~n1201;
  assign n1748 = ~n1746 & ~n1747;
  assign n1749 = ~n57 & n1113;
  assign n1750 = n57 & n1111;
  assign n1751 = ~n1749 & ~n1750;
  assign n1752 = ~n1748 & n1751;
  assign n1753 = n1745 & n1752;
  assign n1754 = ~n1743 & ~n1753;
  assign n1755 = n1729 & ~n1754;
  assign n1756 = ~n1729 & n1754;
  assign n1757 = ~n1755 & ~n1756;
  assign n1758 = ~n1709 & ~n1716;
  assign n1759 = ~n1717 & ~n1758;
  assign n1760 = n1757 & n1759;
  assign n1761 = ~n1755 & ~n1760;
  assign n1762 = n1052 & n1280;
  assign n1763 = n860 & ~n1762;
  assign n1764 = ~n867 & n1316;
  assign n1765 = ~n867 & ~n1315;
  assign n1766 = n989 & ~n1765;
  assign n1767 = n747 & n1315;
  assign n1768 = ~n1764 & ~n1767;
  assign n1769 = ~n1766 & n1768;
  assign n1770 = n1763 & n1769;
  assign n1771 = n1663 & n1770;
  assign n1772 = n57 & ~n1207;
  assign n1773 = ~n57 & n1209;
  assign n1774 = ~n1045 & n1211;
  assign n1775 = n1045 & n1213;
  assign n1776 = ~n1772 & ~n1773;
  assign n1777 = ~n1774 & ~n1775;
  assign n1778 = n1776 & n1777;
  assign n1779 = ~n1108 & n1280;
  assign n1780 = ~n1106 & ~n1280;
  assign n1781 = ~n1779 & ~n1780;
  assign n1782 = n1113 & n1201;
  assign n1783 = n1111 & ~n1201;
  assign n1784 = ~n1782 & ~n1783;
  assign n1785 = ~n1781 & n1784;
  assign n1786 = n1778 & n1785;
  assign n1787 = ~n1763 & ~n1769;
  assign n1788 = ~n1770 & ~n1787;
  assign n1789 = ~n1778 & ~n1785;
  assign n1790 = ~n1786 & ~n1789;
  assign n1791 = n1788 & n1790;
  assign n1792 = ~n1786 & ~n1791;
  assign n1793 = ~n1663 & ~n1770;
  assign n1794 = ~n1771 & ~n1793;
  assign n1795 = ~n1792 & n1794;
  assign n1796 = ~n1771 & ~n1795;
  assign n1797 = n1792 & ~n1794;
  assign n1798 = ~n1795 & ~n1797;
  assign n1799 = n747 & n1316;
  assign n1800 = n747 & ~n1315;
  assign n1801 = n989 & ~n1800;
  assign n1802 = ~n1045 & n1315;
  assign n1803 = ~n1799 & ~n1802;
  assign n1804 = ~n1801 & n1803;
  assign n1805 = n1201 & ~n1209;
  assign n1806 = ~n1201 & n1207;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = n57 & n1211;
  assign n1809 = ~n57 & n1213;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = ~n1807 & n1810;
  assign n1812 = n1804 & n1811;
  assign n1813 = n1157 & n1280;
  assign n1814 = n1040 & ~n1813;
  assign n1815 = ~n1045 & n1316;
  assign n1816 = ~n1045 & ~n1315;
  assign n1817 = n989 & ~n1816;
  assign n1818 = n57 & n1315;
  assign n1819 = ~n1815 & ~n1818;
  assign n1820 = ~n1817 & n1819;
  assign n1821 = n1814 & n1820;
  assign n1822 = ~n1804 & ~n1811;
  assign n1823 = ~n1812 & ~n1822;
  assign n1824 = n1821 & n1823;
  assign n1825 = ~n1812 & ~n1824;
  assign n1826 = ~n1788 & ~n1790;
  assign n1827 = ~n1791 & ~n1826;
  assign n1828 = n1825 & ~n1827;
  assign n1829 = ~n1825 & n1827;
  assign n1830 = ~n1814 & ~n1820;
  assign n1831 = ~n1821 & ~n1830;
  assign n1832 = ~n1201 & ~n1315;
  assign n1833 = ~n989 & ~n1280;
  assign n1834 = ~n1832 & n1833;
  assign n1835 = n57 & n1316;
  assign n1836 = n57 & ~n1315;
  assign n1837 = n989 & ~n1836;
  assign n1838 = ~n1201 & n1315;
  assign n1839 = ~n1835 & ~n1838;
  assign n1840 = ~n1837 & n1839;
  assign n1841 = n1813 & n1840;
  assign n1842 = ~n1834 & ~n1841;
  assign n1843 = ~n1813 & ~n1840;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845 = ~n1831 & ~n1844;
  assign n1846 = n1831 & n1844;
  assign n1847 = ~n1209 & ~n1280;
  assign n1848 = n1207 & n1280;
  assign n1849 = ~n1847 & ~n1848;
  assign n1850 = ~n1201 & n1211;
  assign n1851 = n1201 & n1213;
  assign n1852 = ~n1850 & ~n1851;
  assign n1853 = ~n1849 & n1852;
  assign n1854 = ~n1846 & ~n1853;
  assign n1855 = ~n1845 & ~n1854;
  assign n1856 = n1762 & n1855;
  assign n1857 = ~n1762 & ~n1855;
  assign n1858 = ~n1821 & ~n1823;
  assign n1859 = ~n1824 & ~n1858;
  assign n1860 = ~n1857 & n1859;
  assign n1861 = ~n1829 & ~n1856;
  assign n1862 = ~n1860 & n1861;
  assign n1863 = ~n1828 & ~n1862;
  assign n1864 = ~n1798 & ~n1863;
  assign n1865 = n1798 & n1863;
  assign n1866 = ~n1745 & ~n1752;
  assign n1867 = ~n1753 & ~n1866;
  assign n1868 = ~n1865 & ~n1867;
  assign n1869 = ~n1864 & ~n1868;
  assign n1870 = n1796 & ~n1869;
  assign n1871 = ~n1796 & n1869;
  assign n1872 = ~n1757 & ~n1759;
  assign n1873 = ~n1760 & ~n1872;
  assign n1874 = ~n1871 & ~n1873;
  assign n1875 = ~n1870 & ~n1874;
  assign n1876 = n1761 & ~n1875;
  assign n1877 = ~n1761 & n1875;
  assign n1878 = ~n1723 & ~n1725;
  assign n1879 = ~n1726 & ~n1878;
  assign n1880 = ~n1877 & ~n1879;
  assign n1881 = ~n1876 & ~n1880;
  assign n1882 = n1727 & ~n1881;
  assign n1883 = ~n1727 & n1881;
  assign n1884 = ~n1688 & ~n1690;
  assign n1885 = ~n1691 & ~n1884;
  assign n1886 = ~n1883 & ~n1885;
  assign n1887 = ~n1882 & ~n1886;
  assign n1888 = n1692 & ~n1887;
  assign n1889 = ~n1692 & n1887;
  assign n1890 = ~n1658 & ~n1660;
  assign n1891 = ~n1661 & ~n1890;
  assign n1892 = ~n1889 & ~n1891;
  assign n1893 = ~n1888 & ~n1892;
  assign n1894 = n1662 & ~n1893;
  assign n1895 = ~n1662 & n1893;
  assign n1896 = ~n1605 & ~n1607;
  assign n1897 = ~n1608 & ~n1896;
  assign n1898 = ~n1895 & ~n1897;
  assign n1899 = ~n1894 & ~n1898;
  assign n1900 = n1614 & n1899;
  assign n1901 = ~n1612 & ~n1900;
  assign n1902 = n1563 & ~n1565;
  assign n1903 = ~n1566 & ~n1902;
  assign n1904 = ~n1901 & n1903;
  assign n1905 = ~n1566 & ~n1904;
  assign n1906 = n1491 & ~n1493;
  assign n1907 = ~n1494 & ~n1906;
  assign n1908 = ~n1905 & n1907;
  assign n1909 = ~n1494 & ~n1908;
  assign n1910 = n1449 & ~n1451;
  assign n1911 = ~n1452 & ~n1910;
  assign n1912 = ~n1909 & n1911;
  assign n1913 = ~n1452 & ~n1912;
  assign n1914 = n1381 & ~n1383;
  assign n1915 = ~n1384 & ~n1914;
  assign n1916 = ~n1913 & n1915;
  assign n1917 = ~n1384 & ~n1916;
  assign n1918 = n1268 & ~n1270;
  assign n1919 = ~n1271 & ~n1918;
  assign n1920 = ~n1917 & n1919;
  assign n1921 = ~n1271 & ~n1920;
  assign n1922 = n1136 & ~n1138;
  assign n1923 = ~n1139 & ~n1922;
  assign n1924 = ~n1921 & n1923;
  assign n1925 = ~n1139 & ~n1924;
  assign n1926 = n1085 & ~n1087;
  assign n1927 = ~n1088 & ~n1926;
  assign n1928 = ~n1925 & n1927;
  assign n1929 = ~n1088 & ~n1928;
  assign n1930 = n920 & ~n922;
  assign n1931 = ~n923 & ~n1930;
  assign n1932 = ~n1929 & n1931;
  assign n1933 = ~n923 & ~n1932;
  assign n1934 = n721 & ~n742;
  assign n1935 = ~n743 & ~n1934;
  assign n1936 = ~n1933 & n1935;
  assign n1937 = ~n743 & ~n1936;
  assign n1938 = ~n731 & ~n740;
  assign n1939 = ~n734 & ~n737;
  assign n1940 = n582 & n726;
  assign n1941 = ~n587 & ~n1940;
  assign n1942 = n581 & ~n604;
  assign n1943 = ~n1941 & ~n1942;
  assign n1944 = ~n709 & n1943;
  assign n1945 = n709 & ~n1943;
  assign n1946 = ~n1944 & ~n1945;
  assign n1947 = ~n1939 & n1946;
  assign n1948 = n1939 & ~n1946;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = ~n1938 & n1949;
  assign n1951 = n1938 & ~n1949;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = ~n1937 & n1952;
  assign n1954 = n1937 & ~n1952;
  assign n1955 = ~n1953 & ~n1954;
  assign n1956 = ~n309 & ~n343;
  assign n1957 = ~n370 & ~n412;
  assign n1958 = n1956 & n1957;
  assign n1959 = n786 & n1958;
  assign n1960 = n277 & n1959;
  assign n1961 = ~n140 & ~n560;
  assign n1962 = n840 & n1961;
  assign n1963 = ~n210 & ~n218;
  assign n1964 = ~n311 & n1963;
  assign n1965 = n626 & n1964;
  assign n1966 = n146 & ~n317;
  assign n1967 = n379 & n1966;
  assign n1968 = n184 & n819;
  assign n1969 = n945 & n1962;
  assign n1970 = n1968 & n1969;
  assign n1971 = n1965 & n1967;
  assign n1972 = n1970 & n1971;
  assign n1973 = ~n176 & ~n294;
  assign n1974 = ~n310 & ~n318;
  assign n1975 = ~n520 & n1974;
  assign n1976 = n1973 & n1975;
  assign n1977 = ~n152 & ~n188;
  assign n1978 = ~n192 & ~n209;
  assign n1979 = ~n299 & ~n342;
  assign n1980 = ~n775 & n1979;
  assign n1981 = n1977 & n1978;
  assign n1982 = n114 & n1981;
  assign n1983 = n1980 & n1982;
  assign n1984 = n1976 & n1983;
  assign n1985 = ~n222 & ~n282;
  assign n1986 = ~n554 & n1985;
  assign n1987 = ~n149 & ~n207;
  assign n1988 = ~n262 & ~n377;
  assign n1989 = n1987 & n1988;
  assign n1990 = n135 & n305;
  assign n1991 = n408 & n459;
  assign n1992 = n1990 & n1991;
  assign n1993 = n1986 & n1989;
  assign n1994 = n1992 & n1993;
  assign n1995 = n245 & n1994;
  assign n1996 = n1960 & n1995;
  assign n1997 = n1972 & n1984;
  assign n1998 = n1996 & n1997;
  assign n1999 = ~n1955 & ~n1998;
  assign n2000 = n1933 & ~n1935;
  assign n2001 = ~n1936 & ~n2000;
  assign n2002 = ~n210 & ~n238;
  assign n2003 = ~n248 & ~n294;
  assign n2004 = ~n343 & n2003;
  assign n2005 = n312 & n2002;
  assign n2006 = n414 & n639;
  assign n2007 = n2005 & n2006;
  assign n2008 = n195 & n2004;
  assign n2009 = n270 & n759;
  assign n2010 = n2008 & n2009;
  assign n2011 = n2007 & n2010;
  assign n2012 = n621 & n838;
  assign n2013 = n2011 & n2012;
  assign n2014 = n955 & n2013;
  assign n2015 = ~n2001 & ~n2014;
  assign n2016 = n1929 & ~n1931;
  assign n2017 = ~n1932 & ~n2016;
  assign n2018 = ~n185 & ~n267;
  assign n2019 = ~n157 & ~n176;
  assign n2020 = ~n241 & n2019;
  assign n2021 = n749 & n2018;
  assign n2022 = n2020 & n2021;
  assign n2023 = ~n190 & ~n314;
  assign n2024 = ~n188 & ~n279;
  assign n2025 = n2023 & n2024;
  assign n2026 = n628 & n2025;
  assign n2027 = n407 & n2026;
  assign n2028 = n2022 & n2027;
  assign n2029 = ~n171 & ~n454;
  assign n2030 = ~n197 & ~n372;
  assign n2031 = ~n262 & ~n318;
  assign n2032 = ~n481 & n2031;
  assign n2033 = ~n209 & ~n306;
  assign n2034 = n347 & n2033;
  assign n2035 = n639 & n2029;
  assign n2036 = n2030 & n2035;
  assign n2037 = n1962 & n2034;
  assign n2038 = n1986 & n2032;
  assign n2039 = n2037 & n2038;
  assign n2040 = n402 & n2036;
  assign n2041 = n2039 & n2040;
  assign n2042 = ~n198 & ~n236;
  assign n2043 = ~n284 & n2042;
  assign n2044 = ~n127 & ~n233;
  assign n2045 = ~n251 & n2044;
  assign n2046 = ~n378 & n409;
  assign n2047 = n521 & n637;
  assign n2048 = n956 & n2047;
  assign n2049 = n2043 & n2046;
  assign n2050 = n2045 & n2049;
  assign n2051 = n440 & n2048;
  assign n2052 = n2050 & n2051;
  assign n2053 = n2028 & n2052;
  assign n2054 = n2041 & n2053;
  assign n2055 = ~n2017 & ~n2054;
  assign n2056 = n1925 & ~n1927;
  assign n2057 = ~n1928 & ~n2056;
  assign n2058 = ~n208 & ~n224;
  assign n2059 = ~n377 & ~n571;
  assign n2060 = ~n623 & n2059;
  assign n2061 = n308 & n2058;
  assign n2062 = n456 & n2061;
  assign n2063 = n534 & n2060;
  assign n2064 = n2043 & n2063;
  assign n2065 = n2062 & n2064;
  assign n2066 = ~n142 & ~n241;
  assign n2067 = ~n248 & n2066;
  assign n2068 = ~n134 & ~n297;
  assign n2069 = ~n327 & n2068;
  assign n2070 = n2041 & n2069;
  assign n2071 = ~n192 & ~n427;
  assign n2072 = ~n233 & ~n268;
  assign n2073 = n2071 & n2072;
  assign n2074 = n781 & n813;
  assign n2075 = n2073 & n2074;
  assign n2076 = n1282 & n2067;
  assign n2077 = n2075 & n2076;
  assign n2078 = n1960 & n2077;
  assign n2079 = n2065 & n2078;
  assign n2080 = n2070 & n2079;
  assign n2081 = ~n2057 & ~n2080;
  assign n2082 = n1921 & ~n1923;
  assign n2083 = ~n1924 & ~n2082;
  assign n2084 = ~n200 & ~n241;
  assign n2085 = ~n223 & ~n263;
  assign n2086 = ~n274 & ~n343;
  assign n2087 = n413 & n2086;
  assign n2088 = n637 & n957;
  assign n2089 = n2084 & n2085;
  assign n2090 = n2088 & n2089;
  assign n2091 = n2087 & n2090;
  assign n2092 = n802 & n2091;
  assign n2093 = ~n186 & ~n310;
  assign n2094 = n774 & n2093;
  assign n2095 = ~n189 & ~n372;
  assign n2096 = ~n147 & ~n180;
  assign n2097 = ~n238 & ~n309;
  assign n2098 = n2096 & n2097;
  assign n2099 = n2023 & n2095;
  assign n2100 = n2098 & n2099;
  assign n2101 = ~n131 & ~n149;
  assign n2102 = ~n182 & ~n345;
  assign n2103 = ~n405 & n2102;
  assign n2104 = n2101 & n2103;
  assign n2105 = ~n127 & ~n145;
  assign n2106 = ~n222 & ~n247;
  assign n2107 = ~n262 & ~n325;
  assign n2108 = n2106 & n2107;
  assign n2109 = n533 & n2105;
  assign n2110 = n2108 & n2109;
  assign n2111 = n2100 & n2110;
  assign n2112 = n2104 & n2111;
  assign n2113 = n2092 & n2112;
  assign n2114 = n2094 & n2113;
  assign n2115 = ~n2083 & ~n2114;
  assign n2116 = n1917 & ~n1919;
  assign n2117 = ~n1920 & ~n2116;
  assign n2118 = ~n188 & ~n220;
  assign n2119 = ~n542 & n2118;
  assign n2120 = n562 & n2119;
  assign n2121 = ~n147 & ~n345;
  assign n2122 = ~n158 & n187;
  assign n2123 = ~n310 & ~n405;
  assign n2124 = ~n271 & ~n403;
  assign n2125 = n765 & n2124;
  assign n2126 = n785 & n2123;
  assign n2127 = n2125 & n2126;
  assign n2128 = n136 & n2127;
  assign n2129 = ~n182 & ~n201;
  assign n2130 = ~n356 & n2129;
  assign n2131 = n455 & n622;
  assign n2132 = n974 & n2121;
  assign n2133 = n2131 & n2132;
  assign n2134 = n328 & n2130;
  assign n2135 = n2122 & n2134;
  assign n2136 = n790 & n2133;
  assign n2137 = n2120 & n2136;
  assign n2138 = n2128 & n2135;
  assign n2139 = n2137 & n2138;
  assign n2140 = n827 & n2139;
  assign n2141 = ~n2117 & ~n2140;
  assign n2142 = n1913 & ~n1915;
  assign n2143 = ~n1916 & ~n2142;
  assign n2144 = ~n378 & ~n429;
  assign n2145 = ~n481 & n2144;
  assign n2146 = ~n248 & ~n325;
  assign n2147 = ~n119 & ~n181;
  assign n2148 = ~n196 & ~n458;
  assign n2149 = n2147 & n2148;
  assign n2150 = n319 & n2146;
  assign n2151 = n2149 & n2150;
  assign n2152 = n2145 & n2151;
  assign n2153 = n753 & n2152;
  assign n2154 = ~n264 & ~n377;
  assign n2155 = n2085 & n2154;
  assign n2156 = ~n272 & ~n280;
  assign n2157 = ~n345 & ~n384;
  assign n2158 = n2156 & n2157;
  assign n2159 = n615 & n2158;
  assign n2160 = n2155 & n2159;
  assign n2161 = n402 & n1029;
  assign n2162 = n2160 & n2161;
  assign n2163 = ~n155 & n409;
  assign n2164 = n2162 & n2163;
  assign n2165 = ~n197 & ~n279;
  assign n2166 = ~n370 & ~n537;
  assign n2167 = n2165 & n2166;
  assign n2168 = n413 & n760;
  assign n2169 = n2167 & n2168;
  assign n2170 = ~n113 & ~n240;
  assign n2171 = ~n192 & ~n274;
  assign n2172 = ~n306 & ~n355;
  assign n2173 = ~n454 & n2172;
  assign n2174 = n2170 & n2171;
  assign n2175 = n146 & n2174;
  assign n2176 = n2173 & n2175;
  assign n2177 = n2169 & n2176;
  assign n2178 = n2153 & n2177;
  assign n2179 = n2164 & n2178;
  assign n2180 = ~n2143 & ~n2179;
  assign n2181 = n1909 & ~n1911;
  assign n2182 = ~n1912 & ~n2181;
  assign n2183 = ~n149 & ~n299;
  assign n2184 = ~n272 & ~n310;
  assign n2185 = ~n403 & ~n436;
  assign n2186 = n2184 & n2185;
  assign n2187 = n749 & n2186;
  assign n2188 = n376 & n475;
  assign n2189 = n2045 & n2188;
  assign n2190 = n2187 & n2189;
  assign n2191 = ~n145 & ~n377;
  assign n2192 = n482 & n2191;
  assign n2193 = n522 & n973;
  assign n2194 = n2192 & n2193;
  assign n2195 = ~n222 & ~n297;
  assign n2196 = ~n303 & ~n341;
  assign n2197 = ~n372 & ~n378;
  assign n2198 = ~n520 & n2197;
  assign n2199 = n2195 & n2196;
  assign n2200 = n346 & n426;
  assign n2201 = n2183 & n2200;
  assign n2202 = n2198 & n2199;
  assign n2203 = n819 & n2202;
  assign n2204 = n2194 & n2201;
  assign n2205 = n2203 & n2204;
  assign n2206 = n217 & n2205;
  assign n2207 = n2190 & n2206;
  assign n2208 = ~n2182 & ~n2207;
  assign n2209 = n1905 & ~n1907;
  assign n2210 = ~n1908 & ~n2209;
  assign n2211 = ~n199 & ~n207;
  assign n2212 = ~n294 & n615;
  assign n2213 = ~n113 & ~n224;
  assign n2214 = ~n297 & ~n429;
  assign n2215 = ~n370 & ~n623;
  assign n2216 = ~n267 & ~n298;
  assign n2217 = ~n571 & n2216;
  assign n2218 = n2215 & n2217;
  assign n2219 = ~n272 & n839;
  assign n2220 = n2213 & n2214;
  assign n2221 = n2219 & n2220;
  assign n2222 = n784 & n2067;
  assign n2223 = n2212 & n2222;
  assign n2224 = n2120 & n2221;
  assign n2225 = n2218 & n2224;
  assign n2226 = n2223 & n2225;
  assign n2227 = ~n125 & ~n185;
  assign n2228 = ~n249 & ~n262;
  assign n2229 = ~n436 & n2228;
  assign n2230 = n296 & n2227;
  assign n2231 = n456 & n781;
  assign n2232 = n2211 & n2231;
  assign n2233 = n2229 & n2230;
  assign n2234 = n2232 & n2233;
  assign n2235 = n816 & n2194;
  assign n2236 = n2234 & n2235;
  assign n2237 = n764 & n2236;
  assign n2238 = n421 & n2237;
  assign n2239 = n2226 & n2238;
  assign n2240 = ~n2210 & ~n2239;
  assign n2241 = n1901 & ~n1903;
  assign n2242 = ~n1904 & ~n2241;
  assign n2243 = ~n282 & ~n461;
  assign n2244 = ~n303 & ~n412;
  assign n2245 = ~n274 & ~n313;
  assign n2246 = ~n378 & n2245;
  assign n2247 = n2244 & n2246;
  assign n2248 = n121 & ~n499;
  assign n2249 = ~n144 & ~n268;
  assign n2250 = ~n560 & ~n2248;
  assign n2251 = n2249 & n2250;
  assign n2252 = ~n142 & ~n224;
  assign n2253 = ~n317 & ~n343;
  assign n2254 = ~n428 & n2253;
  assign n2255 = n2252 & n2254;
  assign n2256 = n2251 & n2255;
  assign n2257 = n2247 & n2256;
  assign n2258 = ~n127 & ~n190;
  assign n2259 = ~n200 & ~n309;
  assign n2260 = ~n399 & ~n537;
  assign n2261 = n2259 & n2260;
  assign n2262 = n312 & n2258;
  assign n2263 = n605 & n2214;
  assign n2264 = n2243 & n2263;
  assign n2265 = n2261 & n2262;
  assign n2266 = n302 & n2265;
  assign n2267 = n2264 & n2266;
  assign n2268 = n2128 & n2267;
  assign n2269 = n2257 & n2268;
  assign n2270 = ~n2242 & ~n2269;
  assign n2271 = ~n1614 & ~n1899;
  assign n2272 = ~n1900 & ~n2271;
  assign n2273 = ~n399 & ~n775;
  assign n2274 = ~n279 & ~n623;
  assign n2275 = n2273 & n2274;
  assign n2276 = n178 & n2275;
  assign n2277 = n195 & n943;
  assign n2278 = n2212 & n2277;
  assign n2279 = n756 & n2276;
  assign n2280 = n2278 & n2279;
  assign n2281 = n1972 & n2280;
  assign n2282 = n2190 & n2281;
  assign n2283 = n2272 & n2282;
  assign n2284 = n2242 & n2269;
  assign n2285 = ~n2270 & ~n2284;
  assign n2286 = ~n2283 & n2285;
  assign n2287 = ~n2270 & ~n2286;
  assign n2288 = n2210 & n2239;
  assign n2289 = ~n2240 & ~n2288;
  assign n2290 = ~n2287 & n2289;
  assign n2291 = ~n2240 & ~n2290;
  assign n2292 = n2182 & n2207;
  assign n2293 = ~n2208 & ~n2292;
  assign n2294 = ~n2291 & n2293;
  assign n2295 = ~n2208 & ~n2294;
  assign n2296 = n2143 & n2179;
  assign n2297 = ~n2180 & ~n2296;
  assign n2298 = ~n2295 & n2297;
  assign n2299 = ~n2180 & ~n2298;
  assign n2300 = n2117 & n2140;
  assign n2301 = ~n2141 & ~n2300;
  assign n2302 = ~n2299 & n2301;
  assign n2303 = ~n2141 & ~n2302;
  assign n2304 = n2083 & n2114;
  assign n2305 = ~n2115 & ~n2304;
  assign n2306 = ~n2303 & n2305;
  assign n2307 = ~n2115 & ~n2306;
  assign n2308 = n2057 & n2080;
  assign n2309 = ~n2081 & ~n2308;
  assign n2310 = ~n2307 & n2309;
  assign n2311 = ~n2081 & ~n2310;
  assign n2312 = n2017 & n2054;
  assign n2313 = ~n2055 & ~n2312;
  assign n2314 = ~n2311 & n2313;
  assign n2315 = ~n2055 & ~n2314;
  assign n2316 = n2001 & n2014;
  assign n2317 = ~n2015 & ~n2316;
  assign n2318 = ~n2315 & n2317;
  assign n2319 = ~n2015 & ~n2318;
  assign n2320 = n1955 & n1998;
  assign n2321 = ~n1999 & ~n2320;
  assign n2322 = ~n2319 & n2321;
  assign n2323 = ~n1999 & ~n2322;
  assign n2324 = ~n125 & ~n341;
  assign n2325 = ~n220 & ~n329;
  assign n2326 = ~n238 & ~n310;
  assign n2327 = ~n458 & n2326;
  assign n2328 = n2032 & n2327;
  assign n2329 = ~n119 & ~n303;
  assign n2330 = ~n571 & n2329;
  assign n2331 = n828 & n2330;
  assign n2332 = n543 & n622;
  assign n2333 = n781 & n2243;
  assign n2334 = n2324 & n2325;
  assign n2335 = n2333 & n2334;
  assign n2336 = n2332 & n2335;
  assign n2337 = n2328 & n2331;
  assign n2338 = n2336 & n2337;
  assign n2339 = n764 & n972;
  assign n2340 = n2338 & n2339;
  assign n2341 = n2164 & n2340;
  assign n2342 = ~n604 & ~n663;
  assign n2343 = n604 & n663;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = ~n582 & ~n2344;
  assign n2346 = n582 & n2344;
  assign n2347 = ~n504 & ~n2345;
  assign n2348 = ~n2346 & n2347;
  assign n2349 = ~n1950 & ~n1953;
  assign n2350 = ~n1944 & ~n1947;
  assign n2351 = n2349 & ~n2350;
  assign n2352 = ~n2349 & n2350;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = n2348 & n2353;
  assign n2355 = ~n2348 & ~n2353;
  assign n2356 = ~n2354 & ~n2355;
  assign n2357 = ~n2341 & ~n2356;
  assign n2358 = n2341 & n2356;
  assign n2359 = ~n2357 & ~n2358;
  assign n2360 = ~n2323 & n2359;
  assign n2361 = n2323 & ~n2359;
  assign n2362 = ~n2360 & ~n2361;
  assign n2363 = pi2  & pi22 ;
  assign n2364 = pi2  & ~n50;
  assign n2365 = n1277 & ~n2364;
  assign n2366 = ~n2363 & ~n2365;
  assign n2367 = ~n1280 & ~n2366;
  assign n2368 = n1280 & n2366;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = ~n57 & ~n1201;
  assign n2371 = n57 & n1201;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = ~n2369 & n2372;
  assign n2374 = n2362 & n2373;
  assign n2375 = n2319 & ~n2321;
  assign n2376 = ~n2322 & ~n2375;
  assign n2377 = ~n1201 & ~n1280;
  assign n2378 = n1201 & n1280;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = n2369 & ~n2379;
  assign n2381 = n2376 & n2380;
  assign n2382 = n2315 & ~n2317;
  assign n2383 = ~n2318 & ~n2382;
  assign n2384 = n2369 & ~n2372;
  assign n2385 = n2379 & n2384;
  assign n2386 = n2383 & n2385;
  assign n2387 = ~n2369 & ~n2372;
  assign n2388 = n2376 & n2383;
  assign n2389 = n2311 & ~n2313;
  assign n2390 = ~n2314 & ~n2389;
  assign n2391 = n2383 & n2390;
  assign n2392 = n2307 & ~n2309;
  assign n2393 = ~n2310 & ~n2392;
  assign n2394 = n2390 & n2393;
  assign n2395 = n2303 & ~n2305;
  assign n2396 = ~n2306 & ~n2395;
  assign n2397 = n2393 & n2396;
  assign n2398 = n2299 & ~n2301;
  assign n2399 = ~n2302 & ~n2398;
  assign n2400 = n2396 & n2399;
  assign n2401 = n2295 & ~n2297;
  assign n2402 = ~n2298 & ~n2401;
  assign n2403 = n2399 & n2402;
  assign n2404 = n2291 & ~n2293;
  assign n2405 = ~n2294 & ~n2404;
  assign n2406 = n2402 & n2405;
  assign n2407 = n2287 & ~n2289;
  assign n2408 = ~n2290 & ~n2407;
  assign n2409 = n2405 & n2408;
  assign n2410 = ~n2405 & ~n2408;
  assign n2411 = ~n2409 & ~n2410;
  assign n2412 = ~n2272 & ~n2282;
  assign n2413 = ~n2283 & ~n2412;
  assign n2414 = ~n2408 & n2413;
  assign n2415 = n2283 & ~n2285;
  assign n2416 = ~n2286 & ~n2415;
  assign n2417 = ~n2414 & n2416;
  assign n2418 = n2411 & n2417;
  assign n2419 = ~n2409 & ~n2418;
  assign n2420 = ~n2402 & ~n2405;
  assign n2421 = ~n2406 & ~n2420;
  assign n2422 = ~n2419 & n2421;
  assign n2423 = ~n2406 & ~n2422;
  assign n2424 = ~n2399 & ~n2402;
  assign n2425 = ~n2403 & ~n2424;
  assign n2426 = ~n2423 & n2425;
  assign n2427 = ~n2403 & ~n2426;
  assign n2428 = ~n2396 & ~n2399;
  assign n2429 = ~n2400 & ~n2428;
  assign n2430 = ~n2427 & n2429;
  assign n2431 = ~n2400 & ~n2430;
  assign n2432 = ~n2393 & ~n2396;
  assign n2433 = ~n2397 & ~n2432;
  assign n2434 = ~n2431 & n2433;
  assign n2435 = ~n2397 & ~n2434;
  assign n2436 = ~n2390 & ~n2393;
  assign n2437 = ~n2394 & ~n2436;
  assign n2438 = ~n2435 & n2437;
  assign n2439 = ~n2394 & ~n2438;
  assign n2440 = ~n2383 & ~n2390;
  assign n2441 = ~n2391 & ~n2440;
  assign n2442 = ~n2439 & n2441;
  assign n2443 = ~n2391 & ~n2442;
  assign n2444 = ~n2376 & ~n2383;
  assign n2445 = ~n2388 & ~n2444;
  assign n2446 = ~n2443 & n2445;
  assign n2447 = ~n2388 & ~n2446;
  assign n2448 = n2362 & n2376;
  assign n2449 = ~n2362 & ~n2376;
  assign n2450 = ~n2448 & ~n2449;
  assign n2451 = ~n2447 & n2450;
  assign n2452 = n2447 & ~n2450;
  assign n2453 = ~n2451 & ~n2452;
  assign n2454 = n2387 & n2453;
  assign n2455 = ~n2381 & ~n2386;
  assign n2456 = ~n2374 & n2455;
  assign n2457 = ~n2454 & n2456;
  assign n2458 = n57 & ~n2457;
  assign n2459 = ~n57 & n2457;
  assign n2460 = ~n2458 & ~n2459;
  assign n2461 = ~n57 & ~n1045;
  assign n2462 = n57 & n1045;
  assign n2463 = ~n2461 & ~n2462;
  assign n2464 = ~n747 & ~n867;
  assign n2465 = n747 & n867;
  assign n2466 = ~n2464 & ~n2465;
  assign n2467 = ~n2463 & n2466;
  assign n2468 = n2393 & n2467;
  assign n2469 = ~n747 & ~n1045;
  assign n2470 = n747 & n1045;
  assign n2471 = ~n2469 & ~n2470;
  assign n2472 = n2463 & ~n2471;
  assign n2473 = n2396 & n2472;
  assign n2474 = n2463 & n2471;
  assign n2475 = ~n2466 & n2474;
  assign n2476 = n2399 & n2475;
  assign n2477 = ~n2463 & ~n2466;
  assign n2478 = n2431 & ~n2433;
  assign n2479 = ~n2434 & ~n2478;
  assign n2480 = n2477 & n2479;
  assign n2481 = ~n2473 & ~n2476;
  assign n2482 = ~n2468 & n2481;
  assign n2483 = ~n2480 & n2482;
  assign n2484 = n867 & ~n2483;
  assign n2485 = ~n867 & n2483;
  assign n2486 = ~n2484 & ~n2485;
  assign n2487 = ~n519 & ~n594;
  assign n2488 = n519 & n594;
  assign n2489 = ~n2487 & ~n2488;
  assign n2490 = ~n2413 & ~n2489;
  assign n2491 = ~n453 & ~n867;
  assign n2492 = n453 & n867;
  assign n2493 = ~n2491 & ~n2492;
  assign n2494 = ~n2413 & ~n2493;
  assign n2495 = ~n2413 & ~n2416;
  assign n2496 = ~n2285 & n2413;
  assign n2497 = ~n2495 & ~n2496;
  assign n2498 = ~n511 & ~n519;
  assign n2499 = n511 & n519;
  assign n2500 = ~n2498 & ~n2499;
  assign n2501 = ~n2493 & ~n2500;
  assign n2502 = ~n2497 & n2501;
  assign n2503 = ~n453 & ~n511;
  assign n2504 = n453 & n511;
  assign n2505 = ~n2503 & ~n2504;
  assign n2506 = n2493 & ~n2505;
  assign n2507 = ~n2413 & n2506;
  assign n2508 = ~n2493 & n2500;
  assign n2509 = n2416 & n2508;
  assign n2510 = ~n2507 & ~n2509;
  assign n2511 = ~n2502 & n2510;
  assign n2512 = n519 & ~n2494;
  assign n2513 = n2511 & n2512;
  assign n2514 = n2408 & n2508;
  assign n2515 = n2493 & ~n2500;
  assign n2516 = n2505 & n2515;
  assign n2517 = ~n2413 & n2516;
  assign n2518 = n2416 & n2506;
  assign n2519 = n2408 & ~n2496;
  assign n2520 = ~n2408 & n2496;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = n2501 & ~n2521;
  assign n2523 = ~n2517 & ~n2518;
  assign n2524 = ~n2514 & n2523;
  assign n2525 = ~n2522 & n2524;
  assign n2526 = n2513 & n2525;
  assign n2527 = n2490 & n2526;
  assign n2528 = n2405 & n2508;
  assign n2529 = n2416 & n2516;
  assign n2530 = n2408 & n2506;
  assign n2531 = ~n2411 & ~n2417;
  assign n2532 = ~n2418 & ~n2531;
  assign n2533 = n2501 & n2532;
  assign n2534 = ~n2529 & ~n2530;
  assign n2535 = ~n2528 & n2534;
  assign n2536 = ~n2533 & n2535;
  assign n2537 = n519 & ~n2536;
  assign n2538 = ~n519 & n2536;
  assign n2539 = ~n2537 & ~n2538;
  assign n2540 = ~n2490 & ~n2526;
  assign n2541 = ~n2527 & ~n2540;
  assign n2542 = n2539 & n2541;
  assign n2543 = ~n2527 & ~n2542;
  assign n2544 = n2402 & n2508;
  assign n2545 = n2405 & n2506;
  assign n2546 = n2408 & n2516;
  assign n2547 = n2419 & ~n2421;
  assign n2548 = ~n2422 & ~n2547;
  assign n2549 = n2501 & n2548;
  assign n2550 = ~n2545 & ~n2546;
  assign n2551 = ~n2544 & n2550;
  assign n2552 = ~n2549 & n2551;
  assign n2553 = ~n519 & n2552;
  assign n2554 = n519 & ~n2552;
  assign n2555 = ~n2553 & ~n2554;
  assign n2556 = ~n2344 & ~n2489;
  assign n2557 = ~n2497 & n2556;
  assign n2558 = ~n594 & ~n663;
  assign n2559 = n594 & n663;
  assign n2560 = ~n2558 & ~n2559;
  assign n2561 = n2489 & ~n2560;
  assign n2562 = ~n2413 & n2561;
  assign n2563 = n2344 & ~n2489;
  assign n2564 = n2416 & n2563;
  assign n2565 = ~n2562 & ~n2564;
  assign n2566 = ~n2557 & n2565;
  assign n2567 = ~n604 & ~n2413;
  assign n2568 = ~n2489 & n2567;
  assign n2569 = ~n2566 & n2568;
  assign n2570 = n2566 & ~n2568;
  assign n2571 = ~n2569 & ~n2570;
  assign n2572 = n2555 & n2571;
  assign n2573 = ~n2555 & ~n2571;
  assign n2574 = ~n2572 & ~n2573;
  assign n2575 = ~n2543 & n2574;
  assign n2576 = n2543 & ~n2574;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = ~n2486 & n2577;
  assign n2579 = n2396 & n2467;
  assign n2580 = n2399 & n2472;
  assign n2581 = n2402 & n2475;
  assign n2582 = n2427 & ~n2429;
  assign n2583 = ~n2430 & ~n2582;
  assign n2584 = n2477 & n2583;
  assign n2585 = ~n2580 & ~n2581;
  assign n2586 = ~n2579 & n2585;
  assign n2587 = ~n2584 & n2586;
  assign n2588 = n867 & n2587;
  assign n2589 = ~n867 & ~n2587;
  assign n2590 = ~n2588 & ~n2589;
  assign n2591 = ~n2539 & ~n2541;
  assign n2592 = ~n2542 & ~n2591;
  assign n2593 = n2590 & n2592;
  assign n2594 = n2399 & n2467;
  assign n2595 = n2402 & n2472;
  assign n2596 = n2405 & n2475;
  assign n2597 = n2423 & ~n2425;
  assign n2598 = ~n2426 & ~n2597;
  assign n2599 = n2477 & n2598;
  assign n2600 = ~n2595 & ~n2596;
  assign n2601 = ~n2594 & n2600;
  assign n2602 = ~n2599 & n2601;
  assign n2603 = n867 & ~n2602;
  assign n2604 = ~n867 & n2602;
  assign n2605 = ~n2603 & ~n2604;
  assign n2606 = n519 & ~n2513;
  assign n2607 = ~n2525 & n2606;
  assign n2608 = n2525 & ~n2606;
  assign n2609 = ~n2607 & ~n2608;
  assign n2610 = ~n2605 & n2609;
  assign n2611 = n2402 & n2467;
  assign n2612 = n2405 & n2472;
  assign n2613 = n2408 & n2475;
  assign n2614 = n2477 & n2548;
  assign n2615 = ~n2612 & ~n2613;
  assign n2616 = ~n2611 & n2615;
  assign n2617 = ~n2614 & n2616;
  assign n2618 = n867 & n2617;
  assign n2619 = ~n867 & ~n2617;
  assign n2620 = ~n2618 & ~n2619;
  assign n2621 = n519 & n2494;
  assign n2622 = ~n2511 & n2621;
  assign n2623 = n2511 & ~n2621;
  assign n2624 = ~n2622 & ~n2623;
  assign n2625 = n2620 & n2624;
  assign n2626 = ~n2413 & ~n2463;
  assign n2627 = n2477 & ~n2497;
  assign n2628 = ~n2413 & n2472;
  assign n2629 = n2416 & n2467;
  assign n2630 = ~n2628 & ~n2629;
  assign n2631 = ~n2627 & n2630;
  assign n2632 = ~n867 & ~n2626;
  assign n2633 = n2631 & n2632;
  assign n2634 = n2408 & n2467;
  assign n2635 = ~n2413 & n2475;
  assign n2636 = n2416 & n2472;
  assign n2637 = n2477 & ~n2521;
  assign n2638 = ~n2635 & ~n2636;
  assign n2639 = ~n2634 & n2638;
  assign n2640 = ~n2637 & n2639;
  assign n2641 = n2633 & n2640;
  assign n2642 = n2494 & n2641;
  assign n2643 = n2405 & n2467;
  assign n2644 = n2416 & n2475;
  assign n2645 = n2408 & n2472;
  assign n2646 = n2477 & n2532;
  assign n2647 = ~n2644 & ~n2645;
  assign n2648 = ~n2643 & n2647;
  assign n2649 = ~n2646 & n2648;
  assign n2650 = ~n867 & n2649;
  assign n2651 = n867 & ~n2649;
  assign n2652 = ~n2650 & ~n2651;
  assign n2653 = ~n2494 & ~n2641;
  assign n2654 = ~n2642 & ~n2653;
  assign n2655 = ~n2652 & n2654;
  assign n2656 = ~n2642 & ~n2655;
  assign n2657 = ~n2620 & ~n2624;
  assign n2658 = ~n2625 & ~n2657;
  assign n2659 = ~n2656 & n2658;
  assign n2660 = ~n2625 & ~n2659;
  assign n2661 = n2605 & ~n2609;
  assign n2662 = ~n2610 & ~n2661;
  assign n2663 = ~n2660 & n2662;
  assign n2664 = ~n2610 & ~n2663;
  assign n2665 = ~n2590 & ~n2592;
  assign n2666 = ~n2593 & ~n2665;
  assign n2667 = ~n2664 & n2666;
  assign n2668 = ~n2593 & ~n2667;
  assign n2669 = n2486 & ~n2577;
  assign n2670 = ~n2578 & ~n2669;
  assign n2671 = ~n2668 & n2670;
  assign n2672 = ~n2578 & ~n2671;
  assign n2673 = ~n2572 & ~n2575;
  assign n2674 = n2399 & n2508;
  assign n2675 = n2402 & n2506;
  assign n2676 = n2405 & n2516;
  assign n2677 = n2501 & n2598;
  assign n2678 = ~n2675 & ~n2676;
  assign n2679 = ~n2674 & n2678;
  assign n2680 = ~n2677 & n2679;
  assign n2681 = n519 & ~n2680;
  assign n2682 = ~n519 & n2680;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = ~n604 & ~n2490;
  assign n2685 = n2566 & n2684;
  assign n2686 = ~n604 & ~n2685;
  assign n2687 = n2408 & n2563;
  assign n2688 = n2489 & n2560;
  assign n2689 = ~n2344 & n2688;
  assign n2690 = ~n2413 & n2689;
  assign n2691 = n2416 & n2561;
  assign n2692 = ~n2521 & n2556;
  assign n2693 = ~n2690 & ~n2691;
  assign n2694 = ~n2687 & n2693;
  assign n2695 = ~n2692 & n2694;
  assign n2696 = n2686 & ~n2695;
  assign n2697 = ~n2686 & n2695;
  assign n2698 = ~n2696 & ~n2697;
  assign n2699 = n2683 & n2698;
  assign n2700 = ~n2683 & ~n2698;
  assign n2701 = ~n2699 & ~n2700;
  assign n2702 = n2673 & ~n2701;
  assign n2703 = ~n2673 & n2701;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = n2390 & n2467;
  assign n2706 = n2396 & n2475;
  assign n2707 = n2393 & n2472;
  assign n2708 = n2435 & ~n2437;
  assign n2709 = ~n2438 & ~n2708;
  assign n2710 = n2477 & n2709;
  assign n2711 = ~n2706 & ~n2707;
  assign n2712 = ~n2705 & n2711;
  assign n2713 = ~n2710 & n2712;
  assign n2714 = n867 & n2713;
  assign n2715 = ~n867 & ~n2713;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = n2704 & n2716;
  assign n2718 = ~n2704 & ~n2716;
  assign n2719 = ~n2717 & ~n2718;
  assign n2720 = ~n2672 & n2719;
  assign n2721 = n2672 & ~n2719;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = n2460 & n2722;
  assign n2724 = n2373 & n2376;
  assign n2725 = n2385 & n2390;
  assign n2726 = n2380 & n2383;
  assign n2727 = n2443 & ~n2445;
  assign n2728 = ~n2446 & ~n2727;
  assign n2729 = n2387 & n2728;
  assign n2730 = ~n2725 & ~n2726;
  assign n2731 = ~n2724 & n2730;
  assign n2732 = ~n2729 & n2731;
  assign n2733 = ~n57 & n2732;
  assign n2734 = n57 & ~n2732;
  assign n2735 = ~n2733 & ~n2734;
  assign n2736 = n2668 & ~n2670;
  assign n2737 = ~n2671 & ~n2736;
  assign n2738 = n2735 & n2737;
  assign n2739 = n2373 & n2383;
  assign n2740 = n2380 & n2390;
  assign n2741 = n2385 & n2393;
  assign n2742 = n2439 & ~n2441;
  assign n2743 = ~n2442 & ~n2742;
  assign n2744 = n2387 & n2743;
  assign n2745 = ~n2740 & ~n2741;
  assign n2746 = ~n2739 & n2745;
  assign n2747 = ~n2744 & n2746;
  assign n2748 = ~n57 & n2747;
  assign n2749 = n57 & ~n2747;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = n2664 & ~n2666;
  assign n2752 = ~n2667 & ~n2751;
  assign n2753 = n2750 & n2752;
  assign n2754 = n2373 & n2390;
  assign n2755 = n2385 & n2396;
  assign n2756 = n2380 & n2393;
  assign n2757 = n2387 & n2709;
  assign n2758 = ~n2755 & ~n2756;
  assign n2759 = ~n2754 & n2758;
  assign n2760 = ~n2757 & n2759;
  assign n2761 = ~n57 & n2760;
  assign n2762 = n57 & ~n2760;
  assign n2763 = ~n2761 & ~n2762;
  assign n2764 = n2660 & ~n2662;
  assign n2765 = ~n2663 & ~n2764;
  assign n2766 = n2763 & n2765;
  assign n2767 = n2373 & n2393;
  assign n2768 = n2380 & n2396;
  assign n2769 = n2385 & n2399;
  assign n2770 = n2387 & n2479;
  assign n2771 = ~n2768 & ~n2769;
  assign n2772 = ~n2767 & n2771;
  assign n2773 = ~n2770 & n2772;
  assign n2774 = n57 & ~n2773;
  assign n2775 = ~n57 & n2773;
  assign n2776 = ~n2774 & ~n2775;
  assign n2777 = n2656 & ~n2658;
  assign n2778 = ~n2659 & ~n2777;
  assign n2779 = n2776 & n2778;
  assign n2780 = n2373 & n2396;
  assign n2781 = n2380 & n2399;
  assign n2782 = n2385 & n2402;
  assign n2783 = n2387 & n2583;
  assign n2784 = ~n2781 & ~n2782;
  assign n2785 = ~n2780 & n2784;
  assign n2786 = ~n2783 & n2785;
  assign n2787 = ~n57 & n2786;
  assign n2788 = n57 & ~n2786;
  assign n2789 = ~n2787 & ~n2788;
  assign n2790 = n2652 & ~n2654;
  assign n2791 = ~n2655 & ~n2790;
  assign n2792 = n2789 & n2791;
  assign n2793 = n2373 & n2399;
  assign n2794 = n2380 & n2402;
  assign n2795 = n2385 & n2405;
  assign n2796 = n2387 & n2598;
  assign n2797 = ~n2794 & ~n2795;
  assign n2798 = ~n2793 & n2797;
  assign n2799 = ~n2796 & n2798;
  assign n2800 = n57 & ~n2799;
  assign n2801 = ~n57 & n2799;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = ~n867 & ~n2633;
  assign n2804 = ~n2640 & n2803;
  assign n2805 = n2640 & ~n2803;
  assign n2806 = ~n2804 & ~n2805;
  assign n2807 = n2802 & n2806;
  assign n2808 = n2373 & n2402;
  assign n2809 = n2380 & n2405;
  assign n2810 = n2385 & n2408;
  assign n2811 = n2387 & n2548;
  assign n2812 = ~n2809 & ~n2810;
  assign n2813 = ~n2808 & n2812;
  assign n2814 = ~n2811 & n2813;
  assign n2815 = ~n57 & n2814;
  assign n2816 = n57 & ~n2814;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = ~n867 & n2626;
  assign n2819 = ~n2631 & n2818;
  assign n2820 = n2631 & ~n2818;
  assign n2821 = ~n2819 & ~n2820;
  assign n2822 = n2817 & n2821;
  assign n2823 = ~n2369 & ~n2413;
  assign n2824 = n2387 & ~n2497;
  assign n2825 = n2380 & ~n2413;
  assign n2826 = n2373 & n2416;
  assign n2827 = ~n2825 & ~n2826;
  assign n2828 = ~n2824 & n2827;
  assign n2829 = n57 & ~n2823;
  assign n2830 = n2828 & n2829;
  assign n2831 = n2373 & n2408;
  assign n2832 = n2385 & ~n2413;
  assign n2833 = n2380 & n2416;
  assign n2834 = n2387 & ~n2521;
  assign n2835 = ~n2832 & ~n2833;
  assign n2836 = ~n2831 & n2835;
  assign n2837 = ~n2834 & n2836;
  assign n2838 = n2830 & n2837;
  assign n2839 = n2626 & n2838;
  assign n2840 = n2373 & n2405;
  assign n2841 = n2385 & n2416;
  assign n2842 = n2380 & n2408;
  assign n2843 = n2387 & n2532;
  assign n2844 = ~n2841 & ~n2842;
  assign n2845 = ~n2840 & n2844;
  assign n2846 = ~n2843 & n2845;
  assign n2847 = n57 & ~n2846;
  assign n2848 = ~n57 & n2846;
  assign n2849 = ~n2847 & ~n2848;
  assign n2850 = ~n2626 & ~n2838;
  assign n2851 = ~n2839 & ~n2850;
  assign n2852 = n2849 & n2851;
  assign n2853 = ~n2839 & ~n2852;
  assign n2854 = ~n2817 & ~n2821;
  assign n2855 = ~n2822 & ~n2854;
  assign n2856 = ~n2853 & n2855;
  assign n2857 = ~n2822 & ~n2856;
  assign n2858 = ~n2802 & ~n2806;
  assign n2859 = ~n2807 & ~n2858;
  assign n2860 = ~n2857 & n2859;
  assign n2861 = ~n2807 & ~n2860;
  assign n2862 = ~n2789 & ~n2791;
  assign n2863 = ~n2792 & ~n2862;
  assign n2864 = ~n2861 & n2863;
  assign n2865 = ~n2792 & ~n2864;
  assign n2866 = ~n2776 & ~n2778;
  assign n2867 = ~n2779 & ~n2866;
  assign n2868 = ~n2865 & n2867;
  assign n2869 = ~n2779 & ~n2868;
  assign n2870 = ~n2763 & ~n2765;
  assign n2871 = ~n2766 & ~n2870;
  assign n2872 = ~n2869 & n2871;
  assign n2873 = ~n2766 & ~n2872;
  assign n2874 = ~n2750 & ~n2752;
  assign n2875 = ~n2753 & ~n2874;
  assign n2876 = ~n2873 & n2875;
  assign n2877 = ~n2753 & ~n2876;
  assign n2878 = ~n2735 & ~n2737;
  assign n2879 = ~n2738 & ~n2878;
  assign n2880 = ~n2877 & n2879;
  assign n2881 = ~n2738 & ~n2880;
  assign n2882 = ~n2460 & ~n2722;
  assign n2883 = ~n2723 & ~n2882;
  assign n2884 = ~n2881 & n2883;
  assign n2885 = ~n2723 & ~n2884;
  assign n2886 = ~n2357 & ~n2360;
  assign n2887 = ~n119 & ~n223;
  assign n2888 = ~n247 & ~n314;
  assign n2889 = ~n384 & n2888;
  assign n2890 = n2887 & n2889;
  assign n2891 = n286 & n2890;
  assign n2892 = ~n272 & ~n378;
  assign n2893 = n346 & n521;
  assign n2894 = n776 & n1009;
  assign n2895 = n2892 & n2894;
  assign n2896 = n945 & n2893;
  assign n2897 = n2895 & n2896;
  assign n2898 = n610 & n2897;
  assign n2899 = n2128 & n2891;
  assign n2900 = n2898 & n2899;
  assign n2901 = n1290 & n2900;
  assign n2902 = n2886 & n2901;
  assign n2903 = ~n2886 & ~n2901;
  assign n2904 = ~n2902 & ~n2903;
  assign n2905 = n2373 & ~n2904;
  assign n2906 = n2376 & n2385;
  assign n2907 = n2362 & n2380;
  assign n2908 = ~n2448 & ~n2451;
  assign n2909 = n2362 & ~n2904;
  assign n2910 = ~n2362 & n2904;
  assign n2911 = ~n2909 & ~n2910;
  assign n2912 = ~n2908 & n2911;
  assign n2913 = n2908 & ~n2911;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = n2387 & n2914;
  assign n2916 = ~n2906 & ~n2907;
  assign n2917 = ~n2905 & n2916;
  assign n2918 = ~n2915 & n2917;
  assign n2919 = n57 & ~n2918;
  assign n2920 = ~n57 & n2918;
  assign n2921 = ~n2919 & ~n2920;
  assign n2922 = ~n2717 & ~n2720;
  assign n2923 = ~n2699 & ~n2703;
  assign n2924 = n2396 & n2508;
  assign n2925 = n2399 & n2506;
  assign n2926 = n2402 & n2516;
  assign n2927 = n2501 & n2583;
  assign n2928 = ~n2925 & ~n2926;
  assign n2929 = ~n2924 & n2928;
  assign n2930 = ~n2927 & n2929;
  assign n2931 = n519 & ~n2930;
  assign n2932 = ~n519 & n2930;
  assign n2933 = ~n2931 & ~n2932;
  assign n2934 = n2405 & n2563;
  assign n2935 = n2416 & n2689;
  assign n2936 = n2408 & n2561;
  assign n2937 = n2532 & n2556;
  assign n2938 = ~n2935 & ~n2936;
  assign n2939 = ~n2934 & n2938;
  assign n2940 = ~n2937 & n2939;
  assign n2941 = n604 & ~n2940;
  assign n2942 = ~n604 & n2940;
  assign n2943 = ~n2941 & ~n2942;
  assign n2944 = n2685 & n2695;
  assign n2945 = ~n2567 & ~n2944;
  assign n2946 = n2567 & n2944;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = ~n2943 & n2947;
  assign n2949 = n2943 & ~n2947;
  assign n2950 = ~n2948 & ~n2949;
  assign n2951 = n2933 & n2950;
  assign n2952 = ~n2933 & ~n2950;
  assign n2953 = ~n2951 & ~n2952;
  assign n2954 = n2923 & ~n2953;
  assign n2955 = ~n2923 & n2953;
  assign n2956 = ~n2954 & ~n2955;
  assign n2957 = n2383 & n2467;
  assign n2958 = n2390 & n2472;
  assign n2959 = n2393 & n2475;
  assign n2960 = n2477 & n2743;
  assign n2961 = ~n2958 & ~n2959;
  assign n2962 = ~n2957 & n2961;
  assign n2963 = ~n2960 & n2962;
  assign n2964 = n867 & n2963;
  assign n2965 = ~n867 & ~n2963;
  assign n2966 = ~n2964 & ~n2965;
  assign n2967 = n2956 & n2966;
  assign n2968 = ~n2956 & ~n2966;
  assign n2969 = ~n2967 & ~n2968;
  assign n2970 = ~n2922 & n2969;
  assign n2971 = n2922 & ~n2969;
  assign n2972 = ~n2970 & ~n2971;
  assign n2973 = n2921 & n2972;
  assign n2974 = ~n2921 & ~n2972;
  assign n2975 = ~n2973 & ~n2974;
  assign n2976 = n2885 & ~n2975;
  assign n2977 = ~n2885 & n2975;
  assign n2978 = ~n2976 & ~n2977;
  assign n2979 = ~n209 & ~n457;
  assign n2980 = ~n461 & n2979;
  assign n2981 = ~n520 & ~n571;
  assign n2982 = ~n186 & ~n403;
  assign n2983 = ~n181 & ~n325;
  assign n2984 = ~n355 & n2983;
  assign n2985 = n2273 & n2984;
  assign n2986 = ~n174 & ~n310;
  assign n2987 = n305 & n2986;
  assign n2988 = ~n218 & ~n241;
  assign n2989 = ~n264 & ~n294;
  assign n2990 = ~n299 & ~n542;
  assign n2991 = n2989 & n2990;
  assign n2992 = n2981 & n2988;
  assign n2993 = n2982 & n2992;
  assign n2994 = n1986 & n2991;
  assign n2995 = n2987 & n2994;
  assign n2996 = n2985 & n2993;
  assign n2997 = n2995 & n2996;
  assign n2998 = ~n273 & ~n329;
  assign n2999 = ~n268 & ~n298;
  assign n3000 = ~n314 & ~n433;
  assign n3001 = ~n546 & ~n560;
  assign n3002 = n3000 & n3001;
  assign n3003 = n409 & n2999;
  assign n3004 = n2998 & n3003;
  assign n3005 = n2145 & n3002;
  assign n3006 = n2980 & n3005;
  assign n3007 = n206 & n3004;
  assign n3008 = n3006 & n3007;
  assign n3009 = n169 & n3008;
  assign n3010 = n2997 & n3009;
  assign n3011 = n2902 & n3010;
  assign n3012 = ~n108 & ~n207;
  assign n3013 = ~n210 & ~n248;
  assign n3014 = n3012 & n3013;
  assign n3015 = n344 & n847;
  assign n3016 = n1006 & n2215;
  assign n3017 = n3015 & n3016;
  assign n3018 = n3014 & n3017;
  assign n3019 = n2022 & n2120;
  assign n3020 = n3018 & n3019;
  assign n3021 = n528 & n3020;
  assign n3022 = n498 & n3021;
  assign n3023 = n3011 & n3022;
  assign n3024 = ~n250 & ~n282;
  assign n3025 = n455 & n543;
  assign n3026 = n3024 & n3025;
  assign n3027 = n460 & n472;
  assign n3028 = n1026 & n3027;
  assign n3029 = n536 & n3026;
  assign n3030 = n3028 & n3029;
  assign n3031 = n490 & n528;
  assign n3032 = n578 & n3031;
  assign n3033 = n3030 & n3032;
  assign n3034 = n3023 & n3033;
  assign n3035 = ~n3023 & ~n3033;
  assign n3036 = ~n3034 & ~n3035;
  assign n3037 = pi0  & ~pi22 ;
  assign n3038 = pi1  & ~n3037;
  assign n3039 = ~pi1  & n3037;
  assign n3040 = ~n3038 & ~n3039;
  assign n3041 = n2366 & n3040;
  assign n3042 = ~n2366 & ~n3040;
  assign n3043 = ~n3041 & ~n3042;
  assign n3044 = pi0  & ~n3043;
  assign n3045 = ~n3036 & n3044;
  assign n3046 = ~n3011 & ~n3022;
  assign n3047 = ~n3023 & ~n3046;
  assign n3048 = ~pi0  & ~n3040;
  assign n3049 = ~n3047 & n3048;
  assign n3050 = ~n2902 & ~n3010;
  assign n3051 = ~n3011 & ~n3050;
  assign n3052 = pi2  & n50;
  assign n3053 = ~n3051 & n3052;
  assign n3054 = pi0  & n3043;
  assign n3055 = ~n3047 & ~n3051;
  assign n3056 = ~n2904 & ~n3051;
  assign n3057 = ~n2909 & ~n2912;
  assign n3058 = n2904 & n3010;
  assign n3059 = ~n3056 & ~n3058;
  assign n3060 = ~n3057 & n3059;
  assign n3061 = ~n3056 & ~n3060;
  assign n3062 = n3022 & n3051;
  assign n3063 = ~n3055 & ~n3062;
  assign n3064 = ~n3061 & n3063;
  assign n3065 = ~n3055 & ~n3064;
  assign n3066 = ~n3036 & ~n3047;
  assign n3067 = n3033 & n3047;
  assign n3068 = ~n3066 & ~n3067;
  assign n3069 = ~n3065 & n3068;
  assign n3070 = n3065 & ~n3068;
  assign n3071 = ~n3069 & ~n3070;
  assign n3072 = n3054 & n3071;
  assign n3073 = ~n3049 & ~n3053;
  assign n3074 = ~n3045 & n3073;
  assign n3075 = ~n3072 & n3074;
  assign n3076 = n2366 & n3075;
  assign n3077 = ~n2366 & ~n3075;
  assign n3078 = ~n3076 & ~n3077;
  assign n3079 = n2978 & n3078;
  assign n3080 = n2881 & ~n2883;
  assign n3081 = ~n2884 & ~n3080;
  assign n3082 = n3044 & ~n3047;
  assign n3083 = n3048 & ~n3051;
  assign n3084 = ~n2904 & n3052;
  assign n3085 = n3061 & ~n3063;
  assign n3086 = ~n3064 & ~n3085;
  assign n3087 = n3054 & n3086;
  assign n3088 = ~n3083 & ~n3084;
  assign n3089 = ~n3082 & n3088;
  assign n3090 = ~n3087 & n3089;
  assign n3091 = n2366 & n3090;
  assign n3092 = ~n2366 & ~n3090;
  assign n3093 = ~n3091 & ~n3092;
  assign n3094 = n3081 & n3093;
  assign n3095 = ~n3081 & ~n3093;
  assign n3096 = ~n3094 & ~n3095;
  assign n3097 = n2877 & ~n2879;
  assign n3098 = ~n2880 & ~n3097;
  assign n3099 = n2873 & ~n2875;
  assign n3100 = ~n2876 & ~n3099;
  assign n3101 = n2869 & ~n2871;
  assign n3102 = ~n2872 & ~n3101;
  assign n3103 = n2865 & ~n2867;
  assign n3104 = ~n2868 & ~n3103;
  assign n3105 = n2861 & ~n2863;
  assign n3106 = ~n2864 & ~n3105;
  assign n3107 = n2857 & ~n2859;
  assign n3108 = ~n2860 & ~n3107;
  assign n3109 = n2853 & ~n2855;
  assign n3110 = ~n2856 & ~n3109;
  assign n3111 = n2396 & n3044;
  assign n3112 = n2399 & n3048;
  assign n3113 = n2402 & n3052;
  assign n3114 = n2583 & n3054;
  assign n3115 = ~n3112 & ~n3113;
  assign n3116 = ~n3111 & n3115;
  assign n3117 = ~n3114 & n3116;
  assign n3118 = n2366 & ~n3117;
  assign n3119 = ~n2366 & n3117;
  assign n3120 = ~n3118 & ~n3119;
  assign n3121 = n57 & ~n2830;
  assign n3122 = ~n2837 & n3121;
  assign n3123 = n2837 & ~n3121;
  assign n3124 = ~n3122 & ~n3123;
  assign n3125 = n57 & n2823;
  assign n3126 = ~n2828 & n3125;
  assign n3127 = n2828 & ~n3125;
  assign n3128 = ~n3126 & ~n3127;
  assign n3129 = n2416 & n3048;
  assign n3130 = ~n2408 & n2497;
  assign n3131 = n3054 & ~n3130;
  assign n3132 = ~n2408 & ~n2416;
  assign n3133 = n3044 & ~n3132;
  assign n3134 = ~n51 & ~n2413;
  assign n3135 = ~n2366 & ~n3134;
  assign n3136 = ~n3129 & n3135;
  assign n3137 = ~n3131 & n3136;
  assign n3138 = ~n3133 & n3137;
  assign n3139 = n2823 & n3138;
  assign n3140 = ~n2823 & ~n3138;
  assign n3141 = n2532 & n3054;
  assign n3142 = n2405 & n3044;
  assign n3143 = n2408 & n3048;
  assign n3144 = ~n3142 & ~n3143;
  assign n3145 = ~n3141 & n3144;
  assign n3146 = n2366 & ~n3145;
  assign n3147 = n2416 & n3052;
  assign n3148 = ~n2366 & ~n3147;
  assign n3149 = n3145 & n3148;
  assign n3150 = ~n3146 & ~n3149;
  assign n3151 = ~n3140 & ~n3150;
  assign n3152 = ~n3139 & ~n3151;
  assign n3153 = n3128 & ~n3152;
  assign n3154 = ~n3128 & n3152;
  assign n3155 = n2402 & n3044;
  assign n3156 = n2405 & n3048;
  assign n3157 = n2408 & n3052;
  assign n3158 = n2548 & n3054;
  assign n3159 = ~n3156 & ~n3157;
  assign n3160 = ~n3155 & n3159;
  assign n3161 = ~n3158 & n3160;
  assign n3162 = ~n2366 & ~n3161;
  assign n3163 = n2366 & n3161;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = ~n3154 & n3164;
  assign n3166 = ~n3153 & ~n3165;
  assign n3167 = ~n3124 & n3166;
  assign n3168 = n3124 & ~n3166;
  assign n3169 = n2399 & n3044;
  assign n3170 = n2402 & n3048;
  assign n3171 = n2405 & n3052;
  assign n3172 = n2598 & n3054;
  assign n3173 = ~n3170 & ~n3171;
  assign n3174 = ~n3169 & n3173;
  assign n3175 = ~n3172 & n3174;
  assign n3176 = n2366 & ~n3175;
  assign n3177 = ~n2366 & n3175;
  assign n3178 = ~n3176 & ~n3177;
  assign n3179 = ~n3168 & n3178;
  assign n3180 = ~n3167 & ~n3179;
  assign n3181 = ~n3120 & n3180;
  assign n3182 = n3120 & ~n3180;
  assign n3183 = ~n2849 & ~n2851;
  assign n3184 = ~n2852 & ~n3183;
  assign n3185 = ~n3182 & n3184;
  assign n3186 = ~n3181 & ~n3185;
  assign n3187 = ~n3110 & n3186;
  assign n3188 = n3110 & ~n3186;
  assign n3189 = n2393 & n3044;
  assign n3190 = n2396 & n3048;
  assign n3191 = n2399 & n3052;
  assign n3192 = n2479 & n3054;
  assign n3193 = ~n3190 & ~n3191;
  assign n3194 = ~n3189 & n3193;
  assign n3195 = ~n3192 & n3194;
  assign n3196 = n2366 & ~n3195;
  assign n3197 = ~n2366 & n3195;
  assign n3198 = ~n3196 & ~n3197;
  assign n3199 = ~n3188 & n3198;
  assign n3200 = ~n3187 & ~n3199;
  assign n3201 = n3108 & n3200;
  assign n3202 = ~n3108 & ~n3200;
  assign n3203 = n2390 & n3044;
  assign n3204 = n2393 & n3048;
  assign n3205 = n2709 & n3054;
  assign n3206 = ~n3203 & ~n3204;
  assign n3207 = ~n3205 & n3206;
  assign n3208 = n2366 & ~n3207;
  assign n3209 = n50 & n2396;
  assign n3210 = ~n2366 & ~n3209;
  assign n3211 = n3207 & n3210;
  assign n3212 = ~n3208 & ~n3211;
  assign n3213 = ~n3202 & ~n3212;
  assign n3214 = ~n3201 & ~n3213;
  assign n3215 = n3106 & ~n3214;
  assign n3216 = ~n3106 & n3214;
  assign n3217 = n2383 & n3044;
  assign n3218 = n2390 & n3048;
  assign n3219 = n2393 & n3052;
  assign n3220 = n2743 & n3054;
  assign n3221 = ~n3218 & ~n3219;
  assign n3222 = ~n3217 & n3221;
  assign n3223 = ~n3220 & n3222;
  assign n3224 = ~n2366 & ~n3223;
  assign n3225 = n2366 & n3223;
  assign n3226 = ~n3224 & ~n3225;
  assign n3227 = ~n3216 & n3226;
  assign n3228 = ~n3215 & ~n3227;
  assign n3229 = n3104 & ~n3228;
  assign n3230 = ~n3104 & n3228;
  assign n3231 = n2376 & n3044;
  assign n3232 = n2383 & n3048;
  assign n3233 = n2728 & n3054;
  assign n3234 = ~n3231 & ~n3232;
  assign n3235 = ~n3233 & n3234;
  assign n3236 = n2366 & ~n3235;
  assign n3237 = n50 & n2390;
  assign n3238 = ~n2366 & ~n3237;
  assign n3239 = n3235 & n3238;
  assign n3240 = ~n3236 & ~n3239;
  assign n3241 = ~n3230 & ~n3240;
  assign n3242 = ~n3229 & ~n3241;
  assign n3243 = ~n3102 & n3242;
  assign n3244 = n3102 & ~n3242;
  assign n3245 = n2362 & n3044;
  assign n3246 = n2376 & n3048;
  assign n3247 = n2383 & n3052;
  assign n3248 = n2453 & n3054;
  assign n3249 = ~n3246 & ~n3247;
  assign n3250 = ~n3245 & n3249;
  assign n3251 = ~n3248 & n3250;
  assign n3252 = n2366 & ~n3251;
  assign n3253 = ~n2366 & n3251;
  assign n3254 = ~n3252 & ~n3253;
  assign n3255 = ~n3244 & n3254;
  assign n3256 = ~n3243 & ~n3255;
  assign n3257 = n3100 & n3256;
  assign n3258 = ~n3100 & ~n3256;
  assign n3259 = ~n2904 & n3044;
  assign n3260 = n2362 & n3048;
  assign n3261 = n2914 & n3054;
  assign n3262 = ~n3259 & ~n3260;
  assign n3263 = ~n3261 & n3262;
  assign n3264 = n2366 & ~n3263;
  assign n3265 = n50 & n2376;
  assign n3266 = ~n2366 & ~n3265;
  assign n3267 = n3263 & n3266;
  assign n3268 = ~n3264 & ~n3267;
  assign n3269 = ~n3258 & ~n3268;
  assign n3270 = ~n3257 & ~n3269;
  assign n3271 = ~n3098 & n3270;
  assign n3272 = n3098 & ~n3270;
  assign n3273 = n3044 & ~n3051;
  assign n3274 = ~n2904 & n3048;
  assign n3275 = n2362 & n3052;
  assign n3276 = n3057 & ~n3059;
  assign n3277 = ~n3060 & ~n3276;
  assign n3278 = n3054 & n3277;
  assign n3279 = ~n3274 & ~n3275;
  assign n3280 = ~n3273 & n3279;
  assign n3281 = ~n3278 & n3280;
  assign n3282 = n2366 & ~n3281;
  assign n3283 = ~n2366 & n3281;
  assign n3284 = ~n3282 & ~n3283;
  assign n3285 = ~n3272 & n3284;
  assign n3286 = ~n3271 & ~n3285;
  assign n3287 = n3096 & n3286;
  assign n3288 = ~n3094 & ~n3287;
  assign n3289 = ~n2978 & ~n3078;
  assign n3290 = ~n3079 & ~n3289;
  assign n3291 = ~n3288 & n3290;
  assign n3292 = ~n3079 & ~n3291;
  assign n3293 = ~n2973 & ~n2977;
  assign n3294 = n2373 & ~n3051;
  assign n3295 = n2380 & ~n2904;
  assign n3296 = n2362 & n2385;
  assign n3297 = n2387 & n3277;
  assign n3298 = ~n3295 & ~n3296;
  assign n3299 = ~n3294 & n3298;
  assign n3300 = ~n3297 & n3299;
  assign n3301 = n57 & ~n3300;
  assign n3302 = ~n57 & n3300;
  assign n3303 = ~n3301 & ~n3302;
  assign n3304 = ~n2967 & ~n2970;
  assign n3305 = n2376 & n2467;
  assign n3306 = n2390 & n2475;
  assign n3307 = n2383 & n2472;
  assign n3308 = n2477 & n2728;
  assign n3309 = ~n3306 & ~n3307;
  assign n3310 = ~n3305 & n3309;
  assign n3311 = ~n3308 & n3310;
  assign n3312 = n867 & n3311;
  assign n3313 = ~n867 & ~n3311;
  assign n3314 = ~n3312 & ~n3313;
  assign n3315 = ~n2951 & ~n2955;
  assign n3316 = n2393 & n2508;
  assign n3317 = n2396 & n2506;
  assign n3318 = n2399 & n2516;
  assign n3319 = n2479 & n2501;
  assign n3320 = ~n3317 & ~n3318;
  assign n3321 = ~n3316 & n3320;
  assign n3322 = ~n3319 & n3321;
  assign n3323 = n519 & ~n3322;
  assign n3324 = ~n519 & n3322;
  assign n3325 = ~n3323 & ~n3324;
  assign n3326 = ~n2946 & ~n2948;
  assign n3327 = ~n604 & ~n2416;
  assign n3328 = n2402 & n2563;
  assign n3329 = n2405 & n2561;
  assign n3330 = n2408 & n2689;
  assign n3331 = n2548 & n2556;
  assign n3332 = ~n3329 & ~n3330;
  assign n3333 = ~n3328 & n3332;
  assign n3334 = ~n3331 & n3333;
  assign n3335 = n3327 & ~n3334;
  assign n3336 = ~n3327 & n3334;
  assign n3337 = ~n3335 & ~n3336;
  assign n3338 = ~n3326 & n3337;
  assign n3339 = n3326 & ~n3337;
  assign n3340 = ~n3338 & ~n3339;
  assign n3341 = n3325 & n3340;
  assign n3342 = ~n3325 & ~n3340;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = ~n3315 & n3343;
  assign n3345 = n3315 & ~n3343;
  assign n3346 = ~n3344 & ~n3345;
  assign n3347 = n3314 & n3346;
  assign n3348 = ~n3314 & ~n3346;
  assign n3349 = ~n3347 & ~n3348;
  assign n3350 = ~n3304 & n3349;
  assign n3351 = n3304 & ~n3349;
  assign n3352 = ~n3350 & ~n3351;
  assign n3353 = n3303 & n3352;
  assign n3354 = ~n3303 & ~n3352;
  assign n3355 = ~n3353 & ~n3354;
  assign n3356 = ~n3293 & n3355;
  assign n3357 = n3293 & ~n3355;
  assign n3358 = ~n3356 & ~n3357;
  assign n3359 = n115 & n118;
  assign n3360 = n159 & n578;
  assign n3361 = ~n537 & ~n3359;
  assign n3362 = n468 & n3361;
  assign n3363 = n480 & n528;
  assign n3364 = n567 & n3363;
  assign n3365 = n3360 & n3362;
  assign n3366 = n3364 & n3365;
  assign n3367 = ~n3034 & ~n3366;
  assign n3368 = n3034 & n3366;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = n3044 & ~n3369;
  assign n3371 = ~n3036 & n3048;
  assign n3372 = ~n3047 & n3052;
  assign n3373 = ~n3066 & ~n3069;
  assign n3374 = ~n3036 & ~n3369;
  assign n3375 = n3036 & n3366;
  assign n3376 = ~n3374 & ~n3375;
  assign n3377 = ~n3373 & n3376;
  assign n3378 = n3373 & ~n3376;
  assign n3379 = ~n3377 & ~n3378;
  assign n3380 = n3054 & n3379;
  assign n3381 = ~n3371 & ~n3372;
  assign n3382 = ~n3370 & n3381;
  assign n3383 = ~n3380 & n3382;
  assign n3384 = n2366 & n3383;
  assign n3385 = ~n2366 & ~n3383;
  assign n3386 = ~n3384 & ~n3385;
  assign n3387 = n3358 & n3386;
  assign n3388 = ~n3358 & ~n3386;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = ~n3292 & n3389;
  assign n3391 = n3292 & ~n3389;
  assign n3392 = ~n3390 & ~n3391;
  assign n3393 = ~n192 & ~n225;
  assign n3394 = n483 & n3393;
  assign n3395 = n390 & n3394;
  assign n3396 = n2985 & n3395;
  assign n3397 = ~n108 & ~n542;
  assign n3398 = ~n185 & ~n248;
  assign n3399 = ~n171 & ~n272;
  assign n3400 = ~n314 & ~n537;
  assign n3401 = n3399 & n3400;
  assign n3402 = n2183 & n3401;
  assign n3403 = ~n134 & ~n152;
  assign n3404 = ~n219 & ~n222;
  assign n3405 = ~n433 & ~n454;
  assign n3406 = n3404 & n3405;
  assign n3407 = n398 & n3403;
  assign n3408 = n2030 & n3398;
  assign n3409 = n3407 & n3408;
  assign n3410 = n3406 & n3409;
  assign n3411 = n3402 & n3410;
  assign n3412 = ~n131 & ~n249;
  assign n3413 = n3397 & n3412;
  assign n3414 = n3411 & n3413;
  assign n3415 = ~n190 & ~n263;
  assign n3416 = ~n267 & ~n307;
  assign n3417 = ~n356 & n3416;
  assign n3418 = n605 & n3415;
  assign n3419 = n2324 & n2982;
  assign n3420 = n3418 & n3419;
  assign n3421 = n2980 & n3417;
  assign n3422 = n3420 & n3421;
  assign n3423 = n421 & n3422;
  assign n3424 = n3396 & n3423;
  assign n3425 = n3414 & n3424;
  assign n3426 = n3392 & ~n3425;
  assign n3427 = ~n3392 & n3425;
  assign n3428 = ~n3426 & ~n3427;
  assign n3429 = n3288 & ~n3290;
  assign n3430 = ~n3291 & ~n3429;
  assign n3431 = ~n188 & ~n198;
  assign n3432 = ~n297 & ~n317;
  assign n3433 = ~n403 & n3432;
  assign n3434 = n3431 & n3433;
  assign n3435 = ~n140 & ~n208;
  assign n3436 = ~n224 & ~n233;
  assign n3437 = n3435 & n3436;
  assign n3438 = n281 & n296;
  assign n3439 = n2998 & n3438;
  assign n3440 = n3437 & n3439;
  assign n3441 = n3434 & n3440;
  assign n3442 = ~n127 & ~n134;
  assign n3443 = ~n236 & ~n370;
  assign n3444 = ~n481 & n3443;
  assign n3445 = n2129 & n3442;
  assign n3446 = n330 & n3445;
  assign n3447 = n2155 & n3444;
  assign n3448 = n3446 & n3447;
  assign n3449 = n995 & n3448;
  assign n3450 = ~n145 & ~n279;
  assign n3451 = n302 & n3450;
  assign n3452 = n3449 & n3451;
  assign n3453 = ~n176 & ~n210;
  assign n3454 = ~n226 & ~n237;
  assign n3455 = ~n345 & n3454;
  assign n3456 = n813 & n3453;
  assign n3457 = n842 & n2981;
  assign n3458 = n3456 & n3457;
  assign n3459 = n3455 & n3458;
  assign n3460 = n2247 & n3459;
  assign n3461 = n3441 & n3460;
  assign n3462 = n3452 & n3461;
  assign n3463 = ~n3430 & n3462;
  assign n3464 = n3430 & ~n3462;
  assign n3465 = ~n298 & ~n304;
  assign n3466 = n1292 & n3465;
  assign n3467 = n459 & n3466;
  assign n3468 = n2067 & n3467;
  assign n3469 = n2100 & n3468;
  assign n3470 = ~n237 & ~n324;
  assign n3471 = n351 & n3470;
  assign n3472 = n2331 & n3471;
  assign n3473 = ~n152 & ~n218;
  assign n3474 = ~n222 & ~n251;
  assign n3475 = ~n315 & ~n329;
  assign n3476 = ~n384 & n3475;
  assign n3477 = n3473 & n3474;
  assign n3478 = n544 & n622;
  assign n3479 = n2211 & n2214;
  assign n3480 = n3478 & n3479;
  assign n3481 = n3476 & n3477;
  assign n3482 = n3480 & n3481;
  assign n3483 = n2169 & n3482;
  assign n3484 = n3469 & n3483;
  assign n3485 = n3472 & n3484;
  assign n3486 = ~n3096 & ~n3286;
  assign n3487 = ~n3287 & ~n3485;
  assign n3488 = ~n3486 & n3487;
  assign n3489 = ~n3464 & ~n3488;
  assign n3490 = ~n3463 & ~n3489;
  assign n3491 = n3428 & n3490;
  assign n3492 = ~n3426 & ~n3491;
  assign n3493 = ~n3387 & ~n3390;
  assign n3494 = ~n155 & ~n190;
  assign n3495 = ~n405 & ~n457;
  assign n3496 = n3494 & n3495;
  assign n3497 = n426 & n2044;
  assign n3498 = n3398 & n3497;
  assign n3499 = n3496 & n3498;
  assign n3500 = ~n131 & ~n133;
  assign n3501 = ~n144 & ~n152;
  assign n3502 = ~n219 & ~n315;
  assign n3503 = ~n554 & n3502;
  assign n3504 = n3500 & n3501;
  assign n3505 = n2215 & n2892;
  assign n3506 = n3504 & n3505;
  assign n3507 = n401 & n3503;
  assign n3508 = n3506 & n3507;
  assign n3509 = n2328 & n3508;
  assign n3510 = n3499 & n3509;
  assign n3511 = n1023 & n3510;
  assign n3512 = n3368 & n3511;
  assign n3513 = ~n3368 & ~n3511;
  assign n3514 = ~n3512 & ~n3513;
  assign n3515 = n3044 & ~n3514;
  assign n3516 = n3048 & ~n3369;
  assign n3517 = ~n3036 & n3052;
  assign n3518 = ~n3374 & ~n3377;
  assign n3519 = ~n3369 & ~n3514;
  assign n3520 = n3369 & n3511;
  assign n3521 = ~n3519 & ~n3520;
  assign n3522 = ~n3518 & n3521;
  assign n3523 = n3518 & ~n3521;
  assign n3524 = ~n3522 & ~n3523;
  assign n3525 = n3054 & n3524;
  assign n3526 = ~n3516 & ~n3517;
  assign n3527 = ~n3515 & n3526;
  assign n3528 = ~n3525 & n3527;
  assign n3529 = n2366 & ~n3528;
  assign n3530 = ~n2366 & n3528;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = ~n3353 & ~n3356;
  assign n3533 = ~n3347 & ~n3350;
  assign n3534 = n2362 & n2467;
  assign n3535 = n2376 & n2472;
  assign n3536 = n2383 & n2475;
  assign n3537 = n2453 & n2477;
  assign n3538 = ~n3535 & ~n3536;
  assign n3539 = ~n3534 & n3538;
  assign n3540 = ~n3537 & n3539;
  assign n3541 = n867 & ~n3540;
  assign n3542 = ~n867 & n3540;
  assign n3543 = ~n3541 & ~n3542;
  assign n3544 = ~n3341 & ~n3344;
  assign n3545 = ~n604 & ~n2408;
  assign n3546 = n2399 & n2563;
  assign n3547 = n2402 & n2561;
  assign n3548 = n2405 & n2689;
  assign n3549 = n2556 & n2598;
  assign n3550 = ~n3547 & ~n3548;
  assign n3551 = ~n3546 & n3550;
  assign n3552 = ~n3549 & n3551;
  assign n3553 = n3545 & ~n3552;
  assign n3554 = ~n3545 & n3552;
  assign n3555 = ~n3553 & ~n3554;
  assign n3556 = ~n604 & n2416;
  assign n3557 = n3334 & n3556;
  assign n3558 = ~n3338 & ~n3557;
  assign n3559 = n3555 & ~n3558;
  assign n3560 = ~n3555 & n3558;
  assign n3561 = ~n3559 & ~n3560;
  assign n3562 = n2390 & n2508;
  assign n3563 = n2396 & n2516;
  assign n3564 = n2393 & n2506;
  assign n3565 = n2501 & n2709;
  assign n3566 = ~n3563 & ~n3564;
  assign n3567 = ~n3562 & n3566;
  assign n3568 = ~n3565 & n3567;
  assign n3569 = ~n519 & n3568;
  assign n3570 = n519 & ~n3568;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = n3561 & n3571;
  assign n3573 = ~n3561 & ~n3571;
  assign n3574 = ~n3572 & ~n3573;
  assign n3575 = ~n3544 & n3574;
  assign n3576 = n3544 & ~n3574;
  assign n3577 = ~n3575 & ~n3576;
  assign n3578 = ~n3543 & n3577;
  assign n3579 = n3543 & ~n3577;
  assign n3580 = ~n3578 & ~n3579;
  assign n3581 = n3533 & ~n3580;
  assign n3582 = ~n3533 & n3580;
  assign n3583 = ~n3581 & ~n3582;
  assign n3584 = n2373 & ~n3047;
  assign n3585 = n2380 & ~n3051;
  assign n3586 = n2385 & ~n2904;
  assign n3587 = n2387 & n3086;
  assign n3588 = ~n3585 & ~n3586;
  assign n3589 = ~n3584 & n3588;
  assign n3590 = ~n3587 & n3589;
  assign n3591 = ~n57 & n3590;
  assign n3592 = n57 & ~n3590;
  assign n3593 = ~n3591 & ~n3592;
  assign n3594 = n3583 & n3593;
  assign n3595 = ~n3583 & ~n3593;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = ~n3532 & n3596;
  assign n3598 = n3532 & ~n3596;
  assign n3599 = ~n3597 & ~n3598;
  assign n3600 = ~n3531 & n3599;
  assign n3601 = n3531 & ~n3599;
  assign n3602 = ~n3600 & ~n3601;
  assign n3603 = n3493 & ~n3602;
  assign n3604 = ~n3493 & n3602;
  assign n3605 = ~n3603 & ~n3604;
  assign n3606 = ~n171 & ~n220;
  assign n3607 = ~n481 & n3606;
  assign n3608 = n786 & n3398;
  assign n3609 = n3607 & n3608;
  assign n3610 = n947 & n1282;
  assign n3611 = n2980 & n3610;
  assign n3612 = n645 & n3609;
  assign n3613 = n3611 & n3612;
  assign n3614 = n338 & n3613;
  assign n3615 = n2092 & n3614;
  assign n3616 = ~n3605 & n3615;
  assign n3617 = n3605 & ~n3615;
  assign n3618 = ~n3616 & ~n3617;
  assign n3619 = ~n3492 & n3618;
  assign n3620 = n3492 & ~n3618;
  assign n3621 = ~n3619 & ~n3620;
  assign n3622 = ~n3428 & ~n3490;
  assign n3623 = ~n3491 & ~n3622;
  assign n3624 = n3621 & n3623;
  assign n3625 = ~n3621 & ~n3623;
  assign po0  = ~n3624 & ~n3625;
  assign n3627 = ~n3617 & ~n3619;
  assign n3628 = ~n3600 & ~n3604;
  assign n3629 = ~n225 & ~n356;
  assign n3630 = n146 & n3629;
  assign n3631 = n383 & n2030;
  assign n3632 = n2211 & n3631;
  assign n3633 = n3630 & n3632;
  assign n3634 = n541 & n3633;
  assign n3635 = n761 & n847;
  assign n3636 = ~n201 & ~n226;
  assign n3637 = ~n310 & ~n377;
  assign n3638 = n3636 & n3637;
  assign n3639 = n379 & n3638;
  assign n3640 = n3635 & n3639;
  assign n3641 = n352 & n3640;
  assign n3642 = n1298 & n3641;
  assign n3643 = n3634 & n3642;
  assign n3644 = n2226 & n3643;
  assign n3645 = n3512 & ~n3644;
  assign n3646 = ~n3512 & n3644;
  assign n3647 = ~n3645 & ~n3646;
  assign n3648 = n3044 & n3647;
  assign n3649 = n3048 & ~n3514;
  assign n3650 = n3052 & ~n3369;
  assign n3651 = ~n3519 & ~n3522;
  assign n3652 = ~n3514 & ~n3647;
  assign n3653 = n3514 & ~n3644;
  assign n3654 = ~n3652 & ~n3653;
  assign n3655 = ~n3651 & ~n3654;
  assign n3656 = n3651 & n3654;
  assign n3657 = ~n3655 & ~n3656;
  assign n3658 = n3054 & n3657;
  assign n3659 = ~n3649 & ~n3650;
  assign n3660 = ~n3648 & n3659;
  assign n3661 = ~n3658 & n3660;
  assign n3662 = n2366 & ~n3661;
  assign n3663 = ~n2366 & n3661;
  assign n3664 = ~n3662 & ~n3663;
  assign n3665 = ~n3594 & ~n3597;
  assign n3666 = ~n3578 & ~n3582;
  assign n3667 = n2467 & ~n2904;
  assign n3668 = n2376 & n2475;
  assign n3669 = n2362 & n2472;
  assign n3670 = n2477 & n2914;
  assign n3671 = ~n3668 & ~n3669;
  assign n3672 = ~n3667 & n3671;
  assign n3673 = ~n3670 & n3672;
  assign n3674 = n867 & ~n3673;
  assign n3675 = ~n867 & n3673;
  assign n3676 = ~n3674 & ~n3675;
  assign n3677 = ~n3572 & ~n3575;
  assign n3678 = n2383 & n2508;
  assign n3679 = n2390 & n2506;
  assign n3680 = n2393 & n2516;
  assign n3681 = n2501 & n2743;
  assign n3682 = ~n3679 & ~n3680;
  assign n3683 = ~n3678 & n3682;
  assign n3684 = ~n3681 & n3683;
  assign n3685 = ~n519 & n3684;
  assign n3686 = n519 & ~n3684;
  assign n3687 = ~n3685 & ~n3686;
  assign n3688 = ~n604 & ~n2405;
  assign n3689 = n2396 & n2563;
  assign n3690 = n2399 & n2561;
  assign n3691 = n2402 & n2689;
  assign n3692 = n2556 & n2583;
  assign n3693 = ~n3690 & ~n3691;
  assign n3694 = ~n3689 & n3693;
  assign n3695 = ~n3692 & n3694;
  assign n3696 = n3688 & ~n3695;
  assign n3697 = ~n3688 & n3695;
  assign n3698 = ~n3696 & ~n3697;
  assign n3699 = ~n604 & n2408;
  assign n3700 = n3552 & n3699;
  assign n3701 = ~n3559 & ~n3700;
  assign n3702 = n3698 & ~n3701;
  assign n3703 = ~n3698 & n3701;
  assign n3704 = ~n3702 & ~n3703;
  assign n3705 = n3687 & n3704;
  assign n3706 = ~n3687 & ~n3704;
  assign n3707 = ~n3705 & ~n3706;
  assign n3708 = ~n3677 & n3707;
  assign n3709 = n3677 & ~n3707;
  assign n3710 = ~n3708 & ~n3709;
  assign n3711 = ~n3676 & n3710;
  assign n3712 = n3676 & ~n3710;
  assign n3713 = ~n3711 & ~n3712;
  assign n3714 = n3666 & ~n3713;
  assign n3715 = ~n3666 & n3713;
  assign n3716 = ~n3714 & ~n3715;
  assign n3717 = n2373 & ~n3036;
  assign n3718 = n2380 & ~n3047;
  assign n3719 = n2385 & ~n3051;
  assign n3720 = n2387 & n3071;
  assign n3721 = ~n3718 & ~n3719;
  assign n3722 = ~n3717 & n3721;
  assign n3723 = ~n3720 & n3722;
  assign n3724 = ~n57 & n3723;
  assign n3725 = n57 & ~n3723;
  assign n3726 = ~n3724 & ~n3725;
  assign n3727 = n3716 & n3726;
  assign n3728 = ~n3716 & ~n3726;
  assign n3729 = ~n3727 & ~n3728;
  assign n3730 = ~n3665 & n3729;
  assign n3731 = n3665 & ~n3729;
  assign n3732 = ~n3730 & ~n3731;
  assign n3733 = ~n3664 & n3732;
  assign n3734 = n3664 & ~n3732;
  assign n3735 = ~n3733 & ~n3734;
  assign n3736 = n3628 & ~n3735;
  assign n3737 = ~n3628 & n3735;
  assign n3738 = ~n3736 & ~n3737;
  assign n3739 = n958 & n1299;
  assign n3740 = ~n458 & n2121;
  assign n3741 = ~n127 & ~n181;
  assign n3742 = ~n324 & ~n353;
  assign n3743 = n3741 & n3742;
  assign n3744 = n146 & n639;
  assign n3745 = n1300 & n2979;
  assign n3746 = n3744 & n3745;
  assign n3747 = n2987 & n3743;
  assign n3748 = n3739 & n3740;
  assign n3749 = n3747 & n3748;
  assign n3750 = n3746 & n3749;
  assign n3751 = n2065 & n3750;
  assign n3752 = n3411 & n3751;
  assign n3753 = ~n3738 & n3752;
  assign n3754 = n3738 & ~n3752;
  assign n3755 = ~n3753 & ~n3754;
  assign n3756 = ~n3627 & n3755;
  assign n3757 = n3627 & ~n3755;
  assign n3758 = ~n3756 & ~n3757;
  assign n3759 = ~pi22  & ~pi23 ;
  assign n3760 = pi22  & pi23 ;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = po0  & n3761;
  assign n3763 = ~n3758 & n3762;
  assign n3764 = n3624 & n3758;
  assign n3765 = ~n3624 & ~n3758;
  assign n3766 = ~n3764 & ~n3765;
  assign n3767 = ~n3762 & n3766;
  assign po1  = n3763 | n3767;
  assign n3769 = ~n3754 & ~n3756;
  assign n3770 = ~n3733 & ~n3737;
  assign n3771 = ~n3727 & ~n3730;
  assign n3772 = ~n3711 & ~n3715;
  assign n3773 = n2467 & ~n3051;
  assign n3774 = n2472 & ~n2904;
  assign n3775 = n2362 & n2475;
  assign n3776 = n2477 & n3277;
  assign n3777 = ~n3774 & ~n3775;
  assign n3778 = ~n3773 & n3777;
  assign n3779 = ~n3776 & n3778;
  assign n3780 = n867 & ~n3779;
  assign n3781 = ~n867 & n3779;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = ~n3705 & ~n3708;
  assign n3784 = n2376 & n2508;
  assign n3785 = n2390 & n2516;
  assign n3786 = n2383 & n2506;
  assign n3787 = n2501 & n2728;
  assign n3788 = ~n3785 & ~n3786;
  assign n3789 = ~n3784 & n3788;
  assign n3790 = ~n3787 & n3789;
  assign n3791 = ~n519 & n3790;
  assign n3792 = n519 & ~n3790;
  assign n3793 = ~n3791 & ~n3792;
  assign n3794 = ~n604 & ~n2402;
  assign n3795 = n2393 & n2563;
  assign n3796 = n2396 & n2561;
  assign n3797 = n2399 & n2689;
  assign n3798 = n2479 & n2556;
  assign n3799 = ~n3796 & ~n3797;
  assign n3800 = ~n3795 & n3799;
  assign n3801 = ~n3798 & n3800;
  assign n3802 = n3794 & ~n3801;
  assign n3803 = ~n3794 & n3801;
  assign n3804 = ~n3802 & ~n3803;
  assign n3805 = ~n604 & n2405;
  assign n3806 = n3695 & n3805;
  assign n3807 = ~n3702 & ~n3806;
  assign n3808 = n3804 & ~n3807;
  assign n3809 = ~n3804 & n3807;
  assign n3810 = ~n3808 & ~n3809;
  assign n3811 = n3793 & n3810;
  assign n3812 = ~n3793 & ~n3810;
  assign n3813 = ~n3811 & ~n3812;
  assign n3814 = ~n3783 & n3813;
  assign n3815 = n3783 & ~n3813;
  assign n3816 = ~n3814 & ~n3815;
  assign n3817 = ~n3782 & n3816;
  assign n3818 = n3782 & ~n3816;
  assign n3819 = ~n3817 & ~n3818;
  assign n3820 = n3772 & ~n3819;
  assign n3821 = ~n3772 & n3819;
  assign n3822 = ~n3820 & ~n3821;
  assign n3823 = n2373 & ~n3369;
  assign n3824 = n2380 & ~n3036;
  assign n3825 = n2385 & ~n3047;
  assign n3826 = n2387 & n3379;
  assign n3827 = ~n3824 & ~n3825;
  assign n3828 = ~n3823 & n3827;
  assign n3829 = ~n3826 & n3828;
  assign n3830 = ~n57 & n3829;
  assign n3831 = n57 & ~n3829;
  assign n3832 = ~n3830 & ~n3831;
  assign n3833 = n3822 & n3832;
  assign n3834 = ~n3822 & ~n3832;
  assign n3835 = ~n3833 & ~n3834;
  assign n3836 = ~n3771 & n3835;
  assign n3837 = n3771 & ~n3835;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = n3048 & n3647;
  assign n3840 = ~n3647 & n3655;
  assign n3841 = n3653 & ~n3655;
  assign n3842 = ~n3840 & ~n3841;
  assign n3843 = n3054 & ~n3842;
  assign n3844 = ~n3839 & ~n3843;
  assign n3845 = n3052 & ~n3514;
  assign n3846 = ~n2366 & ~n3845;
  assign n3847 = n3844 & ~n3846;
  assign n3848 = ~n2366 & ~n3844;
  assign n3849 = ~n3847 & ~n3848;
  assign n3850 = n3838 & n3849;
  assign n3851 = ~n3838 & ~n3849;
  assign n3852 = ~n3850 & ~n3851;
  assign n3853 = ~n3770 & n3852;
  assign n3854 = n3770 & ~n3852;
  assign n3855 = ~n3853 & ~n3854;
  assign n3856 = ~n144 & ~n149;
  assign n3857 = ~n307 & n3856;
  assign n3858 = n1024 & n2325;
  assign n3859 = n3857 & n3858;
  assign n3860 = ~n207 & ~n233;
  assign n3861 = ~n310 & ~n343;
  assign n3862 = ~n345 & n3861;
  assign n3863 = n482 & n3860;
  assign n3864 = n614 & n3863;
  assign n3865 = n625 & n3862;
  assign n3866 = n3864 & n3865;
  assign n3867 = n3859 & n3866;
  assign n3868 = n293 & n3867;
  assign n3869 = n3469 & n3868;
  assign n3870 = n3855 & ~n3869;
  assign n3871 = ~n3855 & n3869;
  assign n3872 = ~n3870 & ~n3871;
  assign n3873 = ~n3769 & n3872;
  assign n3874 = n3769 & ~n3872;
  assign n3875 = ~n3873 & ~n3874;
  assign n3876 = ~n3764 & ~n3875;
  assign n3877 = n3764 & n3875;
  assign n3878 = ~n3876 & ~n3877;
  assign n3879 = ~po0  & ~n3766;
  assign n3880 = n3761 & ~n3879;
  assign n3881 = n3878 & ~n3880;
  assign n3882 = ~n3878 & n3880;
  assign po2  = n3881 | n3882;
  assign n3884 = ~n3878 & n3879;
  assign n3885 = n3761 & ~n3884;
  assign n3886 = ~n3870 & ~n3873;
  assign n3887 = ~n3850 & ~n3853;
  assign n3888 = ~n3833 & ~n3836;
  assign n3889 = n3514 & ~n3655;
  assign n3890 = n3054 & ~n3889;
  assign n3891 = ~n3052 & ~n3890;
  assign n3892 = n3647 & ~n3891;
  assign n3893 = n2366 & n3892;
  assign n3894 = ~n2366 & ~n3892;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = ~n3817 & ~n3821;
  assign n3897 = n2467 & ~n3047;
  assign n3898 = n2472 & ~n3051;
  assign n3899 = n2475 & ~n2904;
  assign n3900 = n2477 & n3086;
  assign n3901 = ~n3898 & ~n3899;
  assign n3902 = ~n3897 & n3901;
  assign n3903 = ~n3900 & n3902;
  assign n3904 = n867 & ~n3903;
  assign n3905 = ~n867 & n3903;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = ~n3811 & ~n3814;
  assign n3908 = n2362 & n2508;
  assign n3909 = n2376 & n2506;
  assign n3910 = n2383 & n2516;
  assign n3911 = n2453 & n2501;
  assign n3912 = ~n3909 & ~n3910;
  assign n3913 = ~n3908 & n3912;
  assign n3914 = ~n3911 & n3913;
  assign n3915 = ~n519 & n3914;
  assign n3916 = n519 & ~n3914;
  assign n3917 = ~n3915 & ~n3916;
  assign n3918 = ~n604 & ~n2399;
  assign n3919 = n2390 & n2563;
  assign n3920 = n2396 & n2689;
  assign n3921 = n2393 & n2561;
  assign n3922 = n2556 & n2709;
  assign n3923 = ~n3920 & ~n3921;
  assign n3924 = ~n3919 & n3923;
  assign n3925 = ~n3922 & n3924;
  assign n3926 = n3918 & ~n3925;
  assign n3927 = ~n3918 & n3925;
  assign n3928 = ~n3926 & ~n3927;
  assign n3929 = ~n604 & n2402;
  assign n3930 = n3801 & n3929;
  assign n3931 = ~n3808 & ~n3930;
  assign n3932 = n3928 & ~n3931;
  assign n3933 = ~n3928 & n3931;
  assign n3934 = ~n3932 & ~n3933;
  assign n3935 = n3917 & n3934;
  assign n3936 = ~n3917 & ~n3934;
  assign n3937 = ~n3935 & ~n3936;
  assign n3938 = ~n3907 & n3937;
  assign n3939 = n3907 & ~n3937;
  assign n3940 = ~n3938 & ~n3939;
  assign n3941 = ~n3906 & n3940;
  assign n3942 = n3906 & ~n3940;
  assign n3943 = ~n3941 & ~n3942;
  assign n3944 = n3896 & ~n3943;
  assign n3945 = ~n3896 & n3943;
  assign n3946 = ~n3944 & ~n3945;
  assign n3947 = n2373 & ~n3514;
  assign n3948 = n2380 & ~n3369;
  assign n3949 = n2385 & ~n3036;
  assign n3950 = n2387 & n3524;
  assign n3951 = ~n3948 & ~n3949;
  assign n3952 = ~n3947 & n3951;
  assign n3953 = ~n3950 & n3952;
  assign n3954 = ~n57 & n3953;
  assign n3955 = n57 & ~n3953;
  assign n3956 = ~n3954 & ~n3955;
  assign n3957 = n3946 & n3956;
  assign n3958 = ~n3946 & ~n3956;
  assign n3959 = ~n3957 & ~n3958;
  assign n3960 = ~n3895 & n3959;
  assign n3961 = n3895 & ~n3959;
  assign n3962 = ~n3960 & ~n3961;
  assign n3963 = ~n3888 & n3962;
  assign n3964 = n3888 & ~n3962;
  assign n3965 = ~n3963 & ~n3964;
  assign n3966 = ~n3887 & n3965;
  assign n3967 = n3887 & ~n3965;
  assign n3968 = ~n3966 & ~n3967;
  assign n3969 = ~n264 & ~n315;
  assign n3970 = ~n341 & ~n353;
  assign n3971 = ~n457 & n3970;
  assign n3972 = n2018 & n3969;
  assign n3973 = n3971 & n3972;
  assign n3974 = n777 & n3740;
  assign n3975 = n3973 & n3974;
  assign n3976 = n232 & n402;
  assign n3977 = n3434 & n3976;
  assign n3978 = n1960 & n3975;
  assign n3979 = n3977 & n3978;
  assign n3980 = n1290 & n3979;
  assign n3981 = n3968 & ~n3980;
  assign n3982 = ~n3968 & n3980;
  assign n3983 = ~n3981 & ~n3982;
  assign n3984 = ~n3886 & n3983;
  assign n3985 = n3886 & ~n3983;
  assign n3986 = ~n3984 & ~n3985;
  assign n3987 = n3877 & n3986;
  assign n3988 = ~n3877 & ~n3986;
  assign n3989 = ~n3987 & ~n3988;
  assign n3990 = n3885 & n3989;
  assign n3991 = ~n3885 & ~n3989;
  assign po3  = ~n3990 & ~n3991;
  assign n3993 = ~n3981 & ~n3984;
  assign n3994 = ~n3963 & ~n3966;
  assign n3995 = ~n3957 & ~n3960;
  assign n3996 = ~n3941 & ~n3945;
  assign n3997 = n2467 & ~n3036;
  assign n3998 = n2472 & ~n3047;
  assign n3999 = n2475 & ~n3051;
  assign n4000 = n2477 & n3071;
  assign n4001 = ~n3998 & ~n3999;
  assign n4002 = ~n3997 & n4001;
  assign n4003 = ~n4000 & n4002;
  assign n4004 = ~n867 & n4003;
  assign n4005 = n867 & ~n4003;
  assign n4006 = ~n4004 & ~n4005;
  assign n4007 = ~n3935 & ~n3938;
  assign n4008 = n2383 & n2563;
  assign n4009 = n2390 & n2561;
  assign n4010 = n2393 & n2689;
  assign n4011 = n2556 & n2743;
  assign n4012 = ~n4009 & ~n4010;
  assign n4013 = ~n4008 & n4012;
  assign n4014 = ~n4011 & n4013;
  assign n4015 = n604 & ~n4014;
  assign n4016 = ~n604 & n4014;
  assign n4017 = ~n4015 & ~n4016;
  assign n4018 = ~n604 & n2396;
  assign n4019 = ~n2366 & n4018;
  assign n4020 = n2366 & ~n4018;
  assign n4021 = ~n4019 & ~n4020;
  assign n4022 = ~n4017 & n4021;
  assign n4023 = n4017 & ~n4021;
  assign n4024 = ~n4022 & ~n4023;
  assign n4025 = ~n604 & n2399;
  assign n4026 = n3925 & n4025;
  assign n4027 = ~n3932 & ~n4026;
  assign n4028 = n4024 & ~n4027;
  assign n4029 = ~n4024 & n4027;
  assign n4030 = ~n4028 & ~n4029;
  assign n4031 = n2508 & ~n2904;
  assign n4032 = n2376 & n2516;
  assign n4033 = n2362 & n2506;
  assign n4034 = n2501 & n2914;
  assign n4035 = ~n4032 & ~n4033;
  assign n4036 = ~n4031 & n4035;
  assign n4037 = ~n4034 & n4036;
  assign n4038 = n519 & ~n4037;
  assign n4039 = ~n519 & n4037;
  assign n4040 = ~n4038 & ~n4039;
  assign n4041 = n4030 & n4040;
  assign n4042 = ~n4030 & ~n4040;
  assign n4043 = ~n4041 & ~n4042;
  assign n4044 = ~n4007 & n4043;
  assign n4045 = n4007 & ~n4043;
  assign n4046 = ~n4044 & ~n4045;
  assign n4047 = ~n4006 & n4046;
  assign n4048 = n4006 & ~n4046;
  assign n4049 = ~n4047 & ~n4048;
  assign n4050 = ~n3996 & n4049;
  assign n4051 = n3996 & ~n4049;
  assign n4052 = ~n4050 & ~n4051;
  assign n4053 = n2373 & n3647;
  assign n4054 = n2380 & ~n3514;
  assign n4055 = n2385 & ~n3369;
  assign n4056 = n2387 & n3657;
  assign n4057 = ~n4054 & ~n4055;
  assign n4058 = ~n4053 & n4057;
  assign n4059 = ~n4056 & n4058;
  assign n4060 = n57 & ~n4059;
  assign n4061 = ~n57 & n4059;
  assign n4062 = ~n4060 & ~n4061;
  assign n4063 = n4052 & n4062;
  assign n4064 = ~n4052 & ~n4062;
  assign n4065 = ~n4063 & ~n4064;
  assign n4066 = ~n3995 & n4065;
  assign n4067 = n3995 & ~n4065;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = n3994 & ~n4068;
  assign n4070 = ~n3994 & n4068;
  assign n4071 = ~n4069 & ~n4070;
  assign n4072 = ~n284 & ~n325;
  assign n4073 = ~n342 & n4072;
  assign n4074 = n347 & n572;
  assign n4075 = n637 & n2215;
  assign n4076 = n2325 & n4075;
  assign n4077 = n4073 & n4074;
  assign n4078 = n4076 & n4077;
  assign n4079 = n846 & n4078;
  assign n4080 = n217 & n4079;
  assign n4081 = n2257 & n4080;
  assign n4082 = ~n4071 & n4081;
  assign n4083 = n4071 & ~n4081;
  assign n4084 = ~n4082 & ~n4083;
  assign n4085 = ~n3993 & n4084;
  assign n4086 = n3993 & ~n4084;
  assign n4087 = ~n4085 & ~n4086;
  assign n4088 = ~n3987 & ~n4087;
  assign n4089 = n3987 & n4087;
  assign n4090 = ~n4088 & ~n4089;
  assign n4091 = n3884 & ~n3989;
  assign n4092 = n3761 & ~n4091;
  assign n4093 = n4090 & ~n4092;
  assign n4094 = ~n4090 & n4092;
  assign po4  = n4093 | n4094;
  assign n4096 = ~n4083 & ~n4085;
  assign n4097 = ~n4066 & ~n4070;
  assign n4098 = ~n4050 & ~n4063;
  assign n4099 = n2387 & ~n3842;
  assign n4100 = n2385 & ~n3514;
  assign n4101 = n2380 & n3647;
  assign n4102 = ~n4100 & ~n4101;
  assign n4103 = ~n4099 & n4102;
  assign n4104 = n57 & ~n4103;
  assign n4105 = ~n57 & n4103;
  assign n4106 = ~n4104 & ~n4105;
  assign n4107 = ~n4044 & ~n4047;
  assign n4108 = n2467 & ~n3369;
  assign n4109 = n2472 & ~n3036;
  assign n4110 = n2475 & ~n3047;
  assign n4111 = n2477 & n3379;
  assign n4112 = ~n4109 & ~n4110;
  assign n4113 = ~n4108 & n4112;
  assign n4114 = ~n4111 & n4113;
  assign n4115 = n867 & ~n4114;
  assign n4116 = ~n867 & n4114;
  assign n4117 = ~n4115 & ~n4116;
  assign n4118 = ~n4028 & ~n4041;
  assign n4119 = n2508 & ~n3051;
  assign n4120 = n2506 & ~n2904;
  assign n4121 = n2362 & n2516;
  assign n4122 = n2501 & n3277;
  assign n4123 = ~n4120 & ~n4121;
  assign n4124 = ~n4119 & n4123;
  assign n4125 = ~n4122 & n4124;
  assign n4126 = n519 & ~n4125;
  assign n4127 = ~n519 & n4125;
  assign n4128 = ~n4126 & ~n4127;
  assign n4129 = n2376 & n2563;
  assign n4130 = n2390 & n2689;
  assign n4131 = n2383 & n2561;
  assign n4132 = n2556 & n2728;
  assign n4133 = ~n4130 & ~n4131;
  assign n4134 = ~n4129 & n4133;
  assign n4135 = ~n4132 & n4134;
  assign n4136 = n604 & n4135;
  assign n4137 = ~n604 & ~n4135;
  assign n4138 = ~n4136 & ~n4137;
  assign n4139 = ~n4019 & ~n4022;
  assign n4140 = ~n604 & n2393;
  assign n4141 = ~n2366 & n4140;
  assign n4142 = n2366 & ~n4140;
  assign n4143 = ~n4141 & ~n4142;
  assign n4144 = ~n4139 & n4143;
  assign n4145 = n4139 & ~n4143;
  assign n4146 = ~n4144 & ~n4145;
  assign n4147 = n4138 & n4146;
  assign n4148 = ~n4138 & ~n4146;
  assign n4149 = ~n4147 & ~n4148;
  assign n4150 = n4128 & n4149;
  assign n4151 = ~n4128 & ~n4149;
  assign n4152 = ~n4150 & ~n4151;
  assign n4153 = ~n4118 & n4152;
  assign n4154 = n4118 & ~n4152;
  assign n4155 = ~n4153 & ~n4154;
  assign n4156 = ~n4117 & n4155;
  assign n4157 = n4117 & ~n4155;
  assign n4158 = ~n4156 & ~n4157;
  assign n4159 = ~n4107 & n4158;
  assign n4160 = n4107 & ~n4158;
  assign n4161 = ~n4159 & ~n4160;
  assign n4162 = n4106 & n4161;
  assign n4163 = ~n4106 & ~n4161;
  assign n4164 = ~n4162 & ~n4163;
  assign n4165 = ~n4098 & n4164;
  assign n4166 = n4098 & ~n4164;
  assign n4167 = ~n4165 & ~n4166;
  assign n4168 = ~n4097 & n4167;
  assign n4169 = n4097 & ~n4167;
  assign n4170 = ~n4168 & ~n4169;
  assign n4171 = ~n315 & n2213;
  assign n4172 = n483 & n2085;
  assign n4173 = ~n248 & ~n279;
  assign n4174 = ~n284 & ~n295;
  assign n4175 = n4173 & n4174;
  assign n4176 = n354 & n455;
  assign n4177 = n4175 & n4176;
  assign n4178 = n3739 & n4171;
  assign n4179 = n4172 & n4178;
  assign n4180 = n2104 & n4177;
  assign n4181 = n4179 & n4180;
  assign n4182 = n2997 & n4181;
  assign n4183 = n3634 & n4182;
  assign n4184 = ~n4170 & n4183;
  assign n4185 = n4170 & ~n4183;
  assign n4186 = ~n4184 & ~n4185;
  assign n4187 = ~n4096 & n4186;
  assign n4188 = n4096 & ~n4186;
  assign n4189 = ~n4187 & ~n4188;
  assign n4190 = ~n4089 & ~n4189;
  assign n4191 = n4089 & n4189;
  assign n4192 = ~n4190 & ~n4191;
  assign n4193 = ~n4090 & n4091;
  assign n4194 = n3761 & ~n4193;
  assign n4195 = n4192 & ~n4194;
  assign n4196 = ~n4192 & n4194;
  assign po5  = n4195 | n4196;
  assign n4198 = ~n4185 & ~n4187;
  assign n4199 = ~n4165 & ~n4168;
  assign n4200 = ~n4159 & ~n4162;
  assign n4201 = ~n4153 & ~n4156;
  assign n4202 = n2387 & ~n3889;
  assign n4203 = ~n2385 & ~n4202;
  assign n4204 = n3647 & ~n4203;
  assign n4205 = ~n57 & n4204;
  assign n4206 = n57 & ~n4204;
  assign n4207 = ~n4205 & ~n4206;
  assign n4208 = ~n4201 & ~n4207;
  assign n4209 = n4201 & n4207;
  assign n4210 = ~n4208 & ~n4209;
  assign n4211 = n2467 & ~n3514;
  assign n4212 = n2472 & ~n3369;
  assign n4213 = n2475 & ~n3036;
  assign n4214 = n2477 & n3524;
  assign n4215 = ~n4212 & ~n4213;
  assign n4216 = ~n4211 & n4215;
  assign n4217 = ~n4214 & n4216;
  assign n4218 = n867 & ~n4217;
  assign n4219 = ~n867 & n4217;
  assign n4220 = ~n4218 & ~n4219;
  assign n4221 = ~n4147 & ~n4150;
  assign n4222 = n2508 & ~n3047;
  assign n4223 = n2506 & ~n3051;
  assign n4224 = n2516 & ~n2904;
  assign n4225 = n2501 & n3086;
  assign n4226 = ~n4223 & ~n4224;
  assign n4227 = ~n4222 & n4226;
  assign n4228 = ~n4225 & n4227;
  assign n4229 = n519 & ~n4228;
  assign n4230 = ~n519 & n4228;
  assign n4231 = ~n4229 & ~n4230;
  assign n4232 = n2362 & n2563;
  assign n4233 = n2376 & n2561;
  assign n4234 = n2383 & n2689;
  assign n4235 = n2453 & n2556;
  assign n4236 = ~n4233 & ~n4234;
  assign n4237 = ~n4232 & n4236;
  assign n4238 = ~n4235 & n4237;
  assign n4239 = n604 & n4238;
  assign n4240 = ~n604 & ~n4238;
  assign n4241 = ~n4239 & ~n4240;
  assign n4242 = ~n4141 & ~n4144;
  assign n4243 = ~n604 & n2390;
  assign n4244 = ~n2366 & n4243;
  assign n4245 = n2366 & ~n4243;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = ~n4242 & n4246;
  assign n4248 = n4242 & ~n4246;
  assign n4249 = ~n4247 & ~n4248;
  assign n4250 = n4241 & n4249;
  assign n4251 = ~n4241 & ~n4249;
  assign n4252 = ~n4250 & ~n4251;
  assign n4253 = n4231 & n4252;
  assign n4254 = ~n4231 & ~n4252;
  assign n4255 = ~n4253 & ~n4254;
  assign n4256 = ~n4221 & n4255;
  assign n4257 = n4221 & ~n4255;
  assign n4258 = ~n4256 & ~n4257;
  assign n4259 = ~n4220 & n4258;
  assign n4260 = n4220 & ~n4258;
  assign n4261 = ~n4259 & ~n4260;
  assign n4262 = n4210 & n4261;
  assign n4263 = ~n4210 & ~n4261;
  assign n4264 = ~n4262 & ~n4263;
  assign n4265 = ~n4200 & n4264;
  assign n4266 = n4200 & ~n4264;
  assign n4267 = ~n4265 & ~n4266;
  assign n4268 = ~n4199 & n4267;
  assign n4269 = n4199 & ~n4267;
  assign n4270 = ~n4268 & ~n4269;
  assign n4271 = ~n309 & n409;
  assign n4272 = n2085 & n2121;
  assign n4273 = n2244 & n4272;
  assign n4274 = n425 & n4271;
  assign n4275 = n3635 & n4274;
  assign n4276 = n2218 & n4273;
  assign n4277 = n4275 & n4276;
  assign n4278 = ~n157 & ~n180;
  assign n4279 = ~n271 & ~n329;
  assign n4280 = n4278 & n4279;
  assign n4281 = n839 & n2084;
  assign n4282 = n3024 & n4281;
  assign n4283 = n2251 & n4280;
  assign n4284 = n4282 & n4283;
  assign n4285 = n4277 & n4284;
  assign n4286 = n3414 & n4285;
  assign n4287 = ~n4270 & n4286;
  assign n4288 = n4270 & ~n4286;
  assign n4289 = ~n4287 & ~n4288;
  assign n4290 = ~n4198 & n4289;
  assign n4291 = n4198 & ~n4289;
  assign n4292 = ~n4290 & ~n4291;
  assign n4293 = ~n4191 & ~n4292;
  assign n4294 = n4191 & n4292;
  assign n4295 = ~n4293 & ~n4294;
  assign n4296 = ~n4192 & n4193;
  assign n4297 = n3761 & ~n4296;
  assign n4298 = n4295 & ~n4297;
  assign n4299 = ~n4295 & n4297;
  assign po6  = n4298 | n4299;
  assign n4301 = ~n4288 & ~n4290;
  assign n4302 = ~n4265 & ~n4268;
  assign n4303 = ~n4208 & ~n4262;
  assign n4304 = ~n4256 & ~n4259;
  assign n4305 = n2467 & n3647;
  assign n4306 = n2472 & ~n3514;
  assign n4307 = n2475 & ~n3369;
  assign n4308 = n2477 & n3657;
  assign n4309 = ~n4306 & ~n4307;
  assign n4310 = ~n4305 & n4309;
  assign n4311 = ~n4308 & n4310;
  assign n4312 = n867 & n4311;
  assign n4313 = ~n867 & ~n4311;
  assign n4314 = ~n4312 & ~n4313;
  assign n4315 = ~n4304 & n4314;
  assign n4316 = n4304 & ~n4314;
  assign n4317 = ~n4315 & ~n4316;
  assign n4318 = ~n4250 & ~n4253;
  assign n4319 = ~n4244 & ~n4247;
  assign n4320 = n2563 & ~n2904;
  assign n4321 = n2376 & n2689;
  assign n4322 = n2362 & n2561;
  assign n4323 = n2556 & n2914;
  assign n4324 = ~n4321 & ~n4322;
  assign n4325 = ~n4320 & n4324;
  assign n4326 = ~n4323 & n4325;
  assign n4327 = n604 & ~n4326;
  assign n4328 = ~n604 & n4326;
  assign n4329 = ~n4327 & ~n4328;
  assign n4330 = ~n604 & n2383;
  assign n4331 = ~n57 & n2366;
  assign n4332 = n57 & ~n2366;
  assign n4333 = ~n4331 & ~n4332;
  assign n4334 = n4330 & n4333;
  assign n4335 = ~n4330 & ~n4333;
  assign n4336 = ~n4334 & ~n4335;
  assign n4337 = ~n4329 & n4336;
  assign n4338 = n4329 & ~n4336;
  assign n4339 = ~n4337 & ~n4338;
  assign n4340 = ~n4319 & n4339;
  assign n4341 = n4319 & ~n4339;
  assign n4342 = ~n4340 & ~n4341;
  assign n4343 = n2508 & ~n3036;
  assign n4344 = n2506 & ~n3047;
  assign n4345 = n2516 & ~n3051;
  assign n4346 = n2501 & n3071;
  assign n4347 = ~n4344 & ~n4345;
  assign n4348 = ~n4343 & n4347;
  assign n4349 = ~n4346 & n4348;
  assign n4350 = ~n519 & n4349;
  assign n4351 = n519 & ~n4349;
  assign n4352 = ~n4350 & ~n4351;
  assign n4353 = n4342 & n4352;
  assign n4354 = ~n4342 & ~n4352;
  assign n4355 = ~n4353 & ~n4354;
  assign n4356 = ~n4318 & n4355;
  assign n4357 = n4318 & ~n4355;
  assign n4358 = ~n4356 & ~n4357;
  assign n4359 = n4317 & n4358;
  assign n4360 = ~n4317 & ~n4358;
  assign n4361 = ~n4359 & ~n4360;
  assign n4362 = ~n4303 & n4361;
  assign n4363 = n4303 & ~n4361;
  assign n4364 = ~n4362 & ~n4363;
  assign n4365 = n4302 & ~n4364;
  assign n4366 = ~n4302 & n4364;
  assign n4367 = ~n4365 & ~n4366;
  assign n4368 = ~n152 & ~n325;
  assign n4369 = ~n127 & ~n307;
  assign n4370 = n239 & n4369;
  assign n4371 = n344 & n785;
  assign n4372 = n944 & n4368;
  assign n4373 = n4371 & n4372;
  assign n4374 = n4171 & n4370;
  assign n4375 = n4373 & n4374;
  assign n4376 = n4277 & n4375;
  assign n4377 = n2070 & n4376;
  assign n4378 = n4367 & ~n4377;
  assign n4379 = ~n4367 & n4377;
  assign n4380 = ~n4378 & ~n4379;
  assign n4381 = ~n4301 & n4380;
  assign n4382 = n4301 & ~n4380;
  assign n4383 = ~n4381 & ~n4382;
  assign n4384 = n4294 & n4383;
  assign n4385 = ~n4294 & ~n4383;
  assign n4386 = ~n4384 & ~n4385;
  assign n4387 = ~n4295 & n4296;
  assign n4388 = n3761 & ~n4387;
  assign n4389 = n4386 & ~n4388;
  assign n4390 = ~n4386 & n4388;
  assign po7  = n4389 | n4390;
  assign n4392 = ~n4378 & ~n4381;
  assign n4393 = ~n4362 & ~n4366;
  assign n4394 = ~n4315 & ~n4359;
  assign n4395 = n2477 & ~n3842;
  assign n4396 = n2475 & ~n3514;
  assign n4397 = n2472 & n3647;
  assign n4398 = ~n4396 & ~n4397;
  assign n4399 = ~n4395 & n4398;
  assign n4400 = n867 & ~n4399;
  assign n4401 = ~n867 & n4399;
  assign n4402 = ~n4400 & ~n4401;
  assign n4403 = ~n4353 & ~n4356;
  assign n4404 = n2508 & ~n3369;
  assign n4405 = n2506 & ~n3036;
  assign n4406 = n2516 & ~n3047;
  assign n4407 = n2501 & n3379;
  assign n4408 = ~n4405 & ~n4406;
  assign n4409 = ~n4404 & n4408;
  assign n4410 = ~n4407 & n4409;
  assign n4411 = n519 & ~n4410;
  assign n4412 = ~n519 & n4410;
  assign n4413 = ~n4411 & ~n4412;
  assign n4414 = ~n4337 & ~n4340;
  assign n4415 = n2563 & ~n3051;
  assign n4416 = n2561 & ~n2904;
  assign n4417 = n2362 & n2689;
  assign n4418 = n2556 & n3277;
  assign n4419 = ~n4416 & ~n4417;
  assign n4420 = ~n4415 & n4419;
  assign n4421 = ~n4418 & n4420;
  assign n4422 = n604 & n4421;
  assign n4423 = ~n604 & ~n4421;
  assign n4424 = ~n4422 & ~n4423;
  assign n4425 = ~n604 & n2376;
  assign n4426 = ~n4331 & ~n4334;
  assign n4427 = ~n4425 & ~n4426;
  assign n4428 = n4425 & n4426;
  assign n4429 = ~n4427 & ~n4428;
  assign n4430 = n4424 & n4429;
  assign n4431 = ~n4424 & ~n4429;
  assign n4432 = ~n4430 & ~n4431;
  assign n4433 = ~n4414 & n4432;
  assign n4434 = n4414 & ~n4432;
  assign n4435 = ~n4433 & ~n4434;
  assign n4436 = n4413 & n4435;
  assign n4437 = ~n4413 & ~n4435;
  assign n4438 = ~n4436 & ~n4437;
  assign n4439 = ~n4403 & n4438;
  assign n4440 = n4403 & ~n4438;
  assign n4441 = ~n4439 & ~n4440;
  assign n4442 = ~n4402 & n4441;
  assign n4443 = n4402 & ~n4441;
  assign n4444 = ~n4442 & ~n4443;
  assign n4445 = ~n4394 & n4444;
  assign n4446 = n4394 & ~n4444;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = ~n4393 & n4447;
  assign n4449 = n4393 & ~n4447;
  assign n4450 = ~n4448 & ~n4449;
  assign n4451 = ~n131 & ~n192;
  assign n4452 = ~n222 & n4451;
  assign n4453 = n316 & n547;
  assign n4454 = n2029 & n4453;
  assign n4455 = n4452 & n4454;
  assign n4456 = n1965 & n4455;
  assign n4457 = n421 & n4456;
  assign n4458 = ~n125 & ~n247;
  assign n4459 = ~n457 & ~n537;
  assign n4460 = ~n560 & n4459;
  assign n4461 = n2123 & n4458;
  assign n4462 = n4460 & n4461;
  assign n4463 = n834 & n2122;
  assign n4464 = n4462 & n4463;
  assign n4465 = n850 & n4464;
  assign n4466 = n3452 & n4465;
  assign n4467 = n4457 & n4466;
  assign n4468 = ~n4450 & n4467;
  assign n4469 = n4450 & ~n4467;
  assign n4470 = ~n4468 & ~n4469;
  assign n4471 = ~n4392 & n4470;
  assign n4472 = n4392 & ~n4470;
  assign n4473 = ~n4471 & ~n4472;
  assign n4474 = ~n4384 & ~n4473;
  assign n4475 = n4384 & n4473;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = ~n4386 & n4387;
  assign n4478 = n3761 & ~n4477;
  assign n4479 = n4476 & ~n4478;
  assign n4480 = ~n4476 & n4478;
  assign po8  = n4479 | n4480;
  assign n4482 = ~n4469 & ~n4471;
  assign n4483 = ~n4445 & ~n4448;
  assign n4484 = ~n4439 & ~n4442;
  assign n4485 = ~n4433 & ~n4436;
  assign n4486 = n2477 & ~n3889;
  assign n4487 = ~n2475 & ~n4486;
  assign n4488 = n3647 & ~n4487;
  assign n4489 = ~n867 & ~n4488;
  assign n4490 = n867 & n4488;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = ~n4485 & ~n4491;
  assign n4493 = n4485 & n4491;
  assign n4494 = ~n4492 & ~n4493;
  assign n4495 = ~n4427 & ~n4430;
  assign n4496 = n2563 & ~n3047;
  assign n4497 = n2561 & ~n3051;
  assign n4498 = n2689 & ~n2904;
  assign n4499 = n2556 & n3086;
  assign n4500 = ~n4497 & ~n4498;
  assign n4501 = ~n4496 & n4500;
  assign n4502 = ~n4499 & n4501;
  assign n4503 = n604 & ~n4502;
  assign n4504 = ~n604 & n4502;
  assign n4505 = ~n4503 & ~n4504;
  assign n4506 = ~n604 & n2450;
  assign n4507 = ~n4505 & ~n4506;
  assign n4508 = n4505 & n4506;
  assign n4509 = ~n4507 & ~n4508;
  assign n4510 = ~n4495 & n4509;
  assign n4511 = n4495 & ~n4509;
  assign n4512 = ~n4510 & ~n4511;
  assign n4513 = n2508 & ~n3514;
  assign n4514 = n2506 & ~n3369;
  assign n4515 = n2516 & ~n3036;
  assign n4516 = n2501 & n3524;
  assign n4517 = ~n4514 & ~n4515;
  assign n4518 = ~n4513 & n4517;
  assign n4519 = ~n4516 & n4518;
  assign n4520 = n519 & ~n4519;
  assign n4521 = ~n519 & n4519;
  assign n4522 = ~n4520 & ~n4521;
  assign n4523 = n4512 & n4522;
  assign n4524 = ~n4512 & ~n4522;
  assign n4525 = ~n4523 & ~n4524;
  assign n4526 = n4494 & n4525;
  assign n4527 = ~n4494 & ~n4525;
  assign n4528 = ~n4526 & ~n4527;
  assign n4529 = ~n4484 & n4528;
  assign n4530 = n4484 & ~n4528;
  assign n4531 = ~n4529 & ~n4530;
  assign n4532 = n4483 & ~n4531;
  assign n4533 = ~n4483 & n4531;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = ~n171 & ~n200;
  assign n4536 = ~n280 & ~n311;
  assign n4537 = ~n458 & n4536;
  assign n4538 = n344 & n4535;
  assign n4539 = n2095 & n3024;
  assign n4540 = n4538 & n4539;
  assign n4541 = n2987 & n4537;
  assign n4542 = n4540 & n4541;
  assign n4543 = n161 & n4542;
  assign n4544 = n3396 & n4543;
  assign n4545 = n2226 & n4544;
  assign n4546 = ~n4534 & n4545;
  assign n4547 = n4534 & ~n4545;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = ~n4482 & n4548;
  assign n4550 = n4482 & ~n4548;
  assign n4551 = ~n4549 & ~n4550;
  assign n4552 = ~n4475 & ~n4551;
  assign n4553 = n4475 & n4551;
  assign n4554 = ~n4552 & ~n4553;
  assign n4555 = ~n4476 & n4477;
  assign n4556 = n3761 & ~n4555;
  assign n4557 = n4554 & ~n4556;
  assign n4558 = ~n4554 & n4556;
  assign po9  = n4557 | n4558;
  assign n4560 = ~n4547 & ~n4549;
  assign n4561 = ~n4529 & ~n4533;
  assign n4562 = ~n4492 & ~n4526;
  assign n4563 = ~n4510 & ~n4523;
  assign n4564 = n2508 & n3647;
  assign n4565 = n2506 & ~n3514;
  assign n4566 = n2516 & ~n3369;
  assign n4567 = n2501 & n3657;
  assign n4568 = ~n4565 & ~n4566;
  assign n4569 = ~n4564 & n4568;
  assign n4570 = ~n4567 & n4569;
  assign n4571 = ~n519 & n4570;
  assign n4572 = n519 & ~n4570;
  assign n4573 = ~n4571 & ~n4572;
  assign n4574 = ~n4563 & n4573;
  assign n4575 = n4563 & ~n4573;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = n2563 & ~n3036;
  assign n4578 = n2561 & ~n3047;
  assign n4579 = n2689 & ~n3051;
  assign n4580 = n2556 & n3071;
  assign n4581 = ~n4578 & ~n4579;
  assign n4582 = ~n4577 & n4581;
  assign n4583 = ~n4580 & n4582;
  assign n4584 = ~n604 & n4583;
  assign n4585 = n604 & ~n4583;
  assign n4586 = ~n4584 & ~n4585;
  assign n4587 = ~n604 & ~n2904;
  assign n4588 = ~n867 & ~n4587;
  assign n4589 = n867 & n4587;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = n4425 & ~n4590;
  assign n4592 = ~n4425 & n4590;
  assign n4593 = ~n4591 & ~n4592;
  assign n4594 = ~n604 & ~n2376;
  assign n4595 = n2362 & n4594;
  assign n4596 = ~n4507 & ~n4595;
  assign n4597 = ~n4593 & ~n4596;
  assign n4598 = n4593 & n4596;
  assign n4599 = ~n4597 & ~n4598;
  assign n4600 = n4586 & ~n4599;
  assign n4601 = ~n4586 & n4599;
  assign n4602 = ~n4600 & ~n4601;
  assign n4603 = n4576 & n4602;
  assign n4604 = ~n4576 & ~n4602;
  assign n4605 = ~n4603 & ~n4604;
  assign n4606 = ~n4562 & n4605;
  assign n4607 = n4562 & ~n4605;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = ~n4561 & n4608;
  assign n4610 = n4561 & ~n4608;
  assign n4611 = ~n4609 & ~n4610;
  assign n4612 = ~n234 & ~n399;
  assign n4613 = ~n469 & n4612;
  assign n4614 = n330 & n2324;
  assign n4615 = n3024 & n4614;
  assign n4616 = n184 & n4613;
  assign n4617 = n848 & n2980;
  assign n4618 = n4616 & n4617;
  assign n4619 = n4615 & n4618;
  assign n4620 = n612 & n4619;
  assign n4621 = n955 & n3441;
  assign n4622 = n4620 & n4621;
  assign n4623 = ~n4611 & n4622;
  assign n4624 = n4611 & ~n4622;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = ~n4560 & n4625;
  assign n4627 = n4560 & ~n4625;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = ~n4553 & ~n4628;
  assign n4630 = n4553 & n4628;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = ~n4554 & n4555;
  assign n4633 = n3761 & ~n4632;
  assign n4634 = n4631 & ~n4633;
  assign n4635 = ~n4631 & n4633;
  assign po10  = n4634 | n4635;
  assign n4637 = ~n4624 & ~n4626;
  assign n4638 = ~n4606 & ~n4609;
  assign n4639 = ~n4574 & ~n4603;
  assign n4640 = n2501 & ~n3842;
  assign n4641 = n2516 & ~n3514;
  assign n4642 = n2506 & n3647;
  assign n4643 = ~n4641 & ~n4642;
  assign n4644 = ~n4640 & n4643;
  assign n4645 = n519 & ~n4644;
  assign n4646 = ~n519 & n4644;
  assign n4647 = ~n4645 & ~n4646;
  assign n4648 = n2563 & ~n3369;
  assign n4649 = n2561 & ~n3036;
  assign n4650 = n2689 & ~n3047;
  assign n4651 = n2556 & n3379;
  assign n4652 = ~n4649 & ~n4650;
  assign n4653 = ~n4648 & n4652;
  assign n4654 = ~n4651 & n4653;
  assign n4655 = n604 & n4654;
  assign n4656 = ~n604 & ~n4654;
  assign n4657 = ~n4655 & ~n4656;
  assign n4658 = ~n604 & ~n3051;
  assign n4659 = ~n4425 & ~n4589;
  assign n4660 = ~n4588 & ~n4659;
  assign n4661 = ~n4658 & n4660;
  assign n4662 = n4658 & ~n4660;
  assign n4663 = ~n4661 & ~n4662;
  assign n4664 = n4657 & n4663;
  assign n4665 = ~n4657 & ~n4663;
  assign n4666 = ~n4664 & ~n4665;
  assign n4667 = n4586 & ~n4597;
  assign n4668 = ~n4598 & ~n4667;
  assign n4669 = n4666 & n4668;
  assign n4670 = ~n4666 & ~n4668;
  assign n4671 = ~n4669 & ~n4670;
  assign n4672 = n4647 & n4671;
  assign n4673 = ~n4647 & ~n4671;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = ~n4639 & n4674;
  assign n4676 = n4639 & ~n4674;
  assign n4677 = ~n4675 & ~n4676;
  assign n4678 = ~n4638 & n4677;
  assign n4679 = n4638 & ~n4677;
  assign n4680 = ~n4678 & ~n4679;
  assign n4681 = ~n303 & n754;
  assign n4682 = n841 & n4681;
  assign n4683 = n536 & n4682;
  assign n4684 = n575 & n4683;
  assign n4685 = n3499 & n4684;
  assign n4686 = n636 & n4685;
  assign n4687 = ~n4680 & n4686;
  assign n4688 = n4680 & ~n4686;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = ~n4637 & n4689;
  assign n4691 = n4637 & ~n4689;
  assign n4692 = ~n4690 & ~n4691;
  assign n4693 = ~n4630 & ~n4692;
  assign n4694 = n4630 & n4692;
  assign n4695 = ~n4693 & ~n4694;
  assign n4696 = ~n4631 & n4632;
  assign n4697 = n3761 & ~n4696;
  assign n4698 = n4695 & ~n4697;
  assign n4699 = ~n4695 & n4697;
  assign po11  = n4698 | n4699;
  assign n4701 = ~n4688 & ~n4690;
  assign n4702 = ~n4675 & ~n4678;
  assign n4703 = ~n4669 & ~n4672;
  assign n4704 = ~n4661 & ~n4664;
  assign n4705 = ~n604 & n3063;
  assign n4706 = ~n4704 & ~n4705;
  assign n4707 = n4704 & n4705;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = n2563 & ~n3514;
  assign n4710 = n2561 & ~n3369;
  assign n4711 = n2689 & ~n3036;
  assign n4712 = n2556 & n3524;
  assign n4713 = ~n4710 & ~n4711;
  assign n4714 = ~n4709 & n4713;
  assign n4715 = ~n4712 & n4714;
  assign n4716 = ~n604 & n4715;
  assign n4717 = n604 & ~n4715;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = n2501 & ~n3889;
  assign n4720 = ~n2516 & ~n4719;
  assign n4721 = n3647 & ~n4720;
  assign n4722 = ~n519 & n4721;
  assign n4723 = n519 & ~n4721;
  assign n4724 = ~n4722 & ~n4723;
  assign n4725 = ~n4718 & ~n4724;
  assign n4726 = n4718 & n4724;
  assign n4727 = ~n4725 & ~n4726;
  assign n4728 = n4708 & n4727;
  assign n4729 = ~n4708 & ~n4727;
  assign n4730 = ~n4728 & ~n4729;
  assign n4731 = ~n4703 & n4730;
  assign n4732 = n4703 & ~n4730;
  assign n4733 = ~n4731 & ~n4732;
  assign n4734 = ~n4702 & n4733;
  assign n4735 = n4702 & ~n4733;
  assign n4736 = ~n4734 & ~n4735;
  assign n4737 = n115 & n126;
  assign n4738 = ~n133 & ~n273;
  assign n4739 = ~n372 & ~n457;
  assign n4740 = ~n571 & n4739;
  assign n4741 = n4738 & n4740;
  assign n4742 = ~n131 & ~n4737;
  assign n4743 = n2146 & n4742;
  assign n4744 = n777 & n4743;
  assign n4745 = n3859 & n4744;
  assign n4746 = n4741 & n4745;
  assign n4747 = n2028 & n4746;
  assign n4748 = n2162 & n4747;
  assign n4749 = ~n4736 & n4748;
  assign n4750 = n4736 & ~n4748;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = ~n4701 & n4751;
  assign n4753 = n4701 & ~n4751;
  assign n4754 = ~n4752 & ~n4753;
  assign n4755 = ~n4694 & ~n4754;
  assign n4756 = n4694 & n4754;
  assign n4757 = ~n4755 & ~n4756;
  assign n4758 = ~n4695 & n4696;
  assign n4759 = n3761 & ~n4758;
  assign n4760 = n4757 & ~n4759;
  assign n4761 = ~n4757 & n4759;
  assign po12  = n4760 | n4761;
  assign n4763 = ~n4750 & ~n4752;
  assign n4764 = ~n4731 & ~n4734;
  assign n4765 = ~n4725 & ~n4728;
  assign n4766 = n3047 & n4658;
  assign n4767 = ~n4706 & ~n4766;
  assign n4768 = n2563 & n3647;
  assign n4769 = n2561 & ~n3514;
  assign n4770 = n2689 & ~n3369;
  assign n4771 = n2556 & n3657;
  assign n4772 = ~n4769 & ~n4770;
  assign n4773 = ~n4768 & n4772;
  assign n4774 = ~n4771 & n4773;
  assign n4775 = n604 & ~n4774;
  assign n4776 = ~n604 & n4774;
  assign n4777 = ~n4775 & ~n4776;
  assign n4778 = ~n604 & ~n3047;
  assign n4779 = ~n519 & n4778;
  assign n4780 = n519 & ~n4778;
  assign n4781 = ~n4779 & ~n4780;
  assign n4782 = ~n604 & ~n3036;
  assign n4783 = n4781 & n4782;
  assign n4784 = ~n4781 & ~n4782;
  assign n4785 = ~n4783 & ~n4784;
  assign n4786 = ~n4777 & n4785;
  assign n4787 = n4777 & ~n4785;
  assign n4788 = ~n4786 & ~n4787;
  assign n4789 = ~n4767 & n4788;
  assign n4790 = n4767 & ~n4788;
  assign n4791 = ~n4789 & ~n4790;
  assign n4792 = ~n4765 & n4791;
  assign n4793 = n4765 & ~n4791;
  assign n4794 = ~n4792 & ~n4793;
  assign n4795 = ~n4764 & n4794;
  assign n4796 = n4764 & ~n4794;
  assign n4797 = ~n4795 & ~n4796;
  assign n4798 = ~n306 & ~n325;
  assign n4799 = ~n356 & ~n436;
  assign n4800 = ~n481 & n4799;
  assign n4801 = n4798 & n4800;
  assign n4802 = ~n125 & ~n140;
  assign n4803 = ~n199 & ~n226;
  assign n4804 = ~n428 & n4803;
  assign n4805 = n409 & n4802;
  assign n4806 = n813 & n991;
  assign n4807 = n4805 & n4806;
  assign n4808 = n3739 & n4804;
  assign n4809 = n4807 & n4808;
  assign n4810 = n4801 & n4809;
  assign n4811 = n972 & n4810;
  assign n4812 = n1984 & n3469;
  assign n4813 = n4811 & n4812;
  assign n4814 = n4797 & ~n4813;
  assign n4815 = ~n4797 & n4813;
  assign n4816 = ~n4814 & ~n4815;
  assign n4817 = ~n4763 & n4816;
  assign n4818 = n4763 & ~n4816;
  assign n4819 = ~n4817 & ~n4818;
  assign n4820 = ~n4756 & ~n4819;
  assign n4821 = n4756 & n4819;
  assign n4822 = ~n4820 & ~n4821;
  assign n4823 = ~n4757 & n4758;
  assign n4824 = n3761 & ~n4823;
  assign n4825 = n4822 & ~n4824;
  assign n4826 = ~n4822 & n4824;
  assign po13  = n4825 | n4826;
  assign n4828 = ~n4814 & ~n4817;
  assign n4829 = ~n4792 & ~n4795;
  assign n4830 = ~n4786 & ~n4789;
  assign n4831 = n2556 & ~n3842;
  assign n4832 = n2689 & ~n3514;
  assign n4833 = n2561 & n3647;
  assign n4834 = ~n4832 & ~n4833;
  assign n4835 = ~n4831 & n4834;
  assign n4836 = n604 & n4835;
  assign n4837 = ~n604 & ~n4835;
  assign n4838 = ~n4836 & ~n4837;
  assign n4839 = ~n604 & ~n3369;
  assign n4840 = ~n4779 & ~n4783;
  assign n4841 = ~n4839 & ~n4840;
  assign n4842 = n4839 & n4840;
  assign n4843 = ~n4841 & ~n4842;
  assign n4844 = n4838 & n4843;
  assign n4845 = ~n4838 & ~n4843;
  assign n4846 = ~n4844 & ~n4845;
  assign n4847 = ~n4830 & n4846;
  assign n4848 = n4830 & ~n4846;
  assign n4849 = ~n4847 & ~n4848;
  assign n4850 = ~n4829 & n4849;
  assign n4851 = n4829 & ~n4849;
  assign n4852 = ~n4850 & ~n4851;
  assign n4853 = ~n147 & ~n198;
  assign n4854 = ~n268 & ~n303;
  assign n4855 = ~n428 & n4854;
  assign n4856 = n265 & n4853;
  assign n4857 = n522 & n2146;
  assign n4858 = n2211 & n3024;
  assign n4859 = n4857 & n4858;
  assign n4860 = n4855 & n4856;
  assign n4861 = n4859 & n4860;
  assign n4862 = n816 & n4861;
  assign n4863 = n838 & n1306;
  assign n4864 = n4862 & n4863;
  assign n4865 = n1972 & n4864;
  assign n4866 = ~n4852 & n4865;
  assign n4867 = n4852 & ~n4865;
  assign n4868 = ~n4866 & ~n4867;
  assign n4869 = ~n4828 & n4868;
  assign n4870 = n4828 & ~n4868;
  assign n4871 = ~n4869 & ~n4870;
  assign n4872 = ~n4821 & ~n4871;
  assign n4873 = n4821 & n4871;
  assign n4874 = ~n4872 & ~n4873;
  assign n4875 = ~n4822 & n4823;
  assign n4876 = n3761 & ~n4875;
  assign n4877 = n4874 & ~n4876;
  assign n4878 = ~n4874 & n4876;
  assign po14  = n4877 | n4878;
  assign n4880 = ~n4867 & ~n4869;
  assign n4881 = ~n4841 & ~n4844;
  assign n4882 = n2556 & ~n3889;
  assign n4883 = ~n2689 & ~n4882;
  assign n4884 = n3647 & ~n4883;
  assign n4885 = n604 & n4884;
  assign n4886 = ~n604 & ~n4884;
  assign n4887 = ~n4885 & ~n4886;
  assign n4888 = ~n604 & n3521;
  assign n4889 = ~n4887 & ~n4888;
  assign n4890 = n4884 & n4888;
  assign n4891 = ~n4889 & ~n4890;
  assign n4892 = n4881 & ~n4891;
  assign n4893 = ~n4881 & n4891;
  assign n4894 = ~n4892 & ~n4893;
  assign n4895 = ~n4847 & ~n4850;
  assign n4896 = ~n4894 & n4895;
  assign n4897 = n4894 & ~n4895;
  assign n4898 = ~n4896 & ~n4897;
  assign n4899 = ~n176 & ~n200;
  assign n4900 = ~n262 & n4899;
  assign n4901 = n1005 & n4900;
  assign n4902 = ~n182 & ~n263;
  assign n4903 = ~n299 & ~n311;
  assign n4904 = n4902 & n4903;
  assign n4905 = n622 & n839;
  assign n4906 = n3431 & n4905;
  assign n4907 = n4904 & n4906;
  assign n4908 = n4741 & n4907;
  assign n4909 = n964 & n4908;
  assign n4910 = n2153 & n4909;
  assign n4911 = n4901 & n4910;
  assign n4912 = n4898 & ~n4911;
  assign n4913 = ~n4898 & n4911;
  assign n4914 = ~n4912 & ~n4913;
  assign n4915 = ~n4880 & n4914;
  assign n4916 = n4880 & ~n4914;
  assign n4917 = ~n4915 & ~n4916;
  assign n4918 = ~n4873 & ~n4917;
  assign n4919 = n4873 & n4917;
  assign n4920 = ~n4918 & ~n4919;
  assign n4921 = ~n4874 & n4875;
  assign n4922 = n3761 & ~n4921;
  assign n4923 = n4920 & ~n4922;
  assign n4924 = ~n4920 & n4922;
  assign po15  = n4923 | n4924;
  assign n4926 = ~n4912 & ~n4915;
  assign n4927 = ~n241 & ~n298;
  assign n4928 = ~n461 & n4927;
  assign n4929 = n183 & n640;
  assign n4930 = n4928 & n4929;
  assign n4931 = n2043 & n4930;
  assign n4932 = n3402 & n4801;
  assign n4933 = n4931 & n4932;
  assign n4934 = n3472 & n4933;
  assign n4935 = n2094 & n4934;
  assign n4936 = ~n604 & ~n3511;
  assign n4937 = n3369 & n4936;
  assign n4938 = ~n4889 & ~n4937;
  assign n4939 = ~n4893 & ~n4897;
  assign n4940 = ~n3369 & ~n3647;
  assign n4941 = n3369 & ~n3644;
  assign n4942 = ~n604 & ~n4941;
  assign n4943 = ~n4940 & n4942;
  assign n4944 = n4939 & ~n4943;
  assign n4945 = ~n4939 & n4943;
  assign n4946 = ~n4944 & ~n4945;
  assign n4947 = n4938 & n4946;
  assign n4948 = ~n4938 & ~n4946;
  assign n4949 = ~n4947 & ~n4948;
  assign n4950 = ~n4935 & n4949;
  assign n4951 = n4935 & ~n4949;
  assign n4952 = ~n4950 & ~n4951;
  assign n4953 = n4926 & n4952;
  assign n4954 = ~n4926 & ~n4952;
  assign n4955 = ~n4953 & ~n4954;
  assign n4956 = ~n4919 & n4955;
  assign n4957 = n4919 & ~n4955;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = ~n4920 & n4921;
  assign n4960 = n3761 & ~n4959;
  assign n4961 = n4958 & ~n4960;
  assign n4962 = ~n4958 & n4960;
  assign po16  = n4961 | n4962;
  assign n4964 = ~n4958 & n4959;
  assign n4965 = n3761 & ~n4964;
  assign n4966 = n4926 & ~n4950;
  assign n4967 = ~n4951 & ~n4966;
  assign n4968 = ~n208 & ~n210;
  assign n4969 = ~n457 & n4968;
  assign n4970 = n749 & n813;
  assign n4971 = n1007 & n2324;
  assign n4972 = n4970 & n4971;
  assign n4973 = n253 & n4969;
  assign n4974 = n4972 & n4973;
  assign n4975 = n411 & n4974;
  assign n4976 = n397 & n4975;
  assign n4977 = n2997 & n4976;
  assign n4978 = n4967 & ~n4977;
  assign n4979 = ~n4967 & n4977;
  assign n4980 = ~n4978 & ~n4979;
  assign n4981 = n4957 & n4980;
  assign n4982 = ~n4957 & ~n4980;
  assign n4983 = ~n4981 & ~n4982;
  assign n4984 = n4965 & n4983;
  assign n4985 = ~n4965 & ~n4983;
  assign po17  = ~n4984 & ~n4985;
  assign n4987 = n4964 & ~n4983;
  assign n4988 = n3761 & ~n4987;
  assign n4989 = ~n4978 & ~n4981;
  assign n4990 = ~n185 & ~n268;
  assign n4991 = ~n309 & ~n314;
  assign n4992 = ~n457 & n4991;
  assign n4993 = n4990 & n4992;
  assign n4994 = n625 & n819;
  assign n4995 = n4993 & n4994;
  assign n4996 = n976 & n1976;
  assign n4997 = n4995 & n4996;
  assign n4998 = n1014 & n4997;
  assign n4999 = n3449 & n4998;
  assign n5000 = n423 & n4999;
  assign n5001 = ~n4989 & n5000;
  assign n5002 = n4989 & ~n5000;
  assign n5003 = ~n5001 & ~n5002;
  assign n5004 = n4988 & n5003;
  assign n5005 = ~n4988 & ~n5003;
  assign po18  = n5004 | n5005;
  assign n5007 = n4978 & ~n5000;
  assign n5008 = ~n145 & ~n209;
  assign n5009 = ~n304 & ~n327;
  assign n5010 = ~n412 & ~n461;
  assign n5011 = ~n546 & n5010;
  assign n5012 = n5008 & n5009;
  assign n5013 = n615 & n5012;
  assign n5014 = n4171 & n5011;
  assign n5015 = n5013 & n5014;
  assign n5016 = n2891 & n5015;
  assign n5017 = n796 & n5016;
  assign n5018 = n4901 & n5017;
  assign n5019 = ~n5007 & n5018;
  assign n5020 = n5007 & ~n5018;
  assign n5021 = ~n5019 & ~n5020;
  assign n5022 = n4981 & ~n5000;
  assign n5023 = ~n5021 & ~n5022;
  assign n5024 = n5021 & n5022;
  assign n5025 = ~n5023 & ~n5024;
  assign n5026 = n4987 & n5003;
  assign n5027 = n3761 & ~n5026;
  assign n5028 = n5025 & ~n5027;
  assign n5029 = ~n5025 & n5027;
  assign po19  = n5028 | n5029;
  assign n5031 = ~n5025 & n5026;
  assign n5032 = n3761 & ~n5031;
  assign n5033 = ~n5020 & ~n5024;
  assign n5034 = ~n378 & n470;
  assign n5035 = n545 & n3397;
  assign n5036 = n4368 & n5035;
  assign n5037 = n4172 & n5034;
  assign n5038 = n5036 & n5037;
  assign n5039 = n578 & n5038;
  assign n5040 = n831 & n5039;
  assign n5041 = n4457 & n5040;
  assign n5042 = ~n5033 & n5041;
  assign n5043 = n5033 & ~n5041;
  assign n5044 = ~n5042 & ~n5043;
  assign n5045 = n5032 & n5044;
  assign n5046 = ~n5032 & ~n5044;
  assign po20  = n5045 | n5046;
  assign n5048 = n5020 & ~n5041;
  assign n5049 = ~n427 & n532;
  assign n5050 = n3360 & n5049;
  assign n5051 = n504 & n5050;
  assign n5052 = ~n5048 & n5051;
  assign n5053 = n5048 & ~n5051;
  assign n5054 = ~n5052 & ~n5053;
  assign n5055 = n5024 & ~n5041;
  assign n5056 = ~n5054 & ~n5055;
  assign n5057 = n5054 & n5055;
  assign n5058 = ~n5056 & ~n5057;
  assign n5059 = n5031 & n5044;
  assign n5060 = n3761 & ~n5059;
  assign n5061 = n5058 & ~n5060;
  assign n5062 = ~n5058 & n5060;
  assign po21  = n5061 | n5062;
  assign n5064 = ~n5058 & n5059;
  assign n5065 = n3761 & ~n5064;
  assign n5066 = n504 & n570;
  assign n5067 = ~n5053 & ~n5057;
  assign n5068 = ~n5066 & ~n5067;
  assign n5069 = n5066 & n5067;
  assign n5070 = ~n5068 & ~n5069;
  assign n5071 = ~n5065 & n5070;
  assign n5072 = n5065 & ~n5070;
  assign po22  = n5071 | n5072;
  assign n5074 = n5064 & ~n5070;
  assign n5075 = n3761 & ~n5074;
  assign n5076 = n5053 & n5057;
  assign n5077 = n5068 & ~n5076;
  assign n5078 = ~n5075 & n5077;
  assign n5079 = n98 & n103;
  assign n5080 = n5075 & ~n5077;
  assign n5081 = ~n5078 & ~n5079;
  assign po23  = n5080 | ~n5081;
  assign n5083 = ~n5066 & n5076;
  assign n5084 = ~n5074 & ~n5083;
  assign n5085 = n5064 & n5068;
  assign n5086 = ~n5079 & ~n5085;
  assign n5087 = ~n5084 & n5086;
  assign po24  = n3761 & ~n5087;
endmodule
