module mem_ctrl ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17,
    pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26,
    pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44,
    pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53,
    pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62,
    pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80,
    pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107,
    pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116,
    pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125,
    pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134,
    pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143,
    pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152,
    pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161,
    pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170,
    pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197,
    pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206,
    pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215,
    pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224,
    pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233,
    pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242,
    pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251,
    pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260,
    pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287,
    pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296,
    pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305,
    pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314,
    pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323,
    pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332,
    pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341,
    pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350,
    pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377,
    pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386,
    pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395,
    pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404,
    pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413,
    pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422,
    pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431,
    pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440,
    pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467,
    pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476,
    pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485,
    pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494,
    pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503,
    pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, pi512,
    pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520, pi521,
    pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529, pi530,
    pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539,
    pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548,
    pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557,
    pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566,
    pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574, pi575,
    pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583, pi584,
    pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592, pi593,
    pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601, pi602,
    pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610, pi611,
    pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619, pi620,
    pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629,
    pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638,
    pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647,
    pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656,
    pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664, pi665,
    pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673, pi674,
    pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682, pi683,
    pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691, pi692,
    pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700, pi701,
    pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709, pi710,
    pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719,
    pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728,
    pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737,
    pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746,
    pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754, pi755,
    pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763, pi764,
    pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772, pi773,
    pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781, pi782,
    pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790, pi791,
    pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799, pi800,
    pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808, pi809,
    pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818,
    pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827,
    pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835, pi836,
    pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844, pi845,
    pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853, pi854,
    pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862, pi863,
    pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871, pi872,
    pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880, pi881,
    pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889, pi890,
    pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898, pi899,
    pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907, pi908,
    pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916, pi917,
    pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925, pi926,
    pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934, pi935,
    pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943, pi944,
    pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952, pi953,
    pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961, pi962,
    pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970, pi971,
    pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979, pi980,
    pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988, pi989,
    pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997, pi998,
    pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0, po1, po2, po3, po4, po5, po6, po7, po8,
    po9, po10, po11, po12, po13, po14, po15, po16, po17,
    po18, po19, po20, po21, po22, po23, po24, po25, po26,
    po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44,
    po45, po46, po47, po48, po49, po50, po51, po52, po53,
    po54, po55, po56, po57, po58, po59, po60, po61, po62,
    po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80,
    po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98,
    po99, po100, po101, po102, po103, po104, po105, po106, po107,
    po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125,
    po126, po127, po128, po129, po130, po131, po132, po133, po134,
    po135, po136, po137, po138, po139, po140, po141, po142, po143,
    po144, po145, po146, po147, po148, po149, po150, po151, po152,
    po153, po154, po155, po156, po157, po158, po159, po160, po161,
    po162, po163, po164, po165, po166, po167, po168, po169, po170,
    po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188,
    po189, po190, po191, po192, po193, po194, po195, po196, po197,
    po198, po199, po200, po201, po202, po203, po204, po205, po206,
    po207, po208, po209, po210, po211, po212, po213, po214, po215,
    po216, po217, po218, po219, po220, po221, po222, po223, po224,
    po225, po226, po227, po228, po229, po230, po231, po232, po233,
    po234, po235, po236, po237, po238, po239, po240, po241, po242,
    po243, po244, po245, po246, po247, po248, po249, po250, po251,
    po252, po253, po254, po255, po256, po257, po258, po259, po260,
    po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278,
    po279, po280, po281, po282, po283, po284, po285, po286, po287,
    po288, po289, po290, po291, po292, po293, po294, po295, po296,
    po297, po298, po299, po300, po301, po302, po303, po304, po305,
    po306, po307, po308, po309, po310, po311, po312, po313, po314,
    po315, po316, po317, po318, po319, po320, po321, po322, po323,
    po324, po325, po326, po327, po328, po329, po330, po331, po332,
    po333, po334, po335, po336, po337, po338, po339, po340, po341,
    po342, po343, po344, po345, po346, po347, po348, po349, po350,
    po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368,
    po369, po370, po371, po372, po373, po374, po375, po376, po377,
    po378, po379, po380, po381, po382, po383, po384, po385, po386,
    po387, po388, po389, po390, po391, po392, po393, po394, po395,
    po396, po397, po398, po399, po400, po401, po402, po403, po404,
    po405, po406, po407, po408, po409, po410, po411, po412, po413,
    po414, po415, po416, po417, po418, po419, po420, po421, po422,
    po423, po424, po425, po426, po427, po428, po429, po430, po431,
    po432, po433, po434, po435, po436, po437, po438, po439, po440,
    po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458,
    po459, po460, po461, po462, po463, po464, po465, po466, po467,
    po468, po469, po470, po471, po472, po473, po474, po475, po476,
    po477, po478, po479, po480, po481, po482, po483, po484, po485,
    po486, po487, po488, po489, po490, po491, po492, po493, po494,
    po495, po496, po497, po498, po499, po500, po501, po502, po503,
    po504, po505, po506, po507, po508, po509, po510, po511, po512,
    po513, po514, po515, po516, po517, po518, po519, po520, po521,
    po522, po523, po524, po525, po526, po527, po528, po529, po530,
    po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548,
    po549, po550, po551, po552, po553, po554, po555, po556, po557,
    po558, po559, po560, po561, po562, po563, po564, po565, po566,
    po567, po568, po569, po570, po571, po572, po573, po574, po575,
    po576, po577, po578, po579, po580, po581, po582, po583, po584,
    po585, po586, po587, po588, po589, po590, po591, po592, po593,
    po594, po595, po596, po597, po598, po599, po600, po601, po602,
    po603, po604, po605, po606, po607, po608, po609, po610, po611,
    po612, po613, po614, po615, po616, po617, po618, po619, po620,
    po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638,
    po639, po640, po641, po642, po643, po644, po645, po646, po647,
    po648, po649, po650, po651, po652, po653, po654, po655, po656,
    po657, po658, po659, po660, po661, po662, po663, po664, po665,
    po666, po667, po668, po669, po670, po671, po672, po673, po674,
    po675, po676, po677, po678, po679, po680, po681, po682, po683,
    po684, po685, po686, po687, po688, po689, po690, po691, po692,
    po693, po694, po695, po696, po697, po698, po699, po700, po701,
    po702, po703, po704, po705, po706, po707, po708, po709, po710,
    po711, po712, po713, po714, po715, po716, po717, po718, po719,
    po720, po721, po722, po723, po724, po725, po726, po727, po728,
    po729, po730, po731, po732, po733, po734, po735, po736, po737,
    po738, po739, po740, po741, po742, po743, po744, po745, po746,
    po747, po748, po749, po750, po751, po752, po753, po754, po755,
    po756, po757, po758, po759, po760, po761, po762, po763, po764,
    po765, po766, po767, po768, po769, po770, po771, po772, po773,
    po774, po775, po776, po777, po778, po779, po780, po781, po782,
    po783, po784, po785, po786, po787, po788, po789, po790, po791,
    po792, po793, po794, po795, po796, po797, po798, po799, po800,
    po801, po802, po803, po804, po805, po806, po807, po808, po809,
    po810, po811, po812, po813, po814, po815, po816, po817, po818,
    po819, po820, po821, po822, po823, po824, po825, po826, po827,
    po828, po829, po830, po831, po832, po833, po834, po835, po836,
    po837, po838, po839, po840, po841, po842, po843, po844, po845,
    po846, po847, po848, po849, po850, po851, po852, po853, po854,
    po855, po856, po857, po858, po859, po860, po861, po862, po863,
    po864, po865, po866, po867, po868, po869, po870, po871, po872,
    po873, po874, po875, po876, po877, po878, po879, po880, po881,
    po882, po883, po884, po885, po886, po887, po888, po889, po890,
    po891, po892, po893, po894, po895, po896, po897, po898, po899,
    po900, po901, po902, po903, po904, po905, po906, po907, po908,
    po909, po910, po911, po912, po913, po914, po915, po916, po917,
    po918, po919, po920, po921, po922, po923, po924, po925, po926,
    po927, po928, po929, po930, po931, po932, po933, po934, po935,
    po936, po937, po938, po939, po940, po941, po942, po943, po944,
    po945, po946, po947, po948, po949, po950, po951, po952, po953,
    po954, po955, po956, po957, po958, po959, po960, po961, po962,
    po963, po964, po965, po966, po967, po968, po969, po970, po971,
    po972, po973, po974, po975, po976, po977, po978, po979, po980,
    po981, po982, po983, po984, po985, po986, po987, po988, po989,
    po990, po991, po992, po993, po994, po995, po996, po997, po998,
    po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7,
    pi8, pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16,
    pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25,
    pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34,
    pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43,
    pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52,
    pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61,
    pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70,
    pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97,
    pi98, pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106,
    pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115,
    pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124,
    pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133,
    pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142,
    pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151,
    pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160,
    pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187,
    pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196,
    pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205,
    pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214,
    pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223,
    pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232,
    pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241,
    pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250,
    pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277,
    pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286,
    pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295,
    pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304,
    pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313,
    pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322,
    pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331,
    pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340,
    pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367,
    pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376,
    pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385,
    pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394,
    pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403,
    pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412,
    pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421,
    pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430,
    pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457,
    pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466,
    pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475,
    pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484,
    pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493,
    pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502,
    pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511,
    pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520,
    pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529,
    pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538,
    pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547,
    pi548, pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556,
    pi557, pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565,
    pi566, pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574,
    pi575, pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583,
    pi584, pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592,
    pi593, pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601,
    pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610,
    pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619,
    pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628,
    pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637,
    pi638, pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646,
    pi647, pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655,
    pi656, pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664,
    pi665, pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673,
    pi674, pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682,
    pi683, pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691,
    pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700,
    pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709,
    pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718,
    pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727,
    pi728, pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736,
    pi737, pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745,
    pi746, pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754,
    pi755, pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763,
    pi764, pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772,
    pi773, pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781,
    pi782, pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790,
    pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799,
    pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808,
    pi809, pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817,
    pi818, pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826,
    pi827, pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835,
    pi836, pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844,
    pi845, pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853,
    pi854, pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862,
    pi863, pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871,
    pi872, pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880,
    pi881, pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889,
    pi890, pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898,
    pi899, pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907,
    pi908, pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916,
    pi917, pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925,
    pi926, pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934,
    pi935, pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943,
    pi944, pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952,
    pi953, pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961,
    pi962, pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970,
    pi971, pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979,
    pi980, pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988,
    pi989, pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997,
    pi998, pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0, po1, po2, po3, po4, po5, po6, po7,
    po8, po9, po10, po11, po12, po13, po14, po15, po16,
    po17, po18, po19, po20, po21, po22, po23, po24, po25,
    po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43,
    po44, po45, po46, po47, po48, po49, po50, po51, po52,
    po53, po54, po55, po56, po57, po58, po59, po60, po61,
    po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88,
    po89, po90, po91, po92, po93, po94, po95, po96, po97,
    po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115,
    po116, po117, po118, po119, po120, po121, po122, po123, po124,
    po125, po126, po127, po128, po129, po130, po131, po132, po133,
    po134, po135, po136, po137, po138, po139, po140, po141, po142,
    po143, po144, po145, po146, po147, po148, po149, po150, po151,
    po152, po153, po154, po155, po156, po157, po158, po159, po160,
    po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178,
    po179, po180, po181, po182, po183, po184, po185, po186, po187,
    po188, po189, po190, po191, po192, po193, po194, po195, po196,
    po197, po198, po199, po200, po201, po202, po203, po204, po205,
    po206, po207, po208, po209, po210, po211, po212, po213, po214,
    po215, po216, po217, po218, po219, po220, po221, po222, po223,
    po224, po225, po226, po227, po228, po229, po230, po231, po232,
    po233, po234, po235, po236, po237, po238, po239, po240, po241,
    po242, po243, po244, po245, po246, po247, po248, po249, po250,
    po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268,
    po269, po270, po271, po272, po273, po274, po275, po276, po277,
    po278, po279, po280, po281, po282, po283, po284, po285, po286,
    po287, po288, po289, po290, po291, po292, po293, po294, po295,
    po296, po297, po298, po299, po300, po301, po302, po303, po304,
    po305, po306, po307, po308, po309, po310, po311, po312, po313,
    po314, po315, po316, po317, po318, po319, po320, po321, po322,
    po323, po324, po325, po326, po327, po328, po329, po330, po331,
    po332, po333, po334, po335, po336, po337, po338, po339, po340,
    po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358,
    po359, po360, po361, po362, po363, po364, po365, po366, po367,
    po368, po369, po370, po371, po372, po373, po374, po375, po376,
    po377, po378, po379, po380, po381, po382, po383, po384, po385,
    po386, po387, po388, po389, po390, po391, po392, po393, po394,
    po395, po396, po397, po398, po399, po400, po401, po402, po403,
    po404, po405, po406, po407, po408, po409, po410, po411, po412,
    po413, po414, po415, po416, po417, po418, po419, po420, po421,
    po422, po423, po424, po425, po426, po427, po428, po429, po430,
    po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448,
    po449, po450, po451, po452, po453, po454, po455, po456, po457,
    po458, po459, po460, po461, po462, po463, po464, po465, po466,
    po467, po468, po469, po470, po471, po472, po473, po474, po475,
    po476, po477, po478, po479, po480, po481, po482, po483, po484,
    po485, po486, po487, po488, po489, po490, po491, po492, po493,
    po494, po495, po496, po497, po498, po499, po500, po501, po502,
    po503, po504, po505, po506, po507, po508, po509, po510, po511,
    po512, po513, po514, po515, po516, po517, po518, po519, po520,
    po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538,
    po539, po540, po541, po542, po543, po544, po545, po546, po547,
    po548, po549, po550, po551, po552, po553, po554, po555, po556,
    po557, po558, po559, po560, po561, po562, po563, po564, po565,
    po566, po567, po568, po569, po570, po571, po572, po573, po574,
    po575, po576, po577, po578, po579, po580, po581, po582, po583,
    po584, po585, po586, po587, po588, po589, po590, po591, po592,
    po593, po594, po595, po596, po597, po598, po599, po600, po601,
    po602, po603, po604, po605, po606, po607, po608, po609, po610,
    po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628,
    po629, po630, po631, po632, po633, po634, po635, po636, po637,
    po638, po639, po640, po641, po642, po643, po644, po645, po646,
    po647, po648, po649, po650, po651, po652, po653, po654, po655,
    po656, po657, po658, po659, po660, po661, po662, po663, po664,
    po665, po666, po667, po668, po669, po670, po671, po672, po673,
    po674, po675, po676, po677, po678, po679, po680, po681, po682,
    po683, po684, po685, po686, po687, po688, po689, po690, po691,
    po692, po693, po694, po695, po696, po697, po698, po699, po700,
    po701, po702, po703, po704, po705, po706, po707, po708, po709,
    po710, po711, po712, po713, po714, po715, po716, po717, po718,
    po719, po720, po721, po722, po723, po724, po725, po726, po727,
    po728, po729, po730, po731, po732, po733, po734, po735, po736,
    po737, po738, po739, po740, po741, po742, po743, po744, po745,
    po746, po747, po748, po749, po750, po751, po752, po753, po754,
    po755, po756, po757, po758, po759, po760, po761, po762, po763,
    po764, po765, po766, po767, po768, po769, po770, po771, po772,
    po773, po774, po775, po776, po777, po778, po779, po780, po781,
    po782, po783, po784, po785, po786, po787, po788, po789, po790,
    po791, po792, po793, po794, po795, po796, po797, po798, po799,
    po800, po801, po802, po803, po804, po805, po806, po807, po808,
    po809, po810, po811, po812, po813, po814, po815, po816, po817,
    po818, po819, po820, po821, po822, po823, po824, po825, po826,
    po827, po828, po829, po830, po831, po832, po833, po834, po835,
    po836, po837, po838, po839, po840, po841, po842, po843, po844,
    po845, po846, po847, po848, po849, po850, po851, po852, po853,
    po854, po855, po856, po857, po858, po859, po860, po861, po862,
    po863, po864, po865, po866, po867, po868, po869, po870, po871,
    po872, po873, po874, po875, po876, po877, po878, po879, po880,
    po881, po882, po883, po884, po885, po886, po887, po888, po889,
    po890, po891, po892, po893, po894, po895, po896, po897, po898,
    po899, po900, po901, po902, po903, po904, po905, po906, po907,
    po908, po909, po910, po911, po912, po913, po914, po915, po916,
    po917, po918, po919, po920, po921, po922, po923, po924, po925,
    po926, po927, po928, po929, po930, po931, po932, po933, po934,
    po935, po936, po937, po938, po939, po940, po941, po942, po943,
    po944, po945, po946, po947, po948, po949, po950, po951, po952,
    po953, po954, po955, po956, po957, po958, po959, po960, po961,
    po962, po963, po964, po965, po966, po967, po968, po969, po970,
    po971, po972, po973, po974, po975, po976, po977, po978, po979,
    po980, po981, po982, po983, po984, po985, po986, po987, po988,
    po989, po990, po991, po992, po993, po994, po995, po996, po997,
    po998, po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904,
    n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282,
    n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300,
    n3301, n3302, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686,
    n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927,
    n3928, n3930, n3931, n3932, n3933, n3934,
    n3935, n3936, n3937, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006,
    n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036,
    n4037, n4038, n4039, n4040, n4041, n4042,
    n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072,
    n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114,
    n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144,
    n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4157,
    n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181,
    n4182, n4183, n4184, n4185, n4186, n4187,
    n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217,
    n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235,
    n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4243, n4244, n4245, n4246, n4247,
    n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277,
    n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307,
    n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331,
    n4332, n4333, n4334, n4335, n4336, n4337,
    n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367,
    n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392,
    n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422,
    n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476,
    n4477, n4478, n4479, n4480, n4481, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596,
    n4597, n4598, n4599, n4600, n4601, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747,
    n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036,
    n5037, n5038, n5039, n5040, n5041, n5042,
    n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061,
    n5062, n5063, n5064, n5065, n5066, n5067,
    n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151,
    n5152, n5153, n5154, n5155, n5156, n5157,
    n5158, n5159, n5160, n5161, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181,
    n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211,
    n5212, n5213, n5214, n5215, n5216, n5217,
    n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241,
    n5242, n5243, n5244, n5245, n5246, n5247,
    n5248, n5249, n5250, n5251, n5252, n5253,
    n5254, n5255, n5256, n5257, n5258, n5259,
    n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271,
    n5272, n5273, n5274, n5276, n5277, n5278,
    n5279, n5280, n5281, n5282, n5283, n5284,
    n5285, n5286, n5287, n5288, n5289, n5290,
    n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302,
    n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314,
    n5315, n5316, n5317, n5318, n5319, n5320,
    n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332,
    n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5344,
    n5345, n5346, n5347, n5348, n5349, n5350,
    n5351, n5352, n5353, n5354, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362,
    n5363, n5364, n5365, n5366, n5367, n5368,
    n5369, n5370, n5371, n5372, n5373, n5374,
    n5375, n5376, n5377, n5378, n5379, n5380,
    n5381, n5382, n5383, n5384, n5385, n5386,
    n5387, n5388, n5389, n5390, n5391, n5392,
    n5393, n5394, n5395, n5396, n5397, n5398,
    n5399, n5400, n5401, n5402, n5403, n5404,
    n5405, n5406, n5407, n5408, n5409, n5410,
    n5411, n5412, n5413, n5414, n5415, n5416,
    n5417, n5418, n5419, n5420, n5421, n5422,
    n5423, n5424, n5425, n5426, n5427, n5428,
    n5429, n5430, n5431, n5432, n5433, n5434,
    n5435, n5436, n5437, n5438, n5439, n5440,
    n5441, n5442, n5443, n5444, n5445, n5446,
    n5447, n5448, n5449, n5450, n5451, n5452,
    n5453, n5454, n5455, n5456, n5457, n5458,
    n5459, n5460, n5461, n5462, n5463, n5464,
    n5465, n5466, n5467, n5468, n5469, n5470,
    n5471, n5472, n5473, n5474, n5475, n5476,
    n5477, n5478, n5479, n5480, n5481, n5482,
    n5483, n5484, n5485, n5486, n5487, n5488,
    n5489, n5490, n5491, n5492, n5493, n5494,
    n5495, n5496, n5497, n5498, n5499, n5500,
    n5501, n5502, n5503, n5504, n5505, n5506,
    n5507, n5508, n5510, n5511, n5512, n5513,
    n5514, n5515, n5516, n5517, n5518, n5519,
    n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531,
    n5532, n5533, n5534, n5535, n5536, n5537,
    n5538, n5539, n5540, n5541, n5542, n5543,
    n5544, n5545, n5546, n5547, n5548, n5549,
    n5550, n5551, n5552, n5553, n5554, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561,
    n5562, n5563, n5564, n5565, n5566, n5567,
    n5568, n5569, n5570, n5571, n5572, n5573,
    n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591,
    n5592, n5593, n5594, n5595, n5596, n5597,
    n5598, n5599, n5600, n5601, n5602, n5603,
    n5604, n5605, n5606, n5607, n5608, n5609,
    n5610, n5611, n5612, n5613, n5614, n5615,
    n5616, n5617, n5618, n5619, n5620, n5621,
    n5622, n5623, n5624, n5625, n5626, n5627,
    n5628, n5629, n5630, n5631, n5632, n5633,
    n5634, n5635, n5636, n5637, n5638, n5639,
    n5640, n5641, n5642, n5643, n5644, n5645,
    n5646, n5647, n5648, n5649, n5650, n5651,
    n5652, n5653, n5654, n5655, n5656, n5657,
    n5658, n5659, n5660, n5661, n5662, n5663,
    n5664, n5665, n5666, n5667, n5668, n5669,
    n5670, n5671, n5672, n5673, n5674, n5675,
    n5676, n5677, n5678, n5679, n5680, n5681,
    n5682, n5683, n5684, n5685, n5686, n5687,
    n5688, n5689, n5690, n5691, n5692, n5693,
    n5694, n5695, n5696, n5697, n5698, n5699,
    n5700, n5701, n5702, n5703, n5704, n5705,
    n5706, n5707, n5708, n5709, n5710, n5711,
    n5712, n5713, n5714, n5715, n5716, n5717,
    n5718, n5719, n5720, n5721, n5722, n5723,
    n5724, n5725, n5726, n5727, n5728, n5729,
    n5730, n5731, n5732, n5733, n5734, n5735,
    n5736, n5737, n5738, n5739, n5740, n5741,
    n5742, n5744, n5745, n5746, n5747, n5748,
    n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760,
    n5761, n5762, n5763, n5764, n5765, n5766,
    n5767, n5768, n5769, n5770, n5771, n5772,
    n5773, n5774, n5775, n5776, n5777, n5778,
    n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790,
    n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802,
    n5803, n5804, n5805, n5806, n5807, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814,
    n5815, n5816, n5817, n5818, n5819, n5820,
    n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5830, n5831, n5832,
    n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844,
    n5845, n5846, n5847, n5848, n5849, n5850,
    n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874,
    n5875, n5876, n5877, n5878, n5879, n5880,
    n5881, n5882, n5883, n5884, n5885, n5886,
    n5887, n5888, n5889, n5890, n5891, n5892,
    n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904,
    n5905, n5906, n5907, n5908, n5909, n5910,
    n5911, n5912, n5913, n5914, n5915, n5916,
    n5917, n5918, n5919, n5920, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934,
    n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946,
    n5947, n5948, n5949, n5950, n5951, n5952,
    n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964,
    n5965, n5966, n5967, n5968, n5969, n5970,
    n5971, n5972, n5973, n5974, n5975, n5976,
    n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994,
    n5995, n5996, n5997, n5998, n5999, n6000,
    n6001, n6002, n6003, n6004, n6005, n6006,
    n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6022, n6023, n6024,
    n6025, n6026, n6027, n6028, n6029, n6030,
    n6031, n6032, n6033, n6034, n6035, n6036,
    n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060,
    n6061, n6062, n6063, n6064, n6065, n6066,
    n6067, n6068, n6069, n6070, n6071, n6072,
    n6073, n6074, n6075, n6076, n6077, n6078,
    n6079, n6080, n6081, n6082, n6083, n6084,
    n6085, n6086, n6087, n6088, n6089, n6090,
    n6091, n6092, n6093, n6094, n6095, n6097,
    n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6126, n6127,
    n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145,
    n6146, n6147, n6148, n6149, n6150, n6151,
    n6152, n6153, n6154, n6155, n6156, n6157,
    n6158, n6159, n6160, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170,
    n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236,
    n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6255,
    n6256, n6257, n6258, n6260, n6261, n6262,
    n6263, n6264, n6265, n6266, n6267, n6268,
    n6269, n6270, n6271, n6272, n6273, n6274,
    n6275, n6276, n6277, n6278, n6279, n6280,
    n6281, n6282, n6283, n6285, n6286, n6287,
    n6288, n6289, n6290, n6291, n6292, n6293,
    n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6302, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310, n6311,
    n6312, n6313, n6314, n6315, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372,
    n6373, n6374, n6375, n6376, n6377, n6378,
    n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462,
    n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546,
    n6547, n6548, n6549, n6550, n6551, n6552,
    n6554, n6555, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571,
    n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601,
    n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631,
    n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649,
    n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661,
    n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782,
    n6783, n6784, n6785, n6786, n6787, n6788,
    n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6804, n6805, n6806, n6807,
    n6808, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831,
    n6832, n6833, n6834, n6835, n6836, n6837,
    n6838, n6839, n6840, n6841, n6842, n6843,
    n6844, n6845, n6846, n6847, n6848, n6849,
    n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861,
    n6862, n6863, n6864, n6865, n6866, n6867,
    n6868, n6869, n6870, n6871, n6872, n6873,
    n6874, n6875, n6876, n6877, n6878, n6879,
    n6880, n6881, n6882, n6883, n6884, n6885,
    n6886, n6887, n6888, n6889, n6890, n6891,
    n6892, n6893, n6894, n6895, n6897, n6898,
    n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952,
    n6953, n6954, n6955, n6956, n6957, n6958,
    n6959, n6960, n6961, n6962, n6963, n6964,
    n6965, n6966, n6967, n6968, n6969, n6970,
    n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982,
    n6983, n6984, n6985, n6986, n6987, n6988,
    n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7001,
    n7002, n7003, n7004, n7005, n7006, n7007,
    n7008, n7009, n7010, n7011, n7012, n7013,
    n7014, n7015, n7016, n7017, n7018, n7019,
    n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031,
    n7032, n7033, n7034, n7035, n7036, n7037,
    n7038, n7039, n7040, n7041, n7042, n7043,
    n7044, n7045, n7046, n7047, n7048, n7049,
    n7050, n7051, n7052, n7053, n7054, n7055,
    n7056, n7057, n7058, n7059, n7060, n7061,
    n7062, n7063, n7064, n7065, n7066, n7067,
    n7068, n7069, n7070, n7071, n7072, n7073,
    n7074, n7075, n7076, n7077, n7078, n7079,
    n7080, n7081, n7083, n7084, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092,
    n7093, n7094, n7095, n7096, n7097, n7098,
    n7099, n7100, n7101, n7102, n7103, n7104,
    n7105, n7106, n7107, n7108, n7109, n7110,
    n7111, n7112, n7113, n7114, n7115, n7116,
    n7117, n7118, n7119, n7120, n7121, n7122,
    n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7133, n7134,
    n7135, n7136, n7137, n7138, n7139, n7140,
    n7141, n7142, n7143, n7144, n7145, n7146,
    n7147, n7148, n7149, n7150, n7151, n7152,
    n7153, n7154, n7155, n7156, n7157, n7158,
    n7159, n7160, n7161, n7162, n7163, n7164,
    n7165, n7166, n7167, n7168, n7169, n7170,
    n7171, n7172, n7173, n7174, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7194, n7195,
    n7196, n7197, n7198, n7199, n7200, n7201,
    n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7227, n7228, n7229, n7230, n7231,
    n7232, n7233, n7234, n7235, n7236, n7237,
    n7238, n7239, n7240, n7241, n7242, n7243,
    n7244, n7245, n7246, n7247, n7248, n7249,
    n7250, n7251, n7252, n7253, n7254, n7255,
    n7256, n7257, n7258, n7259, n7260, n7261,
    n7262, n7263, n7264, n7265, n7266, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7320, n7321, n7323, n7324,
    n7325, n7326, n7327, n7328, n7329, n7330,
    n7331, n7332, n7333, n7334, n7335, n7336,
    n7337, n7338, n7339, n7340, n7341, n7342,
    n7343, n7344, n7345, n7346, n7347, n7348,
    n7349, n7350, n7351, n7352, n7353, n7354,
    n7355, n7356, n7357, n7358, n7359, n7360,
    n7361, n7362, n7363, n7364, n7365, n7366,
    n7367, n7368, n7369, n7370, n7371, n7373,
    n7374, n7375, n7376, n7378, n7380, n7382,
    n7384, n7385, n7386, n7387, n7388, n7389,
    n7390, n7391, n7392, n7393, n7394, n7395,
    n7396, n7397, n7398, n7399, n7400, n7401,
    n7402, n7403, n7404, n7405, n7406, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431,
    n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443,
    n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7461,
    n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473,
    n7474, n7475, n7476, n7477, n7478, n7479,
    n7480, n7481, n7482, n7483, n7484, n7485,
    n7486, n7487, n7488, n7489, n7490, n7491,
    n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503,
    n7504, n7505, n7506, n7507, n7508, n7509,
    n7510, n7511, n7512, n7513, n7514, n7515,
    n7516, n7517, n7518, n7519, n7520, n7521,
    n7522, n7523, n7524, n7525, n7526, n7527,
    n7528, n7529, n7530, n7531, n7532, n7533,
    n7534, n7535, n7536, n7537, n7538, n7539,
    n7540, n7541, n7542, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551,
    n7552, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563,
    n7564, n7565, n7566, n7567, n7568, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581,
    n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611,
    n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653,
    n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683,
    n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713,
    n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7721, n7722, n7723, n7724, n7725,
    n7726, n7727, n7728, n7729, n7730, n7731,
    n7732, n7733, n7734, n7735, n7736, n7737,
    n7738, n7739, n7740, n7741, n7742, n7743,
    n7744, n7745, n7746, n7747, n7748, n7749,
    n7750, n7751, n7752, n7753, n7754, n7755,
    n7756, n7757, n7758, n7759, n7760, n7761,
    n7762, n7763, n7764, n7765, n7766, n7767,
    n7768, n7769, n7770, n7771, n7772, n7773,
    n7774, n7775, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785,
    n7786, n7787, n7788, n7789, n7790, n7791,
    n7792, n7793, n7794, n7795, n7796, n7797,
    n7798, n7799, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821,
    n7822, n7823, n7824, n7825, n7826, n7827,
    n7828, n7829, n7830, n7831, n7832, n7833,
    n7834, n7835, n7836, n7837, n7838, n7839,
    n7840, n7841, n7842, n7843, n7844, n7845,
    n7846, n7847, n7848, n7849, n7850, n7851,
    n7852, n7853, n7854, n7855, n7856, n7857,
    n7858, n7859, n7860, n7861, n7862, n7863,
    n7864, n7865, n7866, n7867, n7868, n7869,
    n7870, n7871, n7872, n7873, n7874, n7875,
    n7876, n7877, n7878, n7879, n7880, n7881,
    n7882, n7883, n7884, n7885, n7886, n7887,
    n7888, n7889, n7890, n7891, n7892, n7893,
    n7894, n7895, n7896, n7897, n7898, n7899,
    n7900, n7901, n7902, n7903, n7904, n7905,
    n7906, n7907, n7908, n7909, n7910, n7911,
    n7912, n7913, n7914, n7915, n7916, n7917,
    n7918, n7919, n7920, n7921, n7922, n7923,
    n7924, n7925, n7926, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935,
    n7936, n7937, n7938, n7939, n7940, n7941,
    n7942, n7943, n7944, n7945, n7946, n7947,
    n7948, n7949, n7950, n7951, n7952, n7953,
    n7954, n7955, n7956, n7957, n7958, n7959,
    n7960, n7961, n7962, n7963, n7964, n7965,
    n7966, n7967, n7968, n7969, n7970, n7971,
    n7972, n7973, n7974, n7975, n7976, n7977,
    n7978, n7979, n7980, n7981, n7982, n7983,
    n7984, n7985, n7986, n7987, n7988, n7989,
    n7990, n7991, n7992, n7993, n7994, n7995,
    n7996, n7997, n7998, n7999, n8000, n8001,
    n8002, n8003, n8004, n8005, n8006, n8007,
    n8008, n8009, n8010, n8011, n8012, n8013,
    n8014, n8015, n8016, n8017, n8018, n8019,
    n8020, n8021, n8022, n8023, n8024, n8025,
    n8026, n8027, n8028, n8029, n8030, n8031,
    n8032, n8033, n8034, n8035, n8036, n8037,
    n8038, n8039, n8040, n8041, n8042, n8043,
    n8044, n8045, n8046, n8047, n8048, n8049,
    n8050, n8051, n8052, n8053, n8054, n8055,
    n8056, n8057, n8058, n8059, n8060, n8061,
    n8062, n8063, n8064, n8065, n8066, n8067,
    n8068, n8069, n8070, n8071, n8072, n8073,
    n8074, n8075, n8076, n8077, n8078, n8079,
    n8080, n8081, n8082, n8083, n8084, n8085,
    n8086, n8087, n8088, n8089, n8090, n8091,
    n8092, n8093, n8094, n8095, n8096, n8097,
    n8098, n8099, n8100, n8101, n8102, n8103,
    n8104, n8105, n8106, n8107, n8108, n8109,
    n8110, n8111, n8112, n8113, n8114, n8115,
    n8116, n8117, n8118, n8119, n8120, n8121,
    n8122, n8123, n8124, n8125, n8126, n8127,
    n8128, n8129, n8130, n8131, n8132, n8133,
    n8134, n8135, n8136, n8137, n8138, n8139,
    n8140, n8141, n8142, n8143, n8144, n8145,
    n8146, n8147, n8148, n8149, n8150, n8151,
    n8152, n8153, n8154, n8155, n8156, n8157,
    n8158, n8159, n8160, n8161, n8162, n8163,
    n8164, n8165, n8166, n8167, n8168, n8169,
    n8170, n8171, n8172, n8173, n8174, n8175,
    n8176, n8177, n8178, n8179, n8180, n8181,
    n8182, n8183, n8184, n8185, n8186, n8187,
    n8188, n8189, n8190, n8191, n8192, n8193,
    n8194, n8195, n8196, n8197, n8198, n8199,
    n8200, n8201, n8202, n8203, n8204, n8205,
    n8206, n8207, n8208, n8209, n8210, n8211,
    n8212, n8213, n8214, n8215, n8216, n8217,
    n8218, n8219, n8220, n8221, n8222, n8223,
    n8224, n8225, n8226, n8227, n8228, n8229,
    n8230, n8231, n8232, n8233, n8234, n8235,
    n8236, n8237, n8238, n8239, n8240, n8241,
    n8242, n8243, n8244, n8245, n8246, n8247,
    n8248, n8249, n8250, n8251, n8252, n8253,
    n8254, n8255, n8256, n8257, n8258, n8259,
    n8260, n8261, n8262, n8263, n8264, n8265,
    n8266, n8267, n8268, n8269, n8270, n8271,
    n8272, n8273, n8274, n8275, n8276, n8277,
    n8278, n8279, n8280, n8281, n8282, n8283,
    n8284, n8285, n8286, n8287, n8288, n8289,
    n8290, n8291, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301,
    n8302, n8303, n8304, n8305, n8306, n8307,
    n8308, n8309, n8310, n8311, n8312, n8313,
    n8314, n8315, n8316, n8317, n8318, n8319,
    n8320, n8321, n8322, n8323, n8324, n8325,
    n8326, n8327, n8328, n8329, n8330, n8331,
    n8332, n8333, n8334, n8335, n8336, n8337,
    n8338, n8339, n8340, n8341, n8342, n8343,
    n8344, n8345, n8346, n8347, n8348, n8349,
    n8350, n8351, n8352, n8353, n8354, n8355,
    n8356, n8357, n8358, n8359, n8360, n8361,
    n8362, n8363, n8364, n8365, n8366, n8367,
    n8368, n8369, n8370, n8371, n8372, n8373,
    n8374, n8375, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385,
    n8386, n8387, n8388, n8389, n8390, n8391,
    n8392, n8393, n8394, n8395, n8396, n8397,
    n8398, n8399, n8400, n8401, n8402, n8403,
    n8404, n8405, n8406, n8407, n8408, n8409,
    n8410, n8411, n8412, n8413, n8414, n8415,
    n8416, n8417, n8418, n8419, n8421, n8422,
    n8423, n8424, n8425, n8426, n8427, n8428,
    n8429, n8430, n8431, n8432, n8433, n8434,
    n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446,
    n8447, n8448, n8449, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8463, n8464,
    n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476,
    n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494,
    n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8505, n8506,
    n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518,
    n8519, n8520, n8521, n8522, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530,
    n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548,
    n8549, n8550, n8551, n8552, n8553, n8554,
    n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8564, n8565, n8566,
    n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590,
    n8591, n8592, n8593, n8594, n8595, n8596,
    n8597, n8598, n8599, n8600, n8601, n8602,
    n8603, n8604, n8605, n8606, n8607, n8608,
    n8609, n8610, n8611, n8612, n8613, n8614,
    n8615, n8616, n8617, n8618, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626,
    n8627, n8628, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8636, n8637, n8638,
    n8639, n8640, n8641, n8642, n8643, n8644,
    n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656,
    n8657, n8658, n8659, n8660, n8661, n8662,
    n8663, n8664, n8665, n8666, n8667, n8668,
    n8669, n8670, n8671, n8672, n8673, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686,
    n8687, n8688, n8689, n8690, n8691, n8692,
    n8693, n8694, n8695, n8696, n8697, n8698,
    n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722,
    n8723, n8724, n8725, n8726, n8727, n8728,
    n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746,
    n8747, n8748, n8749, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8757, n8758,
    n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776,
    n8777, n8778, n8779, n8780, n8781, n8782,
    n8783, n8784, n8785, n8786, n8787, n8788,
    n8789, n8790, n8791, n8792, n8793, n8794,
    n8795, n8796, n8797, n8798, n8799, n8800,
    n8801, n8802, n8803, n8804, n8805, n8806,
    n8807, n8808, n8809, n8810, n8811, n8812,
    n8813, n8814, n8815, n8816, n8817, n8818,
    n8819, n8820, n8821, n8822, n8823, n8824,
    n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836,
    n8838, n8839, n8840, n8841, n8842, n8843,
    n8844, n8845, n8846, n8847, n8848, n8849,
    n8850, n8851, n8852, n8853, n8854, n8855,
    n8856, n8857, n8858, n8859, n8860, n8861,
    n8862, n8863, n8864, n8866, n8867, n8868,
    n8869, n8870, n8871, n8872, n8873, n8874,
    n8875, n8876, n8877, n8878, n8879, n8880,
    n8881, n8882, n8883, n8884, n8885, n8886,
    n8887, n8888, n8889, n8890, n8891, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898,
    n8899, n8900, n8901, n8902, n8903, n8904,
    n8905, n8906, n8907, n8908, n8909, n8910,
    n8911, n8912, n8913, n8914, n8915, n8916,
    n8917, n8918, n8919, n8920, n8921, n8922,
    n8923, n8924, n8925, n8926, n8927, n8928,
    n8929, n8930, n8931, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8940, n8941,
    n8942, n8943, n8944, n8945, n8946, n8947,
    n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8956, n8957, n8958, n8959,
    n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971,
    n8972, n8973, n8974, n8975, n8976, n8977,
    n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989,
    n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001,
    n9002, n9003, n9004, n9005, n9006, n9007,
    n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019,
    n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031,
    n9032, n9033, n9034, n9035, n9036, n9037,
    n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061,
    n9062, n9063, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073,
    n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121,
    n9122, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151,
    n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259,
    n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271,
    n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289,
    n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301,
    n9302, n9303, n9304, n9305, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9313,
    n9314, n9315, n9316, n9317, n9318, n9319,
    n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331,
    n9332, n9333, n9334, n9335, n9336, n9337,
    n9338, n9339, n9340, n9341, n9342, n9343,
    n9344, n9345, n9346, n9347, n9348, n9349,
    n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361,
    n9362, n9363, n9364, n9365, n9366, n9367,
    n9368, n9369, n9370, n9371, n9372, n9373,
    n9374, n9375, n9376, n9377, n9378, n9379,
    n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391,
    n9392, n9393, n9394, n9395, n9396, n9397,
    n9398, n9399, n9400, n9401, n9402, n9403,
    n9404, n9405, n9406, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421,
    n9422, n9423, n9424, n9425, n9426, n9427,
    n9428, n9429, n9430, n9431, n9432, n9433,
    n9434, n9435, n9436, n9437, n9438, n9439,
    n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451,
    n9452, n9453, n9454, n9455, n9456, n9457,
    n9458, n9459, n9460, n9461, n9462, n9463,
    n9464, n9465, n9466, n9467, n9468, n9469,
    n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481,
    n9482, n9483, n9484, n9485, n9486, n9487,
    n9488, n9489, n9490, n9491, n9492, n9493,
    n9494, n9495, n9496, n9497, n9498, n9499,
    n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511,
    n9512, n9513, n9514, n9515, n9516, n9517,
    n9518, n9519, n9520, n9521, n9522, n9523,
    n9524, n9525, n9526, n9527, n9528, n9529,
    n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541,
    n9542, n9543, n9544, n9545, n9546, n9547,
    n9548, n9549, n9550, n9551, n9552, n9553,
    n9554, n9555, n9556, n9557, n9558, n9559,
    n9560, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9570, n9571,
    n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583,
    n9584, n9585, n9586, n9587, n9588, n9589,
    n9590, n9591, n9592, n9593, n9594, n9595,
    n9596, n9597, n9598, n9599, n9600, n9601,
    n9602, n9603, n9604, n9605, n9606, n9607,
    n9608, n9609, n9610, n9611, n9612, n9613,
    n9614, n9615, n9616, n9617, n9618, n9619,
    n9620, n9621, n9622, n9623, n9624, n9625,
    n9626, n9627, n9628, n9629, n9630, n9631,
    n9632, n9633, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10017,
    n10018, n10019, n10020, n10021, n10022, n10023,
    n10024, n10025, n10026, n10027, n10028, n10029,
    n10030, n10031, n10032, n10033, n10034, n10035,
    n10036, n10037, n10038, n10039, n10040, n10041,
    n10042, n10043, n10044, n10045, n10046, n10047,
    n10048, n10049, n10050, n10051, n10052, n10053,
    n10054, n10055, n10056, n10057, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065,
    n10066, n10067, n10068, n10069, n10070, n10071,
    n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083,
    n10084, n10085, n10086, n10087, n10088, n10089,
    n10090, n10091, n10093, n10094, n10095, n10096,
    n10097, n10098, n10099, n10100, n10101, n10102,
    n10103, n10104, n10105, n10106, n10107, n10108,
    n10109, n10110, n10111, n10112, n10113, n10115,
    n10116, n10117, n10118, n10119, n10120, n10121,
    n10122, n10123, n10124, n10125, n10126, n10127,
    n10128, n10129, n10130, n10131, n10132, n10133,
    n10134, n10135, n10136, n10137, n10138, n10139,
    n10140, n10141, n10142, n10143, n10144, n10146,
    n10147, n10148, n10149, n10150, n10151, n10152,
    n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170,
    n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188,
    n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200,
    n10201, n10202, n10203, n10204, n10205, n10206,
    n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218,
    n10219, n10220, n10221, n10222, n10223, n10224,
    n10225, n10227, n10228, n10229, n10230, n10231,
    n10232, n10233, n10234, n10235, n10236, n10237,
    n10238, n10240, n10241, n10242, n10243, n10244,
    n10245, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256,
    n10257, n10258, n10259, n10260, n10261, n10262,
    n10263, n10264, n10265, n10266, n10267, n10268,
    n10269, n10270, n10271, n10272, n10273, n10274,
    n10275, n10276, n10277, n10278, n10279, n10280,
    n10281, n10282, n10283, n10284, n10285, n10286,
    n10287, n10288, n10289, n10290, n10291, n10292,
    n10293, n10294, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10303, n10304,
    n10305, n10306, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10315, n10316,
    n10317, n10318, n10319, n10320, n10321, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328,
    n10329, n10330, n10331, n10332, n10333, n10334,
    n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346,
    n10347, n10348, n10349, n10350, n10351, n10352,
    n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364,
    n10365, n10366, n10367, n10368, n10369, n10370,
    n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382,
    n10383, n10384, n10385, n10386, n10387, n10388,
    n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406,
    n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424,
    n10426, n10427, n10428, n10429, n10430, n10431,
    n10432, n10433, n10434, n10435, n10436, n10437,
    n10438, n10439, n10440, n10441, n10442, n10443,
    n10444, n10445, n10446, n10447, n10448, n10449,
    n10450, n10451, n10452, n10453, n10454, n10455,
    n10456, n10457, n10458, n10459, n10460, n10461,
    n10462, n10463, n10464, n10465, n10466, n10467,
    n10468, n10469, n10470, n10471, n10472, n10473,
    n10474, n10475, n10476, n10477, n10478, n10479,
    n10480, n10481, n10482, n10483, n10484, n10485,
    n10486, n10487, n10488, n10489, n10490, n10491,
    n10492, n10493, n10494, n10495, n10496, n10497,
    n10498, n10499, n10500, n10501, n10502, n10503,
    n10504, n10505, n10506, n10507, n10508, n10509,
    n10510, n10511, n10512, n10513, n10514, n10515,
    n10516, n10517, n10518, n10519, n10520, n10521,
    n10522, n10523, n10524, n10525, n10526, n10527,
    n10528, n10529, n10530, n10531, n10532, n10533,
    n10534, n10535, n10536, n10537, n10538, n10539,
    n10540, n10541, n10542, n10543, n10544, n10545,
    n10546, n10547, n10548, n10549, n10550, n10551,
    n10552, n10553, n10554, n10555, n10556, n10557,
    n10558, n10559, n10560, n10561, n10562, n10563,
    n10564, n10565, n10566, n10567, n10568, n10569,
    n10570, n10571, n10572, n10573, n10574, n10575,
    n10576, n10577, n10578, n10579, n10580, n10581,
    n10582, n10583, n10584, n10585, n10586, n10587,
    n10588, n10589, n10590, n10591, n10592, n10593,
    n10594, n10595, n10596, n10597, n10598, n10599,
    n10600, n10601, n10602, n10603, n10604, n10605,
    n10606, n10607, n10608, n10609, n10610, n10611,
    n10612, n10613, n10614, n10615, n10616, n10617,
    n10618, n10619, n10620, n10621, n10622, n10623,
    n10624, n10625, n10626, n10627, n10628, n10629,
    n10630, n10631, n10632, n10633, n10634, n10635,
    n10636, n10637, n10638, n10639, n10640, n10641,
    n10642, n10643, n10644, n10645, n10646, n10647,
    n10648, n10649, n10650, n10651, n10652, n10653,
    n10654, n10655, n10656, n10657, n10658, n10659,
    n10660, n10661, n10662, n10663, n10664, n10665,
    n10666, n10667, n10669, n10670, n10671, n10672,
    n10673, n10674, n10675, n10676, n10677, n10678,
    n10679, n10680, n10681, n10682, n10683, n10684,
    n10685, n10686, n10687, n10688, n10689, n10690,
    n10691, n10692, n10693, n10694, n10695, n10696,
    n10697, n10698, n10699, n10700, n10701, n10702,
    n10703, n10704, n10705, n10706, n10707, n10708,
    n10709, n10710, n10711, n10712, n10713, n10714,
    n10715, n10716, n10717, n10718, n10719, n10720,
    n10721, n10722, n10723, n10724, n10725, n10726,
    n10727, n10728, n10729, n10730, n10731, n10732,
    n10733, n10734, n10735, n10736, n10737, n10738,
    n10739, n10740, n10741, n10742, n10743, n10744,
    n10745, n10746, n10747, n10748, n10749, n10750,
    n10751, n10752, n10753, n10754, n10755, n10756,
    n10757, n10758, n10759, n10760, n10761, n10762,
    n10763, n10764, n10765, n10766, n10767, n10768,
    n10769, n10770, n10771, n10772, n10773, n10774,
    n10775, n10776, n10777, n10778, n10779, n10780,
    n10781, n10782, n10783, n10784, n10785, n10786,
    n10787, n10788, n10789, n10790, n10791, n10792,
    n10793, n10794, n10795, n10796, n10797, n10798,
    n10799, n10800, n10801, n10802, n10803, n10804,
    n10805, n10806, n10807, n10808, n10809, n10810,
    n10811, n10812, n10813, n10814, n10815, n10816,
    n10817, n10818, n10819, n10820, n10821, n10822,
    n10823, n10824, n10825, n10826, n10827, n10828,
    n10829, n10830, n10831, n10832, n10833, n10834,
    n10835, n10836, n10837, n10838, n10839, n10840,
    n10841, n10842, n10843, n10844, n10845, n10846,
    n10848, n10849, n10850, n10851, n10852, n10853,
    n10854, n10855, n10856, n10857, n10858, n10859,
    n10860, n10861, n10862, n10863, n10864, n10865,
    n10866, n10867, n10868, n10869, n10870, n10871,
    n10872, n10873, n10874, n10875, n10876, n10877,
    n10878, n10879, n10880, n10881, n10882, n10883,
    n10884, n10885, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10894, n10895,
    n10896, n10897, n10898, n10899, n10900, n10901,
    n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10911, n10912, n10913,
    n10914, n10915, n10916, n10917, n10918, n10919,
    n10920, n10922, n10923, n10924, n10926, n10927,
    n10928, n10929, n10930, n10931, n10932, n10933,
    n10934, n10935, n10936, n10937, n10938, n10939,
    n10940, n10941, n10942, n10943, n10944, n10946,
    n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958,
    n10959, n10960, n10961, n10962, n10963, n10964,
    n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10981, n10982,
    n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10991, n10992, n10993, n10994, n10995,
    n10997, n10998, n10999, n11000, n11001, n11002,
    n11003, n11004, n11005, n11006, n11007, n11008,
    n11009, n11010, n11011, n11012, n11013, n11014,
    n11016, n11017, n11018, n11019, n11020, n11021,
    n11022, n11023, n11024, n11025, n11026, n11027,
    n11028, n11029, n11030, n11031, n11032, n11033,
    n11034, n11035, n11036, n11037, n11038, n11039,
    n11040, n11042, n11043, n11044, n11045, n11046,
    n11047, n11048, n11050, n11051, n11052, n11053,
    n11054, n11055, n11056, n11057, n11058, n11059,
    n11060, n11061, n11062, n11063, n11064, n11065,
    n11066, n11067, n11068, n11069, n11070, n11071,
    n11072, n11073, n11074, n11075, n11076, n11077,
    n11078, n11079, n11080, n11081, n11082, n11083,
    n11084, n11085, n11086, n11087, n11088, n11089,
    n11090, n11091, n11092, n11093, n11094, n11095,
    n11096, n11097, n11098, n11099, n11100, n11101,
    n11102, n11103, n11104, n11105, n11106, n11107,
    n11108, n11109, n11110, n11111, n11112, n11113,
    n11114, n11115, n11116, n11117, n11118, n11119,
    n11120, n11121, n11122, n11123, n11124, n11125,
    n11126, n11127, n11128, n11129, n11130, n11131,
    n11132, n11133, n11134, n11135, n11136, n11137,
    n11138, n11139, n11140, n11141, n11142, n11143,
    n11144, n11145, n11146, n11147, n11148, n11149,
    n11150, n11151, n11152, n11153, n11154, n11155,
    n11156, n11157, n11158, n11159, n11160, n11161,
    n11162, n11163, n11164, n11165, n11166, n11167,
    n11168, n11169, n11170, n11171, n11172, n11173,
    n11174, n11175, n11176, n11177, n11178, n11179,
    n11180, n11181, n11182, n11183, n11184, n11185,
    n11186, n11187, n11188, n11189, n11190, n11191,
    n11192, n11193, n11194, n11195, n11196, n11197,
    n11198, n11199, n11201, n11202, n11203, n11204,
    n11205, n11206, n11207, n11208, n11209, n11210,
    n11211, n11213, n11214, n11215, n11216, n11217,
    n11218, n11219, n11220, n11221, n11222, n11223,
    n11224, n11225, n11226, n11227, n11228, n11229,
    n11230, n11231, n11233, n11234, n11235, n11236,
    n11237, n11238, n11239, n11240, n11241, n11242,
    n11243, n11244, n11245, n11247, n11248, n11249,
    n11250, n11251, n11252, n11253, n11255, n11256,
    n11257, n11258, n11259, n11260, n11261, n11262,
    n11263, n11265, n11266, n11268, n11269, n11270,
    n11271, n11272, n11274, n11275, n11276, n11277,
    n11278, n11279, n11280, n11281, n11283, n11284,
    n11285, n11286, n11288, n11289, n11290, n11291,
    n11293, n11294, n11295, n11296, n11297, n11299,
    n11300, n11301, n11302, n11303, n11304, n11305,
    n11307, n11308, n11309, n11311, n11312, n11313,
    n11314, n11315, n11316, n11317, n11318, n11319,
    n11320, n11321, n11322, n11323, n11324, n11325,
    n11326, n11328, n11329, n11330, n11331, n11333,
    n11334, n11335, n11336, n11337, n11338, n11339,
    n11341, n11342, n11343, n11344, n11345, n11346,
    n11347, n11348, n11349, n11350, n11351, n11353,
    n11354, n11355, n11356, n11357, n11358, n11359,
    n11360, n11361, n11362, n11363, n11364, n11365,
    n11366, n11367, n11368, n11369, n11370, n11371,
    n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11386, n11387, n11388, n11389, n11390,
    n11391, n11392, n11393, n11395, n11396, n11397,
    n11398, n11399, n11400, n11401, n11402, n11403,
    n11404, n11405, n11406, n11407, n11408, n11410,
    n11411, n11412, n11413, n11414, n11415, n11416,
    n11417, n11418, n11419, n11420, n11422, n11423,
    n11424, n11425, n11426, n11427, n11428, n11429,
    n11430, n11431, n11432, n11433, n11434, n11435,
    n11437, n11438, n11439, n11440, n11441, n11442,
    n11443, n11444, n11445, n11446, n11448, n11449,
    n11450, n11451, n11452, n11453, n11454, n11455,
    n11456, n11457, n11458, n11459, n11460, n11461,
    n11462, n11463, n11464, n11465, n11466, n11467,
    n11468, n11469, n11470, n11471, n11472, n11473,
    n11474, n11475, n11476, n11477, n11478, n11479,
    n11480, n11481, n11482, n11483, n11484, n11485,
    n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497,
    n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509,
    n11510, n11511, n11512, n11513, n11514, n11515,
    n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527,
    n11528, n11529, n11530, n11531, n11532, n11533,
    n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545,
    n11546, n11547, n11548, n11549, n11550, n11551,
    n11552, n11553, n11554, n11555, n11556, n11557,
    n11558, n11559, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569,
    n11570, n11571, n11572, n11573, n11574, n11575,
    n11576, n11577, n11578, n11579, n11580, n11581,
    n11582, n11583, n11584, n11585, n11586, n11587,
    n11588, n11589, n11590, n11591, n11592, n11593,
    n11594, n11595, n11596, n11597, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606,
    n11607, n11609, n11611, n11612, n11613, n11614,
    n11615, n11616, n11617, n11618, n11619, n11620,
    n11621, n11622, n11623, n11624, n11625, n11626,
    n11627, n11628, n11629, n11630, n11631, n11632,
    n11633, n11634, n11635, n11636, n11637, n11638,
    n11639, n11640, n11641, n11642, n11643, n11644,
    n11645, n11646, n11647, n11648, n11649, n11650,
    n11651, n11652, n11653, n11654, n11655, n11656,
    n11657, n11658, n11659, n11660, n11661, n11662,
    n11663, n11664, n11665, n11666, n11667, n11668,
    n11669, n11670, n11671, n11672, n11673, n11674,
    n11675, n11676, n11677, n11678, n11679, n11680,
    n11681, n11682, n11683, n11684, n11685, n11686,
    n11687, n11688, n11689, n11690, n11691, n11692,
    n11693, n11694, n11695, n11696, n11697, n11698,
    n11699, n11700, n11701, n11702, n11703, n11704,
    n11705, n11706, n11707, n11708, n11709, n11710,
    n11711, n11712, n11713, n11714, n11715, n11716,
    n11717, n11718, n11719, n11720, n11721, n11722,
    n11723, n11724, n11725, n11726, n11727, n11728,
    n11729, n11730, n11731, n11732, n11733, n11734,
    n11735, n11736, n11737, n11738, n11739, n11740,
    n11741, n11742, n11743, n11744, n11745, n11746,
    n11747, n11748, n11749, n11750, n11751, n11752,
    n11753, n11754, n11755, n11756, n11757, n11758,
    n11759, n11760, n11761, n11762, n11763, n11764,
    n11765, n11766, n11767, n11768, n11769, n11770,
    n11771, n11772, n11773, n11774, n11775, n11776,
    n11777, n11778, n11779, n11780, n11781, n11782,
    n11783, n11784, n11785, n11786, n11787, n11788,
    n11789, n11790, n11791, n11792, n11793, n11794,
    n11795, n11796, n11797, n11798, n11799, n11800,
    n11801, n11802, n11803, n11804, n11805, n11806,
    n11807, n11808, n11809, n11810, n11811, n11812,
    n11813, n11814, n11815, n11816, n11817, n11818,
    n11819, n11820, n11821, n11822, n11823, n11824,
    n11825, n11826, n11827, n11828, n11829, n11830,
    n11831, n11832, n11833, n11834, n11835, n11836,
    n11837, n11838, n11839, n11840, n11841, n11842,
    n11843, n11844, n11845, n11846, n11847, n11848,
    n11849, n11850, n11851, n11852, n11853, n11854,
    n11855, n11856, n11857, n11858, n11859, n11860,
    n11861, n11862, n11863, n11864, n11865, n11866,
    n11867, n11868, n11869, n11870, n11871, n11872,
    n11873, n11874, n11875, n11876, n11877, n11878,
    n11879, n11880, n11881, n11882, n11883, n11884,
    n11885, n11886, n11887, n11888, n11889, n11890,
    n11891, n11892, n11893, n11894, n11895, n11896,
    n11897, n11898, n11899, n11900, n11901, n11902,
    n11903, n11904, n11905, n11906, n11907, n11908,
    n11909, n11910, n11911, n11912, n11913, n11914,
    n11915, n11916, n11917, n11918, n11919, n11920,
    n11921, n11922, n11923, n11924, n11925, n11926,
    n11927, n11928, n11929, n11930, n11931, n11932,
    n11933, n11934, n11935, n11936, n11937, n11938,
    n11939, n11940, n11941, n11942, n11943, n11944,
    n11945, n11946, n11947, n11948, n11949, n11950,
    n11951, n11952, n11953, n11954, n11955, n11956,
    n11957, n11958, n11959, n11960, n11961, n11962,
    n11963, n11964, n11965, n11966, n11967, n11968,
    n11969, n11970, n11971, n11972, n11973, n11974,
    n11975, n11976, n11977, n11978, n11979, n11980,
    n11981, n11982, n11983, n11984, n11985, n11986,
    n11987, n11988, n11989, n11990, n11991, n11992,
    n11993, n11994, n11995, n11996, n11997, n11998,
    n11999, n12000, n12001, n12002, n12003, n12004,
    n12005, n12006, n12007, n12008, n12009, n12010,
    n12011, n12012, n12013, n12014, n12015, n12016,
    n12017, n12018, n12019, n12020, n12021, n12022,
    n12023, n12024, n12025, n12026, n12027, n12028,
    n12029, n12030, n12031, n12032, n12033, n12034,
    n12035, n12036, n12037, n12038, n12039, n12040,
    n12041, n12042, n12043, n12044, n12045, n12046,
    n12047, n12048, n12049, n12050, n12051, n12052,
    n12053, n12054, n12055, n12056, n12057, n12058,
    n12059, n12060, n12061, n12062, n12063, n12064,
    n12065, n12066, n12067, n12068, n12069, n12070,
    n12071, n12072, n12073, n12074, n12075, n12076,
    n12077, n12078, n12079, n12080, n12081, n12082,
    n12083, n12084, n12085, n12086, n12087, n12088,
    n12089, n12090, n12091, n12092, n12093, n12094,
    n12095, n12096, n12097, n12098, n12099, n12100,
    n12101, n12102, n12103, n12104, n12105, n12106,
    n12107, n12108, n12109, n12111, n12112, n12113,
    n12114, n12115, n12116, n12117, n12118, n12119,
    n12120, n12121, n12122, n12123, n12124, n12125,
    n12126, n12127, n12128, n12129, n12130, n12131,
    n12132, n12133, n12134, n12135, n12136, n12137,
    n12138, n12139, n12140, n12141, n12142, n12143,
    n12144, n12145, n12146, n12147, n12148, n12149,
    n12150, n12151, n12152, n12153, n12154, n12155,
    n12156, n12157, n12158, n12159, n12160, n12161,
    n12162, n12163, n12164, n12165, n12166, n12167,
    n12168, n12169, n12170, n12171, n12172, n12173,
    n12174, n12175, n12176, n12177, n12178, n12179,
    n12180, n12181, n12182, n12183, n12184, n12185,
    n12186, n12187, n12188, n12189, n12190, n12191,
    n12192, n12193, n12194, n12195, n12196, n12197,
    n12198, n12199, n12200, n12201, n12202, n12203,
    n12204, n12205, n12206, n12207, n12208, n12209,
    n12210, n12211, n12212, n12213, n12214, n12215,
    n12216, n12217, n12218, n12219, n12220, n12221,
    n12222, n12223, n12224, n12225, n12226, n12227,
    n12228, n12229, n12230, n12231, n12232, n12233,
    n12234, n12235, n12236, n12237, n12238, n12239,
    n12240, n12241, n12242, n12243, n12244, n12245,
    n12246, n12247, n12248, n12249, n12250, n12251,
    n12252, n12253, n12254, n12255, n12256, n12257,
    n12258, n12259, n12260, n12261, n12262, n12263,
    n12264, n12265, n12266, n12267, n12268, n12269,
    n12270, n12271, n12272, n12273, n12274, n12275,
    n12276, n12277, n12278, n12279, n12280, n12281,
    n12282, n12283, n12284, n12285, n12286, n12287,
    n12288, n12289, n12290, n12291, n12292, n12293,
    n12294, n12295, n12296, n12297, n12298, n12299,
    n12300, n12301, n12302, n12303, n12304, n12305,
    n12306, n12307, n12308, n12309, n12310, n12311,
    n12312, n12313, n12314, n12315, n12316, n12317,
    n12318, n12319, n12320, n12321, n12322, n12323,
    n12324, n12325, n12326, n12327, n12328, n12329,
    n12330, n12331, n12332, n12333, n12334, n12335,
    n12336, n12337, n12338, n12339, n12340, n12341,
    n12342, n12343, n12344, n12345, n12346, n12347,
    n12348, n12349, n12350, n12351, n12352, n12353,
    n12354, n12355, n12356, n12357, n12358, n12359,
    n12360, n12361, n12362, n12363, n12364, n12365,
    n12366, n12367, n12368, n12369, n12370, n12371,
    n12372, n12373, n12374, n12375, n12376, n12377,
    n12378, n12379, n12380, n12381, n12382, n12383,
    n12384, n12385, n12386, n12387, n12388, n12389,
    n12390, n12391, n12392, n12393, n12394, n12395,
    n12396, n12397, n12398, n12399, n12400, n12401,
    n12402, n12403, n12404, n12405, n12406, n12407,
    n12408, n12409, n12410, n12411, n12412, n12413,
    n12414, n12415, n12416, n12417, n12418, n12419,
    n12420, n12421, n12422, n12423, n12424, n12425,
    n12426, n12427, n12428, n12429, n12430, n12431,
    n12432, n12433, n12434, n12435, n12436, n12437,
    n12438, n12439, n12440, n12441, n12442, n12443,
    n12444, n12445, n12446, n12447, n12448, n12449,
    n12450, n12451, n12452, n12453, n12454, n12455,
    n12456, n12457, n12458, n12459, n12460, n12461,
    n12462, n12463, n12464, n12465, n12466, n12467,
    n12468, n12469, n12470, n12471, n12472, n12473,
    n12474, n12475, n12476, n12477, n12478, n12479,
    n12480, n12481, n12482, n12483, n12484, n12485,
    n12486, n12487, n12488, n12489, n12490, n12491,
    n12492, n12493, n12494, n12495, n12496, n12497,
    n12498, n12499, n12500, n12501, n12502, n12503,
    n12504, n12505, n12506, n12507, n12508, n12509,
    n12510, n12511, n12512, n12513, n12514, n12515,
    n12516, n12517, n12518, n12519, n12520, n12521,
    n12522, n12523, n12524, n12525, n12526, n12527,
    n12528, n12529, n12530, n12531, n12532, n12533,
    n12534, n12535, n12536, n12537, n12538, n12539,
    n12540, n12541, n12542, n12543, n12544, n12545,
    n12546, n12547, n12548, n12549, n12550, n12551,
    n12552, n12553, n12554, n12555, n12556, n12557,
    n12558, n12559, n12560, n12561, n12562, n12563,
    n12564, n12565, n12566, n12567, n12568, n12569,
    n12570, n12571, n12572, n12573, n12574, n12575,
    n12576, n12577, n12578, n12579, n12580, n12581,
    n12582, n12583, n12584, n12585, n12586, n12587,
    n12588, n12589, n12590, n12591, n12592, n12593,
    n12594, n12595, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12604, n12605,
    n12606, n12607, n12608, n12609, n12610, n12611,
    n12612, n12613, n12614, n12615, n12616, n12617,
    n12618, n12619, n12620, n12621, n12622, n12623,
    n12624, n12625, n12626, n12627, n12628, n12629,
    n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641,
    n12642, n12643, n12644, n12645, n12646, n12647,
    n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659,
    n12660, n12661, n12662, n12663, n12664, n12665,
    n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677,
    n12678, n12679, n12680, n12681, n12682, n12683,
    n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12691, n12692, n12693, n12694, n12695,
    n12696, n12697, n12698, n12699, n12700, n12701,
    n12702, n12703, n12704, n12705, n12706, n12707,
    n12708, n12709, n12710, n12711, n12712, n12713,
    n12714, n12715, n12716, n12717, n12718, n12719,
    n12720, n12721, n12722, n12723, n12724, n12725,
    n12726, n12727, n12728, n12729, n12730, n12731,
    n12732, n12733, n12734, n12735, n12736, n12737,
    n12738, n12739, n12740, n12741, n12742, n12743,
    n12744, n12745, n12746, n12747, n12748, n12749,
    n12750, n12751, n12752, n12753, n12754, n12755,
    n12756, n12757, n12758, n12759, n12760, n12761,
    n12762, n12763, n12764, n12765, n12766, n12767,
    n12768, n12769, n12770, n12771, n12772, n12773,
    n12774, n12775, n12776, n12777, n12778, n12779,
    n12780, n12781, n12782, n12783, n12784, n12785,
    n12786, n12787, n12788, n12789, n12790, n12791,
    n12792, n12793, n12794, n12795, n12796, n12797,
    n12798, n12799, n12800, n12801, n12802, n12803,
    n12804, n12805, n12806, n12807, n12808, n12809,
    n12810, n12811, n12812, n12813, n12814, n12815,
    n12816, n12817, n12818, n12819, n12820, n12821,
    n12822, n12823, n12824, n12825, n12826, n12827,
    n12828, n12829, n12830, n12831, n12832, n12833,
    n12834, n12835, n12836, n12837, n12838, n12839,
    n12840, n12841, n12842, n12843, n12844, n12845,
    n12846, n12847, n12848, n12849, n12850, n12851,
    n12852, n12853, n12854, n12855, n12856, n12857,
    n12858, n12859, n12860, n12861, n12862, n12863,
    n12864, n12865, n12866, n12867, n12868, n12869,
    n12870, n12871, n12872, n12873, n12874, n12875,
    n12876, n12877, n12878, n12879, n12880, n12881,
    n12882, n12883, n12884, n12885, n12886, n12887,
    n12888, n12889, n12890, n12891, n12892, n12893,
    n12894, n12895, n12896, n12897, n12898, n12899,
    n12900, n12901, n12902, n12903, n12904, n12905,
    n12906, n12907, n12908, n12909, n12910, n12911,
    n12912, n12913, n12914, n12915, n12916, n12917,
    n12918, n12919, n12920, n12921, n12922, n12923,
    n12924, n12925, n12926, n12927, n12928, n12929,
    n12930, n12931, n12932, n12933, n12934, n12935,
    n12936, n12937, n12938, n12939, n12940, n12941,
    n12942, n12943, n12944, n12946, n12947, n12948,
    n12949, n12950, n12951, n12952, n12953, n12954,
    n12956, n12957, n12958, n12959, n12960, n12961,
    n12962, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974,
    n12975, n12976, n12978, n12979, n12980, n12981,
    n12982, n12984, n12985, n12986, n12987, n12989,
    n12990, n12991, n12993, n12994, n12995, n12997,
    n12998, n12999, n13000, n13001, n13002, n13003,
    n13004, n13005, n13006, n13007, n13008, n13009,
    n13010, n13011, n13012, n13013, n13014, n13015,
    n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13027, n13028, n13029,
    n13030, n13032, n13033, n13034, n13035, n13036,
    n13037, n13038, n13039, n13040, n13041, n13042,
    n13044, n13045, n13046, n13047, n13048, n13049,
    n13050, n13051, n13052, n13053, n13054, n13056,
    n13057, n13058, n13059, n13060, n13061, n13063,
    n13064, n13065, n13066, n13067, n13068, n13069,
    n13070, n13071, n13072, n13073, n13074, n13075,
    n13076, n13077, n13078, n13079, n13081, n13082,
    n13083, n13084, n13085, n13086, n13087, n13088,
    n13089, n13090, n13091, n13092, n13093, n13094,
    n13095, n13097, n13098, n13099, n13100, n13101,
    n13102, n13103, n13104, n13105, n13106, n13108,
    n13109, n13110, n13111, n13112, n13113, n13114,
    n13115, n13116, n13118, n13119, n13120, n13121,
    n13123, n13124, n13125, n13126, n13127, n13128,
    n13129, n13130, n13131, n13132, n13133, n13134,
    n13135, n13136, n13137, n13138, n13139, n13140,
    n13141, n13142, n13143, n13144, n13145, n13146,
    n13147, n13148, n13149, n13150, n13151, n13152,
    n13153, n13154, n13155, n13156, n13157, n13158,
    n13159, n13160, n13161, n13162, n13163, n13164,
    n13165, n13166, n13167, n13168, n13169, n13170,
    n13171, n13172, n13173, n13174, n13175, n13176,
    n13177, n13178, n13179, n13180, n13181, n13182,
    n13183, n13184, n13185, n13186, n13187, n13188,
    n13189, n13190, n13191, n13192, n13193, n13194,
    n13195, n13196, n13197, n13199, n13200, n13201,
    n13202, n13203, n13204, n13205, n13206, n13207,
    n13208, n13209, n13210, n13211, n13212, n13213,
    n13214, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232,
    n13233, n13234, n13235, n13236, n13237, n13238,
    n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250,
    n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13297, n13299, n13300,
    n13301, n13302, n13303, n13304, n13305, n13307,
    n13308, n13309, n13310, n13311, n13312, n13313,
    n13314, n13315, n13316, n13317, n13318, n13319,
    n13320, n13321, n13322, n13323, n13325, n13326,
    n13327, n13328, n13329, n13330, n13331, n13332,
    n13333, n13335, n13337, n13338, n13339, n13340,
    n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352,
    n13353, n13355, n13357, n13358, n13359, n13360,
    n13361, n13362, n13363, n13364, n13366, n13367,
    n13368, n13369, n13370, n13373, n13374, n13375,
    n13376, n13377, n13378, n13379, n13380, n13381,
    n13382, n13383, n13384, n13385, n13386, n13387,
    n13388, n13389, n13390, n13391, n13392, n13393,
    n13394, n13395, n13396, n13397, n13398, n13399,
    n13400, n13401, n13402, n13403, n13404, n13405,
    n13406, n13407, n13408, n13409, n13410, n13411,
    n13412, n13413, n13414, n13415, n13416, n13417,
    n13418, n13419, n13420, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430,
    n13431, n13432, n13433, n13434, n13435, n13436,
    n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448,
    n13449, n13450, n13451, n13452, n13453, n13454,
    n13455, n13456, n13457, n13458, n13459, n13460,
    n13461, n13462, n13463, n13465, n13466, n13467,
    n13468, n13469, n13470, n13471, n13472, n13473,
    n13474, n13475, n13476, n13477, n13478, n13479,
    n13480, n13481, n13482, n13483, n13484, n13485,
    n13486, n13487, n13488, n13489, n13490, n13491,
    n13492, n13493, n13494, n13495, n13496, n13497,
    n13498, n13499, n13500, n13501, n13502, n13503,
    n13504, n13505, n13507, n13508, n13509, n13510,
    n13511, n13512, n13513, n13514, n13515, n13516,
    n13517, n13518, n13519, n13520, n13521, n13522,
    n13523, n13524, n13525, n13526, n13527, n13528,
    n13529, n13530, n13531, n13532, n13533, n13534,
    n13535, n13536, n13537, n13538, n13539, n13540,
    n13541, n13542, n13543, n13544, n13545, n13546,
    n13547, n13548, n13549, n13550, n13551, n13552,
    n13553, n13554, n13555, n13557, n13558, n13559,
    n13560, n13561, n13562, n13563, n13564, n13565,
    n13566, n13567, n13568, n13569, n13570, n13571,
    n13573, n13574, n13575, n13576, n13577, n13578,
    n13579, n13580, n13581, n13582, n13583, n13584,
    n13585, n13586, n13587, n13588, n13589, n13590,
    n13591, n13592, n13593, n13594, n13595, n13596,
    n13597, n13598, n13599, n13600, n13601, n13602,
    n13603, n13604, n13605, n13606, n13607, n13608,
    n13609, n13610, n13611, n13612, n13613, n13614,
    n13615, n13616, n13617, n13618, n13619, n13620,
    n13621, n13622, n13623, n13624, n13625, n13626,
    n13627, n13628, n13629, n13630, n13631, n13632,
    n13633, n13634, n13635, n13636, n13637, n13638,
    n13639, n13640, n13641, n13642, n13643, n13644,
    n13645, n13646, n13647, n13648, n13649, n13650,
    n13651, n13652, n13653, n13654, n13655, n13656,
    n13657, n13658, n13659, n13660, n13661, n13662,
    n13663, n13664, n13665, n13666, n13667, n13668,
    n13669, n13670, n13671, n13672, n13673, n13674,
    n13675, n13676, n13677, n13678, n13679, n13680,
    n13681, n13682, n13683, n13684, n13685, n13686,
    n13687, n13688, n13689, n13690, n13691, n13692,
    n13693, n13694, n13695, n13696, n13697, n13698,
    n13699, n13700, n13701, n13702, n13703, n13704,
    n13705, n13706, n13707, n13708, n13709, n13710,
    n13711, n13712, n13713, n13714, n13715, n13716,
    n13717, n13718, n13719, n13720, n13721, n13722,
    n13723, n13724, n13725, n13726, n13727, n13728,
    n13729, n13730, n13731, n13732, n13733, n13734,
    n13735, n13736, n13737, n13738, n13739, n13740,
    n13741, n13742, n13743, n13744, n13745, n13746,
    n13747, n13748, n13749, n13750, n13751, n13752,
    n13753, n13754, n13755, n13756, n13757, n13758,
    n13759, n13760, n13761, n13762, n13763, n13764,
    n13765, n13766, n13767, n13768, n13769, n13770,
    n13771, n13772, n13773, n13774, n13775, n13776,
    n13777, n13778, n13779, n13780, n13781, n13782,
    n13783, n13784, n13785, n13786, n13787, n13788,
    n13789, n13790, n13791, n13792, n13793, n13794,
    n13795, n13796, n13797, n13798, n13799, n13800,
    n13801, n13802, n13803, n13804, n13805, n13806,
    n13807, n13808, n13809, n13810, n13811, n13812,
    n13813, n13814, n13815, n13816, n13817, n13818,
    n13819, n13820, n13821, n13822, n13823, n13824,
    n13825, n13826, n13827, n13828, n13829, n13830,
    n13831, n13832, n13833, n13834, n13835, n13836,
    n13837, n13838, n13839, n13840, n13841, n13842,
    n13843, n13844, n13845, n13846, n13847, n13848,
    n13849, n13850, n13851, n13852, n13853, n13854,
    n13855, n13856, n13857, n13858, n13859, n13860,
    n13861, n13862, n13863, n13864, n13865, n13866,
    n13867, n13868, n13869, n13870, n13871, n13872,
    n13873, n13874, n13875, n13877, n13878, n13879,
    n13880, n13881, n13882, n13883, n13884, n13885,
    n13886, n13887, n13888, n13889, n13890, n13891,
    n13892, n13893, n13894, n13895, n13896, n13897,
    n13898, n13899, n13900, n13901, n13902, n13903,
    n13904, n13905, n13906, n13907, n13908, n13909,
    n13910, n13911, n13912, n13913, n13914, n13915,
    n13916, n13917, n13918, n13919, n13920, n13921,
    n13922, n13923, n13924, n13925, n13926, n13927,
    n13928, n13929, n13930, n13932, n13933, n13934,
    n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952,
    n13953, n13954, n13955, n13956, n13957, n13958,
    n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970,
    n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988,
    n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006,
    n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14041, n14042,
    n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054,
    n14055, n14056, n14057, n14058, n14059, n14060,
    n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078,
    n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14095, n14096,
    n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108,
    n14109, n14110, n14111, n14112, n14113, n14114,
    n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126,
    n14127, n14128, n14129, n14130, n14131, n14132,
    n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144,
    n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162,
    n14163, n14164, n14165, n14166, n14167, n14168,
    n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180,
    n14181, n14182, n14183, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198,
    n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216,
    n14217, n14218, n14219, n14220, n14221, n14222,
    n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240,
    n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252,
    n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14330, n14331,
    n14332, n14333, n14334, n14335, n14336, n14337,
    n14338, n14339, n14340, n14341, n14342, n14343,
    n14344, n14345, n14346, n14347, n14348, n14349,
    n14350, n14351, n14352, n14353, n14354, n14355,
    n14356, n14357, n14358, n14359, n14360, n14361,
    n14362, n14363, n14364, n14365, n14366, n14367,
    n14368, n14369, n14370, n14371, n14372, n14373,
    n14374, n14375, n14376, n14377, n14378, n14379,
    n14380, n14381, n14382, n14383, n14384, n14385,
    n14386, n14387, n14388, n14389, n14390, n14391,
    n14392, n14393, n14394, n14395, n14396, n14397,
    n14398, n14399, n14400, n14401, n14402, n14403,
    n14404, n14405, n14406, n14407, n14408, n14409,
    n14410, n14411, n14412, n14413, n14414, n14415,
    n14416, n14417, n14418, n14419, n14420, n14421,
    n14422, n14423, n14424, n14425, n14426, n14427,
    n14428, n14429, n14430, n14431, n14432, n14433,
    n14434, n14435, n14436, n14437, n14438, n14439,
    n14440, n14441, n14442, n14443, n14444, n14445,
    n14446, n14447, n14448, n14449, n14450, n14451,
    n14452, n14453, n14454, n14455, n14456, n14457,
    n14458, n14459, n14460, n14461, n14462, n14463,
    n14464, n14465, n14466, n14467, n14468, n14469,
    n14470, n14471, n14472, n14473, n14474, n14475,
    n14476, n14477, n14478, n14479, n14480, n14481,
    n14482, n14483, n14484, n14485, n14486, n14487,
    n14488, n14489, n14490, n14491, n14492, n14493,
    n14494, n14495, n14496, n14497, n14498, n14499,
    n14500, n14501, n14502, n14503, n14504, n14505,
    n14506, n14507, n14508, n14509, n14510, n14511,
    n14512, n14513, n14514, n14515, n14516, n14517,
    n14518, n14519, n14520, n14521, n14522, n14523,
    n14524, n14525, n14526, n14527, n14528, n14529,
    n14530, n14531, n14532, n14533, n14534, n14535,
    n14536, n14537, n14538, n14539, n14540, n14541,
    n14542, n14543, n14544, n14545, n14546, n14547,
    n14548, n14549, n14550, n14551, n14552, n14553,
    n14554, n14555, n14556, n14557, n14558, n14559,
    n14560, n14561, n14562, n14563, n14564, n14565,
    n14566, n14567, n14568, n14569, n14570, n14571,
    n14572, n14573, n14574, n14575, n14576, n14577,
    n14578, n14579, n14580, n14581, n14582, n14583,
    n14584, n14585, n14586, n14587, n14588, n14589,
    n14590, n14591, n14592, n14593, n14594, n14595,
    n14596, n14597, n14598, n14599, n14600, n14601,
    n14602, n14603, n14604, n14605, n14606, n14607,
    n14608, n14609, n14610, n14611, n14612, n14613,
    n14614, n14615, n14616, n14617, n14618, n14619,
    n14620, n14621, n14622, n14623, n14624, n14625,
    n14626, n14627, n14628, n14629, n14630, n14631,
    n14632, n14633, n14634, n14635, n14636, n14637,
    n14638, n14639, n14640, n14641, n14642, n14643,
    n14644, n14645, n14646, n14647, n14648, n14649,
    n14650, n14651, n14652, n14653, n14654, n14655,
    n14656, n14657, n14658, n14659, n14660, n14661,
    n14662, n14663, n14664, n14665, n14666, n14667,
    n14668, n14669, n14670, n14671, n14672, n14673,
    n14674, n14675, n14676, n14677, n14678, n14679,
    n14680, n14681, n14682, n14683, n14684, n14685,
    n14686, n14687, n14688, n14689, n14690, n14691,
    n14692, n14693, n14694, n14695, n14696, n14697,
    n14698, n14699, n14700, n14701, n14702, n14703,
    n14704, n14705, n14706, n14707, n14708, n14709,
    n14710, n14711, n14712, n14713, n14714, n14715,
    n14716, n14717, n14718, n14719, n14720, n14721,
    n14722, n14723, n14724, n14725, n14726, n14727,
    n14728, n14729, n14730, n14731, n14732, n14733,
    n14734, n14735, n14737, n14738, n14739, n14740,
    n14741, n14742, n14743, n14745, n14746, n14747,
    n14748, n14749, n14750, n14751, n14752, n14753,
    n14754, n14755, n14756, n14757, n14758, n14759,
    n14760, n14761, n14762, n14763, n14764, n14765,
    n14766, n14767, n14768, n14769, n14770, n14771,
    n14772, n14773, n14774, n14775, n14776, n14777,
    n14778, n14779, n14780, n14781, n14782, n14783,
    n14784, n14785, n14786, n14787, n14788, n14789,
    n14790, n14791, n14792, n14793, n14794, n14795,
    n14796, n14797, n14799, n14800, n14801, n14802,
    n14803, n14804, n14805, n14806, n14807, n14808,
    n14809, n14810, n14811, n14812, n14813, n14814,
    n14815, n14816, n14817, n14818, n14819, n14820,
    n14821, n14822, n14823, n14824, n14825, n14826,
    n14827, n14828, n14829, n14830, n14831, n14832,
    n14833, n14834, n14835, n14836, n14837, n14838,
    n14839, n14840, n14841, n14842, n14843, n14844,
    n14845, n14846, n14847, n14848, n14849, n14850,
    n14851, n14852, n14853, n14854, n14855, n14856,
    n14857, n14858, n14859, n14860, n14861, n14862,
    n14863, n14864, n14865, n14866, n14867, n14868,
    n14869, n14870, n14871, n14872, n14873, n14874,
    n14875, n14876, n14877, n14878, n14879, n14880,
    n14881, n14882, n14883, n14884, n14885, n14886,
    n14887, n14888, n14889, n14890, n14891, n14892,
    n14893, n14894, n14895, n14896, n14897, n14898,
    n14899, n14900, n14901, n14902, n14903, n14904,
    n14905, n14906, n14907, n14908, n14909, n14910,
    n14911, n14912, n14913, n14914, n14915, n14916,
    n14917, n14918, n14919, n14920, n14921, n14922,
    n14923, n14924, n14925, n14926, n14927, n14928,
    n14929, n14930, n14931, n14932, n14933, n14934,
    n14935, n14936, n14937, n14938, n14939, n14940,
    n14941, n14942, n14943, n14944, n14945, n14946,
    n14947, n14948, n14949, n14950, n14951, n14952,
    n14953, n14954, n14955, n14956, n14957, n14958,
    n14959, n14960, n14961, n14962, n14963, n14964,
    n14965, n14966, n14967, n14968, n14969, n14970,
    n14971, n14972, n14973, n14974, n14975, n14976,
    n14977, n14978, n14979, n14980, n14981, n14982,
    n14983, n14984, n14985, n14986, n14987, n14988,
    n14989, n14990, n14991, n14992, n14993, n14994,
    n14995, n14996, n14997, n14998, n14999, n15000,
    n15001, n15002, n15003, n15004, n15005, n15006,
    n15007, n15008, n15009, n15010, n15011, n15012,
    n15013, n15014, n15015, n15016, n15017, n15018,
    n15019, n15020, n15021, n15022, n15023, n15024,
    n15025, n15026, n15027, n15028, n15029, n15030,
    n15031, n15032, n15033, n15034, n15035, n15036,
    n15037, n15038, n15039, n15040, n15041, n15042,
    n15043, n15044, n15045, n15046, n15047, n15048,
    n15049, n15050, n15051, n15052, n15053, n15054,
    n15055, n15056, n15057, n15058, n15059, n15060,
    n15061, n15062, n15063, n15064, n15065, n15066,
    n15067, n15068, n15069, n15070, n15071, n15072,
    n15073, n15074, n15075, n15076, n15077, n15078,
    n15079, n15080, n15081, n15082, n15083, n15084,
    n15085, n15086, n15087, n15088, n15089, n15090,
    n15091, n15092, n15093, n15094, n15095, n15096,
    n15097, n15098, n15099, n15100, n15101, n15102,
    n15103, n15104, n15105, n15106, n15107, n15108,
    n15109, n15110, n15111, n15112, n15113, n15114,
    n15115, n15116, n15117, n15118, n15119, n15120,
    n15121, n15122, n15123, n15124, n15125, n15126,
    n15127, n15128, n15129, n15130, n15131, n15132,
    n15133, n15134, n15135, n15136, n15137, n15138,
    n15139, n15140, n15141, n15142, n15143, n15144,
    n15145, n15146, n15147, n15148, n15149, n15150,
    n15151, n15152, n15153, n15154, n15155, n15156,
    n15157, n15158, n15159, n15160, n15161, n15162,
    n15163, n15164, n15165, n15166, n15167, n15168,
    n15169, n15170, n15171, n15172, n15173, n15174,
    n15175, n15176, n15177, n15178, n15179, n15180,
    n15181, n15182, n15183, n15184, n15185, n15186,
    n15187, n15188, n15189, n15190, n15191, n15192,
    n15193, n15194, n15195, n15196, n15197, n15198,
    n15199, n15200, n15201, n15202, n15203, n15205,
    n15206, n15207, n15208, n15209, n15210, n15211,
    n15212, n15213, n15214, n15215, n15216, n15217,
    n15218, n15219, n15220, n15221, n15222, n15223,
    n15224, n15225, n15226, n15227, n15228, n15229,
    n15230, n15231, n15232, n15233, n15234, n15235,
    n15236, n15237, n15238, n15239, n15240, n15241,
    n15242, n15243, n15244, n15245, n15246, n15247,
    n15248, n15249, n15250, n15251, n15252, n15253,
    n15254, n15255, n15256, n15257, n15258, n15259,
    n15260, n15261, n15262, n15263, n15264, n15265,
    n15266, n15267, n15268, n15269, n15270, n15271,
    n15272, n15273, n15274, n15275, n15276, n15277,
    n15278, n15279, n15280, n15281, n15282, n15283,
    n15284, n15285, n15286, n15287, n15288, n15289,
    n15290, n15291, n15292, n15293, n15294, n15295,
    n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307,
    n15308, n15309, n15310, n15311, n15312, n15313,
    n15314, n15315, n15316, n15317, n15318, n15319,
    n15320, n15321, n15322, n15323, n15324, n15325,
    n15326, n15327, n15328, n15329, n15330, n15331,
    n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343,
    n15344, n15345, n15346, n15347, n15348, n15349,
    n15350, n15351, n15352, n15353, n15354, n15355,
    n15356, n15357, n15358, n15359, n15360, n15361,
    n15362, n15363, n15364, n15365, n15366, n15367,
    n15368, n15369, n15370, n15371, n15372, n15373,
    n15374, n15375, n15376, n15377, n15378, n15379,
    n15380, n15381, n15382, n15383, n15384, n15385,
    n15386, n15387, n15388, n15389, n15390, n15391,
    n15392, n15393, n15394, n15395, n15396, n15397,
    n15398, n15399, n15400, n15401, n15402, n15403,
    n15404, n15405, n15406, n15407, n15408, n15409,
    n15410, n15411, n15412, n15413, n15414, n15415,
    n15416, n15417, n15418, n15419, n15420, n15421,
    n15422, n15423, n15424, n15425, n15426, n15427,
    n15428, n15429, n15430, n15431, n15432, n15433,
    n15434, n15435, n15436, n15437, n15438, n15439,
    n15440, n15441, n15442, n15443, n15444, n15445,
    n15446, n15447, n15448, n15449, n15450, n15451,
    n15452, n15453, n15454, n15455, n15456, n15457,
    n15458, n15459, n15460, n15461, n15462, n15463,
    n15464, n15465, n15466, n15467, n15468, n15469,
    n15470, n15471, n15472, n15473, n15474, n15475,
    n15476, n15477, n15478, n15479, n15480, n15481,
    n15482, n15483, n15484, n15485, n15486, n15487,
    n15488, n15489, n15490, n15491, n15492, n15493,
    n15494, n15495, n15496, n15497, n15498, n15499,
    n15500, n15501, n15502, n15503, n15504, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512,
    n15513, n15514, n15515, n15516, n15517, n15518,
    n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530,
    n15531, n15532, n15533, n15534, n15535, n15536,
    n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548,
    n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566,
    n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15599, n15600, n15601, n15602, n15603,
    n15604, n15605, n15606, n15607, n15608, n15609,
    n15610, n15611, n15612, n15613, n15614, n15615,
    n15616, n15617, n15618, n15619, n15620, n15621,
    n15622, n15624, n15625, n15626, n15627, n15628,
    n15629, n15630, n15631, n15632, n15633, n15634,
    n15635, n15636, n15637, n15638, n15639, n15640,
    n15641, n15642, n15643, n15644, n15645, n15646,
    n15647, n15648, n15649, n15650, n15651, n15652,
    n15653, n15654, n15655, n15656, n15657, n15658,
    n15659, n15660, n15661, n15662, n15663, n15664,
    n15665, n15666, n15667, n15668, n15669, n15670,
    n15671, n15672, n15673, n15674, n15675, n15676,
    n15677, n15678, n15679, n15680, n15681, n15682,
    n15683, n15684, n15685, n15686, n15687, n15688,
    n15689, n15690, n15691, n15692, n15693, n15694,
    n15695, n15696, n15697, n15698, n15699, n15700,
    n15701, n15702, n15703, n15704, n15705, n15706,
    n15707, n15708, n15709, n15710, n15711, n15712,
    n15713, n15714, n15715, n15716, n15717, n15718,
    n15719, n15720, n15721, n15722, n15723, n15724,
    n15725, n15726, n15727, n15728, n15729, n15730,
    n15731, n15732, n15733, n15734, n15735, n15736,
    n15737, n15738, n15739, n15740, n15741, n15742,
    n15743, n15744, n15745, n15746, n15747, n15748,
    n15749, n15750, n15751, n15752, n15753, n15754,
    n15755, n15756, n15757, n15759, n15760, n15761,
    n15762, n15763, n15764, n15765, n15767, n15768,
    n15769, n15770, n15771, n15772, n15773, n15774,
    n15775, n15776, n15777, n15778, n15779, n15780,
    n15781, n15782, n15783, n15784, n15785, n15786,
    n15787, n15788, n15789, n15790, n15791, n15792,
    n15793, n15794, n15795, n15796, n15797, n15798,
    n15799, n15800, n15801, n15802, n15803, n15804,
    n15805, n15806, n15807, n15808, n15809, n15810,
    n15811, n15812, n15813, n15814, n15815, n15816,
    n15817, n15818, n15819, n15820, n15821, n15822,
    n15823, n15824, n15825, n15826, n15827, n15828,
    n15829, n15830, n15831, n15832, n15833, n15834,
    n15835, n15836, n15837, n15838, n15839, n15840,
    n15841, n15842, n15843, n15844, n15845, n15846,
    n15847, n15848, n15849, n15850, n15851, n15852,
    n15853, n15854, n15855, n15856, n15857, n15858,
    n15859, n15860, n15861, n15862, n15863, n15864,
    n15865, n15866, n15867, n15868, n15869, n15870,
    n15871, n15872, n15873, n15874, n15875, n15876,
    n15877, n15878, n15879, n15880, n15881, n15882,
    n15883, n15884, n15885, n15886, n15887, n15888,
    n15889, n15890, n15891, n15892, n15893, n15894,
    n15895, n15896, n15897, n15898, n15899, n15900,
    n15901, n15902, n15903, n15904, n15905, n15906,
    n15907, n15908, n15909, n15910, n15911, n15912,
    n15913, n15914, n15915, n15916, n15917, n15918,
    n15919, n15920, n15921, n15922, n15923, n15924,
    n15925, n15926, n15927, n15928, n15929, n15930,
    n15931, n15932, n15933, n15934, n15935, n15936,
    n15937, n15938, n15939, n15940, n15941, n15942,
    n15943, n15944, n15945, n15946, n15947, n15948,
    n15949, n15950, n15951, n15952, n15953, n15954,
    n15955, n15956, n15957, n15958, n15959, n15960,
    n15961, n15962, n15963, n15964, n15965, n15966,
    n15967, n15968, n15969, n15970, n15971, n15972,
    n15973, n15974, n15975, n15976, n15977, n15978,
    n15979, n15981, n15982, n15983, n15984, n15985,
    n15986, n15987, n15988, n15989, n15990, n15991,
    n15992, n15993, n15994, n15995, n15996, n15997,
    n15998, n15999, n16000, n16001, n16002, n16003,
    n16004, n16005, n16006, n16007, n16008, n16009,
    n16010, n16011, n16012, n16013, n16014, n16015,
    n16016, n16017, n16018, n16019, n16020, n16021,
    n16022, n16023, n16024, n16025, n16026, n16027,
    n16028, n16029, n16030, n16031, n16032, n16033,
    n16034, n16035, n16036, n16037, n16038, n16039,
    n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088,
    n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106,
    n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16155,
    n16156, n16157, n16158, n16159, n16160, n16161,
    n16162, n16163, n16164, n16165, n16166, n16167,
    n16168, n16169, n16170, n16171, n16172, n16173,
    n16174, n16175, n16176, n16177, n16178, n16179,
    n16180, n16181, n16182, n16183, n16184, n16185,
    n16186, n16187, n16188, n16189, n16190, n16191,
    n16192, n16193, n16194, n16195, n16196, n16197,
    n16198, n16199, n16200, n16201, n16202, n16203,
    n16204, n16205, n16206, n16207, n16208, n16209,
    n16210, n16211, n16212, n16213, n16214, n16215,
    n16216, n16217, n16218, n16219, n16220, n16221,
    n16222, n16223, n16224, n16225, n16226, n16227,
    n16228, n16229, n16230, n16231, n16232, n16233,
    n16234, n16235, n16236, n16237, n16238, n16239,
    n16240, n16241, n16242, n16243, n16244, n16245,
    n16246, n16247, n16248, n16249, n16250, n16251,
    n16252, n16253, n16254, n16255, n16256, n16257,
    n16258, n16259, n16260, n16261, n16262, n16263,
    n16264, n16265, n16266, n16267, n16268, n16269,
    n16270, n16271, n16272, n16274, n16275, n16276,
    n16277, n16278, n16279, n16280, n16281, n16282,
    n16283, n16284, n16285, n16286, n16287, n16288,
    n16289, n16290, n16291, n16292, n16293, n16294,
    n16295, n16296, n16297, n16298, n16299, n16300,
    n16301, n16302, n16303, n16304, n16305, n16306,
    n16307, n16308, n16309, n16310, n16311, n16312,
    n16313, n16314, n16315, n16316, n16317, n16318,
    n16319, n16320, n16321, n16322, n16323, n16324,
    n16325, n16326, n16327, n16328, n16329, n16330,
    n16331, n16332, n16333, n16334, n16335, n16336,
    n16337, n16338, n16339, n16340, n16341, n16342,
    n16343, n16344, n16345, n16346, n16347, n16348,
    n16349, n16350, n16351, n16352, n16353, n16354,
    n16355, n16356, n16358, n16359, n16360, n16361,
    n16362, n16363, n16364, n16365, n16366, n16367,
    n16368, n16369, n16371, n16372, n16373, n16374,
    n16375, n16376, n16377, n16378, n16379, n16380,
    n16381, n16382, n16383, n16384, n16385, n16386,
    n16387, n16388, n16389, n16390, n16391, n16392,
    n16393, n16394, n16395, n16396, n16397, n16398,
    n16399, n16400, n16401, n16402, n16403, n16404,
    n16405, n16406, n16407, n16408, n16409, n16410,
    n16411, n16412, n16413, n16414, n16415, n16416,
    n16417, n16418, n16419, n16420, n16421, n16422,
    n16423, n16424, n16425, n16426, n16427, n16428,
    n16429, n16430, n16431, n16432, n16433, n16434,
    n16435, n16436, n16437, n16438, n16439, n16440,
    n16441, n16442, n16443, n16444, n16445, n16446,
    n16447, n16448, n16449, n16450, n16451, n16452,
    n16453, n16454, n16456, n16457, n16458, n16459,
    n16460, n16461, n16462, n16463, n16464, n16465,
    n16466, n16467, n16468, n16469, n16470, n16471,
    n16472, n16473, n16474, n16475, n16476, n16477,
    n16478, n16479, n16480, n16481, n16482, n16483,
    n16484, n16485, n16486, n16487, n16488, n16489,
    n16490, n16491, n16492, n16493, n16494, n16495,
    n16496, n16497, n16498, n16499, n16500, n16501,
    n16502, n16503, n16504, n16505, n16506, n16507,
    n16508, n16510, n16511, n16512, n16513, n16514,
    n16515, n16516, n16517, n16518, n16519, n16520,
    n16521, n16522, n16523, n16524, n16525, n16526,
    n16527, n16528, n16529, n16530, n16531, n16532,
    n16533, n16534, n16535, n16536, n16537, n16538,
    n16539, n16540, n16541, n16542, n16543, n16544,
    n16545, n16546, n16547, n16548, n16549, n16550,
    n16551, n16552, n16553, n16554, n16555, n16556,
    n16557, n16558, n16559, n16560, n16561, n16562,
    n16563, n16564, n16565, n16566, n16567, n16568,
    n16569, n16570, n16571, n16572, n16573, n16574,
    n16575, n16576, n16577, n16578, n16579, n16580,
    n16581, n16582, n16583, n16584, n16585, n16586,
    n16587, n16588, n16589, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598,
    n16599, n16600, n16601, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622,
    n16623, n16624, n16625, n16626, n16627, n16628,
    n16629, n16630, n16631, n16632, n16633, n16634,
    n16635, n16636, n16637, n16638, n16639, n16640,
    n16641, n16642, n16643, n16644, n16645, n16646,
    n16647, n16648, n16649, n16650, n16651, n16652,
    n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664,
    n16665, n16666, n16667, n16668, n16669, n16670,
    n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682,
    n16683, n16684, n16685, n16686, n16687, n16688,
    n16689, n16690, n16691, n16692, n16693, n16694,
    n16695, n16696, n16697, n16698, n16699, n16700,
    n16701, n16702, n16703, n16704, n16705, n16706,
    n16707, n16708, n16709, n16710, n16711, n16712,
    n16713, n16714, n16715, n16716, n16717, n16718,
    n16719, n16720, n16721, n16722, n16723, n16724,
    n16725, n16726, n16727, n16728, n16729, n16730,
    n16731, n16732, n16733, n16734, n16735, n16736,
    n16737, n16738, n16739, n16740, n16741, n16742,
    n16743, n16744, n16745, n16746, n16747, n16748,
    n16749, n16750, n16751, n16752, n16753, n16754,
    n16755, n16756, n16757, n16758, n16759, n16760,
    n16761, n16762, n16763, n16764, n16765, n16766,
    n16767, n16768, n16769, n16770, n16771, n16772,
    n16773, n16774, n16775, n16776, n16777, n16778,
    n16779, n16780, n16781, n16782, n16783, n16784,
    n16785, n16786, n16787, n16788, n16789, n16790,
    n16791, n16792, n16793, n16794, n16795, n16796,
    n16797, n16798, n16799, n16800, n16801, n16802,
    n16803, n16804, n16805, n16806, n16807, n16808,
    n16809, n16810, n16811, n16812, n16813, n16814,
    n16815, n16816, n16817, n16818, n16819, n16820,
    n16821, n16822, n16823, n16824, n16825, n16826,
    n16827, n16828, n16829, n16830, n16831, n16832,
    n16833, n16834, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844,
    n16845, n16846, n16847, n16848, n16849, n16850,
    n16851, n16852, n16853, n16854, n16855, n16856,
    n16857, n16858, n16859, n16860, n16861, n16862,
    n16863, n16864, n16865, n16866, n16867, n16868,
    n16869, n16870, n16871, n16872, n16873, n16874,
    n16875, n16876, n16877, n16878, n16879, n16880,
    n16881, n16882, n16883, n16884, n16885, n16886,
    n16887, n16888, n16889, n16890, n16891, n16892,
    n16893, n16894, n16895, n16896, n16897, n16898,
    n16899, n16900, n16901, n16902, n16903, n16904,
    n16905, n16906, n16907, n16908, n16909, n16910,
    n16911, n16912, n16913, n16914, n16915, n16916,
    n16917, n16918, n16919, n16920, n16921, n16922,
    n16923, n16924, n16925, n16926, n16927, n16928,
    n16929, n16930, n16931, n16932, n16933, n16934,
    n16935, n16936, n16937, n16938, n16939, n16940,
    n16941, n16942, n16943, n16944, n16945, n16946,
    n16947, n16948, n16949, n16950, n16951, n16952,
    n16953, n16954, n16955, n16956, n16957, n16958,
    n16959, n16960, n16961, n16962, n16963, n16964,
    n16965, n16966, n16967, n16968, n16969, n16970,
    n16971, n16972, n16973, n16974, n16975, n16976,
    n16977, n16978, n16979, n16980, n16981, n16982,
    n16983, n16984, n16985, n16986, n16987, n16988,
    n16989, n16990, n16991, n16992, n16993, n16995,
    n16996, n16997, n16998, n16999, n17000, n17001,
    n17002, n17003, n17004, n17005, n17006, n17007,
    n17008, n17009, n17010, n17011, n17012, n17013,
    n17014, n17015, n17016, n17017, n17018, n17019,
    n17020, n17021, n17022, n17023, n17024, n17025,
    n17026, n17027, n17028, n17029, n17030, n17031,
    n17032, n17033, n17034, n17035, n17036, n17037,
    n17038, n17039, n17040, n17041, n17042, n17043,
    n17044, n17045, n17046, n17047, n17048, n17049,
    n17050, n17051, n17052, n17053, n17054, n17055,
    n17056, n17057, n17058, n17059, n17060, n17061,
    n17062, n17063, n17064, n17065, n17066, n17067,
    n17068, n17069, n17070, n17071, n17072, n17073,
    n17074, n17075, n17076, n17077, n17078, n17079,
    n17080, n17081, n17082, n17083, n17084, n17085,
    n17086, n17087, n17088, n17089, n17090, n17091,
    n17092, n17093, n17094, n17095, n17096, n17097,
    n17098, n17099, n17100, n17101, n17102, n17103,
    n17104, n17105, n17106, n17107, n17108, n17109,
    n17110, n17111, n17112, n17113, n17114, n17115,
    n17116, n17117, n17118, n17119, n17120, n17121,
    n17122, n17123, n17124, n17125, n17126, n17127,
    n17128, n17129, n17130, n17131, n17132, n17133,
    n17134, n17135, n17136, n17137, n17138, n17139,
    n17140, n17141, n17142, n17143, n17144, n17145,
    n17146, n17147, n17148, n17149, n17150, n17151,
    n17152, n17153, n17154, n17155, n17156, n17157,
    n17158, n17159, n17160, n17161, n17162, n17163,
    n17164, n17165, n17166, n17167, n17168, n17169,
    n17170, n17171, n17172, n17173, n17174, n17175,
    n17176, n17177, n17178, n17179, n17180, n17181,
    n17182, n17183, n17184, n17185, n17186, n17187,
    n17188, n17189, n17190, n17191, n17192, n17193,
    n17194, n17195, n17196, n17197, n17198, n17199,
    n17200, n17201, n17202, n17203, n17204, n17205,
    n17206, n17207, n17208, n17209, n17210, n17211,
    n17212, n17213, n17214, n17215, n17216, n17217,
    n17218, n17219, n17220, n17221, n17222, n17223,
    n17224, n17225, n17226, n17227, n17228, n17229,
    n17230, n17231, n17232, n17233, n17234, n17235,
    n17236, n17237, n17238, n17239, n17240, n17241,
    n17242, n17243, n17244, n17245, n17246, n17247,
    n17248, n17249, n17250, n17251, n17252, n17253,
    n17254, n17255, n17256, n17257, n17258, n17259,
    n17260, n17261, n17262, n17263, n17264, n17265,
    n17266, n17267, n17268, n17269, n17270, n17271,
    n17272, n17273, n17274, n17275, n17276, n17277,
    n17278, n17279, n17280, n17281, n17282, n17283,
    n17284, n17285, n17286, n17287, n17288, n17289,
    n17290, n17291, n17292, n17293, n17294, n17295,
    n17296, n17297, n17298, n17299, n17300, n17301,
    n17302, n17303, n17304, n17305, n17306, n17307,
    n17308, n17309, n17310, n17311, n17312, n17313,
    n17314, n17315, n17316, n17317, n17318, n17319,
    n17320, n17321, n17322, n17323, n17324, n17325,
    n17326, n17327, n17328, n17329, n17330, n17331,
    n17332, n17333, n17334, n17335, n17336, n17337,
    n17338, n17339, n17340, n17341, n17342, n17343,
    n17344, n17345, n17346, n17347, n17348, n17349,
    n17350, n17351, n17352, n17353, n17354, n17355,
    n17356, n17357, n17358, n17359, n17360, n17361,
    n17362, n17363, n17364, n17365, n17366, n17367,
    n17368, n17369, n17370, n17371, n17372, n17373,
    n17374, n17375, n17376, n17377, n17378, n17379,
    n17380, n17381, n17382, n17383, n17384, n17385,
    n17386, n17387, n17388, n17389, n17390, n17391,
    n17392, n17393, n17394, n17395, n17396, n17397,
    n17398, n17399, n17400, n17401, n17402, n17403,
    n17404, n17405, n17406, n17407, n17408, n17409,
    n17410, n17411, n17412, n17413, n17414, n17415,
    n17416, n17417, n17418, n17419, n17420, n17421,
    n17422, n17423, n17424, n17425, n17426, n17427,
    n17428, n17429, n17430, n17431, n17432, n17433,
    n17434, n17435, n17436, n17437, n17438, n17439,
    n17440, n17441, n17442, n17443, n17444, n17445,
    n17446, n17447, n17448, n17449, n17450, n17451,
    n17452, n17453, n17454, n17455, n17456, n17457,
    n17458, n17459, n17460, n17461, n17462, n17463,
    n17464, n17465, n17466, n17467, n17468, n17469,
    n17470, n17471, n17472, n17473, n17474, n17475,
    n17476, n17477, n17478, n17479, n17480, n17481,
    n17482, n17483, n17484, n17485, n17486, n17487,
    n17488, n17489, n17490, n17491, n17492, n17493,
    n17494, n17495, n17496, n17497, n17498, n17499,
    n17500, n17501, n17502, n17503, n17504, n17505,
    n17506, n17507, n17508, n17509, n17510, n17511,
    n17512, n17513, n17514, n17515, n17516, n17517,
    n17518, n17519, n17520, n17521, n17522, n17523,
    n17524, n17525, n17526, n17527, n17528, n17529,
    n17530, n17531, n17532, n17533, n17534, n17535,
    n17536, n17537, n17538, n17539, n17540, n17541,
    n17542, n17543, n17544, n17545, n17546, n17547,
    n17548, n17549, n17550, n17551, n17552, n17553,
    n17554, n17555, n17556, n17557, n17558, n17559,
    n17560, n17561, n17562, n17563, n17564, n17565,
    n17566, n17567, n17568, n17569, n17570, n17571,
    n17572, n17573, n17574, n17575, n17576, n17577,
    n17578, n17579, n17580, n17581, n17582, n17583,
    n17584, n17585, n17586, n17587, n17588, n17589,
    n17590, n17591, n17592, n17593, n17594, n17595,
    n17596, n17597, n17598, n17599, n17600, n17601,
    n17602, n17603, n17604, n17605, n17606, n17607,
    n17608, n17609, n17610, n17611, n17612, n17613,
    n17614, n17615, n17616, n17617, n17618, n17619,
    n17620, n17621, n17622, n17623, n17624, n17625,
    n17626, n17627, n17628, n17629, n17630, n17631,
    n17632, n17633, n17634, n17635, n17636, n17637,
    n17638, n17639, n17640, n17641, n17642, n17643,
    n17644, n17645, n17646, n17647, n17648, n17649,
    n17650, n17651, n17652, n17653, n17654, n17655,
    n17656, n17657, n17658, n17659, n17660, n17661,
    n17662, n17663, n17664, n17665, n17666, n17667,
    n17668, n17669, n17670, n17671, n17672, n17673,
    n17674, n17675, n17676, n17677, n17678, n17679,
    n17680, n17681, n17682, n17683, n17684, n17685,
    n17686, n17687, n17688, n17689, n17690, n17691,
    n17692, n17693, n17694, n17695, n17696, n17697,
    n17698, n17699, n17700, n17701, n17702, n17703,
    n17704, n17705, n17706, n17707, n17708, n17709,
    n17710, n17711, n17712, n17713, n17714, n17715,
    n17716, n17717, n17718, n17719, n17720, n17721,
    n17722, n17723, n17724, n17725, n17726, n17727,
    n17728, n17729, n17730, n17731, n17732, n17733,
    n17734, n17735, n17736, n17737, n17738, n17739,
    n17740, n17741, n17742, n17743, n17744, n17745,
    n17746, n17747, n17748, n17749, n17750, n17751,
    n17752, n17753, n17754, n17755, n17756, n17757,
    n17758, n17759, n17760, n17761, n17762, n17763,
    n17764, n17765, n17766, n17767, n17768, n17769,
    n17770, n17771, n17772, n17773, n17774, n17775,
    n17776, n17777, n17778, n17779, n17780, n17781,
    n17782, n17783, n17784, n17785, n17786, n17787,
    n17788, n17789, n17790, n17791, n17792, n17793,
    n17794, n17795, n17796, n17797, n17798, n17799,
    n17800, n17801, n17802, n17803, n17804, n17805,
    n17806, n17807, n17808, n17809, n17810, n17811,
    n17812, n17813, n17814, n17815, n17816, n17817,
    n17818, n17819, n17820, n17821, n17822, n17823,
    n17824, n17825, n17826, n17827, n17828, n17829,
    n17830, n17831, n17832, n17833, n17834, n17835,
    n17836, n17837, n17838, n17839, n17840, n17841,
    n17842, n17843, n17844, n17845, n17846, n17847,
    n17848, n17849, n17850, n17851, n17852, n17853,
    n17854, n17855, n17856, n17857, n17858, n17859,
    n17860, n17861, n17862, n17863, n17864, n17865,
    n17866, n17867, n17868, n17869, n17870, n17871,
    n17872, n17873, n17874, n17875, n17876, n17877,
    n17878, n17879, n17880, n17881, n17882, n17883,
    n17884, n17885, n17886, n17887, n17888, n17889,
    n17890, n17891, n17892, n17893, n17894, n17895,
    n17896, n17897, n17898, n17899, n17900, n17901,
    n17902, n17903, n17904, n17905, n17906, n17907,
    n17908, n17909, n17910, n17911, n17912, n17914,
    n17915, n17916, n17917, n17918, n17919, n17920,
    n17921, n17922, n17923, n17924, n17925, n17926,
    n17927, n17928, n17929, n17930, n17931, n17932,
    n17933, n17934, n17935, n17936, n17937, n17938,
    n17939, n17940, n17941, n17942, n17943, n17944,
    n17945, n17946, n17947, n17948, n17949, n17950,
    n17951, n17952, n17953, n17954, n17955, n17956,
    n17957, n17958, n17959, n17960, n17961, n17962,
    n17963, n17964, n17965, n17966, n17967, n17968,
    n17969, n17970, n17971, n17972, n17973, n17974,
    n17975, n17976, n17977, n17978, n17979, n17980,
    n17981, n17982, n17983, n17984, n17985, n17986,
    n17987, n17988, n17989, n17990, n17991, n17992,
    n17993, n17994, n17995, n17996, n17997, n17998,
    n17999, n18000, n18001, n18002, n18003, n18004,
    n18005, n18006, n18007, n18008, n18009, n18010,
    n18011, n18012, n18013, n18014, n18015, n18016,
    n18017, n18018, n18019, n18020, n18021, n18022,
    n18023, n18024, n18025, n18026, n18027, n18028,
    n18029, n18030, n18031, n18032, n18033, n18034,
    n18035, n18036, n18037, n18038, n18039, n18040,
    n18041, n18042, n18043, n18044, n18045, n18046,
    n18047, n18048, n18049, n18050, n18051, n18052,
    n18053, n18054, n18055, n18056, n18057, n18058,
    n18059, n18060, n18061, n18062, n18063, n18064,
    n18065, n18066, n18067, n18068, n18069, n18070,
    n18071, n18072, n18073, n18074, n18075, n18076,
    n18077, n18078, n18079, n18080, n18081, n18082,
    n18083, n18084, n18085, n18086, n18087, n18088,
    n18089, n18090, n18091, n18092, n18093, n18094,
    n18095, n18096, n18097, n18098, n18099, n18100,
    n18101, n18102, n18103, n18104, n18105, n18106,
    n18107, n18108, n18109, n18110, n18111, n18112,
    n18113, n18114, n18115, n18116, n18117, n18118,
    n18119, n18120, n18121, n18122, n18123, n18124,
    n18125, n18126, n18127, n18128, n18129, n18130,
    n18131, n18132, n18133, n18134, n18135, n18136,
    n18137, n18138, n18139, n18140, n18141, n18142,
    n18143, n18144, n18145, n18146, n18147, n18148,
    n18149, n18150, n18151, n18152, n18153, n18154,
    n18155, n18156, n18157, n18158, n18159, n18160,
    n18161, n18162, n18163, n18164, n18165, n18166,
    n18167, n18168, n18169, n18170, n18171, n18172,
    n18173, n18174, n18175, n18176, n18177, n18178,
    n18179, n18180, n18181, n18182, n18183, n18184,
    n18185, n18186, n18187, n18188, n18189, n18190,
    n18191, n18192, n18193, n18194, n18195, n18196,
    n18197, n18198, n18199, n18200, n18201, n18202,
    n18203, n18204, n18205, n18206, n18207, n18208,
    n18209, n18210, n18211, n18212, n18213, n18214,
    n18215, n18216, n18217, n18218, n18219, n18220,
    n18221, n18222, n18223, n18224, n18225, n18226,
    n18227, n18228, n18229, n18230, n18231, n18232,
    n18233, n18234, n18235, n18236, n18237, n18238,
    n18239, n18240, n18241, n18242, n18243, n18244,
    n18245, n18246, n18247, n18248, n18249, n18250,
    n18251, n18252, n18253, n18254, n18255, n18256,
    n18257, n18258, n18259, n18260, n18261, n18262,
    n18263, n18264, n18265, n18266, n18267, n18268,
    n18269, n18270, n18271, n18272, n18273, n18274,
    n18275, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18283, n18284, n18285, n18286,
    n18287, n18288, n18289, n18290, n18291, n18292,
    n18293, n18294, n18295, n18296, n18297, n18298,
    n18299, n18300, n18301, n18302, n18303, n18304,
    n18305, n18306, n18307, n18308, n18309, n18310,
    n18311, n18312, n18313, n18314, n18315, n18316,
    n18317, n18318, n18319, n18320, n18321, n18322,
    n18323, n18324, n18325, n18326, n18327, n18328,
    n18329, n18330, n18331, n18332, n18333, n18334,
    n18335, n18336, n18337, n18338, n18339, n18340,
    n18341, n18342, n18343, n18344, n18345, n18346,
    n18347, n18348, n18349, n18350, n18351, n18352,
    n18353, n18354, n18355, n18356, n18357, n18358,
    n18359, n18360, n18361, n18362, n18363, n18364,
    n18365, n18366, n18367, n18368, n18369, n18370,
    n18371, n18372, n18373, n18374, n18375, n18376,
    n18377, n18378, n18379, n18380, n18381, n18382,
    n18383, n18384, n18385, n18386, n18387, n18388,
    n18389, n18390, n18391, n18392, n18393, n18394,
    n18395, n18396, n18397, n18398, n18399, n18400,
    n18401, n18402, n18403, n18404, n18405, n18406,
    n18407, n18408, n18409, n18410, n18411, n18412,
    n18413, n18414, n18415, n18416, n18417, n18418,
    n18419, n18420, n18421, n18422, n18423, n18424,
    n18425, n18426, n18427, n18428, n18429, n18430,
    n18431, n18432, n18433, n18434, n18435, n18436,
    n18437, n18439, n18440, n18441, n18442, n18443,
    n18444, n18445, n18446, n18447, n18448, n18449,
    n18450, n18451, n18452, n18453, n18454, n18455,
    n18456, n18457, n18458, n18459, n18460, n18461,
    n18462, n18463, n18464, n18465, n18466, n18467,
    n18468, n18469, n18470, n18471, n18472, n18473,
    n18474, n18475, n18476, n18477, n18478, n18479,
    n18480, n18481, n18482, n18483, n18484, n18485,
    n18486, n18487, n18488, n18489, n18490, n18491,
    n18492, n18493, n18494, n18495, n18496, n18497,
    n18498, n18499, n18500, n18501, n18502, n18503,
    n18504, n18505, n18506, n18507, n18508, n18509,
    n18510, n18511, n18512, n18513, n18514, n18515,
    n18516, n18517, n18518, n18519, n18520, n18521,
    n18522, n18523, n18524, n18525, n18526, n18527,
    n18528, n18529, n18530, n18531, n18532, n18533,
    n18534, n18535, n18536, n18537, n18538, n18539,
    n18540, n18541, n18542, n18543, n18544, n18545,
    n18546, n18547, n18548, n18549, n18550, n18551,
    n18552, n18553, n18554, n18555, n18556, n18557,
    n18558, n18559, n18560, n18561, n18562, n18563,
    n18564, n18565, n18566, n18567, n18568, n18569,
    n18570, n18571, n18572, n18573, n18574, n18575,
    n18576, n18577, n18578, n18579, n18580, n18581,
    n18582, n18583, n18584, n18585, n18586, n18587,
    n18588, n18589, n18590, n18591, n18592, n18593,
    n18594, n18595, n18596, n18597, n18598, n18599,
    n18600, n18601, n18602, n18603, n18604, n18605,
    n18606, n18607, n18608, n18609, n18610, n18611,
    n18612, n18613, n18614, n18615, n18616, n18617,
    n18618, n18619, n18620, n18621, n18622, n18623,
    n18624, n18625, n18626, n18627, n18628, n18629,
    n18630, n18631, n18632, n18633, n18634, n18635,
    n18636, n18637, n18638, n18639, n18640, n18641,
    n18642, n18643, n18644, n18645, n18646, n18647,
    n18648, n18649, n18650, n18651, n18652, n18653,
    n18654, n18655, n18656, n18657, n18658, n18659,
    n18660, n18661, n18662, n18663, n18664, n18665,
    n18666, n18667, n18668, n18669, n18670, n18671,
    n18672, n18673, n18674, n18675, n18676, n18677,
    n18678, n18679, n18680, n18681, n18682, n18683,
    n18684, n18685, n18686, n18687, n18688, n18689,
    n18690, n18691, n18692, n18693, n18694, n18695,
    n18696, n18697, n18698, n18699, n18700, n18701,
    n18702, n18703, n18704, n18705, n18706, n18707,
    n18708, n18709, n18710, n18711, n18712, n18713,
    n18714, n18715, n18716, n18717, n18718, n18719,
    n18720, n18721, n18722, n18723, n18724, n18725,
    n18726, n18727, n18728, n18729, n18730, n18731,
    n18732, n18733, n18734, n18735, n18736, n18737,
    n18738, n18739, n18740, n18741, n18742, n18743,
    n18744, n18745, n18746, n18747, n18748, n18749,
    n18750, n18751, n18752, n18753, n18754, n18755,
    n18756, n18757, n18758, n18759, n18760, n18761,
    n18762, n18763, n18764, n18765, n18766, n18767,
    n18768, n18769, n18770, n18771, n18772, n18773,
    n18774, n18775, n18776, n18777, n18778, n18779,
    n18780, n18781, n18782, n18783, n18784, n18785,
    n18786, n18787, n18788, n18789, n18790, n18791,
    n18792, n18793, n18794, n18795, n18796, n18797,
    n18798, n18799, n18800, n18801, n18802, n18803,
    n18804, n18805, n18806, n18807, n18808, n18809,
    n18810, n18811, n18812, n18813, n18814, n18815,
    n18816, n18817, n18818, n18819, n18820, n18821,
    n18822, n18823, n18824, n18825, n18826, n18827,
    n18828, n18829, n18830, n18831, n18832, n18833,
    n18834, n18835, n18836, n18837, n18838, n18839,
    n18840, n18841, n18842, n18843, n18844, n18845,
    n18846, n18847, n18848, n18849, n18850, n18851,
    n18852, n18853, n18854, n18855, n18856, n18857,
    n18858, n18859, n18860, n18861, n18862, n18863,
    n18864, n18865, n18866, n18867, n18868, n18869,
    n18870, n18871, n18872, n18873, n18874, n18875,
    n18876, n18877, n18878, n18879, n18880, n18881,
    n18882, n18883, n18884, n18885, n18886, n18887,
    n18888, n18889, n18890, n18891, n18892, n18893,
    n18894, n18895, n18896, n18897, n18898, n18899,
    n18900, n18901, n18902, n18903, n18904, n18905,
    n18906, n18907, n18908, n18909, n18910, n18911,
    n18912, n18913, n18914, n18915, n18916, n18917,
    n18918, n18919, n18920, n18921, n18922, n18923,
    n18924, n18925, n18926, n18927, n18928, n18929,
    n18930, n18931, n18932, n18933, n18934, n18935,
    n18936, n18937, n18938, n18939, n18940, n18941,
    n18942, n18943, n18944, n18945, n18946, n18947,
    n18948, n18949, n18950, n18951, n18952, n18953,
    n18954, n18955, n18956, n18957, n18958, n18959,
    n18960, n18961, n18962, n18963, n18964, n18965,
    n18966, n18967, n18968, n18969, n18970, n18971,
    n18972, n18973, n18974, n18975, n18976, n18977,
    n18978, n18979, n18980, n18981, n18982, n18983,
    n18984, n18985, n18986, n18987, n18988, n18989,
    n18990, n18991, n18992, n18993, n18994, n18995,
    n18996, n18997, n18998, n18999, n19000, n19001,
    n19002, n19003, n19004, n19005, n19006, n19007,
    n19008, n19009, n19010, n19011, n19012, n19013,
    n19014, n19015, n19016, n19017, n19018, n19019,
    n19020, n19021, n19022, n19023, n19024, n19025,
    n19026, n19027, n19028, n19029, n19030, n19031,
    n19032, n19033, n19034, n19035, n19036, n19037,
    n19038, n19039, n19040, n19041, n19042, n19043,
    n19044, n19045, n19046, n19047, n19048, n19049,
    n19050, n19051, n19052, n19053, n19054, n19055,
    n19056, n19057, n19058, n19059, n19060, n19061,
    n19062, n19063, n19064, n19065, n19066, n19067,
    n19068, n19069, n19070, n19071, n19072, n19073,
    n19074, n19075, n19076, n19077, n19078, n19079,
    n19080, n19081, n19082, n19083, n19084, n19085,
    n19086, n19087, n19088, n19089, n19090, n19091,
    n19092, n19093, n19094, n19095, n19096, n19097,
    n19098, n19099, n19100, n19101, n19102, n19103,
    n19104, n19105, n19106, n19107, n19108, n19109,
    n19110, n19111, n19112, n19113, n19114, n19115,
    n19116, n19117, n19118, n19119, n19120, n19121,
    n19122, n19123, n19124, n19125, n19126, n19127,
    n19128, n19129, n19130, n19131, n19132, n19133,
    n19134, n19135, n19136, n19137, n19138, n19139,
    n19140, n19141, n19142, n19143, n19144, n19145,
    n19146, n19147, n19148, n19149, n19150, n19151,
    n19152, n19153, n19154, n19155, n19156, n19157,
    n19158, n19159, n19160, n19161, n19162, n19163,
    n19164, n19165, n19166, n19167, n19168, n19169,
    n19170, n19171, n19172, n19173, n19174, n19175,
    n19176, n19177, n19178, n19179, n19180, n19181,
    n19182, n19183, n19184, n19185, n19186, n19187,
    n19188, n19189, n19190, n19191, n19192, n19193,
    n19194, n19195, n19196, n19197, n19198, n19199,
    n19200, n19201, n19202, n19203, n19204, n19205,
    n19206, n19207, n19208, n19209, n19210, n19211,
    n19213, n19214, n19215, n19216, n19217, n19218,
    n19219, n19220, n19221, n19222, n19223, n19224,
    n19225, n19226, n19227, n19228, n19229, n19230,
    n19231, n19232, n19233, n19234, n19235, n19236,
    n19237, n19238, n19239, n19240, n19241, n19242,
    n19243, n19244, n19245, n19246, n19247, n19248,
    n19249, n19250, n19251, n19252, n19253, n19254,
    n19255, n19256, n19257, n19258, n19259, n19260,
    n19261, n19262, n19263, n19264, n19265, n19266,
    n19267, n19268, n19269, n19270, n19271, n19272,
    n19273, n19274, n19275, n19276, n19277, n19278,
    n19279, n19280, n19281, n19282, n19283, n19284,
    n19285, n19286, n19287, n19288, n19289, n19290,
    n19291, n19292, n19293, n19294, n19295, n19296,
    n19297, n19298, n19299, n19300, n19301, n19302,
    n19303, n19304, n19305, n19306, n19307, n19308,
    n19309, n19310, n19311, n19312, n19313, n19314,
    n19315, n19316, n19317, n19318, n19319, n19320,
    n19321, n19322, n19323, n19324, n19325, n19326,
    n19327, n19328, n19329, n19330, n19331, n19332,
    n19333, n19334, n19335, n19336, n19337, n19338,
    n19339, n19340, n19341, n19342, n19343, n19344,
    n19345, n19346, n19347, n19348, n19349, n19350,
    n19351, n19352, n19353, n19354, n19355, n19356,
    n19357, n19358, n19359, n19360, n19361, n19362,
    n19363, n19364, n19365, n19366, n19367, n19368,
    n19369, n19370, n19371, n19372, n19373, n19374,
    n19375, n19376, n19377, n19378, n19379, n19380,
    n19381, n19382, n19383, n19384, n19385, n19386,
    n19387, n19388, n19389, n19390, n19391, n19392,
    n19393, n19394, n19395, n19396, n19397, n19398,
    n19399, n19400, n19401, n19402, n19403, n19404,
    n19405, n19406, n19407, n19408, n19409, n19410,
    n19411, n19412, n19413, n19414, n19415, n19416,
    n19417, n19418, n19419, n19420, n19421, n19422,
    n19423, n19424, n19425, n19426, n19427, n19428,
    n19429, n19430, n19431, n19432, n19433, n19434,
    n19435, n19436, n19437, n19438, n19439, n19440,
    n19441, n19442, n19443, n19444, n19445, n19446,
    n19447, n19448, n19449, n19450, n19451, n19452,
    n19453, n19454, n19455, n19456, n19457, n19458,
    n19459, n19460, n19461, n19462, n19463, n19464,
    n19465, n19466, n19467, n19468, n19469, n19470,
    n19471, n19472, n19473, n19474, n19475, n19476,
    n19477, n19478, n19479, n19480, n19481, n19482,
    n19483, n19484, n19485, n19486, n19487, n19488,
    n19489, n19490, n19491, n19492, n19493, n19494,
    n19495, n19496, n19497, n19498, n19499, n19500,
    n19501, n19502, n19503, n19504, n19505, n19506,
    n19507, n19508, n19509, n19510, n19511, n19512,
    n19513, n19514, n19515, n19516, n19517, n19518,
    n19519, n19520, n19521, n19522, n19523, n19524,
    n19525, n19526, n19527, n19528, n19529, n19530,
    n19531, n19532, n19533, n19534, n19535, n19536,
    n19537, n19538, n19539, n19540, n19541, n19542,
    n19543, n19544, n19545, n19546, n19547, n19548,
    n19549, n19550, n19551, n19552, n19553, n19554,
    n19555, n19556, n19557, n19558, n19559, n19560,
    n19561, n19562, n19563, n19564, n19565, n19566,
    n19567, n19568, n19569, n19570, n19571, n19572,
    n19573, n19574, n19575, n19576, n19577, n19578,
    n19579, n19580, n19581, n19582, n19583, n19584,
    n19585, n19586, n19587, n19588, n19589, n19590,
    n19591, n19592, n19593, n19594, n19595, n19596,
    n19597, n19598, n19599, n19600, n19601, n19602,
    n19603, n19604, n19605, n19606, n19607, n19608,
    n19609, n19610, n19611, n19612, n19613, n19614,
    n19615, n19616, n19617, n19618, n19619, n19620,
    n19621, n19622, n19623, n19624, n19625, n19626,
    n19627, n19628, n19629, n19630, n19631, n19632,
    n19633, n19634, n19635, n19636, n19637, n19638,
    n19639, n19640, n19641, n19642, n19643, n19644,
    n19645, n19646, n19647, n19648, n19649, n19650,
    n19651, n19652, n19653, n19654, n19655, n19656,
    n19657, n19658, n19659, n19660, n19661, n19662,
    n19663, n19664, n19665, n19666, n19667, n19668,
    n19669, n19670, n19671, n19672, n19673, n19674,
    n19675, n19676, n19677, n19678, n19679, n19680,
    n19681, n19682, n19683, n19684, n19685, n19686,
    n19687, n19688, n19689, n19690, n19691, n19692,
    n19693, n19694, n19695, n19696, n19697, n19698,
    n19699, n19700, n19701, n19702, n19703, n19704,
    n19705, n19706, n19707, n19708, n19709, n19710,
    n19711, n19712, n19713, n19714, n19715, n19716,
    n19717, n19718, n19719, n19720, n19721, n19722,
    n19723, n19724, n19725, n19726, n19727, n19728,
    n19729, n19730, n19731, n19732, n19733, n19734,
    n19735, n19736, n19737, n19739, n19740, n19741,
    n19742, n19743, n19744, n19745, n19746, n19747,
    n19748, n19749, n19750, n19751, n19752, n19753,
    n19754, n19755, n19756, n19757, n19758, n19759,
    n19760, n19761, n19762, n19763, n19764, n19765,
    n19766, n19767, n19768, n19769, n19770, n19771,
    n19772, n19773, n19774, n19775, n19776, n19777,
    n19778, n19779, n19780, n19781, n19782, n19783,
    n19784, n19785, n19786, n19787, n19788, n19789,
    n19790, n19791, n19792, n19793, n19794, n19795,
    n19796, n19797, n19798, n19799, n19800, n19801,
    n19802, n19803, n19804, n19805, n19806, n19807,
    n19808, n19809, n19810, n19811, n19812, n19813,
    n19814, n19815, n19816, n19817, n19818, n19819,
    n19820, n19821, n19822, n19823, n19824, n19825,
    n19826, n19827, n19828, n19829, n19830, n19831,
    n19832, n19833, n19834, n19835, n19836, n19837,
    n19838, n19839, n19840, n19841, n19842, n19843,
    n19844, n19845, n19846, n19847, n19848, n19849,
    n19850, n19851, n19852, n19853, n19854, n19855,
    n19856, n19857, n19858, n19859, n19860, n19861,
    n19862, n19863, n19864, n19865, n19866, n19867,
    n19868, n19869, n19870, n19871, n19872, n19873,
    n19874, n19875, n19876, n19877, n19878, n19879,
    n19880, n19881, n19882, n19883, n19884, n19885,
    n19886, n19887, n19888, n19889, n19890, n19891,
    n19892, n19893, n19894, n19895, n19896, n19897,
    n19898, n19899, n19900, n19901, n19902, n19903,
    n19904, n19905, n19906, n19907, n19908, n19909,
    n19910, n19911, n19912, n19913, n19914, n19915,
    n19916, n19917, n19918, n19919, n19920, n19921,
    n19922, n19923, n19924, n19925, n19926, n19927,
    n19928, n19929, n19930, n19931, n19932, n19933,
    n19934, n19935, n19936, n19937, n19938, n19939,
    n19940, n19941, n19942, n19943, n19944, n19945,
    n19946, n19947, n19948, n19949, n19950, n19951,
    n19952, n19953, n19954, n19955, n19956, n19957,
    n19958, n19959, n19960, n19961, n19962, n19963,
    n19964, n19965, n19966, n19967, n19968, n19969,
    n19970, n19971, n19972, n19973, n19974, n19975,
    n19976, n19977, n19978, n19979, n19980, n19981,
    n19982, n19983, n19984, n19985, n19986, n19987,
    n19988, n19989, n19990, n19991, n19992, n19993,
    n19994, n19995, n19996, n19997, n19998, n19999,
    n20000, n20001, n20002, n20003, n20004, n20005,
    n20006, n20007, n20008, n20009, n20010, n20011,
    n20012, n20013, n20014, n20015, n20016, n20017,
    n20018, n20019, n20020, n20021, n20022, n20023,
    n20024, n20025, n20026, n20027, n20028, n20029,
    n20030, n20031, n20032, n20033, n20034, n20035,
    n20036, n20037, n20038, n20039, n20040, n20041,
    n20042, n20043, n20044, n20045, n20046, n20047,
    n20048, n20049, n20050, n20051, n20052, n20053,
    n20054, n20055, n20056, n20057, n20058, n20059,
    n20060, n20061, n20062, n20063, n20064, n20065,
    n20066, n20067, n20068, n20069, n20070, n20071,
    n20072, n20073, n20074, n20075, n20076, n20077,
    n20078, n20079, n20080, n20081, n20082, n20083,
    n20084, n20085, n20086, n20087, n20088, n20089,
    n20090, n20091, n20092, n20093, n20094, n20095,
    n20096, n20097, n20098, n20099, n20100, n20101,
    n20102, n20103, n20104, n20105, n20106, n20107,
    n20108, n20109, n20110, n20111, n20112, n20113,
    n20114, n20115, n20116, n20117, n20118, n20119,
    n20120, n20121, n20122, n20123, n20124, n20125,
    n20126, n20127, n20128, n20129, n20130, n20131,
    n20132, n20133, n20134, n20135, n20136, n20137,
    n20138, n20139, n20140, n20141, n20142, n20143,
    n20144, n20145, n20146, n20147, n20148, n20149,
    n20150, n20151, n20152, n20153, n20154, n20155,
    n20156, n20157, n20158, n20159, n20160, n20161,
    n20162, n20163, n20164, n20165, n20166, n20167,
    n20168, n20169, n20170, n20171, n20172, n20173,
    n20174, n20175, n20176, n20177, n20178, n20179,
    n20180, n20181, n20182, n20183, n20184, n20185,
    n20186, n20187, n20188, n20189, n20190, n20191,
    n20192, n20193, n20194, n20195, n20196, n20197,
    n20198, n20199, n20200, n20201, n20202, n20203,
    n20204, n20205, n20206, n20207, n20208, n20209,
    n20210, n20211, n20212, n20213, n20214, n20215,
    n20216, n20217, n20218, n20219, n20220, n20221,
    n20222, n20223, n20224, n20225, n20226, n20227,
    n20228, n20229, n20230, n20231, n20232, n20233,
    n20234, n20235, n20236, n20237, n20238, n20239,
    n20240, n20241, n20242, n20243, n20244, n20245,
    n20246, n20247, n20248, n20249, n20250, n20251,
    n20253, n20254, n20255, n20256, n20257, n20258,
    n20259, n20260, n20261, n20262, n20263, n20264,
    n20265, n20266, n20267, n20268, n20269, n20270,
    n20271, n20272, n20273, n20274, n20275, n20276,
    n20277, n20278, n20279, n20280, n20281, n20282,
    n20283, n20284, n20285, n20286, n20287, n20288,
    n20289, n20290, n20291, n20292, n20293, n20294,
    n20295, n20296, n20297, n20298, n20299, n20300,
    n20301, n20302, n20303, n20304, n20305, n20306,
    n20307, n20308, n20309, n20310, n20311, n20312,
    n20313, n20314, n20315, n20316, n20317, n20318,
    n20319, n20320, n20321, n20322, n20323, n20324,
    n20325, n20326, n20327, n20328, n20329, n20330,
    n20331, n20332, n20333, n20334, n20335, n20336,
    n20337, n20338, n20339, n20340, n20341, n20342,
    n20343, n20344, n20345, n20346, n20347, n20348,
    n20349, n20350, n20351, n20352, n20353, n20354,
    n20355, n20356, n20357, n20358, n20359, n20360,
    n20361, n20362, n20363, n20364, n20365, n20366,
    n20367, n20368, n20369, n20370, n20371, n20372,
    n20373, n20374, n20375, n20376, n20377, n20378,
    n20379, n20380, n20381, n20382, n20383, n20384,
    n20385, n20386, n20387, n20388, n20389, n20390,
    n20391, n20392, n20393, n20394, n20395, n20396,
    n20397, n20398, n20399, n20400, n20401, n20402,
    n20403, n20404, n20405, n20406, n20407, n20408,
    n20409, n20410, n20411, n20412, n20413, n20414,
    n20415, n20416, n20417, n20418, n20419, n20420,
    n20421, n20422, n20423, n20424, n20425, n20426,
    n20427, n20428, n20429, n20430, n20431, n20432,
    n20433, n20434, n20435, n20436, n20437, n20438,
    n20439, n20440, n20441, n20442, n20443, n20444,
    n20445, n20446, n20447, n20448, n20449, n20450,
    n20451, n20452, n20453, n20454, n20455, n20456,
    n20457, n20458, n20459, n20460, n20461, n20462,
    n20463, n20464, n20465, n20466, n20467, n20468,
    n20469, n20470, n20471, n20472, n20473, n20474,
    n20475, n20476, n20477, n20478, n20479, n20480,
    n20481, n20482, n20483, n20484, n20485, n20486,
    n20487, n20488, n20489, n20490, n20491, n20492,
    n20493, n20494, n20495, n20496, n20497, n20498,
    n20499, n20500, n20501, n20502, n20503, n20504,
    n20505, n20506, n20507, n20508, n20509, n20510,
    n20511, n20512, n20513, n20514, n20515, n20516,
    n20517, n20518, n20519, n20520, n20521, n20522,
    n20523, n20524, n20525, n20526, n20527, n20528,
    n20529, n20530, n20531, n20532, n20533, n20534,
    n20535, n20536, n20537, n20538, n20539, n20540,
    n20541, n20542, n20543, n20544, n20545, n20546,
    n20547, n20548, n20549, n20550, n20551, n20552,
    n20553, n20554, n20555, n20556, n20557, n20558,
    n20559, n20560, n20561, n20562, n20563, n20564,
    n20565, n20566, n20567, n20568, n20569, n20570,
    n20571, n20572, n20573, n20574, n20575, n20576,
    n20577, n20578, n20579, n20580, n20581, n20582,
    n20583, n20584, n20585, n20586, n20587, n20588,
    n20589, n20590, n20591, n20592, n20593, n20594,
    n20595, n20596, n20597, n20598, n20599, n20600,
    n20601, n20602, n20603, n20604, n20605, n20606,
    n20607, n20608, n20609, n20610, n20611, n20612,
    n20613, n20614, n20615, n20616, n20617, n20618,
    n20619, n20620, n20621, n20622, n20623, n20624,
    n20625, n20626, n20627, n20628, n20629, n20630,
    n20631, n20632, n20633, n20634, n20635, n20636,
    n20637, n20638, n20639, n20640, n20641, n20642,
    n20643, n20644, n20645, n20646, n20647, n20648,
    n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20658, n20659, n20660,
    n20661, n20662, n20663, n20664, n20665, n20666,
    n20667, n20668, n20669, n20670, n20671, n20672,
    n20673, n20674, n20675, n20676, n20677, n20678,
    n20679, n20680, n20681, n20682, n20683, n20684,
    n20685, n20686, n20687, n20688, n20689, n20690,
    n20691, n20692, n20693, n20694, n20695, n20696,
    n20697, n20698, n20699, n20700, n20701, n20702,
    n20703, n20704, n20705, n20706, n20707, n20708,
    n20709, n20710, n20711, n20712, n20713, n20714,
    n20715, n20716, n20717, n20718, n20719, n20720,
    n20721, n20722, n20723, n20724, n20725, n20726,
    n20727, n20728, n20729, n20730, n20731, n20732,
    n20733, n20734, n20735, n20736, n20737, n20739,
    n20740, n20741, n20742, n20743, n20744, n20745,
    n20746, n20747, n20748, n20749, n20750, n20751,
    n20752, n20753, n20754, n20755, n20756, n20757,
    n20758, n20759, n20760, n20761, n20762, n20763,
    n20764, n20765, n20766, n20767, n20768, n20769,
    n20770, n20771, n20772, n20773, n20774, n20775,
    n20776, n20777, n20778, n20779, n20780, n20781,
    n20782, n20783, n20784, n20785, n20786, n20787,
    n20788, n20789, n20790, n20791, n20792, n20793,
    n20794, n20795, n20796, n20797, n20798, n20799,
    n20800, n20801, n20802, n20803, n20804, n20805,
    n20806, n20807, n20808, n20809, n20810, n20811,
    n20812, n20813, n20814, n20815, n20816, n20817,
    n20818, n20820, n20821, n20822, n20823, n20824,
    n20825, n20826, n20827, n20828, n20829, n20830,
    n20831, n20832, n20833, n20834, n20835, n20836,
    n20837, n20838, n20839, n20840, n20841, n20842,
    n20843, n20844, n20845, n20846, n20847, n20848,
    n20849, n20850, n20851, n20852, n20853, n20854,
    n20855, n20856, n20857, n20858, n20859, n20860,
    n20861, n20862, n20863, n20864, n20865, n20866,
    n20867, n20868, n20869, n20870, n20871, n20872,
    n20873, n20874, n20875, n20876, n20877, n20878,
    n20879, n20880, n20881, n20882, n20883, n20884,
    n20885, n20886, n20887, n20888, n20889, n20890,
    n20891, n20892, n20893, n20894, n20895, n20896,
    n20897, n20898, n20899, n20900, n20901, n20902,
    n20903, n20904, n20905, n20906, n20907, n20908,
    n20909, n20910, n20911, n20912, n20913, n20914,
    n20915, n20916, n20917, n20918, n20919, n20920,
    n20921, n20922, n20923, n20924, n20925, n20926,
    n20927, n20928, n20929, n20930, n20931, n20932,
    n20933, n20934, n20935, n20936, n20937, n20938,
    n20939, n20940, n20941, n20942, n20943, n20944,
    n20945, n20946, n20947, n20948, n20949, n20950,
    n20951, n20952, n20953, n20954, n20955, n20956,
    n20957, n20959, n20960, n20961, n20962, n20963,
    n20964, n20965, n20966, n20967, n20968, n20969,
    n20970, n20971, n20972, n20973, n20974, n20975,
    n20976, n20977, n20978, n20979, n20980, n20981,
    n20982, n20983, n20984, n20985, n20986, n20987,
    n20988, n20989, n20990, n20991, n20992, n20993,
    n20994, n20995, n20996, n20997, n20998, n20999,
    n21000, n21001, n21002, n21003, n21004, n21005,
    n21006, n21007, n21008, n21009, n21010, n21011,
    n21012, n21013, n21014, n21015, n21016, n21017,
    n21018, n21019, n21020, n21021, n21023, n21024,
    n21025, n21026, n21027, n21028, n21029, n21030,
    n21031, n21032, n21033, n21034, n21035, n21036,
    n21037, n21038, n21039, n21040, n21041, n21042,
    n21043, n21044, n21045, n21046, n21047, n21048,
    n21049, n21050, n21051, n21052, n21053, n21054,
    n21055, n21056, n21057, n21058, n21059, n21060,
    n21061, n21062, n21063, n21064, n21065, n21066,
    n21067, n21068, n21069, n21070, n21071, n21072,
    n21073, n21074, n21075, n21076, n21077, n21078,
    n21079, n21080, n21082, n21083, n21084, n21085,
    n21086, n21087, n21088, n21089, n21090, n21091,
    n21092, n21093, n21094, n21095, n21096, n21097,
    n21098, n21099, n21100, n21101, n21102, n21103,
    n21104, n21105, n21106, n21107, n21108, n21109,
    n21110, n21111, n21112, n21113, n21114, n21115,
    n21116, n21117, n21118, n21119, n21120, n21121,
    n21122, n21123, n21124, n21125, n21126, n21127,
    n21128, n21129, n21130, n21131, n21132, n21133,
    n21134, n21135, n21136, n21138, n21139, n21140,
    n21141, n21142, n21143, n21144, n21145, n21146,
    n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158,
    n21159, n21160, n21161, n21162, n21163, n21164,
    n21165, n21166, n21167, n21168, n21169, n21170,
    n21171, n21172, n21173, n21174, n21175, n21176,
    n21177, n21178, n21179, n21180, n21181, n21182,
    n21183, n21184, n21185, n21186, n21187, n21188,
    n21189, n21190, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200,
    n21201, n21202, n21203, n21204, n21205, n21206,
    n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21216, n21217, n21218, n21219,
    n21220, n21221, n21222, n21223, n21224, n21225,
    n21226, n21227, n21228, n21229, n21230, n21231,
    n21232, n21233, n21234, n21235, n21236, n21237,
    n21238, n21239, n21240, n21241, n21242, n21243,
    n21244, n21245, n21246, n21247, n21248, n21249,
    n21250, n21251, n21252, n21253, n21254, n21255,
    n21256, n21257, n21258, n21259, n21260, n21261,
    n21262, n21263, n21264, n21265, n21266, n21267,
    n21268, n21269, n21270, n21271, n21272, n21273,
    n21274, n21275, n21276, n21277, n21278, n21279,
    n21280, n21281, n21282, n21283, n21284, n21285,
    n21286, n21287, n21288, n21289, n21290, n21291,
    n21292, n21293, n21294, n21295, n21296, n21297,
    n21298, n21299, n21300, n21301, n21302, n21303,
    n21304, n21305, n21306, n21307, n21308, n21309,
    n21310, n21311, n21312, n21313, n21314, n21315,
    n21316, n21317, n21318, n21319, n21320, n21321,
    n21323, n21324, n21325, n21326, n21327, n21328,
    n21329, n21330, n21331, n21332, n21333, n21334,
    n21335, n21336, n21337, n21338, n21339, n21340,
    n21341, n21342, n21343, n21344, n21345, n21346,
    n21347, n21348, n21349, n21350, n21351, n21352,
    n21353, n21354, n21355, n21356, n21357, n21358,
    n21359, n21360, n21361, n21362, n21363, n21364,
    n21365, n21366, n21367, n21368, n21369, n21370,
    n21371, n21372, n21373, n21374, n21375, n21376,
    n21377, n21378, n21379, n21380, n21381, n21382,
    n21383, n21384, n21385, n21386, n21387, n21388,
    n21389, n21390, n21391, n21392, n21393, n21394,
    n21395, n21396, n21397, n21398, n21399, n21400,
    n21401, n21402, n21404, n21405, n21406, n21407,
    n21408, n21409, n21410, n21411, n21412, n21413,
    n21414, n21415, n21416, n21417, n21418, n21419,
    n21420, n21421, n21422, n21423, n21424, n21425,
    n21426, n21427, n21428, n21429, n21430, n21431,
    n21432, n21433, n21434, n21435, n21436, n21437,
    n21438, n21439, n21440, n21441, n21442, n21443,
    n21444, n21445, n21446, n21447, n21448, n21449,
    n21450, n21451, n21452, n21453, n21454, n21456,
    n21457, n21458, n21459, n21460, n21461, n21462,
    n21463, n21464, n21465, n21466, n21467, n21468,
    n21469, n21470, n21471, n21472, n21473, n21474,
    n21475, n21476, n21477, n21478, n21479, n21480,
    n21481, n21482, n21483, n21484, n21485, n21486,
    n21487, n21488, n21489, n21490, n21491, n21492,
    n21493, n21494, n21496, n21497, n21498, n21499,
    n21500, n21501, n21502, n21503, n21504, n21505,
    n21506, n21507, n21508, n21509, n21510, n21511,
    n21512, n21513, n21514, n21515, n21516, n21517,
    n21518, n21519, n21520, n21521, n21522, n21523,
    n21524, n21526, n21527, n21528, n21529, n21530,
    n21531, n21532, n21533, n21534, n21535, n21536,
    n21537, n21538, n21539, n21540, n21541, n21542,
    n21543, n21544, n21545, n21546, n21547, n21548,
    n21549, n21550, n21551, n21552, n21553, n21554,
    n21555, n21556, n21557, n21558, n21559, n21560,
    n21561, n21562, n21563, n21564, n21565, n21566,
    n21567, n21568, n21569, n21570, n21571, n21572,
    n21573, n21574, n21575, n21576, n21577, n21578,
    n21579, n21580, n21581, n21583, n21584, n21585,
    n21586, n21587, n21588, n21589, n21590, n21591,
    n21592, n21593, n21594, n21595, n21596, n21597,
    n21598, n21599, n21600, n21601, n21602, n21603,
    n21604, n21605, n21606, n21607, n21608, n21609,
    n21610, n21611, n21612, n21613, n21614, n21615,
    n21616, n21617, n21618, n21619, n21620, n21621,
    n21622, n21623, n21624, n21625, n21626, n21627,
    n21628, n21629, n21630, n21631, n21632, n21633,
    n21634, n21635, n21636, n21637, n21639, n21640,
    n21641, n21642, n21643, n21644, n21645, n21646,
    n21647, n21648, n21649, n21650, n21651, n21652,
    n21653, n21654, n21655, n21656, n21657, n21658,
    n21659, n21660, n21661, n21662, n21663, n21664,
    n21665, n21666, n21667, n21668, n21669, n21670,
    n21671, n21672, n21673, n21674, n21675, n21676,
    n21677, n21678, n21679, n21680, n21681, n21682,
    n21683, n21684, n21685, n21686, n21687, n21688,
    n21689, n21690, n21691, n21692, n21693, n21695,
    n21696, n21697, n21698, n21699, n21700, n21701,
    n21702, n21703, n21704, n21705, n21706, n21707,
    n21708, n21709, n21710, n21711, n21712, n21713,
    n21714, n21715, n21716, n21717, n21718, n21719,
    n21720, n21721, n21722, n21723, n21724, n21725,
    n21726, n21727, n21728, n21729, n21730, n21731,
    n21732, n21733, n21734, n21735, n21736, n21737,
    n21738, n21739, n21740, n21741, n21742, n21743,
    n21744, n21745, n21746, n21747, n21748, n21749,
    n21750, n21751, n21752, n21754, n21755, n21756,
    n21757, n21758, n21759, n21760, n21761, n21762,
    n21763, n21764, n21765, n21766, n21767, n21768,
    n21769, n21770, n21771, n21772, n21773, n21774,
    n21775, n21776, n21777, n21778, n21779, n21780,
    n21781, n21782, n21783, n21784, n21785, n21786,
    n21787, n21788, n21789, n21790, n21791, n21792,
    n21793, n21794, n21795, n21796, n21797, n21798,
    n21799, n21800, n21801, n21802, n21803, n21804,
    n21805, n21806, n21807, n21808, n21809, n21810,
    n21811, n21812, n21813, n21814, n21815, n21816,
    n21817, n21818, n21819, n21820, n21821, n21822,
    n21823, n21824, n21825, n21826, n21827, n21828,
    n21829, n21830, n21831, n21832, n21833, n21834,
    n21835, n21836, n21837, n21838, n21839, n21840,
    n21841, n21842, n21843, n21844, n21845, n21846,
    n21848, n21849, n21850, n21851, n21852, n21853,
    n21854, n21855, n21856, n21857, n21858, n21859,
    n21860, n21861, n21862, n21863, n21864, n21865,
    n21866, n21867, n21868, n21869, n21870, n21871,
    n21872, n21873, n21874, n21875, n21876, n21877,
    n21878, n21879, n21880, n21881, n21882, n21883,
    n21884, n21885, n21886, n21887, n21888, n21889,
    n21890, n21891, n21892, n21893, n21894, n21895,
    n21896, n21897, n21898, n21899, n21900, n21901,
    n21903, n21904, n21905, n21906, n21907, n21908,
    n21909, n21910, n21911, n21912, n21913, n21914,
    n21915, n21916, n21917, n21918, n21919, n21920,
    n21921, n21922, n21923, n21924, n21925, n21926,
    n21927, n21928, n21929, n21930, n21931, n21932,
    n21933, n21934, n21935, n21936, n21937, n21938,
    n21939, n21940, n21941, n21942, n21943, n21944,
    n21945, n21946, n21947, n21948, n21949, n21950,
    n21951, n21952, n21953, n21954, n21955, n21956,
    n21957, n21958, n21959, n21961, n21962, n21963,
    n21964, n21965, n21966, n21967, n21968, n21969,
    n21970, n21971, n21972, n21973, n21974, n21975,
    n21976, n21977, n21978, n21979, n21980, n21981,
    n21982, n21983, n21984, n21985, n21986, n21987,
    n21988, n21989, n21990, n21991, n21992, n21993,
    n21994, n21995, n21996, n21997, n21998, n21999,
    n22001, n22002, n22003, n22004, n22005, n22006,
    n22007, n22008, n22009, n22010, n22011, n22012,
    n22013, n22014, n22015, n22016, n22017, n22018,
    n22019, n22020, n22021, n22022, n22023, n22024,
    n22025, n22026, n22027, n22028, n22029, n22030,
    n22031, n22032, n22033, n22034, n22035, n22036,
    n22037, n22038, n22039, n22041, n22042, n22043,
    n22044, n22045, n22046, n22047, n22048, n22049,
    n22050, n22051, n22052, n22053, n22054, n22055,
    n22056, n22057, n22058, n22059, n22060, n22061,
    n22062, n22063, n22064, n22065, n22066, n22067,
    n22068, n22069, n22070, n22071, n22072, n22073,
    n22074, n22075, n22076, n22077, n22078, n22079,
    n22080, n22081, n22082, n22083, n22084, n22085,
    n22086, n22087, n22088, n22089, n22090, n22091,
    n22092, n22093, n22094, n22095, n22096, n22097,
    n22098, n22099, n22100, n22101, n22102, n22103,
    n22104, n22105, n22106, n22107, n22108, n22109,
    n22110, n22111, n22112, n22113, n22114, n22115,
    n22116, n22117, n22118, n22119, n22120, n22121,
    n22122, n22123, n22124, n22125, n22126, n22127,
    n22128, n22129, n22130, n22131, n22132, n22133,
    n22134, n22135, n22136, n22138, n22139, n22140,
    n22141, n22142, n22143, n22144, n22145, n22146,
    n22147, n22148, n22149, n22150, n22151, n22152,
    n22153, n22154, n22155, n22156, n22157, n22158,
    n22159, n22160, n22161, n22162, n22163, n22164,
    n22165, n22166, n22167, n22168, n22169, n22170,
    n22171, n22172, n22173, n22174, n22175, n22176,
    n22177, n22178, n22179, n22181, n22182, n22183,
    n22184, n22185, n22186, n22187, n22188, n22189,
    n22190, n22191, n22192, n22193, n22194, n22195,
    n22196, n22197, n22198, n22199, n22200, n22201,
    n22202, n22203, n22204, n22205, n22206, n22207,
    n22208, n22209, n22210, n22211, n22212, n22213,
    n22214, n22215, n22216, n22217, n22218, n22219,
    n22220, n22221, n22222, n22223, n22224, n22225,
    n22226, n22227, n22228, n22229, n22230, n22231,
    n22232, n22233, n22234, n22235, n22236, n22237,
    n22238, n22239, n22240, n22241, n22242, n22243,
    n22244, n22245, n22246, n22247, n22248, n22249,
    n22250, n22251, n22252, n22253, n22254, n22255,
    n22256, n22257, n22258, n22259, n22260, n22262,
    n22263, n22264, n22265, n22266, n22267, n22268,
    n22269, n22270, n22271, n22272, n22273, n22274,
    n22275, n22276, n22277, n22278, n22279, n22280,
    n22281, n22282, n22283, n22284, n22285, n22286,
    n22287, n22288, n22289, n22290, n22291, n22292,
    n22293, n22294, n22295, n22296, n22297, n22298,
    n22299, n22300, n22301, n22302, n22303, n22304,
    n22305, n22306, n22307, n22308, n22309, n22310,
    n22311, n22312, n22313, n22314, n22315, n22316,
    n22317, n22318, n22319, n22320, n22321, n22322,
    n22323, n22324, n22325, n22326, n22327, n22328,
    n22329, n22330, n22331, n22332, n22333, n22334,
    n22335, n22336, n22337, n22338, n22339, n22340,
    n22341, n22343, n22344, n22345, n22346, n22347,
    n22348, n22349, n22350, n22351, n22352, n22353,
    n22354, n22355, n22356, n22357, n22358, n22359,
    n22360, n22361, n22362, n22363, n22364, n22365,
    n22366, n22367, n22368, n22369, n22370, n22371,
    n22372, n22373, n22374, n22375, n22376, n22377,
    n22378, n22379, n22380, n22381, n22382, n22383,
    n22384, n22385, n22386, n22387, n22388, n22389,
    n22390, n22391, n22392, n22393, n22394, n22395,
    n22396, n22397, n22398, n22399, n22400, n22401,
    n22402, n22403, n22404, n22405, n22406, n22407,
    n22408, n22409, n22410, n22411, n22412, n22413,
    n22414, n22415, n22416, n22417, n22418, n22419,
    n22420, n22421, n22423, n22424, n22425, n22426,
    n22427, n22428, n22429, n22430, n22431, n22432,
    n22433, n22434, n22435, n22436, n22437, n22438,
    n22439, n22440, n22441, n22442, n22443, n22444,
    n22445, n22446, n22447, n22448, n22449, n22450,
    n22451, n22452, n22453, n22454, n22455, n22456,
    n22457, n22458, n22459, n22460, n22461, n22462,
    n22463, n22464, n22465, n22466, n22467, n22468,
    n22469, n22470, n22471, n22472, n22473, n22474,
    n22475, n22476, n22477, n22478, n22479, n22480,
    n22481, n22482, n22483, n22484, n22485, n22486,
    n22487, n22488, n22489, n22490, n22491, n22492,
    n22493, n22494, n22495, n22496, n22497, n22498,
    n22499, n22500, n22501, n22502, n22504, n22505,
    n22506, n22507, n22508, n22509, n22510, n22511,
    n22512, n22513, n22514, n22515, n22516, n22517,
    n22518, n22519, n22520, n22521, n22522, n22523,
    n22524, n22525, n22526, n22527, n22528, n22529,
    n22530, n22531, n22532, n22533, n22534, n22535,
    n22536, n22537, n22538, n22539, n22540, n22541,
    n22542, n22543, n22544, n22545, n22546, n22547,
    n22548, n22549, n22550, n22551, n22552, n22553,
    n22554, n22555, n22556, n22557, n22558, n22559,
    n22560, n22561, n22562, n22563, n22564, n22565,
    n22566, n22567, n22568, n22569, n22570, n22571,
    n22572, n22573, n22574, n22575, n22576, n22577,
    n22578, n22579, n22580, n22581, n22582, n22583,
    n22585, n22586, n22587, n22588, n22589, n22590,
    n22591, n22592, n22593, n22594, n22595, n22596,
    n22597, n22598, n22599, n22600, n22601, n22602,
    n22603, n22604, n22605, n22606, n22607, n22608,
    n22609, n22610, n22611, n22612, n22613, n22614,
    n22615, n22616, n22617, n22618, n22619, n22620,
    n22621, n22622, n22623, n22624, n22625, n22626,
    n22627, n22628, n22629, n22630, n22631, n22632,
    n22633, n22634, n22635, n22636, n22637, n22638,
    n22639, n22640, n22641, n22642, n22643, n22644,
    n22645, n22646, n22647, n22648, n22649, n22650,
    n22651, n22652, n22653, n22654, n22655, n22656,
    n22657, n22658, n22659, n22660, n22661, n22662,
    n22663, n22664, n22665, n22666, n22667, n22668,
    n22669, n22670, n22671, n22672, n22673, n22674,
    n22675, n22676, n22677, n22678, n22679, n22680,
    n22681, n22682, n22683, n22684, n22685, n22686,
    n22687, n22688, n22689, n22690, n22691, n22692,
    n22693, n22694, n22695, n22696, n22697, n22698,
    n22699, n22700, n22701, n22702, n22703, n22704,
    n22705, n22706, n22707, n22708, n22709, n22710,
    n22711, n22712, n22713, n22714, n22715, n22716,
    n22717, n22718, n22719, n22720, n22721, n22722,
    n22723, n22724, n22725, n22726, n22727, n22728,
    n22729, n22730, n22731, n22732, n22733, n22734,
    n22735, n22736, n22737, n22738, n22739, n22740,
    n22741, n22742, n22743, n22744, n22745, n22746,
    n22747, n22748, n22749, n22750, n22751, n22752,
    n22753, n22754, n22755, n22756, n22757, n22758,
    n22759, n22760, n22761, n22762, n22763, n22764,
    n22765, n22766, n22767, n22768, n22769, n22770,
    n22771, n22772, n22773, n22774, n22775, n22776,
    n22777, n22778, n22779, n22780, n22781, n22782,
    n22783, n22784, n22785, n22786, n22787, n22788,
    n22789, n22790, n22791, n22792, n22793, n22794,
    n22795, n22796, n22797, n22798, n22799, n22800,
    n22801, n22802, n22803, n22804, n22805, n22806,
    n22807, n22808, n22809, n22810, n22811, n22812,
    n22813, n22814, n22815, n22816, n22817, n22818,
    n22819, n22820, n22821, n22822, n22823, n22824,
    n22825, n22826, n22827, n22828, n22829, n22830,
    n22831, n22832, n22833, n22834, n22835, n22836,
    n22837, n22838, n22839, n22840, n22841, n22842,
    n22843, n22844, n22845, n22846, n22847, n22848,
    n22849, n22850, n22851, n22852, n22853, n22854,
    n22855, n22856, n22857, n22858, n22859, n22860,
    n22861, n22862, n22863, n22864, n22865, n22866,
    n22867, n22868, n22869, n22870, n22871, n22872,
    n22873, n22874, n22875, n22876, n22877, n22878,
    n22879, n22880, n22881, n22882, n22883, n22884,
    n22885, n22886, n22887, n22888, n22889, n22890,
    n22891, n22892, n22893, n22894, n22895, n22896,
    n22897, n22898, n22899, n22900, n22901, n22902,
    n22903, n22904, n22905, n22906, n22907, n22908,
    n22909, n22910, n22911, n22912, n22913, n22914,
    n22915, n22916, n22917, n22918, n22919, n22920,
    n22921, n22922, n22923, n22924, n22925, n22926,
    n22927, n22928, n22929, n22930, n22931, n22932,
    n22933, n22934, n22935, n22936, n22937, n22938,
    n22939, n22940, n22941, n22942, n22943, n22944,
    n22945, n22946, n22947, n22948, n22949, n22950,
    n22951, n22952, n22953, n22954, n22955, n22956,
    n22957, n22958, n22959, n22960, n22961, n22962,
    n22963, n22964, n22965, n22966, n22967, n22968,
    n22969, n22970, n22971, n22972, n22973, n22974,
    n22975, n22976, n22977, n22978, n22979, n22980,
    n22981, n22982, n22983, n22984, n22985, n22986,
    n22987, n22988, n22989, n22990, n22991, n22992,
    n22993, n22994, n22995, n22996, n22997, n22998,
    n22999, n23000, n23001, n23002, n23003, n23004,
    n23005, n23006, n23007, n23008, n23009, n23010,
    n23011, n23012, n23013, n23014, n23015, n23016,
    n23017, n23018, n23019, n23020, n23021, n23022,
    n23023, n23024, n23025, n23026, n23027, n23028,
    n23029, n23030, n23031, n23032, n23033, n23034,
    n23035, n23036, n23037, n23038, n23039, n23040,
    n23041, n23042, n23043, n23044, n23045, n23046,
    n23047, n23048, n23049, n23050, n23051, n23052,
    n23053, n23054, n23055, n23056, n23058, n23059,
    n23060, n23061, n23062, n23063, n23064, n23065,
    n23066, n23067, n23068, n23069, n23070, n23071,
    n23072, n23073, n23074, n23075, n23076, n23077,
    n23078, n23079, n23080, n23081, n23082, n23083,
    n23084, n23085, n23086, n23087, n23088, n23089,
    n23090, n23091, n23092, n23093, n23094, n23095,
    n23096, n23097, n23098, n23099, n23100, n23101,
    n23102, n23103, n23104, n23105, n23106, n23107,
    n23108, n23109, n23110, n23111, n23112, n23113,
    n23114, n23115, n23116, n23117, n23118, n23119,
    n23120, n23121, n23122, n23123, n23124, n23125,
    n23126, n23127, n23128, n23129, n23130, n23131,
    n23132, n23133, n23134, n23135, n23136, n23137,
    n23138, n23139, n23140, n23141, n23142, n23143,
    n23144, n23145, n23146, n23147, n23148, n23149,
    n23150, n23151, n23152, n23153, n23154, n23155,
    n23156, n23157, n23158, n23159, n23160, n23161,
    n23162, n23163, n23164, n23165, n23166, n23167,
    n23168, n23169, n23170, n23171, n23172, n23173,
    n23174, n23175, n23176, n23177, n23178, n23179,
    n23180, n23181, n23182, n23183, n23184, n23185,
    n23186, n23187, n23188, n23189, n23190, n23191,
    n23192, n23193, n23194, n23195, n23196, n23197,
    n23198, n23199, n23200, n23201, n23202, n23203,
    n23204, n23205, n23206, n23207, n23208, n23209,
    n23210, n23211, n23212, n23213, n23214, n23215,
    n23216, n23217, n23218, n23219, n23220, n23221,
    n23222, n23223, n23224, n23225, n23226, n23227,
    n23228, n23229, n23230, n23231, n23232, n23233,
    n23234, n23235, n23236, n23237, n23238, n23239,
    n23240, n23241, n23242, n23243, n23244, n23245,
    n23246, n23247, n23248, n23249, n23250, n23251,
    n23252, n23253, n23254, n23255, n23256, n23257,
    n23258, n23259, n23260, n23261, n23262, n23263,
    n23264, n23265, n23266, n23267, n23268, n23269,
    n23270, n23271, n23272, n23273, n23274, n23275,
    n23276, n23277, n23278, n23279, n23280, n23281,
    n23282, n23283, n23284, n23285, n23286, n23287,
    n23288, n23289, n23290, n23291, n23292, n23293,
    n23294, n23295, n23296, n23297, n23298, n23299,
    n23300, n23301, n23302, n23303, n23304, n23305,
    n23306, n23307, n23308, n23309, n23310, n23311,
    n23312, n23313, n23314, n23315, n23316, n23317,
    n23318, n23319, n23320, n23321, n23322, n23323,
    n23324, n23325, n23326, n23327, n23328, n23329,
    n23330, n23331, n23332, n23333, n23334, n23335,
    n23336, n23337, n23338, n23339, n23340, n23341,
    n23342, n23343, n23344, n23345, n23346, n23347,
    n23348, n23349, n23350, n23351, n23352, n23353,
    n23354, n23355, n23356, n23357, n23358, n23359,
    n23360, n23361, n23362, n23363, n23364, n23365,
    n23366, n23367, n23368, n23369, n23370, n23371,
    n23372, n23373, n23374, n23375, n23376, n23377,
    n23378, n23379, n23380, n23381, n23382, n23383,
    n23384, n23385, n23386, n23387, n23388, n23389,
    n23390, n23391, n23392, n23393, n23394, n23395,
    n23396, n23397, n23398, n23399, n23400, n23401,
    n23402, n23403, n23404, n23405, n23406, n23407,
    n23408, n23409, n23410, n23411, n23412, n23413,
    n23414, n23415, n23416, n23417, n23418, n23419,
    n23420, n23421, n23422, n23423, n23424, n23425,
    n23426, n23427, n23428, n23429, n23430, n23431,
    n23432, n23433, n23434, n23435, n23436, n23437,
    n23438, n23439, n23440, n23441, n23442, n23443,
    n23444, n23445, n23446, n23447, n23448, n23449,
    n23450, n23451, n23452, n23453, n23454, n23455,
    n23456, n23457, n23458, n23459, n23460, n23461,
    n23462, n23463, n23464, n23465, n23466, n23467,
    n23468, n23469, n23470, n23471, n23472, n23473,
    n23474, n23475, n23476, n23477, n23478, n23479,
    n23480, n23481, n23482, n23483, n23484, n23485,
    n23486, n23487, n23488, n23489, n23490, n23491,
    n23492, n23493, n23494, n23495, n23496, n23497,
    n23498, n23499, n23500, n23501, n23502, n23503,
    n23504, n23505, n23506, n23507, n23508, n23509,
    n23510, n23511, n23512, n23513, n23514, n23515,
    n23516, n23517, n23518, n23519, n23520, n23521,
    n23522, n23523, n23524, n23525, n23526, n23527,
    n23528, n23529, n23530, n23531, n23532, n23533,
    n23534, n23535, n23536, n23537, n23538, n23540,
    n23541, n23542, n23543, n23544, n23545, n23546,
    n23547, n23548, n23549, n23550, n23551, n23552,
    n23553, n23554, n23555, n23556, n23557, n23558,
    n23559, n23560, n23561, n23562, n23563, n23564,
    n23565, n23566, n23567, n23568, n23569, n23570,
    n23571, n23572, n23573, n23574, n23575, n23576,
    n23577, n23578, n23579, n23580, n23581, n23582,
    n23583, n23584, n23585, n23586, n23587, n23588,
    n23589, n23590, n23591, n23592, n23593, n23594,
    n23595, n23596, n23597, n23598, n23599, n23600,
    n23601, n23602, n23603, n23604, n23605, n23606,
    n23607, n23608, n23609, n23610, n23611, n23612,
    n23613, n23614, n23615, n23616, n23617, n23618,
    n23619, n23620, n23621, n23622, n23623, n23624,
    n23625, n23626, n23627, n23628, n23629, n23630,
    n23631, n23632, n23633, n23634, n23635, n23636,
    n23637, n23638, n23639, n23640, n23641, n23642,
    n23643, n23644, n23645, n23646, n23647, n23648,
    n23649, n23650, n23651, n23652, n23653, n23654,
    n23655, n23656, n23657, n23658, n23659, n23660,
    n23661, n23662, n23663, n23664, n23665, n23666,
    n23667, n23668, n23669, n23670, n23671, n23672,
    n23673, n23674, n23675, n23676, n23677, n23678,
    n23679, n23680, n23681, n23682, n23683, n23684,
    n23685, n23686, n23687, n23688, n23689, n23690,
    n23691, n23692, n23693, n23694, n23695, n23696,
    n23697, n23698, n23699, n23700, n23701, n23702,
    n23703, n23704, n23705, n23706, n23707, n23708,
    n23709, n23710, n23711, n23712, n23713, n23714,
    n23715, n23716, n23717, n23718, n23719, n23720,
    n23721, n23722, n23723, n23724, n23725, n23726,
    n23727, n23728, n23729, n23730, n23731, n23732,
    n23733, n23734, n23735, n23736, n23737, n23738,
    n23739, n23740, n23741, n23742, n23743, n23744,
    n23745, n23746, n23747, n23748, n23749, n23750,
    n23751, n23752, n23753, n23754, n23755, n23756,
    n23757, n23758, n23759, n23760, n23761, n23762,
    n23763, n23764, n23765, n23766, n23767, n23768,
    n23769, n23770, n23771, n23772, n23773, n23774,
    n23775, n23776, n23777, n23778, n23779, n23780,
    n23781, n23782, n23783, n23784, n23785, n23786,
    n23787, n23788, n23789, n23790, n23791, n23792,
    n23793, n23794, n23795, n23796, n23797, n23798,
    n23799, n23800, n23801, n23802, n23803, n23804,
    n23805, n23806, n23807, n23808, n23809, n23810,
    n23811, n23812, n23813, n23814, n23815, n23816,
    n23817, n23818, n23819, n23820, n23821, n23822,
    n23823, n23824, n23825, n23826, n23827, n23828,
    n23829, n23830, n23831, n23832, n23833, n23834,
    n23835, n23836, n23837, n23838, n23839, n23840,
    n23841, n23842, n23843, n23844, n23845, n23846,
    n23847, n23848, n23849, n23850, n23851, n23852,
    n23853, n23854, n23855, n23856, n23857, n23858,
    n23859, n23860, n23861, n23862, n23863, n23864,
    n23865, n23866, n23867, n23868, n23869, n23870,
    n23871, n23872, n23873, n23874, n23875, n23876,
    n23877, n23878, n23879, n23880, n23881, n23882,
    n23883, n23884, n23885, n23886, n23887, n23888,
    n23889, n23890, n23891, n23892, n23893, n23894,
    n23895, n23896, n23897, n23898, n23899, n23900,
    n23901, n23902, n23903, n23904, n23905, n23906,
    n23907, n23908, n23909, n23910, n23911, n23912,
    n23913, n23914, n23915, n23916, n23917, n23918,
    n23919, n23920, n23921, n23922, n23923, n23924,
    n23925, n23926, n23927, n23928, n23929, n23930,
    n23931, n23932, n23933, n23934, n23935, n23936,
    n23937, n23938, n23939, n23940, n23941, n23942,
    n23943, n23944, n23945, n23946, n23947, n23948,
    n23949, n23950, n23951, n23952, n23953, n23954,
    n23955, n23956, n23957, n23958, n23959, n23960,
    n23961, n23962, n23963, n23964, n23965, n23966,
    n23967, n23968, n23969, n23970, n23971, n23972,
    n23973, n23974, n23975, n23976, n23977, n23978,
    n23979, n23980, n23981, n23982, n23983, n23984,
    n23985, n23986, n23987, n23988, n23989, n23990,
    n23991, n23992, n23993, n23994, n23995, n23996,
    n23997, n23998, n23999, n24000, n24001, n24002,
    n24003, n24004, n24005, n24006, n24007, n24008,
    n24009, n24010, n24011, n24012, n24013, n24014,
    n24016, n24017, n24018, n24019, n24020, n24021,
    n24022, n24023, n24024, n24025, n24026, n24027,
    n24028, n24029, n24030, n24031, n24032, n24033,
    n24034, n24035, n24036, n24037, n24038, n24039,
    n24040, n24041, n24042, n24043, n24044, n24045,
    n24046, n24047, n24048, n24049, n24050, n24051,
    n24052, n24053, n24054, n24055, n24056, n24057,
    n24058, n24059, n24060, n24061, n24062, n24063,
    n24064, n24065, n24066, n24067, n24068, n24069,
    n24070, n24071, n24072, n24073, n24074, n24075,
    n24076, n24077, n24078, n24079, n24080, n24081,
    n24082, n24083, n24084, n24085, n24086, n24087,
    n24088, n24089, n24090, n24091, n24092, n24093,
    n24094, n24095, n24096, n24097, n24098, n24099,
    n24100, n24101, n24102, n24103, n24104, n24105,
    n24106, n24107, n24108, n24109, n24110, n24111,
    n24112, n24113, n24114, n24115, n24116, n24117,
    n24118, n24119, n24120, n24121, n24122, n24123,
    n24124, n24125, n24126, n24127, n24128, n24129,
    n24130, n24131, n24132, n24133, n24134, n24135,
    n24136, n24137, n24138, n24139, n24140, n24141,
    n24142, n24143, n24144, n24145, n24146, n24147,
    n24148, n24149, n24150, n24151, n24152, n24153,
    n24154, n24155, n24156, n24157, n24158, n24159,
    n24160, n24161, n24162, n24163, n24164, n24165,
    n24166, n24167, n24168, n24169, n24170, n24171,
    n24172, n24173, n24174, n24175, n24176, n24177,
    n24178, n24179, n24180, n24181, n24182, n24183,
    n24184, n24185, n24186, n24187, n24188, n24189,
    n24190, n24191, n24192, n24193, n24194, n24195,
    n24196, n24197, n24198, n24199, n24200, n24201,
    n24202, n24203, n24204, n24205, n24206, n24207,
    n24208, n24209, n24210, n24211, n24212, n24213,
    n24214, n24215, n24216, n24217, n24218, n24219,
    n24220, n24221, n24222, n24223, n24224, n24225,
    n24226, n24227, n24228, n24229, n24230, n24231,
    n24232, n24233, n24234, n24235, n24236, n24237,
    n24238, n24239, n24240, n24241, n24242, n24243,
    n24244, n24245, n24246, n24247, n24248, n24249,
    n24250, n24251, n24252, n24253, n24254, n24255,
    n24256, n24257, n24258, n24259, n24260, n24261,
    n24262, n24263, n24264, n24265, n24266, n24267,
    n24268, n24269, n24270, n24271, n24272, n24273,
    n24274, n24275, n24276, n24277, n24278, n24279,
    n24280, n24281, n24282, n24283, n24284, n24285,
    n24286, n24287, n24288, n24289, n24290, n24291,
    n24292, n24293, n24294, n24295, n24296, n24297,
    n24298, n24299, n24300, n24301, n24302, n24303,
    n24304, n24305, n24306, n24307, n24308, n24309,
    n24310, n24311, n24312, n24313, n24314, n24315,
    n24316, n24317, n24318, n24319, n24320, n24321,
    n24322, n24323, n24324, n24325, n24326, n24327,
    n24328, n24329, n24330, n24331, n24332, n24333,
    n24334, n24335, n24336, n24337, n24338, n24339,
    n24340, n24341, n24342, n24343, n24344, n24345,
    n24346, n24347, n24348, n24349, n24350, n24351,
    n24352, n24353, n24354, n24355, n24356, n24357,
    n24358, n24359, n24360, n24361, n24362, n24363,
    n24364, n24365, n24366, n24367, n24368, n24369,
    n24370, n24371, n24372, n24373, n24374, n24375,
    n24376, n24377, n24378, n24379, n24380, n24381,
    n24382, n24383, n24384, n24385, n24386, n24387,
    n24388, n24389, n24390, n24391, n24392, n24393,
    n24394, n24395, n24396, n24397, n24398, n24399,
    n24400, n24401, n24402, n24403, n24404, n24405,
    n24406, n24407, n24408, n24409, n24410, n24411,
    n24412, n24413, n24414, n24415, n24416, n24417,
    n24418, n24419, n24420, n24421, n24422, n24423,
    n24424, n24425, n24426, n24427, n24428, n24429,
    n24430, n24431, n24432, n24433, n24434, n24435,
    n24436, n24437, n24438, n24439, n24440, n24441,
    n24442, n24443, n24444, n24445, n24446, n24447,
    n24448, n24449, n24450, n24451, n24452, n24453,
    n24454, n24455, n24456, n24457, n24458, n24459,
    n24460, n24461, n24462, n24464, n24465, n24466,
    n24467, n24468, n24469, n24470, n24471, n24472,
    n24473, n24474, n24475, n24476, n24477, n24478,
    n24479, n24480, n24481, n24482, n24483, n24484,
    n24485, n24486, n24487, n24488, n24489, n24490,
    n24491, n24492, n24493, n24494, n24495, n24496,
    n24497, n24498, n24499, n24500, n24501, n24502,
    n24503, n24504, n24505, n24506, n24507, n24508,
    n24509, n24510, n24511, n24512, n24513, n24514,
    n24515, n24516, n24517, n24518, n24519, n24520,
    n24521, n24522, n24523, n24524, n24525, n24526,
    n24527, n24528, n24529, n24530, n24531, n24532,
    n24533, n24534, n24535, n24536, n24537, n24538,
    n24539, n24540, n24541, n24542, n24543, n24544,
    n24545, n24546, n24547, n24548, n24549, n24550,
    n24551, n24552, n24553, n24554, n24555, n24556,
    n24557, n24558, n24559, n24560, n24561, n24562,
    n24563, n24564, n24565, n24566, n24567, n24568,
    n24569, n24570, n24571, n24572, n24573, n24574,
    n24575, n24576, n24577, n24578, n24579, n24580,
    n24581, n24582, n24583, n24584, n24585, n24586,
    n24587, n24588, n24589, n24590, n24591, n24592,
    n24593, n24594, n24595, n24596, n24597, n24598,
    n24599, n24600, n24601, n24602, n24603, n24604,
    n24605, n24606, n24607, n24608, n24609, n24610,
    n24611, n24612, n24613, n24614, n24615, n24616,
    n24617, n24618, n24619, n24620, n24621, n24622,
    n24623, n24624, n24625, n24626, n24627, n24628,
    n24629, n24630, n24631, n24632, n24633, n24634,
    n24635, n24636, n24637, n24638, n24639, n24640,
    n24641, n24642, n24643, n24644, n24645, n24646,
    n24647, n24648, n24649, n24650, n24651, n24652,
    n24653, n24654, n24655, n24656, n24657, n24658,
    n24659, n24660, n24661, n24662, n24663, n24664,
    n24665, n24666, n24667, n24668, n24669, n24670,
    n24671, n24672, n24673, n24674, n24675, n24676,
    n24677, n24678, n24679, n24680, n24681, n24682,
    n24683, n24684, n24685, n24686, n24687, n24688,
    n24689, n24690, n24691, n24692, n24693, n24694,
    n24695, n24696, n24697, n24698, n24699, n24700,
    n24701, n24702, n24703, n24704, n24705, n24706,
    n24707, n24708, n24709, n24710, n24711, n24712,
    n24713, n24714, n24715, n24716, n24717, n24718,
    n24719, n24720, n24721, n24722, n24723, n24724,
    n24725, n24726, n24727, n24728, n24729, n24730,
    n24731, n24732, n24733, n24734, n24735, n24736,
    n24737, n24738, n24739, n24740, n24741, n24742,
    n24743, n24744, n24745, n24746, n24747, n24748,
    n24749, n24750, n24751, n24752, n24753, n24754,
    n24755, n24756, n24757, n24758, n24759, n24760,
    n24761, n24762, n24763, n24764, n24765, n24766,
    n24767, n24768, n24769, n24770, n24771, n24772,
    n24773, n24774, n24775, n24776, n24777, n24778,
    n24779, n24780, n24781, n24782, n24783, n24784,
    n24785, n24786, n24787, n24788, n24789, n24790,
    n24791, n24792, n24793, n24794, n24795, n24796,
    n24797, n24798, n24799, n24800, n24801, n24802,
    n24803, n24804, n24805, n24806, n24807, n24808,
    n24809, n24810, n24811, n24812, n24813, n24814,
    n24815, n24816, n24817, n24818, n24819, n24820,
    n24821, n24822, n24823, n24824, n24825, n24826,
    n24827, n24828, n24829, n24830, n24831, n24832,
    n24833, n24834, n24835, n24836, n24837, n24838,
    n24839, n24840, n24841, n24842, n24843, n24844,
    n24845, n24846, n24847, n24848, n24849, n24850,
    n24851, n24852, n24853, n24854, n24855, n24856,
    n24857, n24858, n24859, n24860, n24861, n24862,
    n24863, n24864, n24865, n24866, n24867, n24868,
    n24869, n24870, n24871, n24872, n24873, n24874,
    n24875, n24876, n24877, n24878, n24879, n24880,
    n24881, n24882, n24883, n24884, n24885, n24886,
    n24887, n24888, n24889, n24890, n24891, n24892,
    n24893, n24894, n24895, n24896, n24897, n24898,
    n24899, n24900, n24901, n24902, n24903, n24904,
    n24905, n24906, n24907, n24908, n24909, n24910,
    n24911, n24912, n24913, n24914, n24915, n24916,
    n24917, n24918, n24919, n24920, n24921, n24922,
    n24923, n24924, n24925, n24926, n24927, n24928,
    n24929, n24930, n24931, n24932, n24933, n24934,
    n24935, n24936, n24937, n24938, n24939, n24940,
    n24941, n24942, n24943, n24944, n24946, n24947,
    n24948, n24949, n24950, n24951, n24952, n24953,
    n24954, n24955, n24956, n24957, n24958, n24959,
    n24960, n24961, n24962, n24963, n24964, n24965,
    n24966, n24967, n24968, n24969, n24970, n24971,
    n24972, n24973, n24974, n24975, n24976, n24977,
    n24978, n24979, n24980, n24981, n24982, n24983,
    n24984, n24985, n24986, n24987, n24988, n24989,
    n24990, n24991, n24992, n24993, n24994, n24995,
    n24996, n24997, n24998, n24999, n25000, n25001,
    n25002, n25003, n25004, n25005, n25006, n25007,
    n25008, n25009, n25010, n25011, n25012, n25013,
    n25014, n25015, n25016, n25017, n25018, n25019,
    n25020, n25021, n25022, n25023, n25024, n25025,
    n25026, n25027, n25028, n25029, n25030, n25031,
    n25032, n25033, n25034, n25035, n25036, n25037,
    n25038, n25039, n25040, n25041, n25042, n25043,
    n25044, n25045, n25046, n25047, n25048, n25049,
    n25050, n25051, n25052, n25053, n25054, n25055,
    n25056, n25057, n25058, n25059, n25060, n25061,
    n25062, n25063, n25064, n25065, n25066, n25067,
    n25068, n25069, n25070, n25071, n25072, n25073,
    n25074, n25075, n25076, n25077, n25078, n25079,
    n25080, n25081, n25082, n25083, n25084, n25085,
    n25086, n25087, n25088, n25089, n25090, n25091,
    n25092, n25093, n25094, n25095, n25096, n25097,
    n25098, n25099, n25100, n25101, n25102, n25103,
    n25104, n25105, n25106, n25107, n25108, n25109,
    n25110, n25111, n25112, n25113, n25114, n25115,
    n25116, n25117, n25118, n25119, n25120, n25121,
    n25122, n25123, n25124, n25125, n25126, n25127,
    n25128, n25129, n25130, n25131, n25132, n25133,
    n25134, n25135, n25136, n25137, n25138, n25139,
    n25140, n25141, n25142, n25143, n25144, n25145,
    n25146, n25147, n25148, n25149, n25150, n25151,
    n25152, n25153, n25154, n25155, n25156, n25157,
    n25158, n25159, n25160, n25161, n25162, n25163,
    n25164, n25165, n25166, n25167, n25168, n25169,
    n25170, n25171, n25172, n25173, n25174, n25175,
    n25176, n25177, n25178, n25179, n25180, n25181,
    n25182, n25183, n25184, n25185, n25186, n25187,
    n25188, n25189, n25190, n25191, n25192, n25193,
    n25194, n25195, n25196, n25197, n25198, n25199,
    n25200, n25201, n25202, n25203, n25204, n25205,
    n25206, n25207, n25208, n25209, n25210, n25211,
    n25212, n25213, n25214, n25215, n25216, n25217,
    n25218, n25219, n25220, n25221, n25222, n25223,
    n25224, n25225, n25226, n25227, n25228, n25229,
    n25230, n25231, n25232, n25233, n25234, n25235,
    n25236, n25237, n25238, n25239, n25240, n25241,
    n25242, n25243, n25244, n25245, n25246, n25247,
    n25248, n25249, n25250, n25251, n25252, n25253,
    n25254, n25255, n25256, n25257, n25258, n25259,
    n25260, n25261, n25262, n25263, n25264, n25265,
    n25266, n25267, n25268, n25269, n25270, n25271,
    n25272, n25273, n25274, n25275, n25276, n25277,
    n25278, n25279, n25280, n25281, n25282, n25283,
    n25284, n25285, n25286, n25287, n25288, n25289,
    n25290, n25291, n25292, n25293, n25294, n25295,
    n25296, n25297, n25298, n25299, n25300, n25301,
    n25302, n25303, n25304, n25305, n25306, n25307,
    n25308, n25309, n25310, n25311, n25312, n25313,
    n25314, n25315, n25316, n25317, n25318, n25319,
    n25320, n25321, n25322, n25323, n25324, n25325,
    n25326, n25327, n25328, n25329, n25330, n25331,
    n25332, n25333, n25334, n25335, n25336, n25337,
    n25338, n25339, n25340, n25341, n25342, n25343,
    n25344, n25345, n25346, n25347, n25348, n25349,
    n25350, n25351, n25352, n25353, n25354, n25355,
    n25356, n25357, n25358, n25359, n25360, n25361,
    n25362, n25363, n25364, n25365, n25366, n25367,
    n25368, n25369, n25370, n25371, n25372, n25373,
    n25374, n25375, n25376, n25377, n25378, n25379,
    n25380, n25381, n25382, n25383, n25384, n25385,
    n25386, n25387, n25388, n25389, n25390, n25391,
    n25392, n25393, n25394, n25395, n25396, n25397,
    n25398, n25399, n25400, n25401, n25402, n25403,
    n25404, n25405, n25406, n25407, n25408, n25409,
    n25410, n25411, n25412, n25413, n25415, n25416,
    n25417, n25418, n25419, n25420, n25421, n25422,
    n25423, n25424, n25425, n25426, n25427, n25428,
    n25429, n25430, n25431, n25432, n25433, n25434,
    n25435, n25436, n25437, n25438, n25439, n25440,
    n25441, n25442, n25443, n25444, n25445, n25446,
    n25447, n25448, n25449, n25450, n25451, n25452,
    n25453, n25454, n25455, n25456, n25457, n25458,
    n25459, n25460, n25461, n25462, n25463, n25464,
    n25465, n25466, n25467, n25468, n25469, n25470,
    n25471, n25472, n25473, n25474, n25475, n25476,
    n25477, n25478, n25479, n25480, n25481, n25482,
    n25483, n25484, n25485, n25486, n25487, n25488,
    n25489, n25490, n25491, n25492, n25493, n25494,
    n25495, n25496, n25497, n25498, n25499, n25500,
    n25501, n25502, n25503, n25504, n25505, n25506,
    n25507, n25508, n25509, n25510, n25511, n25512,
    n25513, n25514, n25515, n25516, n25517, n25518,
    n25519, n25520, n25521, n25522, n25523, n25524,
    n25525, n25526, n25527, n25528, n25529, n25530,
    n25531, n25532, n25533, n25534, n25535, n25536,
    n25537, n25538, n25539, n25540, n25541, n25542,
    n25543, n25544, n25545, n25546, n25547, n25548,
    n25549, n25550, n25551, n25552, n25553, n25554,
    n25555, n25556, n25557, n25558, n25559, n25560,
    n25561, n25562, n25563, n25564, n25565, n25566,
    n25567, n25568, n25569, n25570, n25571, n25572,
    n25573, n25574, n25575, n25576, n25577, n25578,
    n25579, n25580, n25581, n25582, n25583, n25584,
    n25585, n25586, n25587, n25588, n25589, n25590,
    n25591, n25592, n25593, n25594, n25595, n25596,
    n25597, n25598, n25599, n25600, n25601, n25602,
    n25603, n25604, n25605, n25606, n25607, n25608,
    n25609, n25610, n25611, n25612, n25613, n25614,
    n25615, n25616, n25617, n25618, n25619, n25620,
    n25621, n25622, n25623, n25624, n25625, n25626,
    n25627, n25628, n25629, n25630, n25631, n25632,
    n25633, n25634, n25635, n25636, n25637, n25638,
    n25639, n25640, n25641, n25642, n25643, n25644,
    n25645, n25646, n25647, n25648, n25649, n25650,
    n25651, n25652, n25653, n25654, n25655, n25656,
    n25657, n25658, n25659, n25660, n25661, n25662,
    n25663, n25664, n25665, n25666, n25667, n25668,
    n25669, n25670, n25671, n25672, n25673, n25674,
    n25675, n25676, n25677, n25678, n25679, n25680,
    n25681, n25682, n25683, n25684, n25685, n25686,
    n25687, n25688, n25689, n25690, n25691, n25692,
    n25693, n25694, n25695, n25696, n25697, n25698,
    n25699, n25700, n25701, n25702, n25703, n25704,
    n25705, n25706, n25707, n25708, n25709, n25710,
    n25711, n25712, n25713, n25714, n25715, n25716,
    n25717, n25718, n25719, n25720, n25721, n25722,
    n25723, n25724, n25725, n25726, n25727, n25728,
    n25729, n25730, n25731, n25732, n25733, n25734,
    n25735, n25736, n25737, n25738, n25739, n25740,
    n25741, n25742, n25743, n25744, n25745, n25746,
    n25747, n25748, n25749, n25750, n25751, n25752,
    n25753, n25754, n25755, n25756, n25757, n25758,
    n25759, n25760, n25761, n25762, n25763, n25764,
    n25765, n25766, n25767, n25768, n25769, n25770,
    n25771, n25772, n25773, n25774, n25775, n25776,
    n25777, n25778, n25779, n25780, n25781, n25782,
    n25783, n25784, n25785, n25786, n25787, n25788,
    n25789, n25790, n25791, n25792, n25793, n25794,
    n25795, n25796, n25797, n25798, n25799, n25800,
    n25801, n25802, n25803, n25804, n25805, n25806,
    n25807, n25808, n25809, n25810, n25811, n25812,
    n25813, n25814, n25815, n25816, n25817, n25818,
    n25819, n25820, n25821, n25822, n25823, n25824,
    n25825, n25826, n25827, n25828, n25829, n25830,
    n25831, n25832, n25833, n25834, n25835, n25836,
    n25837, n25838, n25839, n25840, n25841, n25842,
    n25843, n25844, n25845, n25846, n25847, n25848,
    n25849, n25850, n25851, n25852, n25853, n25854,
    n25855, n25856, n25857, n25858, n25859, n25860,
    n25861, n25862, n25863, n25864, n25865, n25866,
    n25867, n25868, n25869, n25870, n25871, n25872,
    n25873, n25874, n25875, n25876, n25877, n25878,
    n25879, n25880, n25881, n25882, n25883, n25884,
    n25885, n25886, n25887, n25888, n25889, n25890,
    n25891, n25892, n25894, n25895, n25896, n25897,
    n25898, n25899, n25900, n25901, n25902, n25903,
    n25904, n25905, n25906, n25907, n25908, n25909,
    n25910, n25911, n25912, n25913, n25914, n25915,
    n25916, n25917, n25918, n25919, n25920, n25921,
    n25922, n25923, n25924, n25925, n25926, n25927,
    n25928, n25929, n25930, n25931, n25932, n25933,
    n25934, n25935, n25936, n25937, n25938, n25939,
    n25940, n25941, n25942, n25943, n25944, n25945,
    n25946, n25947, n25948, n25949, n25950, n25951,
    n25952, n25953, n25954, n25955, n25956, n25957,
    n25958, n25959, n25960, n25961, n25962, n25963,
    n25964, n25965, n25966, n25967, n25968, n25969,
    n25970, n25971, n25972, n25973, n25974, n25975,
    n25976, n25977, n25978, n25979, n25980, n25981,
    n25982, n25983, n25984, n25985, n25986, n25987,
    n25988, n25989, n25990, n25991, n25992, n25993,
    n25994, n25995, n25996, n25997, n25998, n25999,
    n26000, n26001, n26002, n26003, n26004, n26005,
    n26006, n26007, n26008, n26009, n26010, n26011,
    n26012, n26013, n26014, n26015, n26016, n26017,
    n26018, n26019, n26020, n26021, n26022, n26023,
    n26024, n26025, n26026, n26027, n26028, n26029,
    n26030, n26031, n26032, n26033, n26034, n26035,
    n26036, n26037, n26038, n26039, n26040, n26041,
    n26042, n26043, n26044, n26045, n26046, n26047,
    n26048, n26049, n26050, n26051, n26052, n26053,
    n26054, n26055, n26056, n26057, n26058, n26059,
    n26060, n26061, n26062, n26063, n26064, n26065,
    n26066, n26067, n26068, n26069, n26070, n26071,
    n26072, n26073, n26074, n26075, n26076, n26077,
    n26078, n26079, n26080, n26081, n26082, n26083,
    n26084, n26085, n26086, n26087, n26088, n26089,
    n26090, n26091, n26092, n26093, n26094, n26095,
    n26096, n26097, n26098, n26099, n26100, n26101,
    n26102, n26103, n26104, n26105, n26106, n26107,
    n26108, n26109, n26110, n26111, n26112, n26113,
    n26114, n26115, n26116, n26117, n26118, n26119,
    n26120, n26121, n26122, n26123, n26124, n26125,
    n26126, n26127, n26128, n26129, n26130, n26131,
    n26132, n26133, n26134, n26135, n26136, n26137,
    n26138, n26139, n26140, n26141, n26142, n26143,
    n26144, n26145, n26146, n26147, n26148, n26149,
    n26150, n26151, n26152, n26153, n26154, n26155,
    n26156, n26157, n26158, n26159, n26160, n26161,
    n26162, n26163, n26164, n26165, n26166, n26167,
    n26168, n26169, n26170, n26171, n26172, n26173,
    n26174, n26175, n26176, n26177, n26178, n26179,
    n26180, n26181, n26182, n26183, n26184, n26185,
    n26186, n26187, n26188, n26189, n26190, n26191,
    n26192, n26193, n26194, n26195, n26196, n26197,
    n26198, n26199, n26200, n26201, n26202, n26203,
    n26204, n26205, n26206, n26207, n26208, n26209,
    n26210, n26211, n26212, n26213, n26214, n26215,
    n26216, n26217, n26218, n26219, n26220, n26221,
    n26222, n26223, n26224, n26225, n26226, n26227,
    n26228, n26229, n26230, n26231, n26232, n26233,
    n26234, n26235, n26236, n26237, n26238, n26239,
    n26240, n26241, n26242, n26243, n26244, n26245,
    n26246, n26247, n26248, n26249, n26250, n26251,
    n26252, n26253, n26254, n26255, n26256, n26257,
    n26258, n26259, n26260, n26261, n26262, n26263,
    n26264, n26265, n26266, n26267, n26268, n26269,
    n26270, n26271, n26272, n26273, n26274, n26275,
    n26276, n26277, n26278, n26279, n26280, n26281,
    n26282, n26283, n26284, n26285, n26286, n26287,
    n26288, n26289, n26290, n26291, n26292, n26293,
    n26294, n26295, n26296, n26297, n26298, n26299,
    n26300, n26301, n26302, n26303, n26304, n26305,
    n26306, n26307, n26308, n26309, n26310, n26311,
    n26312, n26313, n26314, n26315, n26316, n26317,
    n26318, n26319, n26320, n26321, n26322, n26323,
    n26324, n26325, n26326, n26327, n26328, n26329,
    n26330, n26331, n26332, n26333, n26334, n26335,
    n26336, n26337, n26338, n26339, n26340, n26341,
    n26342, n26343, n26344, n26345, n26346, n26347,
    n26348, n26349, n26350, n26351, n26352, n26353,
    n26354, n26355, n26356, n26357, n26358, n26359,
    n26360, n26361, n26362, n26363, n26364, n26365,
    n26366, n26367, n26369, n26370, n26371, n26372,
    n26373, n26374, n26375, n26376, n26377, n26378,
    n26379, n26380, n26381, n26382, n26383, n26384,
    n26385, n26386, n26387, n26388, n26389, n26390,
    n26391, n26392, n26393, n26394, n26395, n26396,
    n26397, n26398, n26399, n26400, n26401, n26402,
    n26403, n26404, n26405, n26406, n26407, n26408,
    n26409, n26410, n26411, n26412, n26413, n26414,
    n26415, n26416, n26417, n26418, n26419, n26420,
    n26421, n26422, n26423, n26424, n26425, n26426,
    n26427, n26428, n26429, n26430, n26431, n26432,
    n26433, n26434, n26435, n26436, n26437, n26438,
    n26439, n26440, n26441, n26442, n26443, n26444,
    n26445, n26446, n26447, n26448, n26449, n26450,
    n26451, n26452, n26453, n26454, n26455, n26456,
    n26457, n26458, n26459, n26460, n26461, n26462,
    n26463, n26464, n26465, n26466, n26467, n26468,
    n26469, n26470, n26471, n26472, n26473, n26474,
    n26475, n26476, n26477, n26478, n26479, n26480,
    n26481, n26482, n26483, n26484, n26485, n26486,
    n26487, n26488, n26489, n26490, n26491, n26492,
    n26493, n26494, n26495, n26496, n26497, n26498,
    n26499, n26500, n26501, n26502, n26503, n26504,
    n26505, n26506, n26507, n26508, n26509, n26510,
    n26511, n26512, n26513, n26514, n26515, n26516,
    n26517, n26518, n26519, n26520, n26521, n26522,
    n26523, n26524, n26525, n26526, n26527, n26528,
    n26529, n26530, n26531, n26532, n26533, n26534,
    n26535, n26536, n26537, n26538, n26539, n26540,
    n26541, n26542, n26543, n26544, n26545, n26546,
    n26547, n26548, n26549, n26550, n26551, n26552,
    n26553, n26554, n26555, n26556, n26557, n26558,
    n26559, n26560, n26561, n26562, n26563, n26564,
    n26565, n26566, n26567, n26568, n26569, n26570,
    n26571, n26572, n26573, n26574, n26575, n26576,
    n26577, n26578, n26579, n26580, n26581, n26582,
    n26583, n26584, n26585, n26586, n26587, n26588,
    n26589, n26590, n26591, n26592, n26593, n26594,
    n26595, n26596, n26597, n26598, n26599, n26600,
    n26601, n26602, n26603, n26604, n26605, n26606,
    n26607, n26608, n26609, n26610, n26611, n26612,
    n26613, n26614, n26615, n26616, n26617, n26618,
    n26619, n26620, n26621, n26622, n26623, n26624,
    n26625, n26626, n26627, n26628, n26629, n26630,
    n26631, n26632, n26633, n26634, n26635, n26636,
    n26637, n26638, n26639, n26640, n26641, n26642,
    n26643, n26644, n26645, n26646, n26647, n26648,
    n26649, n26650, n26651, n26652, n26653, n26654,
    n26655, n26656, n26657, n26658, n26659, n26660,
    n26661, n26662, n26663, n26664, n26665, n26666,
    n26667, n26668, n26669, n26670, n26671, n26672,
    n26673, n26674, n26675, n26676, n26677, n26678,
    n26679, n26680, n26681, n26682, n26683, n26684,
    n26685, n26686, n26687, n26688, n26689, n26690,
    n26691, n26692, n26693, n26694, n26695, n26696,
    n26697, n26698, n26699, n26700, n26701, n26702,
    n26703, n26704, n26705, n26706, n26707, n26708,
    n26709, n26710, n26711, n26712, n26713, n26714,
    n26715, n26716, n26717, n26718, n26719, n26720,
    n26721, n26722, n26723, n26724, n26725, n26726,
    n26727, n26728, n26729, n26730, n26731, n26732,
    n26733, n26734, n26735, n26736, n26737, n26738,
    n26739, n26740, n26741, n26742, n26743, n26744,
    n26745, n26746, n26747, n26748, n26749, n26750,
    n26751, n26752, n26753, n26754, n26755, n26756,
    n26757, n26758, n26759, n26760, n26761, n26762,
    n26763, n26764, n26765, n26766, n26767, n26768,
    n26769, n26770, n26771, n26772, n26773, n26774,
    n26775, n26776, n26777, n26778, n26779, n26780,
    n26781, n26782, n26783, n26784, n26785, n26786,
    n26787, n26788, n26789, n26790, n26791, n26792,
    n26793, n26794, n26795, n26796, n26797, n26798,
    n26799, n26800, n26801, n26802, n26803, n26804,
    n26805, n26806, n26807, n26808, n26809, n26810,
    n26811, n26812, n26813, n26814, n26815, n26816,
    n26817, n26818, n26819, n26820, n26821, n26822,
    n26823, n26824, n26825, n26826, n26827, n26828,
    n26829, n26830, n26831, n26832, n26833, n26834,
    n26835, n26836, n26837, n26838, n26839, n26840,
    n26841, n26842, n26844, n26845, n26846, n26847,
    n26848, n26849, n26850, n26851, n26852, n26853,
    n26854, n26855, n26856, n26857, n26858, n26859,
    n26860, n26861, n26862, n26863, n26864, n26865,
    n26866, n26867, n26868, n26869, n26870, n26871,
    n26872, n26873, n26874, n26875, n26876, n26877,
    n26878, n26879, n26880, n26881, n26882, n26883,
    n26884, n26885, n26886, n26887, n26888, n26889,
    n26890, n26891, n26892, n26893, n26894, n26895,
    n26896, n26897, n26898, n26899, n26900, n26901,
    n26902, n26903, n26904, n26905, n26906, n26907,
    n26908, n26909, n26910, n26911, n26912, n26913,
    n26914, n26915, n26916, n26917, n26918, n26919,
    n26920, n26921, n26922, n26923, n26924, n26925,
    n26926, n26927, n26928, n26929, n26930, n26931,
    n26932, n26933, n26934, n26935, n26936, n26937,
    n26938, n26939, n26940, n26941, n26942, n26943,
    n26944, n26945, n26946, n26947, n26948, n26949,
    n26950, n26951, n26952, n26953, n26954, n26955,
    n26956, n26957, n26958, n26959, n26960, n26961,
    n26962, n26963, n26964, n26965, n26966, n26967,
    n26968, n26969, n26970, n26971, n26972, n26973,
    n26974, n26975, n26976, n26977, n26978, n26979,
    n26980, n26981, n26982, n26983, n26984, n26985,
    n26986, n26987, n26988, n26989, n26990, n26991,
    n26992, n26993, n26994, n26995, n26996, n26997,
    n26998, n26999, n27000, n27001, n27002, n27003,
    n27004, n27005, n27006, n27007, n27008, n27009,
    n27010, n27011, n27012, n27013, n27014, n27015,
    n27016, n27017, n27018, n27019, n27020, n27021,
    n27022, n27023, n27024, n27025, n27026, n27027,
    n27028, n27029, n27030, n27031, n27032, n27033,
    n27034, n27035, n27036, n27037, n27038, n27039,
    n27040, n27041, n27042, n27043, n27044, n27045,
    n27046, n27047, n27048, n27049, n27050, n27051,
    n27052, n27053, n27054, n27055, n27056, n27057,
    n27058, n27059, n27060, n27061, n27062, n27063,
    n27064, n27065, n27066, n27067, n27068, n27069,
    n27070, n27071, n27072, n27073, n27074, n27075,
    n27076, n27077, n27078, n27079, n27080, n27081,
    n27082, n27083, n27084, n27085, n27086, n27087,
    n27088, n27089, n27090, n27091, n27092, n27093,
    n27094, n27095, n27096, n27097, n27098, n27099,
    n27100, n27101, n27102, n27103, n27104, n27105,
    n27106, n27107, n27108, n27109, n27110, n27111,
    n27112, n27113, n27114, n27115, n27116, n27117,
    n27118, n27119, n27120, n27121, n27122, n27123,
    n27124, n27125, n27126, n27127, n27128, n27129,
    n27130, n27131, n27132, n27133, n27134, n27135,
    n27136, n27137, n27138, n27139, n27140, n27141,
    n27142, n27143, n27144, n27145, n27146, n27147,
    n27148, n27149, n27150, n27151, n27152, n27153,
    n27154, n27155, n27156, n27157, n27158, n27159,
    n27160, n27161, n27162, n27163, n27164, n27165,
    n27166, n27167, n27168, n27169, n27170, n27171,
    n27172, n27173, n27174, n27175, n27176, n27177,
    n27178, n27179, n27180, n27181, n27182, n27183,
    n27184, n27185, n27186, n27187, n27188, n27189,
    n27190, n27191, n27192, n27193, n27194, n27195,
    n27196, n27197, n27198, n27199, n27200, n27201,
    n27202, n27203, n27204, n27205, n27206, n27207,
    n27208, n27209, n27210, n27211, n27212, n27213,
    n27214, n27215, n27216, n27217, n27218, n27219,
    n27220, n27221, n27222, n27223, n27224, n27225,
    n27226, n27227, n27228, n27229, n27230, n27231,
    n27232, n27233, n27234, n27235, n27236, n27237,
    n27238, n27239, n27240, n27241, n27242, n27243,
    n27244, n27245, n27246, n27247, n27248, n27249,
    n27250, n27251, n27252, n27253, n27254, n27255,
    n27256, n27257, n27258, n27259, n27260, n27261,
    n27262, n27263, n27264, n27265, n27266, n27267,
    n27268, n27269, n27270, n27271, n27272, n27273,
    n27274, n27275, n27276, n27277, n27278, n27279,
    n27280, n27281, n27282, n27283, n27284, n27285,
    n27286, n27287, n27288, n27289, n27290, n27291,
    n27292, n27293, n27294, n27295, n27296, n27297,
    n27298, n27299, n27300, n27301, n27302, n27303,
    n27304, n27305, n27306, n27307, n27308, n27309,
    n27310, n27311, n27313, n27314, n27315, n27316,
    n27317, n27318, n27319, n27320, n27321, n27322,
    n27323, n27324, n27325, n27326, n27327, n27328,
    n27329, n27330, n27331, n27332, n27333, n27334,
    n27335, n27336, n27337, n27338, n27339, n27340,
    n27341, n27342, n27343, n27344, n27345, n27346,
    n27347, n27348, n27349, n27350, n27351, n27352,
    n27353, n27354, n27355, n27356, n27357, n27358,
    n27359, n27360, n27361, n27362, n27363, n27364,
    n27365, n27366, n27367, n27368, n27369, n27370,
    n27371, n27372, n27373, n27374, n27375, n27376,
    n27377, n27378, n27379, n27380, n27381, n27382,
    n27383, n27384, n27385, n27386, n27387, n27388,
    n27389, n27390, n27391, n27392, n27393, n27394,
    n27395, n27396, n27397, n27398, n27399, n27400,
    n27401, n27402, n27403, n27404, n27405, n27406,
    n27407, n27408, n27409, n27410, n27411, n27412,
    n27413, n27414, n27415, n27416, n27417, n27418,
    n27419, n27420, n27421, n27422, n27423, n27424,
    n27425, n27426, n27427, n27428, n27429, n27430,
    n27431, n27432, n27433, n27434, n27435, n27436,
    n27437, n27438, n27439, n27440, n27441, n27442,
    n27443, n27444, n27445, n27446, n27447, n27448,
    n27449, n27450, n27451, n27452, n27453, n27454,
    n27455, n27456, n27457, n27458, n27459, n27460,
    n27461, n27462, n27463, n27464, n27465, n27466,
    n27467, n27468, n27469, n27470, n27471, n27472,
    n27473, n27474, n27475, n27476, n27477, n27478,
    n27479, n27480, n27481, n27482, n27483, n27484,
    n27485, n27486, n27487, n27488, n27489, n27490,
    n27491, n27492, n27493, n27494, n27495, n27496,
    n27497, n27498, n27499, n27500, n27501, n27502,
    n27503, n27504, n27505, n27506, n27507, n27508,
    n27509, n27510, n27511, n27512, n27513, n27514,
    n27515, n27516, n27517, n27518, n27519, n27520,
    n27521, n27522, n27523, n27524, n27525, n27526,
    n27527, n27528, n27529, n27530, n27531, n27532,
    n27533, n27534, n27535, n27536, n27537, n27538,
    n27539, n27540, n27541, n27542, n27543, n27544,
    n27545, n27546, n27547, n27548, n27549, n27550,
    n27551, n27552, n27553, n27554, n27555, n27556,
    n27557, n27558, n27559, n27560, n27561, n27562,
    n27563, n27564, n27565, n27566, n27567, n27568,
    n27569, n27570, n27571, n27572, n27573, n27574,
    n27575, n27576, n27577, n27578, n27579, n27580,
    n27581, n27582, n27583, n27584, n27585, n27586,
    n27587, n27588, n27589, n27590, n27591, n27592,
    n27593, n27594, n27595, n27596, n27597, n27598,
    n27599, n27600, n27601, n27602, n27603, n27604,
    n27605, n27606, n27607, n27608, n27609, n27610,
    n27611, n27612, n27613, n27614, n27615, n27616,
    n27617, n27618, n27619, n27620, n27621, n27622,
    n27623, n27624, n27625, n27626, n27627, n27628,
    n27629, n27630, n27631, n27632, n27633, n27634,
    n27635, n27636, n27637, n27638, n27639, n27640,
    n27641, n27642, n27643, n27644, n27645, n27646,
    n27647, n27648, n27649, n27650, n27651, n27652,
    n27653, n27654, n27655, n27656, n27657, n27658,
    n27659, n27660, n27661, n27662, n27663, n27664,
    n27665, n27666, n27667, n27668, n27669, n27670,
    n27671, n27672, n27673, n27674, n27675, n27676,
    n27677, n27678, n27679, n27680, n27681, n27682,
    n27683, n27684, n27685, n27686, n27687, n27688,
    n27689, n27690, n27691, n27692, n27693, n27694,
    n27695, n27696, n27697, n27698, n27699, n27700,
    n27701, n27702, n27703, n27704, n27705, n27706,
    n27707, n27708, n27709, n27710, n27711, n27712,
    n27713, n27714, n27715, n27716, n27717, n27718,
    n27719, n27720, n27721, n27722, n27723, n27724,
    n27725, n27726, n27727, n27728, n27729, n27730,
    n27731, n27732, n27733, n27734, n27735, n27736,
    n27737, n27738, n27739, n27740, n27741, n27742,
    n27743, n27744, n27745, n27746, n27747, n27748,
    n27749, n27750, n27751, n27752, n27753, n27754,
    n27755, n27756, n27757, n27758, n27759, n27760,
    n27761, n27762, n27763, n27764, n27765, n27766,
    n27767, n27768, n27769, n27770, n27771, n27772,
    n27773, n27774, n27775, n27776, n27777, n27778,
    n27779, n27780, n27782, n27783, n27784, n27785,
    n27786, n27787, n27788, n27789, n27790, n27791,
    n27792, n27793, n27794, n27795, n27796, n27797,
    n27798, n27799, n27800, n27801, n27802, n27803,
    n27804, n27805, n27806, n27807, n27808, n27809,
    n27810, n27811, n27812, n27813, n27814, n27815,
    n27816, n27817, n27818, n27819, n27820, n27821,
    n27822, n27823, n27824, n27825, n27826, n27827,
    n27828, n27829, n27830, n27831, n27832, n27833,
    n27834, n27835, n27836, n27837, n27838, n27839,
    n27840, n27841, n27842, n27843, n27844, n27845,
    n27846, n27847, n27848, n27849, n27850, n27851,
    n27852, n27853, n27854, n27855, n27856, n27857,
    n27858, n27859, n27860, n27861, n27862, n27863,
    n27864, n27865, n27866, n27867, n27868, n27869,
    n27870, n27871, n27872, n27873, n27874, n27875,
    n27876, n27877, n27878, n27879, n27880, n27881,
    n27882, n27883, n27884, n27885, n27886, n27887,
    n27888, n27889, n27890, n27891, n27892, n27893,
    n27894, n27895, n27896, n27897, n27898, n27899,
    n27900, n27901, n27902, n27903, n27904, n27905,
    n27906, n27907, n27908, n27909, n27910, n27911,
    n27912, n27913, n27914, n27915, n27916, n27917,
    n27918, n27919, n27920, n27921, n27922, n27923,
    n27924, n27925, n27926, n27927, n27928, n27929,
    n27930, n27931, n27932, n27933, n27934, n27935,
    n27936, n27937, n27938, n27939, n27940, n27941,
    n27942, n27943, n27944, n27945, n27946, n27947,
    n27948, n27949, n27950, n27951, n27952, n27953,
    n27954, n27955, n27956, n27957, n27958, n27959,
    n27960, n27961, n27962, n27963, n27964, n27965,
    n27966, n27967, n27968, n27969, n27970, n27971,
    n27972, n27973, n27974, n27975, n27976, n27977,
    n27978, n27979, n27980, n27981, n27982, n27983,
    n27984, n27985, n27986, n27987, n27988, n27989,
    n27990, n27991, n27992, n27993, n27994, n27995,
    n27996, n27997, n27998, n27999, n28000, n28001,
    n28002, n28003, n28004, n28005, n28006, n28007,
    n28008, n28009, n28010, n28011, n28012, n28013,
    n28014, n28015, n28016, n28017, n28018, n28019,
    n28020, n28021, n28022, n28023, n28024, n28025,
    n28026, n28027, n28028, n28029, n28030, n28031,
    n28032, n28033, n28034, n28035, n28036, n28037,
    n28038, n28039, n28040, n28041, n28042, n28043,
    n28044, n28045, n28046, n28047, n28048, n28049,
    n28050, n28051, n28052, n28053, n28054, n28055,
    n28056, n28057, n28058, n28059, n28060, n28061,
    n28062, n28063, n28064, n28065, n28066, n28067,
    n28068, n28069, n28070, n28071, n28072, n28073,
    n28074, n28075, n28076, n28077, n28078, n28079,
    n28080, n28081, n28082, n28083, n28084, n28085,
    n28086, n28087, n28088, n28089, n28090, n28091,
    n28092, n28093, n28094, n28095, n28096, n28097,
    n28098, n28099, n28100, n28101, n28102, n28103,
    n28104, n28105, n28106, n28107, n28108, n28109,
    n28110, n28111, n28112, n28113, n28114, n28115,
    n28116, n28117, n28118, n28119, n28120, n28121,
    n28122, n28123, n28124, n28125, n28126, n28127,
    n28128, n28129, n28130, n28131, n28132, n28133,
    n28134, n28135, n28136, n28137, n28138, n28139,
    n28140, n28141, n28142, n28143, n28144, n28145,
    n28146, n28147, n28148, n28149, n28150, n28151,
    n28152, n28153, n28154, n28155, n28156, n28157,
    n28158, n28159, n28160, n28161, n28162, n28163,
    n28164, n28165, n28166, n28167, n28168, n28169,
    n28170, n28171, n28172, n28173, n28174, n28175,
    n28176, n28177, n28178, n28179, n28180, n28181,
    n28182, n28183, n28184, n28185, n28186, n28187,
    n28188, n28189, n28190, n28191, n28192, n28193,
    n28194, n28195, n28196, n28197, n28198, n28199,
    n28200, n28201, n28202, n28203, n28204, n28205,
    n28206, n28207, n28208, n28209, n28210, n28211,
    n28212, n28213, n28214, n28215, n28216, n28217,
    n28218, n28219, n28220, n28221, n28222, n28223,
    n28224, n28225, n28226, n28227, n28228, n28229,
    n28230, n28231, n28232, n28233, n28234, n28235,
    n28236, n28237, n28238, n28239, n28240, n28241,
    n28242, n28243, n28244, n28245, n28246, n28247,
    n28248, n28249, n28251, n28252, n28253, n28254,
    n28255, n28256, n28257, n28258, n28259, n28260,
    n28261, n28262, n28263, n28264, n28265, n28266,
    n28267, n28268, n28269, n28270, n28271, n28272,
    n28273, n28274, n28275, n28276, n28277, n28278,
    n28279, n28280, n28281, n28282, n28283, n28284,
    n28285, n28286, n28287, n28288, n28289, n28290,
    n28291, n28292, n28293, n28294, n28295, n28296,
    n28297, n28298, n28299, n28300, n28301, n28302,
    n28303, n28304, n28305, n28306, n28307, n28308,
    n28309, n28310, n28311, n28312, n28313, n28314,
    n28315, n28316, n28317, n28318, n28319, n28320,
    n28321, n28322, n28323, n28324, n28325, n28326,
    n28327, n28328, n28329, n28330, n28331, n28332,
    n28333, n28334, n28335, n28336, n28337, n28338,
    n28339, n28340, n28341, n28342, n28343, n28344,
    n28345, n28346, n28347, n28348, n28349, n28350,
    n28351, n28352, n28353, n28354, n28355, n28356,
    n28357, n28358, n28359, n28360, n28361, n28362,
    n28363, n28364, n28365, n28366, n28367, n28368,
    n28369, n28370, n28371, n28372, n28373, n28374,
    n28375, n28376, n28377, n28378, n28379, n28380,
    n28381, n28382, n28383, n28384, n28385, n28386,
    n28387, n28388, n28389, n28390, n28391, n28392,
    n28393, n28394, n28395, n28396, n28397, n28398,
    n28399, n28400, n28401, n28402, n28403, n28404,
    n28405, n28406, n28407, n28408, n28409, n28410,
    n28411, n28412, n28413, n28414, n28415, n28416,
    n28417, n28418, n28419, n28420, n28421, n28422,
    n28423, n28424, n28425, n28426, n28427, n28428,
    n28429, n28430, n28431, n28432, n28433, n28434,
    n28435, n28436, n28437, n28438, n28439, n28440,
    n28441, n28442, n28443, n28444, n28445, n28446,
    n28447, n28448, n28449, n28450, n28451, n28452,
    n28453, n28454, n28455, n28456, n28457, n28458,
    n28459, n28460, n28461, n28462, n28463, n28464,
    n28465, n28466, n28467, n28468, n28469, n28470,
    n28471, n28472, n28473, n28474, n28475, n28476,
    n28477, n28478, n28479, n28480, n28481, n28482,
    n28483, n28484, n28485, n28486, n28487, n28488,
    n28489, n28490, n28491, n28492, n28493, n28494,
    n28495, n28496, n28497, n28498, n28499, n28500,
    n28501, n28502, n28503, n28504, n28505, n28506,
    n28507, n28508, n28509, n28510, n28511, n28512,
    n28513, n28514, n28515, n28516, n28517, n28518,
    n28519, n28520, n28521, n28522, n28523, n28524,
    n28525, n28526, n28527, n28528, n28529, n28530,
    n28531, n28532, n28533, n28534, n28535, n28536,
    n28537, n28538, n28539, n28540, n28541, n28542,
    n28543, n28544, n28545, n28546, n28547, n28548,
    n28549, n28550, n28551, n28552, n28553, n28554,
    n28555, n28556, n28557, n28558, n28559, n28560,
    n28561, n28562, n28563, n28564, n28565, n28566,
    n28567, n28568, n28569, n28570, n28571, n28572,
    n28573, n28574, n28575, n28576, n28577, n28578,
    n28579, n28580, n28581, n28582, n28583, n28584,
    n28585, n28586, n28587, n28588, n28589, n28590,
    n28591, n28592, n28593, n28594, n28595, n28596,
    n28597, n28598, n28599, n28600, n28601, n28602,
    n28603, n28604, n28605, n28606, n28607, n28608,
    n28609, n28610, n28611, n28612, n28613, n28614,
    n28615, n28616, n28617, n28618, n28619, n28620,
    n28621, n28622, n28623, n28624, n28625, n28626,
    n28627, n28628, n28629, n28630, n28631, n28632,
    n28633, n28634, n28635, n28636, n28637, n28638,
    n28639, n28640, n28641, n28642, n28643, n28644,
    n28645, n28646, n28647, n28648, n28649, n28650,
    n28651, n28652, n28653, n28654, n28655, n28656,
    n28657, n28658, n28659, n28660, n28661, n28662,
    n28663, n28664, n28665, n28666, n28667, n28668,
    n28669, n28670, n28671, n28672, n28673, n28674,
    n28675, n28676, n28677, n28678, n28679, n28680,
    n28681, n28682, n28683, n28684, n28685, n28686,
    n28687, n28688, n28689, n28690, n28691, n28692,
    n28693, n28694, n28695, n28696, n28697, n28698,
    n28699, n28700, n28701, n28702, n28703, n28704,
    n28705, n28706, n28707, n28708, n28709, n28710,
    n28711, n28712, n28713, n28714, n28715, n28716,
    n28717, n28718, n28719, n28720, n28721, n28722,
    n28723, n28724, n28726, n28727, n28728, n28729,
    n28730, n28731, n28732, n28733, n28734, n28735,
    n28736, n28737, n28738, n28739, n28740, n28741,
    n28742, n28743, n28744, n28745, n28746, n28747,
    n28748, n28749, n28750, n28751, n28752, n28753,
    n28754, n28755, n28756, n28757, n28758, n28759,
    n28760, n28761, n28762, n28763, n28764, n28765,
    n28766, n28767, n28768, n28769, n28770, n28771,
    n28772, n28773, n28774, n28775, n28776, n28777,
    n28778, n28779, n28780, n28781, n28782, n28783,
    n28784, n28785, n28786, n28787, n28788, n28789,
    n28790, n28791, n28792, n28793, n28794, n28795,
    n28796, n28797, n28798, n28799, n28800, n28801,
    n28802, n28803, n28804, n28805, n28806, n28807,
    n28808, n28809, n28810, n28811, n28812, n28813,
    n28814, n28815, n28816, n28817, n28818, n28819,
    n28820, n28821, n28822, n28823, n28824, n28825,
    n28826, n28827, n28828, n28829, n28830, n28831,
    n28832, n28833, n28834, n28835, n28836, n28837,
    n28838, n28839, n28840, n28841, n28842, n28843,
    n28844, n28845, n28846, n28847, n28848, n28849,
    n28850, n28851, n28852, n28853, n28854, n28855,
    n28856, n28857, n28858, n28859, n28860, n28861,
    n28862, n28863, n28864, n28865, n28866, n28867,
    n28868, n28869, n28870, n28871, n28872, n28873,
    n28874, n28875, n28876, n28877, n28878, n28879,
    n28880, n28881, n28882, n28883, n28884, n28885,
    n28886, n28887, n28888, n28889, n28890, n28891,
    n28892, n28893, n28894, n28895, n28896, n28897,
    n28898, n28899, n28900, n28901, n28902, n28903,
    n28904, n28905, n28906, n28907, n28908, n28909,
    n28910, n28911, n28912, n28913, n28914, n28915,
    n28916, n28917, n28918, n28919, n28920, n28921,
    n28922, n28923, n28924, n28925, n28926, n28927,
    n28928, n28929, n28930, n28931, n28932, n28933,
    n28934, n28935, n28936, n28937, n28938, n28939,
    n28940, n28941, n28942, n28943, n28944, n28945,
    n28946, n28947, n28948, n28949, n28950, n28951,
    n28952, n28953, n28954, n28955, n28956, n28957,
    n28958, n28959, n28960, n28961, n28962, n28963,
    n28964, n28965, n28966, n28967, n28968, n28969,
    n28970, n28971, n28972, n28973, n28974, n28975,
    n28976, n28977, n28978, n28979, n28980, n28981,
    n28982, n28983, n28984, n28985, n28986, n28987,
    n28988, n28989, n28990, n28991, n28992, n28993,
    n28994, n28995, n28996, n28997, n28998, n28999,
    n29000, n29001, n29002, n29003, n29004, n29005,
    n29006, n29007, n29008, n29009, n29010, n29011,
    n29012, n29013, n29014, n29015, n29016, n29017,
    n29018, n29019, n29020, n29021, n29022, n29023,
    n29024, n29025, n29026, n29027, n29028, n29029,
    n29030, n29031, n29032, n29033, n29034, n29035,
    n29036, n29037, n29038, n29039, n29040, n29041,
    n29042, n29043, n29044, n29045, n29046, n29047,
    n29048, n29049, n29050, n29051, n29052, n29053,
    n29054, n29055, n29056, n29057, n29058, n29059,
    n29060, n29061, n29062, n29063, n29064, n29065,
    n29066, n29067, n29068, n29069, n29070, n29071,
    n29072, n29073, n29074, n29075, n29076, n29077,
    n29078, n29079, n29080, n29081, n29082, n29083,
    n29084, n29085, n29086, n29087, n29088, n29089,
    n29090, n29091, n29092, n29093, n29094, n29095,
    n29096, n29097, n29098, n29099, n29100, n29101,
    n29102, n29103, n29104, n29105, n29106, n29107,
    n29108, n29109, n29110, n29111, n29112, n29113,
    n29114, n29115, n29116, n29117, n29118, n29119,
    n29120, n29121, n29122, n29123, n29124, n29125,
    n29126, n29127, n29128, n29129, n29130, n29131,
    n29132, n29133, n29134, n29135, n29136, n29137,
    n29138, n29139, n29140, n29141, n29142, n29143,
    n29144, n29145, n29146, n29147, n29148, n29149,
    n29150, n29151, n29152, n29153, n29154, n29155,
    n29156, n29157, n29158, n29159, n29160, n29161,
    n29162, n29163, n29164, n29165, n29166, n29167,
    n29168, n29169, n29170, n29171, n29172, n29173,
    n29174, n29175, n29176, n29177, n29178, n29179,
    n29180, n29181, n29182, n29183, n29184, n29185,
    n29186, n29187, n29188, n29189, n29190, n29191,
    n29192, n29193, n29194, n29195, n29196, n29197,
    n29199, n29200, n29201, n29202, n29203, n29204,
    n29205, n29206, n29207, n29208, n29209, n29210,
    n29211, n29212, n29213, n29214, n29215, n29216,
    n29217, n29218, n29219, n29220, n29221, n29222,
    n29223, n29224, n29225, n29226, n29227, n29228,
    n29229, n29230, n29231, n29232, n29233, n29234,
    n29235, n29236, n29237, n29238, n29239, n29240,
    n29241, n29242, n29243, n29244, n29245, n29246,
    n29247, n29248, n29249, n29250, n29251, n29252,
    n29253, n29254, n29255, n29256, n29257, n29258,
    n29259, n29260, n29261, n29262, n29263, n29264,
    n29265, n29266, n29267, n29268, n29269, n29270,
    n29271, n29272, n29273, n29274, n29275, n29276,
    n29277, n29278, n29279, n29280, n29281, n29282,
    n29283, n29284, n29285, n29286, n29287, n29288,
    n29289, n29290, n29291, n29292, n29293, n29294,
    n29295, n29296, n29297, n29298, n29299, n29300,
    n29301, n29302, n29303, n29304, n29305, n29306,
    n29307, n29308, n29309, n29310, n29311, n29312,
    n29313, n29314, n29315, n29316, n29317, n29318,
    n29319, n29320, n29321, n29322, n29323, n29324,
    n29325, n29326, n29327, n29328, n29329, n29330,
    n29331, n29332, n29333, n29334, n29335, n29336,
    n29337, n29338, n29339, n29340, n29341, n29342,
    n29343, n29344, n29345, n29346, n29347, n29348,
    n29349, n29350, n29351, n29352, n29353, n29354,
    n29355, n29356, n29357, n29358, n29359, n29360,
    n29361, n29362, n29363, n29364, n29365, n29366,
    n29367, n29368, n29369, n29370, n29371, n29372,
    n29373, n29374, n29375, n29376, n29377, n29378,
    n29379, n29380, n29381, n29382, n29383, n29384,
    n29385, n29386, n29387, n29388, n29389, n29390,
    n29391, n29392, n29393, n29394, n29395, n29396,
    n29397, n29398, n29399, n29400, n29401, n29402,
    n29403, n29404, n29405, n29406, n29407, n29408,
    n29409, n29410, n29411, n29412, n29413, n29414,
    n29415, n29416, n29417, n29418, n29419, n29420,
    n29421, n29422, n29423, n29424, n29425, n29426,
    n29427, n29428, n29429, n29430, n29431, n29432,
    n29433, n29434, n29435, n29436, n29437, n29438,
    n29439, n29440, n29441, n29442, n29443, n29444,
    n29445, n29446, n29447, n29448, n29449, n29450,
    n29451, n29452, n29453, n29454, n29455, n29456,
    n29457, n29458, n29459, n29460, n29461, n29462,
    n29463, n29464, n29465, n29466, n29467, n29468,
    n29469, n29470, n29471, n29472, n29473, n29474,
    n29475, n29476, n29477, n29478, n29479, n29480,
    n29481, n29482, n29483, n29484, n29485, n29486,
    n29487, n29488, n29489, n29490, n29491, n29492,
    n29493, n29494, n29495, n29496, n29497, n29498,
    n29499, n29500, n29501, n29502, n29503, n29504,
    n29505, n29506, n29507, n29508, n29509, n29510,
    n29511, n29512, n29513, n29514, n29515, n29516,
    n29517, n29518, n29519, n29520, n29521, n29522,
    n29523, n29524, n29525, n29526, n29527, n29528,
    n29529, n29530, n29531, n29532, n29533, n29534,
    n29535, n29536, n29537, n29538, n29539, n29540,
    n29541, n29542, n29543, n29544, n29545, n29546,
    n29547, n29548, n29549, n29550, n29551, n29552,
    n29553, n29554, n29555, n29556, n29557, n29558,
    n29559, n29560, n29561, n29562, n29563, n29564,
    n29565, n29566, n29567, n29568, n29569, n29570,
    n29571, n29572, n29573, n29574, n29575, n29576,
    n29577, n29578, n29579, n29580, n29581, n29582,
    n29583, n29584, n29585, n29586, n29587, n29588,
    n29589, n29590, n29591, n29592, n29593, n29594,
    n29595, n29596, n29597, n29598, n29599, n29600,
    n29601, n29602, n29603, n29604, n29605, n29606,
    n29607, n29608, n29609, n29610, n29611, n29612,
    n29613, n29614, n29615, n29616, n29617, n29618,
    n29619, n29620, n29621, n29622, n29623, n29624,
    n29625, n29626, n29627, n29628, n29629, n29630,
    n29631, n29632, n29633, n29634, n29635, n29636,
    n29637, n29638, n29639, n29640, n29641, n29642,
    n29643, n29644, n29645, n29646, n29647, n29648,
    n29649, n29650, n29651, n29652, n29653, n29654,
    n29655, n29656, n29657, n29658, n29659, n29660,
    n29661, n29662, n29663, n29664, n29665, n29666,
    n29667, n29668, n29669, n29670, n29672, n29673,
    n29674, n29675, n29676, n29677, n29678, n29679,
    n29680, n29681, n29682, n29683, n29684, n29685,
    n29686, n29687, n29688, n29689, n29690, n29691,
    n29692, n29693, n29694, n29695, n29696, n29697,
    n29698, n29699, n29700, n29701, n29702, n29703,
    n29704, n29705, n29706, n29707, n29708, n29709,
    n29710, n29711, n29712, n29713, n29714, n29715,
    n29716, n29717, n29718, n29719, n29720, n29721,
    n29722, n29723, n29724, n29725, n29726, n29727,
    n29728, n29729, n29730, n29731, n29732, n29733,
    n29734, n29735, n29736, n29737, n29738, n29739,
    n29740, n29741, n29742, n29743, n29744, n29745,
    n29746, n29747, n29748, n29749, n29750, n29751,
    n29752, n29753, n29754, n29755, n29756, n29757,
    n29758, n29759, n29760, n29761, n29762, n29763,
    n29764, n29765, n29766, n29767, n29768, n29769,
    n29770, n29771, n29772, n29773, n29774, n29775,
    n29776, n29777, n29778, n29779, n29780, n29781,
    n29782, n29783, n29784, n29785, n29786, n29787,
    n29788, n29789, n29790, n29791, n29792, n29793,
    n29794, n29795, n29796, n29797, n29798, n29799,
    n29800, n29801, n29802, n29803, n29804, n29805,
    n29806, n29807, n29808, n29809, n29810, n29811,
    n29812, n29813, n29814, n29815, n29816, n29817,
    n29818, n29819, n29820, n29821, n29822, n29823,
    n29824, n29825, n29826, n29827, n29828, n29829,
    n29830, n29831, n29832, n29833, n29834, n29835,
    n29836, n29837, n29838, n29839, n29840, n29841,
    n29842, n29843, n29844, n29845, n29846, n29847,
    n29848, n29849, n29850, n29851, n29852, n29853,
    n29854, n29855, n29856, n29857, n29858, n29859,
    n29860, n29861, n29862, n29863, n29864, n29865,
    n29866, n29867, n29868, n29869, n29870, n29871,
    n29872, n29873, n29874, n29875, n29876, n29877,
    n29878, n29879, n29880, n29881, n29882, n29883,
    n29884, n29885, n29886, n29887, n29888, n29889,
    n29890, n29891, n29892, n29893, n29894, n29895,
    n29896, n29897, n29898, n29899, n29900, n29901,
    n29902, n29903, n29904, n29905, n29906, n29907,
    n29908, n29909, n29910, n29911, n29912, n29913,
    n29914, n29915, n29916, n29917, n29918, n29919,
    n29920, n29921, n29922, n29923, n29924, n29925,
    n29926, n29927, n29928, n29929, n29930, n29931,
    n29932, n29933, n29934, n29935, n29936, n29937,
    n29938, n29939, n29940, n29941, n29942, n29943,
    n29944, n29945, n29946, n29947, n29948, n29949,
    n29950, n29951, n29952, n29953, n29954, n29955,
    n29956, n29957, n29958, n29959, n29960, n29961,
    n29962, n29963, n29964, n29965, n29966, n29967,
    n29968, n29969, n29970, n29971, n29972, n29973,
    n29974, n29975, n29976, n29977, n29978, n29979,
    n29980, n29981, n29982, n29983, n29984, n29985,
    n29986, n29987, n29988, n29989, n29990, n29991,
    n29992, n29993, n29994, n29995, n29996, n29997,
    n29998, n29999, n30000, n30001, n30002, n30003,
    n30004, n30005, n30006, n30007, n30008, n30009,
    n30010, n30011, n30012, n30013, n30014, n30015,
    n30016, n30017, n30018, n30019, n30020, n30021,
    n30022, n30023, n30024, n30025, n30026, n30027,
    n30028, n30029, n30030, n30031, n30032, n30033,
    n30034, n30035, n30036, n30037, n30038, n30039,
    n30040, n30041, n30042, n30043, n30044, n30045,
    n30046, n30047, n30048, n30049, n30050, n30051,
    n30052, n30053, n30054, n30055, n30056, n30057,
    n30058, n30059, n30060, n30061, n30062, n30063,
    n30064, n30065, n30066, n30067, n30068, n30069,
    n30070, n30071, n30072, n30073, n30074, n30075,
    n30076, n30077, n30078, n30079, n30080, n30081,
    n30082, n30083, n30084, n30085, n30086, n30087,
    n30088, n30089, n30090, n30091, n30092, n30093,
    n30094, n30095, n30096, n30097, n30098, n30099,
    n30100, n30101, n30102, n30103, n30104, n30105,
    n30106, n30107, n30108, n30109, n30110, n30111,
    n30112, n30113, n30114, n30115, n30116, n30117,
    n30118, n30119, n30120, n30121, n30122, n30123,
    n30124, n30125, n30126, n30127, n30128, n30129,
    n30130, n30131, n30132, n30133, n30134, n30135,
    n30136, n30137, n30138, n30139, n30140, n30141,
    n30142, n30143, n30145, n30146, n30147, n30148,
    n30149, n30150, n30151, n30152, n30153, n30154,
    n30155, n30156, n30157, n30158, n30159, n30160,
    n30161, n30162, n30163, n30164, n30165, n30166,
    n30167, n30168, n30169, n30170, n30171, n30172,
    n30173, n30174, n30175, n30176, n30177, n30178,
    n30179, n30180, n30181, n30182, n30183, n30184,
    n30185, n30186, n30187, n30188, n30189, n30190,
    n30191, n30192, n30193, n30194, n30195, n30196,
    n30197, n30198, n30199, n30200, n30201, n30202,
    n30203, n30204, n30205, n30206, n30207, n30208,
    n30209, n30210, n30211, n30212, n30213, n30214,
    n30215, n30216, n30217, n30218, n30219, n30220,
    n30221, n30222, n30223, n30224, n30225, n30226,
    n30227, n30228, n30229, n30230, n30231, n30232,
    n30233, n30234, n30235, n30236, n30237, n30238,
    n30239, n30240, n30241, n30242, n30243, n30244,
    n30245, n30246, n30247, n30248, n30249, n30250,
    n30251, n30252, n30253, n30254, n30255, n30256,
    n30257, n30258, n30259, n30260, n30261, n30262,
    n30263, n30264, n30265, n30266, n30267, n30268,
    n30269, n30270, n30271, n30272, n30273, n30274,
    n30275, n30276, n30277, n30278, n30279, n30280,
    n30281, n30282, n30283, n30284, n30285, n30286,
    n30287, n30288, n30289, n30290, n30291, n30292,
    n30293, n30294, n30295, n30296, n30297, n30298,
    n30299, n30300, n30301, n30302, n30303, n30304,
    n30305, n30306, n30307, n30308, n30309, n30310,
    n30311, n30312, n30313, n30314, n30315, n30316,
    n30317, n30318, n30319, n30320, n30321, n30322,
    n30323, n30324, n30325, n30326, n30327, n30328,
    n30329, n30330, n30331, n30332, n30333, n30334,
    n30335, n30336, n30337, n30338, n30339, n30340,
    n30341, n30342, n30343, n30344, n30345, n30346,
    n30347, n30348, n30349, n30350, n30351, n30352,
    n30353, n30354, n30355, n30356, n30357, n30358,
    n30359, n30360, n30361, n30362, n30363, n30364,
    n30365, n30366, n30367, n30368, n30369, n30370,
    n30371, n30372, n30373, n30374, n30375, n30376,
    n30377, n30378, n30379, n30380, n30381, n30382,
    n30383, n30384, n30385, n30386, n30387, n30388,
    n30389, n30390, n30391, n30392, n30393, n30394,
    n30395, n30396, n30397, n30398, n30399, n30400,
    n30401, n30402, n30403, n30404, n30405, n30406,
    n30407, n30408, n30409, n30410, n30411, n30412,
    n30413, n30414, n30415, n30416, n30417, n30418,
    n30419, n30420, n30421, n30422, n30423, n30424,
    n30425, n30426, n30427, n30428, n30429, n30430,
    n30431, n30432, n30433, n30434, n30435, n30436,
    n30437, n30438, n30439, n30440, n30441, n30442,
    n30443, n30444, n30445, n30446, n30447, n30448,
    n30449, n30450, n30451, n30452, n30453, n30454,
    n30455, n30456, n30457, n30458, n30459, n30460,
    n30461, n30462, n30463, n30464, n30465, n30466,
    n30467, n30468, n30469, n30470, n30471, n30472,
    n30473, n30474, n30475, n30476, n30477, n30478,
    n30479, n30480, n30481, n30482, n30483, n30484,
    n30485, n30486, n30487, n30488, n30489, n30490,
    n30491, n30492, n30493, n30494, n30495, n30496,
    n30497, n30498, n30499, n30500, n30501, n30502,
    n30503, n30504, n30505, n30506, n30507, n30508,
    n30509, n30510, n30511, n30512, n30513, n30514,
    n30515, n30516, n30517, n30518, n30519, n30520,
    n30521, n30522, n30523, n30524, n30525, n30526,
    n30527, n30528, n30529, n30530, n30531, n30532,
    n30533, n30534, n30535, n30536, n30537, n30538,
    n30539, n30540, n30541, n30542, n30543, n30544,
    n30545, n30546, n30547, n30548, n30549, n30550,
    n30551, n30552, n30553, n30554, n30555, n30556,
    n30557, n30558, n30559, n30560, n30561, n30562,
    n30563, n30564, n30565, n30566, n30567, n30568,
    n30569, n30570, n30571, n30572, n30573, n30574,
    n30575, n30576, n30577, n30578, n30579, n30580,
    n30581, n30582, n30583, n30584, n30585, n30586,
    n30587, n30588, n30589, n30590, n30591, n30592,
    n30593, n30594, n30595, n30596, n30597, n30598,
    n30599, n30600, n30601, n30602, n30603, n30604,
    n30605, n30606, n30607, n30608, n30609, n30610,
    n30611, n30612, n30613, n30614, n30615, n30616,
    n30617, n30618, n30619, n30620, n30622, n30623,
    n30624, n30625, n30626, n30627, n30628, n30629,
    n30630, n30631, n30632, n30633, n30634, n30635,
    n30636, n30637, n30638, n30639, n30640, n30641,
    n30642, n30643, n30644, n30645, n30646, n30647,
    n30648, n30649, n30650, n30651, n30652, n30653,
    n30654, n30655, n30656, n30657, n30658, n30659,
    n30660, n30661, n30662, n30663, n30664, n30665,
    n30666, n30667, n30668, n30669, n30670, n30671,
    n30672, n30673, n30674, n30675, n30676, n30677,
    n30678, n30679, n30680, n30681, n30682, n30683,
    n30684, n30685, n30686, n30687, n30688, n30689,
    n30690, n30691, n30692, n30693, n30694, n30695,
    n30696, n30697, n30698, n30699, n30700, n30701,
    n30702, n30703, n30704, n30705, n30706, n30707,
    n30708, n30709, n30710, n30711, n30712, n30713,
    n30714, n30715, n30716, n30717, n30718, n30719,
    n30720, n30721, n30722, n30723, n30724, n30725,
    n30726, n30727, n30728, n30729, n30730, n30731,
    n30732, n30733, n30734, n30735, n30736, n30737,
    n30738, n30739, n30740, n30741, n30742, n30743,
    n30744, n30745, n30746, n30747, n30748, n30749,
    n30750, n30751, n30752, n30753, n30754, n30755,
    n30756, n30757, n30758, n30759, n30760, n30761,
    n30762, n30763, n30764, n30765, n30766, n30767,
    n30768, n30769, n30770, n30771, n30772, n30773,
    n30774, n30775, n30776, n30777, n30778, n30779,
    n30780, n30781, n30782, n30783, n30784, n30785,
    n30786, n30787, n30788, n30789, n30790, n30791,
    n30792, n30793, n30794, n30795, n30796, n30797,
    n30798, n30799, n30800, n30801, n30802, n30803,
    n30804, n30805, n30806, n30807, n30808, n30809,
    n30810, n30811, n30812, n30813, n30814, n30815,
    n30816, n30817, n30818, n30819, n30820, n30821,
    n30822, n30823, n30824, n30825, n30826, n30827,
    n30828, n30829, n30830, n30831, n30832, n30833,
    n30834, n30835, n30836, n30837, n30838, n30839,
    n30840, n30841, n30842, n30843, n30844, n30845,
    n30846, n30847, n30848, n30849, n30850, n30851,
    n30852, n30853, n30854, n30855, n30856, n30857,
    n30858, n30859, n30860, n30861, n30862, n30863,
    n30864, n30865, n30866, n30867, n30868, n30869,
    n30870, n30871, n30872, n30873, n30874, n30875,
    n30876, n30877, n30878, n30879, n30880, n30881,
    n30882, n30883, n30884, n30885, n30886, n30887,
    n30888, n30889, n30890, n30891, n30892, n30893,
    n30894, n30895, n30896, n30897, n30898, n30899,
    n30900, n30901, n30902, n30903, n30904, n30905,
    n30906, n30907, n30908, n30909, n30910, n30911,
    n30912, n30913, n30914, n30915, n30916, n30917,
    n30918, n30919, n30920, n30921, n30922, n30923,
    n30924, n30925, n30926, n30927, n30928, n30929,
    n30930, n30931, n30932, n30933, n30934, n30935,
    n30936, n30937, n30938, n30939, n30940, n30941,
    n30942, n30943, n30944, n30945, n30946, n30947,
    n30948, n30949, n30950, n30951, n30952, n30953,
    n30954, n30955, n30956, n30957, n30958, n30959,
    n30960, n30961, n30962, n30963, n30964, n30965,
    n30966, n30967, n30968, n30969, n30970, n30971,
    n30972, n30973, n30974, n30975, n30976, n30977,
    n30978, n30979, n30980, n30981, n30982, n30983,
    n30984, n30985, n30986, n30987, n30988, n30989,
    n30990, n30991, n30992, n30993, n30994, n30995,
    n30996, n30997, n30998, n30999, n31000, n31001,
    n31002, n31003, n31004, n31005, n31006, n31007,
    n31008, n31009, n31010, n31011, n31012, n31013,
    n31014, n31015, n31016, n31017, n31018, n31019,
    n31020, n31021, n31022, n31023, n31024, n31025,
    n31026, n31027, n31028, n31029, n31030, n31031,
    n31032, n31033, n31034, n31035, n31036, n31037,
    n31038, n31039, n31040, n31041, n31042, n31043,
    n31044, n31045, n31046, n31047, n31048, n31049,
    n31050, n31051, n31052, n31053, n31054, n31055,
    n31056, n31057, n31058, n31059, n31060, n31061,
    n31062, n31063, n31064, n31065, n31066, n31067,
    n31068, n31069, n31070, n31071, n31072, n31073,
    n31074, n31075, n31076, n31077, n31078, n31079,
    n31080, n31081, n31082, n31083, n31084, n31085,
    n31086, n31087, n31088, n31089, n31090, n31091,
    n31092, n31093, n31094, n31095, n31097, n31098,
    n31099, n31100, n31101, n31102, n31103, n31104,
    n31105, n31106, n31107, n31108, n31109, n31110,
    n31111, n31112, n31113, n31114, n31115, n31116,
    n31117, n31118, n31119, n31120, n31121, n31122,
    n31123, n31124, n31125, n31126, n31127, n31128,
    n31129, n31130, n31131, n31132, n31133, n31134,
    n31135, n31136, n31137, n31138, n31139, n31140,
    n31141, n31142, n31143, n31144, n31145, n31146,
    n31147, n31148, n31149, n31150, n31151, n31152,
    n31153, n31154, n31155, n31156, n31157, n31158,
    n31159, n31160, n31161, n31162, n31163, n31164,
    n31165, n31166, n31167, n31168, n31169, n31170,
    n31171, n31172, n31173, n31174, n31175, n31176,
    n31177, n31178, n31179, n31180, n31181, n31182,
    n31183, n31184, n31185, n31186, n31187, n31188,
    n31189, n31190, n31191, n31192, n31193, n31194,
    n31195, n31196, n31197, n31198, n31199, n31200,
    n31201, n31202, n31203, n31204, n31205, n31206,
    n31207, n31208, n31209, n31210, n31211, n31212,
    n31213, n31214, n31215, n31216, n31217, n31218,
    n31219, n31220, n31221, n31222, n31223, n31224,
    n31225, n31226, n31227, n31228, n31229, n31230,
    n31231, n31232, n31233, n31234, n31235, n31236,
    n31237, n31238, n31239, n31240, n31241, n31242,
    n31243, n31244, n31245, n31246, n31247, n31248,
    n31249, n31250, n31251, n31252, n31253, n31254,
    n31255, n31256, n31257, n31258, n31259, n31260,
    n31261, n31262, n31263, n31264, n31265, n31266,
    n31267, n31268, n31269, n31270, n31271, n31272,
    n31273, n31274, n31275, n31276, n31277, n31278,
    n31279, n31280, n31281, n31282, n31283, n31284,
    n31285, n31286, n31287, n31288, n31289, n31290,
    n31291, n31292, n31293, n31294, n31295, n31296,
    n31297, n31298, n31299, n31300, n31301, n31302,
    n31303, n31304, n31305, n31306, n31307, n31308,
    n31309, n31310, n31311, n31312, n31313, n31314,
    n31315, n31316, n31317, n31318, n31319, n31320,
    n31321, n31322, n31323, n31324, n31325, n31326,
    n31327, n31328, n31329, n31330, n31331, n31332,
    n31333, n31334, n31335, n31336, n31337, n31338,
    n31339, n31340, n31341, n31342, n31343, n31344,
    n31345, n31346, n31347, n31348, n31349, n31350,
    n31351, n31352, n31353, n31354, n31355, n31356,
    n31357, n31358, n31359, n31360, n31361, n31362,
    n31363, n31364, n31365, n31366, n31367, n31368,
    n31369, n31370, n31371, n31372, n31373, n31374,
    n31375, n31376, n31377, n31378, n31379, n31380,
    n31381, n31382, n31383, n31384, n31385, n31386,
    n31387, n31388, n31389, n31390, n31391, n31392,
    n31393, n31394, n31395, n31396, n31397, n31398,
    n31399, n31400, n31401, n31402, n31403, n31404,
    n31405, n31406, n31407, n31408, n31409, n31410,
    n31411, n31412, n31413, n31414, n31415, n31416,
    n31417, n31418, n31419, n31420, n31421, n31422,
    n31423, n31424, n31425, n31426, n31427, n31428,
    n31429, n31430, n31431, n31432, n31433, n31434,
    n31435, n31436, n31437, n31438, n31439, n31440,
    n31441, n31442, n31443, n31444, n31445, n31446,
    n31447, n31448, n31449, n31450, n31451, n31452,
    n31453, n31454, n31455, n31456, n31457, n31458,
    n31459, n31460, n31461, n31462, n31463, n31464,
    n31465, n31466, n31467, n31468, n31469, n31470,
    n31471, n31472, n31473, n31474, n31475, n31476,
    n31477, n31478, n31479, n31480, n31481, n31482,
    n31483, n31484, n31485, n31486, n31487, n31488,
    n31489, n31490, n31491, n31492, n31493, n31494,
    n31495, n31496, n31497, n31498, n31499, n31500,
    n31501, n31502, n31503, n31504, n31505, n31506,
    n31507, n31508, n31509, n31510, n31511, n31512,
    n31513, n31514, n31515, n31516, n31517, n31518,
    n31519, n31520, n31521, n31522, n31523, n31524,
    n31525, n31526, n31527, n31528, n31529, n31530,
    n31531, n31532, n31533, n31534, n31535, n31536,
    n31537, n31538, n31539, n31540, n31541, n31542,
    n31543, n31544, n31545, n31546, n31547, n31548,
    n31549, n31550, n31551, n31552, n31553, n31554,
    n31555, n31556, n31557, n31558, n31559, n31560,
    n31561, n31562, n31563, n31564, n31565, n31566,
    n31567, n31568, n31569, n31570, n31572, n31573,
    n31574, n31575, n31576, n31577, n31578, n31579,
    n31580, n31581, n31582, n31583, n31584, n31585,
    n31586, n31587, n31588, n31589, n31590, n31591,
    n31592, n31593, n31594, n31595, n31596, n31597,
    n31598, n31599, n31600, n31601, n31602, n31603,
    n31604, n31605, n31606, n31607, n31608, n31609,
    n31610, n31611, n31612, n31613, n31614, n31615,
    n31616, n31617, n31618, n31619, n31620, n31621,
    n31622, n31623, n31624, n31625, n31626, n31627,
    n31628, n31629, n31630, n31631, n31632, n31633,
    n31634, n31635, n31636, n31637, n31638, n31639,
    n31640, n31641, n31642, n31643, n31644, n31645,
    n31646, n31647, n31648, n31649, n31650, n31651,
    n31652, n31653, n31654, n31655, n31656, n31657,
    n31658, n31659, n31660, n31661, n31662, n31663,
    n31664, n31665, n31666, n31667, n31668, n31669,
    n31670, n31671, n31672, n31673, n31674, n31675,
    n31676, n31677, n31678, n31679, n31680, n31681,
    n31682, n31683, n31684, n31685, n31686, n31687,
    n31688, n31689, n31690, n31691, n31692, n31693,
    n31694, n31695, n31696, n31697, n31698, n31699,
    n31700, n31701, n31702, n31703, n31704, n31705,
    n31706, n31707, n31708, n31709, n31710, n31711,
    n31712, n31713, n31714, n31715, n31716, n31717,
    n31718, n31719, n31720, n31721, n31722, n31723,
    n31724, n31725, n31726, n31727, n31728, n31729,
    n31730, n31731, n31732, n31733, n31734, n31735,
    n31736, n31737, n31738, n31739, n31740, n31741,
    n31742, n31743, n31744, n31745, n31746, n31747,
    n31748, n31749, n31750, n31751, n31752, n31753,
    n31754, n31755, n31756, n31757, n31758, n31759,
    n31760, n31761, n31762, n31763, n31764, n31765,
    n31766, n31767, n31768, n31769, n31770, n31771,
    n31772, n31773, n31774, n31775, n31776, n31777,
    n31778, n31779, n31780, n31781, n31782, n31783,
    n31784, n31785, n31786, n31787, n31788, n31789,
    n31790, n31791, n31792, n31793, n31794, n31795,
    n31796, n31797, n31798, n31799, n31800, n31801,
    n31802, n31803, n31804, n31805, n31806, n31807,
    n31808, n31809, n31810, n31811, n31812, n31813,
    n31814, n31815, n31816, n31817, n31818, n31819,
    n31820, n31821, n31822, n31823, n31824, n31825,
    n31826, n31827, n31828, n31829, n31830, n31831,
    n31832, n31833, n31834, n31835, n31836, n31837,
    n31838, n31839, n31840, n31841, n31842, n31843,
    n31844, n31845, n31846, n31847, n31848, n31849,
    n31850, n31851, n31852, n31853, n31854, n31855,
    n31856, n31857, n31858, n31859, n31860, n31861,
    n31862, n31863, n31864, n31865, n31866, n31867,
    n31868, n31869, n31870, n31871, n31872, n31873,
    n31874, n31875, n31876, n31877, n31878, n31879,
    n31880, n31881, n31882, n31883, n31884, n31885,
    n31886, n31887, n31888, n31889, n31890, n31891,
    n31892, n31893, n31894, n31895, n31896, n31897,
    n31898, n31899, n31900, n31901, n31902, n31903,
    n31904, n31905, n31906, n31907, n31908, n31909,
    n31910, n31911, n31912, n31913, n31914, n31915,
    n31916, n31917, n31918, n31919, n31920, n31921,
    n31922, n31923, n31924, n31925, n31926, n31927,
    n31928, n31929, n31930, n31931, n31932, n31933,
    n31934, n31935, n31936, n31937, n31938, n31939,
    n31940, n31941, n31942, n31943, n31944, n31945,
    n31946, n31947, n31948, n31949, n31950, n31951,
    n31952, n31953, n31954, n31955, n31956, n31957,
    n31958, n31959, n31960, n31961, n31962, n31963,
    n31964, n31965, n31966, n31967, n31968, n31969,
    n31970, n31971, n31972, n31973, n31974, n31975,
    n31976, n31977, n31978, n31979, n31980, n31981,
    n31982, n31983, n31984, n31985, n31986, n31987,
    n31988, n31989, n31990, n31991, n31992, n31993,
    n31994, n31995, n31996, n31997, n31998, n31999,
    n32000, n32001, n32002, n32003, n32004, n32005,
    n32006, n32007, n32008, n32009, n32010, n32011,
    n32012, n32013, n32014, n32015, n32016, n32017,
    n32018, n32019, n32020, n32021, n32022, n32023,
    n32024, n32025, n32026, n32027, n32028, n32029,
    n32030, n32031, n32032, n32033, n32034, n32035,
    n32036, n32037, n32038, n32039, n32040, n32041,
    n32042, n32043, n32044, n32045, n32047, n32048,
    n32049, n32050, n32051, n32052, n32053, n32054,
    n32055, n32056, n32057, n32058, n32059, n32060,
    n32061, n32062, n32063, n32064, n32065, n32066,
    n32067, n32068, n32069, n32070, n32071, n32072,
    n32073, n32074, n32075, n32076, n32077, n32078,
    n32079, n32080, n32081, n32082, n32083, n32084,
    n32085, n32086, n32087, n32088, n32089, n32090,
    n32091, n32092, n32093, n32094, n32095, n32096,
    n32097, n32098, n32099, n32100, n32101, n32102,
    n32103, n32104, n32105, n32106, n32107, n32108,
    n32109, n32110, n32111, n32112, n32113, n32114,
    n32115, n32116, n32117, n32118, n32119, n32120,
    n32121, n32122, n32123, n32124, n32125, n32126,
    n32127, n32128, n32129, n32130, n32131, n32132,
    n32133, n32134, n32135, n32136, n32137, n32138,
    n32139, n32140, n32141, n32142, n32143, n32144,
    n32145, n32146, n32147, n32148, n32149, n32150,
    n32151, n32152, n32153, n32154, n32155, n32156,
    n32157, n32158, n32159, n32160, n32161, n32162,
    n32163, n32164, n32165, n32166, n32167, n32168,
    n32169, n32170, n32171, n32172, n32173, n32174,
    n32175, n32176, n32177, n32178, n32179, n32180,
    n32181, n32182, n32183, n32184, n32185, n32186,
    n32187, n32188, n32189, n32190, n32191, n32192,
    n32193, n32194, n32195, n32196, n32197, n32198,
    n32199, n32200, n32201, n32202, n32203, n32204,
    n32205, n32206, n32207, n32208, n32209, n32210,
    n32211, n32212, n32213, n32214, n32215, n32216,
    n32217, n32218, n32219, n32220, n32221, n32222,
    n32223, n32224, n32225, n32226, n32227, n32228,
    n32229, n32230, n32231, n32232, n32233, n32234,
    n32235, n32236, n32237, n32238, n32239, n32240,
    n32241, n32242, n32243, n32244, n32245, n32246,
    n32247, n32248, n32249, n32250, n32251, n32252,
    n32253, n32254, n32255, n32256, n32257, n32258,
    n32259, n32260, n32261, n32262, n32263, n32264,
    n32265, n32266, n32267, n32268, n32269, n32270,
    n32271, n32272, n32273, n32274, n32275, n32276,
    n32277, n32278, n32279, n32280, n32281, n32282,
    n32283, n32284, n32285, n32286, n32287, n32288,
    n32289, n32290, n32291, n32292, n32293, n32294,
    n32295, n32296, n32297, n32298, n32299, n32300,
    n32301, n32302, n32303, n32304, n32305, n32306,
    n32307, n32308, n32309, n32310, n32311, n32312,
    n32313, n32314, n32315, n32316, n32317, n32318,
    n32319, n32320, n32321, n32322, n32323, n32324,
    n32325, n32326, n32327, n32328, n32329, n32330,
    n32331, n32332, n32333, n32334, n32335, n32336,
    n32337, n32338, n32339, n32340, n32341, n32342,
    n32343, n32344, n32345, n32346, n32347, n32348,
    n32349, n32350, n32351, n32352, n32353, n32354,
    n32355, n32356, n32357, n32358, n32359, n32360,
    n32361, n32362, n32363, n32364, n32365, n32366,
    n32367, n32368, n32369, n32370, n32371, n32372,
    n32373, n32374, n32375, n32376, n32377, n32378,
    n32379, n32380, n32381, n32382, n32383, n32384,
    n32385, n32386, n32387, n32388, n32389, n32390,
    n32391, n32392, n32393, n32394, n32395, n32396,
    n32397, n32398, n32399, n32400, n32401, n32402,
    n32403, n32404, n32405, n32406, n32407, n32408,
    n32409, n32410, n32411, n32412, n32413, n32414,
    n32415, n32416, n32417, n32418, n32419, n32420,
    n32421, n32422, n32423, n32424, n32425, n32426,
    n32427, n32428, n32429, n32430, n32431, n32432,
    n32433, n32434, n32435, n32436, n32437, n32438,
    n32439, n32440, n32441, n32442, n32443, n32444,
    n32445, n32446, n32447, n32448, n32449, n32450,
    n32451, n32452, n32453, n32454, n32455, n32456,
    n32457, n32458, n32459, n32460, n32461, n32462,
    n32463, n32464, n32465, n32466, n32467, n32468,
    n32469, n32470, n32471, n32472, n32473, n32474,
    n32475, n32476, n32477, n32478, n32479, n32480,
    n32481, n32482, n32483, n32484, n32485, n32486,
    n32487, n32488, n32489, n32490, n32491, n32492,
    n32493, n32494, n32495, n32496, n32497, n32498,
    n32499, n32500, n32501, n32502, n32503, n32504,
    n32505, n32506, n32507, n32508, n32509, n32510,
    n32511, n32512, n32513, n32514, n32515, n32517,
    n32518, n32519, n32520, n32521, n32522, n32523,
    n32524, n32525, n32526, n32527, n32528, n32529,
    n32530, n32531, n32532, n32533, n32534, n32535,
    n32536, n32537, n32538, n32539, n32540, n32541,
    n32542, n32543, n32544, n32545, n32546, n32547,
    n32548, n32549, n32550, n32551, n32552, n32553,
    n32554, n32555, n32556, n32557, n32558, n32559,
    n32560, n32561, n32562, n32563, n32564, n32565,
    n32566, n32567, n32568, n32569, n32570, n32571,
    n32572, n32573, n32574, n32575, n32576, n32577,
    n32578, n32579, n32580, n32581, n32582, n32583,
    n32584, n32585, n32586, n32587, n32588, n32589,
    n32590, n32591, n32592, n32593, n32594, n32595,
    n32596, n32597, n32598, n32599, n32600, n32601,
    n32602, n32603, n32604, n32605, n32606, n32607,
    n32608, n32609, n32610, n32611, n32612, n32613,
    n32614, n32615, n32616, n32617, n32618, n32619,
    n32620, n32621, n32622, n32623, n32624, n32625,
    n32626, n32627, n32628, n32629, n32630, n32631,
    n32632, n32633, n32634, n32635, n32636, n32637,
    n32638, n32639, n32640, n32641, n32642, n32643,
    n32644, n32645, n32646, n32647, n32648, n32649,
    n32650, n32651, n32652, n32653, n32654, n32655,
    n32656, n32657, n32658, n32659, n32660, n32661,
    n32662, n32663, n32664, n32665, n32666, n32667,
    n32668, n32669, n32670, n32671, n32672, n32673,
    n32674, n32675, n32676, n32677, n32678, n32679,
    n32680, n32681, n32682, n32683, n32684, n32685,
    n32686, n32687, n32688, n32689, n32690, n32691,
    n32692, n32693, n32694, n32695, n32696, n32697,
    n32698, n32699, n32700, n32701, n32702, n32703,
    n32704, n32705, n32706, n32707, n32708, n32709,
    n32710, n32711, n32712, n32713, n32714, n32715,
    n32716, n32717, n32718, n32719, n32720, n32721,
    n32722, n32723, n32724, n32725, n32726, n32727,
    n32728, n32729, n32730, n32731, n32732, n32733,
    n32734, n32735, n32736, n32737, n32738, n32739,
    n32740, n32741, n32742, n32743, n32744, n32745,
    n32746, n32747, n32748, n32749, n32750, n32751,
    n32752, n32753, n32754, n32755, n32756, n32757,
    n32758, n32759, n32760, n32761, n32762, n32763,
    n32764, n32765, n32766, n32767, n32768, n32769,
    n32770, n32771, n32772, n32773, n32774, n32775,
    n32776, n32777, n32778, n32779, n32780, n32781,
    n32782, n32783, n32784, n32785, n32786, n32787,
    n32788, n32789, n32790, n32791, n32792, n32793,
    n32794, n32795, n32796, n32797, n32798, n32799,
    n32800, n32801, n32802, n32803, n32804, n32805,
    n32806, n32807, n32808, n32809, n32810, n32811,
    n32812, n32813, n32814, n32815, n32816, n32817,
    n32818, n32819, n32820, n32821, n32822, n32823,
    n32824, n32825, n32826, n32827, n32828, n32829,
    n32830, n32831, n32832, n32833, n32834, n32835,
    n32836, n32837, n32838, n32839, n32840, n32841,
    n32842, n32843, n32844, n32845, n32846, n32847,
    n32848, n32849, n32850, n32851, n32852, n32853,
    n32854, n32855, n32856, n32857, n32858, n32859,
    n32860, n32861, n32862, n32863, n32864, n32865,
    n32866, n32867, n32868, n32869, n32870, n32871,
    n32872, n32873, n32874, n32875, n32876, n32877,
    n32878, n32879, n32880, n32881, n32882, n32883,
    n32884, n32885, n32886, n32887, n32888, n32889,
    n32890, n32891, n32892, n32893, n32894, n32895,
    n32896, n32897, n32898, n32899, n32900, n32901,
    n32902, n32903, n32904, n32905, n32906, n32907,
    n32908, n32909, n32910, n32911, n32912, n32913,
    n32914, n32915, n32916, n32917, n32918, n32919,
    n32920, n32921, n32922, n32923, n32924, n32925,
    n32926, n32927, n32928, n32929, n32930, n32931,
    n32932, n32933, n32934, n32935, n32936, n32937,
    n32938, n32939, n32940, n32941, n32942, n32943,
    n32944, n32945, n32946, n32947, n32948, n32949,
    n32950, n32951, n32952, n32953, n32954, n32955,
    n32956, n32957, n32958, n32959, n32960, n32961,
    n32962, n32963, n32964, n32965, n32966, n32967,
    n32968, n32969, n32970, n32971, n32972, n32973,
    n32974, n32975, n32976, n32977, n32978, n32979,
    n32980, n32981, n32983, n32984, n32985, n32986,
    n32987, n32988, n32989, n32990, n32991, n32992,
    n32993, n32994, n32995, n32996, n32997, n32998,
    n32999, n33000, n33001, n33002, n33003, n33004,
    n33005, n33006, n33007, n33008, n33009, n33010,
    n33011, n33012, n33013, n33014, n33015, n33016,
    n33017, n33018, n33019, n33020, n33021, n33022,
    n33023, n33024, n33025, n33026, n33027, n33028,
    n33029, n33030, n33031, n33033, n33034, n33035,
    n33036, n33037, n33038, n33039, n33040, n33041,
    n33042, n33043, n33044, n33045, n33046, n33047,
    n33048, n33049, n33050, n33051, n33052, n33053,
    n33054, n33055, n33056, n33057, n33058, n33059,
    n33060, n33061, n33062, n33063, n33064, n33065,
    n33066, n33067, n33068, n33069, n33070, n33071,
    n33072, n33073, n33074, n33075, n33076, n33077,
    n33078, n33079, n33080, n33081, n33082, n33083,
    n33084, n33085, n33086, n33087, n33088, n33089,
    n33090, n33091, n33092, n33093, n33094, n33095,
    n33096, n33097, n33098, n33099, n33100, n33102,
    n33103, n33104, n33105, n33106, n33107, n33108,
    n33109, n33110, n33111, n33112, n33113, n33114,
    n33115, n33116, n33117, n33118, n33119, n33120,
    n33121, n33122, n33123, n33124, n33125, n33126,
    n33127, n33128, n33129, n33130, n33131, n33132,
    n33133, n33134, n33135, n33136, n33137, n33138,
    n33139, n33140, n33141, n33142, n33143, n33144,
    n33145, n33146, n33147, n33148, n33149, n33150,
    n33151, n33152, n33153, n33154, n33155, n33156,
    n33157, n33158, n33159, n33160, n33161, n33163,
    n33164, n33165, n33166, n33167, n33168, n33169,
    n33170, n33171, n33172, n33173, n33174, n33175,
    n33176, n33177, n33178, n33179, n33180, n33181,
    n33182, n33183, n33184, n33185, n33186, n33187,
    n33188, n33189, n33190, n33191, n33192, n33193,
    n33194, n33195, n33196, n33197, n33198, n33199,
    n33200, n33201, n33202, n33203, n33204, n33205,
    n33206, n33207, n33208, n33209, n33210, n33211,
    n33212, n33213, n33214, n33215, n33216, n33217,
    n33218, n33219, n33220, n33221, n33222, n33223,
    n33224, n33225, n33226, n33227, n33228, n33229,
    n33230, n33231, n33232, n33233, n33234, n33235,
    n33236, n33237, n33238, n33239, n33240, n33241,
    n33242, n33243, n33244, n33245, n33246, n33247,
    n33248, n33249, n33250, n33251, n33252, n33253,
    n33254, n33255, n33256, n33257, n33258, n33259,
    n33260, n33261, n33262, n33263, n33264, n33265,
    n33266, n33267, n33268, n33269, n33270, n33271,
    n33272, n33273, n33274, n33275, n33276, n33277,
    n33278, n33279, n33280, n33281, n33282, n33283,
    n33284, n33285, n33286, n33287, n33288, n33289,
    n33290, n33291, n33292, n33293, n33294, n33295,
    n33296, n33297, n33298, n33299, n33300, n33301,
    n33302, n33303, n33304, n33305, n33306, n33307,
    n33308, n33309, n33310, n33311, n33312, n33313,
    n33314, n33315, n33316, n33317, n33318, n33319,
    n33320, n33321, n33322, n33323, n33324, n33325,
    n33326, n33327, n33328, n33329, n33330, n33331,
    n33332, n33333, n33334, n33335, n33336, n33337,
    n33338, n33339, n33340, n33341, n33342, n33343,
    n33344, n33345, n33346, n33347, n33348, n33349,
    n33350, n33351, n33352, n33353, n33354, n33355,
    n33356, n33357, n33358, n33359, n33360, n33361,
    n33362, n33363, n33364, n33365, n33366, n33367,
    n33368, n33369, n33370, n33371, n33372, n33373,
    n33374, n33375, n33376, n33377, n33378, n33379,
    n33380, n33381, n33382, n33383, n33384, n33385,
    n33386, n33387, n33388, n33389, n33390, n33391,
    n33392, n33393, n33394, n33395, n33396, n33397,
    n33398, n33399, n33400, n33401, n33402, n33403,
    n33404, n33405, n33406, n33407, n33408, n33409,
    n33410, n33411, n33412, n33413, n33414, n33415,
    n33416, n33417, n33418, n33419, n33420, n33421,
    n33422, n33423, n33424, n33425, n33426, n33427,
    n33428, n33429, n33430, n33431, n33432, n33433,
    n33434, n33435, n33436, n33437, n33438, n33439,
    n33440, n33441, n33442, n33443, n33444, n33445,
    n33446, n33447, n33448, n33449, n33450, n33451,
    n33452, n33453, n33454, n33455, n33456, n33457,
    n33458, n33459, n33460, n33461, n33462, n33463,
    n33464, n33465, n33466, n33467, n33468, n33469,
    n33470, n33471, n33472, n33473, n33474, n33475,
    n33476, n33477, n33478, n33479, n33480, n33481,
    n33482, n33483, n33484, n33485, n33486, n33487,
    n33488, n33489, n33490, n33491, n33492, n33493,
    n33494, n33495, n33496, n33497, n33498, n33499,
    n33500, n33501, n33502, n33503, n33504, n33505,
    n33506, n33507, n33508, n33509, n33510, n33511,
    n33512, n33513, n33514, n33515, n33516, n33517,
    n33518, n33519, n33520, n33521, n33522, n33523,
    n33524, n33525, n33526, n33527, n33528, n33529,
    n33530, n33531, n33532, n33533, n33534, n33535,
    n33536, n33537, n33538, n33539, n33540, n33541,
    n33542, n33543, n33544, n33545, n33546, n33547,
    n33548, n33549, n33550, n33551, n33552, n33553,
    n33554, n33555, n33556, n33557, n33558, n33559,
    n33560, n33561, n33562, n33563, n33564, n33565,
    n33566, n33567, n33568, n33569, n33570, n33571,
    n33572, n33573, n33574, n33575, n33576, n33577,
    n33578, n33579, n33580, n33581, n33582, n33583,
    n33584, n33585, n33586, n33587, n33588, n33589,
    n33590, n33591, n33592, n33593, n33594, n33595,
    n33596, n33597, n33598, n33599, n33600, n33601,
    n33602, n33603, n33604, n33605, n33606, n33607,
    n33608, n33609, n33610, n33611, n33612, n33613,
    n33614, n33615, n33616, n33617, n33618, n33619,
    n33620, n33621, n33622, n33623, n33624, n33625,
    n33626, n33627, n33628, n33629, n33630, n33631,
    n33632, n33633, n33634, n33635, n33636, n33637,
    n33638, n33639, n33640, n33641, n33642, n33643,
    n33644, n33645, n33646, n33647, n33648, n33649,
    n33650, n33651, n33652, n33653, n33654, n33655,
    n33656, n33657, n33658, n33659, n33660, n33661,
    n33662, n33663, n33664, n33665, n33666, n33667,
    n33668, n33669, n33670, n33671, n33672, n33673,
    n33674, n33675, n33676, n33677, n33678, n33679,
    n33680, n33681, n33682, n33683, n33684, n33685,
    n33686, n33687, n33688, n33689, n33690, n33691,
    n33692, n33693, n33694, n33695, n33696, n33697,
    n33698, n33699, n33700, n33701, n33702, n33703,
    n33704, n33705, n33706, n33707, n33708, n33709,
    n33710, n33711, n33712, n33713, n33714, n33715,
    n33716, n33717, n33718, n33719, n33720, n33721,
    n33722, n33723, n33724, n33725, n33726, n33727,
    n33728, n33729, n33730, n33731, n33732, n33733,
    n33734, n33735, n33736, n33737, n33738, n33739,
    n33740, n33741, n33742, n33743, n33744, n33745,
    n33746, n33747, n33748, n33749, n33750, n33751,
    n33752, n33753, n33754, n33755, n33756, n33757,
    n33758, n33759, n33760, n33761, n33762, n33763,
    n33764, n33765, n33766, n33767, n33768, n33769,
    n33770, n33771, n33772, n33773, n33774, n33775,
    n33776, n33777, n33778, n33779, n33780, n33781,
    n33782, n33783, n33784, n33785, n33786, n33787,
    n33788, n33789, n33790, n33791, n33793, n33794,
    n33795, n33796, n33797, n33798, n33799, n33800,
    n33801, n33802, n33803, n33804, n33805, n33806,
    n33807, n33808, n33809, n33810, n33811, n33812,
    n33813, n33814, n33815, n33816, n33817, n33818,
    n33819, n33820, n33821, n33822, n33823, n33824,
    n33825, n33826, n33827, n33828, n33829, n33830,
    n33831, n33832, n33833, n33834, n33835, n33836,
    n33837, n33838, n33839, n33840, n33841, n33842,
    n33843, n33844, n33845, n33846, n33847, n33848,
    n33849, n33850, n33851, n33852, n33853, n33854,
    n33855, n33856, n33857, n33858, n33859, n33860,
    n33861, n33862, n33863, n33864, n33865, n33866,
    n33867, n33868, n33869, n33870, n33871, n33872,
    n33873, n33874, n33875, n33876, n33877, n33878,
    n33879, n33880, n33881, n33882, n33883, n33884,
    n33885, n33886, n33887, n33888, n33889, n33890,
    n33891, n33892, n33893, n33894, n33895, n33896,
    n33897, n33898, n33899, n33900, n33901, n33902,
    n33903, n33904, n33905, n33906, n33907, n33908,
    n33909, n33910, n33911, n33912, n33913, n33914,
    n33915, n33916, n33917, n33918, n33919, n33920,
    n33921, n33922, n33923, n33924, n33925, n33926,
    n33927, n33928, n33929, n33930, n33931, n33932,
    n33933, n33934, n33935, n33936, n33937, n33938,
    n33939, n33940, n33941, n33942, n33943, n33944,
    n33945, n33946, n33947, n33948, n33949, n33950,
    n33951, n33952, n33953, n33954, n33955, n33956,
    n33957, n33958, n33959, n33960, n33961, n33962,
    n33963, n33964, n33965, n33966, n33967, n33968,
    n33969, n33970, n33971, n33972, n33973, n33974,
    n33975, n33976, n33977, n33978, n33979, n33980,
    n33981, n33982, n33983, n33984, n33985, n33986,
    n33987, n33988, n33989, n33990, n33991, n33992,
    n33993, n33994, n33995, n33996, n33997, n33998,
    n33999, n34000, n34001, n34002, n34003, n34004,
    n34005, n34006, n34007, n34008, n34009, n34010,
    n34011, n34012, n34013, n34014, n34015, n34016,
    n34017, n34018, n34019, n34020, n34021, n34022,
    n34023, n34024, n34025, n34026, n34027, n34028,
    n34029, n34030, n34031, n34032, n34033, n34034,
    n34035, n34036, n34037, n34038, n34039, n34040,
    n34041, n34042, n34043, n34044, n34045, n34046,
    n34047, n34048, n34049, n34050, n34051, n34052,
    n34053, n34054, n34055, n34056, n34057, n34058,
    n34059, n34060, n34061, n34062, n34063, n34064,
    n34065, n34066, n34067, n34068, n34069, n34070,
    n34071, n34072, n34073, n34074, n34075, n34076,
    n34077, n34078, n34079, n34080, n34081, n34082,
    n34084, n34085, n34086, n34087, n34088, n34089,
    n34090, n34091, n34092, n34093, n34094, n34095,
    n34096, n34097, n34098, n34099, n34100, n34101,
    n34102, n34103, n34104, n34105, n34106, n34107,
    n34108, n34109, n34110, n34111, n34112, n34113,
    n34114, n34115, n34116, n34117, n34118, n34119,
    n34120, n34121, n34122, n34123, n34124, n34125,
    n34126, n34127, n34128, n34129, n34130, n34131,
    n34132, n34133, n34134, n34135, n34136, n34137,
    n34138, n34139, n34140, n34141, n34142, n34143,
    n34144, n34145, n34146, n34147, n34148, n34149,
    n34150, n34151, n34152, n34153, n34154, n34155,
    n34156, n34157, n34158, n34159, n34160, n34161,
    n34162, n34163, n34164, n34165, n34166, n34167,
    n34168, n34169, n34170, n34171, n34172, n34173,
    n34174, n34175, n34176, n34177, n34178, n34179,
    n34180, n34181, n34182, n34183, n34184, n34185,
    n34186, n34187, n34188, n34189, n34190, n34191,
    n34192, n34193, n34194, n34195, n34196, n34197,
    n34198, n34199, n34200, n34201, n34202, n34203,
    n34204, n34205, n34206, n34207, n34208, n34209,
    n34210, n34211, n34212, n34213, n34214, n34215,
    n34216, n34217, n34218, n34219, n34220, n34221,
    n34222, n34223, n34224, n34225, n34226, n34227,
    n34228, n34229, n34230, n34231, n34232, n34233,
    n34234, n34235, n34236, n34237, n34238, n34239,
    n34240, n34241, n34242, n34243, n34244, n34245,
    n34246, n34247, n34248, n34249, n34250, n34251,
    n34252, n34253, n34254, n34255, n34256, n34257,
    n34258, n34259, n34260, n34261, n34262, n34263,
    n34264, n34265, n34266, n34267, n34268, n34269,
    n34270, n34271, n34272, n34273, n34274, n34275,
    n34276, n34277, n34278, n34279, n34280, n34281,
    n34282, n34283, n34284, n34285, n34286, n34287,
    n34288, n34289, n34290, n34291, n34292, n34293,
    n34294, n34295, n34296, n34297, n34298, n34299,
    n34300, n34301, n34302, n34303, n34304, n34305,
    n34306, n34307, n34308, n34309, n34310, n34311,
    n34312, n34313, n34314, n34315, n34316, n34317,
    n34318, n34319, n34320, n34321, n34322, n34323,
    n34324, n34325, n34326, n34327, n34328, n34329,
    n34330, n34331, n34332, n34333, n34334, n34335,
    n34336, n34337, n34338, n34339, n34340, n34341,
    n34342, n34343, n34344, n34345, n34346, n34347,
    n34348, n34349, n34350, n34351, n34352, n34353,
    n34354, n34355, n34356, n34357, n34358, n34359,
    n34360, n34361, n34362, n34364, n34365, n34366,
    n34367, n34368, n34369, n34370, n34371, n34372,
    n34373, n34374, n34375, n34376, n34377, n34378,
    n34379, n34380, n34381, n34382, n34383, n34384,
    n34385, n34386, n34387, n34388, n34389, n34390,
    n34391, n34392, n34393, n34394, n34395, n34396,
    n34397, n34398, n34399, n34400, n34401, n34402,
    n34403, n34404, n34405, n34406, n34407, n34408,
    n34409, n34410, n34411, n34412, n34413, n34414,
    n34415, n34416, n34417, n34418, n34419, n34420,
    n34421, n34422, n34423, n34424, n34425, n34426,
    n34427, n34428, n34429, n34430, n34431, n34432,
    n34433, n34434, n34435, n34436, n34437, n34438,
    n34439, n34440, n34441, n34442, n34443, n34444,
    n34445, n34446, n34447, n34448, n34449, n34450,
    n34451, n34452, n34453, n34454, n34455, n34456,
    n34457, n34458, n34459, n34460, n34461, n34462,
    n34463, n34464, n34465, n34466, n34467, n34468,
    n34469, n34470, n34471, n34472, n34473, n34474,
    n34475, n34476, n34477, n34478, n34479, n34480,
    n34481, n34482, n34483, n34484, n34485, n34486,
    n34487, n34488, n34489, n34490, n34491, n34492,
    n34493, n34494, n34495, n34496, n34497, n34498,
    n34499, n34500, n34501, n34502, n34503, n34504,
    n34505, n34506, n34507, n34508, n34509, n34510,
    n34511, n34512, n34513, n34514, n34515, n34516,
    n34517, n34518, n34519, n34520, n34521, n34522,
    n34523, n34524, n34525, n34526, n34527, n34528,
    n34529, n34530, n34531, n34532, n34533, n34534,
    n34535, n34536, n34537, n34538, n34539, n34540,
    n34541, n34542, n34543, n34544, n34545, n34546,
    n34547, n34548, n34549, n34550, n34551, n34552,
    n34553, n34554, n34555, n34556, n34557, n34559,
    n34560, n34561, n34562, n34563, n34564, n34565,
    n34567, n34568, n34569, n34570, n34571, n34572,
    n34573, n34575, n34576, n34577, n34578, n34579,
    n34580, n34581, n34582, n34583, n34584, n34585,
    n34586, n34587, n34588, n34589, n34590, n34591,
    n34592, n34593, n34594, n34595, n34596, n34597,
    n34598, n34599, n34600, n34601, n34602, n34603,
    n34604, n34605, n34606, n34607, n34608, n34609,
    n34610, n34611, n34612, n34613, n34614, n34615,
    n34616, n34617, n34618, n34619, n34620, n34621,
    n34622, n34623, n34624, n34625, n34626, n34627,
    n34628, n34629, n34630, n34631, n34632, n34633,
    n34634, n34635, n34636, n34637, n34638, n34639,
    n34640, n34641, n34642, n34643, n34644, n34645,
    n34646, n34647, n34648, n34649, n34650, n34651,
    n34652, n34653, n34654, n34655, n34656, n34657,
    n34658, n34659, n34660, n34661, n34662, n34663,
    n34664, n34665, n34666, n34667, n34668, n34669,
    n34670, n34671, n34672, n34673, n34674, n34675,
    n34676, n34677, n34678, n34679, n34680, n34681,
    n34683, n34684, n34685, n34686, n34687, n34688,
    n34690, n34691, n34692, n34693, n34694, n34695,
    n34696, n34698, n34699, n34700, n34701, n34702,
    n34703, n34704, n34705, n34706, n34707, n34708,
    n34709, n34710, n34711, n34712, n34713, n34714,
    n34715, n34716, n34717, n34718, n34719, n34720,
    n34721, n34722, n34723, n34724, n34725, n34726,
    n34727, n34728, n34729, n34730, n34731, n34732,
    n34733, n34734, n34735, n34736, n34737, n34738,
    n34739, n34740, n34741, n34742, n34743, n34744,
    n34745, n34746, n34747, n34748, n34749, n34750,
    n34751, n34752, n34753, n34754, n34755, n34756,
    n34757, n34758, n34759, n34760, n34761, n34762,
    n34763, n34764, n34765, n34766, n34767, n34768,
    n34769, n34770, n34771, n34772, n34773, n34774,
    n34775, n34776, n34777, n34778, n34779, n34780,
    n34781, n34782, n34783, n34784, n34785, n34786,
    n34787, n34788, n34789, n34790, n34791, n34792,
    n34793, n34794, n34795, n34796, n34797, n34798,
    n34799, n34800, n34801, n34802, n34803, n34804,
    n34805, n34806, n34807, n34808, n34809, n34810,
    n34811, n34812, n34813, n34814, n34815, n34816,
    n34817, n34818, n34819, n34820, n34821, n34822,
    n34823, n34824, n34825, n34826, n34827, n34828,
    n34829, n34830, n34831, n34832, n34833, n34834,
    n34835, n34836, n34837, n34838, n34839, n34840,
    n34841, n34842, n34843, n34844, n34845, n34846,
    n34847, n34848, n34849, n34850, n34851, n34852,
    n34853, n34854, n34855, n34856, n34857, n34858,
    n34859, n34860, n34861, n34862, n34863, n34864,
    n34865, n34866, n34867, n34868, n34869, n34870,
    n34871, n34872, n34873, n34874, n34875, n34876,
    n34877, n34878, n34879, n34880, n34881, n34882,
    n34883, n34884, n34885, n34886, n34887, n34888,
    n34889, n34890, n34891, n34892, n34893, n34894,
    n34895, n34896, n34897, n34898, n34899, n34900,
    n34901, n34902, n34903, n34904, n34905, n34906,
    n34907, n34908, n34909, n34910, n34911, n34912,
    n34913, n34914, n34915, n34916, n34917, n34918,
    n34919, n34920, n34921, n34922, n34923, n34924,
    n34925, n34926, n34927, n34928, n34929, n34930,
    n34931, n34932, n34933, n34934, n34935, n34936,
    n34937, n34938, n34939, n34940, n34941, n34942,
    n34943, n34944, n34945, n34946, n34947, n34948,
    n34949, n34950, n34951, n34952, n34953, n34954,
    n34955, n34956, n34957, n34958, n34959, n34960,
    n34961, n34962, n34963, n34964, n34965, n34966,
    n34967, n34968, n34969, n34970, n34971, n34972,
    n34973, n34974, n34975, n34976, n34977, n34978,
    n34979, n34980, n34981, n34982, n34983, n34984,
    n34985, n34986, n34987, n34988, n34989, n34990,
    n34991, n34992, n34993, n34994, n34995, n34996,
    n34997, n34998, n34999, n35000, n35001, n35002,
    n35003, n35004, n35005, n35006, n35007, n35008,
    n35009, n35010, n35011, n35012, n35013, n35014,
    n35015, n35016, n35017, n35018, n35019, n35020,
    n35021, n35022, n35023, n35024, n35025, n35026,
    n35027, n35028, n35029, n35030, n35031, n35032,
    n35033, n35034, n35035, n35036, n35037, n35038,
    n35039, n35040, n35041, n35042, n35043, n35044,
    n35045, n35046, n35047, n35048, n35049, n35050,
    n35051, n35052, n35053, n35054, n35055, n35056,
    n35057, n35058, n35059, n35060, n35061, n35062,
    n35063, n35064, n35065, n35066, n35067, n35068,
    n35069, n35070, n35071, n35072, n35073, n35074,
    n35075, n35076, n35077, n35078, n35079, n35080,
    n35081, n35082, n35083, n35084, n35085, n35086,
    n35087, n35088, n35089, n35090, n35091, n35092,
    n35093, n35094, n35095, n35096, n35097, n35098,
    n35099, n35100, n35101, n35102, n35103, n35104,
    n35105, n35106, n35107, n35108, n35109, n35110,
    n35111, n35112, n35113, n35114, n35115, n35116,
    n35117, n35118, n35119, n35120, n35121, n35122,
    n35123, n35124, n35125, n35126, n35127, n35128,
    n35129, n35130, n35131, n35132, n35133, n35134,
    n35135, n35136, n35137, n35138, n35139, n35140,
    n35141, n35142, n35143, n35144, n35145, n35146,
    n35147, n35148, n35149, n35150, n35151, n35152,
    n35153, n35154, n35155, n35156, n35157, n35158,
    n35159, n35160, n35161, n35162, n35163, n35164,
    n35165, n35166, n35167, n35168, n35169, n35170,
    n35171, n35172, n35173, n35174, n35175, n35176,
    n35177, n35178, n35179, n35180, n35181, n35182,
    n35183, n35184, n35185, n35186, n35187, n35188,
    n35190, n35191, n35192, n35193, n35194, n35195,
    n35196, n35197, n35198, n35199, n35200, n35201,
    n35202, n35203, n35204, n35205, n35206, n35207,
    n35208, n35209, n35210, n35211, n35212, n35213,
    n35214, n35215, n35216, n35217, n35218, n35219,
    n35220, n35221, n35222, n35223, n35224, n35225,
    n35226, n35227, n35228, n35229, n35230, n35231,
    n35232, n35233, n35234, n35235, n35236, n35237,
    n35238, n35239, n35240, n35241, n35242, n35243,
    n35244, n35245, n35246, n35247, n35248, n35249,
    n35250, n35251, n35252, n35253, n35254, n35255,
    n35256, n35257, n35258, n35259, n35260, n35261,
    n35262, n35263, n35265, n35266, n35267, n35268,
    n35269, n35270, n35271, n35272, n35273, n35274,
    n35275, n35276, n35277, n35278, n35279, n35280,
    n35281, n35282, n35283, n35284, n35285, n35286,
    n35287, n35288, n35289, n35290, n35291, n35292,
    n35293, n35294, n35295, n35296, n35297, n35298,
    n35299, n35300, n35301, n35302, n35303, n35304,
    n35305, n35306, n35307, n35308, n35309, n35310,
    n35311, n35312, n35313, n35314, n35315, n35316,
    n35317, n35318, n35319, n35320, n35321, n35322,
    n35323, n35324, n35325, n35326, n35327, n35328,
    n35329, n35330, n35331, n35332, n35333, n35334,
    n35335, n35336, n35337, n35338, n35339, n35340,
    n35341, n35342, n35343, n35344, n35345, n35346,
    n35347, n35348, n35349, n35350, n35351, n35352,
    n35353, n35354, n35355, n35356, n35357, n35358,
    n35359, n35360, n35361, n35362, n35363, n35364,
    n35365, n35366, n35367, n35368, n35369, n35370,
    n35371, n35372, n35373, n35374, n35375, n35376,
    n35377, n35378, n35379, n35380, n35381, n35382,
    n35383, n35384, n35385, n35386, n35387, n35388,
    n35389, n35390, n35391, n35392, n35393, n35394,
    n35395, n35396, n35397, n35398, n35399, n35400,
    n35401, n35402, n35403, n35404, n35405, n35406,
    n35407, n35408, n35409, n35410, n35411, n35412,
    n35413, n35414, n35415, n35416, n35417, n35418,
    n35419, n35420, n35421, n35422, n35423, n35425,
    n35426, n35427, n35428, n35429, n35430, n35431,
    n35432, n35433, n35434, n35435, n35436, n35437,
    n35438, n35439, n35440, n35441, n35442, n35443,
    n35444, n35445, n35446, n35447, n35448, n35449,
    n35450, n35451, n35452, n35453, n35454, n35455,
    n35456, n35457, n35458, n35459, n35460, n35461,
    n35462, n35463, n35464, n35465, n35466, n35467,
    n35468, n35469, n35470, n35471, n35472, n35473,
    n35474, n35475, n35476, n35477, n35478, n35479,
    n35480, n35481, n35482, n35483, n35484, n35485,
    n35486, n35487, n35488, n35489, n35490, n35491,
    n35492, n35493, n35494, n35495, n35496, n35497,
    n35498, n35499, n35500, n35501, n35502, n35503,
    n35504, n35505, n35506, n35507, n35508, n35509,
    n35510, n35511, n35512, n35513, n35514, n35515,
    n35516, n35517, n35518, n35519, n35520, n35521,
    n35522, n35523, n35524, n35525, n35526, n35527,
    n35528, n35529, n35530, n35531, n35532, n35533,
    n35534, n35535, n35536, n35537, n35538, n35539,
    n35540, n35541, n35542, n35543, n35544, n35545,
    n35546, n35547, n35548, n35549, n35551, n35552,
    n35553, n35554, n35555, n35556, n35557, n35558,
    n35559, n35560, n35561, n35562, n35563, n35564,
    n35565, n35566, n35567, n35568, n35569, n35570,
    n35571, n35572, n35573, n35574, n35575, n35576,
    n35578, n35579, n35580, n35581, n35582, n35583,
    n35584, n35585, n35586, n35587, n35588, n35589,
    n35590, n35591, n35592, n35593, n35594, n35595,
    n35596, n35597, n35599, n35600, n35601, n35602,
    n35603, n35604, n35605, n35606, n35607, n35608,
    n35609, n35610, n35611, n35612, n35613, n35614,
    n35615, n35616, n35617, n35618, n35620, n35621,
    n35622, n35623, n35624, n35625, n35626, n35627,
    n35628, n35629, n35630, n35631, n35632, n35633,
    n35634, n35635, n35636, n35637, n35638, n35639,
    n35641, n35642, n35643, n35644, n35645, n35646,
    n35647, n35648, n35649, n35650, n35651, n35652,
    n35653, n35654, n35655, n35656, n35657, n35658,
    n35659, n35660, n35661, n35662, n35663, n35664,
    n35665, n35666, n35667, n35668, n35669, n35670,
    n35671, n35672, n35673, n35674, n35675, n35676,
    n35677, n35678, n35679, n35680, n35681, n35682,
    n35683, n35684, n35685, n35686, n35687, n35688,
    n35689, n35690, n35691, n35692, n35693, n35694,
    n35695, n35696, n35697, n35698, n35699, n35700,
    n35701, n35702, n35703, n35704, n35705, n35706,
    n35707, n35708, n35709, n35710, n35711, n35712,
    n35713, n35714, n35715, n35716, n35717, n35718,
    n35719, n35720, n35721, n35722, n35723, n35724,
    n35725, n35726, n35727, n35728, n35729, n35730,
    n35731, n35732, n35733, n35734, n35735, n35736,
    n35737, n35738, n35739, n35740, n35741, n35742,
    n35743, n35744, n35745, n35746, n35747, n35748,
    n35749, n35750, n35751, n35752, n35753, n35754,
    n35756, n35757, n35758, n35759, n35760, n35761,
    n35762, n35763, n35764, n35765, n35766, n35767,
    n35768, n35769, n35770, n35771, n35772, n35773,
    n35774, n35775, n35776, n35777, n35778, n35779,
    n35780, n35781, n35782, n35783, n35784, n35785,
    n35786, n35787, n35788, n35789, n35790, n35791,
    n35792, n35793, n35794, n35795, n35796, n35797,
    n35798, n35799, n35800, n35801, n35802, n35803,
    n35804, n35805, n35806, n35807, n35808, n35809,
    n35810, n35811, n35812, n35813, n35814, n35815,
    n35816, n35817, n35818, n35819, n35820, n35821,
    n35822, n35823, n35824, n35825, n35826, n35827,
    n35828, n35829, n35830, n35831, n35832, n35833,
    n35834, n35835, n35836, n35837, n35838, n35839,
    n35840, n35841, n35842, n35843, n35844, n35845,
    n35846, n35847, n35848, n35849, n35850, n35851,
    n35852, n35853, n35854, n35855, n35856, n35857,
    n35858, n35859, n35861, n35862, n35863, n35864,
    n35865, n35866, n35867, n35868, n35869, n35870,
    n35871, n35872, n35873, n35874, n35875, n35876,
    n35877, n35878, n35880, n35881, n35882, n35883,
    n35884, n35885, n35887, n35888, n35889, n35890,
    n35891, n35892, n35893, n35894, n35895, n35896,
    n35897, n35898, n35899, n35900, n35901, n35902,
    n35903, n35904, n35905, n35906, n35908, n35909,
    n35910, n35911, n35912, n35913, n35915, n35916,
    n35917, n35918, n35919, n35920, n35921, n35922,
    n35923, n35924, n35925, n35926, n35927, n35928,
    n35929, n35930, n35931, n35932, n35933, n35934,
    n35935, n35936, n35937, n35938, n35939, n35940,
    n35941, n35942, n35943, n35944, n35945, n35946,
    n35947, n35948, n35949, n35950, n35951, n35952,
    n35953, n35954, n35955, n35956, n35957, n35958,
    n35959, n35960, n35961, n35962, n35963, n35964,
    n35965, n35966, n35967, n35968, n35969, n35970,
    n35971, n35972, n35973, n35974, n35975, n35976,
    n35977, n35978, n35979, n35980, n35981, n35982,
    n35983, n35984, n35985, n35986, n35987, n35988,
    n35989, n35990, n35991, n35992, n35993, n35994,
    n35995, n35996, n35997, n35998, n35999, n36000,
    n36001, n36002, n36003, n36004, n36005, n36006,
    n36007, n36008, n36009, n36010, n36011, n36012,
    n36013, n36014, n36015, n36016, n36017, n36019,
    n36020, n36021, n36022, n36023, n36024, n36025,
    n36026, n36027, n36028, n36029, n36030, n36031,
    n36032, n36033, n36034, n36035, n36036, n36037,
    n36038, n36039, n36040, n36041, n36042, n36043,
    n36044, n36045, n36046, n36047, n36048, n36049,
    n36050, n36051, n36052, n36053, n36054, n36055,
    n36056, n36057, n36058, n36059, n36060, n36061,
    n36062, n36063, n36064, n36065, n36066, n36067,
    n36068, n36069, n36070, n36071, n36072, n36073,
    n36074, n36075, n36076, n36077, n36078, n36079,
    n36080, n36081, n36082, n36083, n36084, n36085,
    n36086, n36087, n36088, n36089, n36090, n36091,
    n36092, n36093, n36094, n36095, n36096, n36097,
    n36098, n36099, n36100, n36101, n36102, n36103,
    n36104, n36105, n36106, n36107, n36108, n36109,
    n36110, n36111, n36112, n36113, n36114, n36115,
    n36116, n36117, n36118, n36119, n36120, n36121,
    n36122, n36123, n36124, n36125, n36126, n36127,
    n36128, n36129, n36130, n36131, n36132, n36133,
    n36134, n36135, n36136, n36137, n36138, n36139,
    n36140, n36141, n36142, n36143, n36144, n36145,
    n36146, n36147, n36148, n36149, n36150, n36151,
    n36152, n36153, n36154, n36155, n36156, n36157,
    n36158, n36159, n36160, n36161, n36162, n36163,
    n36164, n36165, n36166, n36167, n36168, n36169,
    n36170, n36171, n36172, n36173, n36174, n36175,
    n36176, n36177, n36178, n36179, n36180, n36181,
    n36182, n36183, n36184, n36185, n36186, n36187,
    n36188, n36189, n36190, n36191, n36192, n36193,
    n36194, n36195, n36196, n36197, n36198, n36199,
    n36200, n36201, n36202, n36203, n36204, n36205,
    n36206, n36207, n36208, n36209, n36210, n36211,
    n36212, n36213, n36214, n36215, n36216, n36217,
    n36218, n36219, n36220, n36221, n36222, n36223,
    n36224, n36225, n36226, n36227, n36228, n36229,
    n36230, n36231, n36232, n36233, n36234, n36235,
    n36236, n36237, n36238, n36239, n36240, n36241,
    n36242, n36243, n36244, n36245, n36246, n36247,
    n36248, n36249, n36250, n36251, n36252, n36253,
    n36254, n36255, n36256, n36257, n36258, n36259,
    n36260, n36261, n36262, n36263, n36264, n36265,
    n36266, n36267, n36268, n36269, n36270, n36271,
    n36272, n36273, n36274, n36275, n36276, n36277,
    n36278, n36279, n36280, n36281, n36282, n36283,
    n36284, n36285, n36286, n36287, n36288, n36289,
    n36290, n36291, n36292, n36293, n36294, n36295,
    n36296, n36297, n36298, n36299, n36300, n36301,
    n36302, n36303, n36304, n36305, n36306, n36307,
    n36308, n36309, n36310, n36311, n36312, n36313,
    n36314, n36315, n36316, n36317, n36318, n36319,
    n36320, n36321, n36322, n36323, n36324, n36325,
    n36326, n36327, n36328, n36329, n36330, n36331,
    n36332, n36333, n36334, n36335, n36336, n36337,
    n36338, n36339, n36340, n36341, n36342, n36343,
    n36344, n36345, n36346, n36347, n36348, n36349,
    n36350, n36351, n36352, n36353, n36354, n36355,
    n36356, n36357, n36358, n36359, n36360, n36361,
    n36362, n36363, n36364, n36365, n36366, n36367,
    n36368, n36369, n36370, n36371, n36372, n36373,
    n36374, n36375, n36376, n36377, n36378, n36379,
    n36380, n36381, n36382, n36383, n36384, n36385,
    n36386, n36387, n36388, n36389, n36390, n36391,
    n36392, n36393, n36394, n36395, n36396, n36397,
    n36398, n36399, n36400, n36401, n36402, n36403,
    n36404, n36405, n36406, n36407, n36408, n36409,
    n36410, n36411, n36412, n36413, n36414, n36415,
    n36416, n36417, n36418, n36419, n36420, n36421,
    n36422, n36423, n36424, n36425, n36426, n36427,
    n36428, n36429, n36430, n36431, n36432, n36433,
    n36434, n36435, n36436, n36437, n36438, n36439,
    n36440, n36441, n36442, n36443, n36444, n36445,
    n36446, n36447, n36448, n36449, n36450, n36451,
    n36452, n36453, n36454, n36455, n36456, n36457,
    n36458, n36459, n36460, n36461, n36462, n36463,
    n36464, n36465, n36466, n36467, n36468, n36469,
    n36470, n36471, n36472, n36473, n36474, n36475,
    n36476, n36477, n36478, n36479, n36480, n36481,
    n36482, n36483, n36484, n36485, n36486, n36487,
    n36488, n36489, n36490, n36491, n36492, n36493,
    n36494, n36495, n36496, n36497, n36498, n36499,
    n36500, n36501, n36502, n36503, n36504, n36505,
    n36506, n36507, n36508, n36509, n36510, n36511,
    n36512, n36513, n36514, n36515, n36516, n36517,
    n36518, n36519, n36520, n36521, n36522, n36523,
    n36524, n36525, n36526, n36527, n36528, n36529,
    n36530, n36531, n36532, n36533, n36534, n36535,
    n36536, n36537, n36538, n36539, n36540, n36541,
    n36542, n36543, n36544, n36545, n36546, n36547,
    n36548, n36549, n36550, n36551, n36552, n36553,
    n36554, n36555, n36556, n36557, n36558, n36559,
    n36560, n36561, n36562, n36563, n36564, n36565,
    n36566, n36567, n36568, n36569, n36570, n36571,
    n36572, n36573, n36574, n36575, n36576, n36577,
    n36578, n36579, n36580, n36581, n36582, n36583,
    n36584, n36585, n36586, n36587, n36588, n36589,
    n36590, n36591, n36592, n36593, n36594, n36595,
    n36596, n36597, n36598, n36599, n36600, n36601,
    n36602, n36603, n36604, n36605, n36606, n36607,
    n36608, n36609, n36610, n36611, n36612, n36613,
    n36614, n36615, n36616, n36617, n36618, n36619,
    n36620, n36621, n36622, n36623, n36624, n36625,
    n36626, n36627, n36628, n36629, n36630, n36632,
    n36633, n36634, n36635, n36636, n36637, n36638,
    n36639, n36640, n36641, n36642, n36643, n36644,
    n36645, n36646, n36647, n36648, n36649, n36650,
    n36651, n36652, n36653, n36654, n36655, n36656,
    n36657, n36658, n36659, n36660, n36661, n36662,
    n36663, n36664, n36665, n36666, n36667, n36668,
    n36669, n36670, n36671, n36672, n36673, n36674,
    n36675, n36676, n36677, n36678, n36679, n36680,
    n36681, n36682, n36683, n36684, n36685, n36686,
    n36687, n36688, n36689, n36690, n36691, n36692,
    n36693, n36694, n36695, n36696, n36697, n36698,
    n36699, n36700, n36701, n36702, n36703, n36704,
    n36705, n36706, n36707, n36708, n36709, n36710,
    n36711, n36712, n36713, n36714, n36715, n36716,
    n36717, n36718, n36719, n36720, n36721, n36722,
    n36723, n36724, n36725, n36726, n36727, n36728,
    n36729, n36730, n36731, n36732, n36733, n36734,
    n36735, n36736, n36737, n36738, n36739, n36740,
    n36741, n36742, n36743, n36744, n36745, n36746,
    n36747, n36748, n36749, n36750, n36751, n36752,
    n36753, n36754, n36755, n36756, n36757, n36758,
    n36759, n36760, n36761, n36762, n36763, n36764,
    n36765, n36766, n36767, n36768, n36769, n36770,
    n36771, n36772, n36773, n36774, n36775, n36776,
    n36777, n36778, n36779, n36780, n36781, n36782,
    n36783, n36784, n36785, n36786, n36787, n36788,
    n36789, n36790, n36791, n36792, n36793, n36794,
    n36795, n36796, n36797, n36798, n36799, n36800,
    n36801, n36802, n36803, n36804, n36805, n36806,
    n36807, n36808, n36809, n36810, n36811, n36812,
    n36813, n36814, n36815, n36816, n36817, n36818,
    n36819, n36820, n36821, n36822, n36823, n36824,
    n36825, n36826, n36827, n36828, n36829, n36830,
    n36831, n36832, n36833, n36834, n36835, n36836,
    n36837, n36838, n36839, n36840, n36841, n36842,
    n36843, n36844, n36845, n36846, n36847, n36848,
    n36849, n36850, n36851, n36852, n36853, n36854,
    n36855, n36856, n36857, n36858, n36859, n36860,
    n36861, n36862, n36863, n36864, n36865, n36866,
    n36867, n36868, n36869, n36870, n36871, n36872,
    n36873, n36874, n36875, n36876, n36877, n36878,
    n36879, n36880, n36881, n36882, n36883, n36884,
    n36885, n36886, n36887, n36888, n36889, n36890,
    n36891, n36892, n36893, n36894, n36895, n36896,
    n36897, n36898, n36899, n36900, n36901, n36902,
    n36903, n36904, n36905, n36906, n36907, n36908,
    n36909, n36910, n36911, n36912, n36913, n36914,
    n36915, n36916, n36917, n36918, n36919, n36920,
    n36921, n36922, n36923, n36924, n36925, n36926,
    n36927, n36928, n36929, n36930, n36931, n36932,
    n36933, n36934, n36935, n36936, n36937, n36938,
    n36939, n36940, n36941, n36942, n36943, n36944,
    n36945, n36946, n36947, n36948, n36949, n36950,
    n36951, n36952, n36953, n36954, n36955, n36956,
    n36957, n36958, n36959, n36960, n36961, n36962,
    n36963, n36964, n36965, n36966, n36967, n36968,
    n36969, n36970, n36971, n36972, n36973, n36974,
    n36975, n36976, n36977, n36978, n36979, n36980,
    n36981, n36982, n36983, n36984, n36985, n36986,
    n36987, n36988, n36989, n36990, n36991, n36992,
    n36993, n36994, n36995, n36996, n36997, n36998,
    n36999, n37000, n37001, n37002, n37003, n37004,
    n37005, n37006, n37007, n37008, n37009, n37010,
    n37011, n37012, n37013, n37014, n37015, n37016,
    n37017, n37018, n37019, n37020, n37021, n37022,
    n37023, n37024, n37025, n37026, n37027, n37028,
    n37029, n37030, n37031, n37032, n37033, n37034,
    n37035, n37036, n37037, n37038, n37039, n37040,
    n37041, n37042, n37043, n37044, n37045, n37046,
    n37047, n37048, n37049, n37050, n37051, n37052,
    n37053, n37054, n37055, n37056, n37057, n37058,
    n37059, n37060, n37061, n37062, n37063, n37064,
    n37065, n37066, n37067, n37068, n37069, n37070,
    n37071, n37072, n37073, n37074, n37075, n37076,
    n37077, n37078, n37079, n37080, n37081, n37082,
    n37083, n37084, n37085, n37086, n37087, n37088,
    n37089, n37090, n37091, n37092, n37093, n37094,
    n37095, n37096, n37097, n37098, n37099, n37100,
    n37101, n37102, n37103, n37104, n37105, n37106,
    n37107, n37108, n37109, n37110, n37111, n37112,
    n37113, n37114, n37115, n37116, n37117, n37118,
    n37119, n37120, n37121, n37122, n37123, n37124,
    n37125, n37126, n37127, n37128, n37129, n37130,
    n37131, n37132, n37133, n37134, n37135, n37136,
    n37137, n37138, n37139, n37140, n37141, n37142,
    n37143, n37144, n37145, n37146, n37147, n37148,
    n37149, n37150, n37151, n37152, n37153, n37154,
    n37155, n37156, n37157, n37158, n37159, n37160,
    n37161, n37162, n37163, n37164, n37165, n37166,
    n37167, n37168, n37169, n37170, n37171, n37172,
    n37173, n37174, n37175, n37176, n37177, n37178,
    n37179, n37180, n37181, n37182, n37183, n37184,
    n37185, n37186, n37187, n37188, n37189, n37190,
    n37191, n37192, n37193, n37195, n37196, n37197,
    n37198, n37199, n37200, n37201, n37202, n37203,
    n37204, n37205, n37206, n37207, n37208, n37209,
    n37210, n37211, n37212, n37213, n37214, n37215,
    n37216, n37217, n37218, n37219, n37220, n37221,
    n37222, n37223, n37224, n37225, n37226, n37227,
    n37228, n37229, n37230, n37231, n37232, n37233,
    n37234, n37235, n37236, n37237, n37238, n37239,
    n37240, n37241, n37242, n37243, n37244, n37245,
    n37246, n37247, n37248, n37249, n37250, n37251,
    n37252, n37253, n37254, n37255, n37256, n37257,
    n37258, n37259, n37260, n37261, n37262, n37263,
    n37264, n37265, n37266, n37267, n37268, n37269,
    n37270, n37271, n37272, n37273, n37274, n37275,
    n37276, n37277, n37278, n37279, n37280, n37281,
    n37282, n37283, n37284, n37285, n37286, n37287,
    n37288, n37289, n37290, n37291, n37292, n37293,
    n37294, n37295, n37296, n37297, n37298, n37299,
    n37300, n37301, n37302, n37303, n37304, n37305,
    n37306, n37307, n37308, n37309, n37310, n37311,
    n37312, n37313, n37314, n37315, n37316, n37317,
    n37318, n37319, n37320, n37321, n37322, n37323,
    n37324, n37325, n37326, n37327, n37328, n37329,
    n37330, n37331, n37332, n37333, n37334, n37335,
    n37336, n37337, n37338, n37339, n37340, n37341,
    n37342, n37343, n37344, n37345, n37346, n37347,
    n37348, n37349, n37350, n37351, n37352, n37353,
    n37354, n37355, n37356, n37357, n37358, n37359,
    n37360, n37361, n37362, n37363, n37364, n37365,
    n37366, n37367, n37368, n37369, n37370, n37371,
    n37372, n37373, n37374, n37375, n37376, n37377,
    n37378, n37379, n37380, n37381, n37382, n37383,
    n37384, n37385, n37386, n37387, n37388, n37389,
    n37390, n37391, n37392, n37393, n37394, n37395,
    n37396, n37397, n37398, n37399, n37400, n37401,
    n37402, n37403, n37404, n37405, n37406, n37407,
    n37408, n37409, n37410, n37411, n37412, n37413,
    n37414, n37415, n37416, n37417, n37418, n37419,
    n37420, n37421, n37422, n37423, n37424, n37425,
    n37426, n37427, n37428, n37429, n37430, n37431,
    n37432, n37433, n37434, n37435, n37436, n37437,
    n37438, n37439, n37440, n37441, n37442, n37443,
    n37444, n37445, n37446, n37447, n37448, n37449,
    n37450, n37451, n37452, n37453, n37454, n37455,
    n37456, n37457, n37458, n37459, n37460, n37461,
    n37462, n37463, n37464, n37465, n37466, n37467,
    n37468, n37469, n37470, n37471, n37472, n37473,
    n37474, n37475, n37476, n37477, n37478, n37479,
    n37480, n37481, n37482, n37483, n37484, n37485,
    n37486, n37487, n37488, n37489, n37490, n37491,
    n37492, n37493, n37494, n37495, n37496, n37497,
    n37498, n37499, n37500, n37501, n37502, n37503,
    n37504, n37505, n37506, n37507, n37508, n37509,
    n37510, n37511, n37512, n37513, n37514, n37515,
    n37516, n37517, n37518, n37519, n37520, n37521,
    n37522, n37523, n37524, n37525, n37526, n37527,
    n37528, n37529, n37530, n37531, n37532, n37533,
    n37534, n37535, n37536, n37537, n37538, n37539,
    n37540, n37541, n37542, n37543, n37544, n37545,
    n37546, n37547, n37548, n37549, n37550, n37551,
    n37552, n37553, n37554, n37555, n37556, n37557,
    n37558, n37559, n37560, n37561, n37562, n37563,
    n37564, n37565, n37566, n37567, n37568, n37569,
    n37570, n37571, n37572, n37573, n37574, n37575,
    n37576, n37577, n37578, n37579, n37580, n37581,
    n37582, n37583, n37584, n37585, n37586, n37587,
    n37588, n37589, n37590, n37591, n37592, n37593,
    n37594, n37595, n37596, n37597, n37598, n37599,
    n37600, n37601, n37602, n37603, n37604, n37605,
    n37606, n37607, n37608, n37609, n37610, n37611,
    n37612, n37613, n37614, n37615, n37616, n37617,
    n37618, n37619, n37620, n37621, n37622, n37623,
    n37624, n37625, n37626, n37627, n37628, n37629,
    n37630, n37631, n37632, n37633, n37634, n37635,
    n37636, n37637, n37638, n37639, n37640, n37641,
    n37642, n37643, n37644, n37645, n37646, n37647,
    n37648, n37649, n37650, n37651, n37652, n37653,
    n37654, n37655, n37656, n37657, n37658, n37659,
    n37660, n37661, n37662, n37663, n37664, n37665,
    n37666, n37667, n37668, n37669, n37670, n37671,
    n37672, n37673, n37674, n37675, n37676, n37677,
    n37678, n37679, n37680, n37681, n37682, n37683,
    n37684, n37685, n37686, n37687, n37688, n37689,
    n37690, n37691, n37692, n37693, n37694, n37695,
    n37696, n37697, n37698, n37699, n37700, n37701,
    n37702, n37703, n37704, n37705, n37706, n37707,
    n37708, n37709, n37710, n37711, n37712, n37713,
    n37714, n37715, n37716, n37717, n37718, n37719,
    n37720, n37721, n37722, n37723, n37724, n37725,
    n37726, n37727, n37728, n37729, n37730, n37731,
    n37732, n37733, n37734, n37735, n37736, n37737,
    n37738, n37739, n37740, n37741, n37742, n37743,
    n37744, n37745, n37746, n37747, n37748, n37749,
    n37750, n37751, n37752, n37753, n37754, n37755,
    n37756, n37757, n37758, n37759, n37760, n37761,
    n37762, n37763, n37764, n37765, n37766, n37767,
    n37768, n37770, n37771, n37772, n37773, n37774,
    n37775, n37776, n37777, n37778, n37779, n37780,
    n37781, n37782, n37783, n37784, n37785, n37786,
    n37787, n37788, n37789, n37790, n37791, n37792,
    n37793, n37794, n37795, n37796, n37797, n37798,
    n37799, n37800, n37801, n37802, n37803, n37804,
    n37805, n37806, n37807, n37808, n37809, n37810,
    n37811, n37812, n37813, n37814, n37815, n37816,
    n37817, n37818, n37819, n37820, n37821, n37822,
    n37823, n37824, n37825, n37826, n37827, n37828,
    n37829, n37830, n37831, n37832, n37833, n37834,
    n37835, n37836, n37837, n37838, n37839, n37840,
    n37841, n37842, n37843, n37844, n37845, n37846,
    n37847, n37848, n37849, n37850, n37851, n37852,
    n37853, n37854, n37855, n37856, n37857, n37858,
    n37859, n37860, n37861, n37862, n37863, n37864,
    n37865, n37866, n37867, n37868, n37869, n37870,
    n37871, n37872, n37873, n37874, n37875, n37876,
    n37877, n37878, n37879, n37880, n37881, n37882,
    n37883, n37884, n37885, n37886, n37887, n37888,
    n37889, n37890, n37891, n37892, n37893, n37895,
    n37896, n37897, n37898, n37899, n37900, n37901,
    n37902, n37903, n37904, n37905, n37906, n37907,
    n37908, n37909, n37910, n37911, n37912, n37913,
    n37914, n37915, n37916, n37917, n37918, n37919,
    n37920, n37921, n37922, n37923, n37924, n37925,
    n37926, n37927, n37928, n37929, n37930, n37931,
    n37932, n37933, n37934, n37935, n37936, n37937,
    n37938, n37939, n37940, n37941, n37942, n37943,
    n37944, n37945, n37946, n37948, n37949, n37950,
    n37951, n37952, n37953, n37954, n37955, n37956,
    n37957, n37958, n37959, n37960, n37961, n37962,
    n37963, n37964, n37965, n37966, n37967, n37968,
    n37969, n37970, n37971, n37972, n37973, n37974,
    n37975, n37976, n37977, n37979, n37980, n37981,
    n37982, n37983, n37984, n37985, n37986, n37987,
    n37988, n37989, n37991, n37992, n37993, n37994,
    n37995, n37996, n37997, n37998, n37999, n38000,
    n38001, n38002, n38003, n38004, n38005, n38006,
    n38007, n38008, n38009, n38010, n38011, n38012,
    n38013, n38014, n38015, n38016, n38017, n38018,
    n38019, n38020, n38021, n38022, n38023, n38024,
    n38025, n38026, n38027, n38028, n38029, n38030,
    n38031, n38032, n38033, n38034, n38035, n38036,
    n38037, n38038, n38039, n38040, n38041, n38042,
    n38043, n38044, n38045, n38046, n38047, n38048,
    n38049, n38050, n38051, n38052, n38053, n38054,
    n38055, n38056, n38057, n38058, n38059, n38060,
    n38061, n38062, n38063, n38064, n38065, n38066,
    n38067, n38068, n38069, n38070, n38071, n38072,
    n38074, n38075, n38076, n38077, n38078, n38079,
    n38080, n38081, n38082, n38083, n38084, n38085,
    n38086, n38087, n38088, n38089, n38090, n38091,
    n38092, n38093, n38094, n38095, n38096, n38097,
    n38098, n38099, n38100, n38101, n38102, n38103,
    n38104, n38105, n38106, n38107, n38108, n38109,
    n38111, n38112, n38113, n38114, n38115, n38116,
    n38117, n38118, n38119, n38120, n38121, n38122,
    n38123, n38124, n38125, n38126, n38127, n38128,
    n38129, n38130, n38131, n38132, n38134, n38135,
    n38136, n38137, n38138, n38139, n38140, n38141,
    n38142, n38143, n38144, n38145, n38146, n38147,
    n38148, n38149, n38150, n38151, n38152, n38153,
    n38154, n38155, n38156, n38157, n38158, n38159,
    n38160, n38161, n38162, n38163, n38164, n38165,
    n38166, n38167, n38168, n38169, n38170, n38171,
    n38172, n38173, n38174, n38175, n38176, n38177,
    n38178, n38179, n38180, n38181, n38182, n38183,
    n38184, n38185, n38186, n38187, n38188, n38189,
    n38190, n38191, n38192, n38193, n38194, n38195,
    n38196, n38197, n38198, n38199, n38200, n38201,
    n38202, n38203, n38204, n38205, n38206, n38207,
    n38208, n38209, n38210, n38211, n38212, n38213,
    n38214, n38215, n38216, n38217, n38218, n38219,
    n38220, n38221, n38222, n38223, n38224, n38225,
    n38226, n38227, n38228, n38229, n38230, n38231,
    n38232, n38233, n38234, n38235, n38236, n38237,
    n38238, n38239, n38240, n38241, n38242, n38243,
    n38244, n38245, n38246, n38247, n38248, n38249,
    n38250, n38251, n38252, n38253, n38254, n38255,
    n38256, n38257, n38258, n38259, n38260, n38261,
    n38262, n38263, n38264, n38265, n38266, n38267,
    n38268, n38269, n38270, n38271, n38272, n38273,
    n38274, n38275, n38276, n38277, n38278, n38279,
    n38280, n38281, n38282, n38283, n38284, n38285,
    n38286, n38287, n38288, n38289, n38290, n38291,
    n38292, n38293, n38294, n38295, n38296, n38297,
    n38298, n38299, n38300, n38301, n38302, n38303,
    n38304, n38305, n38306, n38307, n38308, n38309,
    n38310, n38311, n38312, n38313, n38314, n38315,
    n38316, n38317, n38318, n38319, n38320, n38321,
    n38322, n38323, n38324, n38325, n38326, n38327,
    n38328, n38329, n38330, n38331, n38332, n38333,
    n38334, n38335, n38336, n38337, n38338, n38339,
    n38340, n38341, n38342, n38343, n38344, n38345,
    n38346, n38347, n38348, n38349, n38350, n38351,
    n38352, n38353, n38354, n38355, n38356, n38357,
    n38358, n38359, n38360, n38361, n38362, n38363,
    n38364, n38365, n38366, n38367, n38368, n38369,
    n38370, n38371, n38372, n38373, n38374, n38375,
    n38376, n38377, n38378, n38379, n38380, n38381,
    n38382, n38383, n38384, n38385, n38386, n38387,
    n38388, n38389, n38390, n38391, n38392, n38393,
    n38394, n38395, n38396, n38397, n38398, n38399,
    n38400, n38401, n38402, n38403, n38404, n38405,
    n38406, n38407, n38408, n38409, n38410, n38411,
    n38412, n38413, n38414, n38415, n38416, n38417,
    n38418, n38419, n38420, n38421, n38422, n38423,
    n38424, n38425, n38426, n38427, n38428, n38429,
    n38430, n38431, n38432, n38433, n38434, n38435,
    n38436, n38437, n38438, n38439, n38440, n38441,
    n38442, n38443, n38444, n38445, n38446, n38447,
    n38448, n38449, n38450, n38451, n38452, n38453,
    n38454, n38455, n38456, n38457, n38458, n38459,
    n38460, n38461, n38462, n38463, n38464, n38465,
    n38466, n38467, n38468, n38469, n38470, n38471,
    n38472, n38473, n38474, n38475, n38476, n38477,
    n38478, n38479, n38480, n38481, n38482, n38483,
    n38484, n38485, n38486, n38487, n38488, n38489,
    n38490, n38491, n38492, n38493, n38494, n38495,
    n38496, n38497, n38498, n38500, n38501, n38502,
    n38503, n38504, n38505, n38506, n38507, n38508,
    n38509, n38510, n38511, n38512, n38513, n38514,
    n38515, n38516, n38517, n38518, n38519, n38520,
    n38521, n38522, n38523, n38524, n38525, n38526,
    n38527, n38528, n38529, n38530, n38531, n38532,
    n38533, n38534, n38535, n38536, n38537, n38538,
    n38539, n38540, n38541, n38542, n38543, n38544,
    n38545, n38546, n38547, n38548, n38549, n38550,
    n38551, n38552, n38553, n38554, n38555, n38556,
    n38557, n38558, n38559, n38560, n38561, n38562,
    n38563, n38564, n38565, n38566, n38567, n38568,
    n38569, n38570, n38571, n38572, n38573, n38574,
    n38575, n38576, n38577, n38578, n38579, n38580,
    n38581, n38582, n38583, n38584, n38585, n38586,
    n38587, n38588, n38589, n38590, n38591, n38592,
    n38593, n38594, n38595, n38596, n38597, n38598,
    n38599, n38600, n38601, n38602, n38603, n38604,
    n38605, n38606, n38607, n38608, n38609, n38610,
    n38611, n38612, n38613, n38614, n38615, n38616,
    n38617, n38618, n38619, n38620, n38621, n38622,
    n38623, n38624, n38625, n38626, n38627, n38628,
    n38629, n38630, n38631, n38632, n38633, n38634,
    n38635, n38636, n38637, n38638, n38639, n38640,
    n38641, n38642, n38643, n38644, n38645, n38646,
    n38647, n38648, n38649, n38650, n38651, n38652,
    n38653, n38654, n38655, n38656, n38657, n38658,
    n38659, n38660, n38661, n38662, n38663, n38664,
    n38665, n38666, n38667, n38668, n38669, n38670,
    n38671, n38672, n38673, n38674, n38675, n38676,
    n38677, n38678, n38679, n38680, n38681, n38682,
    n38683, n38684, n38685, n38686, n38687, n38688,
    n38689, n38690, n38691, n38692, n38693, n38694,
    n38695, n38696, n38697, n38698, n38699, n38700,
    n38701, n38702, n38703, n38704, n38705, n38706,
    n38707, n38708, n38709, n38710, n38711, n38712,
    n38713, n38714, n38715, n38716, n38717, n38718,
    n38719, n38720, n38721, n38722, n38723, n38724,
    n38725, n38726, n38727, n38728, n38729, n38730,
    n38731, n38732, n38733, n38734, n38735, n38736,
    n38737, n38738, n38739, n38740, n38741, n38742,
    n38743, n38744, n38745, n38746, n38747, n38748,
    n38749, n38750, n38751, n38752, n38753, n38754,
    n38755, n38756, n38757, n38758, n38759, n38760,
    n38761, n38762, n38763, n38764, n38765, n38766,
    n38767, n38768, n38769, n38770, n38771, n38772,
    n38773, n38774, n38775, n38776, n38777, n38778,
    n38779, n38781, n38782, n38783, n38784, n38785,
    n38786, n38787, n38788, n38789, n38790, n38791,
    n38792, n38793, n38794, n38795, n38796, n38797,
    n38798, n38799, n38800, n38801, n38802, n38803,
    n38804, n38805, n38806, n38807, n38808, n38809,
    n38810, n38811, n38812, n38813, n38814, n38815,
    n38816, n38817, n38818, n38819, n38820, n38821,
    n38822, n38823, n38824, n38825, n38826, n38827,
    n38828, n38829, n38830, n38831, n38832, n38833,
    n38834, n38835, n38836, n38837, n38838, n38839,
    n38840, n38841, n38842, n38843, n38844, n38845,
    n38846, n38847, n38848, n38849, n38850, n38851,
    n38852, n38853, n38854, n38855, n38856, n38857,
    n38858, n38859, n38860, n38861, n38862, n38863,
    n38864, n38865, n38866, n38867, n38868, n38869,
    n38870, n38871, n38872, n38873, n38874, n38875,
    n38876, n38877, n38878, n38879, n38880, n38881,
    n38882, n38883, n38884, n38885, n38886, n38887,
    n38888, n38889, n38890, n38891, n38892, n38893,
    n38894, n38895, n38896, n38897, n38898, n38899,
    n38900, n38901, n38902, n38903, n38904, n38905,
    n38906, n38907, n38908, n38909, n38910, n38911,
    n38912, n38913, n38914, n38915, n38916, n38917,
    n38918, n38919, n38920, n38921, n38922, n38923,
    n38924, n38925, n38926, n38927, n38928, n38929,
    n38930, n38931, n38932, n38933, n38934, n38935,
    n38936, n38937, n38938, n38939, n38940, n38941,
    n38942, n38943, n38944, n38945, n38946, n38947,
    n38948, n38949, n38950, n38951, n38952, n38953,
    n38954, n38955, n38956, n38957, n38958, n38959,
    n38960, n38961, n38962, n38963, n38964, n38965,
    n38966, n38967, n38968, n38969, n38970, n38971,
    n38972, n38973, n38974, n38975, n38976, n38977,
    n38978, n38979, n38981, n38982, n38983, n38984,
    n38985, n38986, n38987, n38988, n38989, n38990,
    n38991, n38992, n38994, n38995, n38996, n38997,
    n38998, n38999, n39000, n39001, n39002, n39003,
    n39004, n39005, n39006, n39007, n39008, n39009,
    n39010, n39011, n39012, n39013, n39014, n39015,
    n39016, n39017, n39018, n39019, n39020, n39021,
    n39022, n39023, n39024, n39025, n39026, n39027,
    n39028, n39029, n39030, n39031, n39032, n39033,
    n39034, n39035, n39036, n39037, n39038, n39039,
    n39040, n39041, n39042, n39043, n39044, n39045,
    n39046, n39047, n39048, n39049, n39050, n39051,
    n39052, n39053, n39054, n39055, n39056, n39057,
    n39058, n39059, n39060, n39061, n39062, n39063,
    n39064, n39065, n39066, n39067, n39068, n39069,
    n39070, n39071, n39072, n39073, n39074, n39075,
    n39076, n39077, n39078, n39079, n39080, n39081,
    n39082, n39083, n39084, n39085, n39086, n39087,
    n39088, n39089, n39090, n39091, n39092, n39093,
    n39094, n39095, n39096, n39097, n39098, n39099,
    n39100, n39101, n39102, n39103, n39104, n39105,
    n39106, n39107, n39108, n39109, n39110, n39111,
    n39112, n39113, n39114, n39115, n39116, n39117,
    n39118, n39119, n39120, n39121, n39122, n39123,
    n39124, n39125, n39126, n39127, n39128, n39129,
    n39130, n39131, n39132, n39133, n39134, n39135,
    n39136, n39137, n39138, n39139, n39140, n39141,
    n39142, n39143, n39144, n39145, n39146, n39147,
    n39148, n39149, n39150, n39151, n39152, n39153,
    n39154, n39155, n39156, n39157, n39158, n39159,
    n39160, n39161, n39162, n39163, n39164, n39165,
    n39166, n39167, n39168, n39169, n39170, n39171,
    n39172, n39173, n39174, n39175, n39176, n39177,
    n39178, n39179, n39180, n39181, n39182, n39183,
    n39184, n39185, n39186, n39187, n39188, n39189,
    n39190, n39191, n39192, n39193, n39194, n39195,
    n39196, n39197, n39198, n39199, n39200, n39201,
    n39202, n39203, n39204, n39205, n39206, n39207,
    n39208, n39209, n39210, n39211, n39212, n39213,
    n39214, n39215, n39216, n39217, n39218, n39219,
    n39220, n39221, n39222, n39223, n39224, n39225,
    n39226, n39227, n39228, n39229, n39230, n39231,
    n39232, n39233, n39234, n39235, n39236, n39237,
    n39239, n39240, n39241, n39242, n39243, n39244,
    n39245, n39246, n39247, n39248, n39249, n39250,
    n39251, n39252, n39253, n39254, n39255, n39256,
    n39257, n39258, n39259, n39260, n39261, n39262,
    n39263, n39264, n39265, n39266, n39267, n39268,
    n39269, n39270, n39271, n39272, n39273, n39274,
    n39275, n39276, n39277, n39278, n39279, n39280,
    n39281, n39282, n39283, n39284, n39285, n39286,
    n39287, n39288, n39289, n39290, n39291, n39292,
    n39293, n39294, n39295, n39296, n39297, n39298,
    n39299, n39300, n39301, n39302, n39303, n39304,
    n39305, n39306, n39307, n39308, n39309, n39310,
    n39311, n39312, n39313, n39314, n39315, n39316,
    n39317, n39318, n39319, n39320, n39321, n39322,
    n39323, n39324, n39325, n39326, n39327, n39328,
    n39329, n39330, n39331, n39332, n39333, n39334,
    n39335, n39336, n39337, n39338, n39339, n39340,
    n39341, n39342, n39343, n39344, n39345, n39346,
    n39347, n39348, n39349, n39350, n39351, n39352,
    n39353, n39354, n39355, n39356, n39357, n39358,
    n39359, n39360, n39361, n39362, n39363, n39364,
    n39365, n39366, n39367, n39368, n39369, n39370,
    n39371, n39372, n39373, n39374, n39375, n39376,
    n39377, n39378, n39379, n39380, n39381, n39382,
    n39383, n39384, n39385, n39386, n39387, n39388,
    n39389, n39390, n39391, n39392, n39393, n39394,
    n39395, n39396, n39397, n39398, n39399, n39400,
    n39401, n39402, n39403, n39404, n39405, n39406,
    n39407, n39408, n39409, n39410, n39411, n39412,
    n39413, n39414, n39415, n39416, n39417, n39418,
    n39419, n39420, n39421, n39422, n39423, n39424,
    n39425, n39426, n39427, n39428, n39429, n39430,
    n39431, n39432, n39433, n39434, n39435, n39436,
    n39437, n39438, n39439, n39440, n39441, n39442,
    n39443, n39444, n39445, n39446, n39447, n39448,
    n39449, n39450, n39451, n39452, n39453, n39454,
    n39455, n39456, n39457, n39458, n39459, n39460,
    n39461, n39462, n39463, n39464, n39465, n39466,
    n39467, n39468, n39469, n39470, n39471, n39472,
    n39473, n39474, n39475, n39476, n39477, n39478,
    n39479, n39480, n39481, n39482, n39483, n39484,
    n39485, n39486, n39487, n39488, n39489, n39490,
    n39491, n39492, n39493, n39494, n39495, n39496,
    n39497, n39498, n39499, n39500, n39501, n39502,
    n39503, n39504, n39505, n39506, n39507, n39508,
    n39509, n39510, n39511, n39512, n39513, n39514,
    n39515, n39516, n39517, n39518, n39519, n39520,
    n39521, n39522, n39523, n39524, n39525, n39526,
    n39527, n39528, n39529, n39530, n39531, n39532,
    n39533, n39534, n39535, n39536, n39537, n39538,
    n39539, n39540, n39541, n39542, n39543, n39544,
    n39546, n39547, n39548, n39549, n39550, n39551,
    n39552, n39553, n39554, n39555, n39556, n39557,
    n39558, n39559, n39560, n39561, n39562, n39563,
    n39564, n39565, n39566, n39567, n39568, n39569,
    n39570, n39571, n39572, n39573, n39574, n39575,
    n39576, n39577, n39578, n39579, n39580, n39581,
    n39582, n39583, n39584, n39585, n39586, n39587,
    n39588, n39589, n39590, n39591, n39592, n39593,
    n39594, n39595, n39596, n39597, n39598, n39599,
    n39600, n39601, n39602, n39603, n39604, n39605,
    n39606, n39607, n39608, n39609, n39610, n39611,
    n39612, n39613, n39614, n39615, n39616, n39617,
    n39618, n39619, n39620, n39621, n39622, n39623,
    n39624, n39625, n39626, n39627, n39628, n39629,
    n39630, n39631, n39632, n39634, n39635, n39636,
    n39637, n39638, n39639, n39640, n39641, n39642,
    n39643, n39644, n39645, n39646, n39647, n39648,
    n39649, n39650, n39651, n39652, n39653, n39654,
    n39655, n39656, n39657, n39658, n39659, n39660,
    n39661, n39662, n39663, n39664, n39665, n39666,
    n39667, n39668, n39669, n39670, n39671, n39672,
    n39673, n39674, n39675, n39676, n39677, n39678,
    n39679, n39680, n39681, n39682, n39683, n39684,
    n39685, n39686, n39687, n39688, n39689, n39690,
    n39691, n39692, n39693, n39694, n39695, n39696,
    n39697, n39698, n39699, n39700, n39701, n39702,
    n39703, n39704, n39705, n39706, n39707, n39708,
    n39709, n39710, n39711, n39712, n39713, n39714,
    n39715, n39716, n39717, n39718, n39719, n39720,
    n39721, n39722, n39723, n39724, n39725, n39726,
    n39727, n39728, n39729, n39730, n39731, n39732,
    n39733, n39734, n39735, n39736, n39737, n39738,
    n39739, n39740, n39741, n39742, n39743, n39744,
    n39745, n39746, n39747, n39748, n39749, n39750,
    n39751, n39752, n39753, n39754, n39755, n39756,
    n39757, n39758, n39759, n39760, n39761, n39762,
    n39763, n39764, n39765, n39766, n39767, n39768,
    n39769, n39770, n39771, n39772, n39773, n39774,
    n39775, n39776, n39777, n39778, n39779, n39780,
    n39781, n39782, n39783, n39784, n39785, n39786,
    n39787, n39788, n39789, n39790, n39791, n39792,
    n39793, n39794, n39795, n39796, n39797, n39798,
    n39799, n39800, n39801, n39802, n39803, n39804,
    n39805, n39806, n39807, n39808, n39809, n39810,
    n39811, n39812, n39813, n39814, n39815, n39816,
    n39817, n39818, n39819, n39820, n39821, n39822,
    n39823, n39824, n39825, n39826, n39827, n39828,
    n39829, n39830, n39831, n39832, n39833, n39834,
    n39835, n39836, n39837, n39838, n39839, n39840,
    n39841, n39842, n39843, n39844, n39845, n39846,
    n39847, n39848, n39849, n39850, n39851, n39852,
    n39853, n39854, n39855, n39856, n39857, n39858,
    n39859, n39860, n39861, n39862, n39863, n39864,
    n39865, n39866, n39867, n39868, n39869, n39870,
    n39871, n39872, n39873, n39874, n39875, n39876,
    n39877, n39878, n39879, n39880, n39881, n39882,
    n39883, n39884, n39885, n39886, n39887, n39888,
    n39889, n39890, n39891, n39892, n39893, n39894,
    n39895, n39896, n39897, n39898, n39899, n39900,
    n39901, n39902, n39903, n39904, n39905, n39906,
    n39907, n39908, n39909, n39910, n39911, n39912,
    n39913, n39914, n39915, n39916, n39917, n39918,
    n39919, n39920, n39921, n39922, n39923, n39924,
    n39925, n39926, n39927, n39928, n39929, n39930,
    n39931, n39932, n39933, n39934, n39935, n39936,
    n39937, n39938, n39939, n39940, n39941, n39942,
    n39943, n39944, n39945, n39946, n39947, n39948,
    n39949, n39950, n39951, n39952, n39953, n39954,
    n39955, n39956, n39957, n39958, n39959, n39960,
    n39961, n39962, n39963, n39964, n39965, n39966,
    n39967, n39968, n39969, n39970, n39971, n39972,
    n39973, n39974, n39975, n39976, n39977, n39978,
    n39979, n39980, n39981, n39982, n39983, n39984,
    n39985, n39986, n39987, n39988, n39989, n39990,
    n39991, n39992, n39993, n39994, n39995, n39996,
    n39997, n39998, n39999, n40000, n40001, n40002,
    n40003, n40004, n40005, n40006, n40007, n40008,
    n40009, n40010, n40011, n40012, n40013, n40014,
    n40015, n40016, n40017, n40018, n40020, n40021,
    n40022, n40023, n40024, n40025, n40026, n40027,
    n40028, n40029, n40030, n40031, n40032, n40033,
    n40034, n40035, n40036, n40037, n40038, n40039,
    n40040, n40041, n40042, n40043, n40044, n40045,
    n40046, n40047, n40048, n40049, n40050, n40051,
    n40052, n40053, n40054, n40055, n40056, n40057,
    n40058, n40059, n40060, n40061, n40062, n40063,
    n40064, n40065, n40066, n40067, n40068, n40069,
    n40070, n40071, n40072, n40073, n40074, n40075,
    n40076, n40077, n40078, n40079, n40080, n40081,
    n40082, n40083, n40084, n40085, n40086, n40087,
    n40088, n40089, n40090, n40091, n40092, n40093,
    n40094, n40095, n40096, n40097, n40098, n40099,
    n40100, n40101, n40102, n40103, n40104, n40105,
    n40106, n40107, n40108, n40109, n40110, n40111,
    n40112, n40113, n40114, n40115, n40116, n40117,
    n40118, n40119, n40120, n40121, n40122, n40123,
    n40124, n40125, n40126, n40127, n40128, n40129,
    n40130, n40131, n40132, n40133, n40134, n40135,
    n40136, n40137, n40138, n40139, n40140, n40141,
    n40142, n40143, n40144, n40145, n40146, n40147,
    n40148, n40149, n40150, n40151, n40152, n40153,
    n40154, n40155, n40156, n40157, n40158, n40159,
    n40160, n40161, n40162, n40163, n40164, n40165,
    n40166, n40167, n40168, n40169, n40170, n40171,
    n40172, n40173, n40174, n40175, n40176, n40177,
    n40178, n40179, n40180, n40181, n40182, n40183,
    n40184, n40185, n40186, n40187, n40188, n40189,
    n40190, n40191, n40192, n40193, n40194, n40195,
    n40196, n40197, n40198, n40199, n40200, n40201,
    n40202, n40203, n40204, n40205, n40206, n40207,
    n40208, n40209, n40210, n40211, n40212, n40213,
    n40214, n40215, n40216, n40217, n40218, n40219,
    n40220, n40221, n40222, n40223, n40224, n40225,
    n40226, n40227, n40228, n40229, n40230, n40231,
    n40232, n40233, n40234, n40235, n40236, n40237,
    n40238, n40239, n40240, n40241, n40242, n40243,
    n40244, n40245, n40246, n40247, n40248, n40249,
    n40250, n40251, n40252, n40253, n40254, n40255,
    n40256, n40257, n40258, n40259, n40260, n40261,
    n40262, n40263, n40264, n40265, n40266, n40267,
    n40268, n40269, n40270, n40271, n40272, n40273,
    n40274, n40275, n40276, n40278, n40279, n40280,
    n40281, n40282, n40283, n40284, n40285, n40286,
    n40287, n40288, n40289, n40290, n40291, n40292,
    n40293, n40294, n40295, n40296, n40297, n40298,
    n40299, n40300, n40301, n40302, n40303, n40304,
    n40305, n40306, n40307, n40308, n40309, n40310,
    n40311, n40312, n40313, n40314, n40315, n40316,
    n40317, n40318, n40319, n40320, n40321, n40322,
    n40323, n40324, n40325, n40326, n40327, n40328,
    n40329, n40330, n40331, n40332, n40333, n40334,
    n40335, n40336, n40337, n40338, n40339, n40340,
    n40341, n40342, n40343, n40344, n40345, n40346,
    n40347, n40348, n40349, n40350, n40351, n40352,
    n40353, n40354, n40355, n40356, n40358, n40359,
    n40360, n40361, n40362, n40363, n40364, n40365,
    n40366, n40367, n40368, n40369, n40370, n40371,
    n40372, n40373, n40374, n40375, n40376, n40377,
    n40378, n40379, n40380, n40381, n40382, n40383,
    n40384, n40385, n40386, n40387, n40388, n40389,
    n40390, n40391, n40392, n40393, n40394, n40395,
    n40396, n40397, n40398, n40399, n40400, n40401,
    n40402, n40403, n40404, n40405, n40406, n40407,
    n40408, n40409, n40410, n40411, n40412, n40413,
    n40414, n40415, n40416, n40417, n40418, n40419,
    n40420, n40421, n40422, n40423, n40424, n40425,
    n40426, n40427, n40428, n40429, n40430, n40431,
    n40432, n40433, n40434, n40435, n40436, n40437,
    n40438, n40439, n40440, n40441, n40442, n40443,
    n40444, n40445, n40446, n40447, n40448, n40449,
    n40450, n40451, n40452, n40453, n40454, n40455,
    n40456, n40457, n40458, n40459, n40460, n40461,
    n40462, n40463, n40464, n40465, n40466, n40467,
    n40468, n40469, n40470, n40471, n40472, n40473,
    n40474, n40475, n40476, n40477, n40478, n40479,
    n40480, n40481, n40482, n40483, n40484, n40485,
    n40486, n40487, n40488, n40489, n40490, n40491,
    n40492, n40493, n40494, n40495, n40496, n40497,
    n40498, n40499, n40500, n40501, n40502, n40503,
    n40504, n40505, n40506, n40507, n40508, n40509,
    n40510, n40511, n40512, n40513, n40514, n40515,
    n40516, n40517, n40518, n40519, n40520, n40521,
    n40522, n40523, n40524, n40525, n40526, n40527,
    n40528, n40529, n40530, n40531, n40532, n40533,
    n40534, n40535, n40536, n40537, n40538, n40539,
    n40540, n40541, n40542, n40543, n40544, n40545,
    n40546, n40547, n40548, n40549, n40550, n40551,
    n40552, n40553, n40554, n40555, n40556, n40557,
    n40558, n40559, n40560, n40561, n40562, n40563,
    n40564, n40565, n40566, n40567, n40568, n40569,
    n40570, n40571, n40572, n40573, n40574, n40575,
    n40576, n40577, n40578, n40579, n40580, n40581,
    n40582, n40583, n40584, n40585, n40586, n40587,
    n40588, n40589, n40590, n40591, n40592, n40593,
    n40594, n40595, n40596, n40597, n40598, n40599,
    n40600, n40601, n40602, n40603, n40604, n40605,
    n40606, n40607, n40608, n40609, n40610, n40611,
    n40612, n40613, n40614, n40615, n40616, n40617,
    n40618, n40619, n40620, n40621, n40622, n40623,
    n40624, n40625, n40626, n40627, n40628, n40629,
    n40630, n40631, n40632, n40633, n40634, n40635,
    n40636, n40637, n40638, n40639, n40640, n40641,
    n40642, n40643, n40644, n40645, n40646, n40647,
    n40648, n40649, n40650, n40651, n40652, n40653,
    n40654, n40655, n40656, n40657, n40658, n40659,
    n40660, n40661, n40662, n40663, n40665, n40666,
    n40667, n40668, n40669, n40670, n40671, n40672,
    n40673, n40674, n40675, n40676, n40677, n40678,
    n40679, n40680, n40681, n40682, n40683, n40684,
    n40685, n40686, n40687, n40688, n40689, n40690,
    n40691, n40692, n40693, n40694, n40695, n40696,
    n40697, n40698, n40699, n40700, n40701, n40702,
    n40703, n40704, n40705, n40706, n40707, n40708,
    n40709, n40710, n40711, n40713, n40714, n40715,
    n40716, n40717, n40718, n40719, n40720, n40721,
    n40722, n40723, n40724, n40725, n40726, n40727,
    n40728, n40729, n40730, n40731, n40732, n40733,
    n40734, n40735, n40736, n40737, n40738, n40739,
    n40740, n40741, n40742, n40743, n40744, n40745,
    n40746, n40747, n40748, n40749, n40750, n40751,
    n40752, n40753, n40754, n40755, n40756, n40757,
    n40758, n40759, n40760, n40761, n40762, n40763,
    n40764, n40765, n40766, n40767, n40768, n40769,
    n40770, n40771, n40772, n40773, n40774, n40775,
    n40776, n40777, n40778, n40779, n40780, n40781,
    n40782, n40783, n40784, n40785, n40786, n40787,
    n40788, n40789, n40790, n40791, n40792, n40793,
    n40794, n40795, n40796, n40797, n40798, n40799,
    n40800, n40801, n40802, n40803, n40804, n40805,
    n40806, n40807, n40808, n40809, n40810, n40811,
    n40812, n40813, n40814, n40815, n40816, n40817,
    n40818, n40819, n40820, n40821, n40822, n40823,
    n40824, n40825, n40826, n40827, n40828, n40829,
    n40830, n40831, n40832, n40833, n40834, n40835,
    n40836, n40837, n40838, n40839, n40840, n40841,
    n40842, n40843, n40844, n40845, n40846, n40847,
    n40848, n40849, n40850, n40851, n40852, n40853,
    n40854, n40855, n40856, n40857, n40858, n40859,
    n40860, n40861, n40862, n40863, n40864, n40865,
    n40866, n40867, n40868, n40869, n40870, n40871,
    n40872, n40873, n40874, n40875, n40876, n40877,
    n40878, n40879, n40880, n40881, n40882, n40883,
    n40884, n40885, n40886, n40887, n40888, n40889,
    n40890, n40891, n40892, n40893, n40894, n40895,
    n40896, n40897, n40898, n40899, n40900, n40901,
    n40902, n40903, n40904, n40905, n40906, n40907,
    n40908, n40909, n40910, n40911, n40912, n40913,
    n40914, n40915, n40916, n40917, n40918, n40919,
    n40920, n40921, n40922, n40923, n40925, n40926,
    n40927, n40928, n40929, n40930, n40931, n40932,
    n40933, n40934, n40935, n40936, n40937, n40938,
    n40939, n40940, n40941, n40942, n40943, n40944,
    n40945, n40946, n40947, n40948, n40949, n40950,
    n40951, n40952, n40953, n40954, n40955, n40956,
    n40957, n40958, n40959, n40960, n40961, n40962,
    n40963, n40964, n40965, n40966, n40967, n40968,
    n40969, n40970, n40971, n40972, n40973, n40974,
    n40975, n40976, n40977, n40978, n40979, n40980,
    n40981, n40982, n40983, n40984, n40985, n40986,
    n40987, n40988, n40989, n40990, n40991, n40992,
    n40993, n40994, n40995, n40996, n40997, n40998,
    n40999, n41000, n41001, n41002, n41003, n41004,
    n41005, n41006, n41007, n41008, n41009, n41010,
    n41011, n41012, n41013, n41014, n41015, n41016,
    n41017, n41018, n41019, n41020, n41021, n41022,
    n41023, n41024, n41025, n41026, n41027, n41028,
    n41029, n41030, n41031, n41032, n41033, n41034,
    n41035, n41036, n41037, n41038, n41039, n41040,
    n41041, n41042, n41043, n41044, n41045, n41046,
    n41047, n41048, n41049, n41050, n41051, n41052,
    n41053, n41054, n41055, n41056, n41057, n41058,
    n41059, n41060, n41061, n41062, n41063, n41064,
    n41065, n41066, n41067, n41068, n41069, n41070,
    n41071, n41072, n41073, n41074, n41075, n41076,
    n41077, n41078, n41079, n41080, n41081, n41082,
    n41083, n41084, n41085, n41086, n41087, n41088,
    n41089, n41090, n41091, n41092, n41093, n41094,
    n41095, n41096, n41097, n41098, n41099, n41100,
    n41101, n41102, n41103, n41104, n41105, n41106,
    n41107, n41108, n41109, n41110, n41111, n41112,
    n41113, n41114, n41115, n41116, n41117, n41118,
    n41119, n41120, n41121, n41122, n41123, n41124,
    n41125, n41126, n41127, n41128, n41129, n41130,
    n41131, n41132, n41133, n41134, n41135, n41136,
    n41137, n41138, n41139, n41140, n41141, n41142,
    n41143, n41144, n41145, n41146, n41147, n41148,
    n41149, n41150, n41151, n41152, n41153, n41154,
    n41155, n41156, n41157, n41158, n41159, n41160,
    n41161, n41162, n41163, n41164, n41165, n41166,
    n41167, n41168, n41170, n41171, n41172, n41173,
    n41174, n41175, n41176, n41177, n41178, n41179,
    n41180, n41181, n41182, n41183, n41184, n41185,
    n41186, n41187, n41188, n41189, n41190, n41191,
    n41192, n41193, n41194, n41195, n41196, n41197,
    n41198, n41199, n41200, n41201, n41202, n41203,
    n41204, n41205, n41206, n41207, n41208, n41209,
    n41210, n41211, n41212, n41213, n41214, n41215,
    n41216, n41217, n41218, n41219, n41220, n41221,
    n41222, n41223, n41224, n41225, n41226, n41227,
    n41228, n41229, n41230, n41231, n41232, n41233,
    n41234, n41235, n41236, n41237, n41238, n41239,
    n41240, n41241, n41242, n41243, n41244, n41245,
    n41246, n41247, n41248, n41249, n41250, n41251,
    n41252, n41253, n41254, n41255, n41256, n41257,
    n41258, n41259, n41260, n41261, n41262, n41263,
    n41264, n41265, n41266, n41267, n41268, n41269,
    n41270, n41271, n41272, n41273, n41274, n41275,
    n41276, n41277, n41278, n41279, n41280, n41281,
    n41282, n41283, n41284, n41285, n41286, n41287,
    n41288, n41289, n41290, n41291, n41292, n41293,
    n41294, n41295, n41296, n41297, n41298, n41299,
    n41300, n41301, n41302, n41303, n41304, n41305,
    n41306, n41307, n41308, n41309, n41310, n41311,
    n41312, n41313, n41314, n41315, n41316, n41317,
    n41318, n41319, n41320, n41321, n41322, n41323,
    n41324, n41325, n41326, n41327, n41328, n41329,
    n41330, n41331, n41332, n41333, n41334, n41335,
    n41336, n41337, n41338, n41339, n41340, n41341,
    n41342, n41343, n41344, n41345, n41346, n41347,
    n41348, n41349, n41350, n41351, n41352, n41353,
    n41354, n41355, n41356, n41357, n41358, n41359,
    n41360, n41361, n41362, n41363, n41364, n41365,
    n41366, n41367, n41368, n41369, n41370, n41371,
    n41372, n41373, n41374, n41375, n41376, n41377,
    n41378, n41379, n41380, n41381, n41382, n41383,
    n41384, n41385, n41386, n41387, n41388, n41389,
    n41390, n41391, n41393, n41394, n41395, n41396,
    n41397, n41398, n41399, n41400, n41401, n41402,
    n41403, n41404, n41405, n41406, n41407, n41408,
    n41409, n41410, n41411, n41412, n41413, n41414,
    n41415, n41416, n41417, n41418, n41419, n41420,
    n41421, n41422, n41423, n41424, n41425, n41426,
    n41427, n41428, n41429, n41430, n41431, n41432,
    n41433, n41434, n41435, n41436, n41437, n41438,
    n41439, n41440, n41441, n41442, n41443, n41444,
    n41445, n41446, n41447, n41448, n41449, n41450,
    n41451, n41452, n41453, n41454, n41455, n41456,
    n41457, n41458, n41459, n41460, n41461, n41462,
    n41463, n41464, n41465, n41466, n41467, n41468,
    n41469, n41470, n41471, n41472, n41473, n41474,
    n41475, n41476, n41477, n41478, n41479, n41480,
    n41481, n41482, n41483, n41484, n41485, n41486,
    n41487, n41488, n41489, n41490, n41491, n41492,
    n41493, n41494, n41495, n41496, n41497, n41498,
    n41499, n41500, n41501, n41502, n41503, n41504,
    n41505, n41506, n41507, n41508, n41509, n41510,
    n41511, n41512, n41513, n41514, n41515, n41516,
    n41517, n41518, n41519, n41520, n41521, n41522,
    n41523, n41524, n41525, n41526, n41527, n41528,
    n41529, n41530, n41531, n41532, n41533, n41534,
    n41535, n41536, n41537, n41538, n41539, n41540,
    n41541, n41542, n41543, n41544, n41545, n41546,
    n41547, n41548, n41549, n41550, n41551, n41553,
    n41554, n41555, n41556, n41557, n41558, n41559,
    n41560, n41561, n41562, n41563, n41564, n41565,
    n41566, n41567, n41568, n41569, n41570, n41571,
    n41572, n41573, n41574, n41575, n41576, n41577,
    n41578, n41579, n41580, n41581, n41582, n41583,
    n41584, n41585, n41586, n41587, n41588, n41589,
    n41590, n41591, n41592, n41593, n41594, n41595,
    n41596, n41597, n41598, n41599, n41600, n41601,
    n41602, n41603, n41604, n41605, n41606, n41607,
    n41608, n41609, n41610, n41611, n41612, n41613,
    n41614, n41615, n41616, n41617, n41618, n41619,
    n41620, n41621, n41622, n41623, n41624, n41625,
    n41626, n41627, n41628, n41629, n41630, n41631,
    n41632, n41633, n41634, n41635, n41636, n41637,
    n41638, n41639, n41640, n41641, n41642, n41643,
    n41644, n41645, n41646, n41647, n41648, n41649,
    n41650, n41651, n41652, n41653, n41654, n41655,
    n41656, n41657, n41658, n41659, n41660, n41661,
    n41662, n41663, n41664, n41665, n41666, n41667,
    n41668, n41669, n41670, n41671, n41672, n41673,
    n41674, n41675, n41676, n41677, n41678, n41679,
    n41680, n41681, n41682, n41683, n41684, n41685,
    n41686, n41687, n41688, n41689, n41690, n41691,
    n41692, n41693, n41694, n41695, n41696, n41697,
    n41698, n41699, n41700, n41701, n41702, n41703,
    n41704, n41705, n41706, n41707, n41708, n41709,
    n41710, n41711, n41712, n41713, n41714, n41715,
    n41716, n41718, n41719, n41720, n41721, n41722,
    n41723, n41724, n41726, n41727, n41728, n41729,
    n41730, n41731, n41732, n41733, n41734, n41736,
    n41737, n41738, n41739, n41740, n41741, n41742,
    n41743, n41744, n41745, n41746, n41747, n41748,
    n41749, n41750, n41751, n41752, n41753, n41754,
    n41755, n41756, n41757, n41758, n41759, n41760,
    n41761, n41762, n41763, n41764, n41765, n41766,
    n41767, n41768, n41769, n41770, n41771, n41772,
    n41773, n41774, n41775, n41776, n41778, n41779,
    n41780, n41781, n41782, n41783, n41784, n41785,
    n41786, n41787, n41788, n41789, n41790, n41791,
    n41792, n41793, n41794, n41795, n41796, n41797,
    n41798, n41799, n41800, n41801, n41802, n41803,
    n41804, n41805, n41806, n41807, n41808, n41809,
    n41810, n41811, n41812, n41813, n41814, n41815,
    n41816, n41817, n41818, n41819, n41820, n41821,
    n41822, n41823, n41824, n41825, n41826, n41827,
    n41828, n41829, n41830, n41831, n41832, n41833,
    n41834, n41835, n41836, n41837, n41838, n41839,
    n41840, n41841, n41842, n41843, n41844, n41845,
    n41846, n41847, n41848, n41849, n41850, n41851,
    n41852, n41853, n41854, n41855, n41856, n41857,
    n41858, n41859, n41860, n41861, n41862, n41863,
    n41864, n41865, n41866, n41867, n41868, n41869,
    n41870, n41871, n41872, n41873, n41874, n41875,
    n41876, n41877, n41878, n41879, n41880, n41881,
    n41882, n41883, n41884, n41885, n41886, n41887,
    n41888, n41889, n41890, n41891, n41892, n41893,
    n41894, n41895, n41896, n41897, n41898, n41899,
    n41900, n41901, n41902, n41903, n41904, n41905,
    n41906, n41907, n41908, n41909, n41910, n41911,
    n41912, n41913, n41914, n41915, n41916, n41917,
    n41918, n41919, n41920, n41921, n41922, n41923,
    n41924, n41925, n41926, n41927, n41928, n41929,
    n41930, n41931, n41932, n41933, n41934, n41935,
    n41936, n41937, n41938, n41939, n41940, n41941,
    n41942, n41943, n41944, n41945, n41946, n41947,
    n41948, n41949, n41950, n41951, n41952, n41953,
    n41954, n41955, n41956, n41957, n41958, n41959,
    n41960, n41961, n41962, n41963, n41964, n41965,
    n41966, n41967, n41968, n41969, n41970, n41971,
    n41972, n41973, n41974, n41975, n41976, n41977,
    n41978, n41979, n41980, n41981, n41982, n41983,
    n41984, n41985, n41986, n41987, n41988, n41989,
    n41990, n41991, n41992, n41993, n41994, n41995,
    n41996, n41997, n41998, n41999, n42000, n42001,
    n42002, n42003, n42004, n42005, n42006, n42008,
    n42009, n42010, n42011, n42012, n42013, n42014,
    n42015, n42016, n42017, n42018, n42019, n42020,
    n42021, n42022, n42023, n42024, n42025, n42026,
    n42027, n42028, n42029, n42030, n42031, n42032,
    n42033, n42034, n42035, n42036, n42037, n42038,
    n42039, n42040, n42041, n42042, n42043, n42044,
    n42045, n42046, n42047, n42048, n42049, n42050,
    n42051, n42052, n42053, n42054, n42055, n42056,
    n42057, n42058, n42059, n42060, n42061, n42062,
    n42063, n42064, n42065, n42066, n42067, n42068,
    n42069, n42070, n42071, n42072, n42073, n42074,
    n42075, n42076, n42077, n42078, n42079, n42080,
    n42081, n42082, n42083, n42084, n42085, n42086,
    n42087, n42088, n42089, n42090, n42091, n42092,
    n42093, n42094, n42095, n42096, n42097, n42098,
    n42099, n42100, n42101, n42102, n42103, n42104,
    n42105, n42106, n42107, n42108, n42109, n42110,
    n42111, n42112, n42113, n42114, n42115, n42116,
    n42117, n42118, n42119, n42120, n42121, n42122,
    n42123, n42124, n42125, n42126, n42127, n42128,
    n42129, n42130, n42131, n42132, n42133, n42134,
    n42135, n42136, n42137, n42138, n42139, n42140,
    n42141, n42142, n42143, n42144, n42145, n42146,
    n42147, n42148, n42149, n42150, n42151, n42152,
    n42153, n42154, n42155, n42156, n42157, n42158,
    n42159, n42160, n42161, n42162, n42163, n42164,
    n42165, n42166, n42167, n42168, n42169, n42170,
    n42171, n42172, n42173, n42174, n42175, n42176,
    n42177, n42178, n42179, n42180, n42181, n42182,
    n42183, n42184, n42185, n42186, n42187, n42188,
    n42189, n42190, n42191, n42192, n42193, n42194,
    n42195, n42196, n42197, n42198, n42199, n42200,
    n42201, n42202, n42203, n42204, n42205, n42206,
    n42207, n42208, n42209, n42210, n42211, n42212,
    n42213, n42214, n42215, n42216, n42217, n42218,
    n42219, n42220, n42221, n42222, n42223, n42224,
    n42225, n42226, n42227, n42228, n42229, n42230,
    n42231, n42232, n42233, n42235, n42236, n42237,
    n42238, n42239, n42241, n42242, n42243, n42244,
    n42245, n42247, n42248, n42249, n42250, n42251,
    n42253, n42254, n42255, n42256, n42257, n42259,
    n42260, n42261, n42262, n42263, n42265, n42266,
    n42267, n42268, n42269, n42270, n42272, n42273,
    n42274, n42275, n42276, n42277, n42279, n42280,
    n42281, n42282, n42283, n42284, n42285, n42286,
    n42287, n42288, n42289, n42290, n42291, n42292,
    n42293, n42294, n42295, n42296, n42297, n42298,
    n42299, n42300, n42301, n42302, n42303, n42304,
    n42305, n42306, n42307, n42308, n42309, n42310,
    n42311, n42313, n42314, n42315, n42316, n42317,
    n42318, n42319, n42320, n42321, n42322, n42323,
    n42324, n42325, n42326, n42327, n42328, n42329,
    n42330, n42331, n42332, n42333, n42334, n42335,
    n42336, n42337, n42338, n42339, n42340, n42341,
    n42342, n42343, n42344, n42345, n42346, n42347,
    n42348, n42349, n42350, n42351, n42352, n42353,
    n42354, n42355, n42356, n42357, n42358, n42359,
    n42360, n42361, n42362, n42363, n42364, n42365,
    n42366, n42367, n42368, n42369, n42370, n42371,
    n42372, n42373, n42374, n42375, n42376, n42377,
    n42378, n42379, n42380, n42381, n42382, n42383,
    n42384, n42385, n42386, n42387, n42388, n42389,
    n42390, n42391, n42392, n42393, n42394, n42395,
    n42396, n42397, n42398, n42399, n42400, n42401,
    n42402, n42403, n42404, n42405, n42406, n42407,
    n42408, n42409, n42410, n42411, n42412, n42413,
    n42414, n42415, n42416, n42417, n42418, n42419,
    n42420, n42421, n42422, n42423, n42424, n42425,
    n42426, n42427, n42428, n42429, n42430, n42431,
    n42432, n42433, n42434, n42435, n42436, n42437,
    n42438, n42439, n42440, n42441, n42442, n42443,
    n42444, n42445, n42446, n42447, n42448, n42449,
    n42450, n42451, n42452, n42453, n42454, n42455,
    n42456, n42457, n42458, n42459, n42460, n42461,
    n42462, n42463, n42464, n42465, n42466, n42467,
    n42468, n42469, n42470, n42471, n42472, n42473,
    n42474, n42475, n42476, n42477, n42478, n42479,
    n42480, n42481, n42482, n42483, n42484, n42485,
    n42486, n42487, n42488, n42489, n42490, n42491,
    n42492, n42493, n42494, n42495, n42496, n42497,
    n42498, n42499, n42500, n42501, n42502, n42503,
    n42504, n42505, n42506, n42507, n42508, n42509,
    n42510, n42511, n42512, n42513, n42514, n42515,
    n42516, n42517, n42519, n42520, n42521, n42522,
    n42523, n42524, n42525, n42526, n42527, n42528,
    n42529, n42530, n42531, n42532, n42533, n42534,
    n42535, n42536, n42537, n42538, n42539, n42540,
    n42541, n42542, n42543, n42544, n42545, n42546,
    n42547, n42548, n42549, n42550, n42551, n42552,
    n42553, n42554, n42555, n42556, n42557, n42558,
    n42559, n42560, n42561, n42562, n42564, n42565,
    n42566, n42567, n42568, n42569, n42570, n42571,
    n42572, n42573, n42574, n42575, n42576, n42577,
    n42578, n42579, n42580, n42581, n42582, n42583,
    n42584, n42585, n42586, n42587, n42588, n42589,
    n42590, n42591, n42592, n42593, n42594, n42595,
    n42596, n42597, n42598, n42599, n42600, n42601,
    n42602, n42603, n42605, n42606, n42607, n42608,
    n42609, n42610, n42611, n42612, n42613, n42614,
    n42615, n42616, n42617, n42618, n42619, n42620,
    n42621, n42622, n42623, n42624, n42625, n42626,
    n42627, n42628, n42629, n42630, n42631, n42632,
    n42633, n42634, n42635, n42636, n42637, n42638,
    n42639, n42640, n42641, n42642, n42643, n42644,
    n42645, n42646, n42647, n42648, n42649, n42650,
    n42651, n42652, n42653, n42654, n42655, n42656,
    n42657, n42658, n42659, n42660, n42661, n42662,
    n42663, n42664, n42665, n42666, n42667, n42668,
    n42669, n42671, n42672, n42673, n42674, n42675,
    n42676, n42677, n42678, n42679, n42680, n42681,
    n42682, n42683, n42684, n42685, n42686, n42687,
    n42688, n42689, n42690, n42691, n42692, n42693,
    n42694, n42695, n42696, n42697, n42698, n42699,
    n42700, n42701, n42702, n42703, n42704, n42705,
    n42706, n42707, n42708, n42709, n42710, n42711,
    n42712, n42713, n42714, n42715, n42716, n42717,
    n42718, n42719, n42720, n42721, n42722, n42723,
    n42724, n42725, n42726, n42727, n42728, n42729,
    n42730, n42731, n42732, n42733, n42734, n42735,
    n42736, n42737, n42738, n42739, n42740, n42741,
    n42742, n42743, n42744, n42745, n42746, n42747,
    n42748, n42749, n42750, n42751, n42752, n42753,
    n42754, n42755, n42756, n42757, n42758, n42759,
    n42760, n42761, n42762, n42763, n42764, n42765,
    n42766, n42767, n42768, n42769, n42770, n42771,
    n42772, n42773, n42774, n42775, n42776, n42777,
    n42778, n42779, n42780, n42781, n42782, n42783,
    n42784, n42785, n42786, n42787, n42788, n42789,
    n42790, n42791, n42792, n42793, n42794, n42795,
    n42796, n42797, n42798, n42799, n42800, n42801,
    n42802, n42803, n42804, n42805, n42806, n42807,
    n42808, n42809, n42810, n42811, n42812, n42813,
    n42814, n42815, n42816, n42817, n42818, n42819,
    n42820, n42821, n42822, n42823, n42824, n42825,
    n42826, n42827, n42828, n42829, n42830, n42831,
    n42832, n42833, n42834, n42835, n42836, n42837,
    n42838, n42839, n42840, n42841, n42842, n42843,
    n42844, n42845, n42846, n42847, n42848, n42849,
    n42850, n42851, n42852, n42853, n42854, n42855,
    n42856, n42857, n42858, n42859, n42860, n42861,
    n42862, n42863, n42864, n42865, n42866, n42867,
    n42868, n42869, n42871, n42872, n42873, n42874,
    n42875, n42876, n42877, n42878, n42879, n42880,
    n42881, n42882, n42883, n42884, n42885, n42886,
    n42887, n42888, n42889, n42890, n42891, n42892,
    n42893, n42894, n42895, n42896, n42897, n42898,
    n42899, n42900, n42901, n42902, n42903, n42904,
    n42905, n42906, n42907, n42908, n42909, n42910,
    n42911, n42912, n42913, n42914, n42915, n42916,
    n42917, n42918, n42919, n42920, n42921, n42922,
    n42923, n42924, n42925, n42926, n42927, n42928,
    n42929, n42930, n42931, n42932, n42933, n42934,
    n42935, n42936, n42937, n42938, n42939, n42940,
    n42941, n42942, n42943, n42944, n42945, n42946,
    n42947, n42948, n42949, n42950, n42951, n42952,
    n42953, n42954, n42955, n42956, n42957, n42958,
    n42959, n42960, n42961, n42962, n42963, n42964,
    n42965, n42966, n42967, n42968, n42969, n42970,
    n42971, n42972, n42973, n42974, n42975, n42976,
    n42977, n42978, n42979, n42980, n42981, n42982,
    n42983, n42984, n42985, n42986, n42987, n42988,
    n42989, n42990, n42991, n42992, n42993, n42994,
    n42995, n42996, n42997, n42998, n42999, n43000,
    n43001, n43002, n43003, n43004, n43005, n43006,
    n43007, n43008, n43009, n43010, n43011, n43012,
    n43013, n43014, n43015, n43016, n43017, n43018,
    n43019, n43020, n43021, n43023, n43024, n43025,
    n43026, n43027, n43028, n43029, n43030, n43031,
    n43032, n43033, n43034, n43035, n43036, n43037,
    n43038, n43039, n43040, n43041, n43042, n43043,
    n43044, n43045, n43046, n43047, n43048, n43049,
    n43050, n43051, n43052, n43053, n43054, n43055,
    n43056, n43057, n43058, n43059, n43060, n43061,
    n43062, n43063, n43064, n43065, n43066, n43068,
    n43069, n43070, n43071, n43072, n43073, n43074,
    n43075, n43076, n43077, n43078, n43079, n43080,
    n43081, n43082, n43083, n43084, n43085, n43086,
    n43087, n43088, n43089, n43090, n43091, n43092,
    n43093, n43094, n43095, n43096, n43097, n43098,
    n43099, n43100, n43101, n43102, n43103, n43104,
    n43105, n43106, n43107, n43108, n43109, n43110,
    n43112, n43113, n43114, n43115, n43116, n43117,
    n43118, n43119, n43120, n43121, n43122, n43123,
    n43124, n43125, n43126, n43127, n43128, n43129,
    n43130, n43131, n43132, n43133, n43134, n43135,
    n43136, n43137, n43138, n43139, n43140, n43141,
    n43142, n43143, n43144, n43145, n43146, n43147,
    n43148, n43149, n43150, n43151, n43152, n43153,
    n43154, n43155, n43156, n43157, n43159, n43160,
    n43161, n43162, n43163, n43164, n43165, n43166,
    n43167, n43168, n43169, n43170, n43171, n43172,
    n43173, n43174, n43175, n43176, n43177, n43178,
    n43179, n43180, n43181, n43182, n43183, n43184,
    n43185, n43186, n43187, n43188, n43189, n43190,
    n43191, n43192, n43193, n43194, n43195, n43196,
    n43197, n43198, n43199, n43200, n43201, n43202,
    n43203, n43204, n43205, n43206, n43207, n43208,
    n43209, n43210, n43211, n43212, n43213, n43214,
    n43215, n43216, n43217, n43218, n43219, n43220,
    n43221, n43222, n43223, n43224, n43225, n43226,
    n43227, n43228, n43229, n43230, n43231, n43232,
    n43233, n43235, n43236, n43237, n43238, n43239,
    n43240, n43241, n43242, n43243, n43244, n43245,
    n43246, n43247, n43248, n43249, n43250, n43251,
    n43252, n43253, n43254, n43255, n43256, n43257,
    n43258, n43259, n43260, n43261, n43262, n43263,
    n43264, n43265, n43266, n43267, n43268, n43269,
    n43270, n43271, n43272, n43273, n43274, n43275,
    n43276, n43277, n43278, n43279, n43280, n43281,
    n43282, n43283, n43284, n43285, n43286, n43287,
    n43288, n43289, n43290, n43291, n43292, n43293,
    n43294, n43295, n43297, n43298, n43299, n43300,
    n43301, n43302, n43303, n43304, n43305, n43306,
    n43307, n43308, n43309, n43310, n43311, n43312,
    n43313, n43314, n43315, n43316, n43317, n43318,
    n43319, n43320, n43321, n43322, n43323, n43324,
    n43325, n43326, n43327, n43328, n43329, n43330,
    n43331, n43332, n43333, n43334, n43335, n43336,
    n43338, n43339, n43340, n43341, n43342, n43343,
    n43344, n43345, n43346, n43347, n43348, n43349,
    n43350, n43351, n43352, n43353, n43354, n43355,
    n43356, n43357, n43358, n43359, n43360, n43361,
    n43362, n43363, n43364, n43365, n43366, n43367,
    n43368, n43369, n43370, n43371, n43372, n43373,
    n43374, n43375, n43376, n43377, n43378, n43379,
    n43380, n43381, n43382, n43383, n43384, n43385,
    n43386, n43387, n43388, n43389, n43390, n43391,
    n43392, n43393, n43394, n43395, n43397, n43398,
    n43399, n43400, n43401, n43402, n43403, n43404,
    n43405, n43406, n43407, n43408, n43409, n43410,
    n43411, n43412, n43413, n43414, n43415, n43416,
    n43417, n43418, n43419, n43420, n43421, n43422,
    n43423, n43424, n43425, n43427, n43428, n43429,
    n43430, n43431, n43432, n43433, n43434, n43435,
    n43436, n43437, n43438, n43439, n43440, n43441,
    n43442, n43443, n43444, n43445, n43446, n43447,
    n43448, n43449, n43450, n43451, n43452, n43453,
    n43454, n43455, n43456, n43457, n43458, n43459,
    n43460, n43461, n43462, n43463, n43464, n43465,
    n43466, n43467, n43468, n43470, n43471, n43472,
    n43473, n43474, n43475, n43476, n43477, n43478,
    n43479, n43480, n43481, n43482, n43483, n43484,
    n43485, n43486, n43487, n43488, n43489, n43490,
    n43491, n43492, n43493, n43494, n43495, n43496,
    n43497, n43498, n43499, n43500, n43501, n43502,
    n43503, n43504, n43505, n43506, n43507, n43508,
    n43509, n43510, n43511, n43512, n43513, n43514,
    n43515, n43516, n43517, n43518, n43519, n43520,
    n43521, n43522, n43523, n43524, n43525, n43526,
    n43527, n43528, n43529, n43530, n43531, n43532,
    n43533, n43534, n43535, n43536, n43538, n43539,
    n43540, n43541, n43542, n43543, n43544, n43545,
    n43546, n43547, n43548, n43549, n43550, n43551,
    n43552, n43553, n43554, n43555, n43556, n43557,
    n43558, n43559, n43560, n43561, n43562, n43563,
    n43564, n43565, n43566, n43567, n43568, n43569,
    n43570, n43571, n43572, n43573, n43574, n43575,
    n43576, n43577, n43578, n43579, n43580, n43581,
    n43582, n43583, n43584, n43585, n43586, n43587,
    n43588, n43589, n43590, n43591, n43592, n43593,
    n43594, n43595, n43597, n43598, n43599, n43600,
    n43601, n43602, n43603, n43604, n43605, n43606,
    n43607, n43608, n43609, n43610, n43611, n43612,
    n43613, n43614, n43615, n43616, n43617, n43618,
    n43619, n43620, n43621, n43622, n43623, n43624,
    n43625, n43626, n43627, n43628, n43629, n43630,
    n43631, n43632, n43633, n43634, n43635, n43636,
    n43637, n43638, n43639, n43641, n43642, n43643,
    n43644, n43645, n43646, n43647, n43648, n43649,
    n43650, n43651, n43652, n43653, n43654, n43655,
    n43656, n43657, n43658, n43659, n43660, n43661,
    n43662, n43663, n43664, n43665, n43666, n43667,
    n43668, n43669, n43670, n43671, n43672, n43673,
    n43674, n43675, n43676, n43677, n43678, n43680,
    n43681, n43682, n43683, n43684, n43685, n43686,
    n43687, n43688, n43689, n43690, n43691, n43692,
    n43693, n43694, n43695, n43696, n43697, n43698,
    n43699, n43700, n43701, n43702, n43703, n43704,
    n43705, n43706, n43707, n43708, n43709, n43710,
    n43711, n43712, n43713, n43714, n43715, n43716,
    n43717, n43719, n43720, n43721, n43722, n43723,
    n43724, n43725, n43726, n43727, n43728, n43729,
    n43730, n43731, n43732, n43733, n43734, n43735,
    n43736, n43737, n43738, n43739, n43740, n43741,
    n43742, n43743, n43744, n43745, n43746, n43747,
    n43748, n43749, n43750, n43751, n43752, n43753,
    n43754, n43755, n43756, n43757, n43758, n43759,
    n43760, n43761, n43762, n43763, n43764, n43765,
    n43766, n43767, n43768, n43769, n43770, n43771,
    n43772, n43773, n43774, n43775, n43776, n43778,
    n43779, n43780, n43782, n43783, n43784, n43785,
    n43786, n43787, n43788, n43789, n43790, n43791,
    n43792, n43793, n43794, n43795, n43796, n43797,
    n43798, n43799, n43801, n43802, n43803, n43804,
    n43805, n43806, n43807, n43808, n43809, n43810,
    n43811, n43812, n43813, n43814, n43815, n43816,
    n43817, n43819, n43821, n43822, n43824, n43825,
    n43826, n43828, n43829, n43830, n43831, n43832,
    n43833, n43834, n43835, n43836, n43837, n43838,
    n43839, n43841, n43842, n43844, n43845, n43847,
    n43848, n43850, n43851, n43853, n43854, n43856,
    n43857, n43859, n43860, n43862, n43863, n43865,
    n43866, n43868, n43869, n43870, n43871, n43872,
    n43873, n43874, n43876, n43877, n43878, n43879,
    n43880, n43881, n43883, n43884, n43885, n43887,
    n43888, n43889, n43890, n43891, n43892, n43893,
    n43894, n43895, n43896, n43897, n43898, n43899,
    n43900, n43901, n43902, n43903, n43904, n43905,
    n43906, n43907, n43909, n43910, n43912, n43913,
    n43915, n43916, n43918, n43919, n43921, n43922,
    n43924, n43925, n43927, n43928, n43930, n43931,
    n43932, n43933, n43934, n43935, n43936, n43937,
    n43938, n43939, n43940, n43941, n43942, n43943,
    n43944, n43945, n43946, n43947, n43948, n43949,
    n43950, n43951, n43952, n43953, n43954, n43956,
    n43957, n43958, n43960, n43961, n43963, n43964,
    n43965, n43967, n43968, n43970, n43971, n43972,
    n43973, n43974, n43975, n43976, n43977, n43978,
    n43979, n43980, n43982, n43983, n43984, n43985,
    n43987, n43988, n43990, n43991, n43992, n43994,
    n43995, n43996, n43997, n43999, n44000, n44002,
    n44003, n44005, n44006, n44008, n44009, n44011,
    n44012, n44014, n44015, n44017, n44018, n44020,
    n44021, n44023, n44024, n44026, n44027, n44029,
    n44030, n44032, n44033, n44034, n44035, n44036,
    n44037, n44038, n44040, n44041, n44042, n44043,
    n44045, n44046, n44047, n44048, n44049, n44050,
    n44051, n44052, n44053, n44054, n44055, n44057,
    n44058, n44060, n44061, n44063, n44064, n44066,
    n44067, n44069, n44070, n44072, n44073, n44075,
    n44076, n44078, n44079, n44080, n44081, n44082,
    n44084, n44085, n44087, n44088, n44090, n44091,
    n44093, n44094, n44096, n44097, n44099, n44100,
    n44102, n44103, n44105, n44106, n44108, n44109,
    n44111, n44112, n44114, n44115, n44117, n44118,
    n44120, n44121, n44123, n44124, n44126, n44127,
    n44129, n44130, n44132, n44133, n44135, n44136,
    n44138, n44139, n44141, n44142, n44144, n44145,
    n44147, n44148, n44150, n44151, n44153, n44154,
    n44156, n44157, n44159, n44160, n44162, n44163,
    n44165, n44166, n44168, n44169, n44171, n44172,
    n44174, n44175, n44177, n44178, n44180, n44181,
    n44183, n44184, n44186, n44187, n44189, n44190,
    n44192, n44193, n44195, n44196, n44198, n44199,
    n44201, n44202, n44204, n44205, n44207, n44208,
    n44210, n44211, n44213, n44214, n44216, n44217,
    n44219, n44220, n44222, n44223, n44225, n44226,
    n44228, n44229, n44231, n44232, n44234, n44235,
    n44237, n44238, n44240, n44241, n44243, n44244,
    n44246, n44247, n44249, n44250, n44252, n44253,
    n44255, n44256, n44258, n44259, n44261, n44262,
    n44264, n44265, n44267, n44268, n44270, n44271,
    n44273, n44274, n44276, n44277, n44279, n44280,
    n44282, n44283, n44285, n44286, n44288, n44289,
    n44291, n44292, n44294, n44295, n44297, n44298,
    n44300, n44301, n44303, n44304, n44305, n44307,
    n44308, n44310, n44311, n44313, n44314, n44316,
    n44317, n44319, n44320, n44322, n44323, n44325,
    n44326, n44328, n44329, n44331, n44332, n44334,
    n44335, n44337, n44338, n44340, n44341, n44343,
    n44344, n44346, n44347, n44349, n44350, n44352,
    n44353, n44355, n44356, n44358, n44359, n44361,
    n44362, n44364, n44365, n44367, n44368, n44370,
    n44371, n44373, n44374, n44376, n44377, n44379,
    n44380, n44382, n44383, n44385, n44386, n44388,
    n44389, n44391, n44392, n44394, n44395, n44397,
    n44398, n44400, n44401, n44403, n44404, n44406,
    n44407, n44409, n44410, n44412, n44413, n44415,
    n44416, n44418, n44419, n44421, n44422, n44424,
    n44425, n44427, n44428, n44430, n44431, n44433,
    n44434, n44435, n44436, n44437, n44438, n44439,
    n44440, n44441, n44442, n44443, n44444, n44445,
    n44446, n44447, n44448, n44449, n44450, n44451,
    n44452, n44453, n44454, n44455, n44457, n44458,
    n44460, n44461, n44463, n44464, n44466, n44467,
    n44469, n44470, n44472, n44473, n44475, n44476,
    n44478, n44479, n44480, n44481, n44482, n44483,
    n44484, n44485, n44486, n44487, n44488, n44489,
    n44490, n44491, n44492, n44493, n44494, n44495,
    n44496, n44497, n44498, n44499, n44500, n44501,
    n44503, n44504, n44505, n44506, n44507, n44508,
    n44509, n44510, n44511, n44512, n44513, n44514,
    n44515, n44516, n44517, n44518, n44520, n44521,
    n44522, n44523, n44524, n44525, n44526, n44527,
    n44528, n44529, n44530, n44531, n44532, n44533,
    n44534, n44535, n44536, n44537, n44538, n44539,
    n44540, n44541, n44542, n44543, n44544, n44545,
    n44546, n44547, n44548, n44550, n44551, n44552,
    n44553, n44554, n44556, n44557, n44558, n44559,
    n44560, n44561, n44562, n44563, n44564, n44565,
    n44566, n44567, n44568, n44569, n44570, n44571,
    n44572, n44573, n44574, n44576, n44577, n44578,
    n44579, n44580, n44581, n44582, n44583, n44584,
    n44585, n44586, n44587, n44588, n44589, n44590,
    n44591, n44592, n44593, n44594, n44596, n44597,
    n44598, n44599, n44600, n44601, n44602, n44603,
    n44604, n44605, n44606, n44607, n44608, n44609,
    n44610, n44611, n44612, n44613, n44614, n44616,
    n44617, n44618, n44619, n44620, n44621, n44622,
    n44623, n44624, n44625, n44626, n44627, n44628,
    n44629, n44630, n44631, n44632, n44633, n44634,
    n44636, n44637, n44638, n44639, n44640, n44641,
    n44642, n44643, n44644, n44645, n44647, n44648,
    n44649, n44650, n44651, n44652, n44653, n44654,
    n44655, n44656, n44658, n44659, n44660, n44661,
    n44662, n44663, n44664, n44665, n44666, n44667,
    n44669, n44670, n44671, n44672, n44673, n44674,
    n44675, n44676, n44677, n44678, n44679, n44682,
    n44683, n44685, n44686, n44688, n44689, n44691,
    n44692, n44694, n44695, n44697, n44698, n44700,
    n44701, n44703, n44704, n44706, n44707, n44709,
    n44710, n44712, n44713, n44715, n44716, n44718,
    n44719, n44721, n44722, n44724, n44725, n44727,
    n44728, n44730, n44731, n44733, n44734, n44736,
    n44737, n44739, n44740, n44742, n44743, n44745,
    n44746, n44748, n44749, n44751, n44752, n44754,
    n44755, n44756, n44757, n44758, n44759, n44761,
    n44762, n44764, n44765, n44767, n44768, n44770,
    n44771, n44773, n44774, n44776, n44777, n44778,
    n44780, n44781, n44783, n44784, n44786, n44787,
    n44789, n44790, n44792, n44793, n44795, n44796,
    n44798, n44799, n44800, n44801, n44802, n44804,
    n44805, n44807, n44808, n44810, n44811, n44813,
    n44814, n44816, n44817, n44818, n44819, n44821,
    n44822, n44824, n44825, n44827, n44828, n44830,
    n44831, n44833, n44834, n44836, n44837, n44839,
    n44840, n44842, n44843, n44845, n44846, n44848,
    n44849, n44851, n44852, n44854, n44855, n44857,
    n44858, n44860, n44861, n44863, n44864, n44866,
    n44867, n44869, n44870, n44872, n44873, n44875,
    n44876, n44878, n44879, n44881, n44882, n44883,
    n44884, n44886, n44887, n44889, n44890, n44892,
    n44893, n44895, n44896, n44898, n44899, n44901,
    n44902, n44904, n44905, n44907, n44908, n44910,
    n44911, n44913, n44914, n44916, n44917, n44919,
    n44920, n44922, n44923, n44924, n44925, n44927,
    n44928, n44930, n44931, n44933, n44934, n44936,
    n44937, n44939, n44940, n44942, n44943, n44945,
    n44946, n44948, n44949, n44951, n44952, n44954,
    n44955, n44956, n44957, n44958, n44959, n44960,
    n44961, n44962, n44963, n44964, n44965, n44966,
    n44967, n44968, n44969, n44970, n44971, n44972,
    n44973, n44974, n44975, n44976, n44977, n44978,
    n44979, n44980, n44981, n44982, n44983, n44984,
    n44985, n44986, n44987, n44988, n44989, n44990,
    n44991, n44992, n44993, n44994, n44995, n44996,
    n44997, n44998, n44999, n45000, n45001, n45002,
    n45003, n45004, n45005, n45006, n45007, n45008,
    n45009, n45010, n45011, n45012, n45013, n45014,
    n45015, n45016, n45017, n45018, n45019, n45020,
    n45021, n45022, n45023, n45024, n45025, n45026,
    n45027, n45028, n45029, n45030, n45031, n45032,
    n45033, n45034, n45035, n45036, n45037, n45038,
    n45039, n45040, n45041, n45042, n45043, n45044,
    n45045, n45046, n45047, n45048, n45049, n45050,
    n45051, n45052, n45053, n45054, n45055, n45056,
    n45057, n45058, n45059, n45061, n45062, n45064,
    n45065, n45067, n45068, n45069, n45070, n45072,
    n45073, n45075, n45076, n45078, n45079, n45081,
    n45082, n45084, n45085, n45087, n45088, n45090,
    n45091, n45093, n45094, n45096, n45097, n45099,
    n45100, n45102, n45103, n45105, n45106, n45108,
    n45109, n45111, n45112, n45114, n45115, n45117,
    n45118, n45119, n45120, n45121, n45122, n45124,
    n45125, n45126, n45127, n45129, n45130, n45131,
    n45132, n45133, n45134, n45135, n45136, n45137,
    n45138, n45139, n45140, n45141, n45142, n45143,
    n45144, n45145, n45146, n45147, n45148, n45150,
    n45151, n45152, n45154, n45155, n45156, n45158,
    n45159, n45160, n45162, n45163, n45164, n45165,
    n45166, n45167, n45168, n45169, n45170, n45171,
    n45172, n45173, n45174, n45175, n45176, n45177,
    n45178, n45179, n45180, n45181, n45182, n45183,
    n45184, n45185, n45186, n45187, n45188, n45189,
    n45190, n45191, n45192, n45193, n45194, n45195,
    n45196, n45197, n45198, n45199, n45200, n45201,
    n45202, n45203, n45204, n45205, n45206, n45207,
    n45208, n45209, n45210, n45211, n45212, n45213,
    n45214, n45215, n45216, n45217, n45218, n45219,
    n45220, n45221, n45222, n45223, n45224, n45225,
    n45226, n45227, n45228, n45229, n45230, n45231,
    n45232, n45233, n45234, n45235, n45236, n45237,
    n45238, n45239, n45240, n45241, n45242, n45243,
    n45244, n45245, n45246, n45247, n45248, n45249,
    n45250, n45251, n45252, n45253, n45254, n45255,
    n45256, n45257, n45258, n45259, n45260, n45261,
    n45262, n45263, n45264, n45265, n45266, n45267,
    n45268, n45269, n45270, n45271, n45272, n45273,
    n45274, n45275, n45276, n45277, n45278, n45279,
    n45280, n45281, n45282, n45283, n45284, n45285,
    n45286, n45287, n45288, n45289, n45290, n45291,
    n45292, n45293, n45294, n45295, n45296, n45297,
    n45298, n45299, n45300, n45301, n45302, n45303,
    n45304, n45305, n45306, n45307, n45308, n45309,
    n45310, n45311, n45312, n45313, n45314, n45315,
    n45316, n45317, n45318, n45319, n45320, n45321,
    n45322, n45323, n45324, n45325, n45326, n45327,
    n45328, n45329, n45330, n45331, n45332, n45333,
    n45334, n45335, n45336, n45337, n45338, n45339,
    n45340, n45341, n45342, n45343, n45344, n45345,
    n45346, n45347, n45348, n45349, n45350, n45351,
    n45352, n45353, n45354, n45355, n45356, n45357,
    n45358, n45359, n45360, n45361, n45362, n45363,
    n45364, n45365, n45366, n45367, n45368, n45369,
    n45370, n45371, n45372, n45373, n45374, n45375,
    n45376, n45377, n45378, n45379, n45380, n45381,
    n45382, n45383, n45384, n45385, n45386, n45387,
    n45388, n45389, n45390, n45391, n45392, n45393,
    n45394, n45395, n45396, n45397, n45398, n45399,
    n45400, n45401, n45402, n45403, n45404, n45405,
    n45406, n45407, n45408, n45409, n45410, n45411,
    n45412, n45413, n45414, n45415, n45416, n45417,
    n45418, n45419, n45420, n45421, n45422, n45423,
    n45424, n45425, n45426, n45427, n45428, n45429,
    n45430, n45431, n45432, n45433, n45434, n45435,
    n45436, n45437, n45438, n45439, n45440, n45441,
    n45442, n45443, n45444, n45445, n45446, n45447,
    n45448, n45449, n45450, n45451, n45452, n45453,
    n45454, n45455, n45456, n45457, n45458, n45459,
    n45460, n45461, n45462, n45463, n45464, n45465,
    n45466, n45467, n45468, n45469, n45470, n45471,
    n45472, n45473, n45474, n45475, n45476, n45477,
    n45478, n45479, n45480, n45481, n45482, n45483,
    n45484, n45485, n45486, n45487, n45488, n45489,
    n45490, n45491, n45492, n45493, n45494, n45495,
    n45496, n45497, n45498, n45499, n45500, n45501,
    n45502, n45503, n45504, n45505, n45506, n45507,
    n45508, n45509, n45510, n45511, n45512, n45513,
    n45514, n45515, n45516, n45517, n45518, n45519,
    n45520, n45521, n45522, n45523, n45524, n45525,
    n45526, n45527, n45528, n45529, n45530, n45531,
    n45532, n45533, n45534, n45535, n45536, n45537,
    n45538, n45539, n45540, n45541, n45542, n45543,
    n45544, n45545, n45546, n45547, n45548, n45549,
    n45550, n45551, n45552, n45553, n45554, n45555,
    n45556, n45557, n45558, n45559, n45560, n45561,
    n45562, n45563, n45564, n45565, n45566, n45567,
    n45568, n45569, n45570, n45571, n45572, n45573,
    n45574, n45575, n45576, n45577, n45578, n45579,
    n45580, n45581, n45582, n45583, n45584, n45585,
    n45586, n45587, n45588, n45589, n45590, n45591,
    n45592, n45593, n45594, n45595, n45596, n45597,
    n45598, n45599, n45600, n45601, n45602, n45603,
    n45604, n45605, n45606, n45607, n45608, n45609,
    n45610, n45611, n45612, n45613, n45614, n45615,
    n45616, n45617, n45618, n45619, n45620, n45621,
    n45622, n45623, n45624, n45625, n45626, n45627,
    n45628, n45629, n45630, n45631, n45632, n45633,
    n45634, n45635, n45636, n45637, n45638, n45639,
    n45640, n45641, n45642, n45643, n45644, n45645,
    n45646, n45647, n45648, n45649, n45650, n45651,
    n45652, n45653, n45654, n45655, n45656, n45657,
    n45658, n45659, n45660, n45661, n45662, n45663,
    n45664, n45665, n45666, n45667, n45668, n45669,
    n45670, n45671, n45672, n45673, n45674, n45675,
    n45676, n45677, n45678, n45679, n45680, n45681,
    n45682, n45683, n45684, n45685, n45686, n45687,
    n45688, n45689, n45690, n45691, n45692, n45693,
    n45694, n45695, n45696, n45697, n45698, n45699,
    n45700, n45701, n45702, n45703, n45704, n45705,
    n45706, n45707, n45708, n45709, n45710, n45711,
    n45712, n45713, n45714, n45715, n45716, n45717,
    n45718, n45719, n45720, n45721, n45722, n45723,
    n45724, n45725, n45726, n45727, n45728, n45729,
    n45730, n45731, n45732, n45733, n45734, n45735,
    n45736, n45737, n45738, n45739, n45740, n45741,
    n45742, n45743, n45744, n45745, n45746, n45747,
    n45748, n45749, n45750, n45751, n45752, n45753,
    n45754, n45755, n45756, n45757, n45758, n45759,
    n45760, n45761, n45762, n45763, n45764, n45765,
    n45766, n45767, n45769, n45770, n45771, n45772,
    n45773, n45774, n45776, n45777, n45778, n45779,
    n45780, n45782, n45783, n45784, n45785, n45786,
    n45788, n45789, n45790, n45792, n45793, n45794,
    n45795, n45796, n45798, n45799, n45800, n45802,
    n45803, n45805, n45806, n45807, n45809, n45810,
    n45811, n45812, n45813, n45814, n45815, n45816,
    n45817, n45818, n45819, n45821, n45822, n45823,
    n45824, n45826, n45827, n45828, n45829, n45830,
    n45831, n45832, n45833, n45835, n45836, n45837,
    n45838, n45839, n45840, n45842, n45843, n45845,
    n45846, n45847, n45848, n45849, n45851, n45852,
    n45853, n45855, n45856, n45857, n45859, n45860,
    n45861, n45863, n45864, n45865, n45867, n45868,
    n45869, n45871, n45872, n45873, n45875, n45876,
    n45877, n45879, n45880, n45881, n45882, n45884,
    n45885, n45886, n45887, n45889, n45890, n45891,
    n45892, n45894, n45895, n45896, n45897, n45898,
    n45900, n45901, n45902, n45904, n45905, n45906,
    n45908, n45909, n45910, n45912, n45913, n45914,
    n45916, n45917, n45918, n45920, n45921, n45922,
    n45924, n45925, n45926, n45927, n45928, n45930,
    n45931, n45932, n45933, n45935, n45936, n45937,
    n45939, n45940, n45941, n45943, n45944, n45945,
    n45947, n45948, n45949, n45951, n45952, n45953,
    n45955, n45956, n45957, n45959, n45960, n45961,
    n45963, n45964, n45965, n45967, n45968, n45969,
    n45971, n45972, n45973, n45975, n45976, n45977,
    n45979, n45980, n45981, n45983, n45984, n45985,
    n45987, n45988, n45989, n45991, n45992, n45993,
    n45995, n45996, n45997, n45999, n46000, n46001,
    n46003, n46004, n46005, n46007, n46008, n46009,
    n46011, n46012, n46013, n46015, n46016, n46017,
    n46019, n46020, n46021, n46023, n46024, n46025,
    n46027, n46028, n46029, n46031, n46032, n46033,
    n46035, n46036, n46037, n46039, n46040, n46041,
    n46043, n46044, n46045, n46047, n46048, n46049,
    n46051, n46052, n46053, n46055, n46056, n46057,
    n46059, n46060, n46061, n46063, n46064, n46065,
    n46067, n46068, n46069, n46071, n46072, n46073,
    n46074, n46075, n46076, n46077, n46078, n46079,
    n46081, n46083, n46084, n46085, n46087, n46088,
    n46089, n46091, n46092, n46093, n46095, n46096,
    n46097, n46098, n46099, n46100, n46101, n46102,
    n46103, n46104, n46105, n46106, n46107, n46108,
    n46109, n46110, n46111, n46112, n46113, n46114,
    n46115, n46116, n46117, n46118, n46119, n46120,
    n46121, n46122, n46123, n46124, n46125, n46126,
    n46127, n46128, n46129, n46130, n46131, n46132,
    n46133, n46134, n46135, n46136, n46137, n46138,
    n46139, n46140, n46141, n46142, n46144, n46145,
    n46146, n46147, n46148, n46149, n46150, n46151,
    n46152, n46153, n46154, n46155, n46156, n46157,
    n46158, n46159, n46160, n46161, n46162, n46163,
    n46164, n46165, n46166, n46167, n46168, n46169,
    n46170, n46171, n46172, n46173, n46174, n46175,
    n46176, n46177, n46178, n46179, n46180, n46181,
    n46182, n46183, n46184, n46186, n46187, n46188,
    n46190, n46191, n46192, n46193, n46194, n46195,
    n46196, n46197, n46198, n46199, n46200, n46201,
    n46202, n46203, n46204, n46205, n46206, n46207,
    n46208, n46209, n46210, n46211, n46212, n46213,
    n46214, n46215, n46216, n46217, n46218, n46219,
    n46220, n46221, n46222, n46223, n46224, n46226,
    n46227, n46228, n46229, n46230, n46231, n46232,
    n46233, n46234, n46235, n46236, n46237, n46238,
    n46239, n46240, n46241, n46242, n46243, n46244,
    n46245, n46246, n46247, n46248, n46249, n46250,
    n46251, n46252, n46253, n46254, n46255, n46256,
    n46257, n46258, n46259, n46260, n46261, n46263,
    n46264, n46265, n46266, n46267, n46268, n46269,
    n46270, n46271, n46272, n46273, n46274, n46275,
    n46276, n46277, n46278, n46279, n46280, n46281,
    n46282, n46283, n46284, n46285, n46286, n46287,
    n46288, n46289, n46290, n46291, n46292, n46293,
    n46294, n46295, n46296, n46297, n46299, n46300,
    n46301, n46303, n46304, n46305, n46306, n46307,
    n46308, n46309, n46310, n46311, n46312, n46313,
    n46314, n46315, n46316, n46317, n46318, n46319,
    n46320, n46321, n46322, n46323, n46324, n46325,
    n46326, n46327, n46328, n46329, n46330, n46331,
    n46332, n46333, n46334, n46336, n46337, n46338,
    n46339, n46340, n46341, n46342, n46343, n46344,
    n46345, n46346, n46347, n46348, n46349, n46350,
    n46351, n46352, n46353, n46354, n46355, n46356,
    n46357, n46358, n46359, n46360, n46361, n46362,
    n46363, n46364, n46365, n46366, n46368, n46369,
    n46370, n46371, n46372, n46373, n46374, n46375,
    n46376, n46377, n46378, n46379, n46380, n46381,
    n46382, n46383, n46384, n46385, n46386, n46387,
    n46388, n46389, n46390, n46391, n46392, n46393,
    n46394, n46395, n46396, n46397, n46398, n46399,
    n46400, n46401, n46402, n46404, n46405, n46406,
    n46407, n46408, n46409, n46410, n46411, n46412,
    n46413, n46414, n46415, n46416, n46417, n46418,
    n46419, n46420, n46421, n46422, n46423, n46424,
    n46425, n46426, n46427, n46428, n46429, n46430,
    n46431, n46432, n46433, n46434, n46435, n46436,
    n46437, n46438, n46440, n46441, n46442, n46443,
    n46444, n46445, n46446, n46447, n46448, n46449,
    n46450, n46451, n46452, n46453, n46454, n46455,
    n46456, n46457, n46458, n46459, n46460, n46461,
    n46462, n46463, n46464, n46465, n46466, n46467,
    n46468, n46469, n46470, n46471, n46472, n46473,
    n46474, n46475, n46476, n46478, n46479, n46480,
    n46481, n46482, n46483, n46484, n46485, n46486,
    n46487, n46488, n46489, n46490, n46491, n46492,
    n46493, n46494, n46495, n46496, n46497, n46498,
    n46499, n46500, n46501, n46502, n46503, n46504,
    n46505, n46506, n46507, n46508, n46509, n46510,
    n46511, n46512, n46514, n46515, n46516, n46517,
    n46518, n46519, n46520, n46521, n46522, n46523,
    n46524, n46525, n46526, n46527, n46528, n46529,
    n46530, n46531, n46532, n46533, n46534, n46535,
    n46536, n46537, n46538, n46539, n46540, n46541,
    n46542, n46543, n46544, n46545, n46546, n46547,
    n46548, n46550, n46551, n46552, n46553, n46554,
    n46555, n46556, n46557, n46558, n46559, n46560,
    n46561, n46562, n46563, n46564, n46565, n46566,
    n46567, n46568, n46569, n46570, n46571, n46572,
    n46573, n46574, n46575, n46576, n46577, n46578,
    n46579, n46580, n46582, n46583, n46584, n46585,
    n46586, n46587, n46588, n46589, n46590, n46591,
    n46592, n46593, n46594, n46595, n46596, n46597,
    n46598, n46599, n46600, n46601, n46602, n46603,
    n46604, n46605, n46606, n46607, n46608, n46609,
    n46610, n46611, n46612, n46614, n46615, n46616,
    n46617, n46618, n46619, n46620, n46621, n46622,
    n46623, n46624, n46625, n46626, n46627, n46628,
    n46629, n46630, n46631, n46632, n46633, n46634,
    n46635, n46636, n46637, n46638, n46639, n46640,
    n46641, n46642, n46643, n46644, n46645, n46646,
    n46647, n46648, n46649, n46651, n46652, n46653,
    n46655, n46656, n46657, n46659, n46660, n46661,
    n46662, n46663, n46664, n46665, n46666, n46667,
    n46668, n46669, n46670, n46671, n46672, n46673,
    n46674, n46675, n46676, n46677, n46678, n46679,
    n46680, n46681, n46682, n46683, n46684, n46685,
    n46686, n46687, n46688, n46689, n46692, n46693,
    n46694, n46696, n46697, n46698, n46699, n46700,
    n46701, n46702, n46703, n46704, n46705, n46706,
    n46707, n46708, n46709, n46710, n46711, n46712,
    n46713, n46714, n46715, n46716, n46717, n46718,
    n46719, n46720, n46721, n46722, n46723, n46724,
    n46725, n46726, n46727, n46728, n46729, n46730,
    n46731, n46732, n46733, n46735, n46736, n46737,
    n46739, n46740, n46741, n46743, n46744, n46745,
    n46747, n46748, n46749, n46750, n46751, n46752,
    n46753, n46754, n46755, n46756, n46757, n46758,
    n46759, n46760, n46761, n46762, n46763, n46764,
    n46765, n46766, n46767, n46768, n46769, n46770,
    n46771, n46772, n46773, n46774, n46775, n46776,
    n46777, n46778, n46779, n46781, n46782, n46783,
    n46785, n46786, n46787, n46789, n46790, n46791,
    n46792, n46793, n46794, n46795, n46796, n46797,
    n46798, n46799, n46800, n46801, n46802, n46803,
    n46804, n46805, n46806, n46807, n46808, n46809,
    n46810, n46811, n46812, n46813, n46814, n46815,
    n46816, n46817, n46818, n46819, n46820, n46821,
    n46822, n46824, n46825, n46826, n46828, n46829,
    n46830, n46832, n46833, n46834, n46836, n46837,
    n46838, n46840, n46841, n46842, n46844, n46845,
    n46846, n46848, n46849, n46850, n46852, n46853,
    n46854, n46856, n46857, n46858, n46860, n46861,
    n46862, n46864, n46865, n46866, n46868, n46869,
    n46870, n46872, n46873, n46874, n46876, n46877,
    n46878, n46880, n46881, n46882, n46883, n46884,
    n46885, n46886, n46887, n46888, n46889, n46890,
    n46891, n46892, n46893, n46894, n46895, n46896,
    n46897, n46898, n46899, n46900, n46901, n46902,
    n46903, n46904, n46905, n46906, n46907, n46908,
    n46909, n46910, n46911, n46912, n46913, n46914,
    n46916, n46917, n46918, n46919, n46920, n46921,
    n46922, n46923, n46924, n46925, n46926, n46927,
    n46928, n46929, n46930, n46931, n46932, n46933,
    n46934, n46935, n46936, n46937, n46938, n46939,
    n46940, n46941, n46942, n46943, n46944, n46945,
    n46946, n46947, n46948, n46949, n46950, n46951,
    n46952, n46953, n46954, n46956, n46957, n46958,
    n46960, n46961, n46962, n46964, n46965, n46966,
    n46967, n46968, n46969, n46970, n46971, n46972,
    n46973, n46974, n46975, n46976, n46977, n46978,
    n46979, n46980, n46981, n46982, n46983, n46984,
    n46985, n46986, n46987, n46988, n46989, n46990,
    n46991, n46992, n46993, n46994, n46995, n46996,
    n46998, n46999, n47000, n47001, n47002, n47003,
    n47004, n47005, n47006, n47007, n47008, n47009,
    n47010, n47011, n47012, n47013, n47014, n47015,
    n47016, n47017, n47018, n47019, n47020, n47021,
    n47022, n47023, n47024, n47025, n47026, n47027,
    n47028, n47029, n47030, n47031, n47033, n47034,
    n47035, n47036, n47037, n47038, n47039, n47040,
    n47041, n47042, n47043, n47044, n47045, n47046,
    n47047, n47048, n47049, n47050, n47051, n47052,
    n47053, n47054, n47055, n47056, n47057, n47058,
    n47059, n47060, n47061, n47062, n47063, n47064,
    n47065, n47067, n47068, n47069, n47070, n47071,
    n47072, n47073, n47074, n47075, n47076, n47077,
    n47078, n47079, n47080, n47081, n47082, n47083,
    n47084, n47085, n47086, n47087, n47088, n47089,
    n47090, n47091, n47092, n47093, n47094, n47095,
    n47096, n47097, n47098, n47099, n47100, n47102,
    n47103, n47104, n47106, n47107, n47108, n47109,
    n47110, n47111, n47112, n47113, n47114, n47115,
    n47116, n47117, n47118, n47119, n47120, n47121,
    n47122, n47123, n47124, n47125, n47126, n47127,
    n47128, n47129, n47130, n47131, n47132, n47133,
    n47134, n47135, n47136, n47137, n47138, n47139,
    n47140, n47142, n47143, n47144, n47145, n47146,
    n47147, n47148, n47149, n47150, n47151, n47152,
    n47153, n47154, n47155, n47156, n47157, n47158,
    n47159, n47160, n47161, n47162, n47163, n47164,
    n47165, n47166, n47167, n47168, n47169, n47170,
    n47171, n47172, n47173, n47174, n47176, n47177,
    n47178, n47179, n47180, n47181, n47182, n47183,
    n47184, n47185, n47186, n47187, n47188, n47189,
    n47190, n47191, n47192, n47193, n47194, n47195,
    n47196, n47197, n47198, n47199, n47200, n47201,
    n47202, n47203, n47204, n47205, n47206, n47207,
    n47208, n47209, n47210, n47212, n47213, n47214,
    n47215, n47216, n47217, n47218, n47219, n47220,
    n47221, n47222, n47223, n47224, n47225, n47226,
    n47227, n47228, n47229, n47230, n47231, n47232,
    n47233, n47234, n47235, n47236, n47237, n47238,
    n47239, n47240, n47241, n47242, n47243, n47244,
    n47246, n47247, n47248, n47249, n47250, n47251,
    n47252, n47253, n47254, n47255, n47256, n47257,
    n47258, n47259, n47260, n47261, n47262, n47263,
    n47264, n47265, n47266, n47267, n47268, n47269,
    n47270, n47271, n47272, n47273, n47274, n47275,
    n47276, n47277, n47278, n47279, n47281, n47282,
    n47283, n47284, n47285, n47286, n47287, n47288,
    n47289, n47290, n47291, n47292, n47293, n47294,
    n47295, n47296, n47297, n47298, n47299, n47300,
    n47301, n47302, n47303, n47304, n47305, n47306,
    n47307, n47308, n47309, n47310, n47311, n47312,
    n47313, n47314, n47315, n47316, n47317, n47318,
    n47319, n47320, n47321, n47322, n47323, n47324,
    n47325, n47326, n47327, n47328, n47329, n47330,
    n47331, n47332, n47333, n47334, n47335, n47337,
    n47338, n47340, n47341, n47342, n47343, n47344,
    n47345, n47346, n47347, n47348, n47349, n47350,
    n47351, n47352, n47353, n47354, n47355, n47356,
    n47357, n47358, n47359, n47360, n47361, n47362,
    n47363, n47364, n47365, n47366, n47367, n47368,
    n47369, n47370, n47371, n47372, n47373, n47375,
    n47376, n47377, n47379, n47380, n47381, n47383,
    n47384, n47385, n47387, n47388, n47389, n47391,
    n47392, n47393, n47395, n47396, n47397, n47399,
    n47400, n47401, n47403, n47404, n47405, n47407,
    n47408, n47409, n47410, n47411, n47412, n47413,
    n47414, n47415, n47416, n47417, n47418, n47419,
    n47420, n47422, n47423, n47424, n47426, n47427,
    n47428, n47429, n47430, n47431, n47432, n47433,
    n47434, n47435, n47436, n47437, n47438, n47439,
    n47440, n47441, n47442, n47443, n47444, n47445,
    n47446, n47447, n47448, n47449, n47450, n47451,
    n47452, n47453, n47454, n47455, n47456, n47457,
    n47458, n47459, n47460, n47462, n47463, n47464,
    n47466, n47467, n47468, n47470, n47471, n47472,
    n47474, n47475, n47476, n47478, n47479, n47480,
    n47482, n47483, n47485, n47486, n47487, n47489,
    n47490, n47491, n47493, n47494, n47495, n47497,
    n47498, n47499, n47501, n47502, n47503, n47505,
    n47506, n47507, n47509, n47510, n47511, n47513,
    n47514, n47515, n47516, n47517, n47518, n47519,
    n47520, n47521, n47522, n47523, n47525, n47526,
    n47527, n47529, n47530, n47531, n47533, n47534,
    n47535, n47537, n47538, n47539, n47541, n47542,
    n47543, n47545, n47546, n47547, n47549, n47550,
    n47551, n47553, n47554, n47555, n47557, n47558,
    n47559, n47561, n47562, n47563, n47565, n47566,
    n47567, n47569, n47570, n47571, n47573, n47574,
    n47575, n47577, n47578, n47579, n47581, n47582,
    n47583, n47585, n47586, n47587, n47589, n47590,
    n47591, n47593, n47594, n47595, n47596, n47597,
    n47598, n47599, n47600, n47601, n47602, n47603,
    n47604, n47605, n47606, n47608, n47609, n47611,
    n47612, n47613, n47615, n47616, n47617, n47619,
    n47620, n47621, n47623, n47624, n47625, n47626,
    n47627, n47628, n47629, n47630, n47631, n47632,
    n47633, n47634, n47635, n47636, n47637, n47638,
    n47640, n47641, n47642, n47644, n47645, n47646,
    n47647, n47649, n47650, n47651, n47653, n47654,
    n47655, n47656, n47657, n47659, n47660, n47661,
    n47663, n47664, n47665, n47666, n47667, n47668,
    n47669, n47670, n47671, n47672, n47673, n47674,
    n47675, n47676, n47677, n47678, n47680, n47681,
    n47682, n47684, n47685, n47686, n47688, n47689,
    n47690, n47691, n47692, n47693, n47694, n47698,
    n47699, n47701, n47703, n47704, n47706, n47707,
    n47709, n47710, n47712, n47713, n47715, n47716,
    n47718, n47719, n47721, n47722, n47724, n47725,
    n47727, n47728, n47730, n47731, n47733, n47734,
    n47735, n47737, n47738, n47740, n47741, n47742,
    n47743, n47744, n47745, n47746, n47747, n47749,
    n47750, n47752, n47753, n47755, n47756, n47758,
    n47759, n47761, n47762, n47764, n47765, n47767,
    n47768, n47769, n47771, n47772, n47774, n47775,
    n47777, n47778, n47780, n47781, n47783, n47784,
    n47786, n47787, n47789, n47790, n47792, n47793,
    n47795, n47796, n47798, n47799, n47801, n47803,
    n47805, n47807, n47810, n47811, n47812, n47814,
    n47815, n47816, n47817, n47818, n47819, n47820,
    n47821, n47822, n47823, n47824, n47825, n47826,
    n47827, n47828, n47829, n47830, n47831, n47832,
    n47833, n47834, n47835, n47836, n47837, n47838,
    n47839, n47840, n47841, n47843, n47844, n47845,
    n47846, n47847, n47848, n47849, n47850, n47851,
    n47852, n47853, n47854, n47855, n47856, n47857,
    n47858, n47859, n47860, n47861, n47862, n47863,
    n47864, n47865, n47866, n47867, n47868, n47869,
    n47871, n47872, n47873, n47874, n47875, n47876,
    n47877, n47878, n47879, n47880, n47881, n47882,
    n47883, n47884, n47885, n47886, n47887, n47888,
    n47889, n47890, n47891, n47892, n47893, n47894,
    n47895, n47896, n47897, n47899, n47900, n47901,
    n47902, n47903, n47904, n47905, n47906, n47907,
    n47908, n47909, n47910, n47911, n47912, n47913,
    n47914, n47915, n47916, n47917, n47918, n47919,
    n47920, n47921, n47922, n47923, n47924, n47925,
    n47927, n47928, n47930, n47932, n47933, n47935,
    n47938, n47940, n47941, n47943, n47944, n47946,
    n47947, n47949, n47950, n47953, n47954, n47956,
    n47957, n47959, n47960, n47962, n47963, n47965,
    n47966, n47968, n47969, n47971, n47972, n47974,
    n47975, n47977, n47978, n47980, n47981, n47983,
    n47984, n47986, n47987, n47989, n47990, n47992,
    n47993, n47995, n47996, n47998, n47999, n48001,
    n48002, n48004, n48005, n48007, n48008, n48010,
    n48011, n48012, n48013, n48014, n48015, n48016,
    n48017, n48019, n48020, n48022, n48023, n48025,
    n48026, n48028, n48029, n48031, n48032, n48034,
    n48035, n48037, n48038, n48040, n48041, n48042,
    n48043, n48044, n48045, n48046, n48047, n48049,
    n48050, n48052, n48053, n48055, n48056, n48058,
    n48059, n48061, n48062, n48064, n48065, n48066,
    n48067, n48068, n48069, n48070, n48071, n48073,
    n48074, n48076, n48077, n48078, n48079, n48080,
    n48081, n48082, n48083, n48085, n48086, n48087,
    n48088, n48089, n48090, n48091, n48092, n48094,
    n48095, n48096, n48097, n48098, n48099, n48100,
    n48101, n48103, n48104, n48106, n48107, n48109,
    n48111, n48112, n48114, n48115, n48117, n48118,
    n48120, n48122, n48123, n48125, n48126, n48128,
    n48129, n48131, n48132, n48134, n48135, n48137,
    n48138, n48140, n48141, n48143, n48144, n48146,
    n48147, n48149, n48151, n48152, n48154, n48155,
    n48157, n48158, n48160, n48162, n48164, n48165,
    n48167, n48168, n48169, n48170, n48171, n48172,
    n48173, n48174, n48175, n48176, n48178, n48180,
    n48181, n48183, n48184, n48186, n48187, n48189,
    n48191, n48192, n48194, n48196, n48197, n48199,
    n48201, n48202, n48204, n48205, n48207, n48208,
    n48210, n48211, n48213, n48215, n48216, n48218,
    n48219, n48221, n48222, n48224, n48225, n48227,
    n48228, n48230, n48231, n48233, n48235, n48236,
    n48238, n48239, n48241, n48242, n48244, n48246,
    n48248, n48249, n48251, n48253, n48254, n48256,
    n48257, n48259, n48261, n48262, n48264, n48266,
    n48267, n48269, n48270, n48272, n48273, n48275,
    n48276, n48279, n48281, n48283, n48284, n48287;
  assign n2437 = ~pi216 & pi833;
  assign n2438 = pi929 & n2437;
  assign n2439 = pi1144 & ~n2437;
  assign n2440 = ~pi332 & ~n2439;
  assign n2441 = ~n2438 & n2440;
  assign n2442 = pi221 & ~n2441;
  assign n2443 = pi265 & ~pi332;
  assign n2444 = pi216 & ~n2443;
  assign n2445 = pi153 & ~pi332;
  assign n2446 = ~pi105 & ~n2445;
  assign n2447 = ~pi152 & ~pi161;
  assign n2448 = ~pi166 & n2447;
  assign n2449 = pi95 & ~pi479;
  assign n2450 = ~pi40 & ~pi72;
  assign n2451 = ~pi88 & ~pi98;
  assign n2452 = ~pi77 & n2451;
  assign n2453 = ~pi50 & n2452;
  assign n2454 = ~pi102 & n2453;
  assign n2455 = ~pi65 & ~pi71;
  assign n2456 = ~pi83 & ~pi103;
  assign n2457 = ~pi67 & ~pi69;
  assign n2458 = ~pi66 & ~pi73;
  assign n2459 = ~pi61 & ~pi76;
  assign n2460 = ~pi85 & ~pi106;
  assign n2461 = n2459 & n2460;
  assign n2462 = ~pi48 & n2461;
  assign n2463 = ~pi89 & n2462;
  assign n2464 = ~pi49 & n2463;
  assign n2465 = ~pi104 & n2464;
  assign n2466 = ~pi45 & n2465;
  assign n2467 = ~pi68 & ~pi84;
  assign n2468 = ~pi82 & ~pi111;
  assign n2469 = ~pi36 & n2468;
  assign n2470 = n2467 & n2469;
  assign n2471 = n2466 & n2470;
  assign n2472 = n2458 & n2471;
  assign n2473 = n2457 & n2472;
  assign n2474 = n2456 & n2473;
  assign n2475 = n2455 & n2474;
  assign n2476 = ~pi63 & ~pi107;
  assign n2477 = n2475 & n2476;
  assign n2478 = ~pi64 & n2477;
  assign n2479 = ~pi81 & n2478;
  assign n2480 = n2454 & n2479;
  assign n2481 = ~pi97 & ~pi108;
  assign n2482 = ~pi94 & n2481;
  assign n2483 = ~pi53 & ~pi60;
  assign n2484 = ~pi86 & n2483;
  assign n2485 = ~pi46 & n2484;
  assign n2486 = n2482 & n2485;
  assign n2487 = n2480 & n2486;
  assign n2488 = ~pi109 & ~pi110;
  assign n2489 = ~pi58 & ~pi91;
  assign n2490 = ~pi47 & n2489;
  assign n2491 = n2488 & n2490;
  assign n2492 = n2487 & n2491;
  assign n2493 = ~pi90 & ~pi93;
  assign n2494 = ~pi70 & ~pi96;
  assign n2495 = ~pi35 & ~pi51;
  assign n2496 = n2494 & n2495;
  assign n2497 = n2493 & n2496;
  assign n2498 = n2492 & n2497;
  assign n2499 = n2450 & n2498;
  assign n2500 = pi225 & n2499;
  assign n2501 = pi32 & ~n2500;
  assign n2502 = ~pi95 & ~n2501;
  assign n2503 = pi60 & n2480;
  assign n2504 = ~pi53 & ~n2503;
  assign n2505 = ~pi86 & ~pi94;
  assign n2506 = ~pi60 & n2480;
  assign n2507 = pi53 & ~n2506;
  assign n2508 = n2505 & ~n2507;
  assign n2509 = ~n2504 & n2508;
  assign n2510 = ~pi46 & n2488;
  assign n2511 = ~pi47 & ~pi91;
  assign n2512 = n2481 & n2511;
  assign n2513 = n2510 & n2512;
  assign n2514 = ~pi58 & n2513;
  assign n2515 = n2493 & n2514;
  assign n2516 = n2509 & n2515;
  assign n2517 = ~pi35 & ~n2516;
  assign n2518 = ~pi58 & ~pi90;
  assign n2519 = n2486 & n2488;
  assign n2520 = n2511 & n2519;
  assign n2521 = n2480 & n2520;
  assign n2522 = n2518 & n2521;
  assign n2523 = ~pi93 & n2522;
  assign n2524 = pi35 & ~n2523;
  assign n2525 = pi35 & n2523;
  assign n2526 = ~pi225 & n2525;
  assign n2527 = ~pi70 & ~n2526;
  assign n2528 = ~pi51 & n2527;
  assign n2529 = ~n2524 & n2528;
  assign n2530 = ~n2517 & n2529;
  assign n2531 = ~pi96 & ~n2530;
  assign n2532 = ~pi47 & n2519;
  assign n2533 = n2480 & n2532;
  assign n2534 = ~pi35 & ~pi70;
  assign n2535 = ~pi51 & n2534;
  assign n2536 = ~pi93 & n2518;
  assign n2537 = ~pi91 & n2536;
  assign n2538 = n2535 & n2537;
  assign n2539 = n2533 & n2538;
  assign n2540 = pi96 & ~n2539;
  assign n2541 = n2450 & ~n2540;
  assign n2542 = ~n2531 & n2541;
  assign n2543 = ~pi32 & ~n2542;
  assign n2544 = n2502 & ~n2543;
  assign n2545 = ~n2449 & ~n2544;
  assign n2546 = ~pi137 & n2545;
  assign n2547 = ~pi35 & ~pi93;
  assign n2548 = n2522 & n2547;
  assign n2549 = ~pi72 & ~pi96;
  assign n2550 = ~pi51 & ~pi70;
  assign n2551 = n2549 & n2550;
  assign n2552 = n2548 & n2551;
  assign n2553 = pi40 & n2552;
  assign n2554 = ~pi32 & ~n2553;
  assign n2555 = pi72 & ~n2498;
  assign n2556 = ~pi40 & ~n2555;
  assign n2557 = ~pi70 & n2548;
  assign n2558 = pi51 & ~n2557;
  assign n2559 = ~pi96 & ~n2558;
  assign n2560 = ~pi51 & pi70;
  assign n2561 = n2559 & ~n2560;
  assign n2562 = ~n2524 & ~n2526;
  assign n2563 = pi93 & n2522;
  assign n2564 = ~pi35 & ~n2563;
  assign n2565 = pi91 & n2533;
  assign n2566 = n2518 & ~n2565;
  assign n2567 = ~pi109 & n2487;
  assign n2568 = pi110 & ~n2567;
  assign n2569 = pi47 & n2480;
  assign n2570 = n2519 & n2569;
  assign n2571 = pi47 & ~n2570;
  assign n2572 = ~pi91 & ~n2571;
  assign n2573 = ~n2568 & n2572;
  assign n2574 = ~pi47 & ~pi110;
  assign n2575 = pi109 & ~n2487;
  assign n2576 = ~pi102 & n2479;
  assign n2577 = n2451 & n2576;
  assign n2578 = ~pi50 & n2483;
  assign n2579 = ~pi77 & n2578;
  assign n2580 = n2505 & n2579;
  assign n2581 = n2577 & n2580;
  assign n2582 = ~pi97 & n2581;
  assign n2583 = pi108 & ~n2582;
  assign n2584 = ~pi46 & ~n2583;
  assign n2585 = pi97 & ~n2581;
  assign n2586 = n2452 & n2576;
  assign n2587 = n2578 & n2586;
  assign n2588 = ~pi86 & pi94;
  assign n2589 = n2587 & n2588;
  assign n2590 = ~pi97 & ~n2589;
  assign n2591 = pi86 & ~n2587;
  assign n2592 = ~pi94 & ~n2591;
  assign n2593 = pi77 & n2577;
  assign n2594 = ~pi50 & ~n2593;
  assign n2595 = pi81 & ~n2478;
  assign n2596 = pi102 & ~n2479;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = pi64 & ~n2477;
  assign n2599 = pi71 & ~n2474;
  assign n2600 = ~pi65 & ~n2599;
  assign n2601 = ~pi67 & n2472;
  assign n2602 = pi69 & ~n2601;
  assign n2603 = pi83 & ~n2473;
  assign n2604 = ~pi103 & ~n2603;
  assign n2605 = ~n2602 & n2604;
  assign n2606 = ~pi69 & ~pi83;
  assign n2607 = ~pi68 & ~pi111;
  assign n2608 = n2458 & n2466;
  assign n2609 = pi84 & ~n2608;
  assign n2610 = pi85 & pi106;
  assign n2611 = n2459 & ~n2610;
  assign n2612 = pi61 & pi76;
  assign n2613 = n2460 & ~n2612;
  assign n2614 = ~n2611 & ~n2613;
  assign n2615 = ~pi48 & ~n2614;
  assign n2616 = ~n2461 & ~n2615;
  assign n2617 = pi89 & ~n2462;
  assign n2618 = ~pi49 & ~n2617;
  assign n2619 = ~n2616 & n2618;
  assign n2620 = ~n2463 & ~n2619;
  assign n2621 = pi104 & ~n2464;
  assign n2622 = ~pi45 & ~n2621;
  assign n2623 = ~n2620 & n2622;
  assign n2624 = ~n2465 & ~n2623;
  assign n2625 = ~n2466 & ~n2624;
  assign n2626 = n2458 & ~n2625;
  assign n2627 = pi66 & pi73;
  assign n2628 = ~n2458 & ~n2466;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = ~n2626 & n2629;
  assign n2631 = ~pi84 & ~n2630;
  assign n2632 = ~n2609 & ~n2631;
  assign n2633 = n2607 & ~n2632;
  assign n2634 = ~pi84 & n2608;
  assign n2635 = ~pi68 & n2634;
  assign n2636 = pi111 & ~n2635;
  assign n2637 = ~pi82 & ~n2636;
  assign n2638 = pi68 & ~n2634;
  assign n2639 = n2637 & ~n2638;
  assign n2640 = ~n2633 & n2639;
  assign n2641 = ~pi36 & ~pi67;
  assign n2642 = pi82 & n2607;
  assign n2643 = n2634 & n2642;
  assign n2644 = n2641 & ~n2643;
  assign n2645 = ~n2640 & n2644;
  assign n2646 = pi67 & ~n2472;
  assign n2647 = n2468 & n2635;
  assign n2648 = pi36 & ~n2647;
  assign n2649 = ~n2646 & ~n2648;
  assign n2650 = ~n2645 & n2649;
  assign n2651 = n2606 & ~n2650;
  assign n2652 = n2605 & ~n2651;
  assign n2653 = pi103 & n2606;
  assign n2654 = n2601 & n2653;
  assign n2655 = ~pi71 & ~n2654;
  assign n2656 = ~n2652 & n2655;
  assign n2657 = n2600 & ~n2656;
  assign n2658 = ~pi107 & ~n2657;
  assign n2659 = pi65 & ~pi71;
  assign n2660 = n2474 & n2659;
  assign n2661 = n2658 & ~n2660;
  assign n2662 = ~pi63 & pi107;
  assign n2663 = n2475 & n2662;
  assign n2664 = ~n2476 & ~n2663;
  assign n2665 = ~n2661 & ~n2664;
  assign n2666 = ~pi64 & ~n2665;
  assign n2667 = ~n2598 & ~n2666;
  assign n2668 = ~pi81 & ~pi102;
  assign n2669 = ~n2667 & n2668;
  assign n2670 = ~n2658 & ~n2664;
  assign n2671 = pi63 & ~pi107;
  assign n2672 = n2475 & n2671;
  assign n2673 = ~pi64 & ~n2672;
  assign n2674 = ~n2670 & n2673;
  assign n2675 = ~n2598 & ~n2674;
  assign n2676 = n2669 & ~n2675;
  assign n2677 = n2597 & ~n2676;
  assign n2678 = n2451 & ~n2677;
  assign n2679 = ~pi98 & n2576;
  assign n2680 = pi88 & ~n2679;
  assign n2681 = pi98 & ~n2576;
  assign n2682 = ~pi77 & ~n2681;
  assign n2683 = ~n2680 & n2682;
  assign n2684 = ~n2678 & n2683;
  assign n2685 = n2594 & ~n2684;
  assign n2686 = pi50 & ~n2586;
  assign n2687 = ~pi60 & ~n2686;
  assign n2688 = ~n2685 & n2687;
  assign n2689 = n2504 & ~n2688;
  assign n2690 = ~n2507 & ~n2689;
  assign n2691 = ~pi86 & ~n2690;
  assign n2692 = n2592 & ~n2691;
  assign n2693 = n2590 & ~n2692;
  assign n2694 = ~n2585 & ~n2693;
  assign n2695 = ~pi108 & ~n2694;
  assign n2696 = n2584 & ~n2695;
  assign n2697 = pi46 & n2481;
  assign n2698 = n2581 & n2697;
  assign n2699 = ~pi109 & ~n2698;
  assign n2700 = ~n2696 & n2699;
  assign n2701 = ~n2575 & ~n2700;
  assign n2702 = n2574 & ~n2701;
  assign n2703 = n2573 & ~n2702;
  assign n2704 = n2566 & ~n2703;
  assign n2705 = pi58 & ~n2521;
  assign n2706 = pi90 & ~n2492;
  assign n2707 = ~pi93 & ~n2706;
  assign n2708 = ~n2705 & n2707;
  assign n2709 = ~n2704 & n2708;
  assign n2710 = n2564 & ~n2709;
  assign n2711 = n2562 & ~n2710;
  assign n2712 = ~pi51 & ~n2711;
  assign n2713 = n2561 & ~n2712;
  assign n2714 = ~pi72 & ~n2713;
  assign n2715 = n2556 & ~n2714;
  assign n2716 = n2554 & ~n2715;
  assign n2717 = pi96 & n2539;
  assign n2718 = ~pi51 & ~pi72;
  assign n2719 = ~pi40 & n2718;
  assign n2720 = n2548 & n2719;
  assign n2721 = n2717 & n2720;
  assign n2722 = n2716 & ~n2721;
  assign n2723 = ~n2501 & ~n2722;
  assign n2724 = ~pi95 & ~n2723;
  assign n2725 = ~pi32 & ~pi40;
  assign n2726 = n2552 & n2725;
  assign n2727 = pi95 & ~n2726;
  assign n2728 = pi479 & n2727;
  assign n2729 = ~n2724 & ~n2728;
  assign n2730 = pi137 & ~n2729;
  assign n2731 = ~n2546 & ~n2730;
  assign n2732 = pi210 & ~n2731;
  assign n2733 = ~pi833 & pi957;
  assign n2734 = pi1091 & ~n2733;
  assign n2735 = pi841 & n2522;
  assign n2736 = ~pi93 & n2735;
  assign n2737 = n2718 & n2736;
  assign n2738 = ~pi35 & ~pi40;
  assign n2739 = pi225 & n2738;
  assign n2740 = n2494 & n2739;
  assign n2741 = n2737 & n2740;
  assign n2742 = pi32 & ~n2741;
  assign n2743 = ~n2722 & ~n2742;
  assign n2744 = ~pi95 & ~n2743;
  assign n2745 = ~n2728 & ~n2744;
  assign n2746 = pi137 & ~n2745;
  assign n2747 = ~pi95 & ~n2742;
  assign n2748 = ~n2543 & n2747;
  assign n2749 = ~n2449 & ~n2748;
  assign n2750 = ~pi137 & n2749;
  assign n2751 = ~n2746 & ~n2750;
  assign n2752 = ~n2734 & n2751;
  assign n2753 = pi829 & pi950;
  assign n2754 = pi1092 & pi1093;
  assign n2755 = n2753 & n2754;
  assign n2756 = ~n2749 & ~n2755;
  assign n2757 = ~pi97 & ~n2509;
  assign n2758 = ~pi108 & ~n2585;
  assign n2759 = ~pi110 & n2758;
  assign n2760 = ~pi46 & ~pi109;
  assign n2761 = n2511 & n2760;
  assign n2762 = n2536 & n2761;
  assign n2763 = n2759 & n2762;
  assign n2764 = ~n2757 & n2763;
  assign n2765 = ~pi35 & ~n2764;
  assign n2766 = n2529 & ~n2765;
  assign n2767 = ~pi96 & ~n2766;
  assign n2768 = n2541 & ~n2767;
  assign n2769 = ~pi32 & ~n2768;
  assign n2770 = ~n2742 & ~n2769;
  assign n2771 = ~pi95 & ~n2770;
  assign n2772 = pi95 & pi479;
  assign n2773 = n2755 & ~n2772;
  assign n2774 = ~n2771 & n2773;
  assign n2775 = ~pi137 & ~n2774;
  assign n2776 = ~n2756 & n2775;
  assign n2777 = n2734 & ~n2776;
  assign n2778 = ~n2746 & n2777;
  assign n2779 = ~n2752 & ~n2778;
  assign n2780 = ~pi210 & n2779;
  assign n2781 = ~n2732 & ~n2780;
  assign n2782 = pi234 & n2781;
  assign n2783 = ~pi40 & n2549;
  assign n2784 = n2530 & n2783;
  assign n2785 = ~pi32 & ~n2784;
  assign n2786 = n2502 & ~n2785;
  assign n2787 = ~pi137 & ~n2786;
  assign n2788 = ~n2449 & ~n2727;
  assign n2789 = ~n2501 & ~n2716;
  assign n2790 = ~pi95 & ~n2789;
  assign n2791 = n2788 & ~n2790;
  assign n2792 = pi137 & ~n2791;
  assign n2793 = ~n2787 & ~n2792;
  assign n2794 = pi210 & ~n2793;
  assign n2795 = n2734 & n2755;
  assign n2796 = ~n2517 & ~n2795;
  assign n2797 = ~n2765 & n2795;
  assign n2798 = ~n2796 & ~n2797;
  assign n2799 = n2529 & n2783;
  assign n2800 = ~n2798 & n2799;
  assign n2801 = ~pi32 & ~n2800;
  assign n2802 = n2747 & ~n2801;
  assign n2803 = ~pi137 & ~n2802;
  assign n2804 = ~n2716 & ~n2742;
  assign n2805 = ~pi95 & ~n2804;
  assign n2806 = n2788 & ~n2805;
  assign n2807 = pi137 & ~n2806;
  assign n2808 = ~n2803 & ~n2807;
  assign n2809 = ~pi210 & ~n2808;
  assign n2810 = ~n2794 & ~n2809;
  assign n2811 = ~pi234 & n2810;
  assign n2812 = ~pi332 & ~n2811;
  assign n2813 = ~n2782 & n2812;
  assign n2814 = n2448 & ~n2813;
  assign n2815 = pi146 & n2781;
  assign n2816 = pi234 & ~pi332;
  assign n2817 = ~pi210 & ~n2751;
  assign n2818 = ~pi146 & ~n2732;
  assign n2819 = ~n2817 & n2818;
  assign n2820 = n2816 & ~n2819;
  assign n2821 = ~n2815 & n2820;
  assign n2822 = n2747 & ~n2785;
  assign n2823 = ~pi137 & ~n2822;
  assign n2824 = ~n2807 & ~n2823;
  assign n2825 = ~pi210 & ~n2824;
  assign n2826 = ~pi146 & ~n2794;
  assign n2827 = ~n2825 & n2826;
  assign n2828 = ~pi234 & ~pi332;
  assign n2829 = pi146 & n2810;
  assign n2830 = n2828 & ~n2829;
  assign n2831 = ~n2827 & n2830;
  assign n2832 = ~n2448 & ~n2831;
  assign n2833 = ~n2821 & n2832;
  assign n2834 = ~n2814 & ~n2833;
  assign n2835 = pi105 & ~n2834;
  assign n2836 = ~n2446 & ~n2835;
  assign n2837 = pi228 & ~n2836;
  assign n2838 = pi225 & pi841;
  assign n2839 = n2499 & ~n2838;
  assign n2840 = pi32 & ~n2839;
  assign n2841 = ~pi95 & ~n2840;
  assign n2842 = ~pi51 & ~pi96;
  assign n2843 = pi70 & ~n2548;
  assign n2844 = n2842 & ~n2843;
  assign n2845 = n2450 & n2844;
  assign n2846 = ~n2527 & n2845;
  assign n2847 = ~pi32 & ~n2846;
  assign n2848 = n2841 & ~n2847;
  assign n2849 = pi137 & ~n2848;
  assign n2850 = pi93 & ~n2522;
  assign n2851 = ~pi35 & ~n2850;
  assign n2852 = ~n2705 & ~n2706;
  assign n2853 = ~pi53 & n2688;
  assign n2854 = ~pi86 & ~n2853;
  assign n2855 = n2592 & ~n2854;
  assign n2856 = n2590 & ~n2855;
  assign n2857 = ~n2585 & ~n2856;
  assign n2858 = ~pi108 & ~n2857;
  assign n2859 = n2584 & ~n2858;
  assign n2860 = ~pi109 & ~n2859;
  assign n2861 = ~n2575 & ~n2860;
  assign n2862 = n2574 & ~n2861;
  assign n2863 = n2573 & ~n2862;
  assign n2864 = n2566 & ~n2863;
  assign n2865 = n2852 & ~n2864;
  assign n2866 = ~pi93 & ~n2865;
  assign n2867 = n2851 & ~n2866;
  assign n2868 = n2528 & ~n2867;
  assign n2869 = n2559 & ~n2843;
  assign n2870 = ~n2868 & n2869;
  assign n2871 = ~pi72 & ~n2870;
  assign n2872 = n2556 & ~n2871;
  assign n2873 = n2554 & ~n2872;
  assign n2874 = ~n2795 & n2873;
  assign n2875 = n2554 & n2795;
  assign n2876 = ~pi97 & ~n2856;
  assign n2877 = ~pi108 & ~n2876;
  assign n2878 = n2584 & ~n2877;
  assign n2879 = ~pi109 & ~n2878;
  assign n2880 = ~n2575 & ~n2879;
  assign n2881 = n2574 & ~n2880;
  assign n2882 = n2573 & ~n2881;
  assign n2883 = n2566 & ~n2882;
  assign n2884 = n2852 & ~n2883;
  assign n2885 = ~pi93 & ~n2884;
  assign n2886 = n2851 & ~n2885;
  assign n2887 = n2528 & ~n2886;
  assign n2888 = n2869 & ~n2887;
  assign n2889 = ~pi72 & ~n2888;
  assign n2890 = n2556 & ~n2889;
  assign n2891 = n2875 & ~n2890;
  assign n2892 = ~n2840 & ~n2891;
  assign n2893 = ~n2874 & n2892;
  assign n2894 = ~pi95 & ~n2893;
  assign n2895 = n2788 & ~n2894;
  assign n2896 = ~pi137 & ~n2895;
  assign n2897 = ~n2849 & ~n2896;
  assign n2898 = ~pi210 & ~n2897;
  assign n2899 = pi146 & n2898;
  assign n2900 = ~pi225 & n2499;
  assign n2901 = pi32 & ~n2900;
  assign n2902 = ~n2873 & ~n2901;
  assign n2903 = ~pi95 & ~n2902;
  assign n2904 = ~pi137 & n2788;
  assign n2905 = ~n2903 & n2904;
  assign n2906 = ~pi95 & ~n2901;
  assign n2907 = pi137 & n2906;
  assign n2908 = ~n2847 & n2907;
  assign n2909 = pi210 & ~n2908;
  assign n2910 = ~n2905 & n2909;
  assign n2911 = n2816 & ~n2910;
  assign n2912 = ~pi146 & ~pi210;
  assign n2913 = ~n2840 & ~n2873;
  assign n2914 = ~pi95 & ~n2913;
  assign n2915 = n2788 & ~n2914;
  assign n2916 = ~pi137 & ~n2915;
  assign n2917 = ~n2849 & ~n2916;
  assign n2918 = n2912 & ~n2917;
  assign n2919 = n2911 & ~n2918;
  assign n2920 = ~n2899 & n2919;
  assign n2921 = ~pi72 & ~n2717;
  assign n2922 = ~n2870 & n2921;
  assign n2923 = n2556 & ~n2922;
  assign n2924 = n2554 & ~n2923;
  assign n2925 = ~n2795 & n2924;
  assign n2926 = ~n2888 & n2921;
  assign n2927 = n2556 & ~n2926;
  assign n2928 = n2875 & ~n2927;
  assign n2929 = ~n2840 & ~n2928;
  assign n2930 = ~n2925 & n2929;
  assign n2931 = ~pi95 & ~n2930;
  assign n2932 = ~n2727 & ~n2931;
  assign n2933 = ~pi137 & ~n2932;
  assign n2934 = ~pi72 & n2725;
  assign n2935 = n2717 & n2934;
  assign n2936 = n2847 & ~n2935;
  assign n2937 = n2841 & ~n2936;
  assign n2938 = n2449 & n2726;
  assign n2939 = pi137 & ~n2938;
  assign n2940 = ~n2937 & n2939;
  assign n2941 = ~n2933 & ~n2940;
  assign n2942 = ~pi210 & ~n2941;
  assign n2943 = pi146 & n2942;
  assign n2944 = ~pi137 & ~n2727;
  assign n2945 = ~n2901 & ~n2924;
  assign n2946 = ~pi95 & ~n2945;
  assign n2947 = n2944 & ~n2946;
  assign n2948 = n2906 & ~n2936;
  assign n2949 = ~n2938 & ~n2948;
  assign n2950 = pi137 & ~n2949;
  assign n2951 = pi210 & ~n2950;
  assign n2952 = ~n2947 & n2951;
  assign n2953 = n2828 & ~n2952;
  assign n2954 = ~n2840 & ~n2924;
  assign n2955 = ~pi95 & ~n2954;
  assign n2956 = ~n2727 & ~n2955;
  assign n2957 = ~pi137 & ~n2956;
  assign n2958 = ~n2940 & ~n2957;
  assign n2959 = n2912 & ~n2958;
  assign n2960 = n2953 & ~n2959;
  assign n2961 = ~n2943 & n2960;
  assign n2962 = ~n2448 & ~n2961;
  assign n2963 = ~n2920 & n2962;
  assign n2964 = ~n2942 & n2953;
  assign n2965 = ~n2898 & n2911;
  assign n2966 = n2448 & ~n2965;
  assign n2967 = ~n2964 & n2966;
  assign n2968 = ~pi153 & ~n2967;
  assign n2969 = ~n2963 & n2968;
  assign n2970 = ~pi109 & ~n2696;
  assign n2971 = ~n2575 & ~n2970;
  assign n2972 = n2574 & ~n2971;
  assign n2973 = n2573 & ~n2972;
  assign n2974 = n2566 & ~n2973;
  assign n2975 = n2708 & ~n2974;
  assign n2976 = n2564 & ~n2975;
  assign n2977 = n2562 & ~n2976;
  assign n2978 = ~pi51 & ~n2977;
  assign n2979 = n2561 & ~n2978;
  assign n2980 = ~pi72 & ~n2979;
  assign n2981 = n2556 & ~n2980;
  assign n2982 = n2554 & ~n2981;
  assign n2983 = ~n2721 & n2982;
  assign n2984 = ~n2742 & ~n2983;
  assign n2985 = ~pi95 & ~n2984;
  assign n2986 = ~n2727 & ~n2985;
  assign n2987 = pi137 & ~n2986;
  assign n2988 = ~pi146 & ~n2448;
  assign n2989 = n2734 & ~n2988;
  assign n2990 = ~n2756 & n2989;
  assign n2991 = ~n2727 & ~n2749;
  assign n2992 = ~n2990 & n2991;
  assign n2993 = ~n2727 & n2989;
  assign n2994 = n2774 & n2993;
  assign n2995 = ~pi137 & ~n2994;
  assign n2996 = ~n2992 & n2995;
  assign n2997 = ~n2987 & ~n2996;
  assign n2998 = ~pi210 & ~n2997;
  assign n2999 = pi234 & ~n2998;
  assign n3000 = ~n2742 & ~n2982;
  assign n3001 = ~pi95 & ~n3000;
  assign n3002 = n2788 & ~n3001;
  assign n3003 = pi137 & ~n3002;
  assign n3004 = n2803 & ~n2988;
  assign n3005 = n2823 & n2988;
  assign n3006 = ~pi210 & ~pi234;
  assign n3007 = ~n3005 & n3006;
  assign n3008 = ~n3004 & n3007;
  assign n3009 = ~n3003 & n3008;
  assign n3010 = ~n2501 & ~n2982;
  assign n3011 = ~pi95 & ~n3010;
  assign n3012 = n2788 & ~n3011;
  assign n3013 = pi137 & ~n3012;
  assign n3014 = pi210 & ~n2787;
  assign n3015 = ~n3013 & n3014;
  assign n3016 = ~n3009 & ~n3015;
  assign n3017 = ~n2999 & n3016;
  assign n3018 = ~n2501 & ~n2983;
  assign n3019 = ~pi95 & ~n3018;
  assign n3020 = pi137 & ~n2727;
  assign n3021 = ~n3019 & n3020;
  assign n3022 = ~n2545 & n2944;
  assign n3023 = pi210 & pi234;
  assign n3024 = ~n3022 & n3023;
  assign n3025 = ~n3021 & n3024;
  assign n3026 = ~n3017 & ~n3025;
  assign n3027 = n2445 & ~n3026;
  assign n3028 = ~pi228 & ~n3027;
  assign n3029 = ~n2969 & n3028;
  assign n3030 = ~n2837 & ~n3029;
  assign n3031 = ~pi216 & ~n3030;
  assign n3032 = ~n2444 & ~n3031;
  assign n3033 = ~pi221 & ~n3032;
  assign n3034 = ~n2442 & ~n3033;
  assign n3035 = ~pi215 & ~n3034;
  assign n3036 = ~pi332 & ~pi1144;
  assign n3037 = pi215 & ~n3036;
  assign n3038 = pi299 & ~n3037;
  assign n3039 = ~n3035 & n3038;
  assign n3040 = ~pi224 & pi833;
  assign n3041 = pi222 & ~n3040;
  assign n3042 = ~pi223 & ~n3041;
  assign n3043 = n3036 & ~n3042;
  assign n3044 = pi224 & ~n2443;
  assign n3045 = ~pi222 & ~n3044;
  assign n3046 = ~pi332 & ~pi929;
  assign n3047 = n3040 & n3046;
  assign n3048 = ~n3045 & ~n3047;
  assign n3049 = ~pi223 & ~n3048;
  assign n3050 = ~n3043 & ~n3049;
  assign n3051 = ~pi299 & ~n3050;
  assign n3052 = ~pi222 & ~pi224;
  assign n3053 = pi198 & ~n2731;
  assign n3054 = ~pi198 & n2779;
  assign n3055 = ~n3053 & ~n3054;
  assign n3056 = pi142 & n3055;
  assign n3057 = ~pi198 & ~n2751;
  assign n3058 = ~pi142 & ~n3053;
  assign n3059 = ~n3057 & n3058;
  assign n3060 = n2816 & ~n3059;
  assign n3061 = ~n3056 & n3060;
  assign n3062 = ~pi144 & ~pi174;
  assign n3063 = ~pi189 & n3062;
  assign n3064 = ~pi223 & ~n3063;
  assign n3065 = ~pi198 & ~n2824;
  assign n3066 = pi198 & ~n2793;
  assign n3067 = ~pi142 & ~n3066;
  assign n3068 = ~n3065 & n3067;
  assign n3069 = ~pi198 & ~n2808;
  assign n3070 = ~n3066 & ~n3069;
  assign n3071 = pi142 & n3070;
  assign n3072 = n2828 & ~n3071;
  assign n3073 = ~n3068 & n3072;
  assign n3074 = n3064 & ~n3073;
  assign n3075 = ~n3061 & n3074;
  assign n3076 = ~pi223 & n3063;
  assign n3077 = pi234 & n3055;
  assign n3078 = ~pi234 & n3070;
  assign n3079 = ~pi332 & ~n3078;
  assign n3080 = ~n3077 & n3079;
  assign n3081 = n3076 & ~n3080;
  assign n3082 = ~n3075 & ~n3081;
  assign n3083 = n3052 & ~n3082;
  assign n3084 = n3051 & ~n3083;
  assign n3085 = ~pi39 & ~n3084;
  assign n3086 = ~n3039 & n3085;
  assign n3087 = pi234 & n2449;
  assign n3088 = ~pi332 & ~n3087;
  assign n3089 = ~pi95 & n2726;
  assign n3090 = ~n2449 & ~n3089;
  assign n3091 = pi234 & ~n3090;
  assign n3092 = ~pi32 & ~pi95;
  assign n3093 = n2450 & n3092;
  assign n3094 = n2842 & n3093;
  assign n3095 = n2557 & n3094;
  assign n3096 = ~pi234 & n3095;
  assign n3097 = ~n3091 & ~n3096;
  assign n3098 = pi137 & ~n3097;
  assign n3099 = n3088 & ~n3098;
  assign n3100 = ~pi223 & n3052;
  assign n3101 = ~n3099 & n3100;
  assign n3102 = ~n3050 & ~n3101;
  assign n3103 = ~pi299 & ~n3102;
  assign n3104 = pi105 & ~n3099;
  assign n3105 = ~n2446 & ~n3104;
  assign n3106 = pi228 & ~n3105;
  assign n3107 = ~pi332 & n3089;
  assign n3108 = ~pi137 & ~pi153;
  assign n3109 = n3107 & n3108;
  assign n3110 = pi137 & n3095;
  assign n3111 = n2445 & ~n3110;
  assign n3112 = ~pi228 & ~n3111;
  assign n3113 = ~n3109 & n3112;
  assign n3114 = ~n3106 & ~n3113;
  assign n3115 = ~pi216 & ~n3114;
  assign n3116 = ~n2444 & ~n3115;
  assign n3117 = ~pi221 & ~n3116;
  assign n3118 = ~n2442 & ~n3117;
  assign n3119 = ~pi215 & ~n3118;
  assign n3120 = ~n3037 & ~n3119;
  assign n3121 = pi299 & ~n3120;
  assign n3122 = ~n3103 & ~n3121;
  assign n3123 = pi39 & ~n3122;
  assign n3124 = ~pi38 & ~n3123;
  assign n3125 = ~n3086 & n3124;
  assign n3126 = pi105 & pi228;
  assign n3127 = n3088 & n3126;
  assign n3128 = n2445 & ~n3126;
  assign n3129 = ~pi216 & ~n3128;
  assign n3130 = ~n3127 & n3129;
  assign n3131 = ~n2444 & ~n3130;
  assign n3132 = ~pi221 & ~n3131;
  assign n3133 = ~n2442 & ~n3132;
  assign n3134 = ~pi215 & ~n3133;
  assign n3135 = ~n3037 & ~n3134;
  assign n3136 = ~pi215 & ~pi221;
  assign n3137 = n3129 & n3136;
  assign n3138 = ~n3099 & n3137;
  assign n3139 = n3135 & ~n3138;
  assign n3140 = pi299 & ~n3139;
  assign n3141 = ~n3103 & ~n3140;
  assign n3142 = ~pi39 & ~n3141;
  assign n3143 = pi299 & n3135;
  assign n3144 = ~n3088 & n3100;
  assign n3145 = n3051 & ~n3144;
  assign n3146 = ~n3143 & ~n3145;
  assign n3147 = pi39 & n3146;
  assign n3148 = pi38 & ~n3147;
  assign n3149 = ~n3142 & n3148;
  assign n3150 = ~pi100 & ~n3149;
  assign n3151 = ~n3125 & n3150;
  assign n3152 = pi228 & ~n2446;
  assign n3153 = ~pi210 & ~n2988;
  assign n3154 = pi95 & pi234;
  assign n3155 = ~pi137 & ~n3154;
  assign n3156 = ~n3153 & n3155;
  assign n3157 = ~n3097 & ~n3156;
  assign n3158 = ~pi332 & ~n3157;
  assign n3159 = pi105 & ~n3158;
  assign n3160 = n3152 & ~n3159;
  assign n3161 = ~pi137 & pi210;
  assign n3162 = ~pi252 & ~n3161;
  assign n3163 = ~n2988 & n3162;
  assign n3164 = n3107 & n3163;
  assign n3165 = n2988 & n3110;
  assign n3166 = n2445 & ~n3165;
  assign n3167 = ~n3164 & n3166;
  assign n3168 = pi252 & ~n2988;
  assign n3169 = ~n3153 & ~n3168;
  assign n3170 = n3109 & n3169;
  assign n3171 = ~n3167 & ~n3170;
  assign n3172 = ~pi228 & ~n3171;
  assign n3173 = ~pi216 & ~n3172;
  assign n3174 = ~n3160 & n3173;
  assign n3175 = ~n2444 & ~n3174;
  assign n3176 = ~pi221 & ~n3175;
  assign n3177 = ~n2442 & ~n3176;
  assign n3178 = ~pi215 & ~n3177;
  assign n3179 = ~n3037 & ~n3178;
  assign n3180 = pi299 & ~n3179;
  assign n3181 = ~pi38 & ~pi39;
  assign n3182 = pi142 & ~pi198;
  assign n3183 = ~pi137 & ~n3182;
  assign n3184 = ~n3097 & ~n3183;
  assign n3185 = n3088 & ~n3184;
  assign n3186 = n3064 & ~n3185;
  assign n3187 = ~pi137 & pi198;
  assign n3188 = ~pi95 & n3187;
  assign n3189 = ~n3090 & ~n3188;
  assign n3190 = n2816 & ~n3189;
  assign n3191 = n3095 & ~n3187;
  assign n3192 = n2828 & ~n3191;
  assign n3193 = n3076 & ~n3192;
  assign n3194 = ~n3190 & n3193;
  assign n3195 = ~n3186 & ~n3194;
  assign n3196 = n3052 & ~n3195;
  assign n3197 = ~n3050 & ~n3196;
  assign n3198 = ~pi299 & ~n3197;
  assign n3199 = n3181 & ~n3198;
  assign n3200 = ~n3180 & n3199;
  assign n3201 = ~n3146 & ~n3181;
  assign n3202 = pi100 & ~n3201;
  assign n3203 = ~n3200 & n3202;
  assign n3204 = ~pi87 & ~n3203;
  assign n3205 = ~n3151 & n3204;
  assign n3206 = ~pi38 & ~pi100;
  assign n3207 = ~pi39 & n3206;
  assign n3208 = ~n3146 & ~n3207;
  assign n3209 = n3122 & n3207;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = pi87 & ~n3210;
  assign n3212 = ~pi75 & ~n3211;
  assign n3213 = ~n3205 & n3212;
  assign n3214 = n3129 & ~n3160;
  assign n3215 = ~n2444 & ~n3214;
  assign n3216 = ~pi221 & ~n3215;
  assign n3217 = ~n2442 & ~n3216;
  assign n3218 = ~pi215 & ~n3217;
  assign n3219 = ~n3037 & ~n3218;
  assign n3220 = pi299 & ~n3219;
  assign n3221 = ~pi39 & ~pi87;
  assign n3222 = n3206 & n3221;
  assign n3223 = ~n3198 & n3222;
  assign n3224 = ~n3220 & n3223;
  assign n3225 = ~n3146 & ~n3222;
  assign n3226 = pi75 & ~n3225;
  assign n3227 = ~n3224 & n3226;
  assign n3228 = ~n3213 & ~n3227;
  assign n3229 = ~pi92 & ~n3228;
  assign n3230 = ~pi75 & ~pi87;
  assign n3231 = ~n3210 & n3230;
  assign n3232 = ~n3146 & ~n3230;
  assign n3233 = pi92 & ~n3232;
  assign n3234 = ~n3231 & n3233;
  assign n3235 = ~pi54 & ~n3234;
  assign n3236 = ~n3229 & n3235;
  assign n3237 = ~pi75 & ~pi92;
  assign n3238 = n3222 & n3237;
  assign n3239 = n3146 & ~n3238;
  assign n3240 = ~pi87 & ~pi100;
  assign n3241 = ~pi38 & n3240;
  assign n3242 = n3237 & n3241;
  assign n3243 = n3142 & n3242;
  assign n3244 = ~n3239 & ~n3243;
  assign n3245 = pi54 & n3244;
  assign n3246 = ~pi74 & ~n3245;
  assign n3247 = ~n3236 & n3246;
  assign n3248 = ~pi54 & n3244;
  assign n3249 = pi54 & ~n3146;
  assign n3250 = pi74 & ~n3249;
  assign n3251 = ~n3248 & n3250;
  assign n3252 = ~n3247 & ~n3251;
  assign n3253 = ~pi55 & ~n3252;
  assign n3254 = ~pi332 & n3097;
  assign n3255 = pi105 & ~n3254;
  assign n3256 = n3152 & ~n3255;
  assign n3257 = ~pi228 & n2445;
  assign n3258 = ~n3095 & n3257;
  assign n3259 = ~pi216 & ~n3258;
  assign n3260 = ~n3256 & n3259;
  assign n3261 = ~n2444 & ~n3260;
  assign n3262 = ~pi221 & ~n3261;
  assign n3263 = ~n2442 & ~n3262;
  assign n3264 = ~pi215 & ~n3263;
  assign n3265 = ~pi54 & ~pi74;
  assign n3266 = n3237 & n3265;
  assign n3267 = n3240 & n3266;
  assign n3268 = n3181 & n3267;
  assign n3269 = ~n3037 & n3268;
  assign n3270 = ~n3264 & n3269;
  assign n3271 = n3135 & ~n3268;
  assign n3272 = pi55 & ~n3271;
  assign n3273 = ~n3270 & n3272;
  assign n3274 = ~pi56 & ~n3273;
  assign n3275 = ~n3253 & n3274;
  assign n3276 = ~pi100 & n3181;
  assign n3277 = ~pi92 & n3230;
  assign n3278 = n3265 & n3277;
  assign n3279 = ~pi55 & n3278;
  assign n3280 = n3276 & n3279;
  assign n3281 = n3135 & ~n3280;
  assign n3282 = n3120 & n3280;
  assign n3283 = ~n3281 & ~n3282;
  assign n3284 = pi56 & ~n3283;
  assign n3285 = ~pi62 & ~n3284;
  assign n3286 = ~n3275 & n3285;
  assign n3287 = ~pi56 & ~n3283;
  assign n3288 = pi56 & n3135;
  assign n3289 = pi62 & ~n3288;
  assign n3290 = ~n3287 & n3289;
  assign n3291 = ~pi59 & ~n3290;
  assign n3292 = ~n3286 & n3291;
  assign n3293 = ~pi56 & ~pi62;
  assign n3294 = n3280 & n3293;
  assign n3295 = n3138 & n3294;
  assign n3296 = pi59 & n3135;
  assign n3297 = ~n3295 & n3296;
  assign n3298 = ~pi57 & ~n3297;
  assign n3299 = ~n3292 & n3298;
  assign n3300 = ~pi59 & n3295;
  assign n3301 = n3135 & ~n3300;
  assign n3302 = pi57 & ~n3301;
  assign po153 = n3299 | n3302;
  assign n3304 = pi223 & ~pi1146;
  assign n3305 = ~pi299 & ~n3304;
  assign n3306 = ~pi222 & pi224;
  assign n3307 = pi276 & n3306;
  assign n3308 = ~pi939 & n3040;
  assign n3309 = ~pi1146 & ~n3040;
  assign n3310 = pi222 & ~n3309;
  assign n3311 = ~n3308 & n3310;
  assign n3312 = ~pi223 & ~n3311;
  assign n3313 = ~n3307 & n3312;
  assign n3314 = n3305 & ~n3313;
  assign n3315 = pi215 & pi1146;
  assign n3316 = ~pi939 & n2437;
  assign n3317 = ~pi1146 & ~n2437;
  assign n3318 = pi221 & ~n3317;
  assign n3319 = ~n3316 & n3318;
  assign n3320 = ~n3315 & ~n3319;
  assign n3321 = ~pi228 & n3095;
  assign n3322 = ~pi216 & n3321;
  assign n3323 = n3320 & n3322;
  assign n3324 = pi216 & ~pi221;
  assign n3325 = pi276 & n3324;
  assign n3326 = ~n3319 & ~n3325;
  assign n3327 = ~pi215 & ~n3326;
  assign n3328 = ~n3315 & ~n3327;
  assign n3329 = ~pi216 & ~pi221;
  assign n3330 = ~pi215 & n3329;
  assign n3331 = ~n3126 & n3330;
  assign n3332 = n3328 & ~n3331;
  assign n3333 = pi299 & ~n3332;
  assign n3334 = ~n3323 & n3333;
  assign n3335 = ~n3314 & ~n3334;
  assign n3336 = ~pi154 & ~n3335;
  assign n3337 = pi299 & ~n3328;
  assign n3338 = ~n3314 & ~n3337;
  assign n3339 = pi154 & ~n3338;
  assign n3340 = n3207 & ~n3339;
  assign n3341 = ~n3336 & n3340;
  assign n3342 = pi154 & ~n3328;
  assign n3343 = ~pi154 & ~n3332;
  assign n3344 = ~n3342 & ~n3343;
  assign n3345 = pi299 & ~n3344;
  assign n3346 = ~n3314 & ~n3345;
  assign n3347 = ~n3207 & n3346;
  assign n3348 = ~n3341 & ~n3347;
  assign n3349 = pi87 & ~n3348;
  assign n3350 = pi39 & ~n3095;
  assign n3351 = ~pi70 & n2976;
  assign n3352 = ~n2524 & ~n2843;
  assign n3353 = ~n3351 & n3352;
  assign n3354 = ~pi51 & ~n3353;
  assign n3355 = n2559 & ~n3354;
  assign n3356 = n2921 & ~n3355;
  assign n3357 = ~n2555 & ~n3356;
  assign n3358 = n2725 & ~n3357;
  assign n3359 = pi40 & ~n2552;
  assign n3360 = pi32 & ~n2499;
  assign n3361 = ~n3359 & ~n3360;
  assign n3362 = ~n3358 & n3361;
  assign n3363 = ~pi95 & ~n3362;
  assign n3364 = ~n2727 & ~n3363;
  assign n3365 = ~pi39 & ~n3364;
  assign n3366 = ~n3350 & ~n3365;
  assign n3367 = ~pi216 & ~pi228;
  assign n3368 = n3320 & n3367;
  assign n3369 = n3366 & n3368;
  assign n3370 = n3333 & ~n3369;
  assign n3371 = ~n3314 & ~n3370;
  assign n3372 = ~pi154 & ~n3371;
  assign n3373 = ~pi38 & ~n3339;
  assign n3374 = ~n3372 & n3373;
  assign n3375 = pi38 & n3346;
  assign n3376 = ~pi100 & ~n3375;
  assign n3377 = ~n3374 & n3376;
  assign n3378 = ~pi146 & ~n3095;
  assign n3379 = ~pi252 & n3095;
  assign n3380 = pi146 & ~n3379;
  assign n3381 = ~n3378 & ~n3380;
  assign n3382 = pi152 & ~n3381;
  assign n3383 = ~pi161 & ~pi166;
  assign n3384 = n3381 & ~n3383;
  assign n3385 = n3379 & n3383;
  assign n3386 = ~pi152 & ~n3385;
  assign n3387 = ~n3384 & n3386;
  assign n3388 = ~n3382 & ~n3387;
  assign n3389 = ~pi38 & ~pi216;
  assign n3390 = ~pi228 & n3389;
  assign n3391 = ~pi154 & pi299;
  assign n3392 = ~pi39 & n3391;
  assign n3393 = n3390 & n3392;
  assign n3394 = n3320 & n3393;
  assign n3395 = n3388 & n3394;
  assign n3396 = pi100 & ~n3346;
  assign n3397 = ~n3395 & n3396;
  assign n3398 = ~pi87 & ~n3397;
  assign n3399 = ~n3377 & n3398;
  assign n3400 = ~n3349 & ~n3399;
  assign n3401 = ~pi75 & ~n3400;
  assign n3402 = pi75 & n3346;
  assign n3403 = ~pi92 & ~n3402;
  assign n3404 = ~n3401 & n3403;
  assign n3405 = n3230 & n3341;
  assign n3406 = n3230 & n3276;
  assign n3407 = n3346 & ~n3406;
  assign n3408 = pi92 & ~n3407;
  assign n3409 = ~n3405 & n3408;
  assign n3410 = n3265 & ~n3409;
  assign n3411 = ~n3404 & n3410;
  assign n3412 = ~n3265 & n3346;
  assign n3413 = ~pi55 & ~n3412;
  assign n3414 = ~n3411 & n3413;
  assign n3415 = n3323 & ~n3342;
  assign n3416 = n3268 & n3415;
  assign n3417 = pi55 & ~n3344;
  assign n3418 = ~n3416 & n3417;
  assign n3419 = ~pi56 & ~n3418;
  assign n3420 = ~n3414 & n3419;
  assign n3421 = ~pi55 & n3268;
  assign n3422 = ~n3344 & n3421;
  assign n3423 = ~n3415 & n3422;
  assign n3424 = ~n3280 & ~n3344;
  assign n3425 = pi56 & ~n3424;
  assign n3426 = ~n3423 & n3425;
  assign n3427 = ~pi62 & ~n3426;
  assign n3428 = ~n3420 & n3427;
  assign n3429 = ~pi57 & ~pi59;
  assign n3430 = ~pi56 & n3279;
  assign n3431 = n3276 & n3430;
  assign n3432 = ~n3344 & ~n3431;
  assign n3433 = ~n3423 & ~n3432;
  assign n3434 = pi62 & ~n3433;
  assign n3435 = n3429 & ~n3434;
  assign n3436 = ~n3428 & n3435;
  assign n3437 = n3344 & ~n3429;
  assign n3438 = ~pi239 & ~n3437;
  assign n3439 = ~n3436 & n3438;
  assign n3440 = n2717 & n3093;
  assign n3441 = ~n2449 & ~n3440;
  assign n3442 = ~pi224 & n3441;
  assign n3443 = ~n3052 & ~n3307;
  assign n3444 = ~n3442 & ~n3443;
  assign n3445 = n3312 & ~n3444;
  assign n3446 = ~n3304 & ~n3445;
  assign n3447 = ~pi299 & ~n3446;
  assign n3448 = ~pi72 & ~n3355;
  assign n3449 = ~n2555 & ~n3448;
  assign n3450 = n2725 & ~n3449;
  assign n3451 = n3361 & ~n3450;
  assign n3452 = ~pi95 & ~n3451;
  assign n3453 = n2788 & ~n3452;
  assign n3454 = ~pi228 & n3453;
  assign n3455 = n3126 & n3441;
  assign n3456 = ~n3454 & ~n3455;
  assign n3457 = ~pi154 & ~n3456;
  assign n3458 = pi105 & ~n3441;
  assign n3459 = pi228 & ~n3458;
  assign n3460 = ~n2727 & ~n3441;
  assign n3461 = ~pi228 & ~n3460;
  assign n3462 = ~n3459 & ~n3461;
  assign n3463 = pi154 & ~n3462;
  assign n3464 = n3330 & ~n3463;
  assign n3465 = ~n3457 & n3464;
  assign n3466 = pi299 & n3328;
  assign n3467 = ~n3465 & n3466;
  assign n3468 = ~n3447 & ~n3467;
  assign n3469 = ~pi39 & ~n3468;
  assign n3470 = n2449 & n3126;
  assign n3471 = n3330 & n3470;
  assign n3472 = n3344 & ~n3471;
  assign n3473 = pi299 & ~n3472;
  assign n3474 = ~pi223 & ~pi299;
  assign n3475 = n3052 & n3474;
  assign n3476 = n2449 & n3475;
  assign n3477 = ~n3314 & ~n3476;
  assign n3478 = ~n3473 & n3477;
  assign n3479 = pi154 & ~n3472;
  assign n3480 = n3323 & ~n3479;
  assign n3481 = ~n3472 & ~n3480;
  assign n3482 = pi299 & ~n3481;
  assign n3483 = ~n3478 & ~n3482;
  assign n3484 = pi39 & ~n3483;
  assign n3485 = n3206 & ~n3484;
  assign n3486 = ~n3469 & n3485;
  assign n3487 = pi100 & n3395;
  assign n3488 = ~n3206 & ~n3478;
  assign n3489 = ~n3487 & n3488;
  assign n3490 = ~n3486 & ~n3489;
  assign n3491 = ~pi87 & ~n3490;
  assign n3492 = n3207 & n3482;
  assign n3493 = pi87 & ~n3478;
  assign n3494 = ~n3492 & n3493;
  assign n3495 = ~pi75 & ~n3494;
  assign n3496 = ~n3491 & n3495;
  assign n3497 = pi75 & n3478;
  assign n3498 = ~pi92 & ~n3497;
  assign n3499 = ~n3496 & n3498;
  assign n3500 = n3406 & n3482;
  assign n3501 = pi92 & ~n3478;
  assign n3502 = ~n3500 & n3501;
  assign n3503 = n3265 & ~n3502;
  assign n3504 = ~n3499 & n3503;
  assign n3505 = ~n3265 & n3478;
  assign n3506 = ~pi55 & ~n3505;
  assign n3507 = ~n3504 & n3506;
  assign n3508 = n3268 & n3480;
  assign n3509 = pi55 & ~n3472;
  assign n3510 = ~n3508 & n3509;
  assign n3511 = ~pi56 & ~n3510;
  assign n3512 = ~n3507 & n3511;
  assign n3513 = n3421 & n3481;
  assign n3514 = ~n3280 & ~n3472;
  assign n3515 = pi56 & ~n3514;
  assign n3516 = ~n3513 & n3515;
  assign n3517 = ~pi62 & ~n3516;
  assign n3518 = ~n3512 & n3517;
  assign n3519 = ~n3431 & ~n3472;
  assign n3520 = ~pi56 & n3513;
  assign n3521 = ~n3519 & ~n3520;
  assign n3522 = pi62 & ~n3521;
  assign n3523 = n3429 & ~n3522;
  assign n3524 = ~n3518 & n3523;
  assign n3525 = ~n3429 & n3472;
  assign n3526 = pi239 & ~n3525;
  assign n3527 = ~n3524 & n3526;
  assign po154 = n3439 | n3527;
  assign n3529 = ~pi927 & n2437;
  assign n3530 = ~pi1145 & ~n2437;
  assign n3531 = pi221 & ~n3530;
  assign n3532 = ~n3529 & n3531;
  assign n3533 = pi216 & pi274;
  assign n3534 = ~pi221 & ~n3533;
  assign n3535 = ~pi151 & n3456;
  assign n3536 = pi151 & n3462;
  assign n3537 = ~pi216 & ~n3536;
  assign n3538 = ~n3535 & n3537;
  assign n3539 = n3534 & ~n3538;
  assign n3540 = ~n3532 & ~n3539;
  assign n3541 = ~pi215 & ~n3540;
  assign n3542 = pi215 & pi1145;
  assign n3543 = pi299 & ~n3542;
  assign n3544 = ~n3541 & n3543;
  assign n3545 = ~pi927 & n3040;
  assign n3546 = ~pi1145 & ~n3040;
  assign n3547 = pi222 & ~n3546;
  assign n3548 = ~n3545 & n3547;
  assign n3549 = pi224 & pi274;
  assign n3550 = ~pi222 & ~n3549;
  assign n3551 = ~n3442 & n3550;
  assign n3552 = ~n3548 & ~n3551;
  assign n3553 = ~pi223 & ~n3552;
  assign n3554 = pi223 & pi1145;
  assign n3555 = ~pi299 & ~n3554;
  assign n3556 = ~n3553 & n3555;
  assign n3557 = ~pi39 & ~n3556;
  assign n3558 = ~n3544 & n3557;
  assign n3559 = n3306 & ~n3549;
  assign n3560 = ~n3548 & ~n3559;
  assign n3561 = ~pi223 & ~n3560;
  assign n3562 = ~n3554 & ~n3561;
  assign n3563 = ~pi299 & ~n3562;
  assign n3564 = ~n3476 & ~n3563;
  assign n3565 = ~pi151 & ~n3126;
  assign n3566 = ~n3470 & ~n3565;
  assign n3567 = ~pi151 & n3321;
  assign n3568 = ~n3566 & ~n3567;
  assign n3569 = ~pi216 & ~n3568;
  assign n3570 = n3534 & ~n3569;
  assign n3571 = ~n3532 & ~n3570;
  assign n3572 = ~pi215 & ~n3571;
  assign n3573 = ~n3542 & ~n3572;
  assign n3574 = pi299 & ~n3573;
  assign n3575 = n3564 & ~n3574;
  assign n3576 = pi39 & ~n3575;
  assign n3577 = ~pi38 & ~n3576;
  assign n3578 = ~n3558 & n3577;
  assign n3579 = ~pi216 & ~n3565;
  assign n3580 = n3534 & ~n3579;
  assign n3581 = ~n3532 & ~n3580;
  assign n3582 = ~pi215 & ~n3581;
  assign n3583 = ~n3542 & ~n3582;
  assign n3584 = n3136 & n3470;
  assign n3585 = ~n3533 & n3584;
  assign n3586 = n3583 & ~n3585;
  assign n3587 = pi299 & ~n3586;
  assign n3588 = n3564 & ~n3587;
  assign n3589 = pi38 & n3588;
  assign n3590 = ~pi100 & ~n3589;
  assign n3591 = ~n3578 & n3590;
  assign n3592 = ~pi228 & n3388;
  assign n3593 = ~n2449 & n3126;
  assign n3594 = ~n3592 & ~n3593;
  assign n3595 = ~pi151 & n3594;
  assign n3596 = n3569 & ~n3595;
  assign n3597 = n3534 & ~n3596;
  assign n3598 = ~n3532 & ~n3597;
  assign n3599 = ~pi215 & ~n3598;
  assign n3600 = ~n3542 & ~n3599;
  assign n3601 = pi299 & ~n3600;
  assign n3602 = n3181 & n3564;
  assign n3603 = ~n3601 & n3602;
  assign n3604 = ~n3181 & n3588;
  assign n3605 = pi100 & ~n3604;
  assign n3606 = ~n3603 & n3605;
  assign n3607 = ~n3591 & ~n3606;
  assign n3608 = ~pi87 & ~n3607;
  assign n3609 = ~n3207 & n3588;
  assign n3610 = n3207 & n3575;
  assign n3611 = ~n3609 & ~n3610;
  assign n3612 = pi87 & n3611;
  assign n3613 = ~pi75 & ~n3612;
  assign n3614 = ~n3608 & n3613;
  assign n3615 = pi75 & n3588;
  assign n3616 = ~pi92 & ~n3615;
  assign n3617 = ~n3614 & n3616;
  assign n3618 = n3230 & ~n3611;
  assign n3619 = ~n3230 & n3588;
  assign n3620 = pi92 & ~n3619;
  assign n3621 = ~n3618 & n3620;
  assign n3622 = n3265 & ~n3621;
  assign n3623 = ~n3617 & n3622;
  assign n3624 = ~n3265 & n3588;
  assign n3625 = ~pi55 & ~n3624;
  assign n3626 = ~n3623 & n3625;
  assign n3627 = n3268 & n3573;
  assign n3628 = ~n3268 & n3586;
  assign n3629 = pi55 & ~n3628;
  assign n3630 = ~n3627 & n3629;
  assign n3631 = ~pi56 & ~n3630;
  assign n3632 = ~n3626 & n3631;
  assign n3633 = n3280 & ~n3573;
  assign n3634 = ~n3280 & ~n3586;
  assign n3635 = pi56 & ~n3634;
  assign n3636 = ~n3633 & n3635;
  assign n3637 = ~pi62 & ~n3636;
  assign n3638 = ~n3632 & n3637;
  assign n3639 = n3431 & n3573;
  assign n3640 = ~n3431 & n3586;
  assign n3641 = pi62 & ~n3640;
  assign n3642 = ~n3639 & n3641;
  assign n3643 = pi235 & n3429;
  assign n3644 = ~n3642 & n3643;
  assign n3645 = ~n3638 & n3644;
  assign n3646 = ~n3532 & ~n3542;
  assign n3647 = n3322 & n3646;
  assign n3648 = pi299 & ~n3583;
  assign n3649 = ~n3647 & n3648;
  assign n3650 = n3276 & ~n3563;
  assign n3651 = ~n3649 & n3650;
  assign n3652 = ~n3563 & ~n3648;
  assign n3653 = ~n3207 & n3652;
  assign n3654 = ~n3651 & ~n3653;
  assign n3655 = pi87 & ~n3654;
  assign n3656 = ~pi100 & n3366;
  assign n3657 = ~pi39 & pi100;
  assign n3658 = n3388 & n3657;
  assign n3659 = ~n3656 & ~n3658;
  assign n3660 = n3390 & n3646;
  assign n3661 = ~n3659 & n3660;
  assign n3662 = n3648 & ~n3661;
  assign n3663 = ~pi87 & ~n3563;
  assign n3664 = ~n3662 & n3663;
  assign n3665 = ~n3655 & ~n3664;
  assign n3666 = ~pi75 & ~n3665;
  assign n3667 = pi75 & n3652;
  assign n3668 = ~pi92 & ~n3667;
  assign n3669 = ~n3666 & n3668;
  assign n3670 = n3230 & n3651;
  assign n3671 = ~n3406 & n3652;
  assign n3672 = pi92 & ~n3671;
  assign n3673 = ~n3670 & n3672;
  assign n3674 = n3265 & ~n3673;
  assign n3675 = ~n3669 & n3674;
  assign n3676 = ~n3265 & n3652;
  assign n3677 = ~pi55 & ~n3676;
  assign n3678 = ~n3675 & n3677;
  assign n3679 = n3268 & n3647;
  assign n3680 = pi55 & ~n3583;
  assign n3681 = ~n3679 & n3680;
  assign n3682 = ~pi56 & ~n3681;
  assign n3683 = ~n3678 & n3682;
  assign n3684 = n3280 & n3647;
  assign n3685 = ~n3583 & ~n3684;
  assign n3686 = pi56 & ~n3685;
  assign n3687 = ~pi62 & ~n3686;
  assign n3688 = ~n3683 & n3687;
  assign n3689 = ~pi56 & n3684;
  assign n3690 = pi62 & ~n3583;
  assign n3691 = ~n3689 & n3690;
  assign n3692 = ~pi235 & n3429;
  assign n3693 = ~n3691 & n3692;
  assign n3694 = ~n3688 & n3693;
  assign n3695 = pi235 & n3585;
  assign n3696 = ~n3429 & ~n3695;
  assign n3697 = n3583 & n3696;
  assign n3698 = ~n3694 & ~n3697;
  assign po155 = ~n3645 & n3698;
  assign n3700 = pi223 & pi1143;
  assign n3701 = ~pi299 & ~n3700;
  assign n3702 = ~pi944 & n3040;
  assign n3703 = ~pi1143 & ~n3040;
  assign n3704 = pi222 & ~n3703;
  assign n3705 = ~n3702 & n3704;
  assign n3706 = pi224 & pi264;
  assign n3707 = ~pi222 & ~n3706;
  assign n3708 = ~pi284 & n3441;
  assign n3709 = ~pi224 & ~n3708;
  assign n3710 = n3707 & ~n3709;
  assign n3711 = ~n3705 & ~n3710;
  assign n3712 = ~n3441 & n3707;
  assign n3713 = n3711 & ~n3712;
  assign n3714 = ~pi223 & ~n3713;
  assign n3715 = n3701 & ~n3714;
  assign n3716 = ~pi39 & ~n3715;
  assign n3717 = pi215 & pi1143;
  assign n3718 = pi299 & ~n3717;
  assign n3719 = ~pi944 & n2437;
  assign n3720 = ~pi1143 & ~n2437;
  assign n3721 = pi221 & ~n3720;
  assign n3722 = ~n3719 & n3721;
  assign n3723 = pi216 & pi264;
  assign n3724 = ~pi221 & ~n3723;
  assign n3725 = pi284 & ~n2449;
  assign n3726 = pi105 & ~n3725;
  assign n3727 = ~pi105 & pi146;
  assign n3728 = pi228 & ~n3727;
  assign n3729 = ~n3726 & n3728;
  assign n3730 = ~n3458 & n3729;
  assign n3731 = pi146 & ~n3453;
  assign n3732 = ~pi146 & n3460;
  assign n3733 = pi284 & ~n3732;
  assign n3734 = ~n3731 & n3733;
  assign n3735 = ~pi146 & ~pi284;
  assign n3736 = ~n3364 & n3735;
  assign n3737 = ~n3734 & ~n3736;
  assign n3738 = ~pi228 & ~n3737;
  assign n3739 = ~n3730 & ~n3738;
  assign n3740 = ~pi216 & ~n3739;
  assign n3741 = n3724 & ~n3740;
  assign n3742 = ~n3722 & ~n3741;
  assign n3743 = ~pi215 & ~n3742;
  assign n3744 = n3718 & ~n3743;
  assign n3745 = n3716 & ~n3744;
  assign n3746 = ~pi224 & n3725;
  assign n3747 = n3707 & ~n3746;
  assign n3748 = ~n3705 & ~n3747;
  assign n3749 = ~pi223 & ~n3748;
  assign n3750 = ~n3700 & ~n3749;
  assign n3751 = ~pi299 & ~n3750;
  assign n3752 = pi284 & n3095;
  assign n3753 = ~n3378 & ~n3752;
  assign n3754 = ~pi228 & ~n3753;
  assign n3755 = ~n3729 & ~n3754;
  assign n3756 = ~pi216 & ~n3755;
  assign n3757 = n3724 & ~n3756;
  assign n3758 = ~n3722 & ~n3757;
  assign n3759 = ~pi215 & ~n3758;
  assign n3760 = ~n3717 & ~n3759;
  assign n3761 = pi299 & ~n3760;
  assign n3762 = ~n3751 & ~n3761;
  assign n3763 = pi39 & ~n3762;
  assign n3764 = ~pi38 & ~n3763;
  assign n3765 = ~n3745 & n3764;
  assign n3766 = ~n3470 & ~n3729;
  assign n3767 = ~pi146 & ~pi228;
  assign n3768 = n3766 & ~n3767;
  assign n3769 = ~pi216 & ~n3768;
  assign n3770 = n3724 & ~n3769;
  assign n3771 = ~n3722 & ~n3770;
  assign n3772 = ~pi215 & ~n3771;
  assign n3773 = ~n3717 & ~n3772;
  assign n3774 = n3584 & ~n3723;
  assign n3775 = n3773 & ~n3774;
  assign n3776 = pi299 & ~n3775;
  assign n3777 = ~n3751 & ~n3776;
  assign n3778 = pi38 & n3777;
  assign n3779 = ~pi100 & ~n3778;
  assign n3780 = ~n3765 & n3779;
  assign n3781 = pi252 & n2448;
  assign n3782 = ~pi284 & ~n3781;
  assign n3783 = n3095 & n3782;
  assign n3784 = ~pi228 & ~n3783;
  assign n3785 = ~n3380 & n3784;
  assign n3786 = ~n3729 & ~n3785;
  assign n3787 = ~pi216 & ~n3786;
  assign n3788 = n3724 & ~n3787;
  assign n3789 = ~n3722 & ~n3788;
  assign n3790 = ~pi215 & ~n3789;
  assign n3791 = ~n3717 & ~n3790;
  assign n3792 = pi299 & ~n3791;
  assign n3793 = n3181 & ~n3751;
  assign n3794 = ~n3792 & n3793;
  assign n3795 = ~n3181 & n3777;
  assign n3796 = pi100 & ~n3795;
  assign n3797 = ~n3794 & n3796;
  assign n3798 = ~n3780 & ~n3797;
  assign n3799 = ~pi87 & ~n3798;
  assign n3800 = ~n3207 & n3777;
  assign n3801 = n3207 & n3762;
  assign n3802 = ~n3800 & ~n3801;
  assign n3803 = pi87 & n3802;
  assign n3804 = ~pi75 & ~n3803;
  assign n3805 = ~n3799 & n3804;
  assign n3806 = pi75 & n3777;
  assign n3807 = ~pi92 & ~n3806;
  assign n3808 = ~n3805 & n3807;
  assign n3809 = n3230 & ~n3802;
  assign n3810 = ~n3230 & n3777;
  assign n3811 = pi92 & ~n3810;
  assign n3812 = ~n3809 & n3811;
  assign n3813 = n3265 & ~n3812;
  assign n3814 = ~n3808 & n3813;
  assign n3815 = ~n3265 & n3777;
  assign n3816 = ~pi55 & ~n3815;
  assign n3817 = ~n3814 & n3816;
  assign n3818 = n3268 & n3760;
  assign n3819 = ~n3268 & n3775;
  assign n3820 = pi55 & ~n3819;
  assign n3821 = ~n3818 & n3820;
  assign n3822 = ~pi56 & ~n3821;
  assign n3823 = ~n3817 & n3822;
  assign n3824 = n3280 & ~n3760;
  assign n3825 = ~n3280 & ~n3775;
  assign n3826 = pi56 & ~n3825;
  assign n3827 = ~n3824 & n3826;
  assign n3828 = ~pi62 & ~n3827;
  assign n3829 = ~n3823 & n3828;
  assign n3830 = n3431 & n3760;
  assign n3831 = ~n3431 & n3775;
  assign n3832 = pi62 & ~n3831;
  assign n3833 = ~n3830 & n3832;
  assign n3834 = pi238 & n3429;
  assign n3835 = ~n3833 & n3834;
  assign n3836 = ~n3829 & n3835;
  assign n3837 = ~pi146 & ~n3453;
  assign n3838 = pi146 & n3460;
  assign n3839 = ~pi284 & ~n3838;
  assign n3840 = pi146 & pi284;
  assign n3841 = ~n3364 & n3840;
  assign n3842 = ~n3839 & ~n3841;
  assign n3843 = ~n3837 & ~n3842;
  assign n3844 = ~pi228 & ~n3843;
  assign n3845 = n3126 & ~n3441;
  assign n3846 = ~n3729 & ~n3845;
  assign n3847 = ~n3844 & n3846;
  assign n3848 = ~pi216 & ~n3847;
  assign n3849 = n3724 & ~n3848;
  assign n3850 = ~n3722 & ~n3849;
  assign n3851 = ~pi215 & ~n3850;
  assign n3852 = n3718 & ~n3851;
  assign n3853 = n3701 & n3711;
  assign n3854 = n3716 & ~n3853;
  assign n3855 = ~n3852 & n3854;
  assign n3856 = n2449 & n3100;
  assign n3857 = n3751 & ~n3856;
  assign n3858 = ~n3754 & n3766;
  assign n3859 = ~pi216 & ~n3858;
  assign n3860 = n3724 & ~n3859;
  assign n3861 = ~n3722 & ~n3860;
  assign n3862 = ~pi215 & ~n3861;
  assign n3863 = ~n3717 & ~n3862;
  assign n3864 = pi299 & ~n3863;
  assign n3865 = ~n3857 & ~n3864;
  assign n3866 = pi39 & ~n3865;
  assign n3867 = ~pi38 & ~n3866;
  assign n3868 = ~n3855 & n3867;
  assign n3869 = pi299 & ~n3773;
  assign n3870 = ~n3857 & ~n3869;
  assign n3871 = pi38 & n3870;
  assign n3872 = ~pi100 & ~n3871;
  assign n3873 = ~n3868 & n3872;
  assign n3874 = n3766 & ~n3785;
  assign n3875 = ~pi216 & ~n3874;
  assign n3876 = n3724 & ~n3875;
  assign n3877 = ~n3722 & ~n3876;
  assign n3878 = ~pi215 & ~n3877;
  assign n3879 = ~n3717 & ~n3878;
  assign n3880 = pi299 & ~n3879;
  assign n3881 = n3181 & ~n3857;
  assign n3882 = ~n3880 & n3881;
  assign n3883 = ~n3181 & n3870;
  assign n3884 = pi100 & ~n3883;
  assign n3885 = ~n3882 & n3884;
  assign n3886 = ~n3873 & ~n3885;
  assign n3887 = ~pi87 & ~n3886;
  assign n3888 = ~n3207 & n3870;
  assign n3889 = n3207 & n3865;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = pi87 & n3890;
  assign n3892 = ~pi75 & ~n3891;
  assign n3893 = ~n3887 & n3892;
  assign n3894 = pi75 & n3870;
  assign n3895 = ~pi92 & ~n3894;
  assign n3896 = ~n3893 & n3895;
  assign n3897 = n3230 & ~n3890;
  assign n3898 = ~n3230 & n3870;
  assign n3899 = pi92 & ~n3898;
  assign n3900 = ~n3897 & n3899;
  assign n3901 = n3265 & ~n3900;
  assign n3902 = ~n3896 & n3901;
  assign n3903 = ~n3265 & n3870;
  assign n3904 = ~pi55 & ~n3903;
  assign n3905 = ~n3902 & n3904;
  assign n3906 = n3268 & n3863;
  assign n3907 = ~n3268 & n3773;
  assign n3908 = pi55 & ~n3907;
  assign n3909 = ~n3906 & n3908;
  assign n3910 = ~pi56 & ~n3909;
  assign n3911 = ~n3905 & n3910;
  assign n3912 = n3280 & ~n3863;
  assign n3913 = ~n3280 & ~n3773;
  assign n3914 = pi56 & ~n3913;
  assign n3915 = ~n3912 & n3914;
  assign n3916 = ~pi62 & ~n3915;
  assign n3917 = ~n3911 & n3916;
  assign n3918 = n3431 & n3863;
  assign n3919 = ~n3431 & n3773;
  assign n3920 = pi62 & ~n3919;
  assign n3921 = ~n3918 & n3920;
  assign n3922 = ~pi238 & n3429;
  assign n3923 = ~n3921 & n3922;
  assign n3924 = ~n3917 & n3923;
  assign n3925 = pi238 & n3774;
  assign n3926 = ~n3429 & ~n3925;
  assign n3927 = n3773 & n3926;
  assign n3928 = ~n3924 & ~n3927;
  assign po156 = ~n3836 & n3928;
  assign n3930 = pi215 & pi1142;
  assign n3931 = pi299 & ~n3930;
  assign n3932 = ~pi932 & n2437;
  assign n3933 = ~pi1142 & ~n2437;
  assign n3934 = pi221 & ~n3933;
  assign n3935 = ~n3932 & n3934;
  assign n3936 = pi216 & pi277;
  assign n3937 = ~pi221 & ~n3936;
  assign n3938 = ~pi262 & n3460;
  assign n3939 = ~pi172 & ~n3938;
  assign n3940 = pi172 & ~pi262;
  assign n3941 = n3453 & n3940;
  assign n3942 = ~n3939 & ~n3941;
  assign n3943 = pi262 & n3364;
  assign n3944 = ~pi228 & ~n3943;
  assign n3945 = ~n3942 & n3944;
  assign n3946 = pi262 & ~n2449;
  assign n3947 = pi105 & n3946;
  assign n3948 = ~n3440 & n3947;
  assign n3949 = ~pi105 & pi172;
  assign n3950 = pi228 & ~n3949;
  assign n3951 = ~n3948 & n3950;
  assign n3952 = ~n3458 & n3951;
  assign n3953 = ~pi216 & ~n3952;
  assign n3954 = ~n3945 & n3953;
  assign n3955 = n3937 & ~n3954;
  assign n3956 = ~n3935 & ~n3955;
  assign n3957 = ~pi215 & ~n3956;
  assign n3958 = n3931 & ~n3957;
  assign n3959 = pi223 & pi1142;
  assign n3960 = ~pi299 & ~n3959;
  assign n3961 = ~pi932 & n3040;
  assign n3962 = ~pi1142 & ~n3040;
  assign n3963 = pi222 & ~n3962;
  assign n3964 = ~n3961 & n3963;
  assign n3965 = pi224 & pi277;
  assign n3966 = ~pi222 & ~n3965;
  assign n3967 = ~pi262 & n3441;
  assign n3968 = ~pi224 & ~n3967;
  assign n3969 = n3966 & ~n3968;
  assign n3970 = ~n3964 & ~n3969;
  assign n3971 = n3960 & n3970;
  assign n3972 = ~n3441 & n3966;
  assign n3973 = n3970 & ~n3972;
  assign n3974 = ~pi223 & ~n3973;
  assign n3975 = n3960 & ~n3974;
  assign n3976 = ~pi39 & ~n3975;
  assign n3977 = ~n3971 & n3976;
  assign n3978 = ~n3958 & n3977;
  assign n3979 = ~pi224 & n3946;
  assign n3980 = n3966 & ~n3979;
  assign n3981 = ~n3964 & ~n3980;
  assign n3982 = ~pi223 & ~n3981;
  assign n3983 = ~n3959 & ~n3982;
  assign n3984 = ~pi299 & ~n3983;
  assign n3985 = ~n3856 & n3984;
  assign n3986 = ~pi262 & n3095;
  assign n3987 = pi172 & ~pi228;
  assign n3988 = ~n3321 & ~n3987;
  assign n3989 = ~n3986 & ~n3988;
  assign n3990 = ~n3947 & ~n3949;
  assign n3991 = pi228 & ~n3990;
  assign n3992 = ~n3470 & ~n3991;
  assign n3993 = ~n3989 & n3992;
  assign n3994 = ~pi216 & ~n3993;
  assign n3995 = n3937 & ~n3994;
  assign n3996 = ~n3935 & ~n3995;
  assign n3997 = ~pi215 & ~n3996;
  assign n3998 = ~n3930 & ~n3997;
  assign n3999 = pi299 & ~n3998;
  assign n4000 = ~n3985 & ~n3999;
  assign n4001 = pi39 & ~n4000;
  assign n4002 = ~pi38 & ~n4001;
  assign n4003 = ~n3978 & n4002;
  assign n4004 = ~n3987 & ~n3991;
  assign n4005 = ~pi216 & ~n4004;
  assign n4006 = n3937 & ~n4005;
  assign n4007 = ~n3935 & ~n4006;
  assign n4008 = ~pi215 & ~n4007;
  assign n4009 = ~n3930 & ~n4008;
  assign n4010 = ~n3471 & ~n4009;
  assign n4011 = pi299 & n4010;
  assign n4012 = ~n3985 & ~n4011;
  assign n4013 = pi38 & n4012;
  assign n4014 = ~pi100 & ~n4013;
  assign n4015 = ~n4003 & n4014;
  assign n4016 = ~pi262 & n3388;
  assign n4017 = ~n3592 & ~n3987;
  assign n4018 = ~n4016 & ~n4017;
  assign n4019 = n3992 & ~n4018;
  assign n4020 = ~pi216 & ~n4019;
  assign n4021 = n3937 & ~n4020;
  assign n4022 = ~n3935 & ~n4021;
  assign n4023 = ~pi215 & ~n4022;
  assign n4024 = ~n3930 & ~n4023;
  assign n4025 = pi299 & ~n4024;
  assign n4026 = n3181 & ~n3985;
  assign n4027 = ~n4025 & n4026;
  assign n4028 = ~n3181 & n4012;
  assign n4029 = pi100 & ~n4028;
  assign n4030 = ~n4027 & n4029;
  assign n4031 = ~n4015 & ~n4030;
  assign n4032 = ~pi87 & ~n4031;
  assign n4033 = ~n3207 & n4012;
  assign n4034 = n3207 & n4000;
  assign n4035 = ~n4033 & ~n4034;
  assign n4036 = pi87 & n4035;
  assign n4037 = ~pi75 & ~n4036;
  assign n4038 = ~n4032 & n4037;
  assign n4039 = pi75 & n4012;
  assign n4040 = ~pi92 & ~n4039;
  assign n4041 = ~n4038 & n4040;
  assign n4042 = n3230 & ~n4035;
  assign n4043 = ~n3230 & n4012;
  assign n4044 = pi92 & ~n4043;
  assign n4045 = ~n4042 & n4044;
  assign n4046 = n3265 & ~n4045;
  assign n4047 = ~n4041 & n4046;
  assign n4048 = ~n3265 & n4012;
  assign n4049 = ~pi55 & ~n4048;
  assign n4050 = ~n4047 & n4049;
  assign n4051 = n3268 & n3998;
  assign n4052 = ~n3268 & ~n4010;
  assign n4053 = pi55 & ~n4052;
  assign n4054 = ~n4051 & n4053;
  assign n4055 = ~pi56 & ~n4054;
  assign n4056 = ~n4050 & n4055;
  assign n4057 = n3280 & ~n3998;
  assign n4058 = ~n3280 & n4010;
  assign n4059 = pi56 & ~n4058;
  assign n4060 = ~n4057 & n4059;
  assign n4061 = ~pi62 & ~n4060;
  assign n4062 = ~n4056 & n4061;
  assign n4063 = n3431 & n3998;
  assign n4064 = ~n3431 & ~n4010;
  assign n4065 = pi62 & ~n4064;
  assign n4066 = ~n4063 & n4065;
  assign n4067 = n3429 & ~n4066;
  assign n4068 = ~n4062 & n4067;
  assign n4069 = ~n3429 & ~n4010;
  assign n4070 = ~pi249 & ~n4069;
  assign n4071 = ~n4068 & n4070;
  assign n4072 = pi262 & n3453;
  assign n4073 = ~pi172 & ~n4072;
  assign n4074 = ~pi262 & ~n3364;
  assign n4075 = pi262 & ~n3460;
  assign n4076 = pi172 & ~n4075;
  assign n4077 = ~n4074 & n4076;
  assign n4078 = ~n4073 & ~n4077;
  assign n4079 = ~pi228 & ~n4078;
  assign n4080 = ~pi216 & ~n3951;
  assign n4081 = ~n4079 & n4080;
  assign n4082 = n3937 & ~n4081;
  assign n4083 = ~n3935 & ~n4082;
  assign n4084 = ~pi215 & ~n4083;
  assign n4085 = n3931 & ~n4084;
  assign n4086 = n3976 & ~n4085;
  assign n4087 = ~n3989 & ~n3991;
  assign n4088 = ~pi216 & ~n4087;
  assign n4089 = n3937 & ~n4088;
  assign n4090 = ~n3935 & ~n4089;
  assign n4091 = ~pi215 & ~n4090;
  assign n4092 = ~n3930 & ~n4091;
  assign n4093 = pi299 & ~n4092;
  assign n4094 = ~n3984 & ~n4093;
  assign n4095 = pi39 & ~n4094;
  assign n4096 = ~pi38 & ~n4095;
  assign n4097 = ~n4086 & n4096;
  assign n4098 = pi299 & ~n4009;
  assign n4099 = ~n3984 & ~n4098;
  assign n4100 = pi38 & n4099;
  assign n4101 = ~pi100 & ~n4100;
  assign n4102 = ~n4097 & n4101;
  assign n4103 = ~n3991 & ~n4018;
  assign n4104 = ~pi216 & ~n4103;
  assign n4105 = n3937 & ~n4104;
  assign n4106 = ~n3935 & ~n4105;
  assign n4107 = ~pi215 & ~n4106;
  assign n4108 = ~n3930 & ~n4107;
  assign n4109 = pi299 & ~n4108;
  assign n4110 = n3181 & ~n3984;
  assign n4111 = ~n4109 & n4110;
  assign n4112 = ~n3181 & n4099;
  assign n4113 = pi100 & ~n4112;
  assign n4114 = ~n4111 & n4113;
  assign n4115 = ~n4102 & ~n4114;
  assign n4116 = ~pi87 & ~n4115;
  assign n4117 = ~n3207 & n4099;
  assign n4118 = n3207 & n4094;
  assign n4119 = ~n4117 & ~n4118;
  assign n4120 = pi87 & n4119;
  assign n4121 = ~pi75 & ~n4120;
  assign n4122 = ~n4116 & n4121;
  assign n4123 = pi75 & n4099;
  assign n4124 = ~pi92 & ~n4123;
  assign n4125 = ~n4122 & n4124;
  assign n4126 = n3230 & ~n4119;
  assign n4127 = ~n3230 & n4099;
  assign n4128 = pi92 & ~n4127;
  assign n4129 = ~n4126 & n4128;
  assign n4130 = n3265 & ~n4129;
  assign n4131 = ~n4125 & n4130;
  assign n4132 = ~n3265 & n4099;
  assign n4133 = ~pi55 & ~n4132;
  assign n4134 = ~n4131 & n4133;
  assign n4135 = n3268 & n4092;
  assign n4136 = ~n3268 & n4009;
  assign n4137 = pi55 & ~n4136;
  assign n4138 = ~n4135 & n4137;
  assign n4139 = ~pi56 & ~n4138;
  assign n4140 = ~n4134 & n4139;
  assign n4141 = n3280 & ~n4092;
  assign n4142 = ~n3280 & ~n4009;
  assign n4143 = pi56 & ~n4142;
  assign n4144 = ~n4141 & n4143;
  assign n4145 = ~pi62 & ~n4144;
  assign n4146 = ~n4140 & n4145;
  assign n4147 = n3431 & n4092;
  assign n4148 = ~n3431 & n4009;
  assign n4149 = pi62 & ~n4148;
  assign n4150 = ~n4147 & n4149;
  assign n4151 = n3429 & ~n4150;
  assign n4152 = ~n4146 & n4151;
  assign n4153 = ~n3429 & n4009;
  assign n4154 = pi249 & ~n4153;
  assign n4155 = ~n4152 & n4154;
  assign po157 = n4071 | n4155;
  assign n4157 = pi215 & pi1141;
  assign n4158 = pi299 & ~n4157;
  assign n4159 = ~pi935 & n2437;
  assign n4160 = ~pi1141 & ~n2437;
  assign n4161 = pi221 & ~n4160;
  assign n4162 = ~n4159 & n4161;
  assign n4163 = pi216 & pi270;
  assign n4164 = ~pi221 & ~n4163;
  assign n4165 = pi861 & n3460;
  assign n4166 = ~pi171 & ~n4165;
  assign n4167 = pi171 & n3453;
  assign n4168 = ~n4166 & ~n4167;
  assign n4169 = pi861 & ~n4168;
  assign n4170 = ~n3364 & n4166;
  assign n4171 = ~n4169 & ~n4170;
  assign n4172 = ~pi228 & ~n4171;
  assign n4173 = pi861 & ~n2449;
  assign n4174 = pi105 & ~n4173;
  assign n4175 = ~pi105 & pi171;
  assign n4176 = pi228 & ~n4175;
  assign n4177 = ~n4174 & n4176;
  assign n4178 = ~n3458 & n4177;
  assign n4179 = ~pi216 & ~n4178;
  assign n4180 = ~n4172 & n4179;
  assign n4181 = n4164 & ~n4180;
  assign n4182 = ~n4162 & ~n4181;
  assign n4183 = ~pi215 & ~n4182;
  assign n4184 = n4158 & ~n4183;
  assign n4185 = pi223 & pi1141;
  assign n4186 = ~pi299 & ~n4185;
  assign n4187 = ~pi935 & n3040;
  assign n4188 = ~pi1141 & ~n3040;
  assign n4189 = pi222 & ~n4188;
  assign n4190 = ~n4187 & n4189;
  assign n4191 = pi224 & pi270;
  assign n4192 = ~pi222 & ~n4191;
  assign n4193 = pi861 & n3441;
  assign n4194 = ~pi224 & ~n4193;
  assign n4195 = n4192 & ~n4194;
  assign n4196 = ~n4190 & ~n4195;
  assign n4197 = n4186 & n4196;
  assign n4198 = ~n3441 & n4192;
  assign n4199 = n4196 & ~n4198;
  assign n4200 = ~pi223 & ~n4199;
  assign n4201 = n4186 & ~n4200;
  assign n4202 = ~pi39 & ~n4201;
  assign n4203 = ~n4197 & n4202;
  assign n4204 = ~n4184 & n4203;
  assign n4205 = ~pi224 & ~n4173;
  assign n4206 = n4192 & ~n4205;
  assign n4207 = ~n4190 & ~n4206;
  assign n4208 = ~pi223 & ~n4207;
  assign n4209 = ~n4185 & ~n4208;
  assign n4210 = ~pi299 & ~n4209;
  assign n4211 = ~pi216 & ~n4177;
  assign n4212 = pi171 & ~n3095;
  assign n4213 = ~pi861 & n3095;
  assign n4214 = ~pi228 & ~n4213;
  assign n4215 = ~n4212 & n4214;
  assign n4216 = n4211 & ~n4215;
  assign n4217 = n4164 & ~n4216;
  assign n4218 = ~n4162 & ~n4217;
  assign n4219 = ~pi215 & ~n4218;
  assign n4220 = ~n4157 & ~n4219;
  assign n4221 = pi299 & ~n4220;
  assign n4222 = ~n4210 & ~n4221;
  assign n4223 = pi39 & ~n4222;
  assign n4224 = ~pi38 & ~n4223;
  assign n4225 = ~n4204 & n4224;
  assign n4226 = ~pi171 & ~pi228;
  assign n4227 = n4211 & ~n4226;
  assign n4228 = n4164 & ~n4227;
  assign n4229 = ~n4162 & ~n4228;
  assign n4230 = ~pi215 & ~n4229;
  assign n4231 = ~n4157 & ~n4230;
  assign n4232 = pi299 & ~n4231;
  assign n4233 = ~n4210 & ~n4232;
  assign n4234 = pi38 & n4233;
  assign n4235 = ~pi100 & ~n4234;
  assign n4236 = ~n4225 & n4235;
  assign n4237 = pi171 & ~n3388;
  assign n4238 = ~pi861 & n3388;
  assign n4239 = ~pi228 & ~n4238;
  assign n4240 = ~n4237 & n4239;
  assign n4241 = n4211 & ~n4240;
  assign n4242 = n4164 & ~n4241;
  assign n4243 = ~n4162 & ~n4242;
  assign n4244 = ~pi215 & ~n4243;
  assign n4245 = ~n4157 & ~n4244;
  assign n4246 = pi299 & ~n4245;
  assign n4247 = n3181 & ~n4210;
  assign n4248 = ~n4246 & n4247;
  assign n4249 = ~n3181 & n4233;
  assign n4250 = pi100 & ~n4249;
  assign n4251 = ~n4248 & n4250;
  assign n4252 = ~n4236 & ~n4251;
  assign n4253 = ~pi87 & ~n4252;
  assign n4254 = ~n3207 & n4233;
  assign n4255 = n3207 & n4222;
  assign n4256 = ~n4254 & ~n4255;
  assign n4257 = pi87 & n4256;
  assign n4258 = ~pi75 & ~n4257;
  assign n4259 = ~n4253 & n4258;
  assign n4260 = pi75 & n4233;
  assign n4261 = ~pi92 & ~n4260;
  assign n4262 = ~n4259 & n4261;
  assign n4263 = n3230 & ~n4256;
  assign n4264 = ~n3230 & n4233;
  assign n4265 = pi92 & ~n4264;
  assign n4266 = ~n4263 & n4265;
  assign n4267 = n3265 & ~n4266;
  assign n4268 = ~n4262 & n4267;
  assign n4269 = ~n3265 & n4233;
  assign n4270 = ~pi55 & ~n4269;
  assign n4271 = ~n4268 & n4270;
  assign n4272 = n3268 & n4220;
  assign n4273 = ~n3268 & n4231;
  assign n4274 = pi55 & ~n4273;
  assign n4275 = ~n4272 & n4274;
  assign n4276 = ~pi56 & ~n4275;
  assign n4277 = ~n4271 & n4276;
  assign n4278 = n3280 & ~n4220;
  assign n4279 = ~n3280 & ~n4231;
  assign n4280 = pi56 & ~n4279;
  assign n4281 = ~n4278 & n4280;
  assign n4282 = ~pi62 & ~n4281;
  assign n4283 = ~n4277 & n4282;
  assign n4284 = n3431 & n4220;
  assign n4285 = ~n3431 & n4231;
  assign n4286 = pi62 & ~n4285;
  assign n4287 = ~n4284 & n4286;
  assign n4288 = ~pi241 & n3429;
  assign n4289 = ~n4287 & n4288;
  assign n4290 = ~n4283 & n4289;
  assign n4291 = ~pi861 & n3453;
  assign n4292 = ~pi171 & ~n4291;
  assign n4293 = pi861 & ~n3364;
  assign n4294 = ~pi861 & ~n3460;
  assign n4295 = pi171 & ~n4294;
  assign n4296 = ~n4293 & n4295;
  assign n4297 = ~n4292 & ~n4296;
  assign n4298 = ~pi228 & ~n4297;
  assign n4299 = ~n3845 & n4211;
  assign n4300 = ~n4298 & n4299;
  assign n4301 = n4164 & ~n4300;
  assign n4302 = ~n4162 & ~n4301;
  assign n4303 = ~pi215 & ~n4302;
  assign n4304 = n4158 & ~n4303;
  assign n4305 = n4202 & ~n4304;
  assign n4306 = ~n3476 & ~n4210;
  assign n4307 = ~n3470 & n4211;
  assign n4308 = ~n4215 & n4307;
  assign n4309 = n4164 & ~n4308;
  assign n4310 = ~n4162 & ~n4309;
  assign n4311 = ~pi215 & ~n4310;
  assign n4312 = ~n4157 & ~n4311;
  assign n4313 = pi299 & ~n4312;
  assign n4314 = n4306 & ~n4313;
  assign n4315 = pi39 & ~n4314;
  assign n4316 = ~pi38 & ~n4315;
  assign n4317 = ~n4305 & n4316;
  assign n4318 = n3584 & ~n4163;
  assign n4319 = n4231 & ~n4318;
  assign n4320 = pi299 & ~n4319;
  assign n4321 = n4306 & ~n4320;
  assign n4322 = pi38 & n4321;
  assign n4323 = ~pi100 & ~n4322;
  assign n4324 = ~n4317 & n4323;
  assign n4325 = ~n4240 & n4307;
  assign n4326 = n4164 & ~n4325;
  assign n4327 = ~n4162 & ~n4326;
  assign n4328 = ~pi215 & ~n4327;
  assign n4329 = ~n4157 & ~n4328;
  assign n4330 = pi299 & ~n4329;
  assign n4331 = n3181 & n4306;
  assign n4332 = ~n4330 & n4331;
  assign n4333 = ~n3181 & n4321;
  assign n4334 = pi100 & ~n4333;
  assign n4335 = ~n4332 & n4334;
  assign n4336 = ~n4324 & ~n4335;
  assign n4337 = ~pi87 & ~n4336;
  assign n4338 = ~n3207 & n4321;
  assign n4339 = n3207 & n4314;
  assign n4340 = ~n4338 & ~n4339;
  assign n4341 = pi87 & n4340;
  assign n4342 = ~pi75 & ~n4341;
  assign n4343 = ~n4337 & n4342;
  assign n4344 = pi75 & n4321;
  assign n4345 = ~pi92 & ~n4344;
  assign n4346 = ~n4343 & n4345;
  assign n4347 = n3230 & ~n4340;
  assign n4348 = ~n3230 & n4321;
  assign n4349 = pi92 & ~n4348;
  assign n4350 = ~n4347 & n4349;
  assign n4351 = n3265 & ~n4350;
  assign n4352 = ~n4346 & n4351;
  assign n4353 = ~n3265 & n4321;
  assign n4354 = ~pi55 & ~n4353;
  assign n4355 = ~n4352 & n4354;
  assign n4356 = n3268 & n4312;
  assign n4357 = ~n3268 & n4319;
  assign n4358 = pi55 & ~n4357;
  assign n4359 = ~n4356 & n4358;
  assign n4360 = ~pi56 & ~n4359;
  assign n4361 = ~n4355 & n4360;
  assign n4362 = n3280 & ~n4312;
  assign n4363 = ~n3280 & ~n4319;
  assign n4364 = pi56 & ~n4363;
  assign n4365 = ~n4362 & n4364;
  assign n4366 = ~pi62 & ~n4365;
  assign n4367 = ~n4361 & n4366;
  assign n4368 = n3431 & n4312;
  assign n4369 = ~n3431 & n4319;
  assign n4370 = pi62 & ~n4369;
  assign n4371 = ~n4368 & n4370;
  assign n4372 = pi241 & n3429;
  assign n4373 = ~n4371 & n4372;
  assign n4374 = ~n4367 & n4373;
  assign n4375 = pi241 & n4318;
  assign n4376 = ~n3429 & ~n4375;
  assign n4377 = n4231 & n4376;
  assign n4378 = ~n4374 & ~n4377;
  assign po158 = ~n4290 & n4378;
  assign n4380 = pi215 & pi1140;
  assign n4381 = pi299 & ~n4380;
  assign n4382 = ~pi921 & n2437;
  assign n4383 = ~pi1140 & ~n2437;
  assign n4384 = pi221 & ~n4383;
  assign n4385 = ~n4382 & n4384;
  assign n4386 = pi216 & pi282;
  assign n4387 = ~pi221 & ~n4386;
  assign n4388 = pi869 & n3460;
  assign n4389 = ~pi170 & ~n4388;
  assign n4390 = pi170 & n3453;
  assign n4391 = ~n4389 & ~n4390;
  assign n4392 = pi869 & ~n4391;
  assign n4393 = ~n3364 & n4389;
  assign n4394 = ~n4392 & ~n4393;
  assign n4395 = ~pi228 & ~n4394;
  assign n4396 = pi869 & ~n2449;
  assign n4397 = pi105 & ~n4396;
  assign n4398 = ~pi105 & pi170;
  assign n4399 = pi228 & ~n4398;
  assign n4400 = ~n4397 & n4399;
  assign n4401 = ~n3458 & n4400;
  assign n4402 = ~pi216 & ~n4401;
  assign n4403 = ~n4395 & n4402;
  assign n4404 = n4387 & ~n4403;
  assign n4405 = ~n4385 & ~n4404;
  assign n4406 = ~pi215 & ~n4405;
  assign n4407 = n4381 & ~n4406;
  assign n4408 = pi223 & pi1140;
  assign n4409 = ~pi299 & ~n4408;
  assign n4410 = ~pi921 & n3040;
  assign n4411 = ~pi1140 & ~n3040;
  assign n4412 = pi222 & ~n4411;
  assign n4413 = ~n4410 & n4412;
  assign n4414 = pi224 & pi282;
  assign n4415 = ~pi222 & ~n4414;
  assign n4416 = pi869 & n3441;
  assign n4417 = ~pi224 & ~n4416;
  assign n4418 = n4415 & ~n4417;
  assign n4419 = ~n4413 & ~n4418;
  assign n4420 = n4409 & n4419;
  assign n4421 = ~n3441 & n4415;
  assign n4422 = n4419 & ~n4421;
  assign n4423 = ~pi223 & ~n4422;
  assign n4424 = n4409 & ~n4423;
  assign n4425 = ~pi39 & ~n4424;
  assign n4426 = ~n4420 & n4425;
  assign n4427 = ~n4407 & n4426;
  assign n4428 = ~pi224 & ~n4396;
  assign n4429 = n4415 & ~n4428;
  assign n4430 = ~n4413 & ~n4429;
  assign n4431 = ~pi223 & ~n4430;
  assign n4432 = ~n4408 & ~n4431;
  assign n4433 = ~pi299 & ~n4432;
  assign n4434 = ~pi216 & ~n4400;
  assign n4435 = pi170 & ~n3095;
  assign n4436 = ~pi869 & n3095;
  assign n4437 = ~pi228 & ~n4436;
  assign n4438 = ~n4435 & n4437;
  assign n4439 = n4434 & ~n4438;
  assign n4440 = n4387 & ~n4439;
  assign n4441 = ~n4385 & ~n4440;
  assign n4442 = ~pi215 & ~n4441;
  assign n4443 = ~n4380 & ~n4442;
  assign n4444 = pi299 & ~n4443;
  assign n4445 = ~n4433 & ~n4444;
  assign n4446 = pi39 & ~n4445;
  assign n4447 = ~pi38 & ~n4446;
  assign n4448 = ~n4427 & n4447;
  assign n4449 = ~pi170 & ~pi228;
  assign n4450 = n4434 & ~n4449;
  assign n4451 = n4387 & ~n4450;
  assign n4452 = ~n4385 & ~n4451;
  assign n4453 = ~pi215 & ~n4452;
  assign n4454 = ~n4380 & ~n4453;
  assign n4455 = pi299 & ~n4454;
  assign n4456 = ~n4433 & ~n4455;
  assign n4457 = pi38 & n4456;
  assign n4458 = ~pi100 & ~n4457;
  assign n4459 = ~n4448 & n4458;
  assign n4460 = pi170 & ~n3388;
  assign n4461 = ~pi869 & n3388;
  assign n4462 = ~pi228 & ~n4461;
  assign n4463 = ~n4460 & n4462;
  assign n4464 = n4434 & ~n4463;
  assign n4465 = n4387 & ~n4464;
  assign n4466 = ~n4385 & ~n4465;
  assign n4467 = ~pi215 & ~n4466;
  assign n4468 = ~n4380 & ~n4467;
  assign n4469 = pi299 & ~n4468;
  assign n4470 = n3181 & ~n4433;
  assign n4471 = ~n4469 & n4470;
  assign n4472 = ~n3181 & n4456;
  assign n4473 = pi100 & ~n4472;
  assign n4474 = ~n4471 & n4473;
  assign n4475 = ~n4459 & ~n4474;
  assign n4476 = ~pi87 & ~n4475;
  assign n4477 = ~n3207 & n4456;
  assign n4478 = n3207 & n4445;
  assign n4479 = ~n4477 & ~n4478;
  assign n4480 = pi87 & n4479;
  assign n4481 = ~pi75 & ~n4480;
  assign n4482 = ~n4476 & n4481;
  assign n4483 = pi75 & n4456;
  assign n4484 = ~pi92 & ~n4483;
  assign n4485 = ~n4482 & n4484;
  assign n4486 = n3230 & ~n4479;
  assign n4487 = ~n3230 & n4456;
  assign n4488 = pi92 & ~n4487;
  assign n4489 = ~n4486 & n4488;
  assign n4490 = n3265 & ~n4489;
  assign n4491 = ~n4485 & n4490;
  assign n4492 = ~n3265 & n4456;
  assign n4493 = ~pi55 & ~n4492;
  assign n4494 = ~n4491 & n4493;
  assign n4495 = n3268 & n4443;
  assign n4496 = ~n3268 & n4454;
  assign n4497 = pi55 & ~n4496;
  assign n4498 = ~n4495 & n4497;
  assign n4499 = ~pi56 & ~n4498;
  assign n4500 = ~n4494 & n4499;
  assign n4501 = n3280 & ~n4443;
  assign n4502 = ~n3280 & ~n4454;
  assign n4503 = pi56 & ~n4502;
  assign n4504 = ~n4501 & n4503;
  assign n4505 = ~pi62 & ~n4504;
  assign n4506 = ~n4500 & n4505;
  assign n4507 = n3431 & n4443;
  assign n4508 = ~n3431 & n4454;
  assign n4509 = pi62 & ~n4508;
  assign n4510 = ~n4507 & n4509;
  assign n4511 = ~pi248 & n3429;
  assign n4512 = ~n4510 & n4511;
  assign n4513 = ~n4506 & n4512;
  assign n4514 = ~pi869 & n3453;
  assign n4515 = ~pi170 & ~n4514;
  assign n4516 = pi869 & ~n3364;
  assign n4517 = ~pi869 & ~n3460;
  assign n4518 = pi170 & ~n4517;
  assign n4519 = ~n4516 & n4518;
  assign n4520 = ~n4515 & ~n4519;
  assign n4521 = ~pi228 & ~n4520;
  assign n4522 = ~n3845 & n4434;
  assign n4523 = ~n4521 & n4522;
  assign n4524 = n4387 & ~n4523;
  assign n4525 = ~n4385 & ~n4524;
  assign n4526 = ~pi215 & ~n4525;
  assign n4527 = n4381 & ~n4526;
  assign n4528 = n4425 & ~n4527;
  assign n4529 = ~n3476 & ~n4433;
  assign n4530 = ~n3470 & n4434;
  assign n4531 = ~n4438 & n4530;
  assign n4532 = n4387 & ~n4531;
  assign n4533 = ~n4385 & ~n4532;
  assign n4534 = ~pi215 & ~n4533;
  assign n4535 = ~n4380 & ~n4534;
  assign n4536 = pi299 & ~n4535;
  assign n4537 = n4529 & ~n4536;
  assign n4538 = pi39 & ~n4537;
  assign n4539 = ~pi38 & ~n4538;
  assign n4540 = ~n4528 & n4539;
  assign n4541 = n3584 & ~n4386;
  assign n4542 = n4454 & ~n4541;
  assign n4543 = pi299 & ~n4542;
  assign n4544 = n4529 & ~n4543;
  assign n4545 = pi38 & n4544;
  assign n4546 = ~pi100 & ~n4545;
  assign n4547 = ~n4540 & n4546;
  assign n4548 = ~n4463 & n4530;
  assign n4549 = n4387 & ~n4548;
  assign n4550 = ~n4385 & ~n4549;
  assign n4551 = ~pi215 & ~n4550;
  assign n4552 = ~n4380 & ~n4551;
  assign n4553 = pi299 & ~n4552;
  assign n4554 = n3181 & n4529;
  assign n4555 = ~n4553 & n4554;
  assign n4556 = ~n3181 & n4544;
  assign n4557 = pi100 & ~n4556;
  assign n4558 = ~n4555 & n4557;
  assign n4559 = ~n4547 & ~n4558;
  assign n4560 = ~pi87 & ~n4559;
  assign n4561 = ~n3207 & n4544;
  assign n4562 = n3207 & n4537;
  assign n4563 = ~n4561 & ~n4562;
  assign n4564 = pi87 & n4563;
  assign n4565 = ~pi75 & ~n4564;
  assign n4566 = ~n4560 & n4565;
  assign n4567 = pi75 & n4544;
  assign n4568 = ~pi92 & ~n4567;
  assign n4569 = ~n4566 & n4568;
  assign n4570 = n3230 & ~n4563;
  assign n4571 = ~n3230 & n4544;
  assign n4572 = pi92 & ~n4571;
  assign n4573 = ~n4570 & n4572;
  assign n4574 = n3265 & ~n4573;
  assign n4575 = ~n4569 & n4574;
  assign n4576 = ~n3265 & n4544;
  assign n4577 = ~pi55 & ~n4576;
  assign n4578 = ~n4575 & n4577;
  assign n4579 = n3268 & n4535;
  assign n4580 = ~n3268 & n4542;
  assign n4581 = pi55 & ~n4580;
  assign n4582 = ~n4579 & n4581;
  assign n4583 = ~pi56 & ~n4582;
  assign n4584 = ~n4578 & n4583;
  assign n4585 = n3280 & ~n4535;
  assign n4586 = ~n3280 & ~n4542;
  assign n4587 = pi56 & ~n4586;
  assign n4588 = ~n4585 & n4587;
  assign n4589 = ~pi62 & ~n4588;
  assign n4590 = ~n4584 & n4589;
  assign n4591 = n3431 & n4535;
  assign n4592 = ~n3431 & n4542;
  assign n4593 = pi62 & ~n4592;
  assign n4594 = ~n4591 & n4593;
  assign n4595 = pi248 & n3429;
  assign n4596 = ~n4594 & n4595;
  assign n4597 = ~n4590 & n4596;
  assign n4598 = pi248 & n4541;
  assign n4599 = ~n3429 & ~n4598;
  assign n4600 = n4454 & n4599;
  assign n4601 = ~n4597 & ~n4600;
  assign po159 = ~n4513 & n4601;
  assign n4603 = pi215 & pi1139;
  assign n4604 = ~pi148 & ~pi215;
  assign n4605 = pi216 & ~pi1139;
  assign n4606 = ~pi833 & pi1139;
  assign n4607 = pi833 & pi920;
  assign n4608 = ~pi216 & ~n4607;
  assign n4609 = ~n4606 & n4608;
  assign n4610 = pi221 & ~n4609;
  assign n4611 = ~n4605 & n4610;
  assign n4612 = pi216 & pi281;
  assign n4613 = ~pi221 & ~n4612;
  assign n4614 = ~n3126 & ~n3321;
  assign n4615 = pi862 & ~n3470;
  assign n4616 = ~pi216 & ~n4615;
  assign n4617 = ~n4614 & n4616;
  assign n4618 = n4613 & ~n4617;
  assign n4619 = ~n4611 & ~n4618;
  assign n4620 = ~n3126 & ~n3592;
  assign n4621 = n4613 & n4620;
  assign n4622 = n4619 & ~n4621;
  assign n4623 = n4604 & ~n4622;
  assign n4624 = ~n4603 & ~n4623;
  assign n4625 = ~pi216 & ~n4611;
  assign n4626 = n3594 & n4625;
  assign n4627 = ~pi216 & ~pi862;
  assign n4628 = ~n3321 & ~n3593;
  assign n4629 = n4627 & ~n4628;
  assign n4630 = n4613 & ~n4629;
  assign n4631 = ~n4611 & ~n4630;
  assign n4632 = pi148 & ~pi215;
  assign n4633 = ~n4631 & n4632;
  assign n4634 = ~n4626 & n4633;
  assign n4635 = n4624 & ~n4634;
  assign n4636 = pi299 & ~n4635;
  assign n4637 = ~pi920 & n3040;
  assign n4638 = ~pi1139 & ~n3040;
  assign n4639 = pi222 & ~n4638;
  assign n4640 = ~n4637 & n4639;
  assign n4641 = pi223 & pi1139;
  assign n4642 = ~pi224 & ~n4641;
  assign n4643 = ~n4640 & n4642;
  assign n4644 = ~pi862 & n4643;
  assign n4645 = pi224 & pi281;
  assign n4646 = ~pi222 & ~n4645;
  assign n4647 = ~n4640 & ~n4646;
  assign n4648 = ~pi223 & ~n4647;
  assign n4649 = ~n4641 & ~n4648;
  assign n4650 = ~pi299 & ~n4649;
  assign n4651 = ~n4644 & n4650;
  assign n4652 = ~n3856 & n4651;
  assign n4653 = n3181 & ~n4652;
  assign n4654 = ~n4636 & n4653;
  assign n4655 = n3593 & n4627;
  assign n4656 = n4613 & ~n4655;
  assign n4657 = ~n4611 & ~n4656;
  assign n4658 = pi148 & ~n3126;
  assign n4659 = n4625 & n4658;
  assign n4660 = ~pi215 & ~n4659;
  assign n4661 = ~n4657 & n4660;
  assign n4662 = ~n4603 & ~n4661;
  assign n4663 = ~n3471 & ~n4662;
  assign n4664 = pi299 & n4663;
  assign n4665 = ~n4652 & ~n4664;
  assign n4666 = ~n3181 & n4665;
  assign n4667 = pi100 & ~n4666;
  assign n4668 = ~n4654 & n4667;
  assign n4669 = ~pi228 & n3364;
  assign n4670 = ~n3126 & ~n4669;
  assign n4671 = ~pi862 & n4670;
  assign n4672 = pi862 & ~n3462;
  assign n4673 = ~pi216 & ~n4672;
  assign n4674 = ~n4671 & n4673;
  assign n4675 = n4613 & ~n4674;
  assign n4676 = ~n4611 & ~n4675;
  assign n4677 = n4604 & ~n4676;
  assign n4678 = ~n3456 & n4627;
  assign n4679 = n4613 & ~n4678;
  assign n4680 = ~n4611 & ~n4679;
  assign n4681 = n3456 & n4625;
  assign n4682 = n4632 & ~n4681;
  assign n4683 = ~n4680 & n4682;
  assign n4684 = pi299 & ~n4603;
  assign n4685 = ~n4683 & n4684;
  assign n4686 = ~n4677 & n4685;
  assign n4687 = ~n3441 & n4643;
  assign n4688 = ~n4644 & ~n4649;
  assign n4689 = ~n4687 & n4688;
  assign n4690 = ~pi299 & ~n4689;
  assign n4691 = ~pi39 & ~n4690;
  assign n4692 = ~n4686 & n4691;
  assign n4693 = n4604 & ~n4619;
  assign n4694 = n4625 & n4628;
  assign n4695 = n4633 & ~n4694;
  assign n4696 = ~n4603 & ~n4695;
  assign n4697 = ~n4693 & n4696;
  assign n4698 = pi299 & ~n4697;
  assign n4699 = ~n4652 & ~n4698;
  assign n4700 = pi39 & ~n4699;
  assign n4701 = ~pi38 & ~n4700;
  assign n4702 = ~n4692 & n4701;
  assign n4703 = pi38 & n4665;
  assign n4704 = ~pi100 & ~n4703;
  assign n4705 = ~n4702 & n4704;
  assign n4706 = ~n4668 & ~n4705;
  assign n4707 = ~pi87 & ~n4706;
  assign n4708 = ~n3207 & n4665;
  assign n4709 = n3207 & n4699;
  assign n4710 = ~n4708 & ~n4709;
  assign n4711 = pi87 & n4710;
  assign n4712 = ~pi75 & ~n4711;
  assign n4713 = ~n4707 & n4712;
  assign n4714 = pi75 & n4665;
  assign n4715 = ~pi92 & ~n4714;
  assign n4716 = ~n4713 & n4715;
  assign n4717 = n3230 & ~n4710;
  assign n4718 = ~n3230 & n4665;
  assign n4719 = pi92 & ~n4718;
  assign n4720 = ~n4717 & n4719;
  assign n4721 = n3265 & ~n4720;
  assign n4722 = ~n4716 & n4721;
  assign n4723 = ~n3265 & n4665;
  assign n4724 = ~pi55 & ~n4723;
  assign n4725 = ~n4722 & n4724;
  assign n4726 = n3268 & n4697;
  assign n4727 = ~n3268 & ~n4663;
  assign n4728 = pi55 & ~n4727;
  assign n4729 = ~n4726 & n4728;
  assign n4730 = ~pi56 & ~n4729;
  assign n4731 = ~n4725 & n4730;
  assign n4732 = n3280 & ~n4697;
  assign n4733 = ~n3280 & n4663;
  assign n4734 = pi56 & ~n4733;
  assign n4735 = ~n4732 & n4734;
  assign n4736 = ~pi62 & ~n4735;
  assign n4737 = ~n4731 & n4736;
  assign n4738 = n3431 & n4697;
  assign n4739 = ~n3431 & ~n4663;
  assign n4740 = pi62 & ~n4739;
  assign n4741 = ~n4738 & n4740;
  assign n4742 = n3429 & ~n4741;
  assign n4743 = ~n4737 & n4742;
  assign n4744 = ~n3429 & ~n4663;
  assign n4745 = ~pi247 & ~n4744;
  assign n4746 = ~n4743 & n4745;
  assign n4747 = n3594 & n4613;
  assign n4748 = n4631 & ~n4747;
  assign n4749 = n4604 & ~n4748;
  assign n4750 = n4620 & n4625;
  assign n4751 = n4633 & ~n4750;
  assign n4752 = ~n4603 & ~n4751;
  assign n4753 = ~n4749 & n4752;
  assign n4754 = pi299 & ~n4753;
  assign n4755 = ~n3476 & ~n4651;
  assign n4756 = n3181 & n4755;
  assign n4757 = ~n4754 & n4756;
  assign n4758 = pi299 & ~n4662;
  assign n4759 = n4755 & ~n4758;
  assign n4760 = ~n3181 & n4759;
  assign n4761 = pi100 & ~n4760;
  assign n4762 = ~n4757 & n4761;
  assign n4763 = n3441 & n4644;
  assign n4764 = n4650 & ~n4763;
  assign n4765 = pi862 & ~n4670;
  assign n4766 = ~pi862 & n3462;
  assign n4767 = ~pi216 & ~n4766;
  assign n4768 = ~n4765 & n4767;
  assign n4769 = n4613 & ~n4768;
  assign n4770 = ~n4611 & ~n4769;
  assign n4771 = n4632 & ~n4770;
  assign n4772 = n4604 & ~n4680;
  assign n4773 = ~n4603 & ~n4772;
  assign n4774 = ~n4771 & n4773;
  assign n4775 = pi299 & ~n4774;
  assign n4776 = ~n4764 & ~n4775;
  assign n4777 = ~pi39 & ~n4776;
  assign n4778 = ~n4631 & n4660;
  assign n4779 = n4696 & ~n4778;
  assign n4780 = pi299 & ~n4779;
  assign n4781 = n4755 & ~n4780;
  assign n4782 = pi39 & ~n4781;
  assign n4783 = ~pi38 & ~n4782;
  assign n4784 = ~n4777 & n4783;
  assign n4785 = pi38 & n4759;
  assign n4786 = ~pi100 & ~n4785;
  assign n4787 = ~n4784 & n4786;
  assign n4788 = ~n4762 & ~n4787;
  assign n4789 = ~pi87 & ~n4788;
  assign n4790 = ~n3207 & n4759;
  assign n4791 = n3207 & n4781;
  assign n4792 = ~n4790 & ~n4791;
  assign n4793 = pi87 & n4792;
  assign n4794 = ~pi75 & ~n4793;
  assign n4795 = ~n4789 & n4794;
  assign n4796 = pi75 & n4759;
  assign n4797 = ~pi92 & ~n4796;
  assign n4798 = ~n4795 & n4797;
  assign n4799 = n3230 & ~n4792;
  assign n4800 = ~n3230 & n4759;
  assign n4801 = pi92 & ~n4800;
  assign n4802 = ~n4799 & n4801;
  assign n4803 = n3265 & ~n4802;
  assign n4804 = ~n4798 & n4803;
  assign n4805 = ~n3265 & n4759;
  assign n4806 = ~pi55 & ~n4805;
  assign n4807 = ~n4804 & n4806;
  assign n4808 = n3268 & n4779;
  assign n4809 = ~n3268 & n4662;
  assign n4810 = pi55 & ~n4809;
  assign n4811 = ~n4808 & n4810;
  assign n4812 = ~pi56 & ~n4811;
  assign n4813 = ~n4807 & n4812;
  assign n4814 = n3280 & ~n4779;
  assign n4815 = ~n3280 & ~n4662;
  assign n4816 = pi56 & ~n4815;
  assign n4817 = ~n4814 & n4816;
  assign n4818 = ~pi62 & ~n4817;
  assign n4819 = ~n4813 & n4818;
  assign n4820 = n3431 & n4779;
  assign n4821 = ~n3431 & n4662;
  assign n4822 = pi62 & ~n4821;
  assign n4823 = ~n4820 & n4822;
  assign n4824 = n3429 & ~n4823;
  assign n4825 = ~n4819 & n4824;
  assign n4826 = ~n3429 & n4662;
  assign n4827 = pi247 & ~n4826;
  assign n4828 = ~n4825 & n4827;
  assign po160 = n4746 | n4828;
  assign n4830 = pi215 & pi1138;
  assign n4831 = pi299 & ~n4830;
  assign n4832 = ~pi940 & n2437;
  assign n4833 = ~pi1138 & ~n2437;
  assign n4834 = pi221 & ~n4833;
  assign n4835 = ~n4832 & n4834;
  assign n4836 = pi216 & pi269;
  assign n4837 = ~pi221 & ~n4836;
  assign n4838 = pi877 & n3460;
  assign n4839 = ~pi169 & ~n4838;
  assign n4840 = pi169 & n3453;
  assign n4841 = ~n4839 & ~n4840;
  assign n4842 = pi877 & ~n4841;
  assign n4843 = ~n3364 & n4839;
  assign n4844 = ~n4842 & ~n4843;
  assign n4845 = ~pi228 & ~n4844;
  assign n4846 = pi877 & ~n2449;
  assign n4847 = pi105 & ~n4846;
  assign n4848 = ~pi105 & pi169;
  assign n4849 = pi228 & ~n4848;
  assign n4850 = ~n4847 & n4849;
  assign n4851 = ~n3458 & n4850;
  assign n4852 = ~pi216 & ~n4851;
  assign n4853 = ~n4845 & n4852;
  assign n4854 = n4837 & ~n4853;
  assign n4855 = ~n4835 & ~n4854;
  assign n4856 = ~pi215 & ~n4855;
  assign n4857 = n4831 & ~n4856;
  assign n4858 = pi223 & pi1138;
  assign n4859 = ~pi299 & ~n4858;
  assign n4860 = ~pi940 & n3040;
  assign n4861 = ~pi1138 & ~n3040;
  assign n4862 = pi222 & ~n4861;
  assign n4863 = ~n4860 & n4862;
  assign n4864 = pi224 & pi269;
  assign n4865 = ~pi222 & ~n4864;
  assign n4866 = pi877 & n3441;
  assign n4867 = ~pi224 & ~n4866;
  assign n4868 = n4865 & ~n4867;
  assign n4869 = ~n4863 & ~n4868;
  assign n4870 = n4859 & n4869;
  assign n4871 = ~n3441 & n4865;
  assign n4872 = n4869 & ~n4871;
  assign n4873 = ~pi223 & ~n4872;
  assign n4874 = n4859 & ~n4873;
  assign n4875 = ~pi39 & ~n4874;
  assign n4876 = ~n4870 & n4875;
  assign n4877 = ~n4857 & n4876;
  assign n4878 = ~pi224 & ~n4846;
  assign n4879 = n4865 & ~n4878;
  assign n4880 = ~n4863 & ~n4879;
  assign n4881 = ~pi223 & ~n4880;
  assign n4882 = ~n4858 & ~n4881;
  assign n4883 = ~pi299 & ~n4882;
  assign n4884 = ~pi216 & ~n4850;
  assign n4885 = pi169 & ~n3095;
  assign n4886 = ~pi877 & n3095;
  assign n4887 = ~pi228 & ~n4886;
  assign n4888 = ~n4885 & n4887;
  assign n4889 = n4884 & ~n4888;
  assign n4890 = n4837 & ~n4889;
  assign n4891 = ~n4835 & ~n4890;
  assign n4892 = ~pi215 & ~n4891;
  assign n4893 = ~n4830 & ~n4892;
  assign n4894 = pi299 & ~n4893;
  assign n4895 = ~n4883 & ~n4894;
  assign n4896 = pi39 & ~n4895;
  assign n4897 = ~pi38 & ~n4896;
  assign n4898 = ~n4877 & n4897;
  assign n4899 = ~pi169 & ~pi228;
  assign n4900 = n4884 & ~n4899;
  assign n4901 = n4837 & ~n4900;
  assign n4902 = ~n4835 & ~n4901;
  assign n4903 = ~pi215 & ~n4902;
  assign n4904 = ~n4830 & ~n4903;
  assign n4905 = pi299 & ~n4904;
  assign n4906 = ~n4883 & ~n4905;
  assign n4907 = pi38 & n4906;
  assign n4908 = ~pi100 & ~n4907;
  assign n4909 = ~n4898 & n4908;
  assign n4910 = pi169 & ~n3388;
  assign n4911 = ~pi877 & n3388;
  assign n4912 = ~pi228 & ~n4911;
  assign n4913 = ~n4910 & n4912;
  assign n4914 = n4884 & ~n4913;
  assign n4915 = n4837 & ~n4914;
  assign n4916 = ~n4835 & ~n4915;
  assign n4917 = ~pi215 & ~n4916;
  assign n4918 = ~n4830 & ~n4917;
  assign n4919 = pi299 & ~n4918;
  assign n4920 = n3181 & ~n4883;
  assign n4921 = ~n4919 & n4920;
  assign n4922 = ~n3181 & n4906;
  assign n4923 = pi100 & ~n4922;
  assign n4924 = ~n4921 & n4923;
  assign n4925 = ~n4909 & ~n4924;
  assign n4926 = ~pi87 & ~n4925;
  assign n4927 = ~n3207 & n4906;
  assign n4928 = n3207 & n4895;
  assign n4929 = ~n4927 & ~n4928;
  assign n4930 = pi87 & n4929;
  assign n4931 = ~pi75 & ~n4930;
  assign n4932 = ~n4926 & n4931;
  assign n4933 = pi75 & n4906;
  assign n4934 = ~pi92 & ~n4933;
  assign n4935 = ~n4932 & n4934;
  assign n4936 = n3230 & ~n4929;
  assign n4937 = ~n3230 & n4906;
  assign n4938 = pi92 & ~n4937;
  assign n4939 = ~n4936 & n4938;
  assign n4940 = n3265 & ~n4939;
  assign n4941 = ~n4935 & n4940;
  assign n4942 = ~n3265 & n4906;
  assign n4943 = ~pi55 & ~n4942;
  assign n4944 = ~n4941 & n4943;
  assign n4945 = n3268 & n4893;
  assign n4946 = ~n3268 & n4904;
  assign n4947 = pi55 & ~n4946;
  assign n4948 = ~n4945 & n4947;
  assign n4949 = ~pi56 & ~n4948;
  assign n4950 = ~n4944 & n4949;
  assign n4951 = n3280 & ~n4893;
  assign n4952 = ~n3280 & ~n4904;
  assign n4953 = pi56 & ~n4952;
  assign n4954 = ~n4951 & n4953;
  assign n4955 = ~pi62 & ~n4954;
  assign n4956 = ~n4950 & n4955;
  assign n4957 = n3431 & n4893;
  assign n4958 = ~n3431 & n4904;
  assign n4959 = pi62 & ~n4958;
  assign n4960 = ~n4957 & n4959;
  assign n4961 = ~pi246 & n3429;
  assign n4962 = ~n4960 & n4961;
  assign n4963 = ~n4956 & n4962;
  assign n4964 = ~pi877 & n3453;
  assign n4965 = ~pi169 & ~n4964;
  assign n4966 = pi877 & ~n3364;
  assign n4967 = ~pi877 & ~n3460;
  assign n4968 = pi169 & ~n4967;
  assign n4969 = ~n4966 & n4968;
  assign n4970 = ~n4965 & ~n4969;
  assign n4971 = ~pi228 & ~n4970;
  assign n4972 = ~n3845 & n4884;
  assign n4973 = ~n4971 & n4972;
  assign n4974 = n4837 & ~n4973;
  assign n4975 = ~n4835 & ~n4974;
  assign n4976 = ~pi215 & ~n4975;
  assign n4977 = n4831 & ~n4976;
  assign n4978 = n4875 & ~n4977;
  assign n4979 = ~n3476 & ~n4883;
  assign n4980 = ~n3470 & n4884;
  assign n4981 = ~n4888 & n4980;
  assign n4982 = n4837 & ~n4981;
  assign n4983 = ~n4835 & ~n4982;
  assign n4984 = ~pi215 & ~n4983;
  assign n4985 = ~n4830 & ~n4984;
  assign n4986 = pi299 & ~n4985;
  assign n4987 = n4979 & ~n4986;
  assign n4988 = pi39 & ~n4987;
  assign n4989 = ~pi38 & ~n4988;
  assign n4990 = ~n4978 & n4989;
  assign n4991 = n3584 & ~n4836;
  assign n4992 = n4904 & ~n4991;
  assign n4993 = pi299 & ~n4992;
  assign n4994 = n4979 & ~n4993;
  assign n4995 = pi38 & n4994;
  assign n4996 = ~pi100 & ~n4995;
  assign n4997 = ~n4990 & n4996;
  assign n4998 = ~n4913 & n4980;
  assign n4999 = n4837 & ~n4998;
  assign n5000 = ~n4835 & ~n4999;
  assign n5001 = ~pi215 & ~n5000;
  assign n5002 = ~n4830 & ~n5001;
  assign n5003 = pi299 & ~n5002;
  assign n5004 = n3181 & n4979;
  assign n5005 = ~n5003 & n5004;
  assign n5006 = ~n3181 & n4994;
  assign n5007 = pi100 & ~n5006;
  assign n5008 = ~n5005 & n5007;
  assign n5009 = ~n4997 & ~n5008;
  assign n5010 = ~pi87 & ~n5009;
  assign n5011 = ~n3207 & n4994;
  assign n5012 = n3207 & n4987;
  assign n5013 = ~n5011 & ~n5012;
  assign n5014 = pi87 & n5013;
  assign n5015 = ~pi75 & ~n5014;
  assign n5016 = ~n5010 & n5015;
  assign n5017 = pi75 & n4994;
  assign n5018 = ~pi92 & ~n5017;
  assign n5019 = ~n5016 & n5018;
  assign n5020 = n3230 & ~n5013;
  assign n5021 = ~n3230 & n4994;
  assign n5022 = pi92 & ~n5021;
  assign n5023 = ~n5020 & n5022;
  assign n5024 = n3265 & ~n5023;
  assign n5025 = ~n5019 & n5024;
  assign n5026 = ~n3265 & n4994;
  assign n5027 = ~pi55 & ~n5026;
  assign n5028 = ~n5025 & n5027;
  assign n5029 = n3268 & n4985;
  assign n5030 = ~n3268 & n4992;
  assign n5031 = pi55 & ~n5030;
  assign n5032 = ~n5029 & n5031;
  assign n5033 = ~pi56 & ~n5032;
  assign n5034 = ~n5028 & n5033;
  assign n5035 = n3280 & ~n4985;
  assign n5036 = ~n3280 & ~n4992;
  assign n5037 = pi56 & ~n5036;
  assign n5038 = ~n5035 & n5037;
  assign n5039 = ~pi62 & ~n5038;
  assign n5040 = ~n5034 & n5039;
  assign n5041 = n3431 & n4985;
  assign n5042 = ~n3431 & n4992;
  assign n5043 = pi62 & ~n5042;
  assign n5044 = ~n5041 & n5043;
  assign n5045 = pi246 & n3429;
  assign n5046 = ~n5044 & n5045;
  assign n5047 = ~n5040 & n5046;
  assign n5048 = pi246 & n4991;
  assign n5049 = ~n3429 & ~n5048;
  assign n5050 = n4904 & n5049;
  assign n5051 = ~n5047 & ~n5050;
  assign po161 = ~n4963 & n5051;
  assign n5053 = pi215 & pi1137;
  assign n5054 = pi299 & ~n5053;
  assign n5055 = ~pi933 & n2437;
  assign n5056 = ~pi1137 & ~n2437;
  assign n5057 = pi221 & ~n5056;
  assign n5058 = ~n5055 & n5057;
  assign n5059 = pi216 & pi280;
  assign n5060 = ~pi221 & ~n5059;
  assign n5061 = pi878 & n3460;
  assign n5062 = ~pi168 & ~n5061;
  assign n5063 = pi168 & n3453;
  assign n5064 = ~n5062 & ~n5063;
  assign n5065 = pi878 & ~n5064;
  assign n5066 = ~n3364 & n5062;
  assign n5067 = ~n5065 & ~n5066;
  assign n5068 = ~pi228 & ~n5067;
  assign n5069 = pi878 & ~n2449;
  assign n5070 = pi105 & ~n5069;
  assign n5071 = ~pi105 & pi168;
  assign n5072 = pi228 & ~n5071;
  assign n5073 = ~n5070 & n5072;
  assign n5074 = ~n3458 & n5073;
  assign n5075 = ~pi216 & ~n5074;
  assign n5076 = ~n5068 & n5075;
  assign n5077 = n5060 & ~n5076;
  assign n5078 = ~n5058 & ~n5077;
  assign n5079 = ~pi215 & ~n5078;
  assign n5080 = n5054 & ~n5079;
  assign n5081 = pi223 & pi1137;
  assign n5082 = ~pi299 & ~n5081;
  assign n5083 = ~pi933 & n3040;
  assign n5084 = ~pi1137 & ~n3040;
  assign n5085 = pi222 & ~n5084;
  assign n5086 = ~n5083 & n5085;
  assign n5087 = pi224 & pi280;
  assign n5088 = ~pi222 & ~n5087;
  assign n5089 = pi878 & n3441;
  assign n5090 = ~pi224 & ~n5089;
  assign n5091 = n5088 & ~n5090;
  assign n5092 = ~n5086 & ~n5091;
  assign n5093 = n5082 & n5092;
  assign n5094 = ~n3441 & n5088;
  assign n5095 = n5092 & ~n5094;
  assign n5096 = ~pi223 & ~n5095;
  assign n5097 = n5082 & ~n5096;
  assign n5098 = ~pi39 & ~n5097;
  assign n5099 = ~n5093 & n5098;
  assign n5100 = ~n5080 & n5099;
  assign n5101 = ~pi224 & ~n5069;
  assign n5102 = n5088 & ~n5101;
  assign n5103 = ~n5086 & ~n5102;
  assign n5104 = ~pi223 & ~n5103;
  assign n5105 = ~n5081 & ~n5104;
  assign n5106 = ~pi299 & ~n5105;
  assign n5107 = ~pi216 & ~n5073;
  assign n5108 = pi168 & ~n3095;
  assign n5109 = ~pi878 & n3095;
  assign n5110 = ~pi228 & ~n5109;
  assign n5111 = ~n5108 & n5110;
  assign n5112 = n5107 & ~n5111;
  assign n5113 = n5060 & ~n5112;
  assign n5114 = ~n5058 & ~n5113;
  assign n5115 = ~pi215 & ~n5114;
  assign n5116 = ~n5053 & ~n5115;
  assign n5117 = pi299 & ~n5116;
  assign n5118 = ~n5106 & ~n5117;
  assign n5119 = pi39 & ~n5118;
  assign n5120 = ~pi38 & ~n5119;
  assign n5121 = ~n5100 & n5120;
  assign n5122 = ~pi168 & ~pi228;
  assign n5123 = n5107 & ~n5122;
  assign n5124 = n5060 & ~n5123;
  assign n5125 = ~n5058 & ~n5124;
  assign n5126 = ~pi215 & ~n5125;
  assign n5127 = ~n5053 & ~n5126;
  assign n5128 = pi299 & ~n5127;
  assign n5129 = ~n5106 & ~n5128;
  assign n5130 = pi38 & n5129;
  assign n5131 = ~pi100 & ~n5130;
  assign n5132 = ~n5121 & n5131;
  assign n5133 = pi168 & ~n3388;
  assign n5134 = ~pi878 & n3388;
  assign n5135 = ~pi228 & ~n5134;
  assign n5136 = ~n5133 & n5135;
  assign n5137 = n5107 & ~n5136;
  assign n5138 = n5060 & ~n5137;
  assign n5139 = ~n5058 & ~n5138;
  assign n5140 = ~pi215 & ~n5139;
  assign n5141 = ~n5053 & ~n5140;
  assign n5142 = pi299 & ~n5141;
  assign n5143 = n3181 & ~n5106;
  assign n5144 = ~n5142 & n5143;
  assign n5145 = ~n3181 & n5129;
  assign n5146 = pi100 & ~n5145;
  assign n5147 = ~n5144 & n5146;
  assign n5148 = ~n5132 & ~n5147;
  assign n5149 = ~pi87 & ~n5148;
  assign n5150 = ~n3207 & n5129;
  assign n5151 = n3207 & n5118;
  assign n5152 = ~n5150 & ~n5151;
  assign n5153 = pi87 & n5152;
  assign n5154 = ~pi75 & ~n5153;
  assign n5155 = ~n5149 & n5154;
  assign n5156 = pi75 & n5129;
  assign n5157 = ~pi92 & ~n5156;
  assign n5158 = ~n5155 & n5157;
  assign n5159 = n3230 & ~n5152;
  assign n5160 = ~n3230 & n5129;
  assign n5161 = pi92 & ~n5160;
  assign n5162 = ~n5159 & n5161;
  assign n5163 = n3265 & ~n5162;
  assign n5164 = ~n5158 & n5163;
  assign n5165 = ~n3265 & n5129;
  assign n5166 = ~pi55 & ~n5165;
  assign n5167 = ~n5164 & n5166;
  assign n5168 = n3268 & n5116;
  assign n5169 = ~n3268 & n5127;
  assign n5170 = pi55 & ~n5169;
  assign n5171 = ~n5168 & n5170;
  assign n5172 = ~pi56 & ~n5171;
  assign n5173 = ~n5167 & n5172;
  assign n5174 = n3280 & ~n5116;
  assign n5175 = ~n3280 & ~n5127;
  assign n5176 = pi56 & ~n5175;
  assign n5177 = ~n5174 & n5176;
  assign n5178 = ~pi62 & ~n5177;
  assign n5179 = ~n5173 & n5178;
  assign n5180 = n3431 & n5116;
  assign n5181 = ~n3431 & n5127;
  assign n5182 = pi62 & ~n5181;
  assign n5183 = ~n5180 & n5182;
  assign n5184 = ~pi240 & n3429;
  assign n5185 = ~n5183 & n5184;
  assign n5186 = ~n5179 & n5185;
  assign n5187 = ~pi878 & n3453;
  assign n5188 = ~pi168 & ~n5187;
  assign n5189 = pi878 & ~n3364;
  assign n5190 = ~pi878 & ~n3460;
  assign n5191 = pi168 & ~n5190;
  assign n5192 = ~n5189 & n5191;
  assign n5193 = ~n5188 & ~n5192;
  assign n5194 = ~pi228 & ~n5193;
  assign n5195 = ~n3845 & n5107;
  assign n5196 = ~n5194 & n5195;
  assign n5197 = n5060 & ~n5196;
  assign n5198 = ~n5058 & ~n5197;
  assign n5199 = ~pi215 & ~n5198;
  assign n5200 = n5054 & ~n5199;
  assign n5201 = n5098 & ~n5200;
  assign n5202 = ~n3476 & ~n5106;
  assign n5203 = ~n3470 & n5107;
  assign n5204 = ~n5111 & n5203;
  assign n5205 = n5060 & ~n5204;
  assign n5206 = ~n5058 & ~n5205;
  assign n5207 = ~pi215 & ~n5206;
  assign n5208 = ~n5053 & ~n5207;
  assign n5209 = pi299 & ~n5208;
  assign n5210 = n5202 & ~n5209;
  assign n5211 = pi39 & ~n5210;
  assign n5212 = ~pi38 & ~n5211;
  assign n5213 = ~n5201 & n5212;
  assign n5214 = n3584 & ~n5059;
  assign n5215 = n5127 & ~n5214;
  assign n5216 = pi299 & ~n5215;
  assign n5217 = n5202 & ~n5216;
  assign n5218 = pi38 & n5217;
  assign n5219 = ~pi100 & ~n5218;
  assign n5220 = ~n5213 & n5219;
  assign n5221 = ~n5136 & n5203;
  assign n5222 = n5060 & ~n5221;
  assign n5223 = ~n5058 & ~n5222;
  assign n5224 = ~pi215 & ~n5223;
  assign n5225 = ~n5053 & ~n5224;
  assign n5226 = pi299 & ~n5225;
  assign n5227 = n3181 & n5202;
  assign n5228 = ~n5226 & n5227;
  assign n5229 = ~n3181 & n5217;
  assign n5230 = pi100 & ~n5229;
  assign n5231 = ~n5228 & n5230;
  assign n5232 = ~n5220 & ~n5231;
  assign n5233 = ~pi87 & ~n5232;
  assign n5234 = ~n3207 & n5217;
  assign n5235 = n3207 & n5210;
  assign n5236 = ~n5234 & ~n5235;
  assign n5237 = pi87 & n5236;
  assign n5238 = ~pi75 & ~n5237;
  assign n5239 = ~n5233 & n5238;
  assign n5240 = pi75 & n5217;
  assign n5241 = ~pi92 & ~n5240;
  assign n5242 = ~n5239 & n5241;
  assign n5243 = n3230 & ~n5236;
  assign n5244 = ~n3230 & n5217;
  assign n5245 = pi92 & ~n5244;
  assign n5246 = ~n5243 & n5245;
  assign n5247 = n3265 & ~n5246;
  assign n5248 = ~n5242 & n5247;
  assign n5249 = ~n3265 & n5217;
  assign n5250 = ~pi55 & ~n5249;
  assign n5251 = ~n5248 & n5250;
  assign n5252 = n3268 & n5208;
  assign n5253 = ~n3268 & n5215;
  assign n5254 = pi55 & ~n5253;
  assign n5255 = ~n5252 & n5254;
  assign n5256 = ~pi56 & ~n5255;
  assign n5257 = ~n5251 & n5256;
  assign n5258 = n3280 & ~n5208;
  assign n5259 = ~n3280 & ~n5215;
  assign n5260 = pi56 & ~n5259;
  assign n5261 = ~n5258 & n5260;
  assign n5262 = ~pi62 & ~n5261;
  assign n5263 = ~n5257 & n5262;
  assign n5264 = n3431 & n5208;
  assign n5265 = ~n3431 & n5215;
  assign n5266 = pi62 & ~n5265;
  assign n5267 = ~n5264 & n5266;
  assign n5268 = pi240 & n3429;
  assign n5269 = ~n5267 & n5268;
  assign n5270 = ~n5263 & n5269;
  assign n5271 = pi240 & n5214;
  assign n5272 = ~n3429 & ~n5271;
  assign n5273 = n5127 & n5272;
  assign n5274 = ~n5270 & ~n5273;
  assign po162 = ~n5186 & n5274;
  assign n5276 = ~pi928 & n2437;
  assign n5277 = ~pi1136 & ~n2437;
  assign n5278 = pi221 & ~n5277;
  assign n5279 = ~n5276 & n5278;
  assign n5280 = pi216 & pi266;
  assign n5281 = pi875 & ~n2449;
  assign n5282 = pi105 & ~n5281;
  assign n5283 = ~pi105 & ~pi166;
  assign n5284 = ~n5282 & ~n5283;
  assign n5285 = n3459 & ~n5284;
  assign n5286 = ~pi216 & ~n5285;
  assign n5287 = ~pi166 & ~n3453;
  assign n5288 = pi166 & n3460;
  assign n5289 = pi875 & ~n5288;
  assign n5290 = ~n5287 & n5289;
  assign n5291 = pi166 & ~pi875;
  assign n5292 = ~n3364 & n5291;
  assign n5293 = ~n5290 & ~n5292;
  assign n5294 = ~pi228 & ~n5293;
  assign n5295 = ~n3459 & ~n5294;
  assign n5296 = n5286 & ~n5295;
  assign n5297 = ~n5280 & ~n5296;
  assign n5298 = ~pi221 & ~n5297;
  assign n5299 = ~n5279 & ~n5298;
  assign n5300 = ~pi215 & ~n5299;
  assign n5301 = pi215 & pi1136;
  assign n5302 = pi299 & ~n5301;
  assign n5303 = ~n5300 & n5302;
  assign n5304 = ~pi224 & ~pi875;
  assign n5305 = ~n2449 & n5304;
  assign n5306 = pi224 & ~pi266;
  assign n5307 = ~pi222 & ~n5306;
  assign n5308 = ~n5305 & n5307;
  assign n5309 = n3052 & ~n3441;
  assign n5310 = n5308 & ~n5309;
  assign n5311 = ~pi928 & n3040;
  assign n5312 = ~pi1136 & ~n3040;
  assign n5313 = pi222 & ~n5312;
  assign n5314 = ~n5311 & n5313;
  assign n5315 = pi223 & pi1136;
  assign n5316 = ~pi299 & ~n5315;
  assign n5317 = ~n5314 & n5316;
  assign n5318 = ~n5310 & n5317;
  assign n5319 = ~n5308 & ~n5314;
  assign n5320 = ~n5309 & n5319;
  assign n5321 = ~pi223 & ~n5320;
  assign n5322 = n5316 & ~n5321;
  assign n5323 = ~pi39 & ~n5322;
  assign n5324 = ~n5318 & n5323;
  assign n5325 = ~n5303 & n5324;
  assign n5326 = pi228 & n5284;
  assign n5327 = ~pi875 & n3095;
  assign n5328 = pi166 & ~pi228;
  assign n5329 = ~n3321 & ~n5328;
  assign n5330 = ~n5327 & ~n5329;
  assign n5331 = ~n5326 & ~n5330;
  assign n5332 = ~pi216 & ~n5331;
  assign n5333 = ~n5280 & ~n5332;
  assign n5334 = ~pi221 & ~n5333;
  assign n5335 = ~n5279 & ~n5334;
  assign n5336 = ~pi215 & ~n5335;
  assign n5337 = ~n5301 & ~n5336;
  assign n5338 = pi299 & ~n5337;
  assign n5339 = ~pi223 & ~n5319;
  assign n5340 = ~n5315 & ~n5339;
  assign n5341 = ~pi299 & ~n5340;
  assign n5342 = ~n3856 & n5341;
  assign n5343 = ~n5338 & ~n5342;
  assign n5344 = pi39 & ~n5343;
  assign n5345 = ~pi38 & ~n5344;
  assign n5346 = ~n5325 & n5345;
  assign n5347 = ~n5326 & ~n5328;
  assign n5348 = ~pi216 & ~n5347;
  assign n5349 = ~n5280 & ~n5348;
  assign n5350 = ~pi221 & ~n5349;
  assign n5351 = ~n5279 & ~n5350;
  assign n5352 = ~pi215 & ~n5351;
  assign n5353 = ~n5301 & ~n5352;
  assign n5354 = pi299 & ~n5353;
  assign n5355 = ~n5342 & ~n5354;
  assign n5356 = pi38 & n5355;
  assign n5357 = ~pi100 & ~n5356;
  assign n5358 = ~n5346 & n5357;
  assign n5359 = ~pi875 & n3381;
  assign n5360 = pi166 & ~n5359;
  assign n5361 = ~n2447 & ~n3381;
  assign n5362 = n2447 & ~n3379;
  assign n5363 = pi875 & ~n5362;
  assign n5364 = ~n5361 & n5363;
  assign n5365 = ~n5360 & ~n5364;
  assign n5366 = ~pi228 & ~n5365;
  assign n5367 = ~n5326 & ~n5366;
  assign n5368 = ~pi216 & ~n5367;
  assign n5369 = ~n5280 & ~n5368;
  assign n5370 = ~pi221 & ~n5369;
  assign n5371 = ~n5279 & ~n5370;
  assign n5372 = ~pi215 & ~n5371;
  assign n5373 = ~n5301 & ~n5372;
  assign n5374 = pi299 & ~n5373;
  assign n5375 = n3181 & ~n5342;
  assign n5376 = ~n5374 & n5375;
  assign n5377 = ~n3181 & n5355;
  assign n5378 = pi100 & ~n5377;
  assign n5379 = ~n5376 & n5378;
  assign n5380 = ~n5358 & ~n5379;
  assign n5381 = ~pi87 & ~n5380;
  assign n5382 = ~n3207 & n5355;
  assign n5383 = n3207 & n5343;
  assign n5384 = ~n5382 & ~n5383;
  assign n5385 = pi87 & n5384;
  assign n5386 = ~pi75 & ~n5385;
  assign n5387 = ~n5381 & n5386;
  assign n5388 = pi75 & n5355;
  assign n5389 = ~pi92 & ~n5388;
  assign n5390 = ~n5387 & n5389;
  assign n5391 = n3230 & ~n5384;
  assign n5392 = ~n3230 & n5355;
  assign n5393 = pi92 & ~n5392;
  assign n5394 = ~n5391 & n5393;
  assign n5395 = n3265 & ~n5394;
  assign n5396 = ~n5390 & n5395;
  assign n5397 = ~n3265 & n5355;
  assign n5398 = ~pi55 & ~n5397;
  assign n5399 = ~n5396 & n5398;
  assign n5400 = n3268 & n5337;
  assign n5401 = ~n3268 & n5353;
  assign n5402 = pi55 & ~n5401;
  assign n5403 = ~n5400 & n5402;
  assign n5404 = ~pi56 & ~n5403;
  assign n5405 = ~n5399 & n5404;
  assign n5406 = n3280 & ~n5337;
  assign n5407 = ~n3280 & ~n5353;
  assign n5408 = pi56 & ~n5407;
  assign n5409 = ~n5406 & n5408;
  assign n5410 = ~pi62 & ~n5409;
  assign n5411 = ~n5405 & n5410;
  assign n5412 = n3431 & n5337;
  assign n5413 = ~n3431 & n5353;
  assign n5414 = pi62 & ~n5413;
  assign n5415 = ~n5412 & n5414;
  assign n5416 = n3429 & ~n5415;
  assign n5417 = ~n5411 & n5416;
  assign n5418 = ~n3429 & n5353;
  assign n5419 = ~pi245 & ~n5418;
  assign n5420 = ~n5417 & n5419;
  assign n5421 = ~pi166 & ~n3364;
  assign n5422 = pi875 & ~n5421;
  assign n5423 = pi166 & n3453;
  assign n5424 = ~pi166 & ~n3460;
  assign n5425 = ~pi875 & ~n5424;
  assign n5426 = ~n5423 & n5425;
  assign n5427 = ~pi228 & ~n5426;
  assign n5428 = ~n5422 & n5427;
  assign n5429 = n5286 & ~n5428;
  assign n5430 = ~n5280 & ~n5429;
  assign n5431 = ~pi221 & ~n5430;
  assign n5432 = ~n5279 & ~n5431;
  assign n5433 = ~pi215 & ~n5432;
  assign n5434 = n5302 & ~n5433;
  assign n5435 = n5323 & ~n5434;
  assign n5436 = ~n3470 & ~n5326;
  assign n5437 = ~n5330 & n5436;
  assign n5438 = ~pi216 & ~n5437;
  assign n5439 = ~n5280 & ~n5438;
  assign n5440 = ~pi221 & ~n5439;
  assign n5441 = ~n5279 & ~n5440;
  assign n5442 = ~pi215 & ~n5441;
  assign n5443 = ~n5301 & ~n5442;
  assign n5444 = pi299 & ~n5443;
  assign n5445 = ~n5341 & ~n5444;
  assign n5446 = pi39 & ~n5445;
  assign n5447 = ~pi38 & ~n5446;
  assign n5448 = ~n5435 & n5447;
  assign n5449 = ~n3471 & n5353;
  assign n5450 = pi299 & ~n5449;
  assign n5451 = ~n5341 & ~n5450;
  assign n5452 = pi38 & n5451;
  assign n5453 = ~pi100 & ~n5452;
  assign n5454 = ~n5448 & n5453;
  assign n5455 = ~n5366 & n5436;
  assign n5456 = ~pi216 & ~n5455;
  assign n5457 = ~n5280 & ~n5456;
  assign n5458 = ~pi221 & ~n5457;
  assign n5459 = ~n5279 & ~n5458;
  assign n5460 = ~pi215 & ~n5459;
  assign n5461 = ~n5301 & ~n5460;
  assign n5462 = pi299 & ~n5461;
  assign n5463 = n3181 & ~n5341;
  assign n5464 = ~n5462 & n5463;
  assign n5465 = ~n3181 & n5451;
  assign n5466 = pi100 & ~n5465;
  assign n5467 = ~n5464 & n5466;
  assign n5468 = ~n5454 & ~n5467;
  assign n5469 = ~pi87 & ~n5468;
  assign n5470 = ~n3207 & n5451;
  assign n5471 = n3207 & n5445;
  assign n5472 = ~n5470 & ~n5471;
  assign n5473 = pi87 & n5472;
  assign n5474 = ~pi75 & ~n5473;
  assign n5475 = ~n5469 & n5474;
  assign n5476 = pi75 & n5451;
  assign n5477 = ~pi92 & ~n5476;
  assign n5478 = ~n5475 & n5477;
  assign n5479 = n3230 & ~n5472;
  assign n5480 = ~n3230 & n5451;
  assign n5481 = pi92 & ~n5480;
  assign n5482 = ~n5479 & n5481;
  assign n5483 = n3265 & ~n5482;
  assign n5484 = ~n5478 & n5483;
  assign n5485 = ~n3265 & n5451;
  assign n5486 = ~pi55 & ~n5485;
  assign n5487 = ~n5484 & n5486;
  assign n5488 = n3268 & n5443;
  assign n5489 = ~n3268 & n5449;
  assign n5490 = pi55 & ~n5489;
  assign n5491 = ~n5488 & n5490;
  assign n5492 = ~pi56 & ~n5491;
  assign n5493 = ~n5487 & n5492;
  assign n5494 = n3280 & ~n5443;
  assign n5495 = ~n3280 & ~n5449;
  assign n5496 = pi56 & ~n5495;
  assign n5497 = ~n5494 & n5496;
  assign n5498 = ~pi62 & ~n5497;
  assign n5499 = ~n5493 & n5498;
  assign n5500 = n3431 & n5443;
  assign n5501 = ~n3431 & n5449;
  assign n5502 = pi62 & ~n5501;
  assign n5503 = ~n5500 & n5502;
  assign n5504 = n3429 & ~n5503;
  assign n5505 = ~n5499 & n5504;
  assign n5506 = ~n3429 & n5449;
  assign n5507 = pi245 & ~n5506;
  assign n5508 = ~n5505 & n5507;
  assign po163 = n5420 | n5508;
  assign n5510 = ~pi938 & n2437;
  assign n5511 = ~pi1135 & ~n2437;
  assign n5512 = pi221 & ~n5511;
  assign n5513 = ~n5510 & n5512;
  assign n5514 = pi216 & pi279;
  assign n5515 = pi879 & ~n2449;
  assign n5516 = pi105 & ~n5515;
  assign n5517 = ~pi105 & ~pi161;
  assign n5518 = ~n5516 & ~n5517;
  assign n5519 = n3459 & ~n5518;
  assign n5520 = ~pi216 & ~n5519;
  assign n5521 = ~pi161 & ~n3453;
  assign n5522 = pi161 & n3460;
  assign n5523 = pi879 & ~n5522;
  assign n5524 = ~n5521 & n5523;
  assign n5525 = pi161 & ~pi879;
  assign n5526 = ~n3364 & n5525;
  assign n5527 = ~n5524 & ~n5526;
  assign n5528 = ~pi228 & ~n5527;
  assign n5529 = ~n3459 & ~n5528;
  assign n5530 = n5520 & ~n5529;
  assign n5531 = ~n5514 & ~n5530;
  assign n5532 = ~pi221 & ~n5531;
  assign n5533 = ~n5513 & ~n5532;
  assign n5534 = ~pi215 & ~n5533;
  assign n5535 = pi215 & pi1135;
  assign n5536 = pi299 & ~n5535;
  assign n5537 = ~n5534 & n5536;
  assign n5538 = pi223 & pi1135;
  assign n5539 = ~pi299 & ~n5538;
  assign n5540 = ~pi938 & n3040;
  assign n5541 = ~pi1135 & ~n3040;
  assign n5542 = pi222 & ~n5541;
  assign n5543 = ~n5540 & n5542;
  assign n5544 = ~pi224 & ~pi879;
  assign n5545 = ~n2449 & n5544;
  assign n5546 = pi224 & ~pi279;
  assign n5547 = ~pi222 & ~n5546;
  assign n5548 = ~n5545 & n5547;
  assign n5549 = ~n5543 & ~n5548;
  assign n5550 = ~pi223 & ~n5549;
  assign n5551 = n5309 & ~n5543;
  assign n5552 = n5550 & ~n5551;
  assign n5553 = n5539 & ~n5552;
  assign n5554 = ~pi39 & ~n5553;
  assign n5555 = ~n5537 & n5554;
  assign n5556 = pi228 & n5518;
  assign n5557 = ~pi879 & n3095;
  assign n5558 = pi161 & ~pi228;
  assign n5559 = ~n3321 & ~n5558;
  assign n5560 = ~n5557 & ~n5559;
  assign n5561 = ~n5556 & ~n5560;
  assign n5562 = ~pi216 & ~n5561;
  assign n5563 = ~n5514 & ~n5562;
  assign n5564 = ~pi221 & ~n5563;
  assign n5565 = ~n5513 & ~n5564;
  assign n5566 = ~pi215 & ~n5565;
  assign n5567 = ~n5535 & ~n5566;
  assign n5568 = pi299 & ~n5567;
  assign n5569 = ~n5538 & ~n5550;
  assign n5570 = ~pi299 & ~n5569;
  assign n5571 = ~n3856 & n5570;
  assign n5572 = ~n5568 & ~n5571;
  assign n5573 = pi39 & ~n5572;
  assign n5574 = ~pi38 & ~n5573;
  assign n5575 = ~n5555 & n5574;
  assign n5576 = ~n5556 & ~n5558;
  assign n5577 = ~pi216 & ~n5576;
  assign n5578 = ~n5514 & ~n5577;
  assign n5579 = ~pi221 & ~n5578;
  assign n5580 = ~n5513 & ~n5579;
  assign n5581 = ~pi215 & ~n5580;
  assign n5582 = ~n5535 & ~n5581;
  assign n5583 = pi299 & ~n5582;
  assign n5584 = ~n5571 & ~n5583;
  assign n5585 = pi38 & n5584;
  assign n5586 = ~pi100 & ~n5585;
  assign n5587 = ~n5575 & n5586;
  assign n5588 = ~pi879 & n3381;
  assign n5589 = pi161 & ~n5588;
  assign n5590 = ~pi152 & ~pi166;
  assign n5591 = ~n3381 & ~n5590;
  assign n5592 = ~n3379 & n5590;
  assign n5593 = pi879 & ~n5592;
  assign n5594 = ~n5591 & n5593;
  assign n5595 = ~n5589 & ~n5594;
  assign n5596 = ~pi228 & ~n5595;
  assign n5597 = ~n5556 & ~n5596;
  assign n5598 = ~pi216 & ~n5597;
  assign n5599 = ~n5514 & ~n5598;
  assign n5600 = ~pi221 & ~n5599;
  assign n5601 = ~n5513 & ~n5600;
  assign n5602 = ~pi215 & ~n5601;
  assign n5603 = ~n5535 & ~n5602;
  assign n5604 = pi299 & ~n5603;
  assign n5605 = n3181 & ~n5571;
  assign n5606 = ~n5604 & n5605;
  assign n5607 = ~n3181 & n5584;
  assign n5608 = pi100 & ~n5607;
  assign n5609 = ~n5606 & n5608;
  assign n5610 = ~n5587 & ~n5609;
  assign n5611 = ~pi87 & ~n5610;
  assign n5612 = ~n3207 & n5584;
  assign n5613 = n3207 & n5572;
  assign n5614 = ~n5612 & ~n5613;
  assign n5615 = pi87 & n5614;
  assign n5616 = ~pi75 & ~n5615;
  assign n5617 = ~n5611 & n5616;
  assign n5618 = pi75 & n5584;
  assign n5619 = ~pi92 & ~n5618;
  assign n5620 = ~n5617 & n5619;
  assign n5621 = n3230 & ~n5614;
  assign n5622 = ~n3230 & n5584;
  assign n5623 = pi92 & ~n5622;
  assign n5624 = ~n5621 & n5623;
  assign n5625 = n3265 & ~n5624;
  assign n5626 = ~n5620 & n5625;
  assign n5627 = ~n3265 & n5584;
  assign n5628 = ~pi55 & ~n5627;
  assign n5629 = ~n5626 & n5628;
  assign n5630 = n3268 & n5567;
  assign n5631 = ~n3268 & n5582;
  assign n5632 = pi55 & ~n5631;
  assign n5633 = ~n5630 & n5632;
  assign n5634 = ~pi56 & ~n5633;
  assign n5635 = ~n5629 & n5634;
  assign n5636 = n3280 & ~n5567;
  assign n5637 = ~n3280 & ~n5582;
  assign n5638 = pi56 & ~n5637;
  assign n5639 = ~n5636 & n5638;
  assign n5640 = ~pi62 & ~n5639;
  assign n5641 = ~n5635 & n5640;
  assign n5642 = n3431 & n5567;
  assign n5643 = ~n3431 & n5582;
  assign n5644 = pi62 & ~n5643;
  assign n5645 = ~n5642 & n5644;
  assign n5646 = n3429 & ~n5645;
  assign n5647 = ~n5641 & n5646;
  assign n5648 = ~n3429 & n5582;
  assign n5649 = ~pi244 & ~n5648;
  assign n5650 = ~n5647 & n5649;
  assign n5651 = ~pi161 & ~n3364;
  assign n5652 = pi879 & ~n5651;
  assign n5653 = pi161 & n3453;
  assign n5654 = ~pi161 & ~n3460;
  assign n5655 = ~pi879 & ~n5654;
  assign n5656 = ~n5653 & n5655;
  assign n5657 = ~pi228 & ~n5656;
  assign n5658 = ~n5652 & n5657;
  assign n5659 = n5520 & ~n5658;
  assign n5660 = ~n5514 & ~n5659;
  assign n5661 = ~pi221 & ~n5660;
  assign n5662 = ~n5513 & ~n5661;
  assign n5663 = ~pi215 & ~n5662;
  assign n5664 = n5536 & ~n5663;
  assign n5665 = ~n5309 & n5549;
  assign n5666 = ~pi223 & ~n5665;
  assign n5667 = n5539 & ~n5666;
  assign n5668 = ~pi39 & ~n5667;
  assign n5669 = ~n5664 & n5668;
  assign n5670 = ~n3470 & ~n5556;
  assign n5671 = ~n5560 & n5670;
  assign n5672 = ~pi216 & ~n5671;
  assign n5673 = ~n5514 & ~n5672;
  assign n5674 = ~pi221 & ~n5673;
  assign n5675 = ~n5513 & ~n5674;
  assign n5676 = ~pi215 & ~n5675;
  assign n5677 = ~n5535 & ~n5676;
  assign n5678 = pi299 & ~n5677;
  assign n5679 = ~n5570 & ~n5678;
  assign n5680 = pi39 & ~n5679;
  assign n5681 = ~pi38 & ~n5680;
  assign n5682 = ~n5669 & n5681;
  assign n5683 = ~n3471 & n5582;
  assign n5684 = pi299 & ~n5683;
  assign n5685 = ~n5570 & ~n5684;
  assign n5686 = pi38 & n5685;
  assign n5687 = ~pi100 & ~n5686;
  assign n5688 = ~n5682 & n5687;
  assign n5689 = ~n5596 & n5670;
  assign n5690 = ~pi216 & ~n5689;
  assign n5691 = ~n5514 & ~n5690;
  assign n5692 = ~pi221 & ~n5691;
  assign n5693 = ~n5513 & ~n5692;
  assign n5694 = ~pi215 & ~n5693;
  assign n5695 = ~n5535 & ~n5694;
  assign n5696 = pi299 & ~n5695;
  assign n5697 = n3181 & ~n5570;
  assign n5698 = ~n5696 & n5697;
  assign n5699 = ~n3181 & n5685;
  assign n5700 = pi100 & ~n5699;
  assign n5701 = ~n5698 & n5700;
  assign n5702 = ~n5688 & ~n5701;
  assign n5703 = ~pi87 & ~n5702;
  assign n5704 = ~n3207 & n5685;
  assign n5705 = n3207 & n5679;
  assign n5706 = ~n5704 & ~n5705;
  assign n5707 = pi87 & n5706;
  assign n5708 = ~pi75 & ~n5707;
  assign n5709 = ~n5703 & n5708;
  assign n5710 = pi75 & n5685;
  assign n5711 = ~pi92 & ~n5710;
  assign n5712 = ~n5709 & n5711;
  assign n5713 = n3230 & ~n5706;
  assign n5714 = ~n3230 & n5685;
  assign n5715 = pi92 & ~n5714;
  assign n5716 = ~n5713 & n5715;
  assign n5717 = n3265 & ~n5716;
  assign n5718 = ~n5712 & n5717;
  assign n5719 = ~n3265 & n5685;
  assign n5720 = ~pi55 & ~n5719;
  assign n5721 = ~n5718 & n5720;
  assign n5722 = n3268 & n5677;
  assign n5723 = ~n3268 & n5683;
  assign n5724 = pi55 & ~n5723;
  assign n5725 = ~n5722 & n5724;
  assign n5726 = ~pi56 & ~n5725;
  assign n5727 = ~n5721 & n5726;
  assign n5728 = n3280 & ~n5677;
  assign n5729 = ~n3280 & ~n5683;
  assign n5730 = pi56 & ~n5729;
  assign n5731 = ~n5728 & n5730;
  assign n5732 = ~pi62 & ~n5731;
  assign n5733 = ~n5727 & n5732;
  assign n5734 = n3431 & n5677;
  assign n5735 = ~n3431 & n5683;
  assign n5736 = pi62 & ~n5735;
  assign n5737 = ~n5734 & n5736;
  assign n5738 = n3429 & ~n5737;
  assign n5739 = ~n5733 & n5738;
  assign n5740 = ~n3429 & n5683;
  assign n5741 = pi244 & ~n5740;
  assign n5742 = ~n5739 & n5741;
  assign po164 = n5650 | n5742;
  assign n5744 = pi833 & ~pi930;
  assign n5745 = ~pi216 & pi221;
  assign n5746 = n5744 & n5745;
  assign n5747 = pi216 & pi278;
  assign n5748 = ~pi221 & ~n5747;
  assign n5749 = ~pi105 & pi152;
  assign n5750 = pi228 & ~n5749;
  assign n5751 = ~pi846 & n3441;
  assign n5752 = pi105 & ~n5751;
  assign n5753 = n5750 & ~n5752;
  assign n5754 = ~pi216 & ~n5753;
  assign n5755 = pi152 & ~n3453;
  assign n5756 = ~pi152 & n3460;
  assign n5757 = ~pi846 & ~n5756;
  assign n5758 = ~n5755 & n5757;
  assign n5759 = ~pi152 & pi846;
  assign n5760 = ~n3364 & n5759;
  assign n5761 = ~n5758 & ~n5760;
  assign n5762 = ~pi228 & ~n5761;
  assign n5763 = n5754 & ~n5762;
  assign n5764 = n5748 & ~n5763;
  assign n5765 = ~n5746 & ~n5764;
  assign n5766 = pi221 & ~n2437;
  assign n5767 = ~pi215 & pi299;
  assign n5768 = ~n5766 & n5767;
  assign n5769 = n5765 & n5768;
  assign n5770 = pi222 & ~pi224;
  assign n5771 = n5744 & n5770;
  assign n5772 = pi224 & pi278;
  assign n5773 = ~pi222 & ~n5772;
  assign n5774 = ~pi224 & ~n5751;
  assign n5775 = n5773 & ~n5774;
  assign n5776 = ~n5771 & ~n5775;
  assign n5777 = ~n3041 & n3474;
  assign n5778 = n5776 & n5777;
  assign n5779 = ~pi39 & ~n5778;
  assign n5780 = ~n5769 & n5779;
  assign n5781 = pi846 & ~n2449;
  assign n5782 = ~pi224 & n5781;
  assign n5783 = n5773 & ~n5782;
  assign n5784 = n3042 & ~n5771;
  assign n5785 = ~n5783 & n5784;
  assign n5786 = ~pi299 & ~n5785;
  assign n5787 = ~n3856 & n5786;
  assign n5788 = ~pi215 & ~n5766;
  assign n5789 = ~n5746 & n5788;
  assign n5790 = pi105 & n5781;
  assign n5791 = ~n5749 & ~n5790;
  assign n5792 = pi228 & ~n5791;
  assign n5793 = ~n3470 & ~n5792;
  assign n5794 = ~pi846 & n3095;
  assign n5795 = pi152 & ~pi228;
  assign n5796 = ~n3321 & ~n5795;
  assign n5797 = ~n5794 & ~n5796;
  assign n5798 = n5793 & ~n5797;
  assign n5799 = ~pi216 & ~n5798;
  assign n5800 = n5748 & ~n5799;
  assign n5801 = n5789 & ~n5800;
  assign n5802 = pi299 & ~n5801;
  assign n5803 = ~n5787 & ~n5802;
  assign n5804 = pi39 & ~n5803;
  assign n5805 = ~pi38 & ~n5804;
  assign n5806 = ~n5780 & n5805;
  assign n5807 = ~n5792 & ~n5795;
  assign n5808 = ~pi216 & ~n5807;
  assign n5809 = n5748 & ~n5808;
  assign n5810 = n5789 & ~n5809;
  assign n5811 = ~n3471 & ~n5810;
  assign n5812 = pi299 & n5811;
  assign n5813 = ~n5787 & ~n5812;
  assign n5814 = pi38 & n5813;
  assign n5815 = ~pi100 & ~n5814;
  assign n5816 = ~n5806 & n5815;
  assign n5817 = pi846 & ~n3387;
  assign n5818 = ~n3382 & ~n5817;
  assign n5819 = ~pi228 & ~n5818;
  assign n5820 = n5793 & ~n5819;
  assign n5821 = ~pi216 & ~n5820;
  assign n5822 = n5748 & ~n5821;
  assign n5823 = n5789 & ~n5822;
  assign n5824 = pi299 & ~n5823;
  assign n5825 = n3181 & ~n5787;
  assign n5826 = ~n5824 & n5825;
  assign n5827 = ~n3181 & n5813;
  assign n5828 = pi100 & ~n5827;
  assign n5829 = ~n5826 & n5828;
  assign n5830 = ~n5816 & ~n5829;
  assign n5831 = ~pi87 & ~n5830;
  assign n5832 = ~n3207 & n5813;
  assign n5833 = n3207 & n5803;
  assign n5834 = ~n5832 & ~n5833;
  assign n5835 = pi87 & n5834;
  assign n5836 = ~pi75 & ~n5835;
  assign n5837 = ~n5831 & n5836;
  assign n5838 = pi75 & n5813;
  assign n5839 = ~pi92 & ~n5838;
  assign n5840 = ~n5837 & n5839;
  assign n5841 = n3230 & ~n5834;
  assign n5842 = ~n3230 & n5813;
  assign n5843 = pi92 & ~n5842;
  assign n5844 = ~n5841 & n5843;
  assign n5845 = n3265 & ~n5844;
  assign n5846 = ~n5840 & n5845;
  assign n5847 = ~n3265 & n5813;
  assign n5848 = ~pi55 & ~n5847;
  assign n5849 = ~n5846 & n5848;
  assign n5850 = n3268 & n5801;
  assign n5851 = ~n3268 & ~n5811;
  assign n5852 = pi55 & ~n5851;
  assign n5853 = ~n5850 & n5852;
  assign n5854 = ~pi56 & ~n5853;
  assign n5855 = ~n5849 & n5854;
  assign n5856 = n3280 & ~n5801;
  assign n5857 = ~n3280 & n5811;
  assign n5858 = pi56 & ~n5857;
  assign n5859 = ~n5856 & n5858;
  assign n5860 = ~pi62 & ~n5859;
  assign n5861 = ~n5855 & n5860;
  assign n5862 = n3431 & n5801;
  assign n5863 = ~n3431 & ~n5811;
  assign n5864 = pi62 & ~n5863;
  assign n5865 = ~n5862 & n5864;
  assign n5866 = n3429 & ~n5865;
  assign n5867 = ~n5861 & n5866;
  assign n5868 = ~n3429 & ~n5811;
  assign n5869 = pi242 & ~n5868;
  assign n5870 = ~n5867 & n5869;
  assign n5871 = ~pi152 & ~n3453;
  assign n5872 = pi152 & n3460;
  assign n5873 = pi846 & ~n5872;
  assign n5874 = ~n5871 & n5873;
  assign n5875 = pi152 & ~pi846;
  assign n5876 = ~n3364 & n5875;
  assign n5877 = ~pi228 & ~n5876;
  assign n5878 = ~n5874 & n5877;
  assign n5879 = ~n3441 & n5750;
  assign n5880 = n5754 & ~n5879;
  assign n5881 = ~n5878 & n5880;
  assign n5882 = n5748 & ~n5881;
  assign n5883 = ~n5746 & ~n5882;
  assign n5884 = n5768 & n5883;
  assign n5885 = ~n3440 & n5782;
  assign n5886 = n5773 & ~n5885;
  assign n5887 = ~n5771 & n5777;
  assign n5888 = ~n5886 & n5887;
  assign n5889 = ~pi39 & ~n5888;
  assign n5890 = ~n5884 & n5889;
  assign n5891 = ~n5792 & ~n5797;
  assign n5892 = ~pi216 & ~n5891;
  assign n5893 = n5748 & ~n5892;
  assign n5894 = n5789 & ~n5893;
  assign n5895 = pi299 & ~n5894;
  assign n5896 = ~n5786 & ~n5895;
  assign n5897 = pi39 & ~n5896;
  assign n5898 = ~pi38 & ~n5897;
  assign n5899 = ~n5890 & n5898;
  assign n5900 = pi299 & ~n5810;
  assign n5901 = ~n5786 & ~n5900;
  assign n5902 = pi38 & n5901;
  assign n5903 = ~pi100 & ~n5902;
  assign n5904 = ~n5899 & n5903;
  assign n5905 = ~n5792 & ~n5819;
  assign n5906 = ~pi216 & ~n5905;
  assign n5907 = n5748 & ~n5906;
  assign n5908 = n5789 & ~n5907;
  assign n5909 = pi299 & ~n5908;
  assign n5910 = n3181 & ~n5786;
  assign n5911 = ~n5909 & n5910;
  assign n5912 = ~n3181 & n5901;
  assign n5913 = pi100 & ~n5912;
  assign n5914 = ~n5911 & n5913;
  assign n5915 = ~n5904 & ~n5914;
  assign n5916 = ~pi87 & ~n5915;
  assign n5917 = ~n3207 & n5901;
  assign n5918 = n3207 & n5896;
  assign n5919 = ~n5917 & ~n5918;
  assign n5920 = pi87 & n5919;
  assign n5921 = ~pi75 & ~n5920;
  assign n5922 = ~n5916 & n5921;
  assign n5923 = pi75 & n5901;
  assign n5924 = ~pi92 & ~n5923;
  assign n5925 = ~n5922 & n5924;
  assign n5926 = n3230 & ~n5919;
  assign n5927 = ~n3230 & n5901;
  assign n5928 = pi92 & ~n5927;
  assign n5929 = ~n5926 & n5928;
  assign n5930 = n3265 & ~n5929;
  assign n5931 = ~n5925 & n5930;
  assign n5932 = ~n3265 & n5901;
  assign n5933 = ~pi55 & ~n5932;
  assign n5934 = ~n5931 & n5933;
  assign n5935 = n3268 & n5894;
  assign n5936 = ~n3268 & n5810;
  assign n5937 = pi55 & ~n5936;
  assign n5938 = ~n5935 & n5937;
  assign n5939 = ~pi56 & ~n5938;
  assign n5940 = ~n5934 & n5939;
  assign n5941 = n3280 & ~n5894;
  assign n5942 = ~n3280 & ~n5810;
  assign n5943 = pi56 & ~n5942;
  assign n5944 = ~n5941 & n5943;
  assign n5945 = ~pi62 & ~n5944;
  assign n5946 = ~n5940 & n5945;
  assign n5947 = n3431 & n5894;
  assign n5948 = ~n3431 & n5810;
  assign n5949 = pi62 & ~n5948;
  assign n5950 = ~n5947 & n5949;
  assign n5951 = n3429 & ~n5950;
  assign n5952 = ~n5946 & n5951;
  assign n5953 = ~n3429 & n5810;
  assign n5954 = ~pi242 & ~n5953;
  assign n5955 = ~n5952 & n5954;
  assign n5956 = ~n5870 & ~n5955;
  assign n5957 = ~pi1134 & ~n5956;
  assign n5958 = n3474 & ~n5776;
  assign n5959 = ~pi39 & ~n5958;
  assign n5960 = ~n5765 & n5767;
  assign n5961 = n5959 & ~n5960;
  assign n5962 = n3042 & n5787;
  assign n5963 = ~pi299 & ~n5962;
  assign n5964 = ~n5746 & ~n5800;
  assign n5965 = ~pi215 & ~n5964;
  assign n5966 = pi299 & ~n5965;
  assign n5967 = ~n5963 & ~n5966;
  assign n5968 = pi39 & ~n5967;
  assign n5969 = ~pi38 & ~n5968;
  assign n5970 = ~n5961 & n5969;
  assign n5971 = n5788 & ~n5810;
  assign n5972 = ~n3471 & n5971;
  assign n5973 = pi299 & ~n5972;
  assign n5974 = ~n5963 & ~n5973;
  assign n5975 = pi38 & n5974;
  assign n5976 = ~pi100 & ~n5975;
  assign n5977 = ~n5970 & n5976;
  assign n5978 = ~n5746 & ~n5822;
  assign n5979 = ~pi215 & ~n5978;
  assign n5980 = pi299 & ~n5979;
  assign n5981 = n3181 & ~n5963;
  assign n5982 = ~n5980 & n5981;
  assign n5983 = ~n3181 & n5974;
  assign n5984 = pi100 & ~n5983;
  assign n5985 = ~n5982 & n5984;
  assign n5986 = ~n5977 & ~n5985;
  assign n5987 = ~pi87 & ~n5986;
  assign n5988 = ~n3207 & n5974;
  assign n5989 = n3207 & n5967;
  assign n5990 = ~n5988 & ~n5989;
  assign n5991 = pi87 & n5990;
  assign n5992 = ~pi75 & ~n5991;
  assign n5993 = ~n5987 & n5992;
  assign n5994 = pi75 & n5974;
  assign n5995 = ~pi92 & ~n5994;
  assign n5996 = ~n5993 & n5995;
  assign n5997 = n3230 & ~n5990;
  assign n5998 = ~n3230 & n5974;
  assign n5999 = pi92 & ~n5998;
  assign n6000 = ~n5997 & n5999;
  assign n6001 = n3265 & ~n6000;
  assign n6002 = ~n5996 & n6001;
  assign n6003 = ~n3265 & n5974;
  assign n6004 = ~pi55 & ~n6003;
  assign n6005 = ~n6002 & n6004;
  assign n6006 = n3268 & n5965;
  assign n6007 = ~n3268 & n5972;
  assign n6008 = pi55 & ~n6007;
  assign n6009 = ~n6006 & n6008;
  assign n6010 = ~pi56 & ~n6009;
  assign n6011 = ~n6005 & n6010;
  assign n6012 = n3280 & ~n5965;
  assign n6013 = ~n3280 & ~n5972;
  assign n6014 = pi56 & ~n6013;
  assign n6015 = ~n6012 & n6014;
  assign n6016 = ~pi62 & ~n6015;
  assign n6017 = ~n6011 & n6016;
  assign n6018 = n3431 & n5965;
  assign n6019 = ~n3431 & n5972;
  assign n6020 = pi62 & ~n6019;
  assign n6021 = ~n6018 & n6020;
  assign n6022 = n3429 & ~n6021;
  assign n6023 = ~n6017 & n6022;
  assign n6024 = ~n3429 & n5972;
  assign n6025 = pi242 & ~n6024;
  assign n6026 = ~n6023 & n6025;
  assign n6027 = n5767 & ~n5883;
  assign n6028 = n3474 & n5886;
  assign n6029 = n5959 & ~n6028;
  assign n6030 = ~n6027 & n6029;
  assign n6031 = ~pi223 & n5783;
  assign n6032 = n5963 & ~n6031;
  assign n6033 = ~n5746 & ~n5893;
  assign n6034 = ~pi215 & ~n6033;
  assign n6035 = pi299 & ~n6034;
  assign n6036 = ~n6032 & ~n6035;
  assign n6037 = pi39 & ~n6036;
  assign n6038 = ~pi38 & ~n6037;
  assign n6039 = ~n6030 & n6038;
  assign n6040 = pi299 & ~n5971;
  assign n6041 = ~n6032 & ~n6040;
  assign n6042 = pi38 & n6041;
  assign n6043 = ~pi100 & ~n6042;
  assign n6044 = ~n6039 & n6043;
  assign n6045 = ~n5746 & ~n5907;
  assign n6046 = ~pi215 & ~n6045;
  assign n6047 = pi299 & ~n6046;
  assign n6048 = n3181 & ~n6032;
  assign n6049 = ~n6047 & n6048;
  assign n6050 = ~n3181 & n6041;
  assign n6051 = pi100 & ~n6050;
  assign n6052 = ~n6049 & n6051;
  assign n6053 = ~n6044 & ~n6052;
  assign n6054 = ~pi87 & ~n6053;
  assign n6055 = ~n3207 & n6041;
  assign n6056 = n3207 & n6036;
  assign n6057 = ~n6055 & ~n6056;
  assign n6058 = pi87 & n6057;
  assign n6059 = ~pi75 & ~n6058;
  assign n6060 = ~n6054 & n6059;
  assign n6061 = pi75 & n6041;
  assign n6062 = ~pi92 & ~n6061;
  assign n6063 = ~n6060 & n6062;
  assign n6064 = n3230 & ~n6057;
  assign n6065 = ~n3230 & n6041;
  assign n6066 = pi92 & ~n6065;
  assign n6067 = ~n6064 & n6066;
  assign n6068 = n3265 & ~n6067;
  assign n6069 = ~n6063 & n6068;
  assign n6070 = ~n3265 & n6041;
  assign n6071 = ~pi55 & ~n6070;
  assign n6072 = ~n6069 & n6071;
  assign n6073 = n3268 & n6034;
  assign n6074 = ~n3268 & n5971;
  assign n6075 = pi55 & ~n6074;
  assign n6076 = ~n6073 & n6075;
  assign n6077 = ~pi56 & ~n6076;
  assign n6078 = ~n6072 & n6077;
  assign n6079 = n3280 & ~n6034;
  assign n6080 = ~n3280 & ~n5971;
  assign n6081 = pi56 & ~n6080;
  assign n6082 = ~n6079 & n6081;
  assign n6083 = ~pi62 & ~n6082;
  assign n6084 = ~n6078 & n6083;
  assign n6085 = n3431 & n6034;
  assign n6086 = ~n3431 & n5971;
  assign n6087 = pi62 & ~n6086;
  assign n6088 = ~n6085 & n6087;
  assign n6089 = n3429 & ~n6088;
  assign n6090 = ~n6084 & n6089;
  assign n6091 = ~n3429 & n5971;
  assign n6092 = ~pi242 & ~n6091;
  assign n6093 = ~n6090 & n6092;
  assign n6094 = pi1134 & ~n6093;
  assign n6095 = ~n6026 & n6094;
  assign po165 = ~n5957 & ~n6095;
  assign n6097 = pi57 & pi59;
  assign n6098 = n3095 & n3294;
  assign n6099 = ~n3429 & ~n6098;
  assign n6100 = ~n6097 & ~n6099;
  assign n6101 = pi57 & ~n6100;
  assign n6102 = n3089 & n3207;
  assign n6103 = n3279 & n6102;
  assign n6104 = pi56 & ~n6103;
  assign n6105 = ~pi54 & n3277;
  assign n6106 = n6102 & n6105;
  assign n6107 = pi74 & ~n6106;
  assign n6108 = ~pi55 & ~n6107;
  assign n6109 = ~pi39 & n3089;
  assign n6110 = pi38 & ~n6109;
  assign n6111 = ~pi100 & ~n6110;
  assign n6112 = pi58 & n2521;
  assign n6113 = ~pi90 & ~n6112;
  assign n6114 = n2505 & n2578;
  assign n6115 = n2684 & n6114;
  assign n6116 = n2590 & ~n6115;
  assign n6117 = ~n2585 & ~n6116;
  assign n6118 = ~pi108 & ~n6117;
  assign n6119 = n2584 & ~n6118;
  assign n6120 = ~pi110 & n2699;
  assign n6121 = ~n6119 & n6120;
  assign n6122 = ~n2568 & ~n2575;
  assign n6123 = ~n6121 & n6122;
  assign n6124 = ~pi47 & ~n6123;
  assign n6125 = n2489 & ~n2571;
  assign n6126 = ~n6124 & n6125;
  assign n6127 = n6113 & ~n6126;
  assign n6128 = ~n2706 & ~n6127;
  assign n6129 = ~pi93 & ~n6128;
  assign n6130 = ~pi841 & n2522;
  assign n6131 = pi93 & ~n6130;
  assign n6132 = ~n6129 & ~n6131;
  assign n6133 = ~pi35 & ~n6132;
  assign n6134 = ~pi70 & ~n2524;
  assign n6135 = ~n6133 & n6134;
  assign n6136 = ~pi51 & ~n6135;
  assign n6137 = n2559 & ~n6136;
  assign n6138 = n2921 & ~n6137;
  assign n6139 = n2556 & ~n6138;
  assign n6140 = n2554 & ~n6139;
  assign n6141 = ~pi198 & ~pi299;
  assign n6142 = ~pi210 & pi299;
  assign n6143 = ~n6141 & ~n6142;
  assign n6144 = ~pi35 & n2551;
  assign n6145 = ~pi40 & n6144;
  assign n6146 = n2736 & n6145;
  assign n6147 = pi32 & ~n6146;
  assign n6148 = ~n6143 & ~n6147;
  assign n6149 = ~n3360 & n6143;
  assign n6150 = ~n6148 & ~n6149;
  assign n6151 = ~n6140 & ~n6150;
  assign n6152 = ~pi95 & ~n6151;
  assign n6153 = ~n2727 & ~n6152;
  assign n6154 = ~pi39 & ~n6153;
  assign n6155 = pi603 & ~pi642;
  assign n6156 = ~pi614 & ~pi616;
  assign n6157 = n6155 & n6156;
  assign n6158 = ~pi662 & pi680;
  assign n6159 = ~pi661 & n6158;
  assign n6160 = ~pi681 & n6159;
  assign po1101 = n6157 | n6160;
  assign n6162 = ~pi332 & ~pi468;
  assign n6163 = pi835 & pi984;
  assign n6164 = ~pi252 & ~pi1001;
  assign n6165 = ~pi979 & ~n6164;
  assign n6166 = ~n6163 & n6165;
  assign n6167 = ~pi287 & n6166;
  assign n6168 = pi835 & pi950;
  assign n6169 = n6167 & n6168;
  assign n6170 = pi1092 & n6169;
  assign n6171 = ~pi824 & ~pi829;
  assign n6172 = pi824 & ~pi1091;
  assign n6173 = pi1093 & ~n2734;
  assign n6174 = ~n6172 & n6173;
  assign n6175 = ~n6171 & ~n6174;
  assign n6176 = n6170 & n6175;
  assign n6177 = ~n6162 & ~n6176;
  assign n6178 = po1101 & ~n6177;
  assign n6179 = n3095 & ~n6178;
  assign n6180 = n3089 & n6162;
  assign n6181 = po1101 & n6180;
  assign n6182 = ~n6179 & ~n6181;
  assign n6183 = ~pi907 & ~pi947;
  assign n6184 = ~pi960 & ~pi963;
  assign n6185 = ~pi970 & ~pi972;
  assign n6186 = ~pi975 & ~pi978;
  assign n6187 = n6185 & n6186;
  assign n6188 = n6184 & n6187;
  assign n6189 = n6183 & n6188;
  assign n6190 = ~n6182 & n6189;
  assign n6191 = ~n6157 & ~n6162;
  assign n6192 = ~n6160 & n6191;
  assign n6193 = n6176 & ~n6192;
  assign n6194 = n3095 & ~n6193;
  assign n6195 = ~n6189 & n6194;
  assign n6196 = pi215 & ~n6195;
  assign n6197 = ~n6190 & n6196;
  assign n6198 = po1101 & ~n6162;
  assign n6199 = n6162 & ~n6189;
  assign n6200 = ~n6198 & ~n6199;
  assign n6201 = n2795 & n6169;
  assign n6202 = pi216 & pi221;
  assign n6203 = n6201 & n6202;
  assign n6204 = ~n6200 & n6203;
  assign n6205 = n3095 & ~n6204;
  assign n6206 = ~pi215 & ~n6205;
  assign n6207 = pi299 & ~n6206;
  assign n6208 = ~n6197 & n6207;
  assign n6209 = ~pi969 & ~pi971;
  assign n6210 = ~pi974 & ~pi977;
  assign n6211 = n6209 & n6210;
  assign n6212 = ~pi587 & ~pi602;
  assign n6213 = ~pi961 & ~pi967;
  assign n6214 = n6212 & n6213;
  assign n6215 = n6211 & n6214;
  assign n6216 = ~n6182 & n6215;
  assign n6217 = n6194 & ~n6215;
  assign n6218 = pi223 & ~n6217;
  assign n6219 = ~n6216 & n6218;
  assign n6220 = n6162 & ~n6215;
  assign n6221 = ~n6198 & ~n6220;
  assign n6222 = pi222 & pi224;
  assign n6223 = n6201 & n6222;
  assign n6224 = ~n6221 & n6223;
  assign n6225 = n3095 & ~n6224;
  assign n6226 = ~pi223 & ~n6225;
  assign n6227 = ~pi299 & ~n6226;
  assign n6228 = ~n6219 & n6227;
  assign n6229 = pi39 & ~n6228;
  assign n6230 = ~n6208 & n6229;
  assign n6231 = ~n6154 & ~n6230;
  assign n6232 = ~pi38 & ~n6231;
  assign n6233 = n6111 & ~n6232;
  assign n6234 = ~pi39 & n3095;
  assign n6235 = ~pi38 & pi100;
  assign n6236 = n6234 & n6235;
  assign n6237 = ~pi299 & ~n3063;
  assign n6238 = pi299 & ~n2448;
  assign n6239 = ~n6237 & ~n6238;
  assign n6240 = pi146 & n6238;
  assign n6241 = pi142 & n6237;
  assign n6242 = ~n6240 & ~n6241;
  assign n6243 = ~n6239 & n6242;
  assign n6244 = ~n3379 & ~n6243;
  assign n6245 = ~pi41 & ~pi99;
  assign n6246 = ~pi101 & n6245;
  assign n6247 = ~pi42 & ~pi43;
  assign n6248 = ~pi52 & n6247;
  assign n6249 = ~pi113 & ~pi116;
  assign n6250 = ~pi114 & ~pi115;
  assign n6251 = n6249 & n6250;
  assign n6252 = n6248 & n6251;
  assign n6253 = n6246 & n6252;
  assign po1057 = pi44 | ~n6253;
  assign n6255 = ~pi683 & po1057;
  assign n6256 = pi129 & pi250;
  assign n6257 = pi950 & pi1092;
  assign n6258 = ~n6171 & n6257;
  assign po740 = ~pi1093 & n6258;
  assign n6260 = ~pi250 & ~po740;
  assign n6261 = ~n6256 & ~n6260;
  assign n6262 = ~n6255 & ~n6261;
  assign n6263 = n6243 & po1057;
  assign n6264 = n6262 & n6263;
  assign n6265 = ~n6244 & ~n6264;
  assign n6266 = n6236 & n6265;
  assign n6267 = ~pi87 & ~n6266;
  assign n6268 = ~n6233 & n6267;
  assign n6269 = pi87 & ~n6102;
  assign n6270 = ~pi75 & ~n6269;
  assign n6271 = ~pi54 & ~pi92;
  assign n6272 = n6270 & n6271;
  assign n6273 = ~n6268 & n6272;
  assign n6274 = ~pi74 & ~n6273;
  assign n6275 = n6108 & ~n6274;
  assign n6276 = ~pi56 & ~n6275;
  assign n6277 = ~n6104 & ~n6276;
  assign n6278 = ~pi62 & ~n6277;
  assign n6279 = n3430 & n6102;
  assign n6280 = pi62 & ~n6279;
  assign n6281 = ~pi59 & ~n6280;
  assign n6282 = ~n6278 & n6281;
  assign n6283 = ~pi57 & ~n6282;
  assign po167 = ~n6101 & ~n6283;
  assign n6285 = ~pi55 & n3293;
  assign n6286 = ~pi59 & n6285;
  assign n6287 = ~pi228 & ~n6286;
  assign n6288 = pi57 & ~n6287;
  assign n6289 = ~n6160 & ~n6162;
  assign n6290 = ~pi907 & n6162;
  assign n6291 = ~n6289 & ~n6290;
  assign n6292 = ~pi228 & ~n3268;
  assign n6293 = pi30 & pi228;
  assign n6294 = ~n3321 & ~n6293;
  assign n6295 = ~n6292 & ~n6294;
  assign n6296 = n6291 & n6295;
  assign n6297 = n6288 & n6296;
  assign n6298 = ~pi602 & n6162;
  assign n6299 = ~n6289 & ~n6298;
  assign n6300 = ~pi91 & ~pi314;
  assign n6301 = n2574 & ~n2575;
  assign n6302 = pi85 & n2625;
  assign n6303 = n2458 & ~n6302;
  assign n6304 = n2629 & ~n6303;
  assign n6305 = n2467 & ~n6304;
  assign n6306 = ~n2609 & ~n2638;
  assign n6307 = ~n6305 & n6306;
  assign n6308 = n2468 & n6307;
  assign n6309 = ~n2643 & ~n6308;
  assign n6310 = n2641 & ~n6309;
  assign n6311 = pi67 & n2472;
  assign n6312 = n2606 & ~n6311;
  assign n6313 = ~n6310 & n6312;
  assign n6314 = n2605 & ~n6313;
  assign n6315 = ~pi71 & ~n6314;
  assign po1049 = pi64 | ~n2476;
  assign n6317 = n2600 & ~po1049;
  assign n6318 = ~n6315 & n6317;
  assign n6319 = ~pi81 & ~n6318;
  assign n6320 = n2654 & n6317;
  assign n6321 = n6319 & ~n6320;
  assign n6322 = ~pi102 & ~n2595;
  assign n6323 = n2452 & n6322;
  assign n6324 = ~n6321 & n6323;
  assign n6325 = n2594 & ~n6324;
  assign n6326 = n2687 & ~n6325;
  assign n6327 = n2504 & ~n6326;
  assign n6328 = ~n2507 & ~n6327;
  assign n6329 = ~pi86 & ~n6328;
  assign n6330 = ~pi46 & n2481;
  assign n6331 = n2592 & n6330;
  assign n6332 = ~n6329 & n6331;
  assign n6333 = n2699 & ~n6332;
  assign n6334 = n6301 & ~n6333;
  assign n6335 = n6300 & ~n6334;
  assign n6336 = pi91 & ~n2533;
  assign n6337 = ~pi58 & ~n6336;
  assign n6338 = ~pi91 & pi314;
  assign n6339 = ~n6319 & n6323;
  assign n6340 = n2594 & ~n6339;
  assign n6341 = n2687 & ~n6340;
  assign n6342 = n2504 & ~n6341;
  assign n6343 = ~n2507 & ~n6342;
  assign n6344 = ~pi86 & ~n6343;
  assign n6345 = n6331 & ~n6344;
  assign n6346 = n2699 & ~n6345;
  assign n6347 = n6301 & ~n6346;
  assign n6348 = n6338 & ~n6347;
  assign n6349 = n6337 & ~n6348;
  assign n6350 = ~n6335 & n6349;
  assign n6351 = ~pi90 & ~n6350;
  assign n6352 = ~n2706 & ~n6351;
  assign n6353 = ~pi93 & ~n6352;
  assign n6354 = pi93 & ~n2735;
  assign n6355 = ~pi35 & ~n6354;
  assign n6356 = ~n6353 & n6355;
  assign n6357 = ~pi70 & ~n6356;
  assign n6358 = n2844 & ~n6357;
  assign n6359 = ~pi72 & ~n6358;
  assign n6360 = ~pi95 & n2725;
  assign n6361 = ~n2555 & n6360;
  assign n6362 = ~n6359 & n6361;
  assign n6363 = ~n2938 & ~n6362;
  assign n6364 = ~pi841 & n2523;
  assign n6365 = n2535 & n6364;
  assign n6366 = n2783 & n6365;
  assign n6367 = pi32 & n6366;
  assign n6368 = ~pi95 & n6367;
  assign n6369 = ~pi198 & n6368;
  assign n6370 = n6363 & ~n6369;
  assign n6371 = ~pi228 & ~n6370;
  assign n6372 = ~n6293 & ~n6371;
  assign n6373 = n6299 & ~n6372;
  assign n6374 = ~pi299 & ~n6373;
  assign n6375 = pi145 & pi180;
  assign n6376 = pi181 & pi182;
  assign n6377 = n6375 & n6376;
  assign n6378 = ~pi299 & n6377;
  assign n6379 = ~n6374 & ~n6378;
  assign n6380 = n6293 & n6299;
  assign n6381 = ~n6162 & ~n6370;
  assign n6382 = ~pi47 & n2488;
  assign n6383 = ~n2698 & ~n6332;
  assign n6384 = n6382 & ~n6383;
  assign n6385 = n6300 & ~n6384;
  assign n6386 = ~n2698 & ~n6345;
  assign n6387 = n6382 & ~n6386;
  assign n6388 = n6338 & ~n6387;
  assign n6389 = n6337 & ~n6388;
  assign n6390 = ~n6385 & n6389;
  assign n6391 = ~pi90 & ~n6390;
  assign n6392 = ~n2706 & ~n6391;
  assign n6393 = ~pi93 & ~n6392;
  assign n6394 = n6355 & ~n6393;
  assign n6395 = ~pi70 & ~n6394;
  assign n6396 = n2844 & ~n6395;
  assign n6397 = ~pi72 & ~n6396;
  assign n6398 = n6361 & ~n6397;
  assign n6399 = ~n2938 & ~n6398;
  assign n6400 = ~n6369 & n6399;
  assign n6401 = n6162 & ~n6400;
  assign n6402 = ~n6381 & ~n6401;
  assign n6403 = ~pi228 & n6299;
  assign n6404 = ~n6402 & n6403;
  assign n6405 = ~n6380 & ~n6404;
  assign n6406 = n6377 & ~n6405;
  assign n6407 = ~n6379 & ~n6406;
  assign n6408 = n6291 & n6293;
  assign n6409 = pi299 & ~n6408;
  assign n6410 = pi158 & pi159;
  assign n6411 = pi160 & pi197;
  assign n6412 = n6410 & n6411;
  assign n6413 = ~pi210 & n6368;
  assign n6414 = n6363 & ~n6413;
  assign n6415 = ~n6162 & ~n6414;
  assign n6416 = n6399 & ~n6413;
  assign n6417 = n6162 & ~n6416;
  assign n6418 = ~n6415 & ~n6417;
  assign n6419 = n6291 & ~n6418;
  assign n6420 = n6412 & ~n6419;
  assign n6421 = n6291 & ~n6414;
  assign n6422 = ~n6412 & ~n6421;
  assign n6423 = ~pi228 & ~n6422;
  assign n6424 = ~n6420 & n6423;
  assign n6425 = n6409 & ~n6424;
  assign n6426 = pi232 & ~n6425;
  assign n6427 = ~n6407 & n6426;
  assign n6428 = ~pi228 & n6421;
  assign n6429 = n6409 & ~n6428;
  assign n6430 = ~pi232 & ~n6429;
  assign n6431 = ~n6374 & n6430;
  assign n6432 = ~n6427 & ~n6431;
  assign n6433 = ~pi39 & ~n6432;
  assign n6434 = ~pi215 & pi221;
  assign n6435 = ~pi287 & n3095;
  assign n6436 = pi835 & n6166;
  assign n6437 = n6435 & n6436;
  assign n6438 = pi824 & pi1093;
  assign n6439 = n6257 & n6438;
  assign n6440 = n6437 & n6439;
  assign n6441 = ~pi1091 & n6440;
  assign n6442 = pi1091 & n2733;
  assign n6443 = n6439 & ~n6442;
  assign n6444 = ~n2795 & ~n6443;
  assign n6445 = pi1091 & ~n6444;
  assign n6446 = n6437 & n6445;
  assign n6447 = ~n6441 & ~n6446;
  assign n6448 = pi216 & ~n6447;
  assign n6449 = ~pi829 & ~n2733;
  assign n6450 = pi1091 & ~n6449;
  assign n6451 = n6440 & ~n6450;
  assign n6452 = ~pi216 & n6451;
  assign n6453 = ~n6448 & ~n6452;
  assign n6454 = ~pi228 & ~n6453;
  assign n6455 = ~n6293 & ~n6454;
  assign n6456 = n6434 & ~n6455;
  assign n6457 = ~n6293 & ~n6456;
  assign n6458 = n6291 & ~n6457;
  assign n6459 = pi299 & ~n6458;
  assign n6460 = pi224 & n6447;
  assign n6461 = pi222 & ~pi223;
  assign n6462 = ~pi224 & ~n6451;
  assign n6463 = n6461 & ~n6462;
  assign n6464 = ~n6460 & n6463;
  assign n6465 = ~pi228 & n6464;
  assign n6466 = ~n6293 & ~n6465;
  assign n6467 = n6299 & ~n6466;
  assign n6468 = ~pi299 & ~n6467;
  assign n6469 = pi39 & ~n6468;
  assign n6470 = ~n6459 & n6469;
  assign n6471 = ~pi38 & ~n6470;
  assign n6472 = ~n6433 & n6471;
  assign n6473 = pi299 & n6291;
  assign n6474 = ~pi299 & n6299;
  assign n6475 = ~n6473 & ~n6474;
  assign n6476 = ~pi39 & ~n6294;
  assign n6477 = ~n6475 & n6476;
  assign n6478 = n6293 & ~n6475;
  assign n6479 = pi38 & ~n6478;
  assign n6480 = ~n6477 & n6479;
  assign n6481 = ~n6472 & ~n6480;
  assign n6482 = ~pi100 & ~n6481;
  assign n6483 = ~pi142 & ~n3063;
  assign n6484 = n3095 & ~n6261;
  assign n6485 = pi683 & po1057;
  assign n6486 = n6484 & n6485;
  assign n6487 = ~n6289 & n6486;
  assign n6488 = n6483 & n6487;
  assign n6489 = pi252 & ~n6483;
  assign n6490 = pi252 & n6180;
  assign n6491 = ~n6160 & n6490;
  assign n6492 = pi252 & n3095;
  assign n6493 = n6160 & n6492;
  assign n6494 = ~n6491 & ~n6493;
  assign n6495 = n6489 & ~n6494;
  assign n6496 = ~n6488 & ~n6495;
  assign n6497 = ~pi228 & ~n6298;
  assign n6498 = ~n6496 & n6497;
  assign n6499 = ~pi299 & ~n6380;
  assign n6500 = ~n6498 & n6499;
  assign n6501 = ~n2988 & n6494;
  assign n6502 = n2988 & ~n6487;
  assign n6503 = ~pi228 & ~n6290;
  assign n6504 = ~n6502 & n6503;
  assign n6505 = ~n6501 & n6504;
  assign n6506 = n6409 & ~n6505;
  assign n6507 = n3181 & ~n6506;
  assign n6508 = ~n6500 & n6507;
  assign n6509 = ~n3181 & n6478;
  assign n6510 = pi100 & ~n6509;
  assign n6511 = ~n6508 & n6510;
  assign n6512 = ~pi87 & ~n6511;
  assign n6513 = ~n6482 & n6512;
  assign n6514 = pi87 & n6478;
  assign n6515 = ~pi75 & ~n6514;
  assign n6516 = ~n6513 & n6515;
  assign n6517 = ~n3222 & n6478;
  assign n6518 = n3241 & n6477;
  assign n6519 = ~n6517 & ~n6518;
  assign n6520 = pi75 & n6519;
  assign n6521 = ~pi92 & ~n6520;
  assign n6522 = ~n6516 & n6521;
  assign n6523 = ~pi75 & n6519;
  assign n6524 = pi75 & ~n6478;
  assign n6525 = pi92 & ~n6524;
  assign n6526 = ~n6523 & n6525;
  assign n6527 = ~pi54 & ~n6526;
  assign n6528 = ~n6522 & n6527;
  assign n6529 = n3237 & n6519;
  assign n6530 = ~n3237 & ~n6478;
  assign n6531 = ~n6529 & ~n6530;
  assign n6532 = pi54 & ~n6531;
  assign n6533 = ~pi74 & ~n6532;
  assign n6534 = ~n6528 & n6533;
  assign n6535 = ~pi54 & n6529;
  assign n6536 = ~pi54 & n3237;
  assign n6537 = ~n6478 & ~n6536;
  assign n6538 = pi74 & ~n6537;
  assign n6539 = ~n6535 & n6538;
  assign n6540 = ~pi55 & ~n6539;
  assign n6541 = ~n6534 & n6540;
  assign n6542 = pi55 & ~n6296;
  assign n6543 = n3293 & ~n6542;
  assign n6544 = ~n6541 & n6543;
  assign n6545 = ~n3293 & n6408;
  assign n6546 = ~pi59 & ~n6545;
  assign n6547 = ~n6544 & n6546;
  assign n6548 = ~pi228 & ~n6285;
  assign n6549 = n6296 & ~n6548;
  assign n6550 = pi59 & ~n6549;
  assign n6551 = ~pi57 & ~n6550;
  assign n6552 = ~n6547 & n6551;
  assign po171 = ~n6297 & ~n6552;
  assign n6554 = ~pi947 & n6162;
  assign n6555 = ~n6191 & ~n6554;
  assign n6556 = n6295 & n6555;
  assign n6557 = n6288 & n6556;
  assign n6558 = ~pi587 & n6162;
  assign n6559 = ~n6191 & ~n6558;
  assign n6560 = n6293 & n6559;
  assign n6561 = ~pi228 & n6559;
  assign n6562 = ~n6402 & n6561;
  assign n6563 = ~n6560 & ~n6562;
  assign n6564 = n6377 & ~n6563;
  assign n6565 = ~n6372 & n6559;
  assign n6566 = ~n6377 & n6565;
  assign n6567 = ~pi299 & ~n6566;
  assign n6568 = ~n6564 & n6567;
  assign n6569 = n6293 & n6555;
  assign n6570 = pi299 & ~n6569;
  assign n6571 = ~n6418 & n6555;
  assign n6572 = n6412 & ~n6571;
  assign n6573 = ~n6414 & n6555;
  assign n6574 = ~n6412 & ~n6573;
  assign n6575 = ~pi228 & ~n6574;
  assign n6576 = ~n6572 & n6575;
  assign n6577 = n6570 & ~n6576;
  assign n6578 = pi232 & ~n6577;
  assign n6579 = ~n6568 & n6578;
  assign n6580 = ~pi299 & ~n6565;
  assign n6581 = ~pi228 & n6573;
  assign n6582 = n6570 & ~n6581;
  assign n6583 = ~pi232 & ~n6582;
  assign n6584 = ~n6580 & n6583;
  assign n6585 = ~n6579 & ~n6584;
  assign n6586 = ~pi39 & ~n6585;
  assign n6587 = pi299 & n6434;
  assign n6588 = ~n6570 & ~n6587;
  assign n6589 = n6456 & n6555;
  assign n6590 = ~n6588 & ~n6589;
  assign n6591 = ~n6466 & n6559;
  assign n6592 = ~pi299 & ~n6591;
  assign n6593 = pi39 & ~n6592;
  assign n6594 = ~n6590 & n6593;
  assign n6595 = ~pi38 & ~n6594;
  assign n6596 = ~n6586 & n6595;
  assign n6597 = pi299 & ~n6555;
  assign n6598 = ~pi299 & ~n6559;
  assign n6599 = ~n6597 & ~n6598;
  assign n6600 = n6476 & n6599;
  assign n6601 = n6293 & n6599;
  assign n6602 = pi38 & ~n6601;
  assign n6603 = ~n6600 & n6602;
  assign n6604 = ~n6596 & ~n6603;
  assign n6605 = ~pi100 & ~n6604;
  assign n6606 = ~pi228 & n3063;
  assign n6607 = ~n6157 & ~n6490;
  assign n6608 = n6157 & ~n6492;
  assign n6609 = ~n6607 & ~n6608;
  assign n6610 = ~n6558 & n6609;
  assign n6611 = n6606 & ~n6610;
  assign n6612 = pi142 & ~n6609;
  assign n6613 = ~n6191 & n6486;
  assign n6614 = ~pi142 & ~n6613;
  assign n6615 = n6157 & ~n6162;
  assign n6616 = ~pi587 & ~n6615;
  assign n6617 = ~pi228 & ~n6616;
  assign n6618 = ~n6614 & n6617;
  assign n6619 = ~n6612 & n6618;
  assign n6620 = ~n6560 & ~n6606;
  assign n6621 = ~n6619 & n6620;
  assign n6622 = ~n6611 & ~n6621;
  assign n6623 = ~pi299 & ~n6622;
  assign n6624 = n2988 & ~n6554;
  assign n6625 = n6613 & n6624;
  assign n6626 = ~pi947 & ~n6615;
  assign n6627 = ~n2988 & ~n6626;
  assign n6628 = n6609 & n6627;
  assign n6629 = ~n6625 & ~n6628;
  assign n6630 = ~pi228 & ~n6629;
  assign n6631 = n6570 & ~n6630;
  assign n6632 = n3181 & ~n6631;
  assign n6633 = ~n6623 & n6632;
  assign n6634 = ~n3181 & n6601;
  assign n6635 = pi100 & ~n6634;
  assign n6636 = ~n6633 & n6635;
  assign n6637 = ~pi87 & ~n6636;
  assign n6638 = ~n6605 & n6637;
  assign n6639 = pi87 & n6601;
  assign n6640 = ~pi75 & ~n6639;
  assign n6641 = ~n6638 & n6640;
  assign n6642 = ~n3222 & n6601;
  assign n6643 = n3241 & n6600;
  assign n6644 = ~n6642 & ~n6643;
  assign n6645 = pi75 & n6644;
  assign n6646 = ~pi92 & ~n6645;
  assign n6647 = ~n6641 & n6646;
  assign n6648 = ~pi75 & n6644;
  assign n6649 = pi75 & ~n6601;
  assign n6650 = pi92 & ~n6649;
  assign n6651 = ~n6648 & n6650;
  assign n6652 = ~pi54 & ~n6651;
  assign n6653 = ~n6647 & n6652;
  assign n6654 = n3237 & n6644;
  assign n6655 = ~n3237 & ~n6601;
  assign n6656 = ~n6654 & ~n6655;
  assign n6657 = pi54 & ~n6656;
  assign n6658 = ~pi74 & ~n6657;
  assign n6659 = ~n6653 & n6658;
  assign n6660 = ~pi54 & n6654;
  assign n6661 = ~n6536 & ~n6601;
  assign n6662 = pi74 & ~n6661;
  assign n6663 = ~n6660 & n6662;
  assign n6664 = ~pi55 & ~n6663;
  assign n6665 = ~n6659 & n6664;
  assign n6666 = pi55 & ~n6556;
  assign n6667 = n3293 & ~n6666;
  assign n6668 = ~n6665 & n6667;
  assign n6669 = ~n3293 & n6569;
  assign n6670 = ~pi59 & ~n6669;
  assign n6671 = ~n6668 & n6670;
  assign n6672 = ~n6548 & n6556;
  assign n6673 = pi59 & ~n6672;
  assign n6674 = ~pi57 & ~n6673;
  assign n6675 = ~n6671 & n6674;
  assign po172 = ~n6557 & ~n6675;
  assign n6677 = pi30 & n6162;
  assign n6678 = pi228 & n6677;
  assign n6679 = pi970 & n6678;
  assign n6680 = ~pi228 & pi970;
  assign n6681 = n6180 & n6680;
  assign n6682 = n3268 & n6681;
  assign n6683 = n6286 & n6682;
  assign n6684 = ~n6679 & ~n6683;
  assign n6685 = pi57 & ~n6684;
  assign n6686 = pi299 & ~n6679;
  assign n6687 = n6162 & ~n6414;
  assign n6688 = n6680 & n6687;
  assign n6689 = n6686 & ~n6688;
  assign n6690 = pi299 & n6410;
  assign n6691 = ~n6689 & ~n6690;
  assign n6692 = n6411 & ~n6417;
  assign n6693 = ~n6411 & n6414;
  assign n6694 = ~n6692 & ~n6693;
  assign n6695 = n6162 & n6694;
  assign n6696 = n6680 & n6695;
  assign n6697 = ~n6679 & ~n6696;
  assign n6698 = n6410 & ~n6697;
  assign n6699 = ~n6691 & ~n6698;
  assign n6700 = n6162 & ~n6372;
  assign n6701 = ~n6377 & ~n6700;
  assign n6702 = ~pi228 & n6401;
  assign n6703 = ~n6370 & ~n6377;
  assign n6704 = ~n6678 & ~n6703;
  assign n6705 = ~n6702 & n6704;
  assign n6706 = ~n6701 & ~n6705;
  assign n6707 = pi967 & n6706;
  assign n6708 = ~pi299 & ~n6707;
  assign n6709 = pi232 & ~n6708;
  assign n6710 = ~n6699 & n6709;
  assign n6711 = pi967 & n6700;
  assign n6712 = ~pi299 & ~n6711;
  assign n6713 = ~pi232 & ~n6689;
  assign n6714 = ~n6712 & n6713;
  assign n6715 = ~n6710 & ~n6714;
  assign n6716 = ~pi39 & ~n6715;
  assign n6717 = pi299 & pi970;
  assign n6718 = n6434 & ~n6453;
  assign n6719 = n6162 & n6718;
  assign n6720 = ~pi228 & ~n6719;
  assign n6721 = n6717 & ~n6720;
  assign n6722 = ~pi299 & pi967;
  assign n6723 = n6162 & n6464;
  assign n6724 = ~pi228 & ~n6723;
  assign n6725 = n6722 & ~n6724;
  assign n6726 = ~n6721 & ~n6725;
  assign n6727 = pi228 & ~n6677;
  assign n6728 = pi39 & ~n6727;
  assign n6729 = ~n6726 & n6728;
  assign n6730 = ~pi38 & ~n6729;
  assign n6731 = ~n6716 & n6730;
  assign n6732 = ~n6717 & ~n6722;
  assign n6733 = n6678 & ~n6732;
  assign n6734 = pi39 & n6733;
  assign n6735 = pi38 & ~n6734;
  assign n6736 = ~pi228 & ~n6180;
  assign n6737 = ~n6727 & ~n6736;
  assign n6738 = ~pi39 & ~n6732;
  assign n6739 = n6737 & n6738;
  assign n6740 = n6735 & ~n6739;
  assign n6741 = ~n6731 & ~n6740;
  assign n6742 = ~pi100 & ~n6741;
  assign n6743 = n6162 & n6486;
  assign n6744 = n6483 & n6743;
  assign n6745 = ~n6483 & n6490;
  assign n6746 = ~pi228 & ~n6745;
  assign n6747 = ~n6744 & n6746;
  assign n6748 = ~n6727 & ~n6747;
  assign n6749 = pi967 & n6748;
  assign n6750 = ~pi299 & ~n6749;
  assign n6751 = n2988 & ~n6743;
  assign n6752 = ~n2988 & ~n6490;
  assign n6753 = ~pi228 & ~n6752;
  assign n6754 = ~n6751 & n6753;
  assign n6755 = pi970 & n6754;
  assign n6756 = n6686 & ~n6755;
  assign n6757 = n3181 & ~n6756;
  assign n6758 = ~n6750 & n6757;
  assign n6759 = ~n3181 & n6733;
  assign n6760 = pi100 & ~n6759;
  assign n6761 = ~n6758 & n6760;
  assign n6762 = ~pi87 & ~n6761;
  assign n6763 = ~n6742 & n6762;
  assign n6764 = pi87 & n6733;
  assign n6765 = ~pi75 & ~n6764;
  assign n6766 = ~n6763 & n6765;
  assign n6767 = ~n3222 & n6733;
  assign n6768 = n3241 & n6739;
  assign n6769 = ~n6767 & ~n6768;
  assign n6770 = pi75 & n6769;
  assign n6771 = ~pi92 & ~n6770;
  assign n6772 = ~n6766 & n6771;
  assign n6773 = ~pi75 & n6769;
  assign n6774 = pi75 & ~n6733;
  assign n6775 = pi92 & ~n6774;
  assign n6776 = ~n6773 & n6775;
  assign n6777 = ~pi54 & ~n6776;
  assign n6778 = ~n6772 & n6777;
  assign n6779 = n3237 & n6769;
  assign n6780 = ~n3237 & ~n6733;
  assign n6781 = ~n6779 & ~n6780;
  assign n6782 = pi54 & ~n6781;
  assign n6783 = ~pi74 & ~n6782;
  assign n6784 = ~n6778 & n6783;
  assign n6785 = ~pi54 & n6779;
  assign n6786 = ~n6536 & ~n6733;
  assign n6787 = pi74 & ~n6786;
  assign n6788 = ~n6785 & n6787;
  assign n6789 = ~pi55 & ~n6788;
  assign n6790 = ~n6784 & n6789;
  assign n6791 = pi55 & ~n6679;
  assign n6792 = ~n6682 & n6791;
  assign n6793 = n3293 & ~n6792;
  assign n6794 = ~n6790 & n6793;
  assign n6795 = ~n3293 & n6679;
  assign n6796 = ~pi59 & ~n6795;
  assign n6797 = ~n6794 & n6796;
  assign n6798 = n6285 & n6682;
  assign n6799 = pi59 & ~n6679;
  assign n6800 = ~n6798 & n6799;
  assign n6801 = ~pi57 & ~n6800;
  assign n6802 = ~n6797 & n6801;
  assign po173 = ~n6685 & ~n6802;
  assign n6804 = pi972 & n6678;
  assign n6805 = ~pi228 & pi972;
  assign n6806 = n6180 & n6805;
  assign n6807 = n3268 & n6806;
  assign n6808 = n6286 & n6807;
  assign n6809 = ~n6804 & ~n6808;
  assign n6810 = pi57 & ~n6809;
  assign n6811 = pi299 & ~n6804;
  assign n6812 = n6687 & n6805;
  assign n6813 = n6811 & ~n6812;
  assign n6814 = ~n6690 & ~n6813;
  assign n6815 = n6695 & n6805;
  assign n6816 = ~n6804 & ~n6815;
  assign n6817 = n6410 & ~n6816;
  assign n6818 = ~n6814 & ~n6817;
  assign n6819 = pi961 & n6706;
  assign n6820 = ~pi299 & ~n6819;
  assign n6821 = pi232 & ~n6820;
  assign n6822 = ~n6818 & n6821;
  assign n6823 = pi961 & n6700;
  assign n6824 = ~pi299 & ~n6823;
  assign n6825 = ~pi232 & ~n6813;
  assign n6826 = ~n6824 & n6825;
  assign n6827 = ~n6822 & ~n6826;
  assign n6828 = ~pi39 & ~n6827;
  assign n6829 = ~pi299 & pi961;
  assign n6830 = ~n6724 & n6829;
  assign n6831 = pi299 & pi972;
  assign n6832 = ~n6720 & n6831;
  assign n6833 = ~n6830 & ~n6832;
  assign n6834 = n6728 & ~n6833;
  assign n6835 = ~pi38 & ~n6834;
  assign n6836 = ~n6828 & n6835;
  assign n6837 = ~n6829 & ~n6831;
  assign n6838 = n6678 & ~n6837;
  assign n6839 = pi39 & n6838;
  assign n6840 = pi38 & ~n6839;
  assign n6841 = ~pi39 & ~n6837;
  assign n6842 = n6737 & n6841;
  assign n6843 = n6840 & ~n6842;
  assign n6844 = ~n6836 & ~n6843;
  assign n6845 = ~pi100 & ~n6844;
  assign n6846 = pi961 & n6748;
  assign n6847 = ~pi299 & ~n6846;
  assign n6848 = pi972 & n6754;
  assign n6849 = n6811 & ~n6848;
  assign n6850 = n3181 & ~n6849;
  assign n6851 = ~n6847 & n6850;
  assign n6852 = ~n3181 & n6838;
  assign n6853 = pi100 & ~n6852;
  assign n6854 = ~n6851 & n6853;
  assign n6855 = ~pi87 & ~n6854;
  assign n6856 = ~n6845 & n6855;
  assign n6857 = pi87 & n6838;
  assign n6858 = ~pi75 & ~n6857;
  assign n6859 = ~n6856 & n6858;
  assign n6860 = ~n3222 & n6838;
  assign n6861 = n3241 & n6842;
  assign n6862 = ~n6860 & ~n6861;
  assign n6863 = pi75 & n6862;
  assign n6864 = ~pi92 & ~n6863;
  assign n6865 = ~n6859 & n6864;
  assign n6866 = ~pi75 & n6862;
  assign n6867 = pi75 & ~n6838;
  assign n6868 = pi92 & ~n6867;
  assign n6869 = ~n6866 & n6868;
  assign n6870 = ~pi54 & ~n6869;
  assign n6871 = ~n6865 & n6870;
  assign n6872 = n3237 & n6862;
  assign n6873 = ~n3237 & ~n6838;
  assign n6874 = ~n6872 & ~n6873;
  assign n6875 = pi54 & ~n6874;
  assign n6876 = ~pi74 & ~n6875;
  assign n6877 = ~n6871 & n6876;
  assign n6878 = ~pi54 & n6872;
  assign n6879 = ~n6536 & ~n6838;
  assign n6880 = pi74 & ~n6879;
  assign n6881 = ~n6878 & n6880;
  assign n6882 = ~pi55 & ~n6881;
  assign n6883 = ~n6877 & n6882;
  assign n6884 = pi55 & ~n6804;
  assign n6885 = ~n6807 & n6884;
  assign n6886 = n3293 & ~n6885;
  assign n6887 = ~n6883 & n6886;
  assign n6888 = ~n3293 & n6804;
  assign n6889 = ~pi59 & ~n6888;
  assign n6890 = ~n6887 & n6889;
  assign n6891 = n6285 & n6807;
  assign n6892 = pi59 & ~n6804;
  assign n6893 = ~n6891 & n6892;
  assign n6894 = ~pi57 & ~n6893;
  assign n6895 = ~n6890 & n6894;
  assign po174 = ~n6810 & ~n6895;
  assign n6897 = pi960 & n6678;
  assign n6898 = ~pi228 & pi960;
  assign n6899 = n6180 & n6898;
  assign n6900 = n3268 & n6899;
  assign n6901 = n6286 & n6900;
  assign n6902 = ~n6897 & ~n6901;
  assign n6903 = pi57 & ~n6902;
  assign n6904 = pi299 & ~n6897;
  assign n6905 = n6687 & n6898;
  assign n6906 = n6904 & ~n6905;
  assign n6907 = ~n6690 & ~n6906;
  assign n6908 = n6695 & n6898;
  assign n6909 = ~n6897 & ~n6908;
  assign n6910 = n6410 & ~n6909;
  assign n6911 = ~n6907 & ~n6910;
  assign n6912 = pi977 & n6706;
  assign n6913 = ~pi299 & ~n6912;
  assign n6914 = pi232 & ~n6913;
  assign n6915 = ~n6911 & n6914;
  assign n6916 = pi977 & n6700;
  assign n6917 = ~pi299 & ~n6916;
  assign n6918 = ~pi232 & ~n6906;
  assign n6919 = ~n6917 & n6918;
  assign n6920 = ~n6915 & ~n6919;
  assign n6921 = ~pi39 & ~n6920;
  assign n6922 = ~pi299 & pi977;
  assign n6923 = ~n6724 & n6922;
  assign n6924 = pi299 & pi960;
  assign n6925 = ~n6720 & n6924;
  assign n6926 = ~n6923 & ~n6925;
  assign n6927 = n6728 & ~n6926;
  assign n6928 = ~pi38 & ~n6927;
  assign n6929 = ~n6921 & n6928;
  assign n6930 = ~n6922 & ~n6924;
  assign n6931 = n6678 & ~n6930;
  assign n6932 = pi39 & n6931;
  assign n6933 = pi38 & ~n6932;
  assign n6934 = ~pi39 & ~n6930;
  assign n6935 = n6737 & n6934;
  assign n6936 = n6933 & ~n6935;
  assign n6937 = ~n6929 & ~n6936;
  assign n6938 = ~pi100 & ~n6937;
  assign n6939 = pi977 & n6748;
  assign n6940 = ~pi299 & ~n6939;
  assign n6941 = pi960 & n6754;
  assign n6942 = n6904 & ~n6941;
  assign n6943 = n3181 & ~n6942;
  assign n6944 = ~n6940 & n6943;
  assign n6945 = ~n3181 & n6931;
  assign n6946 = pi100 & ~n6945;
  assign n6947 = ~n6944 & n6946;
  assign n6948 = ~pi87 & ~n6947;
  assign n6949 = ~n6938 & n6948;
  assign n6950 = pi87 & n6931;
  assign n6951 = ~pi75 & ~n6950;
  assign n6952 = ~n6949 & n6951;
  assign n6953 = ~n3222 & n6931;
  assign n6954 = n3241 & n6935;
  assign n6955 = ~n6953 & ~n6954;
  assign n6956 = pi75 & n6955;
  assign n6957 = ~pi92 & ~n6956;
  assign n6958 = ~n6952 & n6957;
  assign n6959 = ~pi75 & n6955;
  assign n6960 = pi75 & ~n6931;
  assign n6961 = pi92 & ~n6960;
  assign n6962 = ~n6959 & n6961;
  assign n6963 = ~pi54 & ~n6962;
  assign n6964 = ~n6958 & n6963;
  assign n6965 = n3237 & n6955;
  assign n6966 = ~n3237 & ~n6931;
  assign n6967 = ~n6965 & ~n6966;
  assign n6968 = pi54 & ~n6967;
  assign n6969 = ~pi74 & ~n6968;
  assign n6970 = ~n6964 & n6969;
  assign n6971 = ~pi54 & n6965;
  assign n6972 = ~n6536 & ~n6931;
  assign n6973 = pi74 & ~n6972;
  assign n6974 = ~n6971 & n6973;
  assign n6975 = ~pi55 & ~n6974;
  assign n6976 = ~n6970 & n6975;
  assign n6977 = pi55 & ~n6897;
  assign n6978 = ~n6900 & n6977;
  assign n6979 = n3293 & ~n6978;
  assign n6980 = ~n6976 & n6979;
  assign n6981 = ~n3293 & n6897;
  assign n6982 = ~pi59 & ~n6981;
  assign n6983 = ~n6980 & n6982;
  assign n6984 = n6285 & n6900;
  assign n6985 = pi59 & ~n6897;
  assign n6986 = ~n6984 & n6985;
  assign n6987 = ~pi57 & ~n6986;
  assign n6988 = ~n6983 & n6987;
  assign po175 = ~n6903 & ~n6988;
  assign n6990 = pi963 & n6678;
  assign n6991 = ~pi228 & pi963;
  assign n6992 = n6180 & n6991;
  assign n6993 = n3268 & n6992;
  assign n6994 = n6286 & n6993;
  assign n6995 = ~n6990 & ~n6994;
  assign n6996 = pi57 & ~n6995;
  assign n6997 = pi299 & ~n6990;
  assign n6998 = n6687 & n6991;
  assign n6999 = n6997 & ~n6998;
  assign n7000 = ~n6690 & ~n6999;
  assign n7001 = n6695 & n6991;
  assign n7002 = ~n6990 & ~n7001;
  assign n7003 = n6410 & ~n7002;
  assign n7004 = ~n7000 & ~n7003;
  assign n7005 = pi969 & n6706;
  assign n7006 = ~pi299 & ~n7005;
  assign n7007 = pi232 & ~n7006;
  assign n7008 = ~n7004 & n7007;
  assign n7009 = pi969 & n6700;
  assign n7010 = ~pi299 & ~n7009;
  assign n7011 = ~pi232 & ~n6999;
  assign n7012 = ~n7010 & n7011;
  assign n7013 = ~n7008 & ~n7012;
  assign n7014 = ~pi39 & ~n7013;
  assign n7015 = ~pi299 & pi969;
  assign n7016 = ~n6724 & n7015;
  assign n7017 = pi299 & pi963;
  assign n7018 = ~n6720 & n7017;
  assign n7019 = ~n7016 & ~n7018;
  assign n7020 = n6728 & ~n7019;
  assign n7021 = ~pi38 & ~n7020;
  assign n7022 = ~n7014 & n7021;
  assign n7023 = ~n7015 & ~n7017;
  assign n7024 = n6678 & ~n7023;
  assign n7025 = pi39 & n7024;
  assign n7026 = pi38 & ~n7025;
  assign n7027 = ~pi39 & ~n7023;
  assign n7028 = n6737 & n7027;
  assign n7029 = n7026 & ~n7028;
  assign n7030 = ~n7022 & ~n7029;
  assign n7031 = ~pi100 & ~n7030;
  assign n7032 = pi969 & n6748;
  assign n7033 = ~pi299 & ~n7032;
  assign n7034 = pi963 & n6754;
  assign n7035 = n6997 & ~n7034;
  assign n7036 = n3181 & ~n7035;
  assign n7037 = ~n7033 & n7036;
  assign n7038 = ~n3181 & n7024;
  assign n7039 = pi100 & ~n7038;
  assign n7040 = ~n7037 & n7039;
  assign n7041 = ~pi87 & ~n7040;
  assign n7042 = ~n7031 & n7041;
  assign n7043 = pi87 & n7024;
  assign n7044 = ~pi75 & ~n7043;
  assign n7045 = ~n7042 & n7044;
  assign n7046 = ~n3222 & n7024;
  assign n7047 = n3241 & n7028;
  assign n7048 = ~n7046 & ~n7047;
  assign n7049 = pi75 & n7048;
  assign n7050 = ~pi92 & ~n7049;
  assign n7051 = ~n7045 & n7050;
  assign n7052 = ~pi75 & n7048;
  assign n7053 = pi75 & ~n7024;
  assign n7054 = pi92 & ~n7053;
  assign n7055 = ~n7052 & n7054;
  assign n7056 = ~pi54 & ~n7055;
  assign n7057 = ~n7051 & n7056;
  assign n7058 = n3237 & n7048;
  assign n7059 = ~n3237 & ~n7024;
  assign n7060 = ~n7058 & ~n7059;
  assign n7061 = pi54 & ~n7060;
  assign n7062 = ~pi74 & ~n7061;
  assign n7063 = ~n7057 & n7062;
  assign n7064 = ~pi54 & n7058;
  assign n7065 = ~n6536 & ~n7024;
  assign n7066 = pi74 & ~n7065;
  assign n7067 = ~n7064 & n7066;
  assign n7068 = ~pi55 & ~n7067;
  assign n7069 = ~n7063 & n7068;
  assign n7070 = pi55 & ~n6990;
  assign n7071 = ~n6993 & n7070;
  assign n7072 = n3293 & ~n7071;
  assign n7073 = ~n7069 & n7072;
  assign n7074 = ~n3293 & n6990;
  assign n7075 = ~pi59 & ~n7074;
  assign n7076 = ~n7073 & n7075;
  assign n7077 = n6285 & n6993;
  assign n7078 = pi59 & ~n6990;
  assign n7079 = ~n7077 & n7078;
  assign n7080 = ~pi57 & ~n7079;
  assign n7081 = ~n7076 & n7080;
  assign po176 = ~n6996 & ~n7081;
  assign n7083 = pi975 & n6678;
  assign n7084 = ~pi228 & pi975;
  assign n7085 = n6180 & n7084;
  assign n7086 = n3268 & n7085;
  assign n7087 = n6286 & n7086;
  assign n7088 = ~n7083 & ~n7087;
  assign n7089 = pi57 & ~n7088;
  assign n7090 = pi299 & ~n7083;
  assign n7091 = n6687 & n7084;
  assign n7092 = n7090 & ~n7091;
  assign n7093 = ~n6690 & ~n7092;
  assign n7094 = n6695 & n7084;
  assign n7095 = ~n7083 & ~n7094;
  assign n7096 = n6410 & ~n7095;
  assign n7097 = ~n7093 & ~n7096;
  assign n7098 = pi971 & n6706;
  assign n7099 = ~pi299 & ~n7098;
  assign n7100 = pi232 & ~n7099;
  assign n7101 = ~n7097 & n7100;
  assign n7102 = pi971 & n6700;
  assign n7103 = ~pi299 & ~n7102;
  assign n7104 = ~pi232 & ~n7092;
  assign n7105 = ~n7103 & n7104;
  assign n7106 = ~n7101 & ~n7105;
  assign n7107 = ~pi39 & ~n7106;
  assign n7108 = ~pi299 & pi971;
  assign n7109 = ~n6724 & n7108;
  assign n7110 = pi299 & pi975;
  assign n7111 = ~n6720 & n7110;
  assign n7112 = ~n7109 & ~n7111;
  assign n7113 = n6728 & ~n7112;
  assign n7114 = ~pi38 & ~n7113;
  assign n7115 = ~n7107 & n7114;
  assign n7116 = ~n7108 & ~n7110;
  assign n7117 = n6678 & ~n7116;
  assign n7118 = pi39 & n7117;
  assign n7119 = pi38 & ~n7118;
  assign n7120 = ~pi39 & ~n7116;
  assign n7121 = n6737 & n7120;
  assign n7122 = n7119 & ~n7121;
  assign n7123 = ~n7115 & ~n7122;
  assign n7124 = ~pi100 & ~n7123;
  assign n7125 = pi971 & n6748;
  assign n7126 = ~pi299 & ~n7125;
  assign n7127 = pi975 & n6754;
  assign n7128 = n7090 & ~n7127;
  assign n7129 = n3181 & ~n7128;
  assign n7130 = ~n7126 & n7129;
  assign n7131 = ~n3181 & n7117;
  assign n7132 = pi100 & ~n7131;
  assign n7133 = ~n7130 & n7132;
  assign n7134 = ~pi87 & ~n7133;
  assign n7135 = ~n7124 & n7134;
  assign n7136 = pi87 & n7117;
  assign n7137 = ~pi75 & ~n7136;
  assign n7138 = ~n7135 & n7137;
  assign n7139 = ~n3222 & n7117;
  assign n7140 = n3241 & n7121;
  assign n7141 = ~n7139 & ~n7140;
  assign n7142 = pi75 & n7141;
  assign n7143 = ~pi92 & ~n7142;
  assign n7144 = ~n7138 & n7143;
  assign n7145 = ~pi75 & n7141;
  assign n7146 = pi75 & ~n7117;
  assign n7147 = pi92 & ~n7146;
  assign n7148 = ~n7145 & n7147;
  assign n7149 = ~pi54 & ~n7148;
  assign n7150 = ~n7144 & n7149;
  assign n7151 = n3237 & n7141;
  assign n7152 = ~n3237 & ~n7117;
  assign n7153 = ~n7151 & ~n7152;
  assign n7154 = pi54 & ~n7153;
  assign n7155 = ~pi74 & ~n7154;
  assign n7156 = ~n7150 & n7155;
  assign n7157 = ~pi54 & n7151;
  assign n7158 = ~n6536 & ~n7117;
  assign n7159 = pi74 & ~n7158;
  assign n7160 = ~n7157 & n7159;
  assign n7161 = ~pi55 & ~n7160;
  assign n7162 = ~n7156 & n7161;
  assign n7163 = pi55 & ~n7083;
  assign n7164 = ~n7086 & n7163;
  assign n7165 = n3293 & ~n7164;
  assign n7166 = ~n7162 & n7165;
  assign n7167 = ~n3293 & n7083;
  assign n7168 = ~pi59 & ~n7167;
  assign n7169 = ~n7166 & n7168;
  assign n7170 = n6285 & n7086;
  assign n7171 = pi59 & ~n7083;
  assign n7172 = ~n7170 & n7171;
  assign n7173 = ~pi57 & ~n7172;
  assign n7174 = ~n7169 & n7173;
  assign po177 = ~n7089 & ~n7174;
  assign n7176 = pi978 & n6678;
  assign n7177 = ~pi228 & pi978;
  assign n7178 = n3268 & n7177;
  assign n7179 = n6180 & n7178;
  assign n7180 = n6286 & n7179;
  assign n7181 = ~n7176 & ~n7180;
  assign n7182 = pi57 & ~n7181;
  assign n7183 = ~pi299 & pi974;
  assign n7184 = pi299 & pi978;
  assign n7185 = ~n7183 & ~n7184;
  assign n7186 = n6737 & ~n7185;
  assign n7187 = ~pi39 & n7186;
  assign n7188 = n6678 & ~n7185;
  assign n7189 = pi39 & n7188;
  assign n7190 = pi38 & ~n7189;
  assign n7191 = ~n7187 & n7190;
  assign n7192 = pi299 & ~n7176;
  assign n7193 = n6687 & n7177;
  assign n7194 = n7192 & ~n7193;
  assign n7195 = ~n6690 & ~n7194;
  assign n7196 = n6695 & n7177;
  assign n7197 = ~n7176 & ~n7196;
  assign n7198 = n6410 & ~n7197;
  assign n7199 = ~n7195 & ~n7198;
  assign n7200 = pi974 & n6706;
  assign n7201 = ~pi299 & ~n7200;
  assign n7202 = pi232 & ~n7201;
  assign n7203 = ~n7199 & n7202;
  assign n7204 = pi974 & n6700;
  assign n7205 = ~pi299 & ~n7204;
  assign n7206 = ~pi232 & ~n7194;
  assign n7207 = ~n7205 & n7206;
  assign n7208 = ~n7203 & ~n7207;
  assign n7209 = ~pi39 & ~n7208;
  assign n7210 = ~n6724 & n7183;
  assign n7211 = ~n6720 & n7184;
  assign n7212 = ~n7210 & ~n7211;
  assign n7213 = n6728 & ~n7212;
  assign n7214 = ~pi38 & ~n7213;
  assign n7215 = ~n7209 & n7214;
  assign n7216 = ~n7191 & ~n7215;
  assign n7217 = ~pi100 & ~n7216;
  assign n7218 = pi974 & n6748;
  assign n7219 = ~pi299 & ~n7218;
  assign n7220 = pi978 & n6754;
  assign n7221 = n7192 & ~n7220;
  assign n7222 = n3181 & ~n7221;
  assign n7223 = ~n7219 & n7222;
  assign n7224 = ~n3181 & n7188;
  assign n7225 = pi100 & ~n7224;
  assign n7226 = ~n7223 & n7225;
  assign n7227 = ~pi87 & ~n7226;
  assign n7228 = ~n7217 & n7227;
  assign n7229 = pi87 & n7188;
  assign n7230 = ~pi75 & ~n7229;
  assign n7231 = ~n7228 & n7230;
  assign n7232 = ~pi228 & ~n3222;
  assign n7233 = n7186 & ~n7232;
  assign n7234 = pi75 & ~n7233;
  assign n7235 = ~pi92 & ~n7234;
  assign n7236 = ~n7231 & n7235;
  assign n7237 = ~pi75 & ~n7233;
  assign n7238 = pi75 & ~n7188;
  assign n7239 = pi92 & ~n7238;
  assign n7240 = ~n7237 & n7239;
  assign n7241 = ~pi54 & ~n7240;
  assign n7242 = ~n7236 & n7241;
  assign n7243 = n3237 & ~n7233;
  assign n7244 = ~n3237 & ~n7188;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = pi54 & ~n7245;
  assign n7247 = ~pi74 & ~n7246;
  assign n7248 = ~n7242 & n7247;
  assign n7249 = ~pi54 & n7243;
  assign n7250 = ~n6536 & ~n7188;
  assign n7251 = pi74 & ~n7250;
  assign n7252 = ~n7249 & n7251;
  assign n7253 = ~pi55 & ~n7252;
  assign n7254 = ~n7248 & n7253;
  assign n7255 = pi55 & ~n7176;
  assign n7256 = ~n7179 & n7255;
  assign n7257 = n3293 & ~n7256;
  assign n7258 = ~n7254 & n7257;
  assign n7259 = ~n3293 & n7176;
  assign n7260 = ~pi59 & ~n7259;
  assign n7261 = ~n7258 & n7260;
  assign n7262 = n6285 & n7179;
  assign n7263 = pi59 & ~n7176;
  assign n7264 = ~n7262 & n7263;
  assign n7265 = ~pi57 & ~n7264;
  assign n7266 = ~n7261 & n7265;
  assign po178 = ~n7182 & ~n7266;
  assign n7268 = n3241 & n6234;
  assign n7269 = pi75 & ~n7268;
  assign n7270 = n3206 & n3230;
  assign n7271 = n6234 & n7270;
  assign n7272 = pi92 & ~n7271;
  assign n7273 = ~n7269 & ~n7272;
  assign n7274 = pi299 & ~n6200;
  assign n7275 = n6718 & n7274;
  assign n7276 = ~pi299 & ~n6221;
  assign n7277 = n6464 & n7276;
  assign n7278 = pi39 & ~n7277;
  assign n7279 = ~n7275 & n7278;
  assign n7280 = ~n6415 & n6690;
  assign n7281 = ~n6694 & n7280;
  assign n7282 = n6377 & n6401;
  assign n7283 = ~pi299 & ~n6381;
  assign n7284 = ~n6703 & n7283;
  assign n7285 = ~n7282 & n7284;
  assign n7286 = pi299 & n6414;
  assign n7287 = ~n6410 & n7286;
  assign n7288 = pi232 & ~n7287;
  assign n7289 = ~n7285 & n7288;
  assign n7290 = ~n7281 & n7289;
  assign n7291 = ~pi299 & n6370;
  assign n7292 = ~pi232 & ~n7286;
  assign n7293 = ~n7291 & n7292;
  assign n7294 = ~pi39 & ~n7293;
  assign n7295 = ~n7290 & n7294;
  assign n7296 = ~n7279 & ~n7295;
  assign n7297 = ~pi38 & ~n7296;
  assign n7298 = ~n6110 & ~n7297;
  assign n7299 = ~pi100 & ~n7298;
  assign n7300 = ~pi38 & n6234;
  assign n7301 = pi100 & ~n7300;
  assign n7302 = n6267 & ~n7301;
  assign n7303 = ~n7299 & n7302;
  assign n7304 = n3237 & ~n7303;
  assign n7305 = n7273 & ~n7304;
  assign n7306 = ~pi54 & ~n7305;
  assign n7307 = ~pi92 & n7271;
  assign n7308 = pi54 & ~n7307;
  assign n7309 = ~n7306 & ~n7308;
  assign n7310 = ~pi74 & ~n7309;
  assign n7311 = ~n6107 & ~n7310;
  assign n7312 = ~pi55 & ~n7311;
  assign n7313 = n3278 & n6102;
  assign n7314 = pi55 & ~n7313;
  assign n7315 = ~pi56 & ~n7314;
  assign n7316 = ~pi62 & n7315;
  assign n7317 = ~n7312 & n7316;
  assign n7318 = n3429 & ~n7317;
  assign po195 = n6100 & ~n7318;
  assign n7320 = ~pi954 & ~po195;
  assign n7321 = pi24 & pi954;
  assign po182 = ~n7320 & ~n7321;
  assign n7323 = n3276 & n3321;
  assign n7324 = n3430 & n7323;
  assign n7325 = ~n3126 & ~n7324;
  assign n7326 = pi62 & ~n7325;
  assign n7327 = ~pi100 & n4669;
  assign n7328 = n3095 & ~n6489;
  assign n7329 = ~pi299 & ~n7328;
  assign n7330 = pi299 & ~n3388;
  assign n7331 = ~n7329 & ~n7330;
  assign n7332 = pi100 & n3321;
  assign n7333 = n7331 & n7332;
  assign n7334 = ~pi39 & ~n7333;
  assign n7335 = ~n7327 & n7334;
  assign n7336 = ~pi100 & n3321;
  assign n7337 = pi39 & ~n7336;
  assign n7338 = ~pi38 & ~n7337;
  assign n7339 = ~n7335 & n7338;
  assign n7340 = ~n3126 & ~n7339;
  assign n7341 = ~pi87 & ~n7340;
  assign n7342 = ~n3126 & ~n7323;
  assign n7343 = pi87 & ~n7342;
  assign n7344 = ~pi75 & ~n7343;
  assign n7345 = ~n7341 & n7344;
  assign n7346 = pi75 & ~n3126;
  assign n7347 = ~pi92 & ~n7346;
  assign n7348 = ~n7345 & n7347;
  assign n7349 = n3321 & n3406;
  assign n7350 = ~n3126 & ~n7349;
  assign n7351 = pi92 & ~n7350;
  assign n7352 = n3265 & ~n7351;
  assign n7353 = ~n7348 & n7352;
  assign n7354 = ~n3126 & ~n3265;
  assign n7355 = ~pi55 & ~n7354;
  assign n7356 = ~n7353 & n7355;
  assign n7357 = n3276 & n6105;
  assign n7358 = n3321 & n7357;
  assign n7359 = ~pi74 & n7358;
  assign n7360 = ~n3126 & ~n7359;
  assign n7361 = pi55 & ~n7360;
  assign n7362 = ~pi56 & ~n7361;
  assign n7363 = ~n7356 & n7362;
  assign n7364 = n3280 & n3321;
  assign n7365 = pi56 & ~n3126;
  assign n7366 = ~n7364 & n7365;
  assign n7367 = ~pi62 & ~n7366;
  assign n7368 = ~n7363 & n7367;
  assign n7369 = ~n7326 & ~n7368;
  assign n7370 = n3429 & ~n7369;
  assign n7371 = n3126 & ~n3429;
  assign po183 = n7370 | n7371;
  assign n7373 = pi119 & pi1056;
  assign n7374 = ~pi228 & pi252;
  assign n7375 = ~pi119 & ~n7374;
  assign n7376 = ~pi468 & ~n7375;
  assign po184 = n7373 | ~n7376;
  assign n7378 = pi119 & pi1077;
  assign po185 = ~n7376 | n7378;
  assign n7380 = pi119 & pi1073;
  assign po186 = ~n7376 | n7380;
  assign n7382 = pi119 & pi1041;
  assign po187 = ~n7376 | n7382;
  assign n7384 = pi360 & ~pi462;
  assign n7385 = ~pi360 & pi462;
  assign n7386 = ~n7384 & ~n7385;
  assign n7387 = pi352 & ~pi353;
  assign n7388 = ~pi352 & pi353;
  assign n7389 = ~n7387 & ~n7388;
  assign n7390 = n7386 & n7389;
  assign n7391 = ~n7386 & ~n7389;
  assign n7392 = ~n7390 & ~n7391;
  assign n7393 = pi354 & ~n7392;
  assign n7394 = ~pi354 & n7392;
  assign n7395 = ~n7393 & ~n7394;
  assign n7396 = pi351 & pi1199;
  assign n7397 = pi345 & ~pi346;
  assign n7398 = ~pi345 & pi346;
  assign n7399 = ~n7397 & ~n7398;
  assign n7400 = pi323 & ~n7399;
  assign n7401 = ~pi323 & n7399;
  assign n7402 = ~n7400 & ~n7401;
  assign n7403 = pi358 & ~pi450;
  assign n7404 = ~pi358 & pi450;
  assign n7405 = ~n7403 & ~n7404;
  assign n7406 = n7402 & ~n7405;
  assign n7407 = ~n7402 & n7405;
  assign n7408 = ~n7406 & ~n7407;
  assign n7409 = ~pi327 & ~pi362;
  assign n7410 = pi327 & pi362;
  assign n7411 = ~n7409 & ~n7410;
  assign n7412 = pi343 & ~pi344;
  assign n7413 = ~pi343 & pi344;
  assign n7414 = ~n7412 & ~n7413;
  assign n7415 = n7411 & ~n7414;
  assign n7416 = ~n7411 & n7414;
  assign n7417 = ~n7415 & ~n7416;
  assign n7418 = ~n7408 & ~n7417;
  assign n7419 = n7408 & n7417;
  assign n7420 = pi1197 & ~n7419;
  assign n7421 = ~n7418 & n7420;
  assign n7422 = ~pi74 & n6271;
  assign n7423 = n2534 & ~n6131;
  assign n7424 = ~pi841 & n2492;
  assign n7425 = pi90 & n7424;
  assign n7426 = ~pi93 & ~n7425;
  assign n7427 = n7423 & ~n7426;
  assign n7428 = ~pi51 & ~n7427;
  assign n7429 = ~pi50 & ~pi77;
  assign n7430 = ~pi94 & n7429;
  assign n7431 = n2576 & n7430;
  assign n7432 = ~pi88 & pi98;
  assign n7433 = n2484 & n7432;
  assign n7434 = n7431 & n7433;
  assign n7435 = ~pi97 & ~n7434;
  assign n7436 = n2514 & ~n7435;
  assign n7437 = ~pi35 & n2493;
  assign n7438 = ~pi70 & n7437;
  assign n7439 = n7436 & n7438;
  assign n7440 = n7428 & ~n7439;
  assign n7441 = ~n2558 & ~n7440;
  assign n7442 = ~pi96 & n3093;
  assign n7443 = n7441 & n7442;
  assign n7444 = n6258 & n7443;
  assign n7445 = ~pi96 & ~n7441;
  assign n7446 = pi96 & ~n6365;
  assign n7447 = n3093 & ~n7446;
  assign n7448 = ~pi122 & pi829;
  assign n7449 = n6257 & n7448;
  assign n7450 = n7447 & n7449;
  assign n7451 = ~n7445 & n7450;
  assign n7452 = ~n7444 & ~n7451;
  assign n7453 = ~pi1093 & ~n7452;
  assign n7454 = ~pi87 & ~n7453;
  assign n7455 = n3095 & po740;
  assign n7456 = pi87 & ~n7455;
  assign n7457 = ~pi75 & n3276;
  assign n7458 = ~n7456 & n7457;
  assign n7459 = ~n7454 & n7458;
  assign n7460 = ~pi567 & ~n7459;
  assign n7461 = n7422 & ~n7460;
  assign n7462 = pi232 & n6162;
  assign n7463 = n6239 & n7462;
  assign n7464 = n3222 & ~n7463;
  assign n7465 = ~pi24 & n6492;
  assign n7466 = ~n2733 & po1057;
  assign n7467 = pi1091 & n7466;
  assign n7468 = n7449 & n7467;
  assign n7469 = n7465 & n7468;
  assign n7470 = pi1093 & n7469;
  assign n7471 = n7464 & n7470;
  assign n7472 = pi75 & ~n7471;
  assign n7473 = pi1093 & ~n2733;
  assign n7474 = pi824 & n6257;
  assign n7475 = ~n2558 & n7442;
  assign n7476 = ~n7428 & n7475;
  assign n7477 = n7474 & n7476;
  assign n7478 = ~pi829 & n7477;
  assign n7479 = ~pi24 & n2565;
  assign n7480 = ~pi46 & pi97;
  assign n7481 = ~pi108 & n7480;
  assign n7482 = n6382 & n7481;
  assign n7483 = n2581 & n7482;
  assign n7484 = ~pi91 & n7483;
  assign n7485 = ~n7479 & ~n7484;
  assign n7486 = n2518 & n7423;
  assign n7487 = ~n7485 & n7486;
  assign n7488 = n7428 & ~n7487;
  assign n7489 = ~n2558 & ~n7488;
  assign n7490 = ~pi96 & ~n7489;
  assign n7491 = pi829 & n6257;
  assign n7492 = n7447 & n7491;
  assign n7493 = ~n7490 & n7492;
  assign n7494 = ~n7478 & ~n7493;
  assign n7495 = ~pi122 & ~n7494;
  assign n7496 = pi122 & n6258;
  assign n7497 = n7476 & n7496;
  assign n7498 = ~n7495 & ~n7497;
  assign n7499 = n7473 & ~n7498;
  assign n7500 = pi1091 & ~n7499;
  assign n7501 = ~n7453 & n7500;
  assign n7502 = ~pi1091 & ~n7453;
  assign n7503 = ~n7501 & ~n7502;
  assign n7504 = ~pi39 & ~n7503;
  assign n7505 = ~n2733 & n2753;
  assign n7506 = n6437 & n7505;
  assign n7507 = n2754 & n7506;
  assign n7508 = pi1091 & n7507;
  assign n7509 = ~n6221 & n7508;
  assign n7510 = ~pi299 & n6461;
  assign n7511 = ~pi224 & n7510;
  assign n7512 = n7509 & n7511;
  assign n7513 = ~n6200 & n7508;
  assign n7514 = ~pi216 & n6587;
  assign n7515 = n7513 & n7514;
  assign n7516 = pi39 & ~n7515;
  assign n7517 = ~n7512 & n7516;
  assign n7518 = ~pi38 & ~n7517;
  assign n7519 = ~n7504 & n7518;
  assign n7520 = ~pi100 & ~n7519;
  assign n7521 = n6439 & n7476;
  assign n7522 = n7518 & n7521;
  assign n7523 = ~n7500 & n7522;
  assign n7524 = n7520 & ~n7523;
  assign n7525 = pi1093 & n7449;
  assign n7526 = n7466 & n7525;
  assign n7527 = n3095 & n7526;
  assign n7528 = pi1091 & n7527;
  assign n7529 = pi228 & n7528;
  assign n7530 = n3181 & ~n7463;
  assign n7531 = n7529 & n7530;
  assign n7532 = pi100 & ~n7531;
  assign n7533 = ~n7524 & ~n7532;
  assign n7534 = ~pi87 & ~n7533;
  assign n7535 = n3095 & n7474;
  assign n7536 = ~pi1091 & pi1093;
  assign n7537 = ~n7535 & n7536;
  assign n7538 = pi1093 & n2733;
  assign n7539 = n6258 & ~n7538;
  assign n7540 = n3095 & n7539;
  assign n7541 = ~n7536 & ~n7540;
  assign n7542 = n3207 & ~n7541;
  assign n7543 = ~n7537 & n7542;
  assign n7544 = pi87 & ~n7543;
  assign n7545 = ~n7534 & ~n7544;
  assign n7546 = ~pi75 & ~n7545;
  assign n7547 = ~n7472 & ~n7546;
  assign n7548 = pi567 & ~n7547;
  assign n7549 = n7461 & ~n7548;
  assign n7550 = pi350 & ~pi592;
  assign n7551 = ~n7549 & ~n7550;
  assign n7552 = pi321 & ~pi347;
  assign n7553 = ~pi321 & pi347;
  assign n7554 = ~n7552 & ~n7553;
  assign n7555 = pi316 & ~pi349;
  assign n7556 = ~pi316 & pi349;
  assign n7557 = ~n7555 & ~n7556;
  assign n7558 = pi348 & n7557;
  assign n7559 = ~pi348 & ~n7557;
  assign n7560 = ~n7558 & ~n7559;
  assign n7561 = pi315 & ~pi359;
  assign n7562 = ~pi315 & pi359;
  assign n7563 = ~n7561 & ~n7562;
  assign n7564 = pi322 & n7563;
  assign n7565 = ~pi322 & ~n7563;
  assign n7566 = ~n7564 & ~n7565;
  assign n7567 = n7560 & ~n7566;
  assign n7568 = ~n7560 & n7566;
  assign n7569 = ~n7567 & ~n7568;
  assign n7570 = n7554 & n7569;
  assign n7571 = ~n7554 & ~n7569;
  assign n7572 = ~n7570 & ~n7571;
  assign n7573 = ~pi87 & ~n7532;
  assign n7574 = ~n7520 & n7573;
  assign n7575 = ~pi1091 & ~n7455;
  assign n7576 = pi1091 & ~n7540;
  assign n7577 = pi87 & ~pi100;
  assign n7578 = n3181 & n7577;
  assign n7579 = ~n7576 & n7578;
  assign n7580 = ~n7575 & n7579;
  assign n7581 = ~pi75 & ~n7580;
  assign n7582 = ~n7574 & n7581;
  assign n7583 = ~n7472 & ~n7582;
  assign n7584 = pi567 & ~n7583;
  assign n7585 = n7461 & ~n7584;
  assign n7586 = n7550 & ~n7585;
  assign n7587 = ~n7572 & ~n7586;
  assign n7588 = ~n7551 & n7587;
  assign n7589 = pi452 & ~pi455;
  assign n7590 = ~pi452 & pi455;
  assign n7591 = ~n7589 & ~n7590;
  assign n7592 = pi355 & n7591;
  assign n7593 = ~pi355 & ~n7591;
  assign n7594 = ~n7592 & ~n7593;
  assign n7595 = pi320 & ~pi460;
  assign n7596 = ~pi320 & pi460;
  assign n7597 = ~n7595 & ~n7596;
  assign n7598 = pi342 & ~n7597;
  assign n7599 = ~pi342 & n7597;
  assign n7600 = ~n7598 & ~n7599;
  assign n7601 = pi361 & ~pi441;
  assign n7602 = ~pi361 & pi441;
  assign n7603 = ~n7601 & ~n7602;
  assign n7604 = n7600 & n7603;
  assign n7605 = ~n7600 & ~n7603;
  assign n7606 = ~n7604 & ~n7605;
  assign n7607 = pi458 & n7606;
  assign n7608 = ~pi458 & ~n7606;
  assign n7609 = ~n7607 & ~n7608;
  assign n7610 = n7594 & n7609;
  assign n7611 = ~n7594 & ~n7609;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = pi1196 & n7612;
  assign n7614 = ~pi350 & ~pi592;
  assign n7615 = ~n7549 & ~n7614;
  assign n7616 = ~n7585 & n7614;
  assign n7617 = n7572 & ~n7616;
  assign n7618 = ~n7615 & n7617;
  assign n7619 = ~n7613 & ~n7618;
  assign n7620 = ~n7588 & n7619;
  assign n7621 = ~pi592 & ~n7585;
  assign n7622 = pi592 & ~n7549;
  assign n7623 = ~n7621 & ~n7622;
  assign n7624 = n7613 & ~n7623;
  assign n7625 = pi1198 & ~n7624;
  assign n7626 = ~n7620 & n7625;
  assign n7627 = ~pi455 & ~n7623;
  assign n7628 = pi455 & ~n7549;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = ~pi452 & ~n7629;
  assign n7631 = pi455 & ~n7623;
  assign n7632 = ~pi455 & ~n7549;
  assign n7633 = ~n7631 & ~n7632;
  assign n7634 = pi452 & ~n7633;
  assign n7635 = ~n7630 & ~n7634;
  assign n7636 = ~pi355 & ~n7635;
  assign n7637 = ~pi452 & ~n7633;
  assign n7638 = pi452 & ~n7629;
  assign n7639 = ~n7637 & ~n7638;
  assign n7640 = pi355 & ~n7639;
  assign n7641 = ~n7636 & ~n7640;
  assign n7642 = ~pi458 & ~n7641;
  assign n7643 = ~pi355 & ~n7639;
  assign n7644 = pi355 & ~n7635;
  assign n7645 = ~n7643 & ~n7644;
  assign n7646 = pi458 & ~n7645;
  assign n7647 = ~n7606 & ~n7646;
  assign n7648 = ~n7642 & n7647;
  assign n7649 = ~pi458 & ~n7645;
  assign n7650 = pi458 & ~n7641;
  assign n7651 = n7606 & ~n7650;
  assign n7652 = ~n7649 & n7651;
  assign n7653 = pi1196 & ~n7652;
  assign n7654 = ~n7648 & n7653;
  assign n7655 = ~pi1196 & ~n7549;
  assign n7656 = ~pi1198 & ~n7655;
  assign n7657 = ~n7654 & n7656;
  assign n7658 = ~n7626 & ~n7657;
  assign n7659 = ~n7421 & ~n7658;
  assign n7660 = n7421 & n7623;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = ~n7396 & n7661;
  assign n7663 = pi1199 & ~n7623;
  assign n7664 = pi351 & n7663;
  assign n7665 = ~n7662 & ~n7664;
  assign n7666 = ~pi461 & ~n7665;
  assign n7667 = ~pi351 & pi1199;
  assign n7668 = n7661 & ~n7667;
  assign n7669 = ~pi351 & n7663;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = pi461 & ~n7670;
  assign n7672 = ~n7666 & ~n7671;
  assign n7673 = ~pi357 & ~n7672;
  assign n7674 = ~pi461 & ~n7670;
  assign n7675 = pi461 & ~n7665;
  assign n7676 = ~n7674 & ~n7675;
  assign n7677 = pi357 & ~n7676;
  assign n7678 = ~n7673 & ~n7677;
  assign n7679 = ~pi356 & ~n7678;
  assign n7680 = ~pi357 & ~n7676;
  assign n7681 = pi357 & ~n7672;
  assign n7682 = ~n7680 & ~n7681;
  assign n7683 = pi356 & ~n7682;
  assign n7684 = ~n7679 & ~n7683;
  assign n7685 = n7395 & ~n7684;
  assign n7686 = ~pi356 & ~n7682;
  assign n7687 = pi356 & ~n7678;
  assign n7688 = ~n7686 & ~n7687;
  assign n7689 = ~n7395 & ~n7688;
  assign n7690 = ~pi591 & ~n7689;
  assign n7691 = ~n7685 & n7690;
  assign n7692 = pi591 & n7549;
  assign n7693 = pi590 & ~n7692;
  assign n7694 = ~n7691 & n7693;
  assign n7695 = ~pi285 & ~pi286;
  assign n7696 = ~pi289 & n7695;
  assign n7697 = ~pi288 & n7696;
  assign n7698 = ~pi363 & ~pi372;
  assign n7699 = pi363 & pi372;
  assign n7700 = ~n7698 & ~n7699;
  assign n7701 = pi386 & ~n7700;
  assign n7702 = ~pi386 & n7700;
  assign n7703 = ~n7701 & ~n7702;
  assign n7704 = pi338 & ~pi388;
  assign n7705 = ~pi338 & pi388;
  assign n7706 = ~n7704 & ~n7705;
  assign n7707 = pi337 & ~pi339;
  assign n7708 = ~pi337 & pi339;
  assign n7709 = ~n7707 & ~n7708;
  assign n7710 = pi387 & n7709;
  assign n7711 = ~pi387 & ~n7709;
  assign n7712 = ~n7710 & ~n7711;
  assign n7713 = pi380 & ~n7712;
  assign n7714 = ~pi380 & n7712;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = n7706 & ~n7715;
  assign n7717 = ~n7706 & n7715;
  assign n7718 = ~n7716 & ~n7717;
  assign n7719 = n7703 & n7718;
  assign n7720 = ~n7703 & ~n7718;
  assign n7721 = ~n7719 & ~n7720;
  assign n7722 = pi1196 & ~n7721;
  assign n7723 = ~pi368 & ~pi389;
  assign n7724 = pi368 & pi389;
  assign n7725 = ~n7723 & ~n7724;
  assign n7726 = pi365 & ~pi447;
  assign n7727 = ~pi365 & pi447;
  assign n7728 = ~n7726 & ~n7727;
  assign n7729 = pi336 & ~pi383;
  assign n7730 = ~pi336 & pi383;
  assign n7731 = ~n7729 & ~n7730;
  assign n7732 = pi364 & ~pi366;
  assign n7733 = ~pi364 & pi366;
  assign n7734 = ~n7732 & ~n7733;
  assign n7735 = n7731 & n7734;
  assign n7736 = ~n7731 & ~n7734;
  assign n7737 = ~n7735 & ~n7736;
  assign n7738 = n7728 & n7737;
  assign n7739 = ~n7728 & ~n7737;
  assign n7740 = ~n7738 & ~n7739;
  assign n7741 = n7725 & n7740;
  assign n7742 = ~n7725 & ~n7740;
  assign n7743 = ~n7741 & ~n7742;
  assign n7744 = pi367 & ~n7743;
  assign n7745 = ~pi367 & n7743;
  assign n7746 = ~n7744 & ~n7745;
  assign n7747 = pi1197 & n7746;
  assign n7748 = ~n7722 & ~n7747;
  assign n7749 = pi377 & pi592;
  assign n7750 = ~n7549 & ~n7749;
  assign n7751 = pi379 & ~pi382;
  assign n7752 = ~pi379 & pi382;
  assign n7753 = ~n7751 & ~n7752;
  assign n7754 = pi376 & ~pi439;
  assign n7755 = ~pi376 & pi439;
  assign n7756 = ~n7754 & ~n7755;
  assign n7757 = pi381 & n7756;
  assign n7758 = ~pi381 & ~n7756;
  assign n7759 = ~n7757 & ~n7758;
  assign n7760 = pi317 & ~pi385;
  assign n7761 = ~pi317 & pi385;
  assign n7762 = ~n7760 & ~n7761;
  assign n7763 = pi378 & n7762;
  assign n7764 = ~pi378 & ~n7762;
  assign n7765 = ~n7763 & ~n7764;
  assign n7766 = n7759 & ~n7765;
  assign n7767 = ~n7759 & n7765;
  assign n7768 = ~n7766 & ~n7767;
  assign n7769 = n7753 & n7768;
  assign n7770 = ~n7753 & ~n7768;
  assign n7771 = ~n7769 & ~n7770;
  assign n7772 = ~n7585 & n7749;
  assign n7773 = ~n7771 & ~n7772;
  assign n7774 = ~n7750 & n7773;
  assign n7775 = ~pi377 & pi592;
  assign n7776 = ~n7549 & ~n7775;
  assign n7777 = ~n7585 & n7775;
  assign n7778 = n7771 & ~n7777;
  assign n7779 = ~n7776 & n7778;
  assign n7780 = ~n7774 & ~n7779;
  assign n7781 = n7748 & ~n7780;
  assign n7782 = pi592 & ~n7585;
  assign n7783 = ~pi592 & ~n7549;
  assign n7784 = ~n7782 & ~n7783;
  assign n7785 = ~n7748 & n7784;
  assign n7786 = ~n7781 & ~n7785;
  assign n7787 = pi1199 & n7786;
  assign n7788 = ~pi1196 & ~n7747;
  assign n7789 = n7784 & ~n7788;
  assign n7790 = n7549 & ~n7747;
  assign n7791 = ~pi1196 & n7790;
  assign n7792 = ~n7789 & ~n7791;
  assign n7793 = ~n7721 & ~n7792;
  assign n7794 = n7747 & n7784;
  assign n7795 = ~n7790 & ~n7794;
  assign n7796 = n7721 & ~n7795;
  assign n7797 = ~pi1199 & ~n7796;
  assign n7798 = ~n7793 & n7797;
  assign n7799 = ~n7787 & ~n7798;
  assign n7800 = ~pi374 & ~n7799;
  assign n7801 = ~pi1198 & n7798;
  assign n7802 = ~pi1198 & pi1199;
  assign n7803 = n7786 & n7802;
  assign n7804 = pi1198 & ~n7784;
  assign n7805 = ~n7803 & ~n7804;
  assign n7806 = ~n7801 & n7805;
  assign n7807 = pi374 & ~n7806;
  assign n7808 = ~n7800 & ~n7807;
  assign n7809 = ~pi369 & ~n7808;
  assign n7810 = ~pi374 & ~n7806;
  assign n7811 = pi374 & ~n7799;
  assign n7812 = ~n7810 & ~n7811;
  assign n7813 = pi369 & ~n7812;
  assign n7814 = ~n7809 & ~n7813;
  assign n7815 = ~pi370 & ~n7814;
  assign n7816 = pi369 & ~n7808;
  assign n7817 = ~pi369 & ~n7812;
  assign n7818 = ~n7816 & ~n7817;
  assign n7819 = pi370 & ~n7818;
  assign n7820 = ~n7815 & ~n7819;
  assign n7821 = ~pi371 & ~n7820;
  assign n7822 = ~pi370 & ~n7818;
  assign n7823 = pi370 & ~n7814;
  assign n7824 = ~n7822 & ~n7823;
  assign n7825 = pi371 & ~n7824;
  assign n7826 = ~n7821 & ~n7825;
  assign n7827 = ~pi373 & ~n7826;
  assign n7828 = ~pi371 & ~n7824;
  assign n7829 = pi371 & ~n7820;
  assign n7830 = ~n7828 & ~n7829;
  assign n7831 = pi373 & ~n7830;
  assign n7832 = ~n7827 & ~n7831;
  assign n7833 = ~pi375 & n7832;
  assign n7834 = pi384 & ~pi442;
  assign n7835 = ~pi384 & pi442;
  assign n7836 = ~n7834 & ~n7835;
  assign n7837 = pi440 & ~n7836;
  assign n7838 = ~pi440 & n7836;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = ~pi373 & ~n7830;
  assign n7841 = pi373 & ~n7826;
  assign n7842 = ~n7840 & ~n7841;
  assign n7843 = pi375 & n7842;
  assign n7844 = ~n7839 & ~n7843;
  assign n7845 = ~n7833 & n7844;
  assign n7846 = pi375 & n7832;
  assign n7847 = ~pi375 & n7842;
  assign n7848 = n7839 & ~n7847;
  assign n7849 = ~n7846 & n7848;
  assign n7850 = ~pi591 & ~n7849;
  assign n7851 = ~n7845 & n7850;
  assign n7852 = pi1197 & ~n7623;
  assign n7853 = pi328 & ~pi408;
  assign n7854 = ~pi328 & pi408;
  assign n7855 = ~n7853 & ~n7854;
  assign n7856 = ~pi394 & ~pi396;
  assign n7857 = pi394 & pi396;
  assign n7858 = ~n7856 & ~n7857;
  assign n7859 = n7855 & ~n7858;
  assign n7860 = ~n7855 & n7858;
  assign n7861 = ~n7859 & ~n7860;
  assign n7862 = pi398 & ~pi399;
  assign n7863 = ~pi398 & pi399;
  assign n7864 = ~n7862 & ~n7863;
  assign n7865 = pi395 & n7864;
  assign n7866 = ~pi395 & ~n7864;
  assign n7867 = ~n7865 & ~n7866;
  assign n7868 = pi329 & ~n7867;
  assign n7869 = ~pi329 & n7867;
  assign n7870 = ~n7868 & ~n7869;
  assign n7871 = pi400 & ~n7870;
  assign n7872 = ~pi400 & n7870;
  assign n7873 = ~n7871 & ~n7872;
  assign n7874 = n7861 & n7873;
  assign n7875 = ~n7861 & ~n7873;
  assign n7876 = ~n7874 & ~n7875;
  assign n7877 = pi1198 & ~n7876;
  assign n7878 = n7623 & n7877;
  assign n7879 = pi390 & ~pi410;
  assign n7880 = ~pi390 & pi410;
  assign n7881 = ~n7879 & ~n7880;
  assign n7882 = pi397 & ~pi412;
  assign n7883 = ~pi397 & pi412;
  assign n7884 = ~n7882 & ~n7883;
  assign n7885 = pi404 & n7884;
  assign n7886 = ~pi404 & ~n7884;
  assign n7887 = ~n7885 & ~n7886;
  assign n7888 = pi319 & ~pi324;
  assign n7889 = ~pi319 & pi324;
  assign n7890 = ~n7888 & ~n7889;
  assign n7891 = pi456 & ~n7890;
  assign n7892 = ~pi456 & n7890;
  assign n7893 = ~n7891 & ~n7892;
  assign n7894 = n7887 & ~n7893;
  assign n7895 = ~n7887 & n7893;
  assign n7896 = ~n7894 & ~n7895;
  assign n7897 = n7881 & n7896;
  assign n7898 = ~n7881 & ~n7896;
  assign n7899 = ~n7897 & ~n7898;
  assign n7900 = pi411 & n7899;
  assign n7901 = ~pi411 & ~n7899;
  assign n7902 = ~n7900 & ~n7901;
  assign n7903 = n7523 & n7902;
  assign n7904 = n7520 & ~n7903;
  assign n7905 = n7573 & ~n7904;
  assign n7906 = ~n7541 & n7578;
  assign n7907 = n7535 & n7902;
  assign n7908 = n7536 & ~n7907;
  assign n7909 = n7906 & ~n7908;
  assign n7910 = ~pi75 & ~pi592;
  assign n7911 = pi1196 & n7910;
  assign n7912 = ~n7909 & n7911;
  assign n7913 = ~n7905 & n7912;
  assign n7914 = ~pi1196 & n7546;
  assign n7915 = ~n7913 & ~n7914;
  assign n7916 = ~pi1199 & ~n7915;
  assign n7917 = pi318 & ~pi409;
  assign n7918 = ~pi318 & pi409;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = pi401 & ~pi402;
  assign n7921 = ~pi401 & pi402;
  assign n7922 = ~n7920 & ~n7921;
  assign n7923 = pi406 & n7922;
  assign n7924 = ~pi406 & ~n7922;
  assign n7925 = ~n7923 & ~n7924;
  assign n7926 = ~pi403 & ~pi405;
  assign n7927 = pi403 & pi405;
  assign n7928 = ~n7926 & ~n7927;
  assign n7929 = pi325 & ~pi326;
  assign n7930 = ~pi325 & pi326;
  assign n7931 = ~n7929 & ~n7930;
  assign n7932 = n7928 & n7931;
  assign n7933 = ~n7928 & ~n7931;
  assign n7934 = ~n7932 & ~n7933;
  assign n7935 = n7925 & ~n7934;
  assign n7936 = ~n7925 & n7934;
  assign n7937 = ~n7935 & ~n7936;
  assign n7938 = n7919 & n7937;
  assign n7939 = ~n7919 & ~n7937;
  assign n7940 = ~n7938 & ~n7939;
  assign n7941 = pi1196 & ~n7902;
  assign n7942 = ~pi75 & n7941;
  assign n7943 = ~n7940 & ~n7942;
  assign n7944 = n7523 & n7943;
  assign n7945 = n7520 & ~n7944;
  assign n7946 = n7573 & ~n7945;
  assign n7947 = n7535 & ~n7940;
  assign n7948 = n7536 & ~n7947;
  assign n7949 = n7906 & ~n7948;
  assign n7950 = ~n7908 & n7949;
  assign n7951 = ~pi1196 & n7949;
  assign n7952 = pi1199 & n7910;
  assign n7953 = ~n7951 & n7952;
  assign n7954 = ~n7950 & n7953;
  assign n7955 = ~n7946 & n7954;
  assign n7956 = ~n7547 & ~n7910;
  assign n7957 = ~n7955 & ~n7956;
  assign n7958 = ~n7916 & n7957;
  assign n7959 = pi567 & ~n7958;
  assign n7960 = n7461 & ~n7877;
  assign n7961 = ~n7959 & n7960;
  assign n7962 = ~n7878 & ~n7961;
  assign n7963 = ~pi1197 & n7962;
  assign n7964 = ~n7852 & ~n7963;
  assign n7965 = pi333 & ~n7964;
  assign n7966 = ~pi333 & n7962;
  assign n7967 = ~n7965 & ~n7966;
  assign n7968 = pi391 & ~n7967;
  assign n7969 = pi333 & ~n7962;
  assign n7970 = ~pi333 & n7964;
  assign n7971 = ~n7969 & ~n7970;
  assign n7972 = ~pi391 & n7971;
  assign n7973 = ~n7968 & ~n7972;
  assign n7974 = ~pi392 & ~n7973;
  assign n7975 = ~pi391 & ~n7967;
  assign n7976 = pi391 & n7971;
  assign n7977 = ~n7975 & ~n7976;
  assign n7978 = pi392 & ~n7977;
  assign n7979 = ~n7974 & ~n7978;
  assign n7980 = ~pi393 & ~n7979;
  assign n7981 = ~pi392 & ~n7977;
  assign n7982 = pi392 & ~n7973;
  assign n7983 = ~n7981 & ~n7982;
  assign n7984 = pi393 & ~n7983;
  assign n7985 = ~n7980 & ~n7984;
  assign n7986 = pi334 & n7985;
  assign n7987 = pi407 & ~pi463;
  assign n7988 = ~pi407 & pi463;
  assign n7989 = ~n7987 & ~n7988;
  assign n7990 = pi335 & ~pi413;
  assign n7991 = ~pi335 & pi413;
  assign n7992 = ~n7990 & ~n7991;
  assign n7993 = n7989 & n7992;
  assign n7994 = ~n7989 & ~n7992;
  assign n7995 = ~n7993 & ~n7994;
  assign n7996 = ~pi393 & ~n7983;
  assign n7997 = pi393 & ~n7979;
  assign n7998 = ~n7996 & ~n7997;
  assign n7999 = ~pi334 & n7998;
  assign n8000 = ~n7995 & ~n7999;
  assign n8001 = ~n7986 & n8000;
  assign n8002 = pi334 & n7998;
  assign n8003 = ~pi334 & n7985;
  assign n8004 = n7995 & ~n8003;
  assign n8005 = ~n8002 & n8004;
  assign n8006 = pi591 & ~n8005;
  assign n8007 = ~n8001 & n8006;
  assign n8008 = ~pi590 & ~n8007;
  assign n8009 = ~n7851 & n8008;
  assign n8010 = n7697 & ~n8009;
  assign n8011 = ~n7694 & n8010;
  assign n8012 = n7465 & n7526;
  assign n8013 = pi1091 & ~n8012;
  assign n8014 = n7464 & ~n8013;
  assign n8015 = ~pi122 & pi1093;
  assign n8016 = ~pi98 & n7474;
  assign n8017 = n8015 & n8016;
  assign n8018 = ~pi1091 & ~n8017;
  assign n8019 = n8014 & ~n8018;
  assign n8020 = n7474 & n8015;
  assign n8021 = ~pi1091 & n8020;
  assign n8022 = ~pi98 & n8021;
  assign n8023 = ~n7464 & n8022;
  assign n8024 = pi75 & ~n8023;
  assign n8025 = ~n8019 & n8024;
  assign n8026 = ~pi39 & ~n7501;
  assign n8027 = ~pi122 & n8016;
  assign n8028 = pi122 & n7477;
  assign n8029 = ~n8027 & ~n8028;
  assign n8030 = pi1093 & ~n8029;
  assign n8031 = n7502 & ~n8030;
  assign n8032 = n8026 & ~n8031;
  assign n8033 = pi1091 & ~n7507;
  assign n8034 = ~n8018 & ~n8033;
  assign n8035 = ~n6192 & n8034;
  assign n8036 = n6192 & n8022;
  assign n8037 = ~n8035 & ~n8036;
  assign n8038 = ~n6189 & n8037;
  assign n8039 = ~pi216 & n6434;
  assign n8040 = n6198 & n8034;
  assign n8041 = ~n6198 & n8022;
  assign n8042 = ~n8040 & ~n8041;
  assign n8043 = n6189 & n8042;
  assign n8044 = n8039 & ~n8043;
  assign n8045 = ~n8038 & n8044;
  assign n8046 = n8022 & ~n8039;
  assign n8047 = pi299 & ~n8046;
  assign n8048 = ~n8045 & n8047;
  assign n8049 = ~n6215 & n8037;
  assign n8050 = ~pi223 & n5770;
  assign n8051 = n6215 & n8042;
  assign n8052 = n8050 & ~n8051;
  assign n8053 = ~n8049 & n8052;
  assign n8054 = n8022 & ~n8050;
  assign n8055 = ~pi299 & ~n8054;
  assign n8056 = ~n8053 & n8055;
  assign n8057 = pi39 & ~n8056;
  assign n8058 = ~n8048 & n8057;
  assign n8059 = ~n8032 & ~n8058;
  assign n8060 = ~pi38 & ~n8059;
  assign n8061 = pi38 & n8022;
  assign n8062 = ~pi100 & ~n8061;
  assign n8063 = ~n8060 & n8062;
  assign n8064 = pi228 & ~n7463;
  assign n8065 = pi1091 & ~n7527;
  assign n8066 = ~n8018 & ~n8065;
  assign n8067 = n8064 & ~n8066;
  assign n8068 = ~n8022 & ~n8064;
  assign n8069 = n3181 & ~n8068;
  assign n8070 = ~n8067 & n8069;
  assign n8071 = ~n3181 & n8022;
  assign n8072 = pi100 & ~n8071;
  assign n8073 = ~n8070 & n8072;
  assign n8074 = ~pi87 & ~n8073;
  assign n8075 = ~n8063 & n8074;
  assign n8076 = pi122 & n7535;
  assign n8077 = ~n8027 & ~n8076;
  assign n8078 = pi1093 & ~n8077;
  assign n8079 = n7575 & ~n8078;
  assign n8080 = n3207 & ~n7576;
  assign n8081 = ~n8079 & n8080;
  assign n8082 = ~n8022 & ~n8081;
  assign n8083 = pi87 & ~n8082;
  assign n8084 = ~pi75 & ~n8083;
  assign n8085 = ~n8075 & n8084;
  assign n8086 = ~n8025 & ~n8085;
  assign n8087 = pi567 & ~n8086;
  assign n8088 = n7461 & ~n8087;
  assign n8089 = pi567 & n8022;
  assign n8090 = ~n7422 & n8089;
  assign n8091 = ~n8088 & ~n8090;
  assign n8092 = pi592 & n8091;
  assign n8093 = ~n7621 & ~n8092;
  assign n8094 = n7421 & ~n8093;
  assign n8095 = pi455 & ~n8093;
  assign n8096 = ~pi455 & n8091;
  assign n8097 = ~n8095 & ~n8096;
  assign n8098 = pi452 & ~n8097;
  assign n8099 = pi355 & ~n7609;
  assign n8100 = ~pi355 & n7609;
  assign n8101 = ~n8099 & ~n8100;
  assign n8102 = ~pi455 & ~n8093;
  assign n8103 = pi455 & n8091;
  assign n8104 = ~n8102 & ~n8103;
  assign n8105 = ~pi452 & ~n8104;
  assign n8106 = n8101 & ~n8105;
  assign n8107 = ~n8098 & n8106;
  assign n8108 = pi452 & ~n8104;
  assign n8109 = ~pi452 & ~n8097;
  assign n8110 = ~n8101 & ~n8109;
  assign n8111 = ~n8108 & n8110;
  assign n8112 = pi1196 & ~n8111;
  assign n8113 = ~n8107 & n8112;
  assign n8114 = ~pi1196 & n8091;
  assign n8115 = ~pi1198 & ~n8114;
  assign n8116 = ~n8113 & n8115;
  assign n8117 = ~n7614 & n8091;
  assign n8118 = n7617 & ~n8117;
  assign n8119 = ~n7550 & n8091;
  assign n8120 = n7587 & ~n8119;
  assign n8121 = ~n7613 & ~n8120;
  assign n8122 = ~n8118 & n8121;
  assign n8123 = n7613 & ~n8093;
  assign n8124 = pi1198 & ~n8123;
  assign n8125 = ~n8122 & n8124;
  assign n8126 = ~n7421 & ~n8125;
  assign n8127 = ~n8116 & n8126;
  assign n8128 = ~n8094 & ~n8127;
  assign n8129 = ~n7396 & ~n8128;
  assign n8130 = pi1199 & ~n8093;
  assign n8131 = pi351 & n8130;
  assign n8132 = ~n8129 & ~n8131;
  assign n8133 = ~pi461 & ~n8132;
  assign n8134 = ~n7667 & ~n8128;
  assign n8135 = ~pi351 & n8130;
  assign n8136 = ~n8134 & ~n8135;
  assign n8137 = pi461 & ~n8136;
  assign n8138 = ~n8133 & ~n8137;
  assign n8139 = ~pi357 & ~n8138;
  assign n8140 = ~pi461 & ~n8136;
  assign n8141 = pi461 & ~n8132;
  assign n8142 = ~n8140 & ~n8141;
  assign n8143 = pi357 & ~n8142;
  assign n8144 = ~n8139 & ~n8143;
  assign n8145 = ~pi356 & ~n8144;
  assign n8146 = ~pi357 & ~n8142;
  assign n8147 = pi357 & ~n8138;
  assign n8148 = ~n8146 & ~n8147;
  assign n8149 = pi356 & ~n8148;
  assign n8150 = ~n8145 & ~n8149;
  assign n8151 = n7395 & ~n8150;
  assign n8152 = ~pi356 & ~n8148;
  assign n8153 = pi356 & ~n8144;
  assign n8154 = ~n8152 & ~n8153;
  assign n8155 = ~n7395 & ~n8154;
  assign n8156 = ~pi591 & ~n8155;
  assign n8157 = ~n8151 & n8156;
  assign n8158 = pi591 & ~n8091;
  assign n8159 = pi590 & ~n8158;
  assign n8160 = ~n8157 & n8159;
  assign n8161 = pi375 & n7839;
  assign n8162 = ~pi375 & ~n7839;
  assign n8163 = ~n8161 & ~n8162;
  assign n8164 = pi373 & ~n8163;
  assign n8165 = ~pi373 & n8163;
  assign n8166 = ~n8164 & ~n8165;
  assign n8167 = ~pi592 & n8091;
  assign n8168 = ~n7782 & ~n8167;
  assign n8169 = ~n7748 & n8168;
  assign n8170 = n7748 & ~n8091;
  assign n8171 = ~pi1199 & ~n8170;
  assign n8172 = ~n8169 & n8171;
  assign n8173 = ~n7775 & n8091;
  assign n8174 = n7778 & ~n8173;
  assign n8175 = ~n7749 & n8091;
  assign n8176 = n7773 & ~n8175;
  assign n8177 = ~n8174 & ~n8176;
  assign n8178 = n7748 & ~n8177;
  assign n8179 = pi1199 & ~n8169;
  assign n8180 = ~n8178 & n8179;
  assign n8181 = ~n8172 & ~n8180;
  assign n8182 = ~pi374 & ~n8181;
  assign n8183 = ~pi1198 & ~n8181;
  assign n8184 = pi1198 & ~n8168;
  assign n8185 = ~n8183 & ~n8184;
  assign n8186 = pi374 & ~n8185;
  assign n8187 = ~n8182 & ~n8186;
  assign n8188 = ~pi369 & ~n8187;
  assign n8189 = ~pi374 & ~n8185;
  assign n8190 = pi374 & ~n8181;
  assign n8191 = ~n8189 & ~n8190;
  assign n8192 = pi369 & ~n8191;
  assign n8193 = ~n8188 & ~n8192;
  assign n8194 = ~pi370 & ~n8193;
  assign n8195 = pi369 & ~n8187;
  assign n8196 = ~pi369 & ~n8191;
  assign n8197 = ~n8195 & ~n8196;
  assign n8198 = pi370 & ~n8197;
  assign n8199 = ~n8194 & ~n8198;
  assign n8200 = ~pi371 & ~n8199;
  assign n8201 = ~pi370 & ~n8197;
  assign n8202 = pi370 & ~n8193;
  assign n8203 = ~n8201 & ~n8202;
  assign n8204 = pi371 & ~n8203;
  assign n8205 = ~n8200 & ~n8204;
  assign n8206 = n8166 & ~n8205;
  assign n8207 = ~pi371 & ~n8203;
  assign n8208 = pi371 & ~n8199;
  assign n8209 = ~n8207 & ~n8208;
  assign n8210 = ~n8166 & ~n8209;
  assign n8211 = ~pi591 & ~n8210;
  assign n8212 = ~n8206 & n8211;
  assign n8213 = pi334 & ~n7995;
  assign n8214 = ~pi334 & n7995;
  assign n8215 = ~n8213 & ~n8214;
  assign n8216 = pi393 & n8215;
  assign n8217 = ~pi393 & ~n8215;
  assign n8218 = ~n8216 & ~n8217;
  assign n8219 = ~pi592 & pi1196;
  assign n8220 = n7902 & n8017;
  assign n8221 = ~pi1091 & n8220;
  assign n8222 = pi567 & n8221;
  assign n8223 = ~n7422 & n8222;
  assign n8224 = ~n7940 & n8016;
  assign n8225 = n8223 & n8224;
  assign n8226 = n8219 & ~n8225;
  assign n8227 = ~n8050 & n8221;
  assign n8228 = ~pi299 & ~n8227;
  assign n8229 = ~n7940 & n8017;
  assign n8230 = ~pi1091 & n8229;
  assign n8231 = ~n8050 & n8230;
  assign n8232 = ~pi299 & ~n8231;
  assign n8233 = ~n8228 & ~n8232;
  assign n8234 = ~n6192 & n7508;
  assign n8235 = ~n7940 & n8221;
  assign n8236 = ~n8234 & ~n8235;
  assign n8237 = ~n6215 & n8236;
  assign n8238 = n6198 & n7508;
  assign n8239 = ~n8235 & ~n8238;
  assign n8240 = n6215 & n8239;
  assign n8241 = n8050 & ~n8240;
  assign n8242 = ~n8237 & n8241;
  assign n8243 = ~n8233 & ~n8242;
  assign n8244 = ~n8039 & n8221;
  assign n8245 = pi299 & ~n8244;
  assign n8246 = ~n8039 & n8230;
  assign n8247 = pi299 & ~n8246;
  assign n8248 = ~n8245 & ~n8247;
  assign n8249 = ~n6189 & n8236;
  assign n8250 = n6189 & n8239;
  assign n8251 = n8039 & ~n8250;
  assign n8252 = ~n8249 & n8251;
  assign n8253 = ~n8248 & ~n8252;
  assign n8254 = pi39 & ~n8253;
  assign n8255 = ~n8243 & n8254;
  assign n8256 = n7502 & ~n7902;
  assign n8257 = n8032 & ~n8256;
  assign n8258 = ~n7940 & n8030;
  assign n8259 = n7502 & ~n8258;
  assign n8260 = n8257 & ~n8259;
  assign n8261 = ~n8255 & ~n8260;
  assign n8262 = ~pi38 & ~n8261;
  assign n8263 = pi38 & n8221;
  assign n8264 = ~pi100 & ~n8263;
  assign n8265 = pi38 & n8230;
  assign n8266 = ~pi100 & ~n8265;
  assign n8267 = ~n8264 & ~n8266;
  assign n8268 = ~n8262 & ~n8267;
  assign n8269 = n6237 & n7528;
  assign n8270 = n6162 & ~n6238;
  assign n8271 = ~n6237 & ~n8270;
  assign n8272 = ~pi1091 & ~n8235;
  assign n8273 = n8271 & ~n8272;
  assign n8274 = ~n8065 & n8273;
  assign n8275 = ~n8269 & ~n8274;
  assign n8276 = pi228 & ~n8275;
  assign n8277 = pi228 & n8271;
  assign n8278 = n8235 & ~n8277;
  assign n8279 = pi232 & ~n8278;
  assign n8280 = ~n8276 & n8279;
  assign n8281 = ~pi232 & ~n8235;
  assign n8282 = ~n7529 & n8281;
  assign n8283 = n3181 & ~n8282;
  assign n8284 = ~n8280 & n8283;
  assign n8285 = ~n3181 & n8235;
  assign n8286 = pi100 & ~n8285;
  assign n8287 = ~n8284 & n8286;
  assign n8288 = ~n8268 & ~n8287;
  assign n8289 = ~pi87 & ~n8288;
  assign n8290 = ~n3207 & n8221;
  assign n8291 = pi87 & ~n8290;
  assign n8292 = ~n3207 & n8230;
  assign n8293 = pi87 & ~n8292;
  assign n8294 = ~n8291 & ~n8293;
  assign n8295 = n7575 & ~n7902;
  assign n8296 = n7575 & n7940;
  assign n8297 = n8081 & ~n8296;
  assign n8298 = ~n8295 & n8297;
  assign n8299 = ~n8294 & ~n8298;
  assign n8300 = ~n8289 & ~n8299;
  assign n8301 = ~pi75 & ~n8300;
  assign n8302 = ~n7464 & n8221;
  assign n8303 = pi75 & ~n8302;
  assign n8304 = ~n7464 & n8230;
  assign n8305 = pi75 & ~n8304;
  assign n8306 = ~n8303 & ~n8305;
  assign n8307 = n8014 & ~n8272;
  assign n8308 = ~n8306 & ~n8307;
  assign n8309 = ~n8301 & ~n8308;
  assign n8310 = n8226 & ~n8309;
  assign n8311 = pi567 & n8230;
  assign n8312 = ~n7422 & n8311;
  assign n8313 = ~pi592 & ~pi1196;
  assign n8314 = ~n8312 & n8313;
  assign n8315 = n8293 & ~n8297;
  assign n8316 = n7532 & ~n8230;
  assign n8317 = n8026 & ~n8259;
  assign n8318 = ~n8230 & ~n8238;
  assign n8319 = n6215 & n8318;
  assign n8320 = ~n8230 & ~n8234;
  assign n8321 = ~n6215 & n8320;
  assign n8322 = n8050 & ~n8321;
  assign n8323 = ~n8319 & n8322;
  assign n8324 = n8232 & ~n8323;
  assign n8325 = n6189 & n8318;
  assign n8326 = ~n6189 & n8320;
  assign n8327 = n8039 & ~n8326;
  assign n8328 = ~n8325 & n8327;
  assign n8329 = n8247 & ~n8328;
  assign n8330 = pi39 & ~n8329;
  assign n8331 = ~n8324 & n8330;
  assign n8332 = ~n8317 & ~n8331;
  assign n8333 = ~pi38 & ~n8332;
  assign n8334 = n8266 & ~n8333;
  assign n8335 = ~n8316 & ~n8334;
  assign n8336 = ~pi87 & ~n8335;
  assign n8337 = ~n8315 & ~n8336;
  assign n8338 = ~pi75 & ~n8337;
  assign n8339 = ~pi1091 & ~n8229;
  assign n8340 = n8014 & ~n8339;
  assign n8341 = n8305 & ~n8340;
  assign n8342 = ~n8338 & ~n8341;
  assign n8343 = n8314 & ~n8342;
  assign n8344 = ~n8310 & ~n8343;
  assign n8345 = pi567 & ~n8344;
  assign n8346 = ~n8226 & ~n8314;
  assign n8347 = ~n7461 & ~n8346;
  assign n8348 = pi1199 & ~n8347;
  assign n8349 = ~n8345 & n8348;
  assign n8350 = ~n8221 & ~n8238;
  assign n8351 = n6215 & n8350;
  assign n8352 = ~n8221 & ~n8234;
  assign n8353 = ~n6215 & n8352;
  assign n8354 = n8050 & ~n8353;
  assign n8355 = ~n8351 & n8354;
  assign n8356 = n8228 & ~n8355;
  assign n8357 = n6189 & n8350;
  assign n8358 = ~n6189 & n8352;
  assign n8359 = n8039 & ~n8358;
  assign n8360 = ~n8357 & n8359;
  assign n8361 = n8245 & ~n8360;
  assign n8362 = pi39 & ~n8361;
  assign n8363 = ~n8356 & n8362;
  assign n8364 = ~n8257 & ~n8363;
  assign n8365 = ~pi38 & ~n8364;
  assign n8366 = n8264 & ~n8365;
  assign n8367 = n7532 & ~n8221;
  assign n8368 = ~n8366 & ~n8367;
  assign n8369 = ~pi87 & ~n8368;
  assign n8370 = n8081 & ~n8295;
  assign n8371 = n8291 & ~n8370;
  assign n8372 = ~n8369 & ~n8371;
  assign n8373 = ~pi75 & ~n8372;
  assign n8374 = ~pi1091 & ~n8220;
  assign n8375 = n8014 & ~n8374;
  assign n8376 = n8303 & ~n8375;
  assign n8377 = ~n8373 & ~n8376;
  assign n8378 = pi567 & ~n8377;
  assign n8379 = n7461 & ~n8378;
  assign n8380 = n8219 & ~n8223;
  assign n8381 = ~n8379 & n8380;
  assign n8382 = ~pi1199 & ~n8114;
  assign n8383 = ~n8381 & n8382;
  assign n8384 = ~n7877 & ~n8383;
  assign n8385 = ~n8349 & n8384;
  assign n8386 = n7621 & n7877;
  assign n8387 = ~n8092 & ~n8386;
  assign n8388 = ~n8385 & n8387;
  assign n8389 = ~pi333 & ~n8388;
  assign n8390 = ~pi1197 & ~n8388;
  assign n8391 = pi1197 & ~n8093;
  assign n8392 = ~n8390 & ~n8391;
  assign n8393 = pi333 & ~n8392;
  assign n8394 = ~n8389 & ~n8393;
  assign n8395 = ~pi391 & ~n8394;
  assign n8396 = ~pi333 & ~n8392;
  assign n8397 = pi333 & ~n8388;
  assign n8398 = ~n8396 & ~n8397;
  assign n8399 = pi391 & ~n8398;
  assign n8400 = ~n8395 & ~n8399;
  assign n8401 = ~pi392 & ~n8400;
  assign n8402 = ~pi391 & ~n8398;
  assign n8403 = pi391 & ~n8394;
  assign n8404 = ~n8402 & ~n8403;
  assign n8405 = pi392 & ~n8404;
  assign n8406 = ~n8401 & ~n8405;
  assign n8407 = n8218 & ~n8406;
  assign n8408 = ~pi392 & ~n8404;
  assign n8409 = pi392 & ~n8400;
  assign n8410 = ~n8408 & ~n8409;
  assign n8411 = ~n8218 & ~n8410;
  assign n8412 = pi591 & ~n8411;
  assign n8413 = ~n8407 & n8412;
  assign n8414 = ~pi590 & ~n8413;
  assign n8415 = ~n8212 & n8414;
  assign n8416 = ~n7697 & ~n8415;
  assign n8417 = ~n8160 & n8416;
  assign n8418 = ~pi588 & ~n8417;
  assign n8419 = ~n8011 & n8418;
  assign po1038 = pi57 | ~n6286;
  assign n8421 = pi433 & ~pi451;
  assign n8422 = ~pi433 & pi451;
  assign n8423 = ~n8421 & ~n8422;
  assign n8424 = pi449 & n8423;
  assign n8425 = ~pi449 & ~n8423;
  assign n8426 = ~n8424 & ~n8425;
  assign n8427 = pi448 & ~n8426;
  assign n8428 = ~pi448 & n8426;
  assign n8429 = ~n8427 & ~n8428;
  assign n8430 = ~pi417 & ~pi418;
  assign n8431 = pi417 & pi418;
  assign n8432 = ~n8430 & ~n8431;
  assign n8433 = pi437 & n8432;
  assign n8434 = ~pi437 & ~n8432;
  assign n8435 = ~n8433 & ~n8434;
  assign n8436 = pi453 & ~pi464;
  assign n8437 = ~pi453 & pi464;
  assign n8438 = ~n8436 & ~n8437;
  assign n8439 = n8435 & n8438;
  assign n8440 = ~n8435 & ~n8438;
  assign n8441 = ~n8439 & ~n8440;
  assign n8442 = pi415 & ~pi431;
  assign n8443 = ~pi415 & pi431;
  assign n8444 = ~n8442 & ~n8443;
  assign n8445 = pi416 & ~pi438;
  assign n8446 = ~pi416 & pi438;
  assign n8447 = ~n8445 & ~n8446;
  assign n8448 = n8444 & n8447;
  assign n8449 = ~n8444 & ~n8447;
  assign n8450 = ~n8448 & ~n8449;
  assign n8451 = ~n8441 & n8450;
  assign n8452 = n8441 & ~n8450;
  assign n8453 = pi1197 & ~n8452;
  assign n8454 = ~n8451 & n8453;
  assign n8455 = pi421 & ~pi454;
  assign n8456 = ~pi421 & pi454;
  assign n8457 = ~n8455 & ~n8456;
  assign n8458 = pi432 & ~pi459;
  assign n8459 = ~pi432 & pi459;
  assign n8460 = ~n8458 & ~n8459;
  assign n8461 = n8457 & ~n8460;
  assign n8462 = ~n8457 & n8460;
  assign n8463 = ~n8461 & ~n8462;
  assign n8464 = ~pi419 & ~pi420;
  assign n8465 = pi419 & pi420;
  assign n8466 = ~n8464 & ~n8465;
  assign n8467 = pi423 & ~pi424;
  assign n8468 = ~pi423 & pi424;
  assign n8469 = ~n8467 & ~n8468;
  assign n8470 = n8466 & ~n8469;
  assign n8471 = ~n8466 & n8469;
  assign n8472 = ~n8470 & ~n8471;
  assign n8473 = n8463 & n8472;
  assign n8474 = ~n8463 & ~n8472;
  assign n8475 = ~n8473 & ~n8474;
  assign n8476 = ~pi425 & n8475;
  assign n8477 = pi425 & ~n8475;
  assign n8478 = pi1198 & ~n8477;
  assign n8479 = ~n8476 & n8478;
  assign n8480 = ~n8454 & ~n8479;
  assign n8481 = n7623 & ~n8480;
  assign n8482 = ~pi443 & ~pi592;
  assign n8483 = ~n7549 & ~n8482;
  assign n8484 = ~n7585 & n8482;
  assign n8485 = ~n8483 & ~n8484;
  assign n8486 = ~pi444 & ~n8485;
  assign n8487 = pi443 & ~pi592;
  assign n8488 = ~n7549 & ~n8487;
  assign n8489 = ~n7585 & n8487;
  assign n8490 = ~n8488 & ~n8489;
  assign n8491 = pi444 & ~n8490;
  assign n8492 = ~n8486 & ~n8491;
  assign n8493 = pi436 & ~n8492;
  assign n8494 = ~pi429 & ~pi435;
  assign n8495 = pi429 & pi435;
  assign n8496 = ~n8494 & ~n8495;
  assign n8497 = pi434 & ~pi446;
  assign n8498 = ~pi434 & pi446;
  assign n8499 = ~n8497 & ~n8498;
  assign n8500 = pi414 & ~pi422;
  assign n8501 = ~pi414 & pi422;
  assign n8502 = ~n8500 & ~n8501;
  assign n8503 = n8499 & n8502;
  assign n8504 = ~n8499 & ~n8502;
  assign n8505 = ~n8503 & ~n8504;
  assign n8506 = n8496 & n8505;
  assign n8507 = ~n8496 & ~n8505;
  assign n8508 = ~n8506 & ~n8507;
  assign n8509 = ~pi444 & ~n8490;
  assign n8510 = pi444 & ~n8485;
  assign n8511 = ~n8509 & ~n8510;
  assign n8512 = ~pi436 & ~n8511;
  assign n8513 = ~n8508 & ~n8512;
  assign n8514 = ~n8493 & n8513;
  assign n8515 = pi436 & ~n8511;
  assign n8516 = ~pi436 & ~n8492;
  assign n8517 = n8508 & ~n8516;
  assign n8518 = ~n8515 & n8517;
  assign n8519 = pi1196 & ~n8518;
  assign n8520 = ~n8514 & n8519;
  assign n8521 = ~n7655 & n8480;
  assign n8522 = ~n8520 & n8521;
  assign n8523 = ~n8481 & ~n8522;
  assign n8524 = ~pi428 & ~n8523;
  assign n8525 = pi428 & n7623;
  assign n8526 = ~n8524 & ~n8525;
  assign n8527 = ~pi427 & ~n8526;
  assign n8528 = pi428 & ~n8523;
  assign n8529 = ~pi428 & n7623;
  assign n8530 = ~n8528 & ~n8529;
  assign n8531 = pi427 & ~n8530;
  assign n8532 = ~n8527 & ~n8531;
  assign n8533 = pi430 & ~n8532;
  assign n8534 = ~pi427 & ~n8530;
  assign n8535 = pi427 & ~n8526;
  assign n8536 = ~n8534 & ~n8535;
  assign n8537 = ~pi430 & ~n8536;
  assign n8538 = ~n8533 & ~n8537;
  assign n8539 = pi426 & ~n8538;
  assign n8540 = pi430 & ~n8536;
  assign n8541 = ~pi430 & ~n8532;
  assign n8542 = ~n8540 & ~n8541;
  assign n8543 = ~pi426 & ~n8542;
  assign n8544 = ~n8539 & ~n8543;
  assign n8545 = pi445 & ~n8544;
  assign n8546 = pi426 & ~n8542;
  assign n8547 = ~pi426 & ~n8538;
  assign n8548 = ~n8546 & ~n8547;
  assign n8549 = ~pi445 & ~n8548;
  assign n8550 = ~n8545 & ~n8549;
  assign n8551 = n8429 & ~n8550;
  assign n8552 = pi445 & ~n8548;
  assign n8553 = ~pi445 & ~n8544;
  assign n8554 = ~n8552 & ~n8553;
  assign n8555 = ~n8429 & ~n8554;
  assign n8556 = pi1199 & ~n8555;
  assign n8557 = ~n8551 & n8556;
  assign n8558 = ~pi590 & ~pi591;
  assign n8559 = ~pi1199 & n8523;
  assign n8560 = n8558 & ~n8559;
  assign n8561 = ~n8557 & n8560;
  assign n8562 = n7549 & ~n8558;
  assign n8563 = n7697 & ~n8562;
  assign n8564 = ~n8561 & n8563;
  assign n8565 = n8091 & ~n8487;
  assign n8566 = ~pi436 & pi444;
  assign n8567 = pi436 & ~pi444;
  assign n8568 = ~n8566 & ~n8567;
  assign n8569 = n8508 & ~n8568;
  assign n8570 = ~n8508 & n8568;
  assign n8571 = ~n8569 & ~n8570;
  assign n8572 = ~n8489 & ~n8571;
  assign n8573 = ~n8565 & n8572;
  assign n8574 = n8091 & ~n8482;
  assign n8575 = ~n8484 & n8571;
  assign n8576 = ~n8574 & n8575;
  assign n8577 = pi1196 & ~n8576;
  assign n8578 = ~n8573 & n8577;
  assign n8579 = ~n8114 & ~n8578;
  assign n8580 = n8480 & ~n8579;
  assign n8581 = ~n8093 & ~n8480;
  assign n8582 = ~n8580 & ~n8581;
  assign n8583 = pi428 & n8582;
  assign n8584 = ~pi428 & n8093;
  assign n8585 = pi427 & ~n8584;
  assign n8586 = ~n8583 & n8585;
  assign n8587 = ~pi428 & n8582;
  assign n8588 = pi428 & n8093;
  assign n8589 = ~pi427 & ~n8588;
  assign n8590 = ~n8587 & n8589;
  assign n8591 = ~n8586 & ~n8590;
  assign n8592 = pi430 & ~n8591;
  assign n8593 = ~pi427 & pi428;
  assign n8594 = pi427 & ~pi428;
  assign n8595 = ~n8593 & ~n8594;
  assign n8596 = n8093 & n8595;
  assign n8597 = n8582 & ~n8595;
  assign n8598 = ~n8596 & ~n8597;
  assign n8599 = ~pi430 & n8598;
  assign n8600 = ~n8592 & ~n8599;
  assign n8601 = ~pi426 & ~n8600;
  assign n8602 = ~pi430 & ~n8591;
  assign n8603 = pi430 & n8598;
  assign n8604 = ~n8602 & ~n8603;
  assign n8605 = pi426 & ~n8604;
  assign n8606 = ~n8601 & ~n8605;
  assign n8607 = ~pi445 & ~n8606;
  assign n8608 = ~pi426 & ~n8604;
  assign n8609 = pi426 & ~n8600;
  assign n8610 = ~n8608 & ~n8609;
  assign n8611 = pi445 & ~n8610;
  assign n8612 = ~n8607 & ~n8611;
  assign n8613 = ~pi448 & n8612;
  assign n8614 = ~pi445 & ~n8610;
  assign n8615 = pi445 & ~n8606;
  assign n8616 = ~n8614 & ~n8615;
  assign n8617 = pi448 & n8616;
  assign n8618 = ~n8426 & ~n8617;
  assign n8619 = ~n8613 & n8618;
  assign n8620 = pi448 & n8612;
  assign n8621 = ~pi448 & n8616;
  assign n8622 = n8426 & ~n8621;
  assign n8623 = ~n8620 & n8622;
  assign n8624 = ~n8619 & ~n8623;
  assign n8625 = pi1199 & ~n8624;
  assign n8626 = ~pi1199 & ~n8582;
  assign n8627 = n8558 & ~n8626;
  assign n8628 = ~n8625 & n8627;
  assign n8629 = ~n8091 & ~n8558;
  assign n8630 = ~n7697 & ~n8629;
  assign n8631 = ~n8628 & n8630;
  assign n8632 = ~n8564 & ~n8631;
  assign n8633 = pi588 & ~n8632;
  assign n8634 = ~po1038 & ~n8633;
  assign n8635 = ~n8419 & n8634;
  assign n8636 = ~pi592 & n7612;
  assign n8637 = ~n7600 & n8089;
  assign n8638 = ~n8636 & n8637;
  assign n8639 = pi361 & ~pi458;
  assign n8640 = ~pi361 & pi458;
  assign n8641 = ~n8639 & ~n8640;
  assign n8642 = n7594 & n8641;
  assign n8643 = ~n7594 & ~n8641;
  assign n8644 = ~n8642 & ~n8643;
  assign n8645 = pi441 & ~n8644;
  assign n8646 = ~pi441 & n8644;
  assign n8647 = ~pi592 & ~n8646;
  assign n8648 = ~n8645 & n8647;
  assign n8649 = n7600 & n8089;
  assign n8650 = ~n8648 & n8649;
  assign n8651 = pi1196 & ~n8650;
  assign n8652 = ~n8638 & n8651;
  assign n8653 = ~pi1198 & ~n8652;
  assign n8654 = pi350 & ~n7572;
  assign n8655 = ~pi350 & n7572;
  assign n8656 = ~n8654 & ~n8655;
  assign n8657 = ~n7613 & n8656;
  assign n8658 = ~pi592 & n8089;
  assign n8659 = pi1198 & n8658;
  assign n8660 = n8657 & n8659;
  assign n8661 = ~n8653 & ~n8660;
  assign n8662 = ~n7421 & ~n8661;
  assign n8663 = ~pi592 & ~n8662;
  assign n8664 = n8089 & ~n8663;
  assign n8665 = ~n7667 & ~n8664;
  assign n8666 = pi592 & n8089;
  assign n8667 = pi1199 & ~n8666;
  assign n8668 = ~pi351 & n8667;
  assign n8669 = ~n8665 & ~n8668;
  assign n8670 = ~pi461 & ~n8669;
  assign n8671 = ~n7396 & ~n8664;
  assign n8672 = pi351 & n8667;
  assign n8673 = ~n8671 & ~n8672;
  assign n8674 = pi461 & ~n8673;
  assign n8675 = ~n8670 & ~n8674;
  assign n8676 = ~pi357 & ~n8675;
  assign n8677 = ~pi461 & ~n8673;
  assign n8678 = pi461 & ~n8669;
  assign n8679 = ~n8677 & ~n8678;
  assign n8680 = pi357 & ~n8679;
  assign n8681 = ~n8676 & ~n8680;
  assign n8682 = pi356 & ~n8681;
  assign n8683 = ~pi357 & ~n8679;
  assign n8684 = pi357 & ~n8675;
  assign n8685 = ~n8683 & ~n8684;
  assign n8686 = ~pi356 & ~n8685;
  assign n8687 = n7395 & ~n8686;
  assign n8688 = ~n8682 & n8687;
  assign n8689 = pi356 & ~n8685;
  assign n8690 = ~pi356 & ~n8681;
  assign n8691 = ~n7395 & ~n8690;
  assign n8692 = ~n8689 & n8691;
  assign n8693 = ~n8688 & ~n8692;
  assign n8694 = pi590 & ~n8693;
  assign n8695 = pi592 & ~n7748;
  assign n8696 = ~pi377 & ~n7771;
  assign n8697 = pi377 & n7771;
  assign n8698 = ~n8696 & ~n8697;
  assign n8699 = n7748 & ~n8698;
  assign n8700 = pi592 & ~n8699;
  assign n8701 = n8089 & ~n8700;
  assign n8702 = pi1199 & ~n8701;
  assign n8703 = ~n8695 & ~n8702;
  assign n8704 = n8666 & n8703;
  assign n8705 = ~pi369 & ~pi374;
  assign n8706 = pi369 & pi374;
  assign n8707 = ~n8705 & ~n8706;
  assign n8708 = ~pi370 & ~n8707;
  assign n8709 = pi370 & n8707;
  assign n8710 = ~n8708 & ~n8709;
  assign n8711 = ~pi371 & ~n8710;
  assign n8712 = pi371 & n8710;
  assign n8713 = ~n8711 & ~n8712;
  assign n8714 = ~pi373 & ~n8713;
  assign n8715 = pi373 & n8713;
  assign n8716 = ~n8714 & ~n8715;
  assign n8717 = pi375 & ~n8716;
  assign n8718 = ~pi375 & n8716;
  assign n8719 = ~n8717 & ~n8718;
  assign n8720 = ~n7839 & ~n8719;
  assign n8721 = n7839 & n8719;
  assign n8722 = ~n8720 & ~n8721;
  assign n8723 = n8704 & n8722;
  assign n8724 = ~pi1198 & n8704;
  assign n8725 = ~n8658 & ~n8724;
  assign n8726 = ~n8723 & n8725;
  assign n8727 = ~pi590 & ~n8726;
  assign n8728 = ~pi591 & ~n8727;
  assign n8729 = ~n8694 & n8728;
  assign n8730 = pi1197 & ~n8666;
  assign n8731 = ~pi592 & n8311;
  assign n8732 = ~n7941 & n8731;
  assign n8733 = n8667 & ~n8732;
  assign n8734 = n8219 & n8222;
  assign n8735 = n8089 & ~n8219;
  assign n8736 = ~pi1199 & ~n8735;
  assign n8737 = ~n8734 & n8736;
  assign n8738 = ~n8733 & ~n8737;
  assign n8739 = ~pi1197 & ~n8738;
  assign n8740 = ~n8730 & ~n8739;
  assign n8741 = ~pi333 & ~n8740;
  assign n8742 = pi1198 & ~n8666;
  assign n8743 = n8738 & ~n8742;
  assign n8744 = ~n7876 & ~n8743;
  assign n8745 = n8738 & ~n8744;
  assign n8746 = ~n8741 & n8745;
  assign n8747 = ~pi391 & ~n8746;
  assign n8748 = pi333 & ~n8740;
  assign n8749 = ~pi333 & ~n8738;
  assign n8750 = ~n8744 & ~n8749;
  assign n8751 = ~n8748 & n8750;
  assign n8752 = pi391 & ~n8751;
  assign n8753 = ~n8747 & ~n8752;
  assign n8754 = ~pi392 & ~n8753;
  assign n8755 = ~pi391 & ~n8751;
  assign n8756 = pi391 & ~n8746;
  assign n8757 = ~n8755 & ~n8756;
  assign n8758 = pi392 & ~n8757;
  assign n8759 = ~n8754 & ~n8758;
  assign n8760 = pi393 & ~n8759;
  assign n8761 = ~pi392 & ~n8757;
  assign n8762 = pi392 & ~n8753;
  assign n8763 = ~n8761 & ~n8762;
  assign n8764 = ~pi393 & ~n8763;
  assign n8765 = n8215 & ~n8764;
  assign n8766 = ~n8760 & n8765;
  assign n8767 = pi393 & ~n8763;
  assign n8768 = ~pi393 & ~n8759;
  assign n8769 = ~n8215 & ~n8768;
  assign n8770 = ~n8767 & n8769;
  assign n8771 = ~n8766 & ~n8770;
  assign n8772 = ~pi590 & ~n8771;
  assign n8773 = pi590 & n8089;
  assign n8774 = pi591 & ~n8773;
  assign n8775 = ~n8772 & n8774;
  assign n8776 = ~n8729 & ~n8775;
  assign n8777 = ~pi588 & ~n8776;
  assign n8778 = ~n7697 & po1038;
  assign n8779 = pi436 & ~pi443;
  assign n8780 = ~pi436 & pi443;
  assign n8781 = ~n8779 & ~n8780;
  assign n8782 = ~pi444 & n8781;
  assign n8783 = pi444 & ~n8781;
  assign n8784 = ~n8782 & ~n8783;
  assign n8785 = n8508 & n8784;
  assign n8786 = ~n8508 & ~n8784;
  assign n8787 = n8219 & ~n8786;
  assign n8788 = ~n8785 & n8787;
  assign n8789 = n8480 & ~n8788;
  assign n8790 = n8658 & n8789;
  assign n8791 = pi430 & ~n8595;
  assign n8792 = ~pi430 & n8595;
  assign n8793 = ~n8791 & ~n8792;
  assign n8794 = ~pi426 & ~n8793;
  assign n8795 = pi426 & n8793;
  assign n8796 = ~n8794 & ~n8795;
  assign n8797 = ~pi445 & ~n8796;
  assign n8798 = pi445 & n8796;
  assign n8799 = ~n8797 & ~n8798;
  assign n8800 = ~pi448 & ~n8799;
  assign n8801 = pi448 & n8799;
  assign n8802 = ~n8800 & ~n8801;
  assign n8803 = n8790 & n8802;
  assign n8804 = ~n8666 & ~n8803;
  assign n8805 = ~n8426 & ~n8804;
  assign n8806 = n8790 & ~n8802;
  assign n8807 = ~n8666 & ~n8806;
  assign n8808 = n8426 & ~n8807;
  assign n8809 = pi1199 & ~n8808;
  assign n8810 = ~n8805 & n8809;
  assign n8811 = ~pi1199 & ~n8666;
  assign n8812 = ~n8790 & n8811;
  assign n8813 = n8558 & ~n8812;
  assign n8814 = ~n8810 & n8813;
  assign n8815 = n8089 & ~n8558;
  assign n8816 = pi588 & ~n8815;
  assign n8817 = ~n8814 & n8816;
  assign n8818 = n8778 & ~n8817;
  assign n8819 = ~n8777 & n8818;
  assign n8820 = ~pi217 & ~n8819;
  assign n8821 = ~n8635 & n8820;
  assign n8822 = ~n7549 & n7697;
  assign n8823 = ~n7697 & n8091;
  assign n8824 = ~po1038 & ~n8823;
  assign n8825 = ~n8822 & n8824;
  assign n8826 = n8089 & n8778;
  assign n8827 = pi217 & ~n8826;
  assign n8828 = ~n8825 & n8827;
  assign n8829 = ~pi1161 & ~pi1162;
  assign n8830 = ~pi1163 & n8829;
  assign n8831 = ~n8828 & n8830;
  assign n8832 = ~n8821 & n8831;
  assign n8833 = pi1161 & ~pi1163;
  assign n8834 = n2754 & n8833;
  assign n8835 = ~pi31 & pi1162;
  assign n8836 = n8834 & n8835;
  assign po189 = n8832 | n8836;
  assign n8838 = n3293 & n3429;
  assign n8839 = ~pi55 & ~pi74;
  assign n8840 = n8838 & n8839;
  assign n8841 = n6271 & n8840;
  assign n8842 = pi100 & n3181;
  assign n8843 = n6243 & ~po1057;
  assign n8844 = n6484 & n8843;
  assign n8845 = ~pi137 & n8844;
  assign n8846 = pi129 & n3095;
  assign n8847 = ~pi137 & pi252;
  assign n8848 = po1057 & ~n7463;
  assign n8849 = ~n6243 & ~n8848;
  assign n8850 = n8847 & n8849;
  assign n8851 = n8846 & n8850;
  assign n8852 = ~n8845 & ~n8851;
  assign n8853 = n8842 & ~n8852;
  assign n8854 = ~pi24 & ~pi90;
  assign n8855 = n6145 & n8854;
  assign n8856 = pi50 & n2586;
  assign n8857 = n2484 & n8856;
  assign n8858 = n2482 & n2510;
  assign n8859 = n2490 & n8858;
  assign n8860 = ~pi93 & n8859;
  assign n8861 = n8857 & n8860;
  assign n8862 = n8855 & n8861;
  assign n8863 = pi829 & ~pi1093;
  assign n8864 = n6257 & n8863;
  assign po840 = n2795 | n8864;
  assign n8866 = ~n7697 & ~po840;
  assign n8867 = ~pi137 & ~n8866;
  assign n8868 = n8862 & ~n8867;
  assign n8869 = pi76 & ~pi84;
  assign n8870 = n2468 & n8869;
  assign n8871 = ~pi68 & ~pi73;
  assign n8872 = ~pi49 & ~pi66;
  assign n8873 = n8871 & n8872;
  assign n8874 = n8870 & n8873;
  assign n8875 = ~pi89 & ~pi102;
  assign n8876 = n7429 & n8875;
  assign n8877 = ~pi64 & ~pi81;
  assign n8878 = n2476 & n8877;
  assign n8879 = n8876 & n8878;
  assign n8880 = n8874 & n8879;
  assign n8881 = n2451 & n2641;
  assign n8882 = ~pi103 & n2460;
  assign n8883 = n8881 & n8882;
  assign n8884 = n2455 & n2606;
  assign n8885 = ~pi45 & ~pi48;
  assign n8886 = ~pi61 & ~pi104;
  assign n8887 = n8885 & n8886;
  assign n8888 = n8884 & n8887;
  assign n8889 = n8883 & n8888;
  assign n8890 = n8880 & n8889;
  assign n8891 = ~n8856 & ~n8890;
  assign n8892 = n2486 & n2491;
  assign n8893 = ~n8891 & n8892;
  assign n8894 = ~pi24 & ~n8893;
  assign n8895 = n2484 & n8890;
  assign n8896 = n8859 & n8895;
  assign n8897 = pi24 & ~n8896;
  assign n8898 = n2550 & n2783;
  assign n8899 = n7437 & n8898;
  assign n8900 = n8867 & n8899;
  assign n8901 = ~n8897 & n8900;
  assign n8902 = ~n8894 & n8901;
  assign n8903 = ~n8868 & ~n8902;
  assign n8904 = ~pi32 & ~n8903;
  assign n8905 = ~pi24 & ~pi841;
  assign n8906 = pi32 & ~n8905;
  assign n8907 = n2499 & n8906;
  assign n8908 = ~n8904 & ~n8907;
  assign n8909 = ~n6143 & ~n8908;
  assign n8910 = ~pi32 & ~n8862;
  assign n8911 = n6143 & ~n6147;
  assign n8912 = ~n8910 & n8911;
  assign n8913 = ~n8909 & ~n8912;
  assign n8914 = ~pi95 & n3276;
  assign n8915 = ~n8913 & n8914;
  assign n8916 = ~n8853 & ~n8915;
  assign n8917 = n3230 & ~n8916;
  assign n8918 = ~pi24 & n2548;
  assign n8919 = n2494 & n3093;
  assign n8920 = ~pi51 & n8919;
  assign n8921 = n8918 & n8920;
  assign n8922 = ~po840 & n8921;
  assign n8923 = pi252 & ~n8848;
  assign n8924 = ~pi87 & n3181;
  assign n8925 = pi75 & ~pi100;
  assign n8926 = n8924 & n8925;
  assign n8927 = ~pi137 & n8926;
  assign n8928 = ~n6263 & n8927;
  assign n8929 = ~n8923 & n8928;
  assign n8930 = n8922 & n8929;
  assign n8931 = ~n8917 & ~n8930;
  assign po190 = n8841 & ~n8931;
  assign n8933 = ~pi195 & ~pi196;
  assign n8934 = ~pi138 & n8933;
  assign n8935 = ~pi139 & n8934;
  assign n8936 = ~pi118 & n8935;
  assign n8937 = ~pi79 & n8936;
  assign n8938 = ~pi34 & n8937;
  assign n8939 = ~pi33 & ~n8938;
  assign n8940 = pi149 & pi157;
  assign n8941 = ~pi149 & ~pi157;
  assign n8942 = n6162 & ~n8941;
  assign n8943 = ~n8940 & n8942;
  assign n8944 = pi232 & n8943;
  assign n8945 = pi75 & ~n8944;
  assign n8946 = pi100 & ~n8944;
  assign n8947 = ~n8945 & ~n8946;
  assign n8948 = ~pi75 & ~pi100;
  assign n8949 = n7462 & n8948;
  assign n8950 = pi169 & n8949;
  assign n8951 = n8947 & ~n8950;
  assign n8952 = pi74 & ~n8951;
  assign n8953 = pi164 & n8949;
  assign n8954 = n8947 & ~n8953;
  assign n8955 = ~pi74 & ~n8954;
  assign n8956 = ~n3429 & ~n8955;
  assign n8957 = ~n8952 & n8956;
  assign n8958 = pi178 & pi183;
  assign n8959 = ~pi178 & ~pi183;
  assign n8960 = n6162 & ~n8959;
  assign n8961 = ~n8958 & n8960;
  assign n8962 = ~pi299 & ~n8961;
  assign n8963 = pi299 & ~n8943;
  assign n8964 = pi232 & ~n8963;
  assign n8965 = ~n8962 & n8964;
  assign n8966 = pi100 & ~n8965;
  assign n8967 = pi75 & ~n8965;
  assign n8968 = ~n8966 & ~n8967;
  assign n8969 = pi191 & ~pi299;
  assign n8970 = pi169 & pi299;
  assign n8971 = ~n8969 & ~n8970;
  assign n8972 = n8949 & ~n8971;
  assign n8973 = n8968 & ~n8972;
  assign n8974 = pi74 & ~n8973;
  assign n8975 = ~pi55 & ~n8974;
  assign n8976 = ~pi186 & ~pi299;
  assign n8977 = ~pi164 & pi299;
  assign n8978 = ~n8976 & ~n8977;
  assign n8979 = n7462 & n8978;
  assign n8980 = n8948 & n8979;
  assign n8981 = n8968 & ~n8980;
  assign n8982 = pi54 & ~n8981;
  assign n8983 = pi299 & n7462;
  assign n8984 = ~n6109 & n8983;
  assign n8985 = ~pi186 & ~n8984;
  assign n8986 = ~n6234 & n7462;
  assign n8987 = pi186 & ~n8986;
  assign n8988 = pi164 & ~n8987;
  assign n8989 = ~n8985 & n8988;
  assign n8990 = ~pi299 & n7462;
  assign n8991 = ~n6109 & n8990;
  assign n8992 = ~pi164 & pi186;
  assign n8993 = n8991 & n8992;
  assign n8994 = ~n8989 & ~n8993;
  assign n8995 = pi38 & ~n8994;
  assign n8996 = ~pi176 & pi232;
  assign n8997 = ~pi40 & n2476;
  assign n8998 = ~pi102 & n8877;
  assign n8999 = n2455 & n8998;
  assign n9000 = n2453 & n8999;
  assign n9001 = n2474 & n9000;
  assign n9002 = ~pi60 & n9001;
  assign n9003 = n2505 & n2513;
  assign n9004 = ~pi53 & n9003;
  assign n9005 = n9002 & n9004;
  assign n9006 = ~pi58 & n9005;
  assign n9007 = n7437 & n9006;
  assign n9008 = ~pi32 & n2551;
  assign n9009 = n9007 & n9008;
  assign n9010 = ~pi95 & n9009;
  assign n9011 = n6438 & ~n6450;
  assign n9012 = n6170 & n9011;
  assign n9013 = ~n6201 & ~n9012;
  assign n9014 = n9010 & ~n9013;
  assign n9015 = n6198 & n9014;
  assign n9016 = n8997 & ~n9015;
  assign n9017 = pi224 & n6461;
  assign n9018 = n8997 & ~n9017;
  assign n9019 = ~n9016 & ~n9018;
  assign n9020 = n9010 & n9012;
  assign n9021 = n6162 & n9020;
  assign n9022 = n8997 & ~n9021;
  assign n9023 = ~n6215 & ~n9022;
  assign n9024 = ~n9018 & n9023;
  assign n9025 = pi174 & n9024;
  assign n9026 = ~n9019 & ~n9025;
  assign n9027 = ~pi299 & ~n9026;
  assign n9028 = pi216 & n6434;
  assign n9029 = n8997 & ~n9028;
  assign n9030 = pi299 & ~n9029;
  assign n9031 = n6201 & n9010;
  assign n9032 = ~n6192 & n9031;
  assign n9033 = n8997 & ~n9032;
  assign n9034 = n6162 & n9033;
  assign n9035 = ~pi152 & n9034;
  assign n9036 = n6162 & n9014;
  assign n9037 = n8997 & ~n9036;
  assign n9038 = ~n6189 & ~n9037;
  assign n9039 = n9016 & ~n9038;
  assign n9040 = ~pi154 & ~n9039;
  assign n9041 = ~n9035 & n9040;
  assign n9042 = n8997 & ~n9020;
  assign n9043 = n6199 & ~n9042;
  assign n9044 = pi152 & n9043;
  assign n9045 = n9016 & ~n9044;
  assign n9046 = pi154 & ~n9045;
  assign n9047 = n9028 & ~n9046;
  assign n9048 = ~n9041 & n9047;
  assign n9049 = n9030 & ~n9048;
  assign n9050 = ~n9027 & ~n9049;
  assign n9051 = n6220 & n9031;
  assign n9052 = n8997 & n9017;
  assign n9053 = ~n9051 & n9052;
  assign n9054 = ~n9018 & ~n9053;
  assign n9055 = ~pi299 & n9054;
  assign n9056 = n9050 & ~n9055;
  assign n9057 = n8996 & ~n9056;
  assign n9058 = pi176 & pi232;
  assign n9059 = ~n9050 & n9058;
  assign n9060 = n9030 & ~n9039;
  assign n9061 = ~n6215 & ~n9037;
  assign n9062 = ~n9018 & n9061;
  assign n9063 = ~n9019 & ~n9062;
  assign n9064 = ~pi299 & ~n9063;
  assign n9065 = ~n9060 & ~n9064;
  assign n9066 = ~pi232 & ~n9065;
  assign n9067 = pi39 & ~n9066;
  assign n9068 = ~n9059 & n9067;
  assign n9069 = ~n9057 & n9068;
  assign n9070 = pi95 & ~n8997;
  assign n9071 = ~n2449 & ~n9070;
  assign n9072 = ~pi40 & ~pi479;
  assign n9073 = n2476 & ~n9009;
  assign n9074 = n9072 & n9073;
  assign n9075 = ~n9071 & ~n9074;
  assign n9076 = pi32 & ~n8997;
  assign n9077 = n2476 & ~n2549;
  assign n9078 = n2476 & ~n9007;
  assign n9079 = pi70 & ~n9078;
  assign n9080 = n2476 & ~n9005;
  assign n9081 = pi58 & ~n9080;
  assign n9082 = pi53 & ~n9002;
  assign n9083 = ~pi60 & n8856;
  assign n9084 = n2504 & ~n9083;
  assign n9085 = ~n9082 & ~n9084;
  assign n9086 = ~pi111 & n2456;
  assign n9087 = ~pi68 & n2457;
  assign n9088 = ~pi36 & n9087;
  assign n9089 = n9086 & n9088;
  assign n9090 = ~pi66 & ~pi84;
  assign n9091 = pi73 & ~pi82;
  assign n9092 = n9090 & n9091;
  assign n9093 = n9089 & n9092;
  assign n9094 = n9000 & n9093;
  assign n9095 = n2466 & n9094;
  assign n9096 = n2483 & n9095;
  assign n9097 = n2476 & ~n9096;
  assign n9098 = ~n9085 & n9097;
  assign n9099 = n2505 & ~n9098;
  assign n9100 = ~n2476 & ~n2505;
  assign n9101 = n2513 & ~n9100;
  assign n9102 = ~n9099 & n9101;
  assign n9103 = n2476 & ~n2513;
  assign n9104 = ~pi58 & ~n9103;
  assign n9105 = ~n9102 & n9104;
  assign n9106 = ~n9081 & ~n9105;
  assign n9107 = ~pi90 & ~n9106;
  assign n9108 = ~pi841 & n9006;
  assign n9109 = n2476 & ~n9108;
  assign n9110 = pi90 & ~n9109;
  assign n9111 = n2547 & ~n9110;
  assign n9112 = ~n9107 & n9111;
  assign n9113 = n2476 & ~n2547;
  assign n9114 = ~pi70 & ~n9113;
  assign n9115 = ~n9112 & n9114;
  assign n9116 = ~n9079 & ~n9115;
  assign n9117 = ~pi51 & ~n9116;
  assign n9118 = pi51 & ~n2476;
  assign n9119 = n2549 & ~n9118;
  assign n9120 = ~n9117 & n9119;
  assign n9121 = ~n9077 & ~n9120;
  assign n9122 = ~pi40 & ~n9121;
  assign n9123 = ~pi32 & ~n9122;
  assign n9124 = ~n9076 & ~n9123;
  assign n9125 = ~pi95 & ~n9124;
  assign n9126 = ~n9075 & ~n9125;
  assign n9127 = n2493 & n6144;
  assign n9128 = n9108 & n9127;
  assign n9129 = n8997 & ~n9128;
  assign n9130 = pi32 & ~n9129;
  assign n9131 = ~n9123 & ~n9130;
  assign n9132 = ~pi95 & ~n9131;
  assign n9133 = ~pi198 & n9132;
  assign n9134 = n9126 & ~n9133;
  assign n9135 = ~n6162 & n9134;
  assign n9136 = n9003 & n9085;
  assign n9137 = n2476 & ~n9136;
  assign n9138 = ~pi58 & ~n9137;
  assign n9139 = ~n9081 & ~n9138;
  assign n9140 = ~pi90 & ~n9139;
  assign n9141 = n9111 & ~n9140;
  assign n9142 = n9114 & ~n9141;
  assign n9143 = ~n9079 & ~n9142;
  assign n9144 = ~pi51 & ~n9143;
  assign n9145 = n9119 & ~n9144;
  assign n9146 = ~n9077 & ~n9145;
  assign n9147 = ~pi40 & ~n9146;
  assign n9148 = ~pi32 & ~n9147;
  assign n9149 = ~n9130 & ~n9148;
  assign n9150 = ~pi95 & ~n9149;
  assign n9151 = ~pi198 & n9150;
  assign n9152 = n6162 & ~n9070;
  assign n9153 = ~n9076 & ~n9148;
  assign n9154 = ~pi95 & ~n9153;
  assign n9155 = n9152 & ~n9154;
  assign n9156 = ~n9151 & n9155;
  assign n9157 = ~n9135 & ~n9156;
  assign n9158 = ~pi183 & ~n9157;
  assign n9159 = ~pi40 & ~n9076;
  assign n9160 = n2476 & ~n6144;
  assign n9161 = ~pi32 & ~n9160;
  assign n9162 = pi93 & ~n2476;
  assign n9163 = n6144 & ~n9162;
  assign n9164 = n2476 & ~n9081;
  assign n9165 = ~pi90 & ~n9164;
  assign n9166 = ~n9110 & ~n9165;
  assign n9167 = ~pi93 & ~n9166;
  assign n9168 = n9163 & ~n9167;
  assign n9169 = n9161 & ~n9168;
  assign n9170 = n9159 & ~n9169;
  assign n9171 = ~pi95 & ~n9170;
  assign n9172 = n9152 & ~n9171;
  assign n9173 = ~n9135 & ~n9172;
  assign n9174 = pi183 & ~n9173;
  assign n9175 = ~n9158 & ~n9174;
  assign n9176 = ~pi95 & n9175;
  assign n9177 = ~pi174 & ~n9075;
  assign n9178 = ~n9176 & n9177;
  assign n9179 = pi183 & n6162;
  assign n9180 = ~n9134 & ~n9179;
  assign n9181 = n8892 & n9095;
  assign n9182 = ~pi90 & n9181;
  assign n9183 = n9166 & ~n9182;
  assign n9184 = ~pi93 & ~n9183;
  assign n9185 = n9163 & ~n9184;
  assign n9186 = n9161 & ~n9185;
  assign n9187 = n9159 & ~n9186;
  assign n9188 = ~pi95 & ~n9187;
  assign n9189 = ~n9075 & ~n9188;
  assign n9190 = n6162 & ~n9189;
  assign n9191 = pi183 & n9190;
  assign n9192 = pi174 & ~n9191;
  assign n9193 = ~n9180 & n9192;
  assign n9194 = ~pi180 & ~n9193;
  assign n9195 = ~n9178 & n9194;
  assign n9196 = n9152 & ~n9188;
  assign n9197 = ~n9135 & ~n9196;
  assign n9198 = pi183 & ~n9197;
  assign n9199 = ~pi40 & n6162;
  assign n9200 = ~n9070 & ~n9125;
  assign n9201 = ~n9133 & n9200;
  assign n9202 = n9199 & n9201;
  assign n9203 = ~n9135 & ~n9202;
  assign n9204 = ~pi183 & ~n9203;
  assign n9205 = ~n9198 & ~n9204;
  assign n9206 = pi174 & ~n9205;
  assign n9207 = ~pi174 & ~n9175;
  assign n9208 = pi180 & ~n9207;
  assign n9209 = ~n9206 & n9208;
  assign n9210 = ~n9195 & ~n9209;
  assign n9211 = ~pi193 & ~n9210;
  assign n9212 = ~pi40 & ~n2476;
  assign n9213 = pi95 & ~n9212;
  assign n9214 = pi32 & ~n9212;
  assign n9215 = n2518 & n2547;
  assign n9216 = ~n2476 & ~n9215;
  assign n9217 = n7437 & n9138;
  assign n9218 = ~n9216 & ~n9217;
  assign n9219 = ~pi70 & ~n9218;
  assign n9220 = ~n9079 & ~n9219;
  assign n9221 = ~pi51 & ~n9220;
  assign n9222 = n9119 & ~n9221;
  assign n9223 = ~n9077 & ~n9222;
  assign n9224 = ~pi40 & n9223;
  assign n9225 = ~pi32 & ~n9224;
  assign n9226 = ~n9214 & ~n9225;
  assign n9227 = ~pi95 & ~n9226;
  assign n9228 = ~n9213 & ~n9227;
  assign n9229 = pi198 & ~n9228;
  assign n9230 = ~pi40 & ~n9129;
  assign n9231 = pi32 & ~n9230;
  assign n9232 = ~n9225 & ~n9231;
  assign n9233 = ~pi95 & ~n9232;
  assign n9234 = ~n9213 & ~n9233;
  assign n9235 = ~pi198 & ~n9234;
  assign n9236 = ~n9229 & ~n9235;
  assign n9237 = n9199 & ~n9236;
  assign n9238 = ~n9135 & ~n9237;
  assign n9239 = ~pi183 & ~n9238;
  assign n9240 = n6162 & ~n8997;
  assign n9241 = ~n6162 & ~n9134;
  assign n9242 = ~n9240 & ~n9241;
  assign n9243 = pi183 & n9242;
  assign n9244 = ~pi174 & ~n9243;
  assign n9245 = ~n9239 & n9244;
  assign n9246 = n7437 & n9105;
  assign n9247 = ~n9216 & ~n9246;
  assign n9248 = ~pi70 & ~n9247;
  assign n9249 = ~n9079 & ~n9248;
  assign n9250 = ~pi51 & ~n9249;
  assign n9251 = n9119 & ~n9250;
  assign n9252 = ~pi40 & ~n9077;
  assign n9253 = ~n9251 & n9252;
  assign n9254 = ~pi32 & ~n9253;
  assign n9255 = ~n9214 & ~n9254;
  assign n9256 = ~n2783 & ~n8997;
  assign n9257 = ~n9255 & ~n9256;
  assign n9258 = ~pi95 & ~n9257;
  assign n9259 = ~n9070 & ~n9258;
  assign n9260 = ~n9231 & ~n9254;
  assign n9261 = ~pi95 & ~n9260;
  assign n9262 = ~n9213 & ~n9261;
  assign n9263 = n9259 & ~n9262;
  assign n9264 = ~pi198 & ~n9263;
  assign n9265 = n6162 & ~n9264;
  assign n9266 = n9259 & n9265;
  assign n9267 = ~n9135 & ~n9266;
  assign n9268 = ~pi183 & ~n9267;
  assign n9269 = n8892 & n9127;
  assign n9270 = ~pi32 & n9269;
  assign n9271 = n9095 & n9270;
  assign n9272 = n8997 & ~n9271;
  assign n9273 = ~pi95 & ~n9272;
  assign n9274 = n9152 & ~n9273;
  assign n9275 = ~n9135 & ~n9274;
  assign n9276 = pi183 & ~n9275;
  assign n9277 = pi174 & ~n9276;
  assign n9278 = ~n9268 & n9277;
  assign n9279 = pi180 & ~n9278;
  assign n9280 = ~n9245 & n9279;
  assign n9281 = ~n9075 & ~n9258;
  assign n9282 = ~n9240 & ~n9265;
  assign n9283 = n9281 & ~n9282;
  assign n9284 = ~n9135 & ~n9283;
  assign n9285 = ~pi183 & ~n9284;
  assign n9286 = n6162 & ~n9273;
  assign n9287 = ~n9075 & n9286;
  assign n9288 = ~n9135 & ~n9287;
  assign n9289 = pi183 & ~n9288;
  assign n9290 = pi174 & ~n9289;
  assign n9291 = ~n9285 & n9290;
  assign n9292 = ~pi95 & ~n8997;
  assign n9293 = ~n9075 & ~n9292;
  assign n9294 = n6162 & n9293;
  assign n9295 = ~n9135 & ~n9294;
  assign n9296 = pi183 & ~n9295;
  assign n9297 = ~pi40 & ~n9223;
  assign n9298 = ~pi32 & ~n9297;
  assign n9299 = ~n9076 & ~n9298;
  assign n9300 = ~pi95 & ~n9299;
  assign n9301 = ~n9075 & ~n9300;
  assign n9302 = ~n9130 & ~n9298;
  assign n9303 = ~pi95 & ~n9302;
  assign n9304 = ~pi198 & n9303;
  assign n9305 = n9301 & ~n9304;
  assign n9306 = n6162 & ~n9305;
  assign n9307 = ~n9241 & ~n9306;
  assign n9308 = ~pi183 & n9307;
  assign n9309 = ~pi174 & ~n9308;
  assign n9310 = ~n9296 & n9309;
  assign n9311 = ~pi180 & ~n9310;
  assign n9312 = ~n9291 & n9311;
  assign n9313 = pi193 & ~n9312;
  assign n9314 = ~n9280 & n9313;
  assign n9315 = ~n9211 & ~n9314;
  assign n9316 = ~pi299 & ~n9315;
  assign n9317 = pi158 & pi299;
  assign n9318 = ~pi210 & n9132;
  assign n9319 = n9126 & ~n9318;
  assign n9320 = ~n6162 & ~n9319;
  assign n9321 = n9200 & ~n9318;
  assign n9322 = n6162 & ~n9321;
  assign n9323 = ~n9320 & ~n9322;
  assign n9324 = pi152 & n9323;
  assign n9325 = ~n6162 & n9319;
  assign n9326 = ~pi210 & n9150;
  assign n9327 = n9155 & ~n9326;
  assign n9328 = ~n9325 & ~n9327;
  assign n9329 = ~pi152 & ~n9328;
  assign n9330 = ~pi172 & ~n9329;
  assign n9331 = ~n9324 & n9330;
  assign n9332 = ~pi210 & ~n9263;
  assign n9333 = n6162 & ~n9332;
  assign n9334 = n9259 & n9333;
  assign n9335 = ~n9325 & ~n9334;
  assign n9336 = pi152 & ~n9335;
  assign n9337 = ~n9070 & ~n9303;
  assign n9338 = ~pi210 & ~n9337;
  assign n9339 = n6162 & ~n9338;
  assign n9340 = ~n9070 & ~n9300;
  assign n9341 = n9339 & n9340;
  assign n9342 = ~n9325 & ~n9341;
  assign n9343 = ~pi152 & ~n9342;
  assign n9344 = pi172 & ~n9343;
  assign n9345 = ~n9336 & n9344;
  assign n9346 = ~n9331 & ~n9345;
  assign n9347 = n9317 & ~n9346;
  assign n9348 = ~n9240 & ~n9333;
  assign n9349 = n9281 & ~n9348;
  assign n9350 = pi152 & ~n9349;
  assign n9351 = ~n9240 & ~n9339;
  assign n9352 = n9301 & ~n9351;
  assign n9353 = ~pi152 & ~n9352;
  assign n9354 = pi172 & ~n9353;
  assign n9355 = ~n9350 & n9354;
  assign n9356 = pi152 & ~n9319;
  assign n9357 = ~n9075 & ~n9154;
  assign n9358 = ~n9326 & n9357;
  assign n9359 = n6162 & n9358;
  assign n9360 = ~pi152 & ~n9359;
  assign n9361 = ~pi172 & ~n9360;
  assign n9362 = ~n9356 & n9361;
  assign n9363 = ~pi158 & pi299;
  assign n9364 = ~n9325 & n9363;
  assign n9365 = ~n9362 & n9364;
  assign n9366 = ~n9355 & n9365;
  assign n9367 = ~pi149 & ~n9366;
  assign n9368 = ~n9347 & n9367;
  assign n9369 = ~n9172 & ~n9325;
  assign n9370 = ~pi152 & ~n9369;
  assign n9371 = ~n9196 & ~n9325;
  assign n9372 = pi152 & ~n9371;
  assign n9373 = ~pi172 & ~n9372;
  assign n9374 = ~n9370 & n9373;
  assign n9375 = ~n9240 & ~n9320;
  assign n9376 = ~pi152 & n9375;
  assign n9377 = ~n9274 & ~n9325;
  assign n9378 = pi152 & ~n9377;
  assign n9379 = pi172 & ~n9378;
  assign n9380 = ~n9376 & n9379;
  assign n9381 = ~n9374 & ~n9380;
  assign n9382 = ~pi95 & ~n9381;
  assign n9383 = ~n9075 & ~n9382;
  assign n9384 = n9363 & ~n9383;
  assign n9385 = n9317 & ~n9381;
  assign n9386 = pi149 & ~n9385;
  assign n9387 = ~n9384 & n9386;
  assign n9388 = ~n9368 & ~n9387;
  assign n9389 = ~n9316 & ~n9388;
  assign n9390 = pi232 & ~n9389;
  assign n9391 = ~n6143 & n9132;
  assign n9392 = n9126 & ~n9391;
  assign n9393 = ~pi232 & ~n9392;
  assign n9394 = ~pi39 & ~n9393;
  assign n9395 = ~n9390 & n9394;
  assign n9396 = ~n9069 & ~n9395;
  assign n9397 = ~pi38 & ~n9396;
  assign n9398 = ~n8995 & ~n9397;
  assign n9399 = ~pi100 & ~n9398;
  assign n9400 = ~pi87 & ~n8966;
  assign n9401 = ~n9399 & n9400;
  assign n9402 = pi38 & n8979;
  assign n9403 = ~pi100 & n9402;
  assign n9404 = ~n8966 & ~n9403;
  assign n9405 = n3206 & n8997;
  assign n9406 = pi87 & ~n9405;
  assign n9407 = n9404 & n9406;
  assign n9408 = n3237 & ~n9407;
  assign n9409 = ~n9401 & n9408;
  assign n9410 = ~pi75 & pi92;
  assign n9411 = pi232 & ~n3391;
  assign n9412 = ~pi176 & ~pi299;
  assign n9413 = n6162 & ~n9412;
  assign n9414 = n9411 & n9413;
  assign n9415 = n3221 & n9010;
  assign n9416 = ~n9414 & n9415;
  assign n9417 = n9405 & ~n9416;
  assign n9418 = n9404 & ~n9417;
  assign n9419 = n9410 & ~n9418;
  assign n9420 = ~n8967 & ~n9419;
  assign n9421 = ~n9409 & n9420;
  assign n9422 = ~pi54 & ~n9421;
  assign n9423 = ~n8982 & ~n9422;
  assign n9424 = ~pi74 & ~n9423;
  assign n9425 = n8975 & ~n9424;
  assign n9426 = pi55 & ~n8952;
  assign n9427 = pi54 & ~n8954;
  assign n9428 = ~pi92 & ~n8945;
  assign n9429 = pi164 & n7462;
  assign n9430 = pi38 & ~n9429;
  assign n9431 = n3240 & ~n9430;
  assign n9432 = pi149 & n7462;
  assign n9433 = ~pi39 & ~n9432;
  assign n9434 = n9010 & n9433;
  assign n9435 = n8997 & ~n9434;
  assign n9436 = ~pi38 & ~n9435;
  assign n9437 = n9431 & ~n9436;
  assign n9438 = ~pi38 & ~n8997;
  assign n9439 = ~pi100 & ~n9438;
  assign n9440 = ~n9430 & n9439;
  assign n9441 = pi87 & n9440;
  assign n9442 = ~n8946 & ~n9441;
  assign n9443 = ~n9437 & n9442;
  assign n9444 = ~pi75 & ~n9443;
  assign n9445 = n9428 & ~n9444;
  assign n9446 = ~pi75 & n9440;
  assign n9447 = pi92 & n8947;
  assign n9448 = ~n9446 & n9447;
  assign n9449 = ~pi54 & ~n9448;
  assign n9450 = ~n9445 & n9449;
  assign n9451 = ~n9427 & ~n9450;
  assign n9452 = ~pi74 & ~n9451;
  assign n9453 = n9426 & ~n9452;
  assign n9454 = n3293 & ~n9453;
  assign n9455 = ~n9425 & n9454;
  assign n9456 = pi38 & n9429;
  assign n9457 = n8948 & n9456;
  assign n9458 = n8947 & ~n9457;
  assign n9459 = ~n9427 & n9458;
  assign n9460 = ~pi74 & ~n9459;
  assign n9461 = ~n8952 & ~n9460;
  assign n9462 = ~n3293 & ~n9461;
  assign n9463 = n3429 & ~n9462;
  assign n9464 = ~pi38 & n8997;
  assign n9465 = n8948 & n9464;
  assign n9466 = n3265 & n9465;
  assign n9467 = ~n3293 & n9466;
  assign n9468 = n9463 & ~n9467;
  assign n9469 = ~n9455 & n9468;
  assign n9470 = ~n8957 & ~n9469;
  assign n9471 = ~n8939 & ~n9470;
  assign n9472 = n6220 & n6451;
  assign n9473 = n9017 & n9472;
  assign n9474 = ~pi174 & n9473;
  assign n9475 = ~pi299 & ~n9474;
  assign n9476 = n8996 & ~n9475;
  assign n9477 = ~n6447 & n9017;
  assign n9478 = n6220 & n9477;
  assign n9479 = ~pi174 & n9478;
  assign n9480 = n6220 & n9017;
  assign n9481 = n7508 & n9480;
  assign n9482 = pi174 & n9481;
  assign n9483 = ~pi299 & ~n9482;
  assign n9484 = ~n9479 & n9483;
  assign n9485 = n9058 & ~n9484;
  assign n9486 = ~n9476 & ~n9485;
  assign n9487 = n6199 & ~n6447;
  assign n9488 = pi154 & ~n9487;
  assign n9489 = n6199 & n6451;
  assign n9490 = ~pi154 & ~n9489;
  assign n9491 = ~pi152 & ~n9490;
  assign n9492 = ~n9488 & n9491;
  assign n9493 = n6162 & n7508;
  assign n9494 = ~n6189 & n9493;
  assign n9495 = pi152 & pi154;
  assign n9496 = n9494 & n9495;
  assign n9497 = ~n9492 & ~n9496;
  assign n9498 = n9028 & ~n9497;
  assign n9499 = pi299 & ~n9498;
  assign n9500 = pi39 & ~n9499;
  assign n9501 = ~n9486 & n9500;
  assign n9502 = pi90 & ~n7424;
  assign n9503 = n2547 & ~n6113;
  assign n9504 = ~n9502 & n9503;
  assign n9505 = ~pi90 & n2514;
  assign n9506 = n2547 & n9505;
  assign n9507 = n2508 & n9506;
  assign n9508 = n2476 & n9507;
  assign n9509 = n9099 & n9508;
  assign n9510 = ~pi70 & ~n9509;
  assign n9511 = ~n9504 & n9510;
  assign n9512 = n2844 & n3093;
  assign n9513 = ~n9511 & n9512;
  assign n9514 = ~n9510 & n9512;
  assign n9515 = ~n6368 & ~n9514;
  assign n9516 = ~pi198 & ~n9515;
  assign n9517 = ~n9513 & ~n9516;
  assign n9518 = n9179 & ~n9517;
  assign n9519 = n3092 & n6162;
  assign n9520 = ~pi40 & n9519;
  assign n9521 = ~pi72 & ~pi93;
  assign n9522 = n2496 & n9521;
  assign n9523 = ~n9502 & n9522;
  assign n9524 = ~n6113 & n9523;
  assign n9525 = n2476 & n9181;
  assign n9526 = n9127 & n9525;
  assign n9527 = ~n9524 & ~n9526;
  assign n9528 = n9520 & ~n9527;
  assign n9529 = ~pi183 & n9528;
  assign n9530 = ~pi174 & ~n9529;
  assign n9531 = ~n9518 & n9530;
  assign n9532 = ~n9084 & n9507;
  assign n9533 = ~pi70 & ~n9532;
  assign n9534 = ~n9504 & n9533;
  assign n9535 = n9512 & ~n9534;
  assign n9536 = ~n6369 & ~n9535;
  assign n9537 = n6162 & ~n9536;
  assign n9538 = pi183 & n9537;
  assign n9539 = n9520 & n9524;
  assign n9540 = ~pi183 & n9539;
  assign n9541 = pi174 & ~n9540;
  assign n9542 = ~n9538 & n9541;
  assign n9543 = ~n9531 & ~n9542;
  assign n9544 = pi193 & ~n9543;
  assign n9545 = ~n6369 & ~n9514;
  assign n9546 = ~pi174 & n9545;
  assign n9547 = n9512 & ~n9533;
  assign n9548 = ~n6369 & ~n9547;
  assign n9549 = pi174 & n9548;
  assign n9550 = n9179 & ~n9549;
  assign n9551 = ~n9546 & n9550;
  assign n9552 = n3092 & n9526;
  assign n9553 = n9199 & n9552;
  assign n9554 = ~pi174 & ~pi183;
  assign n9555 = n9553 & n9554;
  assign n9556 = ~pi193 & ~n9555;
  assign n9557 = ~n9551 & n9556;
  assign n9558 = ~n9544 & ~n9557;
  assign n9559 = n2938 & n6162;
  assign n9560 = pi180 & n9559;
  assign n9561 = ~pi299 & ~n9560;
  assign n9562 = ~n9558 & n9561;
  assign n9563 = ~pi39 & pi232;
  assign n9564 = pi172 & n9513;
  assign n9565 = ~n6413 & ~n9514;
  assign n9566 = ~pi152 & n9565;
  assign n9567 = ~n9564 & n9566;
  assign n9568 = ~n6413 & ~n9547;
  assign n9569 = pi172 & n9535;
  assign n9570 = pi152 & ~n9569;
  assign n9571 = n9568 & n9570;
  assign n9572 = pi149 & n6162;
  assign n9573 = ~n9571 & n9572;
  assign n9574 = ~n9567 & n9573;
  assign n9575 = ~pi152 & n9528;
  assign n9576 = ~n9539 & ~n9575;
  assign n9577 = pi172 & ~n9576;
  assign n9578 = ~pi152 & ~pi172;
  assign n9579 = n9553 & n9578;
  assign n9580 = ~n9577 & ~n9579;
  assign n9581 = ~pi149 & ~n9580;
  assign n9582 = pi158 & n9559;
  assign n9583 = pi299 & ~n9582;
  assign n9584 = ~n9581 & n9583;
  assign n9585 = ~n9574 & n9584;
  assign n9586 = n9563 & ~n9585;
  assign n9587 = ~n9562 & n9586;
  assign n9588 = ~n9501 & ~n9587;
  assign n9589 = ~pi38 & ~n9588;
  assign n9590 = ~pi87 & ~n8995;
  assign n9591 = ~n9589 & n9590;
  assign n9592 = pi87 & ~n9402;
  assign n9593 = ~pi100 & ~n9592;
  assign n9594 = ~n9591 & n9593;
  assign n9595 = ~n8966 & ~n9594;
  assign n9596 = n3237 & ~n9595;
  assign n9597 = ~pi38 & ~pi87;
  assign n9598 = ~pi100 & n9597;
  assign n9599 = n9414 & n9598;
  assign n9600 = n6109 & n9599;
  assign n9601 = n9404 & ~n9600;
  assign n9602 = n9410 & ~n9601;
  assign n9603 = ~n8967 & ~n9602;
  assign n9604 = ~n9596 & n9603;
  assign n9605 = ~pi54 & ~n9604;
  assign n9606 = ~n8982 & ~n9605;
  assign n9607 = ~pi74 & ~n9606;
  assign n9608 = n8975 & ~n9607;
  assign n9609 = n6109 & n9432;
  assign n9610 = ~pi38 & ~n9609;
  assign n9611 = n9431 & ~n9610;
  assign n9612 = n7577 & n9456;
  assign n9613 = ~n8946 & ~n9612;
  assign n9614 = ~n9611 & n9613;
  assign n9615 = ~pi75 & ~n9614;
  assign n9616 = n9428 & ~n9615;
  assign n9617 = pi92 & n9458;
  assign n9618 = ~pi54 & ~n9617;
  assign n9619 = ~n9616 & n9618;
  assign n9620 = ~n9427 & ~n9619;
  assign n9621 = ~pi74 & ~n9620;
  assign n9622 = n9426 & ~n9621;
  assign n9623 = n3293 & ~n9622;
  assign n9624 = ~n9608 & n9623;
  assign n9625 = n9463 & ~n9624;
  assign n9626 = ~n8957 & ~n9625;
  assign n9627 = n8939 & ~n9626;
  assign n9628 = ~pi954 & ~n9627;
  assign n9629 = ~n9471 & n9628;
  assign n9630 = ~pi33 & ~n9470;
  assign n9631 = pi33 & ~n9626;
  assign n9632 = pi954 & ~n9631;
  assign n9633 = ~n9630 & n9632;
  assign po191 = ~n9629 & ~n9633;
  assign n9635 = pi197 & n8941;
  assign n9636 = ~pi197 & ~n8941;
  assign n9637 = ~n9635 & ~n9636;
  assign n9638 = pi162 & n6162;
  assign n9639 = n9637 & ~n9638;
  assign n9640 = n9635 & n9638;
  assign n9641 = ~pi162 & ~pi197;
  assign n9642 = n8942 & ~n9641;
  assign n9643 = n6162 & ~n9642;
  assign n9644 = ~n9640 & n9643;
  assign n9645 = ~n9637 & ~n9644;
  assign n9646 = ~n9639 & ~n9645;
  assign n9647 = pi232 & n9646;
  assign n9648 = ~n8948 & n9647;
  assign n9649 = pi167 & n7462;
  assign n9650 = n8948 & n9649;
  assign n9651 = ~n9648 & ~n9650;
  assign n9652 = ~pi74 & n9651;
  assign n9653 = pi148 & n8949;
  assign n9654 = pi74 & ~n9653;
  assign n9655 = ~n9648 & n9654;
  assign n9656 = ~n9652 & ~n9655;
  assign n9657 = ~n3429 & n9656;
  assign n9658 = ~pi54 & ~n9648;
  assign n9659 = pi38 & n9650;
  assign n9660 = n9658 & ~n9659;
  assign n9661 = ~pi74 & n9660;
  assign n9662 = n9656 & ~n9661;
  assign n9663 = ~n3293 & ~n9662;
  assign n9664 = n3429 & ~n9663;
  assign n9665 = ~n3293 & ~n9466;
  assign n9666 = n3429 & ~n9665;
  assign n9667 = ~n9664 & ~n9666;
  assign n9668 = pi299 & ~n9646;
  assign n9669 = pi140 & pi145;
  assign n9670 = ~pi140 & ~pi145;
  assign n9671 = ~n9669 & ~n9670;
  assign n9672 = n8960 & ~n9671;
  assign n9673 = n8959 & ~n9669;
  assign n9674 = n6162 & ~n9670;
  assign n9675 = n9673 & n9674;
  assign n9676 = ~pi299 & ~n9675;
  assign n9677 = ~n9672 & n9676;
  assign n9678 = pi232 & ~n9677;
  assign n9679 = ~n9668 & n9678;
  assign n9680 = pi100 & ~n9679;
  assign n9681 = pi75 & ~n9679;
  assign n9682 = ~n9680 & ~n9681;
  assign n9683 = pi141 & ~pi299;
  assign n9684 = pi148 & pi299;
  assign n9685 = ~n9683 & ~n9684;
  assign n9686 = n7462 & ~n9685;
  assign n9687 = n8948 & ~n9686;
  assign n9688 = n9682 & ~n9687;
  assign n9689 = pi74 & ~n9688;
  assign n9690 = ~pi55 & ~n9689;
  assign n9691 = pi188 & ~pi299;
  assign n9692 = pi167 & pi299;
  assign n9693 = ~n9691 & ~n9692;
  assign n9694 = n7462 & ~n9693;
  assign n9695 = ~pi100 & ~n9694;
  assign n9696 = ~pi75 & n9695;
  assign n9697 = n9682 & ~n9696;
  assign n9698 = pi54 & ~n9697;
  assign n9699 = ~pi142 & ~n9284;
  assign n9700 = pi142 & n9134;
  assign n9701 = ~pi140 & ~n9700;
  assign n9702 = ~n9699 & n9701;
  assign n9703 = ~pi142 & ~n9288;
  assign n9704 = pi142 & ~n9190;
  assign n9705 = ~n9241 & n9704;
  assign n9706 = pi140 & ~n9705;
  assign n9707 = ~n9703 & n9706;
  assign n9708 = ~n9702 & ~n9707;
  assign n9709 = ~pi181 & ~n9708;
  assign n9710 = ~pi142 & ~n9267;
  assign n9711 = pi142 & ~n9203;
  assign n9712 = ~pi140 & ~n9711;
  assign n9713 = ~n9710 & n9712;
  assign n9714 = ~pi142 & ~n9275;
  assign n9715 = pi142 & ~n9197;
  assign n9716 = pi140 & ~n9715;
  assign n9717 = ~n9714 & n9716;
  assign n9718 = ~n9713 & ~n9717;
  assign n9719 = pi181 & ~n9718;
  assign n9720 = pi144 & ~n9719;
  assign n9721 = ~n9709 & n9720;
  assign n9722 = ~pi142 & ~n9238;
  assign n9723 = pi142 & ~n9157;
  assign n9724 = ~pi140 & ~n9723;
  assign n9725 = ~n9722 & n9724;
  assign n9726 = pi142 & ~n9173;
  assign n9727 = ~pi142 & n9242;
  assign n9728 = pi140 & ~n9727;
  assign n9729 = ~n9726 & n9728;
  assign n9730 = ~n9725 & ~n9729;
  assign n9731 = pi181 & ~n9730;
  assign n9732 = ~pi142 & n9307;
  assign n9733 = ~n9151 & n9357;
  assign n9734 = n6162 & ~n9733;
  assign n9735 = pi142 & ~n9734;
  assign n9736 = ~n9241 & n9735;
  assign n9737 = ~pi140 & ~n9736;
  assign n9738 = ~n9732 & n9737;
  assign n9739 = ~pi142 & ~n9295;
  assign n9740 = ~n9075 & ~n9171;
  assign n9741 = n6162 & ~n9740;
  assign n9742 = pi142 & ~n9741;
  assign n9743 = ~n9241 & n9742;
  assign n9744 = pi140 & ~n9743;
  assign n9745 = ~n9739 & n9744;
  assign n9746 = ~n9738 & ~n9745;
  assign n9747 = ~pi181 & ~n9746;
  assign n9748 = ~pi144 & ~n9747;
  assign n9749 = ~n9731 & n9748;
  assign n9750 = ~pi299 & ~n9749;
  assign n9751 = ~n9721 & n9750;
  assign n9752 = ~pi159 & pi299;
  assign n9753 = ~n9294 & ~n9325;
  assign n9754 = ~pi146 & ~n9753;
  assign n9755 = ~n9320 & ~n9741;
  assign n9756 = pi146 & n9755;
  assign n9757 = ~pi161 & ~n9756;
  assign n9758 = ~n9754 & n9757;
  assign n9759 = ~n9287 & ~n9325;
  assign n9760 = ~pi146 & ~n9759;
  assign n9761 = ~n9190 & ~n9320;
  assign n9762 = pi146 & n9761;
  assign n9763 = pi161 & ~n9762;
  assign n9764 = ~n9760 & n9763;
  assign n9765 = ~n9758 & ~n9764;
  assign n9766 = pi162 & ~n9765;
  assign n9767 = pi161 & ~n9349;
  assign n9768 = ~pi161 & ~n9352;
  assign n9769 = ~pi146 & ~n9768;
  assign n9770 = ~n9767 & n9769;
  assign n9771 = pi161 & ~n9319;
  assign n9772 = ~pi161 & ~n9359;
  assign n9773 = pi146 & ~n9772;
  assign n9774 = ~n9771 & n9773;
  assign n9775 = ~pi162 & ~n9325;
  assign n9776 = ~n9774 & n9775;
  assign n9777 = ~n9770 & n9776;
  assign n9778 = ~n9766 & ~n9777;
  assign n9779 = n9752 & ~n9778;
  assign n9780 = ~pi146 & ~n9377;
  assign n9781 = pi146 & ~n9371;
  assign n9782 = pi161 & ~n9781;
  assign n9783 = ~n9780 & n9782;
  assign n9784 = pi146 & ~n9369;
  assign n9785 = ~pi146 & n9375;
  assign n9786 = ~pi161 & ~n9785;
  assign n9787 = ~n9784 & n9786;
  assign n9788 = pi162 & ~n9787;
  assign n9789 = ~n9783 & n9788;
  assign n9790 = pi159 & pi299;
  assign n9791 = ~pi146 & ~n9342;
  assign n9792 = pi146 & ~n9328;
  assign n9793 = ~pi161 & ~n9792;
  assign n9794 = ~n9791 & n9793;
  assign n9795 = ~pi146 & ~n9335;
  assign n9796 = pi146 & n9323;
  assign n9797 = pi161 & ~n9796;
  assign n9798 = ~n9795 & n9797;
  assign n9799 = ~pi162 & ~n9798;
  assign n9800 = ~n9794 & n9799;
  assign n9801 = n9790 & ~n9800;
  assign n9802 = ~n9789 & n9801;
  assign n9803 = ~n9779 & ~n9802;
  assign n9804 = ~n9751 & n9803;
  assign n9805 = pi232 & ~n9804;
  assign n9806 = ~n9393 & ~n9805;
  assign n9807 = n3181 & ~n9806;
  assign n9808 = pi144 & n9063;
  assign n9809 = ~pi177 & ~pi299;
  assign n9810 = ~pi144 & ~n9019;
  assign n9811 = ~n9054 & n9810;
  assign n9812 = n9809 & ~n9811;
  assign n9813 = ~n9808 & n9812;
  assign n9814 = ~n9019 & ~n9024;
  assign n9815 = pi177 & ~pi299;
  assign n9816 = ~n9810 & n9815;
  assign n9817 = ~n9814 & n9816;
  assign n9818 = ~n9813 & ~n9817;
  assign n9819 = pi232 & ~n9818;
  assign n9820 = ~n9066 & ~n9819;
  assign n9821 = ~pi38 & ~n9820;
  assign n9822 = ~pi161 & n9034;
  assign n9823 = ~n9039 & ~n9822;
  assign n9824 = n9028 & ~n9823;
  assign n9825 = ~pi38 & ~pi155;
  assign n9826 = n9030 & n9825;
  assign n9827 = ~n9824 & n9826;
  assign n9828 = pi161 & n9043;
  assign n9829 = n9016 & n9028;
  assign n9830 = ~n9828 & n9829;
  assign n9831 = ~pi38 & pi155;
  assign n9832 = n9030 & n9831;
  assign n9833 = ~n9830 & n9832;
  assign n9834 = ~n9827 & ~n9833;
  assign n9835 = pi232 & ~n9834;
  assign n9836 = ~n9821 & ~n9835;
  assign n9837 = pi39 & ~n9836;
  assign n9838 = pi188 & n8991;
  assign n9839 = ~pi167 & ~n9838;
  assign n9840 = ~pi188 & ~n8984;
  assign n9841 = pi167 & pi188;
  assign n9842 = ~n8986 & n9841;
  assign n9843 = ~n9840 & ~n9842;
  assign n9844 = ~n9839 & n9843;
  assign n9845 = pi38 & ~n9844;
  assign n9846 = ~pi87 & ~n9845;
  assign n9847 = ~n9837 & n9846;
  assign n9848 = ~n9807 & n9847;
  assign n9849 = pi38 & ~n9694;
  assign n9850 = ~n9438 & ~n9849;
  assign n9851 = pi87 & n9850;
  assign n9852 = ~pi100 & ~n9851;
  assign n9853 = ~n9848 & n9852;
  assign n9854 = ~n9680 & ~n9853;
  assign n9855 = n3237 & ~n9854;
  assign n9856 = pi155 & pi299;
  assign n9857 = ~n9815 & ~n9856;
  assign n9858 = ~pi38 & n9857;
  assign n9859 = n7462 & ~n9858;
  assign n9860 = n9415 & ~n9859;
  assign n9861 = n9850 & ~n9860;
  assign n9862 = ~pi100 & ~n9861;
  assign n9863 = ~n9680 & ~n9862;
  assign n9864 = n9410 & ~n9863;
  assign n9865 = ~n9681 & ~n9864;
  assign n9866 = ~n9855 & n9865;
  assign n9867 = ~pi54 & ~n9866;
  assign n9868 = ~n9698 & ~n9867;
  assign n9869 = ~pi74 & ~n9868;
  assign n9870 = n9690 & ~n9869;
  assign n9871 = pi55 & ~n9655;
  assign n9872 = pi54 & n9651;
  assign n9873 = ~n9465 & n9660;
  assign n9874 = ~n6271 & ~n9873;
  assign n9875 = pi100 & ~n9647;
  assign n9876 = pi38 & n9649;
  assign n9877 = n9415 & ~n9638;
  assign n9878 = n9464 & ~n9877;
  assign n9879 = ~pi100 & ~n9878;
  assign n9880 = ~pi232 & n9415;
  assign n9881 = ~n9879 & ~n9880;
  assign n9882 = ~n9876 & ~n9881;
  assign n9883 = ~n9875 & ~n9882;
  assign n9884 = ~pi75 & ~n9883;
  assign n9885 = pi75 & ~n9647;
  assign n9886 = ~pi92 & ~n9885;
  assign n9887 = ~n9884 & n9886;
  assign n9888 = ~n9874 & ~n9887;
  assign n9889 = ~n9872 & ~n9888;
  assign n9890 = ~pi74 & ~n9889;
  assign n9891 = n9871 & ~n9890;
  assign n9892 = n3293 & ~n9891;
  assign n9893 = ~n9870 & n9892;
  assign n9894 = ~n9667 & ~n9893;
  assign n9895 = ~n9657 & ~n9894;
  assign n9896 = ~pi34 & n9895;
  assign n9897 = ~pi142 & n9528;
  assign n9898 = pi142 & n9553;
  assign n9899 = ~pi140 & ~n9898;
  assign n9900 = ~n9897 & n9899;
  assign n9901 = ~pi142 & n9513;
  assign n9902 = pi140 & n9545;
  assign n9903 = ~n9901 & n9902;
  assign n9904 = ~n9900 & ~n9903;
  assign n9905 = ~pi144 & ~n9904;
  assign n9906 = pi140 & ~n6162;
  assign n9907 = ~pi142 & n9539;
  assign n9908 = ~pi140 & ~n9907;
  assign n9909 = ~pi142 & n9535;
  assign n9910 = pi140 & ~n9909;
  assign n9911 = n9548 & n9910;
  assign n9912 = ~n9908 & ~n9911;
  assign n9913 = pi144 & ~n9912;
  assign n9914 = ~n9906 & ~n9913;
  assign n9915 = ~n9905 & n9914;
  assign n9916 = pi181 & n9559;
  assign n9917 = ~pi299 & ~n9916;
  assign n9918 = ~n9915 & n9917;
  assign n9919 = ~pi146 & ~n9528;
  assign n9920 = pi146 & ~n9553;
  assign n9921 = ~pi161 & ~n9920;
  assign n9922 = ~n9919 & n9921;
  assign n9923 = ~pi146 & pi161;
  assign n9924 = n9539 & n9923;
  assign n9925 = ~n9922 & ~n9924;
  assign n9926 = ~pi162 & ~n9925;
  assign n9927 = ~pi162 & n9559;
  assign n9928 = n9790 & ~n9927;
  assign n9929 = ~n9752 & ~n9928;
  assign n9930 = ~n9638 & ~n9929;
  assign n9931 = ~pi146 & n9513;
  assign n9932 = n9565 & ~n9931;
  assign n9933 = ~pi161 & ~n9932;
  assign n9934 = ~pi146 & n9535;
  assign n9935 = n9568 & ~n9934;
  assign n9936 = pi161 & ~n9935;
  assign n9937 = pi159 & n2938;
  assign n9938 = pi299 & ~n9937;
  assign n9939 = ~n9936 & n9938;
  assign n9940 = ~n9933 & n9939;
  assign n9941 = ~n9930 & ~n9940;
  assign n9942 = ~n9926 & ~n9941;
  assign n9943 = pi232 & ~n9942;
  assign n9944 = ~n9918 & n9943;
  assign n9945 = n3181 & ~n9944;
  assign n9946 = pi161 & ~n9494;
  assign n9947 = ~pi161 & ~n9487;
  assign n9948 = n9028 & ~n9947;
  assign n9949 = ~n9946 & n9948;
  assign n9950 = n9831 & ~n9949;
  assign n9951 = ~pi161 & n9028;
  assign n9952 = n9489 & n9951;
  assign n9953 = n9825 & ~n9952;
  assign n9954 = ~n9950 & ~n9953;
  assign n9955 = pi299 & ~n9954;
  assign n9956 = ~pi144 & n9478;
  assign n9957 = pi144 & n9481;
  assign n9958 = n9815 & ~n9957;
  assign n9959 = ~n9956 & n9958;
  assign n9960 = ~pi144 & n9473;
  assign n9961 = n9809 & ~n9960;
  assign n9962 = pi232 & ~n9961;
  assign n9963 = ~n9959 & n9962;
  assign n9964 = ~pi38 & ~n9963;
  assign n9965 = ~n9955 & ~n9964;
  assign n9966 = pi39 & ~n9965;
  assign n9967 = ~n9845 & ~n9966;
  assign n9968 = ~n9945 & n9967;
  assign n9969 = ~pi100 & ~n9968;
  assign n9970 = ~n9680 & ~n9969;
  assign n9971 = ~pi87 & ~n9970;
  assign n9972 = ~n3206 & ~n9695;
  assign n9973 = ~n9680 & n9972;
  assign n9974 = pi87 & ~n9973;
  assign n9975 = ~n9971 & ~n9974;
  assign n9976 = n3237 & ~n9975;
  assign n9977 = pi38 & ~n9693;
  assign n9978 = n3181 & ~n9857;
  assign n9979 = n3089 & n9978;
  assign n9980 = ~n9977 & ~n9979;
  assign n9981 = n7462 & ~n9980;
  assign n9982 = ~pi100 & ~n9981;
  assign n9983 = ~n9680 & ~n9982;
  assign n9984 = ~pi87 & ~n9983;
  assign n9985 = ~n9974 & ~n9984;
  assign n9986 = n9410 & ~n9985;
  assign n9987 = ~n9681 & ~n9986;
  assign n9988 = ~n9976 & n9987;
  assign n9989 = ~pi54 & ~n9988;
  assign n9990 = ~n9698 & ~n9989;
  assign n9991 = ~pi74 & ~n9990;
  assign n9992 = n9690 & ~n9991;
  assign n9993 = ~pi92 & pi162;
  assign n9994 = n9563 & n9993;
  assign n9995 = n9597 & n9994;
  assign n9996 = n6180 & n9995;
  assign n9997 = ~n9876 & ~n9996;
  assign n9998 = n8948 & ~n9997;
  assign n9999 = n9658 & ~n9998;
  assign n10000 = ~n9872 & ~n9999;
  assign n10001 = ~pi74 & ~n10000;
  assign n10002 = n9871 & ~n10001;
  assign n10003 = n3293 & ~n10002;
  assign n10004 = ~n9992 & n10003;
  assign n10005 = n9664 & ~n10004;
  assign n10006 = ~n9657 & ~n10005;
  assign n10007 = pi34 & n10006;
  assign n10008 = ~pi33 & ~pi954;
  assign n10009 = ~n10007 & ~n10008;
  assign n10010 = ~n9896 & n10009;
  assign n10011 = ~pi34 & ~n8937;
  assign n10012 = n9895 & ~n10011;
  assign n10013 = n10006 & n10011;
  assign n10014 = n10008 & ~n10013;
  assign n10015 = ~n10012 & n10014;
  assign po192 = ~n10010 & ~n10015;
  assign n10017 = pi137 & n8844;
  assign n10018 = pi1091 & pi1093;
  assign n10019 = n2733 & n10018;
  assign n10020 = n7474 & ~n10019;
  assign n10021 = pi683 & n10020;
  assign n10022 = pi252 & po1057;
  assign n10023 = ~n10021 & n10022;
  assign n10024 = ~n6243 & ~n10023;
  assign n10025 = ~n7463 & ~n10024;
  assign n10026 = ~n8847 & ~n10025;
  assign n10027 = n8848 & n10024;
  assign n10028 = ~n10026 & ~n10027;
  assign n10029 = n8846 & ~n10028;
  assign n10030 = ~n10017 & ~n10029;
  assign n10031 = n8842 & ~n10030;
  assign n10032 = ~pi90 & n6112;
  assign n10033 = ~pi93 & ~n10032;
  assign n10034 = ~n6131 & ~n10033;
  assign n10035 = ~pi35 & ~n10034;
  assign n10036 = pi35 & ~n2736;
  assign n10037 = n8898 & ~n10036;
  assign n10038 = ~n10035 & n10037;
  assign n10039 = ~pi32 & n10038;
  assign n10040 = pi32 & ~pi93;
  assign n10041 = n8855 & n10040;
  assign n10042 = n7424 & n10041;
  assign n10043 = ~n10039 & ~n10042;
  assign n10044 = ~pi95 & ~n6143;
  assign n10045 = ~n10043 & n10044;
  assign n10046 = ~n2553 & ~n10038;
  assign n10047 = pi1082 & n3092;
  assign n10048 = ~n10046 & n10047;
  assign n10049 = n6143 & ~n10035;
  assign n10050 = n2734 & n7525;
  assign n10051 = ~pi137 & ~n6143;
  assign n10052 = ~n7697 & ~n10051;
  assign n10053 = n10050 & n10052;
  assign n10054 = ~pi122 & ~po740;
  assign n10055 = n7697 & ~n10051;
  assign n10056 = n10054 & n10055;
  assign n10057 = ~n10053 & ~n10056;
  assign n10058 = ~n10049 & n10057;
  assign n10059 = n2493 & n8896;
  assign n10060 = n10035 & ~n10059;
  assign n10061 = n3092 & n10037;
  assign n10062 = ~n10060 & n10061;
  assign n10063 = ~n10058 & n10062;
  assign n10064 = ~pi38 & ~n10063;
  assign n10065 = ~n10048 & n10064;
  assign n10066 = ~n10045 & n10065;
  assign n10067 = pi38 & ~n8921;
  assign n10068 = ~pi39 & ~pi100;
  assign n10069 = ~n10067 & n10068;
  assign n10070 = ~n10066 & n10069;
  assign n10071 = ~n10031 & ~n10070;
  assign n10072 = n3230 & ~n10071;
  assign n10073 = pi137 & ~po840;
  assign n10074 = ~n6263 & n10073;
  assign n10075 = ~n8923 & ~n10074;
  assign n10076 = n8926 & ~n10075;
  assign n10077 = n8921 & n10076;
  assign n10078 = ~n10072 & ~n10077;
  assign n10079 = ~pi92 & ~n10078;
  assign n10080 = ~pi54 & ~n10079;
  assign n10081 = ~pi24 & n7307;
  assign n10082 = pi54 & ~n10081;
  assign n10083 = n3293 & n8839;
  assign n10084 = ~n10082 & n10083;
  assign n10085 = ~n10080 & n10084;
  assign n10086 = ~pi59 & ~n10085;
  assign n10087 = n3268 & n3293;
  assign n10088 = n8921 & n10087;
  assign n10089 = ~pi55 & n10088;
  assign n10090 = pi59 & ~n10089;
  assign n10091 = ~pi57 & ~n10090;
  assign po193 = ~n10086 & n10091;
  assign n10093 = n2514 & n2580;
  assign n10094 = ~pi83 & n2647;
  assign n10095 = ~pi65 & n2451;
  assign n10096 = n2476 & n10095;
  assign n10097 = n8998 & n10096;
  assign n10098 = ~pi69 & n10097;
  assign n10099 = ~pi67 & ~pi71;
  assign n10100 = pi36 & ~pi103;
  assign n10101 = n10099 & n10100;
  assign n10102 = n10098 & n10101;
  assign n10103 = n10094 & n10102;
  assign n10104 = n10093 & n10103;
  assign n10105 = ~pi58 & n7479;
  assign n10106 = ~n10104 & ~n10105;
  assign n10107 = n2493 & n6360;
  assign n10108 = n6144 & n10107;
  assign n10109 = n3265 & ~po1038;
  assign n10110 = n3406 & n10109;
  assign n10111 = ~pi92 & n10110;
  assign n10112 = n10108 & n10111;
  assign n10113 = po740 & n10112;
  assign po194 = ~n10106 & n10113;
  assign n10115 = ~pi39 & n3093;
  assign n10116 = pi24 & n10115;
  assign n10117 = n2498 & n10116;
  assign n10118 = pi38 & ~n10117;
  assign n10119 = ~pi81 & ~n2598;
  assign n10120 = n6360 & n9215;
  assign n10121 = n2520 & n10120;
  assign n10122 = n2551 & n10121;
  assign n10123 = ~pi71 & n2476;
  assign n10124 = ~pi104 & n2461;
  assign n10125 = n10123 & n10124;
  assign n10126 = ~pi45 & ~pi73;
  assign n10127 = n8872 & n10126;
  assign n10128 = ~pi48 & ~pi65;
  assign n10129 = ~pi82 & ~pi84;
  assign n10130 = pi89 & n10129;
  assign n10131 = n10128 & n10130;
  assign n10132 = n10127 & n10131;
  assign n10133 = n9089 & n10132;
  assign n10134 = n10125 & n10133;
  assign n10135 = pi332 & n10134;
  assign n10136 = ~pi64 & ~n10135;
  assign n10137 = ~pi39 & ~pi841;
  assign n10138 = n2454 & n10137;
  assign n10139 = ~n10136 & n10138;
  assign n10140 = n10122 & n10139;
  assign n10141 = n10119 & n10140;
  assign n10142 = ~pi38 & ~n10141;
  assign n10143 = n3267 & ~po1038;
  assign n10144 = ~n10142 & n10143;
  assign po196 = ~n10118 & n10144;
  assign n10146 = ~pi38 & n10143;
  assign n10147 = ~pi984 & ~n6257;
  assign n10148 = pi835 & ~n10147;
  assign n10149 = n6165 & ~n10148;
  assign n10150 = n6175 & ~n10149;
  assign n10151 = pi1093 & n10150;
  assign n10152 = n6166 & n6435;
  assign n10153 = ~n10151 & n10152;
  assign n10154 = ~pi215 & n10153;
  assign n10155 = ~n6192 & n10150;
  assign n10156 = n10152 & ~n10155;
  assign n10157 = ~n6189 & n10156;
  assign n10158 = n6198 & n10150;
  assign n10159 = n10152 & ~n10158;
  assign n10160 = n6189 & n10159;
  assign n10161 = pi299 & ~n10160;
  assign n10162 = ~n10157 & n10161;
  assign n10163 = ~n10154 & n10162;
  assign n10164 = pi786 & ~pi1082;
  assign n10165 = ~pi223 & n10153;
  assign n10166 = ~n6215 & n10156;
  assign n10167 = n6215 & n10159;
  assign n10168 = ~pi299 & ~n10167;
  assign n10169 = ~n10166 & n10168;
  assign n10170 = ~n10165 & n10169;
  assign n10171 = ~n10164 & ~n10170;
  assign n10172 = ~n10163 & n10171;
  assign n10173 = n5767 & ~n6200;
  assign n10174 = n3474 & ~n6221;
  assign n10175 = ~n10173 & ~n10174;
  assign n10176 = po740 & n10164;
  assign n10177 = ~n10175 & n10176;
  assign n10178 = n6437 & n10177;
  assign n10179 = ~n10172 & ~n10178;
  assign n10180 = pi39 & ~n10179;
  assign n10181 = ~pi39 & ~pi95;
  assign n10182 = n6143 & n6367;
  assign n10183 = n2510 & ~n2583;
  assign n10184 = n8876 & n8881;
  assign n10185 = n9086 & n10184;
  assign n10186 = n8877 & n9090;
  assign n10187 = ~pi65 & ~pi69;
  assign n10188 = n10186 & n10187;
  assign n10189 = pi48 & ~pi49;
  assign n10190 = ~pi68 & ~pi82;
  assign n10191 = n10189 & n10190;
  assign n10192 = n10126 & n10191;
  assign n10193 = n10188 & n10192;
  assign n10194 = n10185 & n10193;
  assign n10195 = n10125 & n10194;
  assign n10196 = ~pi841 & n2483;
  assign n10197 = n2505 & n10196;
  assign n10198 = ~pi97 & n10197;
  assign n10199 = n10195 & n10198;
  assign n10200 = n10183 & n10199;
  assign n10201 = pi108 & n2510;
  assign n10202 = n2582 & n10201;
  assign n10203 = ~pi47 & ~n10202;
  assign n10204 = ~n10200 & n10203;
  assign n10205 = ~pi986 & ~po740;
  assign n10206 = pi252 & ~n10205;
  assign n10207 = pi314 & ~n10206;
  assign n10208 = n6125 & n10207;
  assign n10209 = ~n10204 & n10208;
  assign n10210 = ~pi47 & ~pi841;
  assign n10211 = n10195 & n10210;
  assign n10212 = ~n2569 & ~n10211;
  assign n10213 = n2489 & n2519;
  assign n10214 = ~n10207 & n10213;
  assign n10215 = ~n10212 & n10214;
  assign n10216 = ~n10209 & ~n10215;
  assign n10217 = n2493 & ~n10216;
  assign n10218 = ~pi35 & ~n10217;
  assign n10219 = pi35 & ~n6364;
  assign n10220 = n2551 & ~n10219;
  assign n10221 = n2725 & n10220;
  assign n10222 = ~n10218 & n10221;
  assign n10223 = ~n10182 & ~n10222;
  assign n10224 = n10181 & ~n10223;
  assign n10225 = ~n10180 & ~n10224;
  assign po197 = n10146 & ~n10225;
  assign n10227 = n3092 & ~n3359;
  assign n10228 = pi102 & n2536;
  assign n10229 = n2453 & n10228;
  assign n10230 = n6144 & n10229;
  assign n10231 = n2520 & n10230;
  assign n10232 = n2479 & n10231;
  assign n10233 = ~pi40 & ~n10232;
  assign n10234 = n10227 & ~n10233;
  assign n10235 = ~pi1082 & ~n10234;
  assign n10236 = n6360 & n10232;
  assign n10237 = pi1082 & ~n10236;
  assign n10238 = n10111 & ~n10237;
  assign po198 = ~n10235 & n10238;
  assign n10240 = ~pi41 & ~pi72;
  assign n10241 = ~n8064 & ~n10240;
  assign n10242 = ~n2734 & n10240;
  assign n10243 = n8064 & ~n10242;
  assign n10244 = ~pi44 & n3095;
  assign n10245 = ~pi101 & n10244;
  assign n10246 = n7525 & n10245;
  assign n10247 = n7465 & n10246;
  assign n10248 = pi41 & ~n10247;
  assign n10249 = ~pi41 & pi72;
  assign n10250 = n2734 & ~n10249;
  assign n10251 = ~pi99 & n6252;
  assign n10252 = ~pi72 & pi101;
  assign n10253 = ~pi41 & ~n10252;
  assign n10254 = ~pi24 & n2498;
  assign n10255 = pi252 & n6360;
  assign n10256 = n7525 & n10255;
  assign n10257 = n10254 & n10256;
  assign n10258 = ~pi44 & n10257;
  assign n10259 = n10253 & n10258;
  assign n10260 = ~n10251 & n10259;
  assign n10261 = n10250 & ~n10260;
  assign n10262 = ~n10248 & n10261;
  assign n10263 = n10243 & ~n10262;
  assign n10264 = ~n10241 & ~n10263;
  assign n10265 = ~pi39 & ~n10264;
  assign n10266 = ~pi166 & n6162;
  assign n10267 = pi161 & n10266;
  assign n10268 = ~pi152 & n10267;
  assign n10269 = ~n6237 & ~n10268;
  assign n10270 = ~pi189 & n6162;
  assign n10271 = pi144 & n10270;
  assign n10272 = ~pi174 & n10271;
  assign n10273 = ~pi299 & ~n10272;
  assign n10274 = pi232 & ~n10273;
  assign n10275 = ~n10269 & n10274;
  assign n10276 = ~pi72 & ~n10275;
  assign n10277 = pi39 & ~n10276;
  assign n10278 = n3241 & ~n10277;
  assign n10279 = ~n10265 & n10278;
  assign n10280 = ~pi39 & ~n10240;
  assign n10281 = ~n10277 & ~n10280;
  assign n10282 = ~n3241 & n10281;
  assign n10283 = pi75 & ~n10282;
  assign n10284 = ~n10279 & n10283;
  assign n10285 = n7443 & ~n7449;
  assign n10286 = ~pi1093 & ~n7451;
  assign n10287 = ~n10285 & n10286;
  assign n10288 = ~pi44 & ~n10287;
  assign n10289 = n2761 & ~n7435;
  assign n10290 = n2759 & n10289;
  assign n10291 = ~n7479 & ~n10290;
  assign n10292 = n2518 & ~n10291;
  assign n10293 = n7426 & ~n10292;
  assign n10294 = n7423 & ~n10293;
  assign n10295 = ~pi51 & ~n10294;
  assign n10296 = ~n2558 & ~n10295;
  assign n10297 = ~pi96 & ~n10296;
  assign n10298 = n6360 & ~n7446;
  assign n10299 = ~pi72 & n7449;
  assign n10300 = n10298 & n10299;
  assign n10301 = ~n10297 & n10300;
  assign n10302 = ~n10285 & ~n10301;
  assign n10303 = pi1093 & n10302;
  assign n10304 = n10288 & ~n10303;
  assign n10305 = ~pi101 & n10304;
  assign n10306 = pi41 & ~n10305;
  assign n10307 = ~n7445 & n10298;
  assign n10308 = n10299 & ~n10307;
  assign n10309 = ~pi72 & ~n7443;
  assign n10310 = ~n7449 & n10309;
  assign n10311 = ~pi1093 & ~n10310;
  assign n10312 = ~n10308 & n10311;
  assign n10313 = ~pi72 & n10302;
  assign n10314 = pi1093 & ~n10313;
  assign n10315 = ~n10312 & ~n10314;
  assign n10316 = pi44 & ~pi72;
  assign n10317 = ~n10315 & ~n10316;
  assign n10318 = ~pi101 & ~n10317;
  assign n10319 = n10253 & ~n10318;
  assign n10320 = n2734 & ~n10319;
  assign n10321 = ~n10306 & n10320;
  assign n10322 = pi1093 & ~n7443;
  assign n10323 = n10288 & ~n10322;
  assign n10324 = ~pi101 & n10323;
  assign n10325 = pi41 & ~n10324;
  assign n10326 = n10309 & ~n10312;
  assign n10327 = ~n10316 & ~n10326;
  assign n10328 = ~pi101 & ~n10327;
  assign n10329 = n10253 & ~n10328;
  assign n10330 = ~n2734 & ~n10329;
  assign n10331 = ~n10325 & n10330;
  assign n10332 = pi228 & ~n10331;
  assign n10333 = ~n10321 & n10332;
  assign n10334 = ~pi109 & n6330;
  assign n10335 = n2589 & n10334;
  assign n10336 = ~pi110 & ~n10335;
  assign n10337 = n2489 & ~n2568;
  assign n10338 = ~pi480 & pi949;
  assign n10339 = n2497 & n10338;
  assign n10340 = ~pi47 & n10339;
  assign n10341 = n10337 & n10340;
  assign n10342 = ~n10336 & n10341;
  assign n10343 = pi901 & ~pi959;
  assign n10344 = n2514 & n2589;
  assign n10345 = n2497 & n10344;
  assign n10346 = ~n10338 & n10345;
  assign n10347 = n10343 & ~n10346;
  assign n10348 = ~n10342 & n10347;
  assign n10349 = n2490 & n2567;
  assign n10350 = pi110 & n10349;
  assign n10351 = n10339 & n10350;
  assign n10352 = ~n10343 & ~n10351;
  assign n10353 = ~pi250 & pi252;
  assign n10354 = n6360 & n10353;
  assign n10355 = ~n10352 & n10354;
  assign n10356 = ~n10348 & n10355;
  assign n10357 = ~pi72 & n10356;
  assign n10358 = n10108 & n10350;
  assign n10359 = n10338 & ~n10353;
  assign n10360 = n10358 & n10359;
  assign n10361 = ~n10357 & ~n10360;
  assign n10362 = ~pi44 & ~n10361;
  assign n10363 = ~pi101 & n10362;
  assign n10364 = pi41 & ~n10363;
  assign n10365 = n6360 & ~n10353;
  assign n10366 = n10351 & n10365;
  assign n10367 = ~pi72 & ~n10366;
  assign n10368 = ~n10356 & n10367;
  assign n10369 = ~n10316 & ~n10368;
  assign n10370 = ~pi101 & ~n10369;
  assign n10371 = n10253 & ~n10370;
  assign n10372 = ~n10364 & ~n10371;
  assign n10373 = ~pi228 & ~n10372;
  assign n10374 = ~pi39 & ~n10373;
  assign n10375 = ~n10333 & n10374;
  assign n10376 = pi287 & n3095;
  assign n10377 = n10275 & n10376;
  assign n10378 = ~n10276 & ~n10377;
  assign n10379 = pi39 & ~n10378;
  assign n10380 = n3206 & ~n10379;
  assign n10381 = ~n10375 & n10380;
  assign n10382 = n2498 & n6360;
  assign n10383 = ~pi44 & n10382;
  assign n10384 = n10253 & n10383;
  assign n10385 = ~n10249 & ~n10384;
  assign n10386 = ~pi72 & ~n7525;
  assign n10387 = ~n10385 & ~n10386;
  assign n10388 = ~n10251 & n10387;
  assign n10389 = pi41 & ~n10246;
  assign n10390 = n2734 & ~n10251;
  assign n10391 = ~n10250 & ~n10390;
  assign n10392 = ~n10389 & ~n10391;
  assign n10393 = ~n10388 & n10392;
  assign n10394 = n10243 & ~n10393;
  assign n10395 = ~n10241 & ~n10394;
  assign n10396 = ~pi39 & ~n10395;
  assign n10397 = ~n10277 & ~n10396;
  assign n10398 = n6235 & ~n10397;
  assign n10399 = pi38 & ~n10281;
  assign n10400 = ~pi87 & ~n10399;
  assign n10401 = ~n10398 & n10400;
  assign n10402 = ~n10381 & n10401;
  assign n10403 = pi41 & ~n10245;
  assign n10404 = pi228 & n10385;
  assign n10405 = ~n10403 & n10404;
  assign n10406 = ~pi228 & n10240;
  assign n10407 = n3207 & ~n10406;
  assign n10408 = ~n10405 & n10407;
  assign n10409 = ~n3206 & n10280;
  assign n10410 = pi87 & ~n10409;
  assign n10411 = ~n10277 & n10410;
  assign n10412 = ~n10408 & n10411;
  assign n10413 = ~pi75 & ~n10412;
  assign n10414 = ~n10402 & n10413;
  assign n10415 = ~n10284 & ~n10414;
  assign n10416 = n7422 & ~n10415;
  assign n10417 = ~n7422 & ~n10281;
  assign n10418 = ~po1038 & ~n10417;
  assign n10419 = ~n10416 & n10418;
  assign n10420 = pi39 & pi232;
  assign n10421 = n10268 & n10420;
  assign n10422 = ~pi72 & ~n10280;
  assign n10423 = po1038 & n10422;
  assign n10424 = ~n10421 & n10423;
  assign po199 = ~n10419 & ~n10424;
  assign n10426 = pi211 & pi214;
  assign n10427 = pi212 & n10426;
  assign n10428 = ~pi219 & ~n10427;
  assign n10429 = ~pi115 & n2734;
  assign n10430 = pi42 & ~pi114;
  assign n10431 = ~pi72 & pi116;
  assign n10432 = pi72 & pi113;
  assign n10433 = pi72 & ~n6245;
  assign n10434 = ~pi99 & n10319;
  assign n10435 = ~n10433 & ~n10434;
  assign n10436 = ~pi113 & ~n10435;
  assign n10437 = ~n10432 & ~n10436;
  assign n10438 = ~pi116 & n10437;
  assign n10439 = ~n10431 & ~n10438;
  assign n10440 = n10430 & n10439;
  assign n10441 = pi42 & ~pi72;
  assign n10442 = pi114 & ~n10441;
  assign n10443 = n6245 & n10305;
  assign n10444 = n6249 & n10443;
  assign n10445 = ~pi42 & ~n10444;
  assign n10446 = ~n10442 & ~n10445;
  assign n10447 = ~n10440 & n10446;
  assign n10448 = n10429 & ~n10447;
  assign n10449 = ~pi115 & ~n2734;
  assign n10450 = ~pi99 & n10329;
  assign n10451 = ~n10433 & ~n10450;
  assign n10452 = ~pi113 & ~n10451;
  assign n10453 = ~n10432 & ~n10452;
  assign n10454 = ~n10431 & ~n10453;
  assign n10455 = pi42 & ~n10454;
  assign n10456 = n6245 & n10324;
  assign n10457 = n6249 & n10456;
  assign n10458 = ~pi42 & n10457;
  assign n10459 = ~pi114 & ~n10458;
  assign n10460 = ~n10455 & n10459;
  assign n10461 = ~n10442 & ~n10460;
  assign n10462 = n10449 & ~n10461;
  assign n10463 = pi115 & ~n10441;
  assign n10464 = pi228 & ~n10463;
  assign n10465 = ~n10462 & n10464;
  assign n10466 = ~n10448 & n10465;
  assign n10467 = ~pi99 & n10371;
  assign n10468 = ~n10433 & ~n10467;
  assign n10469 = ~pi72 & pi113;
  assign n10470 = ~n10468 & ~n10469;
  assign n10471 = ~n10431 & n10470;
  assign n10472 = n10430 & n10471;
  assign n10473 = n6245 & n10363;
  assign n10474 = ~pi113 & n10473;
  assign n10475 = ~pi116 & n10474;
  assign n10476 = ~pi42 & ~n10475;
  assign n10477 = ~n10442 & ~n10476;
  assign n10478 = ~n10472 & n10477;
  assign n10479 = ~pi115 & ~n10478;
  assign n10480 = ~pi228 & ~n10463;
  assign n10481 = ~n10479 & n10480;
  assign n10482 = ~pi39 & ~n10481;
  assign n10483 = ~n10466 & n10482;
  assign n10484 = ~pi72 & pi199;
  assign n10485 = ~pi232 & ~n10484;
  assign n10486 = ~pi299 & ~n10485;
  assign n10487 = ~pi72 & ~n10270;
  assign n10488 = n6162 & n10376;
  assign n10489 = ~pi189 & n10488;
  assign n10490 = ~n10487 & ~n10489;
  assign n10491 = pi199 & ~n10490;
  assign n10492 = pi232 & ~n10491;
  assign n10493 = n10486 & ~n10492;
  assign n10494 = pi39 & ~n10493;
  assign n10495 = ~n10483 & ~n10494;
  assign n10496 = n3206 & ~n10495;
  assign n10497 = ~n8064 & ~n10441;
  assign n10498 = ~n10429 & n10441;
  assign n10499 = n8064 & ~n10498;
  assign n10500 = n10429 & ~n10442;
  assign n10501 = n6245 & n10245;
  assign n10502 = n6249 & n10501;
  assign n10503 = n7525 & n10502;
  assign n10504 = ~pi114 & ~n6248;
  assign n10505 = n10503 & n10504;
  assign n10506 = ~pi42 & n10505;
  assign n10507 = n6246 & n10383;
  assign n10508 = n6249 & n10507;
  assign n10509 = ~pi72 & ~n10508;
  assign n10510 = ~n10386 & ~n10509;
  assign n10511 = pi42 & ~n10510;
  assign n10512 = ~pi114 & ~n10511;
  assign n10513 = ~n10506 & n10512;
  assign n10514 = n10500 & ~n10513;
  assign n10515 = n10499 & ~n10514;
  assign n10516 = ~n10497 & ~n10515;
  assign n10517 = ~pi39 & ~n10516;
  assign n10518 = pi199 & n10487;
  assign n10519 = pi232 & ~n10518;
  assign n10520 = n10486 & ~n10519;
  assign n10521 = pi39 & ~n10520;
  assign n10522 = ~n10517 & ~n10521;
  assign n10523 = n6235 & ~n10522;
  assign n10524 = ~pi39 & ~n10441;
  assign n10525 = ~n10521 & ~n10524;
  assign n10526 = pi38 & ~n10525;
  assign n10527 = ~pi87 & ~n10526;
  assign n10528 = ~n10523 & n10527;
  assign n10529 = ~n10496 & n10528;
  assign n10530 = pi228 & n10502;
  assign n10531 = ~pi115 & n10530;
  assign n10532 = ~pi114 & n10531;
  assign n10533 = ~pi42 & n10532;
  assign n10534 = pi228 & n10507;
  assign n10535 = n6251 & n10534;
  assign n10536 = n10441 & ~n10535;
  assign n10537 = n3207 & ~n10536;
  assign n10538 = ~n10533 & n10537;
  assign n10539 = ~n3206 & n10524;
  assign n10540 = pi87 & ~n10539;
  assign n10541 = ~n10538 & n10540;
  assign n10542 = ~n10521 & n10541;
  assign n10543 = ~pi75 & ~n10542;
  assign n10544 = ~n10529 & n10543;
  assign n10545 = n7465 & n10505;
  assign n10546 = ~pi42 & n10545;
  assign n10547 = n6246 & n10258;
  assign n10548 = ~pi113 & n10547;
  assign n10549 = ~pi116 & n10548;
  assign n10550 = n10441 & ~n10549;
  assign n10551 = ~pi114 & ~n10550;
  assign n10552 = ~n10546 & n10551;
  assign n10553 = n10500 & ~n10552;
  assign n10554 = n10499 & ~n10553;
  assign n10555 = n3241 & ~n10497;
  assign n10556 = ~n10554 & n10555;
  assign n10557 = ~n3241 & n10441;
  assign n10558 = ~pi39 & ~n10557;
  assign n10559 = ~n10556 & n10558;
  assign n10560 = ~n10521 & ~n10559;
  assign n10561 = pi75 & ~n10560;
  assign n10562 = n7422 & ~n10561;
  assign n10563 = ~n10544 & n10562;
  assign n10564 = pi207 & pi208;
  assign n10565 = ~n7422 & n10525;
  assign n10566 = ~n10564 & ~n10565;
  assign n10567 = ~n10563 & n10566;
  assign n10568 = ~pi72 & pi200;
  assign n10569 = ~pi232 & ~n10568;
  assign n10570 = ~pi299 & ~n10569;
  assign n10571 = pi200 & n10487;
  assign n10572 = pi232 & ~n10571;
  assign n10573 = n10570 & ~n10572;
  assign n10574 = pi39 & ~n10573;
  assign n10575 = ~n10520 & n10574;
  assign n10576 = ~n10524 & ~n10575;
  assign n10577 = ~n7422 & n10576;
  assign n10578 = n10564 & ~n10577;
  assign n10579 = pi200 & ~n10490;
  assign n10580 = n10492 & ~n10579;
  assign n10581 = ~n10486 & ~n10570;
  assign n10582 = ~n10580 & ~n10581;
  assign n10583 = pi39 & ~n10582;
  assign n10584 = ~n10483 & ~n10583;
  assign n10585 = n3206 & ~n10584;
  assign n10586 = pi38 & ~n10576;
  assign n10587 = ~pi87 & ~n10586;
  assign n10588 = ~n10517 & ~n10575;
  assign n10589 = n6235 & ~n10588;
  assign n10590 = n10587 & ~n10589;
  assign n10591 = ~n10585 & n10590;
  assign n10592 = n10541 & ~n10575;
  assign n10593 = ~pi75 & ~n10592;
  assign n10594 = ~n10591 & n10593;
  assign n10595 = ~n10559 & ~n10575;
  assign n10596 = pi75 & ~n10595;
  assign n10597 = n7422 & ~n10596;
  assign n10598 = ~n10594 & n10597;
  assign n10599 = n10578 & ~n10598;
  assign n10600 = ~n10567 & ~n10599;
  assign n10601 = n10428 & ~n10600;
  assign n10602 = pi232 & ~pi299;
  assign n10603 = ~n10491 & n10602;
  assign n10604 = n10266 & n10376;
  assign n10605 = ~pi166 & n7462;
  assign n10606 = ~pi72 & ~n10605;
  assign n10607 = pi232 & pi299;
  assign n10608 = ~n10606 & n10607;
  assign n10609 = ~n10604 & n10608;
  assign n10610 = pi72 & ~pi232;
  assign n10611 = pi299 & ~n10610;
  assign n10612 = n10485 & ~n10611;
  assign n10613 = ~n10609 & ~n10612;
  assign n10614 = ~n10603 & n10613;
  assign n10615 = pi39 & ~n10614;
  assign n10616 = ~n10483 & ~n10615;
  assign n10617 = n3206 & ~n10616;
  assign n10618 = pi299 & n10606;
  assign n10619 = pi39 & ~n10618;
  assign n10620 = ~n10520 & n10619;
  assign n10621 = ~n10517 & ~n10620;
  assign n10622 = n6235 & ~n10621;
  assign n10623 = ~n10524 & ~n10620;
  assign n10624 = pi38 & ~n10623;
  assign n10625 = ~pi87 & ~n10624;
  assign n10626 = ~n10622 & n10625;
  assign n10627 = ~n10617 & n10626;
  assign n10628 = n10541 & ~n10620;
  assign n10629 = ~pi75 & ~n10628;
  assign n10630 = ~n10627 & n10629;
  assign n10631 = ~n10559 & ~n10620;
  assign n10632 = pi75 & ~n10631;
  assign n10633 = n7422 & ~n10632;
  assign n10634 = ~n10630 & n10633;
  assign n10635 = ~n10564 & ~n10634;
  assign n10636 = ~pi299 & n10580;
  assign n10637 = ~n10568 & n10612;
  assign n10638 = ~n10609 & ~n10637;
  assign n10639 = ~n10636 & n10638;
  assign n10640 = pi39 & ~n10639;
  assign n10641 = ~n10483 & ~n10640;
  assign n10642 = n3206 & ~n10641;
  assign n10643 = n10574 & n10620;
  assign n10644 = ~n10517 & ~n10643;
  assign n10645 = n6235 & ~n10644;
  assign n10646 = ~n10587 & ~n10625;
  assign n10647 = ~n10645 & ~n10646;
  assign n10648 = ~n10642 & n10647;
  assign n10649 = n10540 & ~n10643;
  assign n10650 = ~n10538 & n10649;
  assign n10651 = ~pi75 & ~n10650;
  assign n10652 = ~n10648 & n10651;
  assign n10653 = ~n10559 & ~n10643;
  assign n10654 = pi75 & ~n10653;
  assign n10655 = n7422 & ~n10654;
  assign n10656 = ~n10652 & n10655;
  assign n10657 = n10578 & ~n10656;
  assign n10658 = ~n10635 & ~n10657;
  assign n10659 = ~n7422 & n10623;
  assign n10660 = ~n10428 & ~n10659;
  assign n10661 = ~n10658 & n10660;
  assign n10662 = ~po1038 & ~n10661;
  assign n10663 = ~n10601 & n10662;
  assign n10664 = ~n10428 & n10606;
  assign n10665 = pi39 & ~n10664;
  assign n10666 = po1038 & ~n10524;
  assign n10667 = ~n10665 & n10666;
  assign po200 = n10663 | n10667;
  assign n10669 = pi212 & pi214;
  assign n10670 = ~pi211 & ~pi219;
  assign n10671 = n10669 & ~n10670;
  assign n10672 = ~pi211 & ~n10669;
  assign n10673 = ~n10671 & ~n10672;
  assign n10674 = ~n2734 & n10454;
  assign n10675 = n2734 & n10439;
  assign n10676 = ~n10674 & ~n10675;
  assign n10677 = pi228 & ~n10676;
  assign n10678 = ~pi228 & n10471;
  assign n10679 = ~n10677 & ~n10678;
  assign n10680 = ~pi42 & n6250;
  assign n10681 = pi43 & n10680;
  assign n10682 = ~n10679 & n10681;
  assign n10683 = ~n2734 & ~n10456;
  assign n10684 = n2734 & ~n10443;
  assign n10685 = ~n10683 & ~n10684;
  assign n10686 = ~pi113 & n10685;
  assign n10687 = pi228 & ~n10686;
  assign n10688 = ~pi228 & ~n10475;
  assign n10689 = ~pi116 & ~n10688;
  assign n10690 = ~n10687 & n10689;
  assign n10691 = ~pi43 & ~n10690;
  assign n10692 = pi43 & ~pi72;
  assign n10693 = ~n10680 & ~n10692;
  assign n10694 = ~n10691 & ~n10693;
  assign n10695 = ~n10682 & n10694;
  assign n10696 = ~pi39 & ~n10695;
  assign n10697 = ~n10579 & n10602;
  assign n10698 = n10569 & ~n10611;
  assign n10699 = ~n10609 & ~n10698;
  assign n10700 = ~n10697 & n10699;
  assign n10701 = pi39 & ~n10700;
  assign n10702 = ~n10696 & ~n10701;
  assign n10703 = n3206 & ~n10702;
  assign n10704 = ~n8064 & ~n10692;
  assign n10705 = n2734 & n10680;
  assign n10706 = n10692 & ~n10705;
  assign n10707 = n8064 & ~n10706;
  assign n10708 = ~pi43 & pi52;
  assign n10709 = n10503 & n10708;
  assign n10710 = pi43 & ~n10510;
  assign n10711 = ~n10709 & ~n10710;
  assign n10712 = n10705 & ~n10711;
  assign n10713 = n10707 & ~n10712;
  assign n10714 = ~n10704 & ~n10713;
  assign n10715 = ~pi39 & ~n10714;
  assign n10716 = ~n10573 & n10619;
  assign n10717 = ~n10715 & ~n10716;
  assign n10718 = n6235 & ~n10717;
  assign n10719 = ~pi39 & ~n10692;
  assign n10720 = ~n10716 & ~n10719;
  assign n10721 = pi38 & ~n10720;
  assign n10722 = ~pi87 & ~n10721;
  assign n10723 = ~n10718 & n10722;
  assign n10724 = ~n10703 & n10723;
  assign n10725 = ~pi43 & ~n10502;
  assign n10726 = pi43 & ~n10509;
  assign n10727 = pi228 & n10680;
  assign n10728 = ~n10726 & n10727;
  assign n10729 = ~n10725 & n10728;
  assign n10730 = n10692 & ~n10727;
  assign n10731 = n3207 & ~n10730;
  assign n10732 = ~n10729 & n10731;
  assign n10733 = ~n3206 & n10719;
  assign n10734 = pi87 & ~n10733;
  assign n10735 = ~n10732 & n10734;
  assign n10736 = ~n10716 & n10735;
  assign n10737 = ~pi75 & ~n10736;
  assign n10738 = ~n10724 & n10737;
  assign n10739 = ~pi72 & ~n10549;
  assign n10740 = pi43 & n10739;
  assign n10741 = n7465 & n10503;
  assign n10742 = n10708 & n10741;
  assign n10743 = ~n10740 & ~n10742;
  assign n10744 = n10705 & ~n10743;
  assign n10745 = n10707 & ~n10744;
  assign n10746 = ~n10704 & ~n10745;
  assign n10747 = ~pi39 & ~n10746;
  assign n10748 = n3241 & ~n10747;
  assign n10749 = ~n3241 & ~n10719;
  assign n10750 = ~n10748 & ~n10749;
  assign n10751 = ~n10716 & ~n10750;
  assign n10752 = pi75 & ~n10751;
  assign n10753 = n7422 & ~n10752;
  assign n10754 = ~n10738 & n10753;
  assign n10755 = ~n7422 & n10720;
  assign n10756 = ~n10564 & ~n10755;
  assign n10757 = ~n10754 & n10756;
  assign n10758 = ~pi199 & ~pi200;
  assign n10759 = ~n10490 & n10758;
  assign n10760 = n10602 & ~n10759;
  assign n10761 = ~pi299 & ~n10758;
  assign n10762 = ~pi72 & ~n10761;
  assign n10763 = ~pi232 & ~n10762;
  assign n10764 = ~n10609 & ~n10763;
  assign n10765 = ~n10760 & n10764;
  assign n10766 = pi39 & ~n10765;
  assign n10767 = ~n10696 & ~n10766;
  assign n10768 = n3206 & ~n10767;
  assign n10769 = ~pi299 & ~n10763;
  assign n10770 = n10487 & n10758;
  assign n10771 = pi232 & ~n10770;
  assign n10772 = n10769 & ~n10771;
  assign n10773 = pi39 & ~n10772;
  assign n10774 = ~n10618 & n10773;
  assign n10775 = ~n10715 & ~n10774;
  assign n10776 = n6235 & ~n10775;
  assign n10777 = ~n10719 & ~n10774;
  assign n10778 = pi38 & ~n10777;
  assign n10779 = ~pi87 & ~n10778;
  assign n10780 = ~n10776 & n10779;
  assign n10781 = ~n10768 & n10780;
  assign n10782 = n10735 & ~n10774;
  assign n10783 = ~pi75 & ~n10782;
  assign n10784 = ~n10781 & n10783;
  assign n10785 = ~n10750 & ~n10774;
  assign n10786 = pi75 & ~n10785;
  assign n10787 = n7422 & ~n10786;
  assign n10788 = ~n10784 & n10787;
  assign n10789 = ~n7422 & n10777;
  assign n10790 = n10564 & ~n10789;
  assign n10791 = ~n10788 & n10790;
  assign n10792 = ~n10757 & ~n10791;
  assign n10793 = n10673 & ~n10792;
  assign n10794 = pi232 & ~n10579;
  assign n10795 = n10570 & ~n10794;
  assign n10796 = pi39 & ~n10795;
  assign n10797 = ~n10696 & ~n10796;
  assign n10798 = n3206 & ~n10797;
  assign n10799 = ~n10574 & ~n10715;
  assign n10800 = n6235 & ~n10799;
  assign n10801 = ~n10574 & ~n10719;
  assign n10802 = pi38 & ~n10801;
  assign n10803 = ~pi87 & ~n10802;
  assign n10804 = ~n10800 & n10803;
  assign n10805 = ~n10798 & n10804;
  assign n10806 = ~n10574 & n10735;
  assign n10807 = ~pi75 & ~n10806;
  assign n10808 = ~n10805 & n10807;
  assign n10809 = ~n10574 & ~n10750;
  assign n10810 = pi75 & ~n10809;
  assign n10811 = n7422 & ~n10810;
  assign n10812 = ~n10808 & n10811;
  assign n10813 = ~n7422 & n10801;
  assign n10814 = ~n10564 & ~n10813;
  assign n10815 = ~n10812 & n10814;
  assign n10816 = pi232 & ~n10759;
  assign n10817 = n10769 & ~n10816;
  assign n10818 = pi39 & ~n10817;
  assign n10819 = ~n10696 & ~n10818;
  assign n10820 = n3206 & ~n10819;
  assign n10821 = ~n10715 & ~n10773;
  assign n10822 = n6235 & ~n10821;
  assign n10823 = ~n10719 & ~n10773;
  assign n10824 = pi38 & ~n10823;
  assign n10825 = ~pi87 & ~n10824;
  assign n10826 = ~n10822 & n10825;
  assign n10827 = ~n10820 & n10826;
  assign n10828 = ~n3276 & ~n10823;
  assign n10829 = n10735 & ~n10828;
  assign n10830 = ~pi75 & ~n10829;
  assign n10831 = ~n10827 & n10830;
  assign n10832 = ~n10750 & ~n10773;
  assign n10833 = pi75 & ~n10832;
  assign n10834 = n7422 & ~n10833;
  assign n10835 = ~n10831 & n10834;
  assign n10836 = ~n7422 & n10823;
  assign n10837 = n10564 & ~n10836;
  assign n10838 = ~n10835 & n10837;
  assign n10839 = ~n10815 & ~n10838;
  assign n10840 = ~n10673 & ~n10839;
  assign n10841 = ~po1038 & ~n10840;
  assign n10842 = ~n10793 & n10841;
  assign n10843 = n10606 & n10673;
  assign n10844 = pi39 & ~n10843;
  assign n10845 = po1038 & ~n10719;
  assign n10846 = ~n10844 & n10845;
  assign po201 = n10842 | n10846;
  assign n10848 = ~n8064 & ~n10316;
  assign n10849 = ~pi39 & ~n10848;
  assign n10850 = ~n2734 & n10316;
  assign n10851 = n8064 & ~n10850;
  assign n10852 = pi44 & pi72;
  assign n10853 = n7467 & ~n10852;
  assign n10854 = n7525 & n10244;
  assign n10855 = n7465 & n10854;
  assign n10856 = pi44 & ~n10257;
  assign n10857 = ~n10855 & ~n10856;
  assign n10858 = n10853 & ~n10857;
  assign n10859 = n10851 & ~n10858;
  assign n10860 = n10849 & ~n10859;
  assign n10861 = pi39 & n7463;
  assign n10862 = ~pi72 & n10861;
  assign n10863 = ~n10860 & ~n10862;
  assign n10864 = n3241 & ~n10863;
  assign n10865 = ~pi39 & ~n10316;
  assign n10866 = pi39 & ~n10862;
  assign n10867 = ~n10865 & ~n10866;
  assign n10868 = ~n3241 & n10867;
  assign n10869 = pi75 & ~n10868;
  assign n10870 = ~n10864 & n10869;
  assign n10871 = pi44 & n10315;
  assign n10872 = n2734 & ~n10304;
  assign n10873 = ~n10871 & n10872;
  assign n10874 = pi44 & n10326;
  assign n10875 = ~n2734 & ~n10323;
  assign n10876 = ~n10874 & n10875;
  assign n10877 = ~n10873 & ~n10876;
  assign n10878 = pi228 & ~n10877;
  assign n10879 = pi44 & n10368;
  assign n10880 = ~pi228 & ~n10879;
  assign n10881 = ~n10362 & n10880;
  assign n10882 = ~pi39 & ~n10881;
  assign n10883 = ~n10878 & n10882;
  assign n10884 = pi287 & n10382;
  assign n10885 = ~pi72 & ~n10884;
  assign n10886 = n10861 & n10885;
  assign n10887 = n3206 & ~n10886;
  assign n10888 = ~n10883 & n10887;
  assign n10889 = n7525 & n10382;
  assign n10890 = pi44 & ~n10889;
  assign n10891 = ~n10854 & ~n10890;
  assign n10892 = n10853 & ~n10891;
  assign n10893 = n10851 & ~n10892;
  assign n10894 = n10849 & ~n10893;
  assign n10895 = n6235 & ~n10862;
  assign n10896 = ~n10894 & n10895;
  assign n10897 = pi38 & ~n10867;
  assign n10898 = ~pi87 & ~n10897;
  assign n10899 = ~n10896 & n10898;
  assign n10900 = ~n10888 & n10899;
  assign n10901 = pi228 & n3206;
  assign n10902 = n10244 & n10901;
  assign n10903 = n10382 & n10901;
  assign n10904 = n10316 & ~n10903;
  assign n10905 = ~pi39 & ~n10904;
  assign n10906 = ~n10902 & n10905;
  assign n10907 = pi87 & ~n10866;
  assign n10908 = ~n10906 & n10907;
  assign n10909 = ~pi75 & ~n10908;
  assign n10910 = ~n10900 & n10909;
  assign n10911 = ~n10870 & ~n10910;
  assign n10912 = n7422 & ~n10911;
  assign n10913 = ~n7422 & ~n10867;
  assign n10914 = ~po1038 & ~n10913;
  assign n10915 = ~n10912 & n10914;
  assign n10916 = n2448 & n7462;
  assign n10917 = ~pi72 & n10916;
  assign n10918 = pi39 & ~n10917;
  assign n10919 = po1038 & ~n10865;
  assign n10920 = ~n10918 & n10919;
  assign po202 = n10915 | n10920;
  assign n10922 = ~pi38 & pi39;
  assign n10923 = n10143 & n10922;
  assign n10924 = pi979 & n10923;
  assign po203 = n6435 & n10924;
  assign n10926 = ~pi49 & ~pi76;
  assign n10927 = n8871 & n10926;
  assign n10928 = ~pi102 & ~pi104;
  assign n10929 = ~pi111 & n10928;
  assign n10930 = n10123 & n10929;
  assign n10931 = n10927 & n10930;
  assign n10932 = pi61 & ~pi82;
  assign n10933 = ~pi83 & ~pi89;
  assign n10934 = n10932 & n10933;
  assign n10935 = n7429 & n8885;
  assign n10936 = n10934 & n10935;
  assign n10937 = n8883 & n10936;
  assign n10938 = n10188 & n10937;
  assign n10939 = n10931 & n10938;
  assign n10940 = n8892 & n10939;
  assign n10941 = ~pi841 & n10940;
  assign n10942 = n2491 & n2698;
  assign n10943 = pi24 & n10942;
  assign n10944 = ~n10941 & ~n10943;
  assign po204 = n10112 & ~n10944;
  assign n10946 = ~n2680 & n7429;
  assign n10947 = ~pi82 & n2463;
  assign n10948 = ~pi84 & pi104;
  assign n10949 = n2607 & n10948;
  assign n10950 = n10127 & n10949;
  assign n10951 = n10947 & n10950;
  assign n10952 = ~pi36 & ~n10951;
  assign n10953 = n8884 & n8998;
  assign n10954 = ~pi67 & ~pi103;
  assign n10955 = n2476 & n10954;
  assign n10956 = ~pi98 & n10955;
  assign n10957 = n10953 & n10956;
  assign n10958 = ~n10952 & n10957;
  assign n10959 = ~n2648 & n10958;
  assign n10960 = ~pi88 & ~n10959;
  assign n10961 = n2532 & ~n10960;
  assign n10962 = n10946 & n10961;
  assign n10963 = n2489 & n10962;
  assign n10964 = ~n10105 & ~n10963;
  assign n10965 = n10108 & ~n10964;
  assign n10966 = n7538 & ~n10965;
  assign n10967 = ~n6257 & n10965;
  assign n10968 = ~pi36 & n10958;
  assign n10969 = ~pi88 & ~n10968;
  assign n10970 = n10946 & ~n10969;
  assign n10971 = n10122 & n10970;
  assign n10972 = ~pi824 & n6257;
  assign n10973 = n10971 & n10972;
  assign n10974 = pi829 & ~n10973;
  assign n10975 = ~n10967 & n10974;
  assign n10976 = ~n2733 & n10975;
  assign n10977 = ~n10966 & ~n10976;
  assign n10978 = pi1091 & ~n10977;
  assign n10979 = ~n7474 & n10965;
  assign n10980 = ~pi829 & ~n10979;
  assign n10981 = ~n10975 & ~n10980;
  assign n10982 = ~pi1093 & ~n10981;
  assign n10983 = n7474 & n10108;
  assign n10984 = ~n10106 & n10983;
  assign n10985 = ~n6449 & ~n7536;
  assign n10986 = ~n10984 & ~n10985;
  assign n10987 = ~n10979 & n10986;
  assign n10988 = n10111 & ~n10987;
  assign n10989 = ~n10982 & n10988;
  assign po205 = ~n10978 & n10989;
  assign n10991 = ~pi72 & pi841;
  assign n10992 = n2494 & n10991;
  assign n10993 = ~pi51 & n10992;
  assign n10994 = n10195 & n10993;
  assign n10995 = n10111 & n10994;
  assign po206 = n10121 & n10995;
  assign n10997 = pi74 & ~n8921;
  assign n10998 = ~pi103 & n2641;
  assign n10999 = n10186 & n10998;
  assign n11000 = n8871 & n8884;
  assign n11001 = n10999 & n11000;
  assign n11002 = n2453 & n2476;
  assign n11003 = ~pi45 & pi49;
  assign n11004 = n10929 & n11003;
  assign n11005 = n11002 & n11004;
  assign n11006 = n11001 & n11005;
  assign n11007 = n10947 & n11006;
  assign n11008 = n2495 & n8892;
  assign n11009 = n11007 & n11008;
  assign n11010 = n10107 & n10992;
  assign n11011 = n11009 & n11010;
  assign n11012 = ~pi74 & ~n11011;
  assign n11013 = n7357 & ~po1038;
  assign n11014 = ~n11012 & n11013;
  assign po207 = ~n10997 & n11014;
  assign n11016 = pi24 & n8859;
  assign n11017 = ~n10344 & ~n11016;
  assign n11018 = pi24 & ~pi94;
  assign n11019 = ~n8857 & n11018;
  assign n11020 = ~pi252 & ~n8848;
  assign n11021 = pi252 & ~po840;
  assign n11022 = ~n11020 & ~n11021;
  assign n11023 = n10108 & n11022;
  assign n11024 = ~n11019 & n11023;
  assign n11025 = ~n11017 & n11024;
  assign n11026 = n2535 & n7442;
  assign n11027 = pi24 & ~pi90;
  assign n11028 = n11026 & n11027;
  assign n11029 = ~n11022 & n11028;
  assign n11030 = n8861 & n11029;
  assign n11031 = ~n11025 & ~n11030;
  assign n11032 = ~pi100 & ~n11031;
  assign n11033 = pi100 & n6243;
  assign n11034 = n6486 & n11033;
  assign n11035 = ~n11032 & ~n11034;
  assign n11036 = n3181 & n3230;
  assign n11037 = ~n11035 & n11036;
  assign n11038 = n6263 & n8926;
  assign n11039 = n8922 & n11038;
  assign n11040 = ~n11037 & ~n11039;
  assign po208 = n8841 & ~n11040;
  assign n11042 = n2489 & n10112;
  assign n11043 = n2532 & n11042;
  assign n11044 = n8999 & n11002;
  assign n11045 = n2456 & n11044;
  assign n11046 = ~pi69 & n11045;
  assign n11047 = n2641 & n11046;
  assign n11048 = n2643 & n11047;
  assign po209 = n11043 & n11048;
  assign n11050 = ~pi219 & n10672;
  assign n11051 = pi52 & ~pi72;
  assign n11052 = ~pi39 & n11051;
  assign n11053 = pi38 & ~n11052;
  assign n11054 = n6247 & n6250;
  assign n11055 = pi228 & n11054;
  assign n11056 = ~pi52 & n10502;
  assign n11057 = pi52 & n10509;
  assign n11058 = ~n11056 & ~n11057;
  assign n11059 = n11055 & ~n11058;
  assign n11060 = n11051 & ~n11055;
  assign n11061 = ~n11059 & ~n11060;
  assign n11062 = ~pi38 & n11061;
  assign n11063 = ~n11053 & ~n11062;
  assign n11064 = ~pi100 & ~n11063;
  assign n11065 = pi100 & ~n11052;
  assign n11066 = ~pi100 & n10922;
  assign n11067 = pi87 & ~n11066;
  assign n11068 = ~n11065 & n11067;
  assign n11069 = ~n11064 & n11068;
  assign n11070 = ~pi114 & n6247;
  assign n11071 = pi52 & ~n10439;
  assign n11072 = ~pi52 & n10444;
  assign n11073 = n10429 & ~n11072;
  assign n11074 = ~n11071 & n11073;
  assign n11075 = pi52 & ~n10454;
  assign n11076 = ~pi52 & n10457;
  assign n11077 = n10449 & ~n11076;
  assign n11078 = ~n11075 & n11077;
  assign n11079 = ~n11074 & ~n11078;
  assign n11080 = n11070 & ~n11079;
  assign n11081 = ~n11051 & ~n11054;
  assign n11082 = pi228 & ~n11081;
  assign n11083 = ~n11080 & n11082;
  assign n11084 = pi52 & ~n10471;
  assign n11085 = ~pi52 & n10475;
  assign n11086 = n11054 & ~n11085;
  assign n11087 = ~n11084 & n11086;
  assign n11088 = ~pi228 & ~n11081;
  assign n11089 = ~n11087 & n11088;
  assign n11090 = ~pi39 & ~n11089;
  assign n11091 = ~n11083 & n11090;
  assign n11092 = ~pi100 & n11091;
  assign n11093 = n8064 & n10429;
  assign n11094 = n11070 & n11093;
  assign n11095 = n7525 & n11094;
  assign n11096 = n10508 & n11095;
  assign n11097 = n11051 & ~n11096;
  assign n11098 = pi100 & ~n11097;
  assign n11099 = ~pi39 & ~n11098;
  assign n11100 = ~n11092 & n11099;
  assign n11101 = ~pi38 & ~n11100;
  assign n11102 = ~pi87 & ~n11053;
  assign n11103 = ~n11101 & n11102;
  assign n11104 = ~n11069 & ~n11103;
  assign n11105 = ~pi75 & ~n11104;
  assign n11106 = n10549 & n11094;
  assign n11107 = n3241 & n11106;
  assign n11108 = n11052 & ~n11107;
  assign n11109 = pi75 & n11108;
  assign n11110 = n7422 & ~n11109;
  assign n11111 = ~n11105 & n11110;
  assign n11112 = ~n7422 & ~n11052;
  assign n11113 = n10564 & ~n11112;
  assign n11114 = ~n11111 & n11113;
  assign n11115 = ~n10818 & ~n11091;
  assign n11116 = n3206 & ~n11115;
  assign n11117 = ~pi39 & ~n11097;
  assign n11118 = ~n10773 & ~n11117;
  assign n11119 = n6235 & ~n11118;
  assign n11120 = ~pi39 & ~n11051;
  assign n11121 = ~n10773 & ~n11120;
  assign n11122 = pi38 & ~n11121;
  assign n11123 = ~pi87 & ~n11122;
  assign n11124 = ~n11119 & n11123;
  assign n11125 = ~n11116 & n11124;
  assign n11126 = ~n3206 & n11121;
  assign n11127 = ~pi39 & n11061;
  assign n11128 = n3206 & ~n10773;
  assign n11129 = ~n11127 & n11128;
  assign n11130 = ~n11126 & ~n11129;
  assign n11131 = pi87 & ~n11130;
  assign n11132 = ~pi75 & ~n11131;
  assign n11133 = ~n11125 & n11132;
  assign n11134 = n11051 & ~n11106;
  assign n11135 = ~pi39 & ~n11134;
  assign n11136 = n3241 & ~n10773;
  assign n11137 = ~n11135 & n11136;
  assign n11138 = ~n3241 & n11121;
  assign n11139 = pi75 & ~n11138;
  assign n11140 = ~n11137 & n11139;
  assign n11141 = n7422 & ~n10564;
  assign n11142 = ~n11140 & n11141;
  assign n11143 = ~n11133 & n11142;
  assign n11144 = ~n11114 & ~n11143;
  assign n11145 = ~n11050 & ~n11144;
  assign n11146 = ~n10609 & n10611;
  assign n11147 = pi39 & ~n11146;
  assign n11148 = ~n11091 & ~n11147;
  assign n11149 = n3206 & ~n11148;
  assign n11150 = ~n10619 & ~n11120;
  assign n11151 = pi38 & ~n11150;
  assign n11152 = ~n10619 & ~n11117;
  assign n11153 = n6235 & ~n11152;
  assign n11154 = ~n11151 & ~n11153;
  assign n11155 = ~n11149 & n11154;
  assign n11156 = ~pi87 & ~n11155;
  assign n11157 = ~n3206 & n11150;
  assign n11158 = pi87 & ~n11157;
  assign n11159 = n3206 & ~n10619;
  assign n11160 = ~n11127 & n11159;
  assign n11161 = n11158 & ~n11160;
  assign n11162 = n10564 & ~n11161;
  assign n11163 = ~n11156 & n11162;
  assign n11164 = ~n10766 & ~n11091;
  assign n11165 = n3206 & ~n11164;
  assign n11166 = ~n10774 & ~n11117;
  assign n11167 = n6235 & ~n11166;
  assign n11168 = n11122 & ~n11150;
  assign n11169 = ~n11167 & ~n11168;
  assign n11170 = ~n11165 & n11169;
  assign n11171 = ~pi87 & ~n11170;
  assign n11172 = n3206 & ~n10774;
  assign n11173 = ~n11127 & n11172;
  assign n11174 = ~n11126 & n11158;
  assign n11175 = ~n11173 & n11174;
  assign n11176 = ~n10564 & ~n11175;
  assign n11177 = ~n11171 & n11176;
  assign n11178 = ~n11163 & ~n11177;
  assign n11179 = ~pi75 & ~n11178;
  assign n11180 = ~pi39 & ~n11108;
  assign n11181 = ~n10564 & n10774;
  assign n11182 = n10564 & n10619;
  assign n11183 = pi75 & ~n11182;
  assign n11184 = ~n11181 & n11183;
  assign n11185 = ~n11180 & n11184;
  assign n11186 = n7422 & ~n11185;
  assign n11187 = ~n11179 & n11186;
  assign n11188 = ~n7422 & ~n11150;
  assign n11189 = n11050 & ~n11188;
  assign n11190 = ~n11187 & n11189;
  assign n11191 = ~n7422 & ~n10564;
  assign n11192 = n11121 & n11191;
  assign n11193 = ~po1038 & ~n11192;
  assign n11194 = ~n11190 & n11193;
  assign n11195 = ~n11145 & n11194;
  assign n11196 = pi39 & n11050;
  assign n11197 = n10606 & n11196;
  assign n11198 = po1038 & ~n11052;
  assign n11199 = ~n11197 & n11198;
  assign po210 = ~n11195 & ~n11199;
  assign n11201 = pi24 & n10108;
  assign n11202 = pi53 & n2505;
  assign n11203 = n2514 & n11202;
  assign n11204 = n2506 & n11203;
  assign n11205 = n11201 & n11204;
  assign n11206 = ~pi39 & ~n11205;
  assign n11207 = ~pi287 & ~pi979;
  assign n11208 = n6163 & n11207;
  assign n11209 = pi39 & ~n11208;
  assign n11210 = n10146 & ~n11209;
  assign n11211 = ~n11206 & n11210;
  assign po211 = ~n3350 & n11211;
  assign n11213 = n3242 & n10117;
  assign n11214 = pi54 & ~n11213;
  assign n11215 = n8859 & n9004;
  assign n11216 = ~pi60 & ~pi85;
  assign n11217 = pi106 & n11216;
  assign n11218 = n2468 & n8875;
  assign n11219 = n11217 & n11218;
  assign n11220 = n10927 & n11219;
  assign n11221 = n8888 & n10999;
  assign n11222 = n11220 & n11221;
  assign n11223 = n11002 & n11222;
  assign n11224 = n11215 & n11223;
  assign n11225 = ~pi841 & n2493;
  assign n11226 = n8919 & n11225;
  assign n11227 = n2495 & n3238;
  assign n11228 = n11226 & n11227;
  assign n11229 = n11224 & n11228;
  assign n11230 = ~pi54 & ~n11229;
  assign n11231 = n8840 & ~n11230;
  assign po212 = ~n11214 & n11231;
  assign n11233 = ~pi54 & n11213;
  assign n11234 = ~pi74 & n11233;
  assign n11235 = pi55 & ~n11234;
  assign n11236 = pi45 & n2468;
  assign n11237 = n2476 & n11236;
  assign n11238 = n11001 & n11237;
  assign n11239 = n2465 & n11238;
  assign n11240 = n6360 & n9269;
  assign n11241 = n2454 & n3268;
  assign n11242 = n11240 & n11241;
  assign n11243 = n11239 & n11242;
  assign n11244 = ~pi55 & ~n11243;
  assign n11245 = n8838 & ~n11244;
  assign po213 = ~n11235 & n11245;
  assign n11247 = pi56 & ~pi62;
  assign n11248 = pi55 & n10088;
  assign n11249 = ~n11247 & ~n11248;
  assign n11250 = n3092 & n3280;
  assign n11251 = n6146 & n11250;
  assign n11252 = pi56 & ~n11251;
  assign n11253 = n3429 & ~n11252;
  assign po214 = ~n11249 & n11253;
  assign n11255 = n6366 & n11250;
  assign n11256 = ~pi56 & pi62;
  assign n11257 = ~pi924 & n11256;
  assign n11258 = ~n11247 & ~n11257;
  assign n11259 = n11255 & ~n11258;
  assign n11260 = ~pi57 & ~n11259;
  assign n11261 = n6285 & n11234;
  assign n11262 = pi57 & ~n11261;
  assign n11263 = ~pi59 & ~n11262;
  assign po215 = ~n11260 & n11263;
  assign n11265 = ~pi93 & n11026;
  assign n11266 = n10111 & n11265;
  assign po216 = n7425 & n11266;
  assign n11268 = pi924 & n11256;
  assign n11269 = n11255 & n11268;
  assign n11270 = ~pi59 & ~n11269;
  assign n11271 = pi59 & ~n11261;
  assign n11272 = ~pi57 & ~n11271;
  assign po217 = ~n11270 & n11272;
  assign n11274 = pi39 & ~pi979;
  assign n11275 = ~n6163 & n11274;
  assign n11276 = n6164 & n11275;
  assign n11277 = n6435 & n11276;
  assign n11278 = ~pi39 & n11201;
  assign n11279 = n11215 & n11278;
  assign n11280 = n2503 & n11279;
  assign n11281 = ~n11277 & ~n11280;
  assign po218 = n10146 & ~n11281;
  assign n11283 = pi841 & n10940;
  assign n11284 = ~pi24 & n11215;
  assign n11285 = n2503 & n11284;
  assign n11286 = ~n11283 & ~n11285;
  assign po219 = n10112 & ~n11286;
  assign n11288 = n11251 & n11256;
  assign n11289 = ~pi57 & ~n11288;
  assign n11290 = pi57 & ~n10089;
  assign n11291 = ~pi59 & ~n11290;
  assign po220 = ~n11289 & n11291;
  assign n11293 = n2671 & n8892;
  assign n11294 = n9001 & n11293;
  assign n11295 = pi999 & n11294;
  assign n11296 = ~pi24 & n10942;
  assign n11297 = ~n11295 & ~n11296;
  assign po221 = n10112 & ~n11297;
  assign n11299 = ~pi64 & ~n2663;
  assign n11300 = n2454 & ~n11299;
  assign n11301 = n10119 & n11300;
  assign n11302 = pi841 & ~n11301;
  assign n11303 = n2662 & n9001;
  assign n11304 = ~pi841 & ~n11303;
  assign n11305 = n11043 & ~n11304;
  assign po222 = ~n11302 & n11305;
  assign n11307 = pi39 & n10164;
  assign n11308 = n10146 & n11307;
  assign n11309 = ~n10169 & n11308;
  assign po223 = ~n10162 & n11309;
  assign n11311 = ~pi199 & ~pi299;
  assign n11312 = pi314 & n2453;
  assign n11313 = n11240 & n11312;
  assign n11314 = pi81 & ~pi102;
  assign n11315 = n11313 & n11314;
  assign n11316 = n2478 & n11315;
  assign n11317 = n3268 & n11316;
  assign n11318 = ~n11311 & n11317;
  assign n11319 = pi219 & ~n11318;
  assign n11320 = n3206 & n3266;
  assign n11321 = pi199 & ~pi299;
  assign n11322 = n3221 & n11321;
  assign n11323 = n11320 & n11322;
  assign n11324 = n11316 & n11323;
  assign n11325 = ~pi219 & ~n11324;
  assign n11326 = ~po1038 & ~n11325;
  assign po224 = ~n11319 & n11326;
  assign n11328 = pi83 & ~pi103;
  assign n11329 = n11044 & n11328;
  assign n11330 = n10111 & n11329;
  assign n11331 = n11313 & n11330;
  assign po225 = n2473 & n11331;
  assign n11333 = ~n6200 & n6451;
  assign n11334 = n3324 & n5767;
  assign n11335 = n11333 & n11334;
  assign n11336 = ~n6221 & n6451;
  assign n11337 = n3306 & n3474;
  assign n11338 = n11336 & n11337;
  assign n11339 = ~n11335 & ~n11338;
  assign po226 = n10923 & ~n11339;
  assign n11341 = pi69 & n10998;
  assign n11342 = n10094 & n11341;
  assign n11343 = ~pi71 & ~n11342;
  assign n11344 = ~pi81 & ~pi314;
  assign n11345 = n2454 & n11344;
  assign n11346 = n6317 & n11345;
  assign n11347 = ~n11343 & n11346;
  assign n11348 = n10097 & n11312;
  assign n11349 = ~n11044 & n11348;
  assign n11350 = n2474 & n11349;
  assign n11351 = ~n11347 & ~n11350;
  assign po227 = n11043 & ~n11351;
  assign n11353 = n2548 & n2560;
  assign n11354 = ~pi96 & n11353;
  assign n11355 = n10116 & n11354;
  assign n11356 = pi198 & pi589;
  assign n11357 = n3475 & ~n6221;
  assign n11358 = n11356 & n11357;
  assign n11359 = pi210 & pi589;
  assign n11360 = ~pi221 & n5767;
  assign n11361 = ~pi216 & n11360;
  assign n11362 = ~n6200 & n11361;
  assign n11363 = n11359 & n11362;
  assign n11364 = ~n11358 & ~n11363;
  assign n11365 = ~pi593 & n6436;
  assign n11366 = ~n6444 & n11365;
  assign n11367 = ~n11364 & n11366;
  assign n11368 = ~pi287 & ~n11367;
  assign n11369 = pi39 & ~n11368;
  assign n11370 = n3095 & n11369;
  assign n11371 = ~n11355 & ~n11370;
  assign po228 = n10146 & ~n11371;
  assign n11373 = ~pi50 & n8892;
  assign n11374 = n6323 & n11373;
  assign n11375 = n2458 & n2470;
  assign n11376 = n6302 & n11375;
  assign n11377 = n10955 & n11376;
  assign n11378 = ~pi64 & n8884;
  assign n11379 = n11377 & n11378;
  assign n11380 = ~pi81 & ~n11379;
  assign n11381 = ~pi199 & pi200;
  assign n11382 = ~pi299 & n11381;
  assign n11383 = pi211 & ~pi219;
  assign n11384 = pi299 & n11383;
  assign n11385 = ~n11382 & ~n11384;
  assign n11386 = pi314 & ~n11385;
  assign n11387 = n10108 & n11386;
  assign n11388 = ~n11380 & n11387;
  assign n11389 = n11374 & n11388;
  assign n11390 = n10953 & n11385;
  assign n11391 = n11313 & n11390;
  assign n11392 = n11377 & n11391;
  assign n11393 = ~n11389 & ~n11392;
  assign po229 = n10111 & ~n11393;
  assign n11395 = pi24 & n2498;
  assign n11396 = pi72 & n11395;
  assign n11397 = pi88 & n10093;
  assign n11398 = n6443 & n9127;
  assign n11399 = n11397 & n11398;
  assign n11400 = n2679 & n11399;
  assign n11401 = ~n11396 & ~n11400;
  assign n11402 = n6360 & ~n11401;
  assign n11403 = ~pi39 & ~n11402;
  assign n11404 = n7511 & n11336;
  assign n11405 = n7514 & n11333;
  assign n11406 = pi39 & ~n11405;
  assign n11407 = ~n11404 & n11406;
  assign n11408 = n10146 & ~n11407;
  assign po230 = ~n11403 & n11408;
  assign n11410 = n9017 & n11336;
  assign n11411 = ~pi299 & ~n11410;
  assign n11412 = n9028 & n11333;
  assign n11413 = pi299 & ~n11412;
  assign n11414 = ~n11411 & ~n11413;
  assign n11415 = pi39 & ~n11414;
  assign n11416 = ~pi314 & pi1050;
  assign n11417 = n9525 & n10108;
  assign n11418 = n11416 & n11417;
  assign n11419 = ~pi39 & ~n11418;
  assign n11420 = n10146 & ~n11419;
  assign po231 = ~n11415 & n11420;
  assign n11422 = pi74 & n11233;
  assign n11423 = n2538 & n7483;
  assign n11424 = ~pi96 & ~n11423;
  assign n11425 = ~pi96 & ~pi1093;
  assign n11426 = n7474 & n11425;
  assign n11427 = n3406 & n7422;
  assign n11428 = ~n11426 & n11427;
  assign n11429 = ~pi96 & ~n6143;
  assign n11430 = pi479 & ~n11429;
  assign n11431 = ~po840 & ~n11430;
  assign n11432 = n11428 & n11431;
  assign n11433 = ~n11424 & n11432;
  assign n11434 = n7447 & n11433;
  assign n11435 = ~n11422 & ~n11434;
  assign po232 = ~po1038 & ~n11435;
  assign n11437 = pi96 & ~pi1093;
  assign n11438 = ~n2733 & n10018;
  assign n11439 = ~n11424 & n11438;
  assign n11440 = ~n11437 & ~n11439;
  assign n11441 = n3222 & ~n11440;
  assign n11442 = n7492 & n11441;
  assign n11443 = ~pi75 & ~n11442;
  assign n11444 = n3241 & n10117;
  assign n11445 = pi75 & ~n11444;
  assign n11446 = n8841 & ~n11445;
  assign po233 = ~n11443 & n11446;
  assign n11448 = n3093 & n10345;
  assign n11449 = pi252 & n7491;
  assign n11450 = n11448 & ~n11449;
  assign n11451 = ~pi137 & n11450;
  assign n11452 = ~pi137 & n2734;
  assign n11453 = ~n8859 & ~n10344;
  assign n11454 = ~pi94 & ~n8895;
  assign n11455 = n10108 & ~n11454;
  assign n11456 = ~n11453 & n11455;
  assign n11457 = ~n7491 & ~n11456;
  assign n11458 = ~pi252 & n11456;
  assign n11459 = n8890 & n10122;
  assign n11460 = pi252 & n11459;
  assign n11461 = n7491 & ~n11460;
  assign n11462 = ~n11458 & n11461;
  assign n11463 = ~n11457 & ~n11462;
  assign n11464 = pi122 & ~n11463;
  assign n11465 = n7474 & n11457;
  assign n11466 = ~n6258 & ~n11448;
  assign n11467 = ~n11462 & ~n11466;
  assign n11468 = ~n11465 & n11467;
  assign n11469 = ~pi122 & ~n11468;
  assign n11470 = ~n11464 & ~n11469;
  assign n11471 = ~pi1093 & ~n11470;
  assign n11472 = ~pi122 & ~n11450;
  assign n11473 = ~n11464 & ~n11472;
  assign n11474 = pi1093 & ~n11473;
  assign n11475 = ~n11471 & ~n11474;
  assign n11476 = n2734 & ~n11475;
  assign n11477 = ~n11452 & ~n11476;
  assign n11478 = ~n11451 & ~n11477;
  assign n11479 = ~pi122 & n11448;
  assign n11480 = pi1093 & ~n11456;
  assign n11481 = ~n8015 & ~n11480;
  assign n11482 = ~n11479 & ~n11481;
  assign n11483 = ~n11471 & ~n11482;
  assign n11484 = ~n2734 & ~n11483;
  assign n11485 = ~pi137 & ~n2734;
  assign n11486 = ~n11484 & ~n11485;
  assign n11487 = pi252 & pi1092;
  assign n11488 = ~pi1093 & n11487;
  assign n11489 = n2753 & n11488;
  assign n11490 = ~pi137 & ~n11489;
  assign n11491 = n11448 & n11490;
  assign n11492 = ~n11486 & ~n11491;
  assign n11493 = ~n11478 & ~n11492;
  assign n11494 = ~po1057 & ~n11493;
  assign n11495 = ~n10054 & n11459;
  assign n11496 = po1057 & ~n11495;
  assign n11497 = ~pi137 & po1057;
  assign n11498 = ~n11496 & ~n11497;
  assign n11499 = ~n11494 & n11498;
  assign n11500 = ~pi210 & ~n11499;
  assign n11501 = ~n11476 & ~n11484;
  assign n11502 = ~po1057 & ~n11501;
  assign n11503 = ~n11496 & ~n11502;
  assign n11504 = pi210 & ~n11503;
  assign n11505 = ~n11500 & ~n11504;
  assign n11506 = n2447 & n10266;
  assign n11507 = ~n11505 & ~n11506;
  assign n11508 = ~pi210 & ~n11493;
  assign n11509 = pi210 & ~n11501;
  assign n11510 = ~n11508 & ~n11509;
  assign n11511 = n11506 & ~n11510;
  assign n11512 = pi299 & ~n11511;
  assign n11513 = ~n11507 & n11512;
  assign n11514 = ~pi198 & ~n11499;
  assign n11515 = pi198 & ~n11503;
  assign n11516 = ~n11514 & ~n11515;
  assign n11517 = n3063 & n6162;
  assign n11518 = ~n11516 & ~n11517;
  assign n11519 = pi198 & ~n11501;
  assign n11520 = ~pi198 & ~n11493;
  assign n11521 = ~n11519 & ~n11520;
  assign n11522 = n11517 & ~n11521;
  assign n11523 = ~pi299 & ~n11522;
  assign n11524 = ~n11518 & n11523;
  assign n11525 = ~n11513 & ~n11524;
  assign n11526 = pi232 & ~n11525;
  assign n11527 = ~pi299 & ~n11516;
  assign n11528 = pi299 & ~n11505;
  assign n11529 = ~pi232 & ~n11528;
  assign n11530 = ~n11527 & n11529;
  assign n11531 = ~n11526 & ~n11530;
  assign n11532 = n7697 & ~n11531;
  assign n11533 = n7491 & ~n11448;
  assign n11534 = ~n11449 & ~n11457;
  assign n11535 = ~n11533 & n11534;
  assign n11536 = n8015 & ~n11535;
  assign n11537 = ~n11464 & ~n11536;
  assign n11538 = n2734 & ~n11537;
  assign n11539 = ~n2734 & n11480;
  assign n11540 = ~pi1093 & ~n11463;
  assign n11541 = ~n11539 & ~n11540;
  assign n11542 = ~n11538 & n11541;
  assign n11543 = ~po1057 & n11542;
  assign n11544 = po1057 & n11459;
  assign n11545 = ~n10050 & n11544;
  assign n11546 = ~n11543 & ~n11545;
  assign n11547 = pi210 & ~n11546;
  assign n11548 = ~pi137 & ~n11535;
  assign n11549 = pi137 & n11540;
  assign n11550 = ~n11548 & ~n11549;
  assign n11551 = ~pi1093 & ~n11550;
  assign n11552 = ~n11480 & ~n11551;
  assign n11553 = ~po1057 & n11552;
  assign n11554 = ~n11544 & ~n11553;
  assign n11555 = n8864 & n11497;
  assign n11556 = ~n2734 & ~n11555;
  assign n11557 = ~n11554 & n11556;
  assign n11558 = pi137 & ~n11537;
  assign n11559 = n11550 & ~n11558;
  assign n11560 = ~po1057 & ~n11559;
  assign n11561 = pi137 & ~n8015;
  assign n11562 = n7491 & ~n11561;
  assign n11563 = n11459 & ~n11562;
  assign n11564 = po1057 & ~n11563;
  assign n11565 = n2734 & ~n11564;
  assign n11566 = ~n11560 & n11565;
  assign n11567 = ~n11557 & ~n11566;
  assign n11568 = ~pi210 & ~n11567;
  assign n11569 = ~n11547 & ~n11568;
  assign n11570 = ~n11506 & ~n11569;
  assign n11571 = ~n6173 & ~n11559;
  assign n11572 = ~n11539 & ~n11571;
  assign n11573 = ~pi210 & ~n11572;
  assign n11574 = pi210 & ~n11542;
  assign n11575 = n11506 & ~n11574;
  assign n11576 = ~n11573 & n11575;
  assign n11577 = pi299 & ~n11576;
  assign n11578 = ~n11570 & n11577;
  assign n11579 = pi198 & ~n11546;
  assign n11580 = ~pi198 & ~n11567;
  assign n11581 = ~n11579 & ~n11580;
  assign n11582 = ~n11517 & ~n11581;
  assign n11583 = ~pi198 & n11572;
  assign n11584 = pi198 & n11542;
  assign n11585 = ~n11583 & ~n11584;
  assign n11586 = n11517 & ~n11585;
  assign n11587 = ~pi299 & ~n11586;
  assign n11588 = ~n11582 & n11587;
  assign n11589 = ~n11578 & ~n11588;
  assign n11590 = pi232 & ~n11589;
  assign n11591 = pi299 & ~n11569;
  assign n11592 = ~pi299 & ~n11581;
  assign n11593 = ~pi232 & ~n11592;
  assign n11594 = ~n11591 & n11593;
  assign n11595 = ~n7697 & ~n11594;
  assign n11596 = ~n11590 & n11595;
  assign n11597 = ~n11532 & ~n11596;
  assign po234 = n10111 & ~n11597;
  assign n11599 = n2578 & n2593;
  assign n11600 = ~pi86 & ~n11599;
  assign n11601 = n6331 & ~n11600;
  assign n11602 = n2491 & n11601;
  assign n11603 = ~pi314 & ~n11602;
  assign n11604 = pi86 & n8859;
  assign n11605 = n2587 & n11604;
  assign n11606 = pi314 & ~n11605;
  assign n11607 = n10112 & ~n11606;
  assign po235 = ~n11603 & n11607;
  assign n11609 = pi119 & pi232;
  assign po236 = ~pi468 & n11609;
  assign n11611 = pi163 & ~n9644;
  assign n11612 = ~pi163 & ~n9640;
  assign n11613 = ~n9642 & n11612;
  assign n11614 = ~n11611 & ~n11613;
  assign n11615 = pi232 & n11614;
  assign n11616 = pi75 & ~n11615;
  assign n11617 = pi100 & ~n11615;
  assign n11618 = ~n11616 & ~n11617;
  assign n11619 = pi147 & n7462;
  assign n11620 = n8948 & n11619;
  assign n11621 = n11618 & ~n11620;
  assign n11622 = ~n8948 & n11615;
  assign n11623 = pi74 & ~n11622;
  assign n11624 = ~n3429 & ~n11623;
  assign n11625 = n11621 & n11624;
  assign n11626 = pi299 & ~n11614;
  assign n11627 = ~n9673 & n9674;
  assign n11628 = pi184 & n6162;
  assign n11629 = ~n11627 & n11628;
  assign n11630 = ~pi184 & n11627;
  assign n11631 = ~pi299 & ~n11630;
  assign n11632 = ~n11629 & n11631;
  assign n11633 = pi232 & ~n11632;
  assign n11634 = ~n11626 & n11633;
  assign n11635 = ~n8948 & n11634;
  assign n11636 = pi74 & ~n11635;
  assign n11637 = ~pi55 & ~n11636;
  assign n11638 = ~pi187 & ~pi299;
  assign n11639 = ~pi147 & pi299;
  assign n11640 = ~n11638 & ~n11639;
  assign n11641 = n7462 & n11640;
  assign n11642 = n8948 & ~n11641;
  assign n11643 = pi54 & ~n11642;
  assign n11644 = ~n11635 & n11643;
  assign n11645 = ~pi187 & ~n8984;
  assign n11646 = pi187 & ~n8986;
  assign n11647 = pi147 & ~n11646;
  assign n11648 = ~n11645 & n11647;
  assign n11649 = ~pi147 & pi187;
  assign n11650 = n8991 & n11649;
  assign n11651 = ~n11648 & ~n11650;
  assign n11652 = pi38 & ~n11651;
  assign n11653 = ~pi40 & ~n9170;
  assign n11654 = ~pi95 & ~n11653;
  assign n11655 = ~pi40 & ~n9187;
  assign n11656 = pi166 & n11655;
  assign n11657 = n11654 & ~n11656;
  assign n11658 = n6162 & ~n9213;
  assign n11659 = ~n11657 & n11658;
  assign n11660 = ~pi153 & ~n11659;
  assign n11661 = ~pi40 & ~n9272;
  assign n11662 = ~pi95 & ~n11661;
  assign n11663 = pi166 & ~n11662;
  assign n11664 = n11658 & n11663;
  assign n11665 = n9212 & n10266;
  assign n11666 = pi153 & ~n11665;
  assign n11667 = ~n11664 & n11666;
  assign n11668 = pi160 & ~n11667;
  assign n11669 = ~n11660 & n11668;
  assign n11670 = ~pi153 & n11657;
  assign n11671 = ~n2449 & ~n9213;
  assign n11672 = n9072 & ~n9073;
  assign n11673 = ~n11671 & ~n11672;
  assign n11674 = ~n11417 & ~n11662;
  assign n11675 = pi153 & ~n11663;
  assign n11676 = ~n11674 & n11675;
  assign n11677 = ~pi160 & n6162;
  assign n11678 = ~n11676 & n11677;
  assign n11679 = ~n11673 & n11678;
  assign n11680 = ~n11670 & n11679;
  assign n11681 = pi163 & ~n11680;
  assign n11682 = ~n11669 & n11681;
  assign n11683 = ~pi40 & ~n9321;
  assign n11684 = ~pi95 & ~n11683;
  assign n11685 = ~n11673 & ~n11684;
  assign n11686 = pi166 & n11685;
  assign n11687 = ~pi40 & n9146;
  assign n11688 = ~pi32 & ~n11687;
  assign n11689 = ~n9231 & ~n11688;
  assign n11690 = ~pi95 & ~n11689;
  assign n11691 = ~n11673 & ~n11690;
  assign n11692 = ~pi210 & ~n11691;
  assign n11693 = ~n9214 & ~n11688;
  assign n11694 = ~pi95 & ~n11693;
  assign n11695 = ~n11673 & ~n11694;
  assign n11696 = pi210 & ~n11695;
  assign n11697 = n10266 & ~n11696;
  assign n11698 = ~n11692 & n11697;
  assign n11699 = ~pi153 & ~n11698;
  assign n11700 = ~n11686 & n11699;
  assign n11701 = ~n9227 & ~n11673;
  assign n11702 = pi210 & ~n11701;
  assign n11703 = ~n9233 & ~n11673;
  assign n11704 = ~pi210 & ~n11703;
  assign n11705 = n10266 & ~n11704;
  assign n11706 = ~n11702 & n11705;
  assign n11707 = ~n9261 & ~n11673;
  assign n11708 = ~pi210 & ~n11707;
  assign n11709 = pi166 & n6162;
  assign n11710 = ~pi95 & ~n9255;
  assign n11711 = ~n11673 & ~n11710;
  assign n11712 = pi210 & ~n11711;
  assign n11713 = n11709 & ~n11712;
  assign n11714 = ~n11708 & n11713;
  assign n11715 = pi153 & ~n11714;
  assign n11716 = ~n11706 & n11715;
  assign n11717 = ~pi160 & ~n11716;
  assign n11718 = ~n11700 & n11717;
  assign n11719 = n11683 & n11709;
  assign n11720 = ~n9213 & ~n11694;
  assign n11721 = pi210 & ~n11720;
  assign n11722 = ~n9213 & ~n11690;
  assign n11723 = ~pi210 & ~n11722;
  assign n11724 = n10266 & ~n11723;
  assign n11725 = ~n11721 & n11724;
  assign n11726 = ~pi153 & ~n11725;
  assign n11727 = ~n11719 & n11726;
  assign n11728 = ~n9213 & ~n11710;
  assign n11729 = pi210 & ~n11728;
  assign n11730 = ~pi210 & ~n9262;
  assign n11731 = n11709 & ~n11730;
  assign n11732 = ~n11729 & n11731;
  assign n11733 = ~pi210 & ~n9234;
  assign n11734 = pi210 & ~n9228;
  assign n11735 = n10266 & ~n11734;
  assign n11736 = ~n11733 & n11735;
  assign n11737 = pi153 & ~n11736;
  assign n11738 = ~n11732 & n11737;
  assign n11739 = pi160 & ~n11738;
  assign n11740 = ~n11727 & n11739;
  assign n11741 = ~pi163 & ~n11740;
  assign n11742 = ~n11718 & n11741;
  assign n11743 = ~n11682 & ~n11742;
  assign n11744 = ~n6162 & n11685;
  assign n11745 = pi299 & ~n11744;
  assign n11746 = ~n11743 & n11745;
  assign n11747 = ~pi40 & ~n9201;
  assign n11748 = ~pi95 & ~n11747;
  assign n11749 = ~n11673 & ~n11748;
  assign n11750 = ~n6162 & n11749;
  assign n11751 = ~pi175 & ~pi299;
  assign n11752 = pi189 & n11655;
  assign n11753 = n11654 & ~n11752;
  assign n11754 = ~pi182 & n11673;
  assign n11755 = pi182 & n9213;
  assign n11756 = n6162 & ~n11755;
  assign n11757 = ~n11754 & n11756;
  assign n11758 = ~n11753 & n11757;
  assign n11759 = pi184 & ~n11758;
  assign n11760 = pi189 & n6162;
  assign n11761 = n11747 & n11760;
  assign n11762 = pi198 & ~n11720;
  assign n11763 = ~pi198 & ~n11722;
  assign n11764 = n10270 & ~n11763;
  assign n11765 = ~n11762 & n11764;
  assign n11766 = pi182 & ~pi184;
  assign n11767 = ~n11765 & n11766;
  assign n11768 = ~n11761 & n11767;
  assign n11769 = ~n11759 & ~n11768;
  assign n11770 = n11751 & ~n11769;
  assign n11771 = pi198 & ~n11728;
  assign n11772 = ~pi198 & ~n9262;
  assign n11773 = n11760 & ~n11772;
  assign n11774 = ~n11771 & n11773;
  assign n11775 = n9236 & n10270;
  assign n11776 = pi182 & ~n11775;
  assign n11777 = ~n11774 & n11776;
  assign n11778 = pi198 & ~n11711;
  assign n11779 = ~pi198 & ~n11707;
  assign n11780 = n11760 & ~n11779;
  assign n11781 = ~n11778 & n11780;
  assign n11782 = ~pi182 & ~n11781;
  assign n11783 = ~n11777 & ~n11782;
  assign n11784 = pi95 & ~pi182;
  assign n11785 = ~n9236 & ~n11784;
  assign n11786 = n10270 & ~n11673;
  assign n11787 = ~n11785 & n11786;
  assign n11788 = ~n11783 & ~n11787;
  assign n11789 = ~pi184 & ~n11788;
  assign n11790 = pi175 & ~pi299;
  assign n11791 = ~pi95 & pi189;
  assign n11792 = n2476 & ~n11791;
  assign n11793 = n11661 & ~n11792;
  assign n11794 = ~n11784 & ~n11793;
  assign n11795 = n11628 & ~n11794;
  assign n11796 = ~n11754 & n11795;
  assign n11797 = n11790 & ~n11796;
  assign n11798 = ~n11789 & n11797;
  assign n11799 = ~n11770 & ~n11798;
  assign n11800 = ~n11750 & ~n11799;
  assign n11801 = ~n10270 & n11749;
  assign n11802 = ~pi182 & ~pi184;
  assign n11803 = n11751 & n11802;
  assign n11804 = ~pi95 & ~n11765;
  assign n11805 = n11786 & ~n11804;
  assign n11806 = n11803 & ~n11805;
  assign n11807 = ~n11801 & n11806;
  assign n11808 = ~n11800 & ~n11807;
  assign n11809 = ~n11746 & n11808;
  assign n11810 = pi232 & ~n11809;
  assign n11811 = pi299 & n11685;
  assign n11812 = ~pi299 & n11749;
  assign n11813 = ~pi232 & ~n11812;
  assign n11814 = ~n11811 & n11813;
  assign n11815 = ~pi39 & ~n11814;
  assign n11816 = ~n11810 & n11815;
  assign n11817 = ~n9017 & ~n9212;
  assign n11818 = ~pi40 & ~n9016;
  assign n11819 = ~pi189 & ~n11818;
  assign n11820 = n2476 & ~n9020;
  assign n11821 = n9199 & ~n11820;
  assign n11822 = n6192 & n9212;
  assign n11823 = n2476 & ~n9014;
  assign n11824 = ~pi40 & ~n11823;
  assign n11825 = n6198 & n11824;
  assign n11826 = ~n11822 & ~n11825;
  assign n11827 = ~n11821 & n11826;
  assign n11828 = pi189 & ~n6215;
  assign n11829 = n11827 & n11828;
  assign n11830 = ~n11819 & ~n11829;
  assign n11831 = pi179 & ~n11830;
  assign n11832 = n6215 & ~n11818;
  assign n11833 = n9031 & n9199;
  assign n11834 = ~n2476 & n9199;
  assign n11835 = ~n11833 & ~n11834;
  assign n11836 = n11826 & n11835;
  assign n11837 = ~pi189 & ~n11836;
  assign n11838 = ~n6192 & n11824;
  assign n11839 = ~n11822 & ~n11838;
  assign n11840 = pi189 & ~n11839;
  assign n11841 = ~pi179 & ~n6215;
  assign n11842 = ~n11840 & n11841;
  assign n11843 = ~n11837 & n11842;
  assign n11844 = ~n11832 & ~n11843;
  assign n11845 = ~n11831 & n11844;
  assign n11846 = n9017 & ~n11845;
  assign n11847 = ~n11817 & ~n11846;
  assign n11848 = ~pi299 & ~n11847;
  assign n11849 = ~n9028 & n9212;
  assign n11850 = pi299 & ~n11849;
  assign n11851 = pi166 & ~n6189;
  assign n11852 = n11827 & n11851;
  assign n11853 = ~n11818 & ~n11851;
  assign n11854 = n9028 & ~n11853;
  assign n11855 = ~n11852 & n11854;
  assign n11856 = n11850 & ~n11855;
  assign n11857 = ~n11848 & ~n11856;
  assign n11858 = pi156 & pi232;
  assign n11859 = ~n11857 & n11858;
  assign n11860 = n6189 & ~n11818;
  assign n11861 = ~n6189 & n11839;
  assign n11862 = ~n11860 & ~n11861;
  assign n11863 = ~pi166 & ~n6189;
  assign n11864 = ~n11862 & ~n11863;
  assign n11865 = n11836 & n11863;
  assign n11866 = n9028 & ~n11865;
  assign n11867 = ~n11864 & n11866;
  assign n11868 = n11850 & ~n11867;
  assign n11869 = ~n11848 & ~n11868;
  assign n11870 = ~pi156 & pi232;
  assign n11871 = ~n11869 & n11870;
  assign n11872 = ~n6215 & n11839;
  assign n11873 = ~n11832 & ~n11872;
  assign n11874 = n9017 & ~n11873;
  assign n11875 = ~pi299 & ~n11817;
  assign n11876 = ~n11874 & n11875;
  assign n11877 = n9030 & n11862;
  assign n11878 = ~pi232 & ~n11877;
  assign n11879 = ~n11876 & n11878;
  assign n11880 = pi39 & ~n11879;
  assign n11881 = ~n11871 & n11880;
  assign n11882 = ~n11859 & n11881;
  assign n11883 = ~pi38 & ~n11882;
  assign n11884 = ~n11816 & n11883;
  assign n11885 = ~n11652 & ~n11884;
  assign n11886 = n3240 & ~n11885;
  assign n11887 = pi100 & ~n11634;
  assign n11888 = pi38 & ~n11641;
  assign n11889 = ~pi100 & ~n11888;
  assign n11890 = ~pi38 & ~pi40;
  assign n11891 = pi87 & ~n2476;
  assign n11892 = n11890 & n11891;
  assign n11893 = n11889 & ~n11892;
  assign n11894 = pi87 & n11893;
  assign n11895 = ~n11887 & ~n11894;
  assign n11896 = ~n11886 & n11895;
  assign n11897 = n3237 & ~n11896;
  assign n11898 = pi75 & ~n11634;
  assign n11899 = pi39 & ~n9212;
  assign n11900 = n9597 & ~n11899;
  assign n11901 = n2476 & ~n9010;
  assign n11902 = ~pi40 & ~n11901;
  assign n11903 = ~pi179 & ~pi299;
  assign n11904 = ~pi156 & pi299;
  assign n11905 = ~n11903 & ~n11904;
  assign n11906 = n7462 & n11905;
  assign n11907 = n2476 & n11906;
  assign n11908 = n11902 & ~n11907;
  assign n11909 = ~pi39 & ~n11908;
  assign n11910 = n11900 & ~n11909;
  assign n11911 = n11893 & ~n11910;
  assign n11912 = ~n11887 & ~n11911;
  assign n11913 = n9410 & ~n11912;
  assign n11914 = ~n11898 & ~n11913;
  assign n11915 = ~n11897 & n11914;
  assign n11916 = ~pi54 & ~n11915;
  assign n11917 = ~n11644 & ~n11916;
  assign n11918 = ~pi74 & ~n11917;
  assign n11919 = n11637 & ~n11918;
  assign n11920 = pi55 & ~n11623;
  assign n11921 = pi54 & ~n11621;
  assign n11922 = pi163 & pi232;
  assign n11923 = ~n6162 & n9010;
  assign n11924 = n8997 & ~n11923;
  assign n11925 = n11922 & n11924;
  assign n11926 = n11902 & ~n11925;
  assign n11927 = ~pi39 & ~n11926;
  assign n11928 = n11900 & ~n11927;
  assign n11929 = pi38 & ~n11619;
  assign n11930 = ~pi100 & ~n11929;
  assign n11931 = ~n11892 & n11930;
  assign n11932 = ~n11928 & n11931;
  assign n11933 = ~n11617 & ~n11932;
  assign n11934 = n3237 & ~n11933;
  assign n11935 = ~n11890 & n11930;
  assign n11936 = ~n11617 & ~n11935;
  assign n11937 = ~n9405 & n11936;
  assign n11938 = n9410 & ~n11937;
  assign n11939 = ~n11616 & ~n11938;
  assign n11940 = ~n11934 & n11939;
  assign n11941 = ~pi54 & ~n11940;
  assign n11942 = ~n11921 & ~n11941;
  assign n11943 = ~pi74 & ~n11942;
  assign n11944 = n11920 & ~n11943;
  assign n11945 = n3293 & ~n11944;
  assign n11946 = ~n11919 & n11945;
  assign n11947 = ~pi75 & ~n11936;
  assign n11948 = ~n11616 & ~n11947;
  assign n11949 = ~pi54 & ~n11948;
  assign n11950 = ~n11921 & ~n11949;
  assign n11951 = ~pi74 & ~n11950;
  assign n11952 = ~n11623 & ~n11951;
  assign n11953 = ~n3293 & ~n11952;
  assign n11954 = n3429 & ~n11953;
  assign n11955 = ~n9467 & n11954;
  assign n11956 = ~n11946 & n11955;
  assign n11957 = ~n11625 & ~n11956;
  assign n11958 = ~pi79 & n11957;
  assign n11959 = ~pi32 & pi95;
  assign n11960 = ~pi479 & n11959;
  assign n11961 = n2552 & n11960;
  assign n11962 = ~pi40 & ~n11961;
  assign n11963 = n9565 & n11962;
  assign n11964 = n10266 & ~n11963;
  assign n11965 = n9568 & n11962;
  assign n11966 = n11709 & ~n11965;
  assign n11967 = ~pi153 & ~n11966;
  assign n11968 = ~n11964 & n11967;
  assign n11969 = ~pi210 & ~n9515;
  assign n11970 = ~n9513 & n11962;
  assign n11971 = ~n11969 & n11970;
  assign n11972 = n10266 & ~n11971;
  assign n11973 = pi153 & n9535;
  assign n11974 = n9568 & ~n11973;
  assign n11975 = n11709 & ~n11974;
  assign n11976 = ~n11966 & ~n11975;
  assign n11977 = ~n11967 & n11976;
  assign n11978 = ~n11972 & n11977;
  assign n11979 = ~n11968 & ~n11978;
  assign n11980 = pi40 & ~n6162;
  assign n11981 = pi163 & ~n11980;
  assign n11982 = ~n11979 & n11981;
  assign n11983 = pi160 & ~n11982;
  assign n11984 = pi153 & n9513;
  assign n11985 = n9565 & ~n11984;
  assign n11986 = n10266 & ~n11985;
  assign n11987 = ~pi40 & pi163;
  assign n11988 = ~n11975 & n11987;
  assign n11989 = ~n11986 & n11988;
  assign n11990 = pi153 & n9519;
  assign n11991 = n9524 & n11990;
  assign n11992 = n9552 & n10266;
  assign n11993 = ~pi40 & ~pi163;
  assign n11994 = ~n11992 & n11993;
  assign n11995 = ~n11991 & n11994;
  assign n11996 = ~pi160 & ~n11995;
  assign n11997 = ~n11989 & n11996;
  assign n11998 = ~n11983 & ~n11997;
  assign n11999 = n6162 & n11961;
  assign n12000 = n11995 & ~n11999;
  assign n12001 = pi299 & ~n12000;
  assign n12002 = ~n11998 & n12001;
  assign n12003 = pi184 & n9545;
  assign n12004 = ~pi184 & ~n9552;
  assign n12005 = ~pi189 & ~n12004;
  assign n12006 = ~n12003 & n12005;
  assign n12007 = pi182 & n11961;
  assign n12008 = pi184 & pi189;
  assign n12009 = ~n9548 & n12008;
  assign n12010 = ~n12007 & ~n12009;
  assign n12011 = ~n12006 & n12010;
  assign n12012 = n6162 & ~n12011;
  assign n12013 = ~pi40 & ~n12012;
  assign n12014 = n11751 & ~n12013;
  assign n12015 = ~pi189 & n9527;
  assign n12016 = pi189 & ~n9524;
  assign n12017 = n3092 & ~n12016;
  assign n12018 = ~n12015 & n12017;
  assign n12019 = ~n12007 & ~n12018;
  assign n12020 = n6162 & ~n12019;
  assign n12021 = ~pi184 & ~n12020;
  assign n12022 = ~n9517 & n10270;
  assign n12023 = pi189 & n9537;
  assign n12024 = ~pi182 & pi184;
  assign n12025 = ~n12023 & n12024;
  assign n12026 = ~n12022 & n12025;
  assign n12027 = ~n12021 & ~n12026;
  assign n12028 = ~pi40 & ~n12027;
  assign n12029 = ~n9516 & n11970;
  assign n12030 = n10270 & ~n12029;
  assign n12031 = n9536 & n11962;
  assign n12032 = n11760 & ~n12031;
  assign n12033 = pi182 & pi184;
  assign n12034 = ~n11980 & n12033;
  assign n12035 = ~n12032 & n12034;
  assign n12036 = ~n12030 & n12035;
  assign n12037 = n11790 & ~n12036;
  assign n12038 = ~n12028 & n12037;
  assign n12039 = ~n12014 & ~n12038;
  assign n12040 = ~n12002 & n12039;
  assign n12041 = ~pi39 & ~n12040;
  assign n12042 = n2552 & n9519;
  assign n12043 = ~pi189 & n9012;
  assign n12044 = pi179 & n6201;
  assign n12045 = ~n12043 & ~n12044;
  assign n12046 = ~n6215 & n9017;
  assign n12047 = ~n12045 & n12046;
  assign n12048 = n12042 & n12047;
  assign n12049 = ~pi40 & ~pi299;
  assign n12050 = ~n12048 & n12049;
  assign n12051 = ~n6189 & n9028;
  assign n12052 = pi156 & n6201;
  assign n12053 = ~pi166 & n9012;
  assign n12054 = ~n12052 & ~n12053;
  assign n12055 = n12051 & ~n12054;
  assign n12056 = n12042 & n12055;
  assign n12057 = ~pi40 & pi299;
  assign n12058 = ~n12056 & n12057;
  assign n12059 = pi39 & ~n12058;
  assign n12060 = ~n12050 & n12059;
  assign n12061 = pi232 & ~n12060;
  assign n12062 = ~n12041 & n12061;
  assign n12063 = ~pi40 & ~pi232;
  assign n12064 = ~pi38 & ~n12063;
  assign n12065 = ~n12062 & n12064;
  assign n12066 = ~n11652 & ~n12065;
  assign n12067 = n3240 & ~n12066;
  assign n12068 = pi87 & ~n11890;
  assign n12069 = n11889 & n12068;
  assign n12070 = ~n11887 & ~n12069;
  assign n12071 = ~n12067 & n12070;
  assign n12072 = n3237 & ~n12071;
  assign n12073 = n3092 & n3221;
  assign n12074 = n11906 & n12073;
  assign n12075 = n2552 & n12074;
  assign n12076 = n11890 & ~n12075;
  assign n12077 = n11889 & ~n12076;
  assign n12078 = ~n11887 & ~n12077;
  assign n12079 = n9410 & ~n12078;
  assign n12080 = ~n11898 & ~n12079;
  assign n12081 = ~n12072 & n12080;
  assign n12082 = ~pi54 & ~n12081;
  assign n12083 = ~n11644 & ~n12082;
  assign n12084 = ~pi74 & ~n12083;
  assign n12085 = n11637 & ~n12084;
  assign n12086 = ~pi92 & n3221;
  assign n12087 = n11922 & n12086;
  assign n12088 = n12042 & n12087;
  assign n12089 = n11890 & ~n12088;
  assign n12090 = ~pi75 & n11930;
  assign n12091 = ~n12089 & n12090;
  assign n12092 = n11618 & ~n12091;
  assign n12093 = ~pi54 & ~n12092;
  assign n12094 = ~n11921 & ~n12093;
  assign n12095 = ~pi74 & ~n12094;
  assign n12096 = n11920 & ~n12095;
  assign n12097 = n3293 & ~n12096;
  assign n12098 = ~n12085 & n12097;
  assign n12099 = n11954 & ~n12098;
  assign n12100 = ~n11625 & ~n12099;
  assign n12101 = pi79 & n12100;
  assign n12102 = ~pi34 & n10008;
  assign n12103 = ~n12101 & ~n12102;
  assign n12104 = ~n11958 & n12103;
  assign n12105 = ~pi79 & ~n8936;
  assign n12106 = n11957 & ~n12105;
  assign n12107 = n12100 & n12105;
  assign n12108 = n12102 & ~n12107;
  assign n12109 = ~n12106 & n12108;
  assign po237 = n12104 | n12109;
  assign n12111 = pi98 & pi1092;
  assign n12112 = pi1093 & n12111;
  assign n12113 = ~pi567 & n2754;
  assign n12114 = ~n12112 & ~n12113;
  assign n12115 = ~n8558 & n12114;
  assign n12116 = pi588 & ~n12115;
  assign n12117 = pi592 & ~n12114;
  assign n12118 = ~n7422 & n12114;
  assign n12119 = n7422 & ~n12113;
  assign n12120 = pi75 & n12112;
  assign n12121 = pi1091 & n12112;
  assign n12122 = ~pi110 & n2490;
  assign n12123 = ~pi88 & n2484;
  assign n12124 = n10334 & n12123;
  assign n12125 = n12122 & n12124;
  assign n12126 = n7431 & n12125;
  assign n12127 = n7438 & n12126;
  assign n12128 = pi51 & n12127;
  assign n12129 = pi90 & pi93;
  assign n12130 = ~pi841 & ~n2493;
  assign n12131 = ~n12129 & n12130;
  assign n12132 = n2535 & n12131;
  assign n12133 = n12126 & n12132;
  assign n12134 = ~n12128 & ~n12133;
  assign n12135 = pi824 & pi950;
  assign n12136 = n7442 & n12135;
  assign n12137 = ~n12134 & n12136;
  assign n12138 = ~pi98 & ~n12137;
  assign n12139 = pi1092 & ~n12138;
  assign n12140 = ~n12121 & ~n12139;
  assign n12141 = ~n7536 & ~n12121;
  assign n12142 = n3222 & ~n12141;
  assign n12143 = ~n12140 & n12142;
  assign n12144 = n3094 & n12135;
  assign n12145 = n12127 & n12144;
  assign n12146 = ~pi98 & ~n12145;
  assign n12147 = pi1092 & ~n12146;
  assign n12148 = ~n12121 & ~n12147;
  assign n12149 = n7578 & ~n12141;
  assign n12150 = ~n12148 & n12149;
  assign n12151 = ~n3207 & n12112;
  assign n12152 = ~n12150 & ~n12151;
  assign n12153 = ~n12143 & n12152;
  assign n12154 = ~pi75 & ~n12153;
  assign n12155 = ~n12120 & ~n12154;
  assign n12156 = pi567 & ~n12155;
  assign n12157 = n12119 & ~n12156;
  assign n12158 = ~n12118 & ~n12157;
  assign n12159 = ~pi592 & n12158;
  assign n12160 = ~n12117 & ~n12159;
  assign n12161 = ~n8480 & n12160;
  assign n12162 = ~pi1196 & ~n12114;
  assign n12163 = n8480 & ~n12162;
  assign n12164 = ~pi443 & ~n12114;
  assign n12165 = pi443 & ~n12160;
  assign n12166 = ~n12164 & ~n12165;
  assign n12167 = n8568 & n12166;
  assign n12168 = pi443 & ~n12114;
  assign n12169 = ~pi443 & ~n12160;
  assign n12170 = ~n12168 & ~n12169;
  assign n12171 = ~n8568 & n12170;
  assign n12172 = ~n12167 & ~n12171;
  assign n12173 = pi435 & ~n12172;
  assign n12174 = pi444 & n12166;
  assign n12175 = ~pi444 & n12170;
  assign n12176 = ~pi436 & ~n12175;
  assign n12177 = ~n12174 & n12176;
  assign n12178 = pi444 & n12170;
  assign n12179 = ~pi444 & n12166;
  assign n12180 = pi436 & ~n12179;
  assign n12181 = ~n12178 & n12180;
  assign n12182 = ~n12177 & ~n12181;
  assign n12183 = ~pi435 & n12182;
  assign n12184 = ~n12173 & ~n12183;
  assign n12185 = pi429 & n12184;
  assign n12186 = ~pi435 & ~n12172;
  assign n12187 = pi435 & n12182;
  assign n12188 = ~n12186 & ~n12187;
  assign n12189 = ~pi429 & n12188;
  assign n12190 = ~n8505 & ~n12189;
  assign n12191 = ~n12185 & n12190;
  assign n12192 = pi429 & n12188;
  assign n12193 = ~pi429 & n12184;
  assign n12194 = n8505 & ~n12193;
  assign n12195 = ~n12192 & n12194;
  assign n12196 = pi1196 & ~n12195;
  assign n12197 = ~n12191 & n12196;
  assign n12198 = n12163 & ~n12197;
  assign n12199 = ~n12161 & ~n12198;
  assign n12200 = ~pi428 & ~n12199;
  assign n12201 = pi428 & n12160;
  assign n12202 = ~n12200 & ~n12201;
  assign n12203 = ~pi427 & ~n12202;
  assign n12204 = pi428 & ~n12199;
  assign n12205 = ~pi428 & n12160;
  assign n12206 = ~n12204 & ~n12205;
  assign n12207 = pi427 & ~n12206;
  assign n12208 = ~n12203 & ~n12207;
  assign n12209 = pi430 & ~n12208;
  assign n12210 = ~pi427 & ~n12206;
  assign n12211 = pi427 & ~n12202;
  assign n12212 = ~n12210 & ~n12211;
  assign n12213 = ~pi430 & ~n12212;
  assign n12214 = ~n12209 & ~n12213;
  assign n12215 = pi426 & ~n12214;
  assign n12216 = pi430 & ~n12212;
  assign n12217 = ~pi430 & ~n12208;
  assign n12218 = ~n12216 & ~n12217;
  assign n12219 = ~pi426 & ~n12218;
  assign n12220 = ~n12215 & ~n12219;
  assign n12221 = pi445 & ~n12220;
  assign n12222 = pi426 & ~n12218;
  assign n12223 = ~pi426 & ~n12214;
  assign n12224 = ~n12222 & ~n12223;
  assign n12225 = ~pi445 & ~n12224;
  assign n12226 = ~n12221 & ~n12225;
  assign n12227 = ~pi448 & n12226;
  assign n12228 = pi445 & ~n12224;
  assign n12229 = ~pi445 & ~n12220;
  assign n12230 = ~n12228 & ~n12229;
  assign n12231 = pi448 & n12230;
  assign n12232 = ~n8426 & ~n12231;
  assign n12233 = ~n12227 & n12232;
  assign n12234 = ~pi448 & n12230;
  assign n12235 = pi448 & n12226;
  assign n12236 = n8426 & ~n12235;
  assign n12237 = ~n12234 & n12236;
  assign n12238 = pi1199 & ~n12237;
  assign n12239 = ~n12233 & n12238;
  assign n12240 = ~pi1199 & n12199;
  assign n12241 = n8558 & ~n12240;
  assign n12242 = ~n12239 & n12241;
  assign n12243 = n12116 & ~n12242;
  assign n12244 = pi591 & ~n12114;
  assign n12245 = pi590 & ~n12244;
  assign n12246 = n8657 & n12114;
  assign n12247 = ~n8657 & n12160;
  assign n12248 = ~n12246 & ~n12247;
  assign n12249 = pi1198 & ~n12248;
  assign n12250 = ~pi1198 & ~n12162;
  assign n12251 = n7591 & n12114;
  assign n12252 = ~n7591 & n12160;
  assign n12253 = ~n12251 & ~n12252;
  assign n12254 = pi355 & ~n12253;
  assign n12255 = pi455 & ~n12114;
  assign n12256 = ~pi455 & ~n12160;
  assign n12257 = ~n12255 & ~n12256;
  assign n12258 = ~pi452 & ~n12257;
  assign n12259 = ~pi455 & ~n12114;
  assign n12260 = pi455 & ~n12160;
  assign n12261 = ~n12259 & ~n12260;
  assign n12262 = pi452 & ~n12261;
  assign n12263 = ~n12258 & ~n12262;
  assign n12264 = ~pi355 & n12263;
  assign n12265 = ~n12254 & ~n12264;
  assign n12266 = pi458 & n12265;
  assign n12267 = ~pi355 & ~n12253;
  assign n12268 = pi355 & n12263;
  assign n12269 = ~n12267 & ~n12268;
  assign n12270 = ~pi458 & n12269;
  assign n12271 = n7606 & ~n12270;
  assign n12272 = ~n12266 & n12271;
  assign n12273 = pi458 & n12269;
  assign n12274 = ~pi458 & n12265;
  assign n12275 = ~n7606 & ~n12274;
  assign n12276 = ~n12273 & n12275;
  assign n12277 = pi1196 & ~n12276;
  assign n12278 = ~n12272 & n12277;
  assign n12279 = n12250 & ~n12278;
  assign n12280 = ~n12249 & ~n12279;
  assign n12281 = ~n7421 & ~n12280;
  assign n12282 = n7421 & n12160;
  assign n12283 = ~n12281 & ~n12282;
  assign n12284 = ~n7396 & n12283;
  assign n12285 = pi1199 & ~n12160;
  assign n12286 = pi351 & n12285;
  assign n12287 = ~n12284 & ~n12286;
  assign n12288 = ~pi461 & ~n12287;
  assign n12289 = ~n7667 & n12283;
  assign n12290 = ~pi351 & n12285;
  assign n12291 = ~n12289 & ~n12290;
  assign n12292 = pi461 & ~n12291;
  assign n12293 = ~n12288 & ~n12292;
  assign n12294 = ~pi357 & ~n12293;
  assign n12295 = ~pi461 & ~n12291;
  assign n12296 = pi461 & ~n12287;
  assign n12297 = ~n12295 & ~n12296;
  assign n12298 = pi357 & ~n12297;
  assign n12299 = ~n12294 & ~n12298;
  assign n12300 = ~pi356 & ~n12299;
  assign n12301 = ~pi357 & ~n12297;
  assign n12302 = pi357 & ~n12293;
  assign n12303 = ~n12301 & ~n12302;
  assign n12304 = pi356 & ~n12303;
  assign n12305 = ~n12300 & ~n12304;
  assign n12306 = pi354 & ~n12305;
  assign n12307 = ~pi356 & ~n12303;
  assign n12308 = pi356 & ~n12299;
  assign n12309 = ~n12307 & ~n12308;
  assign n12310 = ~pi354 & ~n12309;
  assign n12311 = n7392 & ~n12310;
  assign n12312 = ~n12306 & n12311;
  assign n12313 = pi354 & ~n12309;
  assign n12314 = ~pi354 & ~n12305;
  assign n12315 = ~n7392 & ~n12314;
  assign n12316 = ~n12313 & n12315;
  assign n12317 = ~pi591 & ~n12316;
  assign n12318 = ~n12312 & n12317;
  assign n12319 = n12245 & ~n12318;
  assign n12320 = ~pi1197 & ~n7877;
  assign n12321 = ~n12160 & ~n12320;
  assign n12322 = n8219 & ~n12118;
  assign n12323 = ~pi411 & n12111;
  assign n12324 = n7899 & ~n12323;
  assign n12325 = pi411 & n12139;
  assign n12326 = n12324 & ~n12325;
  assign n12327 = ~n7899 & ~n12111;
  assign n12328 = ~n7901 & ~n12327;
  assign n12329 = ~pi411 & n12139;
  assign n12330 = ~n12328 & ~n12329;
  assign n12331 = ~n12326 & ~n12330;
  assign n12332 = ~n12121 & ~n12331;
  assign n12333 = n12142 & ~n12332;
  assign n12334 = pi411 & n12147;
  assign n12335 = n12324 & ~n12334;
  assign n12336 = ~pi411 & n12147;
  assign n12337 = ~n12328 & ~n12336;
  assign n12338 = ~n12335 & ~n12337;
  assign n12339 = ~n12121 & ~n12338;
  assign n12340 = n12149 & ~n12339;
  assign n12341 = ~n12151 & ~n12340;
  assign n12342 = ~n12333 & n12341;
  assign n12343 = ~pi75 & ~n12342;
  assign n12344 = ~n12120 & ~n12343;
  assign n12345 = pi567 & ~n12344;
  assign n12346 = n12119 & ~n12345;
  assign n12347 = n12322 & ~n12346;
  assign n12348 = ~n12117 & ~n12162;
  assign n12349 = ~pi1199 & n12348;
  assign n12350 = ~n12347 & n12349;
  assign n12351 = n7940 & n12150;
  assign n12352 = n7940 & n12139;
  assign n12353 = ~n7940 & n12111;
  assign n12354 = ~n12352 & ~n12353;
  assign n12355 = n12143 & ~n12354;
  assign n12356 = ~n12351 & ~n12355;
  assign n12357 = n12342 & n12356;
  assign n12358 = n12322 & ~n12357;
  assign n12359 = n7940 & n12147;
  assign n12360 = ~n12353 & ~n12359;
  assign n12361 = n12150 & ~n12360;
  assign n12362 = ~n12151 & ~n12361;
  assign n12363 = ~n12355 & n12362;
  assign n12364 = n8313 & ~n12118;
  assign n12365 = ~n12363 & n12364;
  assign n12366 = ~n12358 & ~n12365;
  assign n12367 = ~pi75 & pi567;
  assign n12368 = ~n12366 & n12367;
  assign n12369 = n7910 & n12119;
  assign n12370 = ~n12114 & ~n12369;
  assign n12371 = pi1199 & ~n12370;
  assign n12372 = ~n12368 & n12371;
  assign n12373 = ~n7877 & ~n12372;
  assign n12374 = ~n12350 & n12373;
  assign n12375 = ~pi1197 & n12374;
  assign n12376 = ~n12321 & ~n12375;
  assign n12377 = ~pi333 & ~n12376;
  assign n12378 = n7877 & ~n12160;
  assign n12379 = ~n12374 & ~n12378;
  assign n12380 = pi333 & ~n12379;
  assign n12381 = ~n12377 & ~n12380;
  assign n12382 = ~pi391 & ~n12381;
  assign n12383 = pi333 & ~n12376;
  assign n12384 = ~pi333 & ~n12379;
  assign n12385 = ~n12383 & ~n12384;
  assign n12386 = pi391 & ~n12385;
  assign n12387 = ~n12382 & ~n12386;
  assign n12388 = ~pi392 & ~n12387;
  assign n12389 = ~pi391 & ~n12385;
  assign n12390 = pi391 & ~n12381;
  assign n12391 = ~n12389 & ~n12390;
  assign n12392 = pi392 & ~n12391;
  assign n12393 = ~n12388 & ~n12392;
  assign n12394 = pi393 & ~n12393;
  assign n12395 = ~pi392 & ~n12391;
  assign n12396 = pi392 & ~n12387;
  assign n12397 = ~n12395 & ~n12396;
  assign n12398 = ~pi393 & ~n12397;
  assign n12399 = n8215 & ~n12398;
  assign n12400 = ~n12394 & n12399;
  assign n12401 = pi393 & ~n12397;
  assign n12402 = ~pi393 & ~n12393;
  assign n12403 = ~n8215 & ~n12402;
  assign n12404 = ~n12401 & n12403;
  assign n12405 = pi591 & ~n12404;
  assign n12406 = ~n12400 & n12405;
  assign n12407 = ~pi592 & ~n12114;
  assign n12408 = pi592 & n12158;
  assign n12409 = ~n12407 & ~n12408;
  assign n12410 = ~n8699 & n12409;
  assign n12411 = n8699 & n12114;
  assign n12412 = pi1199 & ~n12411;
  assign n12413 = ~n12410 & n12412;
  assign n12414 = ~pi1197 & ~n12114;
  assign n12415 = ~n7722 & ~n12414;
  assign n12416 = n7746 & n12409;
  assign n12417 = ~n7746 & n12114;
  assign n12418 = pi1197 & ~n12417;
  assign n12419 = ~n12416 & n12418;
  assign n12420 = n12415 & ~n12419;
  assign n12421 = n7722 & n12409;
  assign n12422 = ~pi1199 & ~n12421;
  assign n12423 = ~n12420 & n12422;
  assign n12424 = ~n12413 & ~n12423;
  assign n12425 = ~pi1198 & ~n12424;
  assign n12426 = pi1198 & ~n12409;
  assign n12427 = ~n12425 & ~n12426;
  assign n12428 = ~pi374 & ~n12427;
  assign n12429 = pi374 & ~n12424;
  assign n12430 = ~n12428 & ~n12429;
  assign n12431 = ~pi369 & ~n12430;
  assign n12432 = pi371 & n8166;
  assign n12433 = ~pi371 & ~n8166;
  assign n12434 = ~n12432 & ~n12433;
  assign n12435 = pi370 & ~n12434;
  assign n12436 = ~pi370 & n12434;
  assign n12437 = ~n12435 & ~n12436;
  assign n12438 = ~pi374 & ~n12424;
  assign n12439 = pi374 & ~n12427;
  assign n12440 = ~n12438 & ~n12439;
  assign n12441 = pi369 & ~n12440;
  assign n12442 = n12437 & ~n12441;
  assign n12443 = ~n12431 & n12442;
  assign n12444 = pi369 & ~n12430;
  assign n12445 = ~pi369 & ~n12440;
  assign n12446 = ~n12437 & ~n12445;
  assign n12447 = ~n12444 & n12446;
  assign n12448 = ~pi591 & ~n12447;
  assign n12449 = ~n12443 & n12448;
  assign n12450 = ~pi590 & ~n12449;
  assign n12451 = ~n12406 & n12450;
  assign n12452 = ~pi588 & ~n12451;
  assign n12453 = ~n12319 & n12452;
  assign n12454 = n7697 & ~n12453;
  assign n12455 = ~n12243 & n12454;
  assign n12456 = ~n8021 & ~n12112;
  assign n12457 = ~pi122 & n12456;
  assign n12458 = n7536 & ~n12457;
  assign n12459 = n3207 & ~n12121;
  assign n12460 = ~n12458 & n12459;
  assign n12461 = ~pi87 & n12459;
  assign n12462 = ~n12139 & n12461;
  assign n12463 = pi87 & n12459;
  assign n12464 = ~n12147 & n12463;
  assign n12465 = ~n12462 & ~n12464;
  assign n12466 = pi122 & ~n12465;
  assign n12467 = ~n12460 & ~n12466;
  assign n12468 = ~pi75 & ~n12467;
  assign n12469 = pi567 & n7422;
  assign n12470 = ~n7457 & n12456;
  assign n12471 = n12469 & ~n12470;
  assign n12472 = ~n12468 & n12471;
  assign n12473 = ~n7422 & ~n12456;
  assign n12474 = ~n12113 & ~n12473;
  assign n12475 = ~n12472 & n12474;
  assign n12476 = ~pi592 & ~n12475;
  assign n12477 = ~n12117 & ~n12476;
  assign n12478 = ~n8480 & n12477;
  assign n12479 = pi443 & ~n12477;
  assign n12480 = ~n12164 & ~n12479;
  assign n12481 = n8568 & n12480;
  assign n12482 = ~pi443 & ~n12477;
  assign n12483 = ~n12168 & ~n12482;
  assign n12484 = ~n8568 & n12483;
  assign n12485 = ~n12481 & ~n12484;
  assign n12486 = pi435 & ~n12485;
  assign n12487 = pi444 & n12480;
  assign n12488 = ~pi444 & n12483;
  assign n12489 = ~pi436 & ~n12488;
  assign n12490 = ~n12487 & n12489;
  assign n12491 = pi444 & n12483;
  assign n12492 = ~pi444 & n12480;
  assign n12493 = pi436 & ~n12492;
  assign n12494 = ~n12491 & n12493;
  assign n12495 = ~n12490 & ~n12494;
  assign n12496 = ~pi435 & n12495;
  assign n12497 = ~n12486 & ~n12496;
  assign n12498 = pi429 & n12497;
  assign n12499 = ~pi435 & ~n12485;
  assign n12500 = pi435 & n12495;
  assign n12501 = ~n12499 & ~n12500;
  assign n12502 = ~pi429 & n12501;
  assign n12503 = ~n8505 & ~n12502;
  assign n12504 = ~n12498 & n12503;
  assign n12505 = pi429 & n12501;
  assign n12506 = ~pi429 & n12497;
  assign n12507 = n8505 & ~n12506;
  assign n12508 = ~n12505 & n12507;
  assign n12509 = pi1196 & ~n12508;
  assign n12510 = ~n12504 & n12509;
  assign n12511 = n12163 & ~n12510;
  assign n12512 = ~n12478 & ~n12511;
  assign n12513 = ~pi428 & ~n12512;
  assign n12514 = pi428 & n12477;
  assign n12515 = ~n12513 & ~n12514;
  assign n12516 = ~pi427 & ~n12515;
  assign n12517 = pi428 & ~n12512;
  assign n12518 = ~pi428 & n12477;
  assign n12519 = ~n12517 & ~n12518;
  assign n12520 = pi427 & ~n12519;
  assign n12521 = ~n12516 & ~n12520;
  assign n12522 = pi430 & ~n12521;
  assign n12523 = ~pi427 & ~n12519;
  assign n12524 = pi427 & ~n12515;
  assign n12525 = ~n12523 & ~n12524;
  assign n12526 = ~pi430 & ~n12525;
  assign n12527 = ~n12522 & ~n12526;
  assign n12528 = pi426 & ~n12527;
  assign n12529 = pi430 & ~n12525;
  assign n12530 = ~pi430 & ~n12521;
  assign n12531 = ~n12529 & ~n12530;
  assign n12532 = ~pi426 & ~n12531;
  assign n12533 = ~n12528 & ~n12532;
  assign n12534 = pi445 & ~n12533;
  assign n12535 = pi426 & ~n12531;
  assign n12536 = ~pi426 & ~n12527;
  assign n12537 = ~n12535 & ~n12536;
  assign n12538 = ~pi445 & ~n12537;
  assign n12539 = ~n12534 & ~n12538;
  assign n12540 = pi448 & n12539;
  assign n12541 = pi445 & ~n12537;
  assign n12542 = ~pi445 & ~n12533;
  assign n12543 = ~n12541 & ~n12542;
  assign n12544 = ~pi448 & n12543;
  assign n12545 = n8426 & ~n12544;
  assign n12546 = ~n12540 & n12545;
  assign n12547 = ~pi448 & n12539;
  assign n12548 = pi448 & n12543;
  assign n12549 = ~n8426 & ~n12548;
  assign n12550 = ~n12547 & n12549;
  assign n12551 = pi1199 & ~n12550;
  assign n12552 = ~n12546 & n12551;
  assign n12553 = ~pi1199 & n12512;
  assign n12554 = n8558 & ~n12553;
  assign n12555 = ~n12552 & n12554;
  assign n12556 = n12116 & ~n12555;
  assign n12557 = ~n8657 & n12477;
  assign n12558 = ~n12246 & ~n12557;
  assign n12559 = pi1198 & ~n12558;
  assign n12560 = ~n7591 & n12477;
  assign n12561 = ~n12251 & ~n12560;
  assign n12562 = ~pi355 & ~n12561;
  assign n12563 = ~pi455 & ~n12477;
  assign n12564 = ~n12255 & ~n12563;
  assign n12565 = ~pi452 & ~n12564;
  assign n12566 = pi455 & ~n12477;
  assign n12567 = ~n12259 & ~n12566;
  assign n12568 = pi452 & ~n12567;
  assign n12569 = ~n12565 & ~n12568;
  assign n12570 = pi355 & n12569;
  assign n12571 = ~n12562 & ~n12570;
  assign n12572 = pi458 & n12571;
  assign n12573 = pi355 & ~n12561;
  assign n12574 = ~pi355 & n12569;
  assign n12575 = ~n12573 & ~n12574;
  assign n12576 = ~pi458 & n12575;
  assign n12577 = ~n7606 & ~n12576;
  assign n12578 = ~n12572 & n12577;
  assign n12579 = pi458 & n12575;
  assign n12580 = ~pi458 & n12571;
  assign n12581 = n7606 & ~n12580;
  assign n12582 = ~n12579 & n12581;
  assign n12583 = pi1196 & ~n12582;
  assign n12584 = ~n12578 & n12583;
  assign n12585 = n12250 & ~n12584;
  assign n12586 = ~n12559 & ~n12585;
  assign n12587 = ~n7421 & ~n12586;
  assign n12588 = n7421 & n12477;
  assign n12589 = ~n12587 & ~n12588;
  assign n12590 = ~n7396 & n12589;
  assign n12591 = pi1199 & ~n12477;
  assign n12592 = pi351 & n12591;
  assign n12593 = ~n12590 & ~n12592;
  assign n12594 = ~pi461 & ~n12593;
  assign n12595 = ~n7667 & n12589;
  assign n12596 = ~pi351 & n12591;
  assign n12597 = ~n12595 & ~n12596;
  assign n12598 = pi461 & ~n12597;
  assign n12599 = ~n12594 & ~n12598;
  assign n12600 = ~pi357 & ~n12599;
  assign n12601 = ~pi461 & ~n12597;
  assign n12602 = pi461 & ~n12593;
  assign n12603 = ~n12601 & ~n12602;
  assign n12604 = pi357 & ~n12603;
  assign n12605 = ~n12600 & ~n12604;
  assign n12606 = ~pi356 & ~n12605;
  assign n12607 = ~pi357 & ~n12603;
  assign n12608 = pi357 & ~n12599;
  assign n12609 = ~n12607 & ~n12608;
  assign n12610 = pi356 & ~n12609;
  assign n12611 = ~n12606 & ~n12610;
  assign n12612 = pi354 & ~n12611;
  assign n12613 = ~pi356 & ~n12609;
  assign n12614 = pi356 & ~n12605;
  assign n12615 = ~n12613 & ~n12614;
  assign n12616 = ~pi354 & ~n12615;
  assign n12617 = n7392 & ~n12616;
  assign n12618 = ~n12612 & n12617;
  assign n12619 = pi354 & ~n12615;
  assign n12620 = ~pi354 & ~n12611;
  assign n12621 = ~n7392 & ~n12620;
  assign n12622 = ~n12619 & n12621;
  assign n12623 = ~pi591 & ~n12622;
  assign n12624 = ~n12618 & n12623;
  assign n12625 = n12245 & ~n12624;
  assign n12626 = pi367 & ~n12114;
  assign n12627 = pi592 & ~n12475;
  assign n12628 = ~n12407 & ~n12627;
  assign n12629 = ~pi367 & ~n12628;
  assign n12630 = ~n12626 & ~n12629;
  assign n12631 = ~n7725 & n12630;
  assign n12632 = ~pi367 & ~n12114;
  assign n12633 = pi367 & ~n12628;
  assign n12634 = ~n12632 & ~n12633;
  assign n12635 = n7725 & n12634;
  assign n12636 = ~n12631 & ~n12635;
  assign n12637 = n7728 & n12636;
  assign n12638 = n7725 & ~n12630;
  assign n12639 = ~n7725 & ~n12634;
  assign n12640 = ~n12638 & ~n12639;
  assign n12641 = ~n7728 & ~n12640;
  assign n12642 = n7737 & ~n12641;
  assign n12643 = ~n12637 & n12642;
  assign n12644 = ~n7728 & n12636;
  assign n12645 = n7728 & ~n12640;
  assign n12646 = ~n7737 & ~n12645;
  assign n12647 = ~n12644 & n12646;
  assign n12648 = pi1197 & ~n12647;
  assign n12649 = ~n12643 & n12648;
  assign n12650 = n12415 & ~n12649;
  assign n12651 = n7722 & n12628;
  assign n12652 = ~pi1199 & ~n12651;
  assign n12653 = ~n12650 & n12652;
  assign n12654 = ~pi1198 & n12653;
  assign n12655 = ~n8699 & n12628;
  assign n12656 = ~n12411 & ~n12655;
  assign n12657 = n7802 & n12656;
  assign n12658 = pi1198 & ~n12628;
  assign n12659 = ~n12657 & ~n12658;
  assign n12660 = ~n12654 & n12659;
  assign n12661 = ~pi374 & ~n12660;
  assign n12662 = pi1199 & n12656;
  assign n12663 = ~n12653 & ~n12662;
  assign n12664 = pi374 & ~n12663;
  assign n12665 = ~n12661 & ~n12664;
  assign n12666 = pi369 & ~n12665;
  assign n12667 = ~pi374 & ~n12663;
  assign n12668 = pi374 & ~n12660;
  assign n12669 = ~n12667 & ~n12668;
  assign n12670 = ~pi369 & ~n12669;
  assign n12671 = ~n12437 & ~n12670;
  assign n12672 = ~n12666 & n12671;
  assign n12673 = ~pi369 & ~n12665;
  assign n12674 = pi369 & ~n12669;
  assign n12675 = n12437 & ~n12674;
  assign n12676 = ~n12673 & n12675;
  assign n12677 = ~pi591 & ~n12676;
  assign n12678 = ~n12672 & n12677;
  assign n12679 = ~n12320 & n12477;
  assign n12680 = pi397 & ~pi404;
  assign n12681 = ~pi397 & pi404;
  assign n12682 = ~n12680 & ~n12681;
  assign n12683 = pi411 & ~n12682;
  assign n12684 = ~pi411 & n12682;
  assign n12685 = ~n12683 & ~n12684;
  assign n12686 = ~n7881 & n12685;
  assign n12687 = n7881 & ~n12685;
  assign n12688 = ~n12686 & ~n12687;
  assign n12689 = n7474 & n12688;
  assign n12690 = ~n12111 & ~n12689;
  assign n12691 = ~pi412 & ~n12690;
  assign n12692 = n7474 & ~n12688;
  assign n12693 = ~n12111 & ~n12692;
  assign n12694 = pi412 & ~n12693;
  assign n12695 = ~n7893 & ~n12694;
  assign n12696 = ~n12691 & n12695;
  assign n12697 = pi412 & ~n12690;
  assign n12698 = ~pi412 & ~n12693;
  assign n12699 = n7893 & ~n12698;
  assign n12700 = ~n12697 & n12699;
  assign n12701 = ~pi122 & ~n12700;
  assign n12702 = ~n12696 & n12701;
  assign n12703 = ~n12111 & ~n12702;
  assign n12704 = n7536 & ~n12703;
  assign n12705 = ~n12121 & ~n12704;
  assign n12706 = pi567 & ~n12705;
  assign n12707 = ~n12113 & ~n12706;
  assign n12708 = ~n12119 & ~n12707;
  assign n12709 = pi122 & n12331;
  assign n12710 = ~n12702 & ~n12709;
  assign n12711 = n7536 & ~n12710;
  assign n12712 = n12461 & ~n12711;
  assign n12713 = pi122 & n12338;
  assign n12714 = ~n12702 & ~n12713;
  assign n12715 = n7536 & ~n12714;
  assign n12716 = n12463 & ~n12715;
  assign n12717 = ~n3207 & n12705;
  assign n12718 = ~n12716 & ~n12717;
  assign n12719 = ~n12712 & n12718;
  assign n12720 = ~pi75 & ~n12719;
  assign n12721 = pi75 & n12705;
  assign n12722 = n12469 & ~n12721;
  assign n12723 = ~n12720 & n12722;
  assign n12724 = ~n12708 & ~n12723;
  assign n12725 = n8219 & ~n12724;
  assign n12726 = ~n12162 & ~n12725;
  assign n12727 = ~pi1199 & ~n12726;
  assign n12728 = n7474 & n7940;
  assign n12729 = ~pi122 & ~n12111;
  assign n12730 = ~n12728 & n12729;
  assign n12731 = ~n12456 & ~n12730;
  assign n12732 = pi567 & n12731;
  assign n12733 = ~n12113 & ~n12732;
  assign n12734 = ~n12706 & n12733;
  assign n12735 = ~n12119 & ~n12734;
  assign n12736 = ~n12141 & ~n12730;
  assign n12737 = n3207 & ~n12736;
  assign n12738 = ~n12704 & n12737;
  assign n12739 = ~n12359 & n12463;
  assign n12740 = ~n12338 & n12739;
  assign n12741 = n12354 & n12461;
  assign n12742 = ~n12331 & n12741;
  assign n12743 = ~n12740 & ~n12742;
  assign n12744 = ~pi122 & n12728;
  assign n12745 = ~n12702 & ~n12744;
  assign n12746 = ~n12743 & n12745;
  assign n12747 = ~n12738 & ~n12746;
  assign n12748 = ~pi75 & ~n12747;
  assign n12749 = ~n7457 & ~n12731;
  assign n12750 = ~n12704 & n12749;
  assign n12751 = n12469 & ~n12750;
  assign n12752 = ~n12748 & n12751;
  assign n12753 = ~n12735 & ~n12752;
  assign n12754 = n8219 & ~n12753;
  assign n12755 = ~n12119 & ~n12733;
  assign n12756 = n12360 & n12463;
  assign n12757 = ~n12741 & ~n12756;
  assign n12758 = pi122 & ~n12757;
  assign n12759 = ~n12737 & ~n12758;
  assign n12760 = ~pi75 & ~n12759;
  assign n12761 = n12469 & ~n12749;
  assign n12762 = ~n12760 & n12761;
  assign n12763 = ~n12755 & ~n12762;
  assign n12764 = n8313 & ~n12763;
  assign n12765 = ~n12754 & ~n12764;
  assign n12766 = pi1199 & ~n12765;
  assign n12767 = ~n12117 & ~n12766;
  assign n12768 = ~n12727 & n12767;
  assign n12769 = n12320 & n12768;
  assign n12770 = ~n12679 & ~n12769;
  assign n12771 = pi333 & ~n12770;
  assign n12772 = n7877 & ~n12477;
  assign n12773 = ~n7877 & ~n12768;
  assign n12774 = ~n12772 & ~n12773;
  assign n12775 = ~pi333 & n12774;
  assign n12776 = ~n12771 & ~n12775;
  assign n12777 = pi391 & ~n12776;
  assign n12778 = pi333 & ~n12774;
  assign n12779 = ~pi333 & n12770;
  assign n12780 = ~n12778 & ~n12779;
  assign n12781 = ~pi391 & n12780;
  assign n12782 = ~n12777 & ~n12781;
  assign n12783 = ~pi392 & ~n12782;
  assign n12784 = ~pi391 & n12776;
  assign n12785 = pi391 & ~n12780;
  assign n12786 = ~n12784 & ~n12785;
  assign n12787 = pi392 & n12786;
  assign n12788 = ~n12783 & ~n12787;
  assign n12789 = pi393 & ~n12788;
  assign n12790 = pi392 & ~n12782;
  assign n12791 = ~pi392 & n12786;
  assign n12792 = ~n12790 & ~n12791;
  assign n12793 = ~pi393 & ~n12792;
  assign n12794 = ~n12789 & ~n12793;
  assign n12795 = n8215 & ~n12794;
  assign n12796 = pi393 & ~n12792;
  assign n12797 = ~pi393 & ~n12788;
  assign n12798 = ~n12796 & ~n12797;
  assign n12799 = ~n8215 & ~n12798;
  assign n12800 = pi591 & ~n12799;
  assign n12801 = ~n12795 & n12800;
  assign n12802 = ~pi590 & ~n12801;
  assign n12803 = ~n12678 & n12802;
  assign n12804 = ~pi588 & ~n12803;
  assign n12805 = ~n12625 & n12804;
  assign n12806 = ~n7697 & ~n12805;
  assign n12807 = ~n12556 & n12806;
  assign n12808 = ~pi80 & ~po1038;
  assign n12809 = ~n12807 & n12808;
  assign n12810 = ~n12455 & n12809;
  assign n12811 = ~n8658 & n12114;
  assign n12812 = ~n12320 & ~n12811;
  assign n12813 = n8219 & ~n12707;
  assign n12814 = n12348 & ~n12813;
  assign n12815 = ~pi1199 & ~n12814;
  assign n12816 = n8219 & ~n12734;
  assign n12817 = n8313 & ~n12733;
  assign n12818 = ~n12117 & ~n12817;
  assign n12819 = ~n12816 & n12818;
  assign n12820 = pi1199 & ~n12819;
  assign n12821 = ~n12815 & ~n12820;
  assign n12822 = n12320 & ~n12821;
  assign n12823 = ~n12812 & ~n12822;
  assign n12824 = pi333 & ~n12823;
  assign n12825 = n7877 & ~n12811;
  assign n12826 = ~n7877 & ~n12821;
  assign n12827 = ~n12825 & ~n12826;
  assign n12828 = ~pi333 & ~n12827;
  assign n12829 = ~n12824 & ~n12828;
  assign n12830 = ~pi391 & ~n12829;
  assign n12831 = pi392 & n8218;
  assign n12832 = ~pi392 & ~n8218;
  assign n12833 = ~n12831 & ~n12832;
  assign n12834 = ~pi333 & ~n12823;
  assign n12835 = pi333 & ~n12827;
  assign n12836 = ~n12834 & ~n12835;
  assign n12837 = pi391 & ~n12836;
  assign n12838 = n12833 & ~n12837;
  assign n12839 = ~n12830 & n12838;
  assign n12840 = ~pi391 & ~n12836;
  assign n12841 = pi391 & ~n12829;
  assign n12842 = ~n12833 & ~n12841;
  assign n12843 = ~n12840 & n12842;
  assign n12844 = pi591 & ~n12843;
  assign n12845 = ~n12839 & n12844;
  assign n12846 = n8089 & n8726;
  assign n12847 = n12114 & ~n12846;
  assign n12848 = ~pi591 & ~n12847;
  assign n12849 = ~pi590 & ~n12848;
  assign n12850 = ~n12845 & n12849;
  assign n12851 = ~n8666 & n12114;
  assign n12852 = n8662 & n12851;
  assign n12853 = ~n7396 & n12852;
  assign n12854 = ~n12811 & ~n12853;
  assign n12855 = pi461 & ~n12854;
  assign n12856 = ~n7667 & n12852;
  assign n12857 = ~n12811 & ~n12856;
  assign n12858 = ~pi461 & ~n12857;
  assign n12859 = ~n12855 & ~n12858;
  assign n12860 = pi357 & ~n12859;
  assign n12861 = pi461 & ~n12857;
  assign n12862 = ~pi461 & ~n12854;
  assign n12863 = ~n12861 & ~n12862;
  assign n12864 = ~pi357 & ~n12863;
  assign n12865 = ~n12860 & ~n12864;
  assign n12866 = pi356 & ~n12865;
  assign n12867 = pi357 & ~n12863;
  assign n12868 = ~pi357 & ~n12859;
  assign n12869 = ~n12867 & ~n12868;
  assign n12870 = ~pi356 & ~n12869;
  assign n12871 = ~n12866 & ~n12870;
  assign n12872 = ~pi354 & n12871;
  assign n12873 = pi356 & ~n12869;
  assign n12874 = ~pi356 & ~n12865;
  assign n12875 = ~n12873 & ~n12874;
  assign n12876 = pi354 & n12875;
  assign n12877 = n7392 & ~n12876;
  assign n12878 = ~n12872 & n12877;
  assign n12879 = ~pi354 & n12875;
  assign n12880 = pi354 & n12871;
  assign n12881 = ~n7392 & ~n12880;
  assign n12882 = ~n12879 & n12881;
  assign n12883 = ~pi591 & ~n12882;
  assign n12884 = ~n12878 & n12883;
  assign n12885 = n12245 & ~n12884;
  assign n12886 = ~pi588 & ~n12885;
  assign n12887 = ~n12850 & n12886;
  assign n12888 = n8658 & ~n8789;
  assign n12889 = n12114 & ~n12888;
  assign n12890 = ~pi428 & ~n12889;
  assign n12891 = pi428 & ~n12811;
  assign n12892 = ~n12890 & ~n12891;
  assign n12893 = ~pi427 & ~n12892;
  assign n12894 = pi428 & ~n12889;
  assign n12895 = ~pi428 & ~n12811;
  assign n12896 = ~n12894 & ~n12895;
  assign n12897 = pi427 & ~n12896;
  assign n12898 = ~n12893 & ~n12897;
  assign n12899 = ~pi430 & ~n12898;
  assign n12900 = ~pi427 & ~n12896;
  assign n12901 = pi427 & ~n12892;
  assign n12902 = ~n12900 & ~n12901;
  assign n12903 = pi430 & ~n12902;
  assign n12904 = ~n12899 & ~n12903;
  assign n12905 = ~pi426 & ~n12904;
  assign n12906 = ~pi430 & ~n12902;
  assign n12907 = pi430 & ~n12898;
  assign n12908 = ~n12906 & ~n12907;
  assign n12909 = pi426 & ~n12908;
  assign n12910 = ~n12905 & ~n12909;
  assign n12911 = ~pi445 & ~n12910;
  assign n12912 = ~pi426 & ~n12908;
  assign n12913 = pi426 & ~n12904;
  assign n12914 = ~n12912 & ~n12913;
  assign n12915 = pi445 & ~n12914;
  assign n12916 = ~n12911 & ~n12915;
  assign n12917 = pi448 & ~n12916;
  assign n12918 = ~pi445 & ~n12914;
  assign n12919 = pi445 & ~n12910;
  assign n12920 = ~n12918 & ~n12919;
  assign n12921 = ~pi448 & ~n12920;
  assign n12922 = ~n8426 & ~n12921;
  assign n12923 = ~n12917 & n12922;
  assign n12924 = ~pi448 & ~n12916;
  assign n12925 = pi448 & ~n12920;
  assign n12926 = n8426 & ~n12925;
  assign n12927 = ~n12924 & n12926;
  assign n12928 = pi1199 & ~n12927;
  assign n12929 = ~n12923 & n12928;
  assign n12930 = ~pi1199 & ~n12889;
  assign n12931 = n8558 & ~n12930;
  assign n12932 = ~n12929 & n12931;
  assign n12933 = n12116 & ~n12932;
  assign n12934 = ~n7697 & ~n12933;
  assign n12935 = ~n12887 & n12934;
  assign n12936 = n7697 & n12114;
  assign n12937 = ~pi80 & po1038;
  assign n12938 = ~n12936 & n12937;
  assign n12939 = ~n12935 & n12938;
  assign n12940 = ~pi217 & ~n12939;
  assign n12941 = ~n12810 & n12940;
  assign n12942 = ~pi80 & ~n12114;
  assign n12943 = pi217 & ~n12942;
  assign n12944 = n8830 & ~n12943;
  assign po238 = ~n12941 & n12944;
  assign n12946 = ~po1038 & n11242;
  assign n12947 = pi81 & ~pi314;
  assign n12948 = n2478 & n12947;
  assign n12949 = pi68 & ~pi81;
  assign n12950 = n2469 & n12949;
  assign n12951 = n10955 & n12950;
  assign n12952 = n11378 & n12951;
  assign n12953 = n2634 & n12952;
  assign n12954 = ~n12948 & ~n12953;
  assign po239 = n12946 & ~n12954;
  assign n12956 = pi69 & pi314;
  assign n12957 = n2601 & n12956;
  assign n12958 = pi66 & ~pi73;
  assign n12959 = n2457 & n12958;
  assign n12960 = n2471 & n12959;
  assign n12961 = ~n12957 & ~n12960;
  assign n12962 = n11043 & n11045;
  assign po240 = ~n12961 & n12962;
  assign n12964 = n2486 & n11044;
  assign n12965 = n2491 & n12964;
  assign n12966 = n2469 & n2608;
  assign n12967 = pi84 & n9087;
  assign n12968 = n12966 & n12967;
  assign n12969 = ~pi83 & ~n12968;
  assign n12970 = n12965 & ~n12969;
  assign n12971 = n2604 & n12970;
  assign n12972 = ~pi314 & ~n12971;
  assign n12973 = n2456 & n12968;
  assign n12974 = n12965 & n12973;
  assign n12975 = pi314 & ~n12974;
  assign n12976 = n10112 & ~n12975;
  assign po241 = ~n12972 & n12976;
  assign n12978 = pi211 & pi299;
  assign n12979 = pi219 & pi299;
  assign n12980 = ~n12978 & ~n12979;
  assign n12981 = ~n10761 & n12980;
  assign n12982 = ~po1038 & n12981;
  assign po242 = n11317 & n12982;
  assign n12984 = n6311 & n11046;
  assign n12985 = ~pi314 & n11047;
  assign n12986 = n11376 & n12985;
  assign n12987 = ~n12984 & ~n12986;
  assign po243 = n11043 & ~n12987;
  assign n12989 = n7513 & n11334;
  assign n12990 = n7509 & n11337;
  assign n12991 = ~n12989 & ~n12990;
  assign po244 = n10923 & ~n12991;
  assign n12993 = n2654 & n12964;
  assign n12994 = pi314 & n10112;
  assign n12995 = n2491 & n12994;
  assign po245 = n12993 & n12995;
  assign n12997 = n7474 & n10971;
  assign n12998 = ~pi1093 & ~n12997;
  assign n12999 = n7430 & n12124;
  assign n13000 = n10968 & n12999;
  assign n13001 = n10983 & n12122;
  assign n13002 = n13000 & n13001;
  assign n13003 = pi1093 & ~n13002;
  assign n13004 = n3268 & ~n10019;
  assign n13005 = ~n13003 & n13004;
  assign n13006 = ~n12998 & n13005;
  assign n13007 = n7697 & ~n13006;
  assign n13008 = n2497 & n7474;
  assign n13009 = ~pi1093 & n3093;
  assign n13010 = n3268 & n13009;
  assign n13011 = n13008 & n13010;
  assign n13012 = n11397 & n13011;
  assign n13013 = n2679 & n13012;
  assign n13014 = ~n7697 & ~n13013;
  assign n13015 = ~po1038 & ~n13014;
  assign po246 = ~n13007 & n13015;
  assign n13017 = pi70 & ~n8918;
  assign n13018 = n2454 & n8877;
  assign n13019 = n8892 & n13018;
  assign n13020 = n10134 & n13019;
  assign n13021 = pi841 & n7437;
  assign n13022 = n13020 & n13021;
  assign n13023 = ~pi70 & ~n13022;
  assign n13024 = n3094 & n10111;
  assign n13025 = ~n13023 & n13024;
  assign po247 = ~n13017 & n13025;
  assign n13027 = ~pi1050 & n9525;
  assign n13028 = ~pi90 & ~n13027;
  assign n13029 = n11266 & ~n13028;
  assign n13030 = ~n2706 & n13029;
  assign po248 = ~n7425 & n13030;
  assign n13032 = ~pi58 & n2565;
  assign n13033 = ~n10104 & ~n13032;
  assign n13034 = n2795 & n10108;
  assign n13035 = ~n13033 & n13034;
  assign n13036 = pi24 & n2536;
  assign n13037 = ~n2795 & n13036;
  assign n13038 = n11026 & n13037;
  assign n13039 = n2565 & n13038;
  assign n13040 = ~pi39 & ~n13039;
  assign n13041 = ~n13035 & n13040;
  assign n13042 = n10143 & ~n13041;
  assign po249 = n7518 & n13042;
  assign n13044 = pi92 & n3095;
  assign n13045 = n3406 & n11416;
  assign n13046 = n13044 & n13045;
  assign n13047 = n5767 & n6202;
  assign n13048 = n7513 & n13047;
  assign n13049 = n3474 & n6222;
  assign n13050 = n7509 & n13049;
  assign n13051 = ~n13048 & ~n13050;
  assign n13052 = n3277 & n11066;
  assign n13053 = ~n13051 & n13052;
  assign n13054 = ~n13046 & ~n13053;
  assign po250 = n10109 & ~n13054;
  assign n13056 = ~pi1050 & n3095;
  assign n13057 = pi92 & ~n13056;
  assign n13058 = pi93 & n11026;
  assign n13059 = n2735 & n13058;
  assign n13060 = ~pi92 & ~n13059;
  assign n13061 = n10110 & ~n13060;
  assign po251 = ~n13057 & n13061;
  assign n13063 = n11009 & n11226;
  assign n13064 = n2734 & n13063;
  assign n13065 = pi1093 & ~n13064;
  assign n13066 = n7491 & ~n13065;
  assign n13067 = n10197 & n11007;
  assign n13068 = ~n2589 & ~n13067;
  assign n13069 = n2514 & n10108;
  assign n13070 = pi252 & n13069;
  assign n13071 = ~n13068 & n13070;
  assign n13072 = ~n13066 & ~n13071;
  assign n13073 = ~po840 & ~n13072;
  assign n13074 = ~n13063 & ~n13073;
  assign n13075 = pi252 & n13072;
  assign n13076 = ~n13074 & ~n13075;
  assign n13077 = n8848 & ~n13076;
  assign n13078 = ~n8848 & ~n13063;
  assign n13079 = n10111 & ~n13078;
  assign po252 = ~n13077 & n13079;
  assign n13081 = ~n6221 & ~n6447;
  assign n13082 = n3475 & ~n11356;
  assign n13083 = n13081 & n13082;
  assign n13084 = ~n11359 & n11362;
  assign n13085 = ~n6447 & n13084;
  assign n13086 = pi39 & ~n13085;
  assign n13087 = ~n13083 & n13086;
  assign n13088 = n2450 & n11959;
  assign n13089 = n11395 & n13088;
  assign n13090 = ~pi332 & n10108;
  assign n13091 = n11225 & n13090;
  assign n13092 = n13020 & n13091;
  assign n13093 = ~pi39 & ~n13092;
  assign n13094 = ~n13089 & n13093;
  assign n13095 = n10146 & ~n13094;
  assign po253 = ~n13087 & n13095;
  assign n13097 = n10254 & n13088;
  assign n13098 = pi479 & ~po840;
  assign n13099 = n2935 & n13098;
  assign n13100 = pi96 & n2725;
  assign n13101 = n2534 & n13100;
  assign n13102 = ~n13098 & n13101;
  assign n13103 = n2737 & n13102;
  assign n13104 = ~n13099 & ~n13103;
  assign n13105 = ~pi95 & ~n13104;
  assign n13106 = ~n13097 & ~n13105;
  assign po254 = n10111 & ~n13106;
  assign n13108 = pi39 & pi593;
  assign n13109 = ~n11364 & n13108;
  assign n13110 = ~n6447 & n13109;
  assign n13111 = n6143 & n13098;
  assign n13112 = ~po740 & ~n13111;
  assign n13113 = ~pi96 & n10115;
  assign n13114 = ~n13112 & n13113;
  assign n13115 = n11423 & n13114;
  assign n13116 = ~n13110 & ~n13115;
  assign po255 = n10146 & ~n13116;
  assign n13118 = ~pi92 & n11417;
  assign n13119 = ~n13044 & ~n13118;
  assign n13120 = pi314 & pi1050;
  assign n13121 = n10110 & n13120;
  assign po256 = ~n13119 & n13121;
  assign n13123 = ~pi72 & pi99;
  assign n13124 = ~n8064 & ~n13123;
  assign n13125 = ~n2734 & n13123;
  assign n13126 = n8064 & ~n13125;
  assign n13127 = ~n10259 & n13123;
  assign n13128 = n6246 & n10855;
  assign n13129 = ~n13127 & ~n13128;
  assign n13130 = n10390 & ~n13129;
  assign n13131 = n13126 & ~n13130;
  assign n13132 = ~n13124 & ~n13131;
  assign n13133 = ~pi39 & ~n13132;
  assign n13134 = ~pi72 & pi152;
  assign n13135 = n10267 & n13134;
  assign n13136 = pi299 & n13135;
  assign n13137 = ~pi72 & n10271;
  assign n13138 = n10273 & n13137;
  assign n13139 = ~n13136 & ~n13138;
  assign n13140 = pi232 & ~n13139;
  assign n13141 = pi39 & ~n13140;
  assign n13142 = n3241 & ~n13141;
  assign n13143 = ~n13133 & n13142;
  assign n13144 = ~pi39 & ~n13123;
  assign n13145 = ~n13141 & ~n13144;
  assign n13146 = ~n3241 & n13145;
  assign n13147 = pi75 & ~n13146;
  assign n13148 = ~n13143 & n13147;
  assign n13149 = pi41 & pi72;
  assign n13150 = pi99 & ~n13149;
  assign n13151 = ~n10319 & n13150;
  assign n13152 = n10684 & ~n13151;
  assign n13153 = ~n10329 & n13150;
  assign n13154 = n10683 & ~n13153;
  assign n13155 = ~n13152 & ~n13154;
  assign n13156 = pi228 & ~n13155;
  assign n13157 = ~n10371 & n13150;
  assign n13158 = ~pi228 & ~n10473;
  assign n13159 = ~n13157 & n13158;
  assign n13160 = ~pi39 & ~n13159;
  assign n13161 = ~n13156 & n13160;
  assign n13162 = n10420 & ~n13139;
  assign n13163 = ~n10884 & n13162;
  assign n13164 = n3206 & ~n13163;
  assign n13165 = ~n13161 & n13164;
  assign n13166 = ~n10387 & n13123;
  assign n13167 = n6245 & n10246;
  assign n13168 = ~n13166 & ~n13167;
  assign n13169 = n10390 & ~n13168;
  assign n13170 = n13126 & ~n13169;
  assign n13171 = ~n13124 & ~n13170;
  assign n13172 = ~pi39 & ~n13171;
  assign n13173 = ~n13141 & ~n13172;
  assign n13174 = n6235 & ~n13173;
  assign n13175 = pi38 & ~n13145;
  assign n13176 = ~pi87 & ~n13175;
  assign n13177 = ~n13174 & n13176;
  assign n13178 = ~n13165 & n13177;
  assign n13179 = pi228 & n10501;
  assign n13180 = pi228 & n10384;
  assign n13181 = n13123 & ~n13180;
  assign n13182 = n3276 & ~n13181;
  assign n13183 = ~n13179 & n13182;
  assign n13184 = ~n3276 & ~n13145;
  assign n13185 = pi87 & ~n13184;
  assign n13186 = ~n13183 & n13185;
  assign n13187 = ~pi75 & ~n13186;
  assign n13188 = ~n13178 & n13187;
  assign n13189 = ~n13148 & ~n13188;
  assign n13190 = n7422 & ~n13189;
  assign n13191 = ~n7422 & ~n13145;
  assign n13192 = ~po1038 & ~n13191;
  assign n13193 = ~n13190 & n13192;
  assign n13194 = pi232 & n13135;
  assign n13195 = pi39 & ~n13194;
  assign n13196 = po1038 & ~n13144;
  assign n13197 = ~n13195 & n13196;
  assign po257 = n13193 | n13197;
  assign n13199 = ~n7462 & n10023;
  assign n13200 = pi129 & ~n13199;
  assign n13201 = n6239 & ~n13200;
  assign n13202 = n6243 & ~n6262;
  assign n13203 = pi129 & ~n10023;
  assign n13204 = ~n6242 & ~n13203;
  assign n13205 = ~n13202 & ~n13204;
  assign n13206 = ~n13201 & n13205;
  assign n13207 = ~pi75 & n3221;
  assign n13208 = n6235 & n13207;
  assign n13209 = ~n13206 & n13208;
  assign n13210 = ~pi24 & n8926;
  assign n13211 = po840 & n13210;
  assign n13212 = ~n8923 & n13211;
  assign n13213 = ~n13209 & ~n13212;
  assign n13214 = n8841 & ~n13213;
  assign po258 = n3095 & n13214;
  assign n13216 = ~n8064 & ~n10252;
  assign n13217 = ~n2734 & n10252;
  assign n13218 = n8064 & ~n13217;
  assign n13219 = n2734 & ~n6253;
  assign n13220 = n10252 & ~n10258;
  assign n13221 = ~n10247 & ~n13220;
  assign n13222 = n13219 & ~n13221;
  assign n13223 = n13218 & ~n13222;
  assign n13224 = ~n13216 & ~n13223;
  assign n13225 = ~pi39 & ~n13224;
  assign n13226 = ~pi144 & pi174;
  assign n13227 = n10270 & n13226;
  assign n13228 = ~pi72 & n13227;
  assign n13229 = ~pi299 & ~n13228;
  assign n13230 = pi152 & n3383;
  assign n13231 = n6162 & n13230;
  assign n13232 = ~pi72 & n13231;
  assign n13233 = pi299 & ~n13232;
  assign n13234 = pi232 & ~n13233;
  assign n13235 = ~n13229 & n13234;
  assign n13236 = pi39 & ~n13235;
  assign n13237 = n3241 & ~n13236;
  assign n13238 = ~n13225 & n13237;
  assign n13239 = ~pi39 & ~n10252;
  assign n13240 = ~n13236 & ~n13239;
  assign n13241 = ~n3241 & n13240;
  assign n13242 = pi75 & ~n13241;
  assign n13243 = ~n13238 & n13242;
  assign n13244 = pi101 & ~n10317;
  assign n13245 = n2734 & ~n10305;
  assign n13246 = ~n13244 & n13245;
  assign n13247 = pi101 & ~n10327;
  assign n13248 = ~n2734 & ~n10324;
  assign n13249 = ~n13247 & n13248;
  assign n13250 = ~n13246 & ~n13249;
  assign n13251 = pi228 & ~n13250;
  assign n13252 = pi101 & ~n10369;
  assign n13253 = ~pi228 & ~n10363;
  assign n13254 = ~n13252 & n13253;
  assign n13255 = ~pi39 & ~n13254;
  assign n13256 = ~n13251 & n13255;
  assign n13257 = n10885 & n13227;
  assign n13258 = ~pi299 & ~n13257;
  assign n13259 = n10885 & n13231;
  assign n13260 = pi299 & ~n13259;
  assign n13261 = n10420 & ~n13260;
  assign n13262 = ~n13258 & n13261;
  assign n13263 = n3206 & ~n13262;
  assign n13264 = ~n13256 & n13263;
  assign n13265 = ~pi44 & n10889;
  assign n13266 = n10252 & ~n13265;
  assign n13267 = ~n10246 & ~n13266;
  assign n13268 = n13219 & ~n13267;
  assign n13269 = n13218 & ~n13268;
  assign n13270 = ~n13216 & ~n13269;
  assign n13271 = ~pi39 & ~n13270;
  assign n13272 = ~n13236 & ~n13271;
  assign n13273 = n6235 & ~n13272;
  assign n13274 = pi38 & ~n13240;
  assign n13275 = ~pi87 & ~n13274;
  assign n13276 = ~n13273 & n13275;
  assign n13277 = ~n13264 & n13276;
  assign n13278 = ~pi101 & n10902;
  assign n13279 = n10383 & n10901;
  assign n13280 = n10252 & ~n13279;
  assign n13281 = ~pi39 & ~n13280;
  assign n13282 = ~n13278 & n13281;
  assign n13283 = pi87 & ~n13236;
  assign n13284 = ~n13282 & n13283;
  assign n13285 = ~pi75 & ~n13284;
  assign n13286 = ~n13277 & n13285;
  assign n13287 = ~n13243 & ~n13286;
  assign n13288 = n7422 & ~n13287;
  assign n13289 = ~n7422 & ~n13240;
  assign n13290 = ~po1038 & ~n13289;
  assign n13291 = ~n13288 & n13290;
  assign n13292 = pi232 & n13232;
  assign n13293 = pi39 & ~n13292;
  assign n13294 = po1038 & ~n13239;
  assign n13295 = ~n13293 & n13294;
  assign po259 = n13291 | n13295;
  assign n13297 = n2660 & n8878;
  assign po260 = n12946 & n13297;
  assign n13299 = ~pi109 & ~n12993;
  assign n13300 = n6301 & ~n13299;
  assign n13301 = ~pi314 & ~n13300;
  assign n13302 = pi109 & n2574;
  assign n13303 = n2487 & n13302;
  assign n13304 = pi314 & ~n13303;
  assign n13305 = n11042 & ~n13304;
  assign po261 = ~n13301 & n13305;
  assign n13307 = n7697 & ~n8848;
  assign n13308 = n10020 & ~n13307;
  assign n13309 = n10358 & ~n13308;
  assign n13310 = ~pi110 & ~n13000;
  assign n13311 = ~pi47 & n10983;
  assign n13312 = ~n13310 & n13311;
  assign n13313 = n10337 & n13312;
  assign n13314 = ~po1057 & ~n13313;
  assign n13315 = po1057 & ~n13002;
  assign n13316 = ~n7463 & ~n10019;
  assign n13317 = ~n13315 & n13316;
  assign n13318 = ~n13314 & n13317;
  assign n13319 = n7463 & ~n10019;
  assign n13320 = n13313 & n13319;
  assign n13321 = ~n13318 & ~n13320;
  assign n13322 = ~n7697 & ~n13321;
  assign n13323 = ~n13309 & ~n13322;
  assign po262 = n10111 & ~n13323;
  assign n13325 = pi24 & n11224;
  assign n13326 = ~pi53 & ~n11223;
  assign n13327 = n2508 & ~n13326;
  assign n13328 = ~pi24 & n2514;
  assign n13329 = n13327 & n13328;
  assign n13330 = ~n13325 & ~n13329;
  assign n13331 = pi841 & ~n13330;
  assign n13332 = n8905 & n11204;
  assign n13333 = ~n13331 & ~n13332;
  assign po264 = n10112 & ~n13333;
  assign n13335 = ~pi999 & n10112;
  assign po265 = n11294 & n13335;
  assign n13337 = ~pi97 & n7434;
  assign n13338 = ~pi108 & ~n13337;
  assign n13339 = n2490 & ~n13338;
  assign n13340 = n10183 & n13339;
  assign n13341 = ~pi314 & ~n13340;
  assign n13342 = pi314 & ~n7436;
  assign n13343 = n7438 & ~n10206;
  assign n13344 = ~n13342 & n13343;
  assign n13345 = ~n13341 & n13344;
  assign n13346 = n7438 & n10206;
  assign n13347 = n13340 & n13346;
  assign n13348 = ~pi51 & ~n13347;
  assign n13349 = ~n13345 & n13348;
  assign n13350 = n3207 & n7475;
  assign n13351 = ~n13349 & n13350;
  assign n13352 = ~pi87 & ~n13351;
  assign n13353 = n6270 & n8841;
  assign po266 = ~n13352 & n13353;
  assign n13355 = n2593 & n11373;
  assign po267 = n12994 & n13355;
  assign n13357 = ~pi82 & pi111;
  assign n13358 = n8892 & n13357;
  assign n13359 = n11047 & n13358;
  assign n13360 = n2635 & n13359;
  assign n13361 = pi314 & n13360;
  assign n13362 = n8848 & n10020;
  assign n13363 = n10350 & n13362;
  assign n13364 = ~n13361 & ~n13363;
  assign po268 = n10112 & ~n13364;
  assign n13366 = pi72 & n10254;
  assign n13367 = ~pi314 & n13360;
  assign n13368 = n9127 & n13367;
  assign n13369 = ~n13366 & ~n13368;
  assign n13370 = n6360 & n10111;
  assign po269 = ~n13369 & n13370;
  assign po270 = ~pi124 | pi468;
  assign n13373 = ~pi99 & ~n10330;
  assign n13374 = ~n10320 & n13373;
  assign n13375 = pi113 & ~n10433;
  assign n13376 = ~n13374 & n13375;
  assign n13377 = n10687 & ~n13376;
  assign n13378 = pi113 & n10468;
  assign n13379 = ~pi228 & ~n10474;
  assign n13380 = ~n13378 & n13379;
  assign n13381 = ~pi39 & ~n13380;
  assign n13382 = ~n13377 & n13381;
  assign n13383 = n3206 & ~n13382;
  assign n13384 = ~pi39 & n10469;
  assign n13385 = pi38 & ~n13384;
  assign n13386 = n2734 & n8064;
  assign n13387 = n7525 & n10507;
  assign n13388 = ~n6252 & ~n13387;
  assign n13389 = n13386 & ~n13388;
  assign n13390 = n10469 & ~n13389;
  assign n13391 = ~n6252 & n13386;
  assign n13392 = ~pi113 & n13391;
  assign n13393 = n13167 & n13392;
  assign n13394 = ~n13390 & ~n13393;
  assign n13395 = ~pi39 & ~n13394;
  assign n13396 = n6235 & ~n13395;
  assign n13397 = ~n13385 & ~n13396;
  assign n13398 = ~n13383 & n13397;
  assign n13399 = ~pi87 & ~n13398;
  assign n13400 = n10469 & ~n10534;
  assign n13401 = ~pi113 & n13179;
  assign n13402 = ~n13400 & ~n13401;
  assign n13403 = n3276 & ~n13402;
  assign n13404 = ~n3206 & n13384;
  assign n13405 = pi87 & ~n13404;
  assign n13406 = ~n13403 & n13405;
  assign n13407 = ~n13399 & ~n13406;
  assign n13408 = ~pi75 & ~n13407;
  assign n13409 = n7465 & n13393;
  assign n13410 = ~n6252 & ~n10547;
  assign n13411 = n13386 & ~n13410;
  assign n13412 = n10469 & ~n13411;
  assign n13413 = ~n13409 & ~n13412;
  assign n13414 = n3222 & ~n13413;
  assign n13415 = ~n3241 & n13384;
  assign n13416 = pi75 & ~n13415;
  assign n13417 = ~n13414 & n13416;
  assign n13418 = ~n13408 & ~n13417;
  assign n13419 = n8841 & ~n13418;
  assign n13420 = ~n8841 & ~n13384;
  assign po271 = ~n13419 & ~n13420;
  assign n13422 = pi114 & n10739;
  assign n13423 = n11093 & ~n13422;
  assign n13424 = ~n10545 & n13423;
  assign n13425 = ~pi72 & pi114;
  assign n13426 = ~n11093 & ~n13425;
  assign n13427 = n3222 & ~n13426;
  assign n13428 = ~n13424 & n13427;
  assign n13429 = ~pi39 & n13425;
  assign n13430 = ~n3241 & n13429;
  assign n13431 = pi75 & ~n13430;
  assign n13432 = ~n13428 & n13431;
  assign n13433 = ~pi114 & ~n10690;
  assign n13434 = pi114 & ~n10679;
  assign n13435 = ~n13433 & ~n13434;
  assign n13436 = ~pi115 & ~n13435;
  assign n13437 = pi115 & ~n13425;
  assign n13438 = ~pi39 & ~n13437;
  assign n13439 = ~n13436 & n13438;
  assign n13440 = n3206 & ~n13439;
  assign n13441 = pi114 & ~n10510;
  assign n13442 = n11093 & ~n13441;
  assign n13443 = ~n10505 & n13442;
  assign n13444 = ~pi39 & ~n13426;
  assign n13445 = ~n13443 & n13444;
  assign n13446 = n6235 & ~n13445;
  assign n13447 = pi38 & ~n13429;
  assign n13448 = ~pi87 & ~n13447;
  assign n13449 = ~n13446 & n13448;
  assign n13450 = ~n13440 & n13449;
  assign n13451 = pi228 & n10508;
  assign n13452 = ~pi115 & n13451;
  assign n13453 = n13425 & ~n13452;
  assign n13454 = n3206 & ~n13453;
  assign n13455 = ~n10532 & n13454;
  assign n13456 = ~n3206 & ~n13429;
  assign n13457 = n11067 & ~n13456;
  assign n13458 = ~n13455 & n13457;
  assign n13459 = ~pi75 & ~n13458;
  assign n13460 = ~n13450 & n13459;
  assign n13461 = ~n13432 & ~n13460;
  assign n13462 = n8841 & ~n13461;
  assign n13463 = ~n8841 & ~n13429;
  assign po272 = ~n13462 & ~n13463;
  assign n13465 = ~pi52 & n11070;
  assign n13466 = ~pi115 & ~n13465;
  assign n13467 = n10503 & n13466;
  assign n13468 = n7465 & n13467;
  assign n13469 = pi115 & n10739;
  assign n13470 = n13386 & ~n13469;
  assign n13471 = ~n13468 & n13470;
  assign n13472 = ~pi72 & pi115;
  assign n13473 = ~n13386 & ~n13472;
  assign n13474 = n3222 & ~n13473;
  assign n13475 = ~n13471 & n13474;
  assign n13476 = ~pi39 & n13472;
  assign n13477 = ~n3241 & n13476;
  assign n13478 = pi75 & ~n13477;
  assign n13479 = ~n13475 & n13478;
  assign n13480 = pi115 & ~n10679;
  assign n13481 = ~pi115 & ~n10690;
  assign n13482 = ~pi39 & ~n13481;
  assign n13483 = ~n13480 & n13482;
  assign n13484 = n3206 & ~n13483;
  assign n13485 = pi115 & ~n10510;
  assign n13486 = n13386 & ~n13485;
  assign n13487 = ~n13467 & n13486;
  assign n13488 = ~pi39 & ~n13473;
  assign n13489 = ~n13487 & n13488;
  assign n13490 = n6235 & ~n13489;
  assign n13491 = pi38 & ~n13476;
  assign n13492 = ~pi87 & ~n13491;
  assign n13493 = ~n13490 & n13492;
  assign n13494 = ~n13484 & n13493;
  assign n13495 = ~n13451 & n13472;
  assign n13496 = n3206 & ~n13495;
  assign n13497 = ~n10531 & n13496;
  assign n13498 = ~n3206 & ~n13476;
  assign n13499 = n11067 & ~n13498;
  assign n13500 = ~n13497 & n13499;
  assign n13501 = ~pi75 & ~n13500;
  assign n13502 = ~n13494 & n13501;
  assign n13503 = ~n13479 & ~n13502;
  assign n13504 = n8841 & ~n13503;
  assign n13505 = ~n8841 & ~n13476;
  assign po273 = ~n13504 & ~n13505;
  assign n13507 = pi116 & n10453;
  assign n13508 = ~n2734 & ~n13507;
  assign n13509 = n2734 & ~n10437;
  assign n13510 = pi116 & ~n13509;
  assign n13511 = ~n10444 & ~n13510;
  assign n13512 = ~n13508 & ~n13511;
  assign n13513 = ~n2734 & n10457;
  assign n13514 = pi228 & ~n13513;
  assign n13515 = ~n13512 & n13514;
  assign n13516 = pi116 & ~n10470;
  assign n13517 = n10688 & ~n13516;
  assign n13518 = ~pi39 & ~n13517;
  assign n13519 = ~n13515 & n13518;
  assign n13520 = n3206 & ~n13519;
  assign n13521 = n10431 & ~n13386;
  assign n13522 = ~pi113 & n13387;
  assign n13523 = n10431 & ~n13522;
  assign n13524 = ~n10503 & ~n13523;
  assign n13525 = n13391 & ~n13524;
  assign n13526 = ~n13521 & ~n13525;
  assign n13527 = ~pi39 & ~n13526;
  assign n13528 = n6235 & ~n13527;
  assign n13529 = ~pi39 & n10431;
  assign n13530 = pi38 & ~n13529;
  assign n13531 = ~pi87 & ~n13530;
  assign n13532 = ~n13528 & n13531;
  assign n13533 = ~n13520 & n13532;
  assign n13534 = ~pi113 & n10534;
  assign n13535 = n10431 & ~n13534;
  assign n13536 = ~pi38 & ~n13535;
  assign n13537 = ~n10530 & n13536;
  assign n13538 = ~n13530 & ~n13537;
  assign n13539 = ~pi100 & ~n13538;
  assign n13540 = pi100 & ~n13529;
  assign n13541 = n11067 & ~n13540;
  assign n13542 = ~n13539 & n13541;
  assign n13543 = ~pi75 & ~n13542;
  assign n13544 = ~n13533 & n13543;
  assign n13545 = n10431 & ~n10548;
  assign n13546 = ~n10741 & ~n13545;
  assign n13547 = n13391 & ~n13546;
  assign n13548 = ~n13521 & ~n13547;
  assign n13549 = n3222 & ~n13548;
  assign n13550 = ~n3241 & n13529;
  assign n13551 = pi75 & ~n13550;
  assign n13552 = ~n13549 & n13551;
  assign n13553 = ~n13544 & ~n13552;
  assign n13554 = n8841 & ~n13553;
  assign n13555 = ~n8841 & ~n13529;
  assign po274 = ~n13554 & ~n13555;
  assign n13557 = n3657 & n7331;
  assign n13558 = ~n3656 & ~n13557;
  assign n13559 = ~pi38 & ~n13558;
  assign n13560 = ~pi87 & ~n13559;
  assign n13561 = n6270 & ~n13560;
  assign n13562 = ~pi92 & ~n13561;
  assign n13563 = ~pi54 & ~n7272;
  assign n13564 = ~pi74 & n13563;
  assign n13565 = ~n13562 & n13564;
  assign n13566 = ~pi55 & ~n13565;
  assign n13567 = ~n7314 & ~n13566;
  assign n13568 = ~pi56 & ~n13567;
  assign n13569 = ~n6104 & ~n13568;
  assign n13570 = ~pi62 & ~n13569;
  assign n13571 = ~pi57 & n6281;
  assign po275 = ~n13570 & n13571;
  assign n13573 = pi163 & n6162;
  assign n13574 = ~n11614 & ~n13573;
  assign n13575 = ~pi150 & ~n13574;
  assign n13576 = pi150 & n9643;
  assign n13577 = n11612 & n13576;
  assign n13578 = ~n13575 & ~n13577;
  assign n13579 = pi232 & ~n13578;
  assign n13580 = ~n8948 & n13579;
  assign n13581 = pi74 & ~n13580;
  assign n13582 = pi165 & n7462;
  assign n13583 = ~pi38 & ~pi54;
  assign n13584 = ~n13582 & ~n13583;
  assign n13585 = n8948 & n13584;
  assign n13586 = ~pi74 & ~n13580;
  assign n13587 = ~n13585 & n13586;
  assign n13588 = ~n13581 & ~n13587;
  assign n13589 = ~n3293 & ~n13588;
  assign n13590 = n3429 & ~n13589;
  assign n13591 = ~n9666 & ~n13590;
  assign n13592 = pi299 & n13578;
  assign n13593 = ~pi184 & ~n11627;
  assign n13594 = ~pi185 & n13593;
  assign n13595 = pi185 & ~n13593;
  assign n13596 = n6162 & ~n13595;
  assign n13597 = ~n13594 & n13596;
  assign n13598 = ~pi299 & ~n13597;
  assign n13599 = pi232 & ~n13598;
  assign n13600 = ~n13592 & n13599;
  assign n13601 = ~n8948 & n13600;
  assign n13602 = pi74 & ~n13601;
  assign n13603 = ~pi55 & ~n13602;
  assign n13604 = ~pi143 & ~pi299;
  assign n13605 = ~pi165 & pi299;
  assign n13606 = ~n13604 & ~n13605;
  assign n13607 = n7462 & n13606;
  assign n13608 = n8948 & ~n13607;
  assign n13609 = pi54 & ~n13608;
  assign n13610 = ~n13601 & n13609;
  assign n13611 = ~pi143 & ~n8984;
  assign n13612 = pi143 & ~n8986;
  assign n13613 = pi165 & ~n13612;
  assign n13614 = ~n13611 & n13613;
  assign n13615 = pi143 & ~pi165;
  assign n13616 = n8991 & n13615;
  assign n13617 = pi38 & ~n13616;
  assign n13618 = ~n13614 & n13617;
  assign n13619 = n3240 & ~n13618;
  assign n13620 = ~n6162 & n9293;
  assign n13621 = pi151 & ~pi168;
  assign n13622 = ~n9359 & n13621;
  assign n13623 = pi168 & n9349;
  assign n13624 = ~pi168 & n9352;
  assign n13625 = ~pi151 & ~n13624;
  assign n13626 = ~n13623 & n13625;
  assign n13627 = ~n13622 & ~n13626;
  assign n13628 = ~n13620 & ~n13627;
  assign n13629 = ~n6162 & ~n9293;
  assign n13630 = n6162 & ~n9319;
  assign n13631 = ~n13629 & ~n13630;
  assign n13632 = pi151 & pi168;
  assign n13633 = ~n13631 & n13632;
  assign n13634 = pi150 & ~n13633;
  assign n13635 = ~n13628 & n13634;
  assign n13636 = ~n9190 & ~n13629;
  assign n13637 = pi168 & n13636;
  assign n13638 = ~n9741 & ~n13629;
  assign n13639 = ~pi168 & n13638;
  assign n13640 = pi151 & ~n13639;
  assign n13641 = ~n13637 & n13640;
  assign n13642 = pi168 & n9287;
  assign n13643 = pi168 & n6162;
  assign n13644 = n9293 & ~n13643;
  assign n13645 = ~pi151 & ~n13644;
  assign n13646 = ~n13642 & n13645;
  assign n13647 = ~pi150 & ~n13646;
  assign n13648 = ~n13641 & n13647;
  assign n13649 = pi299 & ~n13648;
  assign n13650 = ~n13635 & n13649;
  assign n13651 = ~n9283 & ~n13620;
  assign n13652 = ~pi173 & ~n13651;
  assign n13653 = n6162 & ~n9134;
  assign n13654 = pi173 & ~n13629;
  assign n13655 = ~n13653 & n13654;
  assign n13656 = pi185 & ~n13655;
  assign n13657 = ~n13652 & n13656;
  assign n13658 = pi173 & n13636;
  assign n13659 = ~n9287 & ~n13620;
  assign n13660 = ~pi173 & ~n13659;
  assign n13661 = ~pi185 & ~n13660;
  assign n13662 = ~n13658 & n13661;
  assign n13663 = pi190 & ~n13662;
  assign n13664 = ~n13657 & n13663;
  assign n13665 = pi173 & ~n9733;
  assign n13666 = ~pi173 & ~n9305;
  assign n13667 = n6162 & ~n13666;
  assign n13668 = ~n13665 & n13667;
  assign n13669 = pi185 & ~n13620;
  assign n13670 = ~n13668 & n13669;
  assign n13671 = pi173 & n13638;
  assign n13672 = ~pi173 & n9293;
  assign n13673 = ~pi185 & ~n13672;
  assign n13674 = ~n13671 & n13673;
  assign n13675 = ~pi190 & ~n13674;
  assign n13676 = ~n13670 & n13675;
  assign n13677 = ~pi299 & ~n13676;
  assign n13678 = ~n13664 & n13677;
  assign n13679 = pi232 & ~n13678;
  assign n13680 = ~n13650 & n13679;
  assign n13681 = ~pi232 & n9293;
  assign n13682 = ~pi39 & ~n13681;
  assign n13683 = ~n13680 & n13682;
  assign n13684 = ~pi178 & ~pi299;
  assign n13685 = pi168 & n9020;
  assign n13686 = pi157 & n9031;
  assign n13687 = ~n13685 & ~n13686;
  assign n13688 = n6162 & n12051;
  assign n13689 = ~n13687 & n13688;
  assign n13690 = pi299 & ~n13689;
  assign n13691 = ~n13684 & ~n13690;
  assign n13692 = n8997 & ~n13691;
  assign n13693 = pi178 & ~n9054;
  assign n13694 = ~pi190 & ~n13693;
  assign n13695 = ~pi299 & ~n13694;
  assign n13696 = ~n13692 & ~n13695;
  assign n13697 = ~n9052 & ~n12046;
  assign n13698 = pi178 & ~n13697;
  assign n13699 = ~n9061 & n13698;
  assign n13700 = ~pi178 & ~n13697;
  assign n13701 = ~n9023 & n13700;
  assign n13702 = ~pi299 & ~n9018;
  assign n13703 = pi190 & n13702;
  assign n13704 = ~n13701 & n13703;
  assign n13705 = ~n13699 & n13704;
  assign n13706 = pi232 & ~n13705;
  assign n13707 = ~n13696 & n13706;
  assign n13708 = ~pi232 & n8997;
  assign n13709 = pi39 & ~n13708;
  assign n13710 = ~n13707 & n13709;
  assign n13711 = ~pi38 & ~n13710;
  assign n13712 = ~n13683 & n13711;
  assign n13713 = n13619 & ~n13712;
  assign n13714 = pi100 & ~n13600;
  assign n13715 = pi38 & ~n13607;
  assign n13716 = n7577 & ~n13715;
  assign n13717 = ~n9464 & n13716;
  assign n13718 = ~n13714 & ~n13717;
  assign n13719 = ~n13713 & n13718;
  assign n13720 = n3237 & ~n13719;
  assign n13721 = pi75 & ~n13600;
  assign n13722 = ~pi100 & ~n13715;
  assign n13723 = ~pi157 & pi299;
  assign n13724 = ~n13684 & ~n13723;
  assign n13725 = n7462 & n13724;
  assign n13726 = n9415 & n13725;
  assign n13727 = n9464 & ~n13726;
  assign n13728 = n13722 & ~n13727;
  assign n13729 = ~n13714 & ~n13728;
  assign n13730 = n9410 & ~n13729;
  assign n13731 = ~n13721 & ~n13730;
  assign n13732 = ~n13720 & n13731;
  assign n13733 = ~pi54 & ~n13732;
  assign n13734 = ~n13610 & ~n13733;
  assign n13735 = ~pi74 & ~n13734;
  assign n13736 = n13603 & ~n13735;
  assign n13737 = pi55 & ~n13581;
  assign n13738 = pi150 & n7462;
  assign n13739 = ~pi92 & n9415;
  assign n13740 = n13738 & n13739;
  assign n13741 = n8997 & n13583;
  assign n13742 = ~n13740 & n13741;
  assign n13743 = ~n13584 & ~n13742;
  assign n13744 = n8948 & ~n13743;
  assign n13745 = n13586 & ~n13744;
  assign n13746 = n13737 & ~n13745;
  assign n13747 = n3293 & ~n13746;
  assign n13748 = ~n13736 & n13747;
  assign n13749 = ~n13591 & ~n13748;
  assign n13750 = ~n8948 & ~n13579;
  assign n13751 = n8948 & n13582;
  assign n13752 = ~n3429 & ~n13751;
  assign n13753 = ~n13750 & n13752;
  assign n13754 = ~n13581 & n13753;
  assign n13755 = ~n13749 & ~n13754;
  assign n13756 = pi118 & n13755;
  assign n13757 = ~pi79 & n12102;
  assign n13758 = n6198 & ~n6447;
  assign n13759 = ~pi157 & n9494;
  assign n13760 = pi168 & ~n13759;
  assign n13761 = pi157 & ~n9489;
  assign n13762 = ~pi157 & ~pi168;
  assign n13763 = ~n9487 & n13762;
  assign n13764 = ~n13761 & ~n13763;
  assign n13765 = ~n13760 & n13764;
  assign n13766 = ~n13758 & ~n13765;
  assign n13767 = n13047 & ~n13766;
  assign n13768 = ~pi178 & ~n6215;
  assign n13769 = n9493 & n13768;
  assign n13770 = ~n13758 & ~n13769;
  assign n13771 = pi190 & ~n13770;
  assign n13772 = ~pi178 & ~n13081;
  assign n13773 = pi178 & ~n9472;
  assign n13774 = ~n13758 & n13773;
  assign n13775 = ~pi190 & ~n13774;
  assign n13776 = ~n13772 & n13775;
  assign n13777 = ~n13771 & ~n13776;
  assign n13778 = n13049 & ~n13777;
  assign n13779 = pi232 & ~n13778;
  assign n13780 = ~n13767 & n13779;
  assign n13781 = n7276 & n9477;
  assign n13782 = ~n6200 & n13047;
  assign n13783 = ~n6447 & n13782;
  assign n13784 = ~pi232 & ~n13783;
  assign n13785 = ~n13781 & n13784;
  assign n13786 = pi39 & ~n13785;
  assign n13787 = ~n13780 & n13786;
  assign n13788 = n9526 & n13621;
  assign n13789 = ~pi168 & n9527;
  assign n13790 = pi168 & ~n9524;
  assign n13791 = ~pi151 & ~n13790;
  assign n13792 = ~n13789 & n13791;
  assign n13793 = ~n13788 & ~n13792;
  assign n13794 = n9520 & ~n13793;
  assign n13795 = pi150 & ~n13794;
  assign n13796 = ~pi151 & n9513;
  assign n13797 = n9565 & ~n13796;
  assign n13798 = ~pi168 & ~n13797;
  assign n13799 = ~pi151 & n9535;
  assign n13800 = n9568 & ~n13799;
  assign n13801 = n13643 & ~n13800;
  assign n13802 = ~pi150 & ~n13801;
  assign n13803 = ~n13798 & n13802;
  assign n13804 = ~n13795 & ~n13803;
  assign n13805 = ~n9513 & ~n11969;
  assign n13806 = ~n6162 & ~n13805;
  assign n13807 = pi299 & ~n13806;
  assign n13808 = ~n13804 & n13807;
  assign n13809 = n6360 & n9526;
  assign n13810 = pi173 & n13809;
  assign n13811 = ~pi173 & n6360;
  assign n13812 = ~n9527 & n13811;
  assign n13813 = ~n13810 & ~n13812;
  assign n13814 = ~pi190 & n6162;
  assign n13815 = ~n13813 & n13814;
  assign n13816 = ~pi173 & pi190;
  assign n13817 = n9539 & n13816;
  assign n13818 = pi185 & ~n13817;
  assign n13819 = ~n13815 & n13818;
  assign n13820 = ~pi173 & n9513;
  assign n13821 = n9545 & ~n13820;
  assign n13822 = ~pi190 & ~n13821;
  assign n13823 = pi173 & n9548;
  assign n13824 = pi190 & n9537;
  assign n13825 = ~n13823 & n13824;
  assign n13826 = ~pi185 & ~n13825;
  assign n13827 = ~n13822 & n13826;
  assign n13828 = ~n13819 & ~n13827;
  assign n13829 = ~n6162 & ~n9517;
  assign n13830 = ~pi299 & ~n13829;
  assign n13831 = ~n13828 & n13830;
  assign n13832 = ~n13808 & ~n13831;
  assign n13833 = pi232 & ~n13832;
  assign n13834 = ~n6143 & ~n9515;
  assign n13835 = ~pi232 & ~n9513;
  assign n13836 = ~n13834 & n13835;
  assign n13837 = ~pi39 & ~n13836;
  assign n13838 = ~n13833 & n13837;
  assign n13839 = ~n13787 & ~n13838;
  assign n13840 = ~pi38 & ~n13839;
  assign n13841 = n13619 & ~n13840;
  assign n13842 = ~n13714 & ~n13716;
  assign n13843 = ~n13841 & n13842;
  assign n13844 = n3237 & ~n13843;
  assign n13845 = n8924 & ~n13725;
  assign n13846 = n3095 & n13845;
  assign n13847 = n13722 & ~n13846;
  assign n13848 = ~n13714 & ~n13847;
  assign n13849 = n9410 & ~n13848;
  assign n13850 = ~n13721 & ~n13849;
  assign n13851 = ~n13844 & n13850;
  assign n13852 = ~pi54 & ~n13851;
  assign n13853 = ~n13610 & ~n13852;
  assign n13854 = ~pi74 & ~n13853;
  assign n13855 = n13603 & ~n13854;
  assign n13856 = pi54 & n13582;
  assign n13857 = ~pi92 & n8948;
  assign n13858 = n8924 & n13857;
  assign n13859 = ~n13738 & n13858;
  assign n13860 = ~n13856 & n13859;
  assign n13861 = n3095 & n13860;
  assign n13862 = n13587 & ~n13861;
  assign n13863 = n13737 & ~n13862;
  assign n13864 = n3293 & ~n13863;
  assign n13865 = ~n13855 & n13864;
  assign n13866 = n13590 & ~n13865;
  assign n13867 = ~n13754 & ~n13866;
  assign n13868 = ~pi118 & n13867;
  assign n13869 = ~n13757 & ~n13868;
  assign n13870 = ~n13756 & n13869;
  assign n13871 = ~pi118 & ~n8935;
  assign n13872 = n13755 & n13871;
  assign n13873 = n13867 & ~n13871;
  assign n13874 = n13757 & ~n13873;
  assign n13875 = ~n13872 & n13874;
  assign po276 = n13870 | n13875;
  assign n13877 = pi128 & pi228;
  assign n13878 = ~n10109 & n13877;
  assign n13879 = ~n3052 & n3474;
  assign n13880 = n7509 & n13879;
  assign n13881 = ~n3329 & n5767;
  assign n13882 = n7513 & n13881;
  assign n13883 = ~n13880 & ~n13882;
  assign n13884 = pi39 & ~n13883;
  assign n13885 = n2579 & n10103;
  assign n13886 = n11600 & ~n13885;
  assign n13887 = n2592 & ~n13886;
  assign n13888 = ~pi97 & ~n13887;
  assign n13889 = ~pi46 & n2795;
  assign n13890 = n2758 & n13889;
  assign n13891 = ~n13888 & n13890;
  assign n13892 = pi299 & n6412;
  assign n13893 = ~n6378 & ~n13892;
  assign n13894 = n7462 & ~n13893;
  assign n13895 = pi109 & ~n13894;
  assign n13896 = ~n2795 & n11601;
  assign n13897 = ~n13895 & ~n13896;
  assign n13898 = ~n13891 & n13897;
  assign n13899 = ~n6301 & ~n13894;
  assign n13900 = ~n6382 & n13894;
  assign n13901 = ~n13899 & ~n13900;
  assign n13902 = ~n13898 & n13901;
  assign n13903 = ~pi91 & ~n13902;
  assign n13904 = n2536 & ~n6336;
  assign n13905 = ~n13903 & n13904;
  assign n13906 = ~n2563 & ~n13905;
  assign n13907 = ~pi39 & n11026;
  assign n13908 = ~n13906 & n13907;
  assign n13909 = ~n13884 & ~n13908;
  assign n13910 = ~pi38 & ~n13909;
  assign n13911 = ~pi228 & n13910;
  assign n13912 = ~n13877 & ~n13911;
  assign n13913 = ~pi100 & ~n13912;
  assign n13914 = n3181 & n3321;
  assign n13915 = ~n13877 & ~n13914;
  assign n13916 = pi100 & ~n13915;
  assign n13917 = ~pi87 & ~n13916;
  assign n13918 = ~n13913 & n13917;
  assign n13919 = pi87 & ~n13877;
  assign n13920 = ~pi75 & ~n13919;
  assign n13921 = ~n13918 & n13920;
  assign n13922 = n7336 & n8924;
  assign n13923 = ~n13877 & ~n13922;
  assign n13924 = pi75 & ~n13923;
  assign n13925 = ~pi92 & ~n13924;
  assign n13926 = ~n13921 & n13925;
  assign n13927 = pi92 & ~n13877;
  assign n13928 = ~n7349 & n13927;
  assign n13929 = n10109 & ~n13928;
  assign n13930 = ~n13926 & n13929;
  assign po277 = n13878 | n13930;
  assign n13932 = ~pi31 & ~pi80;
  assign n13933 = pi818 & n13932;
  assign n13934 = ~n7422 & n8021;
  assign n13935 = ~n7697 & ~n13934;
  assign n13936 = ~pi120 & ~n7422;
  assign n13937 = ~pi1093 & n13936;
  assign n13938 = n13935 & ~n13937;
  assign n13939 = n3095 & n7468;
  assign n13940 = pi120 & ~n8021;
  assign n13941 = ~n7528 & n13940;
  assign n13942 = n13939 & ~n13941;
  assign n13943 = ~pi120 & pi1093;
  assign n13944 = n7528 & ~n13943;
  assign n13945 = ~n13942 & ~n13944;
  assign n13946 = n3181 & n8064;
  assign n13947 = ~n13945 & n13946;
  assign n13948 = ~n8021 & n13943;
  assign n13949 = ~n13940 & ~n13948;
  assign n13950 = pi100 & ~n13949;
  assign n13951 = ~n13947 & n13950;
  assign n13952 = ~pi1093 & n7452;
  assign n13953 = pi120 & n13952;
  assign n13954 = ~pi39 & ~n13953;
  assign n13955 = n7492 & ~n10297;
  assign n13956 = n7443 & n7474;
  assign n13957 = ~pi829 & n13956;
  assign n13958 = ~pi122 & ~n13957;
  assign n13959 = ~n13955 & n13958;
  assign n13960 = pi122 & ~n7444;
  assign n13961 = ~n2733 & ~n13960;
  assign n13962 = ~n13959 & n13961;
  assign n13963 = n10018 & ~n13962;
  assign n13964 = ~pi122 & n7474;
  assign n13965 = n7536 & ~n13956;
  assign n13966 = ~n13964 & n13965;
  assign n13967 = ~n13963 & ~n13966;
  assign n13968 = n13954 & n13967;
  assign n13969 = n6192 & ~n13949;
  assign n13970 = ~n7508 & n13940;
  assign n13971 = pi1091 & pi1092;
  assign n13972 = n7506 & n13971;
  assign n13973 = n13948 & ~n13972;
  assign n13974 = ~n13970 & ~n13973;
  assign n13975 = ~n6192 & ~n13974;
  assign n13976 = ~n13969 & ~n13975;
  assign n13977 = ~n6215 & ~n13976;
  assign n13978 = ~n6198 & n13949;
  assign n13979 = n6198 & n13974;
  assign n13980 = ~n13978 & ~n13979;
  assign n13981 = n6215 & n13980;
  assign n13982 = n8050 & ~n13981;
  assign n13983 = ~n13977 & n13982;
  assign n13984 = ~n8050 & n13949;
  assign n13985 = ~pi299 & ~n13984;
  assign n13986 = ~n13983 & n13985;
  assign n13987 = ~n6189 & ~n13976;
  assign n13988 = n6189 & n13980;
  assign n13989 = n8039 & ~n13988;
  assign n13990 = ~n13987 & n13989;
  assign n13991 = ~n8039 & n13949;
  assign n13992 = pi299 & ~n13991;
  assign n13993 = ~n13990 & n13992;
  assign n13994 = pi39 & ~n13993;
  assign n13995 = ~n13986 & n13994;
  assign n13996 = ~n13968 & ~n13995;
  assign n13997 = ~pi38 & ~n13996;
  assign n13998 = pi38 & n8021;
  assign n13999 = ~pi120 & ~pi1093;
  assign n14000 = pi38 & n13999;
  assign n14001 = ~pi100 & ~n14000;
  assign n14002 = ~n13998 & n14001;
  assign n14003 = ~n13997 & n14002;
  assign n14004 = ~n13951 & ~n14003;
  assign n14005 = ~pi87 & ~n14004;
  assign n14006 = n7544 & ~n13999;
  assign n14007 = n7536 & ~n13964;
  assign n14008 = ~n8076 & n14007;
  assign n14009 = n7542 & ~n14008;
  assign n14010 = ~n3207 & n8021;
  assign n14011 = pi87 & ~n14010;
  assign n14012 = ~n14009 & n14011;
  assign n14013 = n14006 & n14012;
  assign n14014 = ~n14005 & ~n14013;
  assign n14015 = ~pi75 & ~n14014;
  assign n14016 = n7463 & n13949;
  assign n14017 = ~n7469 & n13948;
  assign n14018 = ~pi1091 & ~n8020;
  assign n14019 = ~n8013 & ~n14018;
  assign n14020 = pi120 & ~n14019;
  assign n14021 = ~n7463 & ~n14020;
  assign n14022 = ~n14017 & n14021;
  assign n14023 = ~n14016 & ~n14022;
  assign n14024 = n3222 & ~n14023;
  assign n14025 = ~n3222 & n13949;
  assign n14026 = pi75 & ~n14025;
  assign n14027 = ~n14024 & n14026;
  assign n14028 = n7422 & ~n14027;
  assign n14029 = ~n14015 & n14028;
  assign n14030 = n13938 & ~n14029;
  assign n14031 = ~n13963 & ~n13965;
  assign n14032 = n13954 & n14031;
  assign n14033 = pi1093 & ~n6198;
  assign n14034 = n6215 & n14033;
  assign n14035 = n6192 & ~n6215;
  assign n14036 = n8050 & ~n14035;
  assign n14037 = ~n14034 & n14036;
  assign n14038 = n7508 & n14037;
  assign n14039 = ~pi299 & ~n13999;
  assign n14040 = ~n14038 & n14039;
  assign n14041 = n6189 & n14033;
  assign n14042 = ~n6189 & n6192;
  assign n14043 = n8039 & ~n14042;
  assign n14044 = ~n14041 & n14043;
  assign n14045 = n7508 & n14044;
  assign n14046 = pi299 & ~n13999;
  assign n14047 = ~n14045 & n14046;
  assign n14048 = pi39 & ~n14047;
  assign n14049 = ~n14040 & n14048;
  assign n14050 = ~n14032 & ~n14049;
  assign n14051 = ~pi38 & ~n14050;
  assign n14052 = n14001 & ~n14051;
  assign n14053 = pi120 & n7528;
  assign n14054 = ~pi120 & n13939;
  assign n14055 = ~n14053 & ~n14054;
  assign n14056 = n13946 & ~n14055;
  assign n14057 = pi100 & ~n13999;
  assign n14058 = ~n14056 & n14057;
  assign n14059 = ~n14052 & ~n14058;
  assign n14060 = ~pi87 & ~n14059;
  assign n14061 = ~n14006 & ~n14060;
  assign n14062 = ~pi75 & ~n14061;
  assign n14063 = n7472 & ~n13999;
  assign n14064 = n7422 & ~n14063;
  assign n14065 = ~n14062 & n14064;
  assign n14066 = n7697 & ~n13937;
  assign n14067 = ~n14065 & n14066;
  assign n14068 = ~n14030 & ~n14067;
  assign n14069 = n13933 & ~n14068;
  assign n14070 = ~po1038 & ~n14069;
  assign n14071 = ~n7697 & n13949;
  assign n14072 = pi120 & ~n14071;
  assign n14073 = n13933 & ~n13999;
  assign n14074 = ~n14071 & n14073;
  assign n14075 = po1038 & ~n14074;
  assign n14076 = ~n14072 & n14075;
  assign n14077 = ~n8830 & ~n14076;
  assign n14078 = pi951 & pi982;
  assign n14079 = pi1092 & n14078;
  assign n14080 = pi1093 & n14079;
  assign n14081 = ~pi120 & ~n14080;
  assign n14082 = ~n14071 & ~n14081;
  assign n14083 = n14075 & ~n14082;
  assign n14084 = n8830 & ~n14083;
  assign n14085 = ~n14077 & ~n14084;
  assign n14086 = ~n14070 & ~n14085;
  assign n14087 = pi120 & n7470;
  assign n14088 = ~pi1091 & n14080;
  assign n14089 = ~pi120 & ~n14088;
  assign n14090 = n10018 & n14079;
  assign n14091 = ~pi93 & ~pi122;
  assign n14092 = n2549 & n14091;
  assign n14093 = n2753 & n8854;
  assign n14094 = n14092 & n14093;
  assign n14095 = n2535 & n14094;
  assign n14096 = n10255 & n14095;
  assign n14097 = n7466 & n14096;
  assign n14098 = n2492 & n14097;
  assign n14099 = n14090 & ~n14098;
  assign n14100 = n14089 & ~n14099;
  assign n14101 = ~n14087 & ~n14100;
  assign n14102 = ~n7463 & ~n14101;
  assign n14103 = n7463 & n14081;
  assign n14104 = n3222 & ~n14103;
  assign n14105 = ~n14102 & n14104;
  assign n14106 = ~n3222 & ~n14081;
  assign n14107 = pi75 & ~n14106;
  assign n14108 = ~n14105 & n14107;
  assign n14109 = pi950 & n3095;
  assign n14110 = n7448 & n7466;
  assign n14111 = n14109 & n14110;
  assign n14112 = n14090 & ~n14111;
  assign n14113 = n14089 & ~n14112;
  assign n14114 = ~n14053 & ~n14113;
  assign n14115 = ~pi39 & n8064;
  assign n14116 = ~n14114 & n14115;
  assign n14117 = pi100 & ~n14116;
  assign n14118 = ~pi38 & ~n14117;
  assign n14119 = ~n13946 & n14081;
  assign n14120 = ~n14118 & ~n14119;
  assign n14121 = ~n8050 & n14081;
  assign n14122 = ~pi299 & ~n14121;
  assign n14123 = ~n8238 & ~n14081;
  assign n14124 = n6215 & n14123;
  assign n14125 = ~n8234 & ~n14081;
  assign n14126 = ~n6215 & n14125;
  assign n14127 = n8050 & ~n14126;
  assign n14128 = ~n14124 & n14127;
  assign n14129 = n14122 & ~n14128;
  assign n14130 = ~n8039 & n14081;
  assign n14131 = pi299 & ~n14130;
  assign n14132 = n6189 & n14123;
  assign n14133 = ~n6189 & n14125;
  assign n14134 = n8039 & ~n14133;
  assign n14135 = ~n14132 & n14134;
  assign n14136 = n14131 & ~n14135;
  assign n14137 = ~n14129 & ~n14136;
  assign n14138 = pi39 & ~n14137;
  assign n14139 = ~n13952 & n14031;
  assign n14140 = pi120 & n14139;
  assign n14141 = n2580 & n7432;
  assign n14142 = n2576 & n14141;
  assign n14143 = ~pi97 & ~n14142;
  assign n14144 = n2761 & ~n14143;
  assign n14145 = n2759 & n14144;
  assign n14146 = ~n7479 & ~n14145;
  assign n14147 = n2518 & ~n14146;
  assign n14148 = n7426 & ~n14147;
  assign n14149 = n7423 & ~n14148;
  assign n14150 = ~pi51 & ~n14149;
  assign n14151 = ~n2558 & ~n14150;
  assign n14152 = ~pi96 & ~n14151;
  assign n14153 = ~pi72 & pi950;
  assign n14154 = n10298 & n14153;
  assign n14155 = ~n14152 & n14154;
  assign n14156 = n7448 & n14079;
  assign n14157 = ~n14155 & n14156;
  assign n14158 = n9505 & n14142;
  assign n14159 = n7423 & n14158;
  assign n14160 = n7428 & ~n14159;
  assign n14161 = pi950 & n7475;
  assign n14162 = ~n14160 & n14161;
  assign n14163 = pi824 & n14162;
  assign n14164 = n14079 & ~n14163;
  assign n14165 = ~pi829 & n14164;
  assign n14166 = pi829 & pi1092;
  assign n14167 = pi122 & n14078;
  assign n14168 = n14166 & n14167;
  assign n14169 = ~n14162 & n14168;
  assign n14170 = ~n14165 & ~n14169;
  assign n14171 = ~n14157 & n14170;
  assign n14172 = n7473 & ~n14171;
  assign n14173 = n2733 & n14080;
  assign n14174 = ~n14172 & ~n14173;
  assign n14175 = pi1091 & ~n14174;
  assign n14176 = n14088 & ~n14163;
  assign n14177 = ~pi120 & ~n14176;
  assign n14178 = ~n14175 & n14177;
  assign n14179 = ~pi39 & ~n14178;
  assign n14180 = ~n14140 & n14179;
  assign n14181 = ~n14138 & ~n14180;
  assign n14182 = n3206 & ~n14181;
  assign n14183 = ~n14120 & ~n14182;
  assign n14184 = ~pi87 & ~n14183;
  assign n14185 = ~n3207 & n14081;
  assign n14186 = pi87 & ~n14185;
  assign n14187 = ~n2733 & ~n6171;
  assign n14188 = n14109 & n14187;
  assign n14189 = n14090 & ~n14188;
  assign n14190 = pi824 & n14109;
  assign n14191 = n14088 & ~n14190;
  assign n14192 = ~n14189 & ~n14191;
  assign n14193 = ~pi120 & ~n14192;
  assign n14194 = ~n7537 & ~n7541;
  assign n14195 = pi120 & ~n14194;
  assign n14196 = n3207 & ~n14195;
  assign n14197 = ~n14193 & n14196;
  assign n14198 = n14186 & ~n14197;
  assign n14199 = ~pi75 & ~n14198;
  assign n14200 = ~n14184 & n14199;
  assign n14201 = ~n14108 & ~n14200;
  assign n14202 = n7422 & ~n14201;
  assign n14203 = n7697 & ~n14202;
  assign n14204 = ~n13964 & n14088;
  assign n14205 = ~n14112 & ~n14204;
  assign n14206 = ~pi120 & ~n14205;
  assign n14207 = ~n13941 & ~n14206;
  assign n14208 = n8064 & ~n14207;
  assign n14209 = ~n13949 & ~n14081;
  assign n14210 = ~n8064 & n14209;
  assign n14211 = n3181 & ~n14210;
  assign n14212 = ~n14208 & n14211;
  assign n14213 = ~n3181 & ~n14209;
  assign n14214 = pi100 & ~n14213;
  assign n14215 = ~n14212 & n14214;
  assign n14216 = ~n13952 & n13967;
  assign n14217 = pi120 & n14216;
  assign n14218 = n14007 & n14164;
  assign n14219 = ~pi120 & ~n14218;
  assign n14220 = ~n14175 & n14219;
  assign n14221 = ~n14217 & ~n14220;
  assign n14222 = ~pi39 & ~n14221;
  assign n14223 = ~n7506 & n14090;
  assign n14224 = ~n14204 & ~n14223;
  assign n14225 = ~pi120 & ~n14224;
  assign n14226 = ~n13970 & ~n14225;
  assign n14227 = ~n6192 & ~n14226;
  assign n14228 = n6192 & n14209;
  assign n14229 = ~n14227 & ~n14228;
  assign n14230 = ~n6189 & ~n14229;
  assign n14231 = n6198 & ~n14226;
  assign n14232 = ~n6198 & n14209;
  assign n14233 = ~n14231 & ~n14232;
  assign n14234 = n6189 & ~n14233;
  assign n14235 = n8039 & ~n14234;
  assign n14236 = ~n14230 & n14235;
  assign n14237 = n8021 & ~n8039;
  assign n14238 = n14131 & ~n14237;
  assign n14239 = ~n14236 & n14238;
  assign n14240 = ~n6215 & ~n14229;
  assign n14241 = n6215 & ~n14233;
  assign n14242 = n8050 & ~n14241;
  assign n14243 = ~n14240 & n14242;
  assign n14244 = ~n13984 & n14122;
  assign n14245 = ~n14243 & n14244;
  assign n14246 = pi39 & ~n14245;
  assign n14247 = ~n14239 & n14246;
  assign n14248 = ~n14222 & ~n14247;
  assign n14249 = ~pi38 & ~n14248;
  assign n14250 = pi38 & ~n14209;
  assign n14251 = ~pi100 & ~n14250;
  assign n14252 = ~n14249 & n14251;
  assign n14253 = ~n14215 & ~n14252;
  assign n14254 = ~pi87 & ~n14253;
  assign n14255 = ~n14009 & ~n14196;
  assign n14256 = ~n14189 & ~n14204;
  assign n14257 = n14193 & ~n14256;
  assign n14258 = ~n14255 & ~n14257;
  assign n14259 = ~n14010 & n14186;
  assign n14260 = ~n14258 & n14259;
  assign n14261 = ~n14254 & ~n14260;
  assign n14262 = ~pi75 & ~n14261;
  assign n14263 = n7463 & ~n14209;
  assign n14264 = ~n14099 & ~n14204;
  assign n14265 = ~pi120 & ~n14264;
  assign n14266 = n14021 & ~n14265;
  assign n14267 = ~n14263 & ~n14266;
  assign n14268 = n3222 & ~n14267;
  assign n14269 = ~n3222 & ~n14209;
  assign n14270 = pi75 & ~n14269;
  assign n14271 = ~n14268 & n14270;
  assign n14272 = n7422 & ~n14271;
  assign n14273 = ~n14262 & n14272;
  assign n14274 = n13938 & ~n14273;
  assign n14275 = ~n14203 & ~n14274;
  assign n14276 = n13936 & ~n14080;
  assign n14277 = n14084 & ~n14276;
  assign n14278 = ~n14275 & n14277;
  assign n14279 = ~pi39 & ~n14139;
  assign n14280 = n7518 & ~n14279;
  assign n14281 = ~pi100 & ~n14280;
  assign n14282 = ~n7532 & ~n14281;
  assign n14283 = ~pi87 & ~n14282;
  assign n14284 = ~n7544 & ~n14283;
  assign n14285 = ~pi75 & ~n14284;
  assign n14286 = ~n7472 & ~n14285;
  assign n14287 = n7697 & ~n13936;
  assign n14288 = ~n14286 & n14287;
  assign n14289 = n7532 & ~n8021;
  assign n14290 = ~pi39 & ~n14216;
  assign n14291 = ~n8021 & ~n8234;
  assign n14292 = ~n6215 & n14291;
  assign n14293 = ~n8021 & ~n8238;
  assign n14294 = n6215 & n14293;
  assign n14295 = n8050 & ~n14294;
  assign n14296 = ~n14292 & n14295;
  assign n14297 = n8021 & ~n8050;
  assign n14298 = ~pi299 & ~n14297;
  assign n14299 = ~n14296 & n14298;
  assign n14300 = ~n6189 & n14291;
  assign n14301 = n6189 & n14293;
  assign n14302 = n8039 & ~n14301;
  assign n14303 = ~n14300 & n14302;
  assign n14304 = pi299 & ~n14237;
  assign n14305 = ~n14303 & n14304;
  assign n14306 = ~n14299 & ~n14305;
  assign n14307 = pi39 & ~n14306;
  assign n14308 = ~pi38 & ~n14307;
  assign n14309 = ~n14290 & n14308;
  assign n14310 = ~pi100 & ~n13998;
  assign n14311 = ~n14309 & n14310;
  assign n14312 = ~n14289 & ~n14311;
  assign n14313 = ~pi87 & ~n14312;
  assign n14314 = ~n14012 & ~n14313;
  assign n14315 = ~pi75 & ~n14314;
  assign n14316 = n7464 & n14019;
  assign n14317 = ~n7464 & n8021;
  assign n14318 = pi75 & ~n14317;
  assign n14319 = ~n14316 & n14318;
  assign n14320 = ~n14315 & ~n14319;
  assign n14321 = n13935 & ~n14320;
  assign n14322 = ~n7422 & ~n14071;
  assign n14323 = ~n14321 & ~n14322;
  assign n14324 = ~n14288 & n14323;
  assign n14325 = pi120 & n14077;
  assign n14326 = ~n14324 & n14325;
  assign n14327 = ~n14278 & ~n14326;
  assign n14328 = ~n13933 & ~n14327;
  assign po278 = n14086 | n14328;
  assign n14330 = n2467 & n10099;
  assign n14331 = ~pi51 & n14330;
  assign n14332 = n6162 & ~n14331;
  assign n14333 = pi51 & pi146;
  assign n14334 = pi51 & n6162;
  assign n14335 = ~pi146 & n14334;
  assign n14336 = pi161 & ~n14335;
  assign n14337 = ~n14333 & ~n14336;
  assign n14338 = n14332 & n14337;
  assign n14339 = ~pi87 & ~n14338;
  assign n14340 = pi87 & ~n13573;
  assign n14341 = pi232 & ~n14340;
  assign n14342 = ~n14339 & n14341;
  assign n14343 = ~pi134 & ~pi135;
  assign n14344 = ~pi136 & n14343;
  assign n14345 = ~pi130 & n14344;
  assign n14346 = ~pi132 & n14345;
  assign n14347 = ~pi126 & n14346;
  assign n14348 = ~pi121 & n14347;
  assign n14349 = ~pi125 & ~pi133;
  assign n14350 = pi121 & ~n14349;
  assign n14351 = ~pi121 & n14349;
  assign n14352 = ~n14350 & ~n14351;
  assign n14353 = ~n14348 & ~n14352;
  assign n14354 = ~pi87 & n14331;
  assign n14355 = ~n14353 & n14354;
  assign n14356 = po1038 & ~n14355;
  assign n14357 = ~n14342 & n14356;
  assign n14358 = pi299 & ~n14338;
  assign n14359 = ~pi142 & n14334;
  assign n14360 = pi144 & ~n14359;
  assign n14361 = pi51 & pi142;
  assign n14362 = n14332 & ~n14361;
  assign n14363 = ~n14360 & n14362;
  assign n14364 = ~pi299 & ~n14363;
  assign n14365 = pi232 & ~n14364;
  assign n14366 = ~n14358 & n14365;
  assign n14367 = pi38 & ~n14366;
  assign n14368 = ~pi100 & ~n14367;
  assign n14369 = pi38 & ~n14331;
  assign n14370 = ~pi100 & ~n14369;
  assign n14371 = ~n14368 & ~n14370;
  assign n14372 = n2456 & n10098;
  assign n14373 = n12966 & n14372;
  assign n14374 = ~pi50 & pi77;
  assign n14375 = n2484 & n14374;
  assign n14376 = n14373 & n14375;
  assign n14377 = n2494 & n7437;
  assign n14378 = ~pi24 & pi314;
  assign n14379 = n14377 & n14378;
  assign n14380 = n8859 & n14379;
  assign n14381 = n14376 & n14380;
  assign n14382 = n3093 & n14381;
  assign n14383 = n2579 & n14373;
  assign n14384 = ~pi58 & n14377;
  assign n14385 = n9003 & n14384;
  assign n14386 = n14383 & n14385;
  assign n14387 = pi72 & n6360;
  assign n14388 = n14386 & n14387;
  assign n14389 = pi86 & n14383;
  assign n14390 = ~n14376 & ~n14389;
  assign n14391 = n11016 & ~n14390;
  assign n14392 = ~pi24 & n11604;
  assign n14393 = n14383 & n14392;
  assign n14394 = n14330 & ~n14393;
  assign n14395 = ~n14391 & n14394;
  assign n14396 = ~pi51 & ~n14330;
  assign n14397 = ~n2497 & ~n14396;
  assign n14398 = ~n14395 & ~n14397;
  assign n14399 = n3093 & n14398;
  assign n14400 = n14331 & ~n14399;
  assign n14401 = ~n14388 & n14400;
  assign n14402 = ~n14382 & n14401;
  assign n14403 = ~n6162 & ~n14402;
  assign n14404 = pi72 & n10382;
  assign n14405 = ~n14334 & ~n14404;
  assign n14406 = n6162 & ~n14405;
  assign n14407 = ~n14403 & ~n14406;
  assign n14408 = ~pi51 & n14379;
  assign n14409 = n13355 & n14408;
  assign n14410 = n3093 & n6162;
  assign n14411 = n14409 & n14410;
  assign n14412 = n14407 & ~n14411;
  assign n14413 = pi142 & n14412;
  assign n14414 = ~n6162 & n14402;
  assign n14415 = ~pi72 & ~n14409;
  assign n14416 = n6361 & ~n14415;
  assign n14417 = n6162 & ~n14416;
  assign n14418 = ~n14414 & ~n14417;
  assign n14419 = ~pi142 & ~n14418;
  assign n14420 = ~pi144 & ~n14419;
  assign n14421 = ~n14413 & n14420;
  assign n14422 = n14331 & ~n14382;
  assign n14423 = ~n14399 & n14422;
  assign n14424 = ~n6162 & ~n14423;
  assign n14425 = ~n14332 & ~n14424;
  assign n14426 = ~n14388 & n14425;
  assign n14427 = ~n14382 & n14426;
  assign n14428 = n14360 & ~n14427;
  assign n14429 = ~pi180 & ~n14428;
  assign n14430 = ~n14421 & n14429;
  assign n14431 = pi144 & ~n14426;
  assign n14432 = ~pi144 & ~n14407;
  assign n14433 = ~n14431 & ~n14432;
  assign n14434 = ~n14359 & ~n14433;
  assign n14435 = pi180 & ~n14434;
  assign n14436 = pi179 & ~n14435;
  assign n14437 = ~n14430 & n14436;
  assign n14438 = ~pi24 & ~n11605;
  assign n14439 = pi24 & ~n11602;
  assign n14440 = ~n14438 & ~n14439;
  assign n14441 = ~pi314 & ~n14440;
  assign n14442 = pi314 & ~n11602;
  assign n14443 = ~n14441 & ~n14442;
  assign n14444 = n2497 & n14443;
  assign n14445 = ~pi72 & ~n14444;
  assign n14446 = n6361 & ~n14445;
  assign n14447 = n6162 & ~n14446;
  assign n14448 = ~n14414 & ~n14447;
  assign n14449 = ~pi142 & ~n14448;
  assign n14450 = n7437 & n8919;
  assign n14451 = n14443 & n14450;
  assign n14452 = ~pi51 & ~n14451;
  assign n14453 = ~n14404 & n14452;
  assign n14454 = n6162 & ~n14453;
  assign n14455 = ~n14403 & ~n14454;
  assign n14456 = pi142 & n14455;
  assign n14457 = ~pi144 & ~n14456;
  assign n14458 = ~n14449 & n14457;
  assign n14459 = n14360 & ~n14402;
  assign n14460 = ~pi180 & ~n14459;
  assign n14461 = ~n14458 & n14460;
  assign n14462 = n2497 & n14440;
  assign n14463 = ~pi72 & ~n14462;
  assign n14464 = n6361 & ~n14463;
  assign n14465 = n6162 & ~n14464;
  assign n14466 = ~n14414 & ~n14465;
  assign n14467 = ~pi142 & ~n14466;
  assign n14468 = n14410 & n14462;
  assign n14469 = ~n14406 & ~n14468;
  assign n14470 = ~n14403 & n14469;
  assign n14471 = pi142 & n14470;
  assign n14472 = ~pi144 & ~n14471;
  assign n14473 = ~n14467 & n14472;
  assign n14474 = ~pi51 & n6162;
  assign n14475 = ~n14401 & n14474;
  assign n14476 = ~n14403 & ~n14475;
  assign n14477 = n6162 & ~n14400;
  assign n14478 = ~pi142 & ~n14477;
  assign n14479 = n6162 & n14396;
  assign n14480 = ~n14410 & ~n14479;
  assign n14481 = n3093 & ~n14398;
  assign n14482 = ~n14480 & ~n14481;
  assign n14483 = pi142 & ~n14482;
  assign n14484 = ~n14478 & ~n14483;
  assign n14485 = ~n14425 & ~n14484;
  assign n14486 = n14476 & ~n14485;
  assign n14487 = pi144 & ~n14486;
  assign n14488 = pi180 & ~n14487;
  assign n14489 = ~n14473 & n14488;
  assign n14490 = ~pi179 & ~n14489;
  assign n14491 = ~n14461 & n14490;
  assign n14492 = ~n14437 & ~n14491;
  assign n14493 = ~pi299 & ~n14492;
  assign n14494 = ~pi161 & ~n14335;
  assign n14495 = ~n14407 & n14494;
  assign n14496 = n14336 & ~n14426;
  assign n14497 = ~n14495 & ~n14496;
  assign n14498 = n9317 & ~n14497;
  assign n14499 = pi146 & n14412;
  assign n14500 = ~pi146 & ~n14418;
  assign n14501 = ~pi161 & ~n14500;
  assign n14502 = ~n14499 & n14501;
  assign n14503 = n14336 & ~n14427;
  assign n14504 = ~n14502 & ~n14503;
  assign n14505 = n9363 & ~n14504;
  assign n14506 = ~n14498 & ~n14505;
  assign n14507 = pi156 & ~n14506;
  assign n14508 = pi146 & n14455;
  assign n14509 = ~pi146 & ~n14448;
  assign n14510 = n9363 & ~n14509;
  assign n14511 = ~n14508 & n14510;
  assign n14512 = ~pi146 & ~n14466;
  assign n14513 = pi146 & n14470;
  assign n14514 = n9317 & ~n14513;
  assign n14515 = ~n14512 & n14514;
  assign n14516 = ~pi161 & ~n14515;
  assign n14517 = ~n14511 & n14516;
  assign n14518 = ~pi146 & ~n14477;
  assign n14519 = pi146 & ~n14482;
  assign n14520 = ~n14518 & ~n14519;
  assign n14521 = ~n14425 & ~n14520;
  assign n14522 = n14476 & ~n14521;
  assign n14523 = n9317 & ~n14522;
  assign n14524 = n9363 & ~n14335;
  assign n14525 = ~n14402 & n14524;
  assign n14526 = pi161 & ~n14525;
  assign n14527 = ~n14523 & n14526;
  assign n14528 = ~pi156 & ~n14527;
  assign n14529 = ~n14517 & n14528;
  assign n14530 = ~n14507 & ~n14529;
  assign n14531 = ~n14493 & n14530;
  assign n14532 = n9563 & ~n14531;
  assign n14533 = n3093 & n14386;
  assign n14534 = n14331 & ~n14533;
  assign n14535 = ~n14335 & ~n14534;
  assign n14536 = pi161 & ~n14535;
  assign n14537 = ~n6162 & ~n14534;
  assign n14538 = n2557 & n7442;
  assign n14539 = ~pi51 & ~n14538;
  assign n14540 = n6162 & ~n14539;
  assign n14541 = ~n14537 & ~n14540;
  assign n14542 = pi146 & ~n14541;
  assign n14543 = ~n6180 & ~n14537;
  assign n14544 = ~pi146 & ~n14543;
  assign n14545 = ~pi161 & ~n14544;
  assign n14546 = ~n14542 & n14545;
  assign n14547 = ~n14536 & ~n14546;
  assign n14548 = n6434 & ~n14547;
  assign n14549 = ~n9028 & ~n14548;
  assign n14550 = ~pi287 & n6162;
  assign n14551 = ~pi51 & n14550;
  assign n14552 = ~n14541 & ~n14551;
  assign n14553 = n14494 & n14552;
  assign n14554 = n14533 & ~n14550;
  assign n14555 = n14331 & ~n14554;
  assign n14556 = n14336 & ~n14555;
  assign n14557 = ~n14553 & ~n14556;
  assign n14558 = pi216 & ~n14557;
  assign n14559 = ~n14549 & ~n14558;
  assign n14560 = ~n14331 & ~n14338;
  assign n14561 = ~n6434 & ~n14560;
  assign n14562 = n9790 & ~n14561;
  assign n14563 = ~n14559 & n14562;
  assign n14564 = pi142 & ~n14541;
  assign n14565 = ~pi142 & ~n14543;
  assign n14566 = n6461 & ~n14565;
  assign n14567 = ~n14564 & n14566;
  assign n14568 = ~n9017 & ~n14567;
  assign n14569 = pi224 & ~n14359;
  assign n14570 = n14552 & n14569;
  assign n14571 = ~n14568 & ~n14570;
  assign n14572 = ~n14331 & ~n14359;
  assign n14573 = ~n6461 & ~n14572;
  assign n14574 = pi144 & ~n14573;
  assign n14575 = ~n6461 & n14479;
  assign n14576 = ~n14573 & ~n14575;
  assign n14577 = ~n14574 & n14576;
  assign n14578 = ~n14571 & n14577;
  assign n14579 = ~pi51 & ~n14534;
  assign n14580 = ~pi287 & ~n14579;
  assign n14581 = ~n14479 & ~n14550;
  assign n14582 = ~n14580 & ~n14581;
  assign n14583 = ~n14362 & ~n14582;
  assign n14584 = n9017 & ~n14583;
  assign n14585 = n14330 & n14584;
  assign n14586 = pi51 & ~n6162;
  assign n14587 = ~n14579 & ~n14586;
  assign n14588 = n6461 & ~n14361;
  assign n14589 = n14587 & n14588;
  assign n14590 = n14574 & ~n14589;
  assign n14591 = ~n14585 & n14590;
  assign n14592 = pi181 & ~n14591;
  assign n14593 = ~n14578 & n14592;
  assign n14594 = ~n14567 & n14577;
  assign n14595 = ~pi181 & ~n14590;
  assign n14596 = ~n14594 & n14595;
  assign n14597 = ~pi299 & ~n14596;
  assign n14598 = ~n14593 & n14597;
  assign n14599 = n9752 & ~n14561;
  assign n14600 = ~n14548 & n14599;
  assign n14601 = pi232 & ~n14600;
  assign n14602 = ~n14598 & n14601;
  assign n14603 = ~n14563 & n14602;
  assign n14604 = ~n6587 & ~n7510;
  assign n14605 = n14533 & ~n14604;
  assign n14606 = ~pi232 & n14331;
  assign n14607 = ~n14605 & n14606;
  assign n14608 = pi39 & ~n14607;
  assign n14609 = ~n14603 & n14608;
  assign n14610 = ~pi39 & ~pi232;
  assign n14611 = ~n14402 & n14610;
  assign n14612 = ~n14609 & ~n14611;
  assign n14613 = ~n14532 & n14612;
  assign n14614 = ~pi38 & ~n14613;
  assign n14615 = ~n14371 & ~n14614;
  assign n14616 = pi100 & n14331;
  assign n14617 = n3278 & ~n14616;
  assign n14618 = pi100 & n14366;
  assign n14619 = n14617 & ~n14618;
  assign n14620 = ~n14615 & n14619;
  assign n14621 = ~pi87 & ~n3266;
  assign n14622 = ~n14331 & n14621;
  assign n14623 = ~n14366 & n14622;
  assign n14624 = ~pi184 & ~pi299;
  assign n14625 = ~pi163 & pi299;
  assign n14626 = ~n14624 & ~n14625;
  assign n14627 = n7462 & n14626;
  assign n14628 = pi87 & ~n14627;
  assign n14629 = ~n14353 & ~n14628;
  assign n14630 = ~n14623 & n14629;
  assign n14631 = ~n14620 & n14630;
  assign n14632 = n6162 & ~n14452;
  assign n14633 = ~n14361 & n14632;
  assign n14634 = pi144 & ~n14633;
  assign n14635 = n14330 & ~n14381;
  assign n14636 = n14377 & n14635;
  assign n14637 = n14395 & n14636;
  assign n14638 = ~n14397 & ~n14637;
  assign n14639 = n3093 & ~n14638;
  assign n14640 = ~n14480 & ~n14639;
  assign n14641 = pi142 & n14640;
  assign n14642 = n6162 & ~n14423;
  assign n14643 = ~pi142 & n14642;
  assign n14644 = ~pi144 & ~n14643;
  assign n14645 = ~n14641 & n14644;
  assign n14646 = pi180 & ~n14645;
  assign n14647 = ~n14634 & n14646;
  assign n14648 = n14360 & ~n14468;
  assign n14649 = ~pi144 & ~n14484;
  assign n14650 = ~pi180 & ~n14649;
  assign n14651 = ~n14648 & n14650;
  assign n14652 = pi179 & ~n14651;
  assign n14653 = ~n14647 & n14652;
  assign n14654 = n14360 & ~n14411;
  assign n14655 = ~pi51 & ~n14635;
  assign n14656 = n3093 & ~n14655;
  assign n14657 = ~n14480 & ~n14656;
  assign n14658 = pi142 & n14657;
  assign n14659 = n6162 & ~n14422;
  assign n14660 = ~pi142 & n14659;
  assign n14661 = ~pi144 & ~n14660;
  assign n14662 = ~n14658 & n14661;
  assign n14663 = pi180 & ~n14662;
  assign n14664 = ~n14654 & n14663;
  assign n14665 = ~pi180 & n14363;
  assign n14666 = ~pi179 & ~n14665;
  assign n14667 = ~n14664 & n14666;
  assign n14668 = ~n14653 & ~n14667;
  assign n14669 = ~pi299 & ~n14668;
  assign n14670 = ~n14333 & n14632;
  assign n14671 = pi161 & ~n14670;
  assign n14672 = pi146 & n14640;
  assign n14673 = ~pi146 & n14642;
  assign n14674 = ~pi161 & ~n14673;
  assign n14675 = ~n14672 & n14674;
  assign n14676 = ~n14671 & ~n14675;
  assign n14677 = n9317 & ~n14676;
  assign n14678 = n14336 & ~n14468;
  assign n14679 = ~pi161 & ~n14520;
  assign n14680 = ~n14678 & ~n14679;
  assign n14681 = n9363 & ~n14680;
  assign n14682 = pi232 & ~n14681;
  assign n14683 = ~n14677 & n14682;
  assign n14684 = pi156 & ~n14683;
  assign n14685 = ~pi39 & ~n14684;
  assign n14686 = ~n14669 & n14685;
  assign n14687 = ~pi142 & ~n14538;
  assign n14688 = n9017 & n14550;
  assign n14689 = pi142 & ~n3095;
  assign n14690 = n14688 & ~n14689;
  assign n14691 = ~n14687 & n14690;
  assign n14692 = n14360 & ~n14691;
  assign n14693 = ~pi144 & ~n14362;
  assign n14694 = ~n14584 & n14693;
  assign n14695 = pi181 & ~n14694;
  assign n14696 = ~n14692 & n14695;
  assign n14697 = ~pi181 & n14363;
  assign n14698 = ~pi299 & ~n14697;
  assign n14699 = ~n14696 & n14698;
  assign n14700 = n6162 & n6435;
  assign n14701 = n14336 & ~n14700;
  assign n14702 = n14494 & ~n14582;
  assign n14703 = n9028 & ~n14702;
  assign n14704 = ~n14701 & n14703;
  assign n14705 = ~n9028 & n14338;
  assign n14706 = n9790 & ~n14705;
  assign n14707 = ~n14704 & n14706;
  assign n14708 = ~pi159 & n14358;
  assign n14709 = n10420 & ~n14708;
  assign n14710 = ~n14707 & n14709;
  assign n14711 = ~n14699 & n14710;
  assign n14712 = ~pi38 & ~n14711;
  assign n14713 = ~n14686 & n14712;
  assign n14714 = n14336 & ~n14411;
  assign n14715 = pi146 & n14657;
  assign n14716 = ~pi146 & n14659;
  assign n14717 = ~pi161 & ~n14716;
  assign n14718 = ~n14715 & n14717;
  assign n14719 = ~n14714 & ~n14718;
  assign n14720 = n9317 & ~n14719;
  assign n14721 = ~pi158 & n14358;
  assign n14722 = pi232 & ~n14721;
  assign n14723 = ~n14720 & n14722;
  assign n14724 = ~pi156 & n3181;
  assign n14725 = ~n14723 & n14724;
  assign n14726 = n14368 & ~n14725;
  assign n14727 = ~n14713 & n14726;
  assign n14728 = n3278 & ~n14618;
  assign n14729 = ~n14727 & n14728;
  assign n14730 = ~n14366 & n14621;
  assign n14731 = n14353 & ~n14628;
  assign n14732 = ~n14730 & n14731;
  assign n14733 = ~n14729 & n14732;
  assign n14734 = ~po1038 & ~n14733;
  assign n14735 = ~n14631 & n14734;
  assign po279 = n14357 | n14735;
  assign n14737 = n8021 & n8778;
  assign n14738 = n7422 & n14286;
  assign n14739 = n7697 & ~n14738;
  assign n14740 = n7422 & n14320;
  assign n14741 = n13935 & ~n14740;
  assign n14742 = ~po1038 & ~n14741;
  assign n14743 = ~n14739 & n14742;
  assign po280 = n14737 | n14743;
  assign n14745 = ~pi110 & n9012;
  assign n14746 = ~n6200 & n6434;
  assign n14747 = n14745 & n14746;
  assign n14748 = pi39 & ~n14747;
  assign n14749 = pi110 & n10020;
  assign n14750 = ~n10916 & n14749;
  assign n14751 = po1057 & n14750;
  assign n14752 = ~pi39 & ~n14751;
  assign n14753 = po1038 & ~n14752;
  assign n14754 = ~n14748 & n14753;
  assign n14755 = ~pi38 & n3267;
  assign n14756 = pi299 & n14747;
  assign n14757 = ~n6221 & n7510;
  assign n14758 = n14745 & n14757;
  assign n14759 = pi39 & ~n14758;
  assign n14760 = ~n14756 & n14759;
  assign n14761 = ~pi111 & ~n6307;
  assign n14762 = ~pi36 & n2637;
  assign n14763 = ~n14761 & n14762;
  assign n14764 = n2457 & ~n14763;
  assign n14765 = ~n2602 & ~n2646;
  assign n14766 = ~n14764 & n14765;
  assign n14767 = ~pi83 & ~n14766;
  assign n14768 = n2604 & ~n14767;
  assign n14769 = ~pi71 & ~n14768;
  assign n14770 = n6317 & ~n14769;
  assign n14771 = ~pi81 & ~n14770;
  assign n14772 = n11374 & ~n14771;
  assign n14773 = ~pi90 & ~n14772;
  assign n14774 = n2496 & ~n14773;
  assign n14775 = pi90 & ~n10349;
  assign n14776 = n9521 & ~n14775;
  assign n14777 = n14774 & n14776;
  assign n14778 = pi72 & n2497;
  assign n14779 = n10349 & n14778;
  assign n14780 = ~n14777 & ~n14779;
  assign n14781 = n6360 & ~n14780;
  assign n14782 = ~pi110 & ~n14781;
  assign n14783 = n13362 & ~n14782;
  assign n14784 = n2707 & n14774;
  assign n14785 = ~pi72 & ~n14784;
  assign n14786 = n6361 & ~n13362;
  assign n14787 = ~n14785 & n14786;
  assign n14788 = ~pi39 & ~n14787;
  assign n14789 = ~n14783 & n14788;
  assign n14790 = ~n14760 & ~n14789;
  assign n14791 = n14755 & ~n14790;
  assign n14792 = pi110 & n13362;
  assign n14793 = ~pi39 & ~n14792;
  assign n14794 = ~n14760 & ~n14793;
  assign n14795 = ~n14755 & ~n14794;
  assign n14796 = ~po1038 & ~n14795;
  assign n14797 = ~n14791 & n14796;
  assign po281 = ~n14754 & ~n14797;
  assign n14799 = ~pi125 & n14348;
  assign n14800 = pi125 & pi133;
  assign n14801 = ~n14349 & ~n14800;
  assign n14802 = ~n14799 & ~n14801;
  assign n14803 = n14331 & ~n14802;
  assign n14804 = pi172 & n14334;
  assign n14805 = ~pi152 & n14479;
  assign n14806 = ~n14804 & ~n14805;
  assign n14807 = pi232 & ~n14806;
  assign n14808 = ~n14803 & ~n14807;
  assign n14809 = ~pi87 & ~n14808;
  assign n14810 = pi87 & n7462;
  assign n14811 = pi162 & n14810;
  assign n14812 = po1038 & ~n14811;
  assign n14813 = ~n14809 & n14812;
  assign n14814 = ~pi152 & n6162;
  assign n14815 = n14404 & ~n14814;
  assign n14816 = n14330 & ~n14388;
  assign n14817 = n14474 & ~n14816;
  assign n14818 = ~pi152 & n14817;
  assign n14819 = ~pi197 & ~n14818;
  assign n14820 = ~n14815 & n14819;
  assign n14821 = n14474 & n14816;
  assign n14822 = ~n14382 & n14821;
  assign n14823 = ~n6162 & n14404;
  assign n14824 = ~n14474 & ~n14823;
  assign n14825 = ~n14822 & ~n14824;
  assign n14826 = ~pi152 & pi197;
  assign n14827 = ~n14825 & n14826;
  assign n14828 = ~n14820 & ~n14827;
  assign n14829 = ~n14804 & ~n14828;
  assign n14830 = ~n6162 & ~n14404;
  assign n14831 = ~n14417 & ~n14830;
  assign n14832 = ~pi172 & n14831;
  assign n14833 = ~n14334 & ~n14411;
  assign n14834 = ~n14404 & n14833;
  assign n14835 = pi172 & ~n14834;
  assign n14836 = pi152 & pi197;
  assign n14837 = ~n14835 & n14836;
  assign n14838 = ~n14832 & n14837;
  assign n14839 = ~n14829 & ~n14838;
  assign n14840 = n9825 & ~n14839;
  assign n14841 = ~n14447 & ~n14830;
  assign n14842 = ~pi172 & n14841;
  assign n14843 = ~n14453 & ~n14830;
  assign n14844 = pi172 & n14843;
  assign n14845 = pi152 & ~n14844;
  assign n14846 = ~n14842 & n14845;
  assign n14847 = n6162 & n14402;
  assign n14848 = ~n14824 & ~n14847;
  assign n14849 = ~pi152 & ~n14804;
  assign n14850 = ~n14848 & n14849;
  assign n14851 = pi197 & ~n14850;
  assign n14852 = ~n14846 & n14851;
  assign n14853 = ~n14465 & ~n14830;
  assign n14854 = pi152 & n14853;
  assign n14855 = ~n14475 & ~n14823;
  assign n14856 = ~pi152 & ~n14855;
  assign n14857 = ~pi172 & ~n14856;
  assign n14858 = ~n14854 & n14857;
  assign n14859 = n14405 & ~n14468;
  assign n14860 = pi152 & ~n14859;
  assign n14861 = n14401 & n14821;
  assign n14862 = ~n14830 & ~n14861;
  assign n14863 = ~pi152 & n14862;
  assign n14864 = pi172 & ~n14863;
  assign n14865 = ~n14860 & n14864;
  assign n14866 = ~pi197 & ~n14865;
  assign n14867 = ~n14858 & n14866;
  assign n14868 = n9831 & ~n14867;
  assign n14869 = ~n14852 & n14868;
  assign n14870 = ~n14840 & ~n14869;
  assign n14871 = pi299 & ~n14870;
  assign n14872 = pi145 & n14831;
  assign n14873 = ~pi145 & n14404;
  assign n14874 = pi174 & ~n14873;
  assign n14875 = ~n14872 & n14874;
  assign n14876 = pi145 & n14825;
  assign n14877 = ~n14817 & ~n14823;
  assign n14878 = ~pi145 & ~n14877;
  assign n14879 = ~pi174 & ~n14878;
  assign n14880 = ~n14876 & n14879;
  assign n14881 = ~n14875 & ~n14880;
  assign n14882 = ~pi193 & ~n14881;
  assign n14883 = ~pi145 & n14411;
  assign n14884 = ~n14833 & ~n14883;
  assign n14885 = ~n14404 & ~n14884;
  assign n14886 = pi174 & ~n14885;
  assign n14887 = ~n14334 & ~n14382;
  assign n14888 = pi145 & ~n14887;
  assign n14889 = n14821 & ~n14888;
  assign n14890 = ~pi174 & ~n14889;
  assign n14891 = ~n14830 & n14890;
  assign n14892 = pi193 & ~n14891;
  assign n14893 = ~n14886 & n14892;
  assign n14894 = ~n14882 & ~n14893;
  assign n14895 = n9809 & ~n14894;
  assign n14896 = pi145 & n14841;
  assign n14897 = ~pi145 & n14853;
  assign n14898 = ~pi193 & ~n14897;
  assign n14899 = ~n14896 & n14898;
  assign n14900 = pi145 & n14843;
  assign n14901 = ~pi145 & ~n14859;
  assign n14902 = pi193 & ~n14901;
  assign n14903 = ~n14900 & n14902;
  assign n14904 = pi174 & ~n14903;
  assign n14905 = ~n14899 & n14904;
  assign n14906 = pi193 & n14334;
  assign n14907 = pi145 & ~n14906;
  assign n14908 = ~n14848 & n14907;
  assign n14909 = ~pi174 & ~n14908;
  assign n14910 = ~pi145 & ~n14906;
  assign n14911 = n14855 & n14910;
  assign n14912 = n14909 & ~n14911;
  assign n14913 = n9815 & ~n14912;
  assign n14914 = ~n14905 & n14913;
  assign n14915 = ~n14895 & ~n14914;
  assign n14916 = ~pi38 & ~n14915;
  assign n14917 = ~n14871 & ~n14916;
  assign n14918 = n9563 & ~n14917;
  assign n14919 = ~n7511 & ~n7514;
  assign n14920 = n3095 & ~n14919;
  assign n14921 = ~pi232 & ~n14920;
  assign n14922 = pi39 & ~n14921;
  assign n14923 = n14538 & n14550;
  assign n14924 = ~n14334 & ~n14923;
  assign n14925 = pi224 & n14924;
  assign n14926 = n6461 & ~n14925;
  assign n14927 = n3095 & ~n6162;
  assign n14928 = ~n14540 & ~n14927;
  assign n14929 = n8050 & n14928;
  assign n14930 = n14926 & ~n14929;
  assign n14931 = ~n14334 & ~n14930;
  assign n14932 = pi174 & ~n14931;
  assign n14933 = n6162 & ~n14534;
  assign n14934 = ~n14927 & ~n14933;
  assign n14935 = n8050 & n14934;
  assign n14936 = n14533 & n14550;
  assign n14937 = pi224 & ~n14936;
  assign n14938 = n6461 & ~n14937;
  assign n14939 = ~n14332 & ~n14938;
  assign n14940 = ~n14935 & ~n14939;
  assign n14941 = ~pi174 & n14940;
  assign n14942 = pi193 & ~n14941;
  assign n14943 = ~n14932 & n14942;
  assign n14944 = n6162 & n14579;
  assign n14945 = ~n14927 & ~n14944;
  assign n14946 = ~pi224 & n14945;
  assign n14947 = pi224 & ~n14582;
  assign n14948 = n6461 & ~n14947;
  assign n14949 = ~n14946 & n14948;
  assign n14950 = ~n14575 & ~n14949;
  assign n14951 = ~pi174 & ~n14950;
  assign n14952 = ~n8050 & ~n14688;
  assign n14953 = n3095 & ~n14952;
  assign n14954 = pi174 & n14953;
  assign n14955 = ~pi193 & ~n14954;
  assign n14956 = ~n14951 & n14955;
  assign n14957 = pi180 & ~n14956;
  assign n14958 = ~n14943 & n14957;
  assign n14959 = ~n8050 & ~n14332;
  assign n14960 = ~n14945 & ~n14959;
  assign n14961 = ~pi174 & n14960;
  assign n14962 = n3095 & n8050;
  assign n14963 = pi174 & n14962;
  assign n14964 = ~n14906 & ~n14963;
  assign n14965 = ~n14961 & n14964;
  assign n14966 = ~pi180 & ~n14965;
  assign n14967 = ~pi299 & ~n14966;
  assign n14968 = ~n14958 & n14967;
  assign n14969 = ~n8039 & n14806;
  assign n14970 = ~pi152 & ~n14934;
  assign n14971 = pi152 & ~n14928;
  assign n14972 = ~n14970 & ~n14971;
  assign n14973 = pi51 & ~pi172;
  assign n14974 = ~n14972 & ~n14973;
  assign n14975 = ~pi216 & ~n14974;
  assign n14976 = n6434 & n14975;
  assign n14977 = ~n14969 & ~n14976;
  assign n14978 = n9363 & ~n14977;
  assign n14979 = pi152 & ~n14700;
  assign n14980 = ~pi152 & ~n14582;
  assign n14981 = ~pi172 & ~n14980;
  assign n14982 = ~n14979 & n14981;
  assign n14983 = pi152 & n14924;
  assign n14984 = ~n14332 & ~n14936;
  assign n14985 = ~pi152 & n14984;
  assign n14986 = pi172 & ~n14985;
  assign n14987 = ~n14983 & n14986;
  assign n14988 = pi216 & ~n14987;
  assign n14989 = ~n14982 & n14988;
  assign n14990 = n6434 & ~n14989;
  assign n14991 = ~n14975 & n14990;
  assign n14992 = ~n6434 & ~n14806;
  assign n14993 = n9317 & ~n14992;
  assign n14994 = ~n14991 & n14993;
  assign n14995 = ~n14978 & ~n14994;
  assign n14996 = ~n14968 & n14995;
  assign n14997 = pi232 & ~n14996;
  assign n14998 = n14922 & ~n14997;
  assign n14999 = ~pi232 & ~n14404;
  assign n15000 = ~pi39 & ~n14999;
  assign n15001 = ~pi38 & ~n15000;
  assign n15002 = ~n14998 & n15001;
  assign n15003 = pi299 & n14806;
  assign n15004 = ~pi174 & n14479;
  assign n15005 = ~pi299 & ~n14906;
  assign n15006 = ~n15004 & n15005;
  assign n15007 = pi232 & ~n15006;
  assign n15008 = ~n15003 & n15007;
  assign n15009 = pi38 & ~n15008;
  assign n15010 = ~pi100 & ~n15009;
  assign n15011 = ~n15002 & n15010;
  assign n15012 = ~n14918 & n15011;
  assign n15013 = pi100 & n15008;
  assign n15014 = n3278 & ~n15013;
  assign n15015 = ~n15012 & n15014;
  assign n15016 = n14621 & ~n15008;
  assign n15017 = pi140 & ~pi299;
  assign n15018 = pi162 & pi299;
  assign n15019 = ~n15017 & ~n15018;
  assign n15020 = n7462 & ~n15019;
  assign n15021 = pi87 & ~n15020;
  assign n15022 = n14802 & ~n15021;
  assign n15023 = ~n15016 & n15022;
  assign n15024 = ~n15015 & n15023;
  assign n15025 = ~pi145 & ~n14424;
  assign n15026 = ~n14632 & n15025;
  assign n15027 = ~n14424 & ~n14468;
  assign n15028 = pi145 & n15027;
  assign n15029 = ~pi51 & n15028;
  assign n15030 = ~pi174 & ~n15029;
  assign n15031 = ~n15026 & n15030;
  assign n15032 = ~pi145 & ~n14422;
  assign n15033 = ~n6162 & ~n14422;
  assign n15034 = ~n14332 & ~n15033;
  assign n15035 = ~n14399 & n15034;
  assign n15036 = ~n15032 & n15035;
  assign n15037 = pi174 & ~n15036;
  assign n15038 = ~pi193 & ~n15037;
  assign n15039 = ~n15031 & n15038;
  assign n15040 = n14410 & n14444;
  assign n15041 = ~n14424 & ~n15040;
  assign n15042 = ~pi145 & n15041;
  assign n15043 = ~pi174 & ~n15028;
  assign n15044 = ~n15042 & n15043;
  assign n15045 = n3093 & n15036;
  assign n15046 = ~n14424 & ~n14640;
  assign n15047 = pi174 & ~n15046;
  assign n15048 = ~n15045 & n15047;
  assign n15049 = pi193 & ~n15048;
  assign n15050 = ~n15044 & n15049;
  assign n15051 = n9809 & ~n15050;
  assign n15052 = ~n15039 & n15051;
  assign n15053 = ~n14334 & ~n14424;
  assign n15054 = ~pi174 & ~n14883;
  assign n15055 = pi145 & n14330;
  assign n15056 = ~n15054 & ~n15055;
  assign n15057 = n15053 & ~n15056;
  assign n15058 = ~n14424 & ~n14659;
  assign n15059 = pi174 & n15058;
  assign n15060 = ~n15057 & ~n15059;
  assign n15061 = ~pi193 & ~n15060;
  assign n15062 = pi145 & ~n14479;
  assign n15063 = ~pi145 & pi174;
  assign n15064 = ~n14657 & n15063;
  assign n15065 = ~n15062 & ~n15064;
  assign n15066 = ~n15054 & n15065;
  assign n15067 = pi193 & ~n14424;
  assign n15068 = ~n15066 & n15067;
  assign n15069 = n9815 & ~n15068;
  assign n15070 = ~n15061 & n15069;
  assign n15071 = ~n15052 & ~n15070;
  assign n15072 = ~pi38 & ~n15071;
  assign n15073 = ~pi152 & ~n15041;
  assign n15074 = pi152 & ~n15046;
  assign n15075 = pi172 & ~n15074;
  assign n15076 = ~n15073 & n15075;
  assign n15077 = ~pi152 & n14632;
  assign n15078 = ~n14423 & ~n14814;
  assign n15079 = ~pi172 & ~n15078;
  assign n15080 = ~n15077 & n15079;
  assign n15081 = ~n15076 & ~n15080;
  assign n15082 = ~pi197 & ~n15081;
  assign n15083 = ~pi152 & ~n15027;
  assign n15084 = ~n14424 & ~n14482;
  assign n15085 = pi172 & n15084;
  assign n15086 = ~pi172 & n15035;
  assign n15087 = pi152 & ~n15086;
  assign n15088 = ~n15085 & n15087;
  assign n15089 = ~pi172 & n14334;
  assign n15090 = pi197 & ~n15089;
  assign n15091 = ~n15088 & n15090;
  assign n15092 = ~n15083 & n15091;
  assign n15093 = pi299 & n9825;
  assign n15094 = ~n15092 & n15093;
  assign n15095 = ~n15082 & n15094;
  assign n15096 = ~n14411 & ~n14424;
  assign n15097 = ~pi152 & n15096;
  assign n15098 = ~n14334 & n15097;
  assign n15099 = pi152 & n15058;
  assign n15100 = ~pi172 & ~n15099;
  assign n15101 = ~n15098 & n15100;
  assign n15102 = ~n14424 & ~n14657;
  assign n15103 = pi152 & n15102;
  assign n15104 = pi172 & ~n15103;
  assign n15105 = ~n15097 & n15104;
  assign n15106 = ~pi197 & ~n15105;
  assign n15107 = ~n15101 & n15106;
  assign n15108 = ~pi172 & ~n14805;
  assign n15109 = ~n14425 & n15108;
  assign n15110 = pi152 & n14479;
  assign n15111 = ~n14424 & ~n15110;
  assign n15112 = pi172 & ~n15111;
  assign n15113 = pi197 & ~n15112;
  assign n15114 = ~n15109 & n15113;
  assign n15115 = pi299 & n9831;
  assign n15116 = ~n15114 & n15115;
  assign n15117 = ~n15107 & n15116;
  assign n15118 = ~n15095 & ~n15117;
  assign n15119 = ~n15072 & n15118;
  assign n15120 = n9563 & ~n15119;
  assign n15121 = ~n14370 & ~n15010;
  assign n15122 = ~n14331 & n14806;
  assign n15123 = ~n9028 & ~n15122;
  assign n15124 = ~pi152 & n14543;
  assign n15125 = pi152 & n14587;
  assign n15126 = pi172 & ~n15125;
  assign n15127 = ~n15124 & n15126;
  assign n15128 = ~n14534 & ~n14814;
  assign n15129 = ~pi152 & n14540;
  assign n15130 = ~n15128 & ~n15129;
  assign n15131 = ~pi172 & ~n15130;
  assign n15132 = n9028 & ~n15131;
  assign n15133 = ~n15127 & n15132;
  assign n15134 = n9363 & ~n15133;
  assign n15135 = n14552 & n14849;
  assign n15136 = pi152 & ~n14804;
  assign n15137 = ~n14555 & n15136;
  assign n15138 = n9028 & ~n15137;
  assign n15139 = ~n15135 & n15138;
  assign n15140 = n9317 & ~n15139;
  assign n15141 = ~n15134 & ~n15140;
  assign n15142 = ~n15123 & ~n15141;
  assign n15143 = ~n6162 & ~n14330;
  assign n15144 = ~n9017 & ~n15143;
  assign n15145 = ~n14586 & n15144;
  assign n15146 = n9017 & n14543;
  assign n15147 = ~n15145 & ~n15146;
  assign n15148 = ~pi174 & ~n15147;
  assign n15149 = n9017 & n14533;
  assign n15150 = n14331 & ~n15149;
  assign n15151 = ~n14334 & ~n15150;
  assign n15152 = pi174 & ~n15151;
  assign n15153 = ~pi180 & ~n15152;
  assign n15154 = ~n15148 & n15153;
  assign n15155 = n9017 & ~n14537;
  assign n15156 = ~n10488 & n15155;
  assign n15157 = ~n15145 & ~n15156;
  assign n15158 = ~pi174 & ~n15157;
  assign n15159 = ~pi51 & ~n14555;
  assign n15160 = n6162 & ~n15159;
  assign n15161 = ~n15150 & ~n15160;
  assign n15162 = pi174 & ~n15161;
  assign n15163 = pi180 & ~n15162;
  assign n15164 = ~n15158 & n15163;
  assign n15165 = pi193 & ~n15164;
  assign n15166 = ~n15154 & n15165;
  assign n15167 = n9017 & n14541;
  assign n15168 = ~pi51 & n15144;
  assign n15169 = ~n15167 & ~n15168;
  assign n15170 = pi180 & n14551;
  assign n15171 = ~pi174 & ~n15170;
  assign n15172 = n15169 & n15171;
  assign n15173 = pi180 & n14555;
  assign n15174 = pi174 & ~n15150;
  assign n15175 = ~n15173 & n15174;
  assign n15176 = ~pi193 & ~n15175;
  assign n15177 = ~n15172 & n15176;
  assign n15178 = ~pi299 & ~n15177;
  assign n15179 = ~n15166 & n15178;
  assign n15180 = ~n15142 & ~n15179;
  assign n15181 = pi232 & ~n15180;
  assign n15182 = ~pi299 & ~n15150;
  assign n15183 = n9028 & n14533;
  assign n15184 = n14331 & ~n15183;
  assign n15185 = pi299 & ~n15184;
  assign n15186 = ~n15182 & ~n15185;
  assign n15187 = ~pi232 & ~n15186;
  assign n15188 = pi39 & ~n15187;
  assign n15189 = ~n15181 & n15188;
  assign n15190 = ~pi232 & ~n14423;
  assign n15191 = ~pi39 & ~n15190;
  assign n15192 = ~pi38 & ~n15191;
  assign n15193 = ~n15189 & n15192;
  assign n15194 = ~n15121 & ~n15193;
  assign n15195 = ~n15120 & n15194;
  assign n15196 = n14617 & ~n15013;
  assign n15197 = ~n15195 & n15196;
  assign n15198 = n14622 & ~n15008;
  assign n15199 = ~n14802 & ~n15021;
  assign n15200 = ~n15198 & n15199;
  assign n15201 = ~n15197 & n15200;
  assign n15202 = ~po1038 & ~n15201;
  assign n15203 = ~n15024 & n15202;
  assign po282 = n14813 | n15203;
  assign n15205 = ~pi189 & n14848;
  assign n15206 = pi189 & n14841;
  assign n15207 = ~n15205 & ~n15206;
  assign n15208 = pi178 & ~n15207;
  assign n15209 = pi189 & ~n14831;
  assign n15210 = ~pi189 & ~n14825;
  assign n15211 = ~pi178 & ~n15210;
  assign n15212 = ~n15209 & n15211;
  assign n15213 = ~n15208 & ~n15212;
  assign n15214 = pi181 & ~n15213;
  assign n15215 = pi189 & n14853;
  assign n15216 = ~pi189 & ~n14855;
  assign n15217 = pi178 & ~n15216;
  assign n15218 = ~n15215 & n15217;
  assign n15219 = ~pi189 & ~n14877;
  assign n15220 = pi189 & n14404;
  assign n15221 = ~pi178 & ~n15220;
  assign n15222 = ~n14334 & n15221;
  assign n15223 = ~n15219 & n15222;
  assign n15224 = ~pi181 & ~n15223;
  assign n15225 = n14877 & n15221;
  assign n15226 = n15224 & ~n15225;
  assign n15227 = ~n15218 & n15226;
  assign n15228 = n11751 & ~n15227;
  assign n15229 = ~n15214 & n15228;
  assign n15230 = ~pi153 & n14841;
  assign n15231 = pi153 & n14843;
  assign n15232 = pi157 & ~n15231;
  assign n15233 = ~n15230 & n15232;
  assign n15234 = ~pi153 & n14831;
  assign n15235 = pi153 & ~n14834;
  assign n15236 = ~pi157 & ~n15235;
  assign n15237 = ~n15234 & n15236;
  assign n15238 = ~n15233 & ~n15237;
  assign n15239 = pi166 & ~n15238;
  assign n15240 = ~pi157 & n14825;
  assign n15241 = pi157 & n14848;
  assign n15242 = pi153 & n14334;
  assign n15243 = ~pi166 & ~n15242;
  assign n15244 = ~n15241 & n15243;
  assign n15245 = ~n15240 & n15244;
  assign n15246 = ~n15239 & ~n15245;
  assign n15247 = n9790 & ~n15246;
  assign n15248 = pi166 & ~n14859;
  assign n15249 = ~pi166 & n14862;
  assign n15250 = pi153 & ~n15249;
  assign n15251 = ~n15248 & n15250;
  assign n15252 = pi166 & n14853;
  assign n15253 = ~pi166 & ~n14855;
  assign n15254 = ~pi153 & ~n15253;
  assign n15255 = ~n15252 & n15254;
  assign n15256 = ~n15251 & ~n15255;
  assign n15257 = pi157 & ~n15256;
  assign n15258 = ~pi166 & ~n14877;
  assign n15259 = pi166 & n14404;
  assign n15260 = ~pi157 & ~n15242;
  assign n15261 = ~n15259 & n15260;
  assign n15262 = ~n15258 & n15261;
  assign n15263 = ~n15257 & ~n15262;
  assign n15264 = n9752 & ~n15263;
  assign n15265 = ~pi189 & n15053;
  assign n15266 = n14843 & ~n15265;
  assign n15267 = pi178 & ~n15205;
  assign n15268 = ~n15266 & n15267;
  assign n15269 = pi189 & n14834;
  assign n15270 = ~n14334 & n15210;
  assign n15271 = ~n15269 & ~n15270;
  assign n15272 = ~pi178 & ~n15271;
  assign n15273 = pi181 & ~n15272;
  assign n15274 = ~n15268 & n15273;
  assign n15275 = pi189 & ~n14859;
  assign n15276 = ~pi189 & n14862;
  assign n15277 = pi178 & ~n15276;
  assign n15278 = ~n15275 & n15277;
  assign n15279 = n15224 & ~n15278;
  assign n15280 = n11790 & ~n15279;
  assign n15281 = ~n15274 & n15280;
  assign n15282 = ~n15264 & ~n15281;
  assign n15283 = ~n15247 & n15282;
  assign n15284 = ~n15229 & n15283;
  assign n15285 = pi232 & ~n15284;
  assign n15286 = n15000 & ~n15285;
  assign n15287 = ~pi126 & n14351;
  assign n15288 = pi126 & ~n14351;
  assign n15289 = ~n15287 & ~n15288;
  assign n15290 = ~n14347 & ~n15289;
  assign n15291 = ~pi166 & ~n14934;
  assign n15292 = pi166 & ~n14928;
  assign n15293 = ~n15291 & ~n15292;
  assign n15294 = pi51 & ~pi153;
  assign n15295 = ~n15293 & ~n15294;
  assign n15296 = ~pi216 & ~n15295;
  assign n15297 = pi166 & ~n14924;
  assign n15298 = ~pi166 & ~n14984;
  assign n15299 = pi153 & ~n15298;
  assign n15300 = ~n15297 & n15299;
  assign n15301 = pi166 & n14700;
  assign n15302 = ~pi166 & n14582;
  assign n15303 = ~pi153 & ~n15302;
  assign n15304 = ~n15301 & n15303;
  assign n15305 = pi160 & ~n15304;
  assign n15306 = ~n15300 & n15305;
  assign n15307 = pi216 & ~n15306;
  assign n15308 = n6434 & ~n15307;
  assign n15309 = ~n15296 & n15308;
  assign n15310 = ~pi51 & ~n14479;
  assign n15311 = ~n10266 & ~n14330;
  assign n15312 = ~pi51 & ~n15311;
  assign n15313 = ~n15242 & ~n15312;
  assign n15314 = ~n15310 & ~n15313;
  assign n15315 = pi299 & ~n15314;
  assign n15316 = ~pi160 & pi216;
  assign n15317 = n6587 & ~n15316;
  assign n15318 = ~n15315 & ~n15317;
  assign n15319 = ~n15309 & ~n15318;
  assign n15320 = ~pi189 & n14960;
  assign n15321 = pi189 & n14962;
  assign n15322 = ~pi182 & ~n15321;
  assign n15323 = ~n15320 & n15322;
  assign n15324 = ~n14334 & n15323;
  assign n15325 = pi189 & ~n14931;
  assign n15326 = ~pi189 & n14940;
  assign n15327 = pi182 & ~n15326;
  assign n15328 = ~n15325 & n15327;
  assign n15329 = ~n15324 & ~n15328;
  assign n15330 = n11790 & ~n15329;
  assign n15331 = ~pi189 & ~n14950;
  assign n15332 = pi189 & n14953;
  assign n15333 = pi182 & ~n15332;
  assign n15334 = ~n15331 & n15333;
  assign n15335 = ~n15323 & ~n15334;
  assign n15336 = n11751 & ~n15335;
  assign n15337 = ~n15330 & ~n15336;
  assign n15338 = ~n15319 & n15337;
  assign n15339 = pi232 & ~n15338;
  assign n15340 = n14922 & ~n15339;
  assign n15341 = n15290 & ~n15340;
  assign n15342 = ~n15286 & n15341;
  assign n15343 = ~pi166 & ~n15041;
  assign n15344 = pi166 & ~n15046;
  assign n15345 = pi153 & ~n15344;
  assign n15346 = ~n15343 & n15345;
  assign n15347 = ~pi166 & n14632;
  assign n15348 = ~n10266 & ~n14423;
  assign n15349 = ~pi153 & ~n15348;
  assign n15350 = ~n15347 & n15349;
  assign n15351 = ~n15346 & ~n15350;
  assign n15352 = ~pi157 & ~n15351;
  assign n15353 = pi51 & n10266;
  assign n15354 = pi166 & ~n15058;
  assign n15355 = ~n15353 & ~n15354;
  assign n15356 = ~pi153 & ~n15355;
  assign n15357 = ~pi166 & ~n15096;
  assign n15358 = pi153 & pi166;
  assign n15359 = ~n15102 & n15358;
  assign n15360 = pi157 & ~n15359;
  assign n15361 = ~n15357 & n15360;
  assign n15362 = ~n15356 & n15361;
  assign n15363 = n9752 & ~n15362;
  assign n15364 = ~n15352 & n15363;
  assign n15365 = ~n10270 & ~n14423;
  assign n15366 = ~pi189 & n14632;
  assign n15367 = ~n15365 & ~n15366;
  assign n15368 = ~pi178 & ~n15367;
  assign n15369 = pi189 & n15058;
  assign n15370 = pi178 & ~n15265;
  assign n15371 = ~pi189 & n15096;
  assign n15372 = pi178 & ~n15371;
  assign n15373 = ~n15370 & ~n15372;
  assign n15374 = ~n15369 & ~n15373;
  assign n15375 = ~pi181 & ~n15374;
  assign n15376 = ~n15368 & n15375;
  assign n15377 = ~n14468 & n15265;
  assign n15378 = pi189 & n15035;
  assign n15379 = ~pi178 & ~n15378;
  assign n15380 = ~n15377 & n15379;
  assign n15381 = ~n14425 & n15370;
  assign n15382 = pi181 & ~n15381;
  assign n15383 = ~n15380 & n15382;
  assign n15384 = n11751 & ~n15383;
  assign n15385 = ~n15376 & n15384;
  assign n15386 = ~pi189 & n15041;
  assign n15387 = pi189 & n15046;
  assign n15388 = ~pi178 & ~n15387;
  assign n15389 = ~n15386 & n15388;
  assign n15390 = pi189 & n15102;
  assign n15391 = n15372 & ~n15390;
  assign n15392 = ~pi181 & ~n15391;
  assign n15393 = ~n15389 & n15392;
  assign n15394 = ~pi189 & ~n14468;
  assign n15395 = pi189 & ~n14482;
  assign n15396 = ~pi178 & ~n15395;
  assign n15397 = ~n15394 & n15396;
  assign n15398 = pi178 & n11760;
  assign n15399 = n14396 & n15398;
  assign n15400 = pi181 & ~n15399;
  assign n15401 = ~n14424 & n15400;
  assign n15402 = ~n15397 & n15401;
  assign n15403 = n11790 & ~n15402;
  assign n15404 = ~n15393 & n15403;
  assign n15405 = ~pi166 & ~n15027;
  assign n15406 = pi166 & ~n15035;
  assign n15407 = ~n15353 & ~n15406;
  assign n15408 = ~pi153 & ~n15407;
  assign n15409 = ~n15084 & n15358;
  assign n15410 = ~pi157 & ~n15409;
  assign n15411 = ~n15408 & n15410;
  assign n15412 = ~n15405 & n15411;
  assign n15413 = ~pi153 & ~n15314;
  assign n15414 = ~n14425 & n15413;
  assign n15415 = pi166 & n14479;
  assign n15416 = ~n14424 & ~n15415;
  assign n15417 = pi153 & ~n15416;
  assign n15418 = pi157 & ~n15417;
  assign n15419 = ~n15414 & n15418;
  assign n15420 = n9790 & ~n15419;
  assign n15421 = ~n15412 & n15420;
  assign n15422 = ~n15404 & ~n15421;
  assign n15423 = ~n15385 & n15422;
  assign n15424 = ~n15364 & n15423;
  assign n15425 = pi232 & ~n15424;
  assign n15426 = n15191 & ~n15425;
  assign n15427 = ~n10266 & ~n14534;
  assign n15428 = ~pi166 & n14540;
  assign n15429 = ~n15427 & ~n15428;
  assign n15430 = ~pi153 & ~n15429;
  assign n15431 = ~pi166 & n14543;
  assign n15432 = pi166 & n14587;
  assign n15433 = pi153 & ~n15432;
  assign n15434 = ~n15431 & n15433;
  assign n15435 = ~n15430 & ~n15434;
  assign n15436 = ~pi160 & ~n15435;
  assign n15437 = ~pi166 & n14552;
  assign n15438 = pi166 & ~n14555;
  assign n15439 = ~n15437 & ~n15438;
  assign n15440 = pi160 & ~n15242;
  assign n15441 = ~n15439 & n15440;
  assign n15442 = n9028 & ~n15441;
  assign n15443 = ~n15436 & n15442;
  assign n15444 = ~n9028 & ~n15313;
  assign n15445 = pi299 & ~n15444;
  assign n15446 = ~n15443 & n15445;
  assign n15447 = pi182 & n14555;
  assign n15448 = pi189 & ~n15150;
  assign n15449 = ~n15447 & n15448;
  assign n15450 = pi182 & n14551;
  assign n15451 = ~pi189 & ~n15450;
  assign n15452 = n15169 & n15451;
  assign n15453 = ~n15449 & ~n15452;
  assign n15454 = n11751 & ~n15453;
  assign n15455 = ~pi189 & ~n15147;
  assign n15456 = pi189 & ~n15151;
  assign n15457 = ~pi182 & ~n15456;
  assign n15458 = ~n15455 & n15457;
  assign n15459 = ~pi189 & ~n15157;
  assign n15460 = pi189 & ~n15161;
  assign n15461 = pi182 & ~n15460;
  assign n15462 = ~n15459 & n15461;
  assign n15463 = ~n15458 & ~n15462;
  assign n15464 = n11790 & ~n15463;
  assign n15465 = ~n15454 & ~n15464;
  assign n15466 = ~n15446 & n15465;
  assign n15467 = pi232 & ~n15466;
  assign n15468 = n15188 & ~n15467;
  assign n15469 = ~n15290 & ~n15468;
  assign n15470 = ~n15426 & n15469;
  assign n15471 = n3206 & ~n15470;
  assign n15472 = ~n15342 & n15471;
  assign n15473 = ~pi189 & n14479;
  assign n15474 = pi175 & n14334;
  assign n15475 = ~pi299 & ~n15474;
  assign n15476 = ~n15473 & n15475;
  assign n15477 = pi232 & ~n15476;
  assign n15478 = ~n15315 & n15477;
  assign n15479 = ~n3206 & n15478;
  assign n15480 = ~n3206 & n14331;
  assign n15481 = ~n15290 & n15480;
  assign n15482 = n3278 & ~n15481;
  assign n15483 = ~n15479 & n15482;
  assign n15484 = ~n15472 & n15483;
  assign n15485 = n14621 & ~n15478;
  assign n15486 = ~pi150 & pi299;
  assign n15487 = ~pi185 & ~pi299;
  assign n15488 = ~n15486 & ~n15487;
  assign n15489 = n7462 & n15488;
  assign n15490 = pi87 & ~n15489;
  assign n15491 = ~n15485 & ~n15490;
  assign n15492 = n14354 & ~n15290;
  assign n15493 = ~n15491 & ~n15492;
  assign n15494 = ~po1038 & ~n15493;
  assign n15495 = ~n15484 & n15494;
  assign n15496 = pi232 & ~n15310;
  assign n15497 = n15290 & ~n15496;
  assign n15498 = ~pi232 & ~n14331;
  assign n15499 = ~n15313 & ~n15498;
  assign n15500 = ~n15497 & n15499;
  assign n15501 = ~pi87 & ~n15500;
  assign n15502 = pi87 & ~n13738;
  assign n15503 = po1038 & ~n15502;
  assign n15504 = ~n15501 & n15503;
  assign po283 = ~n15495 & ~n15504;
  assign n15506 = n3280 & n8846;
  assign n15507 = ~n3293 & ~n15506;
  assign n15508 = pi129 & n6109;
  assign n15509 = pi38 & ~n15508;
  assign n15510 = ~n2524 & ~n2850;
  assign n15511 = n2597 & ~n2669;
  assign n15512 = n2451 & ~n15511;
  assign n15513 = n2683 & ~n15512;
  assign n15514 = n2594 & ~n15513;
  assign n15515 = n2687 & ~n15514;
  assign n15516 = n2504 & ~n15515;
  assign n15517 = ~n2507 & ~n15516;
  assign n15518 = ~pi86 & ~n15517;
  assign n15519 = n2592 & ~n15518;
  assign n15520 = n2590 & ~n15519;
  assign n15521 = ~n2585 & ~n15520;
  assign n15522 = ~pi108 & ~n15521;
  assign n15523 = n2584 & ~n15522;
  assign n15524 = n2699 & ~n15523;
  assign n15525 = ~n2575 & ~n15524;
  assign n15526 = n2574 & ~n15525;
  assign n15527 = n2573 & ~n15526;
  assign n15528 = ~po740 & n15527;
  assign n15529 = ~pi97 & ~n15519;
  assign n15530 = ~n2585 & ~n15529;
  assign n15531 = ~pi108 & ~n15530;
  assign n15532 = n2584 & ~n15531;
  assign n15533 = n2699 & ~n15532;
  assign n15534 = ~n2575 & ~n15533;
  assign n15535 = n2574 & ~n15534;
  assign n15536 = n2573 & ~n15535;
  assign n15537 = po740 & n15536;
  assign n15538 = pi250 & ~n7463;
  assign n15539 = n10022 & n15538;
  assign n15540 = ~n15537 & n15539;
  assign n15541 = ~n15528 & n15540;
  assign n15542 = pi127 & n15527;
  assign n15543 = ~pi127 & n15536;
  assign n15544 = ~n15539 & ~n15543;
  assign n15545 = ~n15542 & n15544;
  assign n15546 = ~n15541 & ~n15545;
  assign n15547 = n2566 & ~n15546;
  assign n15548 = n2852 & ~n15547;
  assign n15549 = n2547 & ~n15548;
  assign n15550 = n15510 & ~n15549;
  assign n15551 = ~pi70 & ~n15550;
  assign n15552 = ~n2843 & ~n15551;
  assign n15553 = ~pi51 & ~n15552;
  assign n15554 = n2559 & ~n15553;
  assign n15555 = n2921 & ~n15554;
  assign n15556 = ~n2555 & ~n15555;
  assign n15557 = n2725 & ~n15556;
  assign n15558 = n3361 & ~n15557;
  assign n15559 = ~pi95 & ~n15558;
  assign n15560 = ~pi39 & pi129;
  assign n15561 = ~n2727 & n15560;
  assign n15562 = ~n15559 & n15561;
  assign n15563 = pi39 & n8846;
  assign n15564 = ~pi38 & ~n15563;
  assign n15565 = ~n15562 & n15564;
  assign n15566 = ~n15509 & ~n15565;
  assign n15567 = n3240 & ~n15566;
  assign n15568 = ~n3207 & ~n8924;
  assign n15569 = n8846 & ~n15568;
  assign n15570 = ~n3240 & ~n15569;
  assign n15571 = ~pi75 & ~n15570;
  assign n15572 = ~n15567 & n15571;
  assign n15573 = pi129 & n7268;
  assign n15574 = pi75 & n15573;
  assign n15575 = ~pi92 & ~n15574;
  assign n15576 = ~n15572 & n15575;
  assign n15577 = pi92 & ~pi129;
  assign n15578 = n13563 & ~n15577;
  assign n15579 = ~n15576 & n15578;
  assign n15580 = pi54 & n3238;
  assign n15581 = n8846 & n15580;
  assign n15582 = ~pi74 & ~n15581;
  assign n15583 = ~n15579 & n15582;
  assign n15584 = n6536 & n15573;
  assign n15585 = pi74 & ~n15584;
  assign n15586 = ~pi55 & ~n15585;
  assign n15587 = ~n15583 & n15586;
  assign n15588 = pi55 & n3266;
  assign n15589 = n15573 & n15588;
  assign n15590 = ~n15587 & ~n15589;
  assign n15591 = ~pi56 & ~n15590;
  assign n15592 = ~n11247 & ~n11256;
  assign n15593 = ~n15591 & n15592;
  assign n15594 = ~n15507 & ~n15593;
  assign n15595 = n3429 & ~n15594;
  assign n15596 = ~pi129 & ~n3429;
  assign n15597 = n6100 & ~n15596;
  assign po284 = ~n15595 & n15597;
  assign n15599 = ~n6107 & ~n7314;
  assign n15600 = ~pi38 & ~n3366;
  assign n15601 = n6111 & ~n15600;
  assign n15602 = n6236 & ~n6261;
  assign n15603 = ~pi87 & ~n15602;
  assign n15604 = ~n15601 & n15603;
  assign n15605 = n6270 & ~n15604;
  assign n15606 = n8848 & n10353;
  assign n15607 = ~pi129 & ~n15606;
  assign n15608 = po740 & n15606;
  assign n15609 = n8926 & ~n15608;
  assign n15610 = ~n15607 & n15609;
  assign n15611 = n3095 & n15610;
  assign n15612 = n6271 & ~n15611;
  assign n15613 = ~n15605 & n15612;
  assign n15614 = ~n7272 & ~n7308;
  assign n15615 = ~n15613 & n15614;
  assign n15616 = n8839 & ~n15615;
  assign n15617 = n15599 & ~n15616;
  assign n15618 = ~pi56 & ~n15617;
  assign n15619 = ~n6104 & ~n15618;
  assign n15620 = ~pi62 & ~n15619;
  assign n15621 = ~n6280 & ~n15620;
  assign n15622 = n3429 & ~n15621;
  assign po286 = n6100 & ~n15622;
  assign n15624 = ~pi51 & ~n15186;
  assign n15625 = ~pi232 & ~n15624;
  assign n15626 = n10922 & ~n15625;
  assign n15627 = ~pi51 & ~n14541;
  assign n15628 = ~n14550 & n15627;
  assign n15629 = pi169 & ~n15628;
  assign n15630 = pi162 & n9028;
  assign n15631 = ~pi169 & ~n15159;
  assign n15632 = n15630 & ~n15631;
  assign n15633 = ~n15629 & n15632;
  assign n15634 = pi169 & n6162;
  assign n15635 = ~n3095 & n15634;
  assign n15636 = ~n14579 & ~n15634;
  assign n15637 = ~pi162 & n9028;
  assign n15638 = ~n15636 & n15637;
  assign n15639 = ~n15635 & n15638;
  assign n15640 = ~n9028 & n14396;
  assign n15641 = ~n15634 & n15640;
  assign n15642 = pi299 & ~n15641;
  assign n15643 = ~n15639 & n15642;
  assign n15644 = ~n15633 & n15643;
  assign n15645 = ~pi191 & ~pi299;
  assign n15646 = ~pi51 & ~n15150;
  assign n15647 = pi140 & n15160;
  assign n15648 = n15646 & ~n15647;
  assign n15649 = n15645 & ~n15648;
  assign n15650 = ~pi51 & n15169;
  assign n15651 = pi140 & n14550;
  assign n15652 = n15650 & ~n15651;
  assign n15653 = n8969 & ~n15652;
  assign n15654 = ~n15649 & ~n15653;
  assign n15655 = ~n15644 & n15654;
  assign n15656 = pi232 & ~n15655;
  assign n15657 = n15626 & ~n15656;
  assign n15658 = n7462 & ~n8971;
  assign n15659 = n14396 & ~n15658;
  assign n15660 = ~n10922 & n15659;
  assign n15661 = ~pi100 & ~n15660;
  assign n15662 = ~n15657 & n15661;
  assign n15663 = ~n15310 & ~n15659;
  assign n15664 = pi100 & n15663;
  assign n15665 = n3278 & ~n15664;
  assign n15666 = ~n14616 & n15665;
  assign n15667 = ~n15662 & n15666;
  assign n15668 = pi87 & ~n9694;
  assign n15669 = n14621 & ~n15663;
  assign n15670 = ~n15668 & ~n15669;
  assign n15671 = ~n14354 & ~n15670;
  assign n15672 = ~pi132 & n15287;
  assign n15673 = pi130 & ~n15672;
  assign n15674 = ~pi130 & n15672;
  assign n15675 = ~n15673 & ~n15674;
  assign n15676 = ~n14345 & ~n15675;
  assign n15677 = ~n15671 & ~n15676;
  assign n15678 = ~n15667 & n15677;
  assign n15679 = ~n14586 & n14984;
  assign n15680 = pi224 & ~n15679;
  assign n15681 = ~n6162 & ~n14539;
  assign n15682 = ~n14933 & ~n15681;
  assign n15683 = ~pi224 & ~n15682;
  assign n15684 = ~n15680 & ~n15683;
  assign n15685 = n6461 & ~n15684;
  assign n15686 = ~n6461 & ~n15310;
  assign n15687 = ~n15685 & ~n15686;
  assign n15688 = pi140 & n15687;
  assign n15689 = n8050 & ~n15682;
  assign n15690 = ~n8050 & ~n15310;
  assign n15691 = ~n15689 & ~n15690;
  assign n15692 = ~pi140 & n15691;
  assign n15693 = n8969 & ~n15692;
  assign n15694 = ~n15688 & n15693;
  assign n15695 = ~n14539 & ~n15634;
  assign n15696 = pi169 & n14933;
  assign n15697 = ~n15695 & ~n15696;
  assign n15698 = ~pi216 & ~n15697;
  assign n15699 = ~pi51 & ~n14923;
  assign n15700 = ~pi169 & n15699;
  assign n15701 = pi169 & n15679;
  assign n15702 = pi162 & pi216;
  assign n15703 = ~n15701 & n15702;
  assign n15704 = ~n15700 & n15703;
  assign n15705 = ~n15698 & ~n15704;
  assign n15706 = n6434 & ~n15705;
  assign n15707 = pi169 & n14479;
  assign n15708 = ~pi51 & ~n15707;
  assign n15709 = ~n8039 & ~n15630;
  assign n15710 = ~n15708 & n15709;
  assign n15711 = ~n15706 & ~n15710;
  assign n15712 = pi299 & ~n15711;
  assign n15713 = n14538 & n14926;
  assign n15714 = ~pi51 & ~n15713;
  assign n15715 = pi140 & n15714;
  assign n15716 = n8050 & n14538;
  assign n15717 = ~pi51 & ~n15716;
  assign n15718 = ~pi140 & n15717;
  assign n15719 = n15645 & ~n15718;
  assign n15720 = ~n15715 & n15719;
  assign n15721 = ~n15712 & ~n15720;
  assign n15722 = ~n15694 & n15721;
  assign n15723 = pi232 & ~n15722;
  assign n15724 = n14538 & ~n14919;
  assign n15725 = ~pi51 & ~n15724;
  assign n15726 = ~pi232 & ~n15725;
  assign n15727 = pi39 & ~n15726;
  assign n15728 = ~n15723 & n15727;
  assign n15729 = ~pi232 & ~n14453;
  assign n15730 = ~pi39 & ~n15729;
  assign n15731 = ~n6162 & n14453;
  assign n15732 = ~n14847 & ~n15731;
  assign n15733 = ~n8971 & ~n15732;
  assign n15734 = n8971 & n14453;
  assign n15735 = pi232 & ~n15734;
  assign n15736 = ~n15733 & n15735;
  assign n15737 = n15730 & ~n15736;
  assign n15738 = ~n15728 & ~n15737;
  assign n15739 = ~pi38 & ~n15738;
  assign n15740 = pi38 & ~n15663;
  assign n15741 = ~pi100 & ~n15740;
  assign n15742 = ~n15739 & n15741;
  assign n15743 = n15665 & ~n15742;
  assign n15744 = n15670 & n15676;
  assign n15745 = ~n15743 & n15744;
  assign n15746 = ~n15678 & ~n15745;
  assign n15747 = ~po1038 & ~n15746;
  assign n15748 = ~pi51 & ~pi87;
  assign n15749 = ~n15707 & n15748;
  assign n15750 = n15676 & n15749;
  assign n15751 = pi169 & n7462;
  assign n15752 = ~pi87 & n14396;
  assign n15753 = ~n15751 & n15752;
  assign n15754 = pi87 & ~n9649;
  assign n15755 = po1038 & ~n15754;
  assign n15756 = ~n15753 & n15755;
  assign n15757 = ~n15750 & n15756;
  assign po287 = ~n15747 & ~n15757;
  assign n15759 = ~pi100 & ~n13910;
  assign n15760 = ~pi87 & ~n7301;
  assign n15761 = ~n15759 & n15760;
  assign n15762 = ~pi75 & ~n15761;
  assign n15763 = ~n7269 & ~n15762;
  assign n15764 = ~pi92 & ~n15763;
  assign n15765 = n8840 & n13563;
  assign po288 = ~n15764 & n15765;
  assign n15767 = pi51 & ~pi151;
  assign n15768 = ~n13643 & ~n14334;
  assign n15769 = ~n15767 & ~n15768;
  assign n15770 = n14332 & n15769;
  assign n15771 = pi232 & n15770;
  assign n15772 = pi132 & ~n15287;
  assign n15773 = ~n15672 & ~n15772;
  assign n15774 = ~n14346 & ~n15773;
  assign n15775 = n14331 & ~n15774;
  assign n15776 = ~n15771 & ~n15775;
  assign n15777 = ~pi87 & ~n15776;
  assign n15778 = pi164 & n14810;
  assign n15779 = po1038 & ~n15778;
  assign n15780 = ~n15777 & n15779;
  assign n15781 = ~pi190 & ~pi299;
  assign n15782 = ~n6162 & ~n14464;
  assign n15783 = pi182 & ~n15782;
  assign n15784 = ~n14447 & n15783;
  assign n15785 = ~pi182 & n14464;
  assign n15786 = ~pi173 & ~n15785;
  assign n15787 = ~n15784 & n15786;
  assign n15788 = ~n6162 & n14464;
  assign n15789 = ~n14454 & ~n15788;
  assign n15790 = pi182 & ~n15789;
  assign n15791 = n14469 & ~n15788;
  assign n15792 = ~pi182 & ~n15791;
  assign n15793 = pi173 & ~n15792;
  assign n15794 = ~n15790 & n15793;
  assign n15795 = ~n15787 & ~n15794;
  assign n15796 = n15781 & ~n15795;
  assign n15797 = ~pi151 & ~n14446;
  assign n15798 = pi151 & n14453;
  assign n15799 = ~pi168 & ~n15798;
  assign n15800 = ~n15797 & n15799;
  assign n15801 = pi168 & ~n15767;
  assign n15802 = ~n14402 & n15801;
  assign n15803 = n6162 & ~n15802;
  assign n15804 = ~n15800 & n15803;
  assign n15805 = pi160 & ~n15782;
  assign n15806 = ~n15804 & n15805;
  assign n15807 = ~pi168 & ~n15791;
  assign n15808 = pi168 & ~n14861;
  assign n15809 = ~n15782 & n15808;
  assign n15810 = pi151 & ~n15809;
  assign n15811 = ~n15807 & n15810;
  assign n15812 = ~n13643 & n14464;
  assign n15813 = pi168 & n14475;
  assign n15814 = ~pi151 & ~n15813;
  assign n15815 = ~n15812 & n15814;
  assign n15816 = ~pi160 & ~n15815;
  assign n15817 = ~n15811 & n15816;
  assign n15818 = pi299 & ~n15817;
  assign n15819 = ~n15806 & n15818;
  assign n15820 = pi190 & ~pi299;
  assign n15821 = pi182 & n14382;
  assign n15822 = n14401 & ~n15821;
  assign n15823 = pi51 & ~pi173;
  assign n15824 = n6162 & ~n15823;
  assign n15825 = ~n15822 & n15824;
  assign n15826 = n15820 & ~n15825;
  assign n15827 = ~n15788 & n15826;
  assign n15828 = pi232 & ~n15827;
  assign n15829 = ~n15819 & n15828;
  assign n15830 = ~n15796 & n15829;
  assign n15831 = ~pi232 & n14464;
  assign n15832 = ~n15830 & ~n15831;
  assign n15833 = ~pi39 & ~n15832;
  assign n15834 = pi168 & ~n14934;
  assign n15835 = ~pi168 & ~n14928;
  assign n15836 = ~n15834 & ~n15835;
  assign n15837 = ~n15767 & ~n15836;
  assign n15838 = ~pi216 & ~n15837;
  assign n15839 = ~pi168 & ~n14924;
  assign n15840 = pi168 & ~n14984;
  assign n15841 = pi151 & ~n15840;
  assign n15842 = ~n15839 & n15841;
  assign n15843 = ~pi168 & n14700;
  assign n15844 = pi168 & n14582;
  assign n15845 = ~pi151 & ~n15844;
  assign n15846 = ~n15843 & n15845;
  assign n15847 = pi149 & ~n15846;
  assign n15848 = ~n15842 & n15847;
  assign n15849 = pi216 & ~n15848;
  assign n15850 = n6434 & ~n15849;
  assign n15851 = ~n15838 & n15850;
  assign n15852 = pi299 & ~n15770;
  assign n15853 = ~pi149 & pi216;
  assign n15854 = n6587 & ~n15853;
  assign n15855 = ~n15852 & ~n15854;
  assign n15856 = ~n15851 & ~n15855;
  assign n15857 = pi183 & ~n14950;
  assign n15858 = ~pi183 & ~n14945;
  assign n15859 = ~pi173 & ~n15858;
  assign n15860 = ~n15857 & n15859;
  assign n15861 = ~pi183 & n14959;
  assign n15862 = ~pi183 & ~n14935;
  assign n15863 = pi173 & ~n14940;
  assign n15864 = ~n15862 & n15863;
  assign n15865 = ~n15861 & ~n15864;
  assign n15866 = ~n15860 & n15865;
  assign n15867 = n15820 & ~n15866;
  assign n15868 = pi183 & n14931;
  assign n15869 = ~pi183 & ~n14334;
  assign n15870 = ~n14962 & n15869;
  assign n15871 = pi173 & ~n15870;
  assign n15872 = ~n15868 & n15871;
  assign n15873 = ~pi183 & ~n8050;
  assign n15874 = ~pi173 & ~n15873;
  assign n15875 = n14953 & n15874;
  assign n15876 = n15781 & ~n15875;
  assign n15877 = ~n15872 & n15876;
  assign n15878 = ~n15867 & ~n15877;
  assign n15879 = ~n15856 & n15878;
  assign n15880 = pi232 & ~n15879;
  assign n15881 = n14922 & ~n15880;
  assign n15882 = ~n15833 & ~n15881;
  assign n15883 = n3206 & ~n15882;
  assign n15884 = pi190 & n14479;
  assign n15885 = pi173 & n14334;
  assign n15886 = ~pi299 & ~n15885;
  assign n15887 = ~n15884 & n15886;
  assign n15888 = pi232 & ~n15887;
  assign n15889 = ~n15852 & n15888;
  assign n15890 = ~n3206 & n15889;
  assign n15891 = n3278 & ~n15890;
  assign n15892 = ~n15883 & n15891;
  assign n15893 = n14621 & ~n15889;
  assign n15894 = pi87 & ~n8979;
  assign n15895 = n15774 & ~n15894;
  assign n15896 = ~n15893 & n15895;
  assign n15897 = ~n15892 & n15896;
  assign n15898 = ~pi183 & ~n15147;
  assign n15899 = pi183 & ~n15157;
  assign n15900 = pi173 & ~n15899;
  assign n15901 = ~n15898 & n15900;
  assign n15902 = pi183 & n14551;
  assign n15903 = ~pi173 & ~n15902;
  assign n15904 = n15169 & n15903;
  assign n15905 = ~n15901 & ~n15904;
  assign n15906 = n15820 & ~n15905;
  assign n15907 = ~n14331 & n15852;
  assign n15908 = ~n13047 & ~n15907;
  assign n15909 = ~n14555 & ~n15769;
  assign n15910 = ~pi168 & ~n15909;
  assign n15911 = pi149 & ~n15910;
  assign n15912 = ~pi151 & n14334;
  assign n15913 = pi168 & ~n15912;
  assign n15914 = ~n14537 & n15913;
  assign n15915 = ~n15628 & n15914;
  assign n15916 = n15911 & ~n15915;
  assign n15917 = pi168 & ~n14543;
  assign n15918 = ~pi168 & ~n14587;
  assign n15919 = pi151 & ~n15918;
  assign n15920 = ~n15917 & n15919;
  assign n15921 = pi168 & n14540;
  assign n15922 = ~n13643 & ~n14534;
  assign n15923 = ~pi151 & ~n15922;
  assign n15924 = ~n15921 & n15923;
  assign n15925 = ~pi149 & ~n15924;
  assign n15926 = ~n15920 & n15925;
  assign n15927 = n9028 & ~n15926;
  assign n15928 = ~n15916 & n15927;
  assign n15929 = ~n15908 & ~n15928;
  assign n15930 = pi183 & n14555;
  assign n15931 = n15781 & ~n15885;
  assign n15932 = ~n15150 & n15931;
  assign n15933 = ~n15930 & n15932;
  assign n15934 = ~n15929 & ~n15933;
  assign n15935 = ~n15906 & n15934;
  assign n15936 = pi232 & ~n15935;
  assign n15937 = ~n15187 & ~n15936;
  assign n15938 = pi39 & ~n15937;
  assign n15939 = pi151 & n14657;
  assign n15940 = ~pi151 & ~n14422;
  assign n15941 = ~pi168 & ~n15940;
  assign n15942 = ~n15939 & n15941;
  assign n15943 = ~n14411 & n15913;
  assign n15944 = ~n15942 & ~n15943;
  assign n15945 = ~pi160 & ~n15033;
  assign n15946 = ~n15944 & n15945;
  assign n15947 = ~pi151 & ~n15770;
  assign n15948 = ~n15034 & n15947;
  assign n15949 = ~pi168 & n14479;
  assign n15950 = ~n15033 & ~n15949;
  assign n15951 = pi151 & ~n15950;
  assign n15952 = pi160 & ~n15951;
  assign n15953 = ~n15948 & n15952;
  assign n15954 = pi299 & ~n15953;
  assign n15955 = ~n15946 & n15954;
  assign n15956 = ~pi182 & n14411;
  assign n15957 = ~n15033 & ~n15823;
  assign n15958 = ~n15956 & n15957;
  assign n15959 = n15820 & ~n15958;
  assign n15960 = pi182 & n15034;
  assign n15961 = ~n14422 & n15931;
  assign n15962 = ~n15960 & n15961;
  assign n15963 = pi232 & ~n15962;
  assign n15964 = ~n15959 & n15963;
  assign n15965 = ~n15955 & n15964;
  assign n15966 = ~pi232 & n14422;
  assign n15967 = ~pi39 & ~n15966;
  assign n15968 = ~n15965 & n15967;
  assign n15969 = n3206 & ~n15968;
  assign n15970 = ~n15938 & n15969;
  assign n15971 = n3278 & ~n15480;
  assign n15972 = ~n15890 & n15971;
  assign n15973 = ~n15970 & n15972;
  assign n15974 = n14622 & ~n15889;
  assign n15975 = ~n15774 & ~n15894;
  assign n15976 = ~n15974 & n15975;
  assign n15977 = ~n15973 & n15976;
  assign n15978 = ~po1038 & ~n15977;
  assign n15979 = ~n15897 & n15978;
  assign po289 = n15780 | n15979;
  assign n15981 = ~n6162 & ~n14416;
  assign n15982 = ~n14447 & ~n15981;
  assign n15983 = pi299 & n9411;
  assign n15984 = n15982 & n15983;
  assign n15985 = n14416 & ~n15983;
  assign n15986 = ~pi39 & ~pi176;
  assign n15987 = ~n15985 & n15986;
  assign n15988 = ~n15984 & n15987;
  assign n15989 = n9411 & n15982;
  assign n15990 = ~n9411 & n14416;
  assign n15991 = ~pi39 & pi176;
  assign n15992 = ~n15990 & n15991;
  assign n15993 = ~n15989 & n15992;
  assign n15994 = pi197 & n14550;
  assign n15995 = ~n5745 & ~n15994;
  assign n15996 = n6587 & ~n15995;
  assign n15997 = ~pi145 & ~n8050;
  assign n15998 = ~pi299 & ~n15997;
  assign n15999 = ~n14952 & n15998;
  assign n16000 = ~n15996 & ~n15999;
  assign n16001 = n3095 & ~n16000;
  assign n16002 = pi232 & ~n16001;
  assign n16003 = ~n14921 & ~n16002;
  assign n16004 = pi39 & ~n16003;
  assign n16005 = n11320 & ~n16004;
  assign n16006 = ~n15993 & n16005;
  assign n16007 = ~n15988 & n16006;
  assign n16008 = ~pi133 & ~n14799;
  assign n16009 = ~pi87 & n16008;
  assign n16010 = ~n16007 & n16009;
  assign n16011 = pi145 & n14555;
  assign n16012 = n15182 & ~n16011;
  assign n16013 = n15183 & ~n15994;
  assign n16014 = n14331 & ~n16013;
  assign n16015 = pi299 & ~n16014;
  assign n16016 = ~n16012 & ~n16015;
  assign n16017 = pi232 & ~n16016;
  assign n16018 = n15188 & ~n16017;
  assign n16019 = ~n9414 & n14399;
  assign n16020 = ~pi39 & n14331;
  assign n16021 = ~n16019 & n16020;
  assign n16022 = ~pi38 & ~n16021;
  assign n16023 = ~n16018 & n16022;
  assign n16024 = n14370 & ~n16023;
  assign n16025 = n14617 & ~n16024;
  assign n16026 = ~n14622 & ~n16025;
  assign n16027 = ~n16008 & ~n16026;
  assign n16028 = ~pi183 & ~pi299;
  assign n16029 = ~pi149 & pi299;
  assign n16030 = ~n16028 & ~n16029;
  assign n16031 = n7462 & n16030;
  assign n16032 = pi87 & ~n16031;
  assign n16033 = ~n16027 & ~n16032;
  assign n16034 = ~n16010 & n16033;
  assign n16035 = ~po1038 & ~n16034;
  assign n16036 = n14354 & ~n16008;
  assign n16037 = pi149 & n14810;
  assign n16038 = po1038 & ~n16037;
  assign n16039 = ~n16036 & n16038;
  assign po290 = n16035 | n16039;
  assign n16041 = ~pi136 & n15674;
  assign n16042 = ~pi135 & n16041;
  assign n16043 = pi134 & ~n16042;
  assign n16044 = n14330 & ~n16043;
  assign n16045 = po1038 & n15748;
  assign n16046 = pi171 & n6162;
  assign n16047 = ~n14330 & n16046;
  assign n16048 = pi232 & n16047;
  assign n16049 = n16045 & ~n16048;
  assign n16050 = ~n16044 & n16049;
  assign n16051 = pi39 & pi186;
  assign n16052 = pi192 & ~pi299;
  assign n16053 = ~n14550 & n15650;
  assign n16054 = n16052 & ~n16053;
  assign n16055 = ~pi192 & ~pi299;
  assign n16056 = ~n15160 & n15646;
  assign n16057 = n16055 & ~n16056;
  assign n16058 = ~n16054 & ~n16057;
  assign n16059 = n15640 & ~n16046;
  assign n16060 = pi299 & ~n16059;
  assign n16061 = pi171 & ~n15628;
  assign n16062 = ~pi171 & ~n15159;
  assign n16063 = n9028 & ~n16062;
  assign n16064 = ~n16061 & n16063;
  assign n16065 = n16060 & ~n16064;
  assign n16066 = n16058 & ~n16065;
  assign n16067 = pi232 & ~n16066;
  assign n16068 = ~n15625 & ~n16067;
  assign n16069 = n16051 & ~n16068;
  assign n16070 = pi39 & ~pi186;
  assign n16071 = ~n15650 & n16052;
  assign n16072 = ~n15646 & n16055;
  assign n16073 = ~n16071 & ~n16072;
  assign n16074 = ~n16065 & n16073;
  assign n16075 = pi232 & ~n16074;
  assign n16076 = ~n15625 & ~n16075;
  assign n16077 = n16070 & ~n16076;
  assign n16078 = pi171 & pi299;
  assign n16079 = ~n16052 & ~n16078;
  assign n16080 = n7462 & ~n16079;
  assign n16081 = n14396 & ~n16080;
  assign n16082 = ~pi39 & ~n16081;
  assign n16083 = pi164 & ~n16082;
  assign n16084 = ~n16077 & n16083;
  assign n16085 = ~n16069 & n16084;
  assign n16086 = n4212 & n6162;
  assign n16087 = ~n14579 & ~n16046;
  assign n16088 = n9028 & ~n16087;
  assign n16089 = ~n16086 & n16088;
  assign n16090 = n16060 & ~n16089;
  assign n16091 = n16058 & ~n16090;
  assign n16092 = pi232 & ~n16091;
  assign n16093 = ~n15625 & ~n16092;
  assign n16094 = n16051 & ~n16093;
  assign n16095 = n16073 & ~n16090;
  assign n16096 = pi232 & ~n16095;
  assign n16097 = ~n15625 & ~n16096;
  assign n16098 = n16070 & ~n16097;
  assign n16099 = ~pi164 & ~n16082;
  assign n16100 = ~n16098 & n16099;
  assign n16101 = ~n16094 & n16100;
  assign n16102 = n3206 & ~n16101;
  assign n16103 = ~n16085 & n16102;
  assign n16104 = ~n15310 & ~n16081;
  assign n16105 = ~n3206 & n16104;
  assign n16106 = n3278 & ~n16105;
  assign n16107 = ~n15480 & n16106;
  assign n16108 = ~n16103 & n16107;
  assign n16109 = n14621 & n16081;
  assign n16110 = ~n16043 & ~n16109;
  assign n16111 = ~n16108 & n16110;
  assign n16112 = pi232 & ~n16079;
  assign n16113 = n15732 & n16112;
  assign n16114 = ~n14453 & ~n16112;
  assign n16115 = ~pi39 & ~n16114;
  assign n16116 = ~n16113 & n16115;
  assign n16117 = ~pi51 & ~n16047;
  assign n16118 = ~pi164 & pi216;
  assign n16119 = n6434 & ~n16118;
  assign n16120 = ~n16117 & ~n16119;
  assign n16121 = ~n14539 & ~n16046;
  assign n16122 = pi171 & n14933;
  assign n16123 = ~n16121 & ~n16122;
  assign n16124 = ~pi216 & ~n16123;
  assign n16125 = ~pi171 & n15699;
  assign n16126 = pi171 & n15679;
  assign n16127 = pi164 & pi216;
  assign n16128 = ~n16126 & n16127;
  assign n16129 = ~n16125 & n16128;
  assign n16130 = ~n16124 & ~n16129;
  assign n16131 = n6434 & ~n16130;
  assign n16132 = ~n16120 & ~n16131;
  assign n16133 = pi299 & ~n16132;
  assign n16134 = ~n15691 & n16052;
  assign n16135 = ~n15717 & n16055;
  assign n16136 = ~n16051 & ~n16135;
  assign n16137 = ~n16134 & n16136;
  assign n16138 = ~n15687 & n16052;
  assign n16139 = ~n15714 & n16055;
  assign n16140 = pi186 & ~n16139;
  assign n16141 = ~n16138 & n16140;
  assign n16142 = ~n16137 & ~n16141;
  assign n16143 = ~n16133 & ~n16142;
  assign n16144 = pi232 & ~n16143;
  assign n16145 = n15727 & ~n16144;
  assign n16146 = n3206 & ~n16145;
  assign n16147 = ~n16116 & n16146;
  assign n16148 = n16106 & ~n16147;
  assign n16149 = n14621 & ~n16104;
  assign n16150 = n16043 & ~n16149;
  assign n16151 = ~n16148 & n16150;
  assign n16152 = ~po1038 & ~n16151;
  assign n16153 = ~n16111 & n16152;
  assign po291 = n16050 | n16153;
  assign n16155 = pi170 & n6162;
  assign n16156 = n10607 & n16155;
  assign n16157 = n14396 & ~n16156;
  assign n16158 = pi194 & n8990;
  assign n16159 = n16157 & ~n16158;
  assign n16160 = ~n15310 & ~n16159;
  assign n16161 = pi100 & n16160;
  assign n16162 = n3278 & ~n16161;
  assign n16163 = ~n14539 & ~n16155;
  assign n16164 = pi170 & n14933;
  assign n16165 = n8039 & ~n16164;
  assign n16166 = ~n16163 & n16165;
  assign n16167 = ~n9028 & ~n16166;
  assign n16168 = ~pi170 & n15699;
  assign n16169 = pi170 & n15679;
  assign n16170 = pi216 & ~n16169;
  assign n16171 = ~n16168 & n16170;
  assign n16172 = ~n16167 & ~n16171;
  assign n16173 = pi150 & pi299;
  assign n16174 = ~n14330 & n16155;
  assign n16175 = ~pi51 & ~n16174;
  assign n16176 = ~n6434 & n16175;
  assign n16177 = n16173 & ~n16176;
  assign n16178 = ~n16172 & n16177;
  assign n16179 = ~n8039 & n16175;
  assign n16180 = n15486 & ~n16179;
  assign n16181 = ~n16166 & n16180;
  assign n16182 = ~n16178 & ~n16181;
  assign n16183 = pi185 & n15714;
  assign n16184 = ~pi185 & n15717;
  assign n16185 = ~pi299 & ~n16184;
  assign n16186 = ~n16183 & n16185;
  assign n16187 = n16182 & ~n16186;
  assign n16188 = pi232 & ~n16187;
  assign n16189 = n15727 & ~n16188;
  assign n16190 = ~pi299 & ~n14453;
  assign n16191 = pi170 & ~n15732;
  assign n16192 = ~pi170 & n14453;
  assign n16193 = n10607 & ~n16192;
  assign n16194 = ~n16191 & n16193;
  assign n16195 = n15730 & ~n16194;
  assign n16196 = ~n16190 & n16195;
  assign n16197 = ~n16189 & ~n16196;
  assign n16198 = ~pi38 & ~n16197;
  assign n16199 = ~n15310 & ~n16157;
  assign n16200 = pi38 & ~n16199;
  assign n16201 = ~pi194 & ~n16200;
  assign n16202 = ~n16198 & n16201;
  assign n16203 = pi185 & n15687;
  assign n16204 = ~pi185 & n15691;
  assign n16205 = ~pi299 & ~n16204;
  assign n16206 = ~n16203 & n16205;
  assign n16207 = n16182 & ~n16206;
  assign n16208 = pi232 & ~n16207;
  assign n16209 = n15727 & ~n16208;
  assign n16210 = n10602 & n15732;
  assign n16211 = n16195 & ~n16210;
  assign n16212 = ~n16209 & ~n16211;
  assign n16213 = ~pi38 & ~n16212;
  assign n16214 = pi170 & n7462;
  assign n16215 = ~n8990 & ~n16214;
  assign n16216 = n14396 & n16215;
  assign n16217 = ~n15310 & ~n16216;
  assign n16218 = pi38 & ~n16217;
  assign n16219 = pi194 & ~n16218;
  assign n16220 = ~n16213 & n16219;
  assign n16221 = ~n16202 & ~n16220;
  assign n16222 = ~pi100 & ~n16221;
  assign n16223 = n16162 & ~n16222;
  assign n16224 = pi135 & ~n16041;
  assign n16225 = pi134 & n16042;
  assign n16226 = ~n16224 & ~n16225;
  assign n16227 = n14621 & ~n16160;
  assign n16228 = ~n16226 & ~n16227;
  assign n16229 = ~n16223 & n16228;
  assign n16230 = pi185 & n15160;
  assign n16231 = n15646 & ~n16230;
  assign n16232 = ~n10922 & n16157;
  assign n16233 = ~pi194 & ~n16232;
  assign n16234 = ~n16231 & n16233;
  assign n16235 = ~pi185 & n15650;
  assign n16236 = ~n10922 & n16216;
  assign n16237 = pi194 & ~n16236;
  assign n16238 = ~n16053 & n16237;
  assign n16239 = ~n16235 & n16238;
  assign n16240 = ~n16234 & ~n16239;
  assign n16241 = ~pi299 & ~n16240;
  assign n16242 = pi170 & ~n15628;
  assign n16243 = ~pi170 & ~n15159;
  assign n16244 = n9028 & ~n16243;
  assign n16245 = ~n16242 & n16244;
  assign n16246 = n16173 & ~n16245;
  assign n16247 = n4435 & n6162;
  assign n16248 = ~n14579 & ~n16155;
  assign n16249 = n9028 & ~n16248;
  assign n16250 = ~n16247 & n16249;
  assign n16251 = n15486 & ~n16250;
  assign n16252 = ~n16246 & ~n16251;
  assign n16253 = n15640 & ~n16155;
  assign n16254 = ~n16233 & ~n16237;
  assign n16255 = ~n16253 & ~n16254;
  assign n16256 = ~n16252 & n16255;
  assign n16257 = ~n16241 & ~n16256;
  assign n16258 = pi232 & ~n16257;
  assign n16259 = ~n15626 & ~n16254;
  assign n16260 = ~n16258 & ~n16259;
  assign n16261 = ~pi100 & ~n16260;
  assign n16262 = ~n14616 & n16162;
  assign n16263 = ~n16261 & n16262;
  assign n16264 = n14621 & n16159;
  assign n16265 = n16226 & ~n16264;
  assign n16266 = ~n16263 & n16265;
  assign n16267 = ~po1038 & ~n16266;
  assign n16268 = ~n16229 & n16267;
  assign n16269 = n14330 & n16226;
  assign n16270 = ~n14330 & n16214;
  assign n16271 = n16045 & ~n16270;
  assign n16272 = ~n16269 & n16271;
  assign po292 = n16268 | n16272;
  assign n16274 = pi136 & ~n15674;
  assign n16275 = ~n16041 & ~n16274;
  assign n16276 = ~n14344 & ~n16275;
  assign n16277 = ~n14396 & n16276;
  assign n16278 = pi148 & n7462;
  assign n16279 = ~n14330 & ~n16278;
  assign n16280 = ~n16277 & ~n16279;
  assign n16281 = n16045 & ~n16280;
  assign n16282 = ~n9685 & ~n15732;
  assign n16283 = n9685 & n14453;
  assign n16284 = pi232 & ~n16283;
  assign n16285 = ~n16282 & n16284;
  assign n16286 = n15730 & ~n16285;
  assign n16287 = pi184 & n15687;
  assign n16288 = ~pi184 & n15691;
  assign n16289 = n9683 & ~n16288;
  assign n16290 = ~n16287 & n16289;
  assign n16291 = pi184 & n15714;
  assign n16292 = ~pi141 & ~pi299;
  assign n16293 = ~pi184 & n15717;
  assign n16294 = n16292 & ~n16293;
  assign n16295 = ~n16291 & n16294;
  assign n16296 = n8039 & ~n15682;
  assign n16297 = pi163 & n6434;
  assign n16298 = n15679 & n16297;
  assign n16299 = ~n8039 & ~n15310;
  assign n16300 = ~n16297 & ~n16299;
  assign n16301 = ~n16298 & ~n16300;
  assign n16302 = pi148 & ~n16301;
  assign n16303 = ~n16296 & n16302;
  assign n16304 = ~pi287 & n13573;
  assign n16305 = pi216 & ~n16304;
  assign n16306 = n6434 & ~n16305;
  assign n16307 = n14538 & n16306;
  assign n16308 = ~pi51 & ~pi148;
  assign n16309 = ~n16307 & n16308;
  assign n16310 = pi299 & ~n16309;
  assign n16311 = ~n16303 & n16310;
  assign n16312 = ~n16295 & ~n16311;
  assign n16313 = ~n16290 & n16312;
  assign n16314 = pi232 & ~n16313;
  assign n16315 = n15727 & ~n16314;
  assign n16316 = n3206 & ~n16315;
  assign n16317 = ~n16286 & n16316;
  assign n16318 = n9686 & ~n14330;
  assign n16319 = ~pi51 & ~n16318;
  assign n16320 = ~n3206 & ~n16319;
  assign n16321 = n3278 & ~n16320;
  assign n16322 = ~n16317 & n16321;
  assign n16323 = n14621 & n16319;
  assign n16324 = n16276 & ~n16323;
  assign n16325 = ~n16322 & n16324;
  assign n16326 = ~n11066 & ~n14330;
  assign n16327 = n16319 & n16326;
  assign n16328 = n9028 & n15627;
  assign n16329 = ~n6162 & n15640;
  assign n16330 = pi148 & ~n16329;
  assign n16331 = ~n16328 & n16330;
  assign n16332 = ~pi51 & n15183;
  assign n16333 = ~pi148 & ~n16332;
  assign n16334 = ~n16304 & ~n16333;
  assign n16335 = ~pi148 & n14396;
  assign n16336 = ~n16334 & ~n16335;
  assign n16337 = ~n16331 & ~n16336;
  assign n16338 = pi299 & ~n16337;
  assign n16339 = pi184 & n15160;
  assign n16340 = n15646 & ~n16339;
  assign n16341 = n16292 & ~n16340;
  assign n16342 = pi184 & n14550;
  assign n16343 = n15650 & ~n16342;
  assign n16344 = n9683 & ~n16343;
  assign n16345 = ~n16341 & ~n16344;
  assign n16346 = ~n16338 & n16345;
  assign n16347 = pi232 & ~n16346;
  assign n16348 = ~pi100 & n15626;
  assign n16349 = ~n16347 & n16348;
  assign n16350 = ~n16327 & ~n16349;
  assign n16351 = n3278 & ~n16350;
  assign n16352 = ~n14330 & n16323;
  assign n16353 = ~n16276 & ~n16352;
  assign n16354 = ~n16351 & n16353;
  assign n16355 = ~po1038 & ~n16354;
  assign n16356 = ~n16325 & n16355;
  assign po293 = n16281 | n16356;
  assign n16358 = ~pi39 & pi137;
  assign n16359 = n10376 & n14755;
  assign n16360 = n6142 & n11506;
  assign n16361 = ~pi299 & ~po1038;
  assign n16362 = ~pi198 & n11517;
  assign n16363 = n16361 & n16362;
  assign n16364 = ~n16360 & ~n16363;
  assign n16365 = ~n16359 & ~n16364;
  assign n16366 = ~pi210 & n11506;
  assign n16367 = po1038 & n16366;
  assign n16368 = ~n16365 & ~n16367;
  assign n16369 = n10420 & ~n16368;
  assign po294 = n16358 | n16369;
  assign n16371 = ~n9415 & n9465;
  assign n16372 = pi92 & ~n16371;
  assign n16373 = n3265 & ~n16372;
  assign n16374 = ~pi75 & ~n9406;
  assign n16375 = ~pi299 & ~n9733;
  assign n16376 = pi299 & ~n9358;
  assign n16377 = ~pi232 & ~n16376;
  assign n16378 = ~n16375 & n16377;
  assign n16379 = ~pi39 & ~n16378;
  assign n16380 = pi148 & n6162;
  assign n16381 = ~n9358 & ~n16380;
  assign n16382 = pi148 & n13630;
  assign n16383 = ~n16381 & ~n16382;
  assign n16384 = pi299 & ~n16383;
  assign n16385 = ~n6162 & ~n9733;
  assign n16386 = ~n13653 & ~n16385;
  assign n16387 = ~pi299 & ~n16386;
  assign n16388 = pi141 & n16387;
  assign n16389 = ~pi141 & n16375;
  assign n16390 = pi232 & ~n16389;
  assign n16391 = ~n16388 & n16390;
  assign n16392 = ~n16384 & n16391;
  assign n16393 = n16379 & ~n16392;
  assign n16394 = ~n9033 & ~n11924;
  assign n16395 = n9053 & ~n16394;
  assign n16396 = n13702 & ~n16395;
  assign n16397 = ~n6189 & ~n9033;
  assign n16398 = n9028 & ~n16394;
  assign n16399 = ~n16397 & n16398;
  assign n16400 = n9030 & ~n16399;
  assign n16401 = ~n16396 & ~n16400;
  assign n16402 = ~pi232 & ~n16401;
  assign n16403 = ~n9038 & ~n16394;
  assign n16404 = ~n9029 & ~n16403;
  assign n16405 = pi148 & ~n16404;
  assign n16406 = ~n9684 & ~n16400;
  assign n16407 = ~n16405 & ~n16406;
  assign n16408 = ~pi141 & n16396;
  assign n16409 = ~n9061 & n16395;
  assign n16410 = n13702 & ~n16409;
  assign n16411 = pi141 & n16410;
  assign n16412 = ~n16408 & ~n16411;
  assign n16413 = ~n16407 & n16412;
  assign n16414 = pi232 & ~n16413;
  assign n16415 = ~n16402 & ~n16414;
  assign n16416 = pi39 & ~n16415;
  assign n16417 = n3206 & ~n16416;
  assign n16418 = ~n16393 & n16417;
  assign n16419 = ~pi87 & ~n16418;
  assign n16420 = n16374 & ~n16419;
  assign n16421 = ~pi92 & ~n16420;
  assign n16422 = n16373 & ~n16421;
  assign n16423 = ~pi55 & ~n16422;
  assign n16424 = n9466 & ~n13739;
  assign n16425 = pi55 & ~n16424;
  assign n16426 = ~n16423 & ~n16425;
  assign n16427 = n3293 & ~n16426;
  assign n16428 = n9666 & ~n16427;
  assign n16429 = pi138 & n16428;
  assign n16430 = ~pi232 & ~n11414;
  assign n16431 = ~n9683 & ~n11414;
  assign n16432 = n6198 & n6451;
  assign n16433 = n9017 & n16432;
  assign n16434 = n9683 & ~n16433;
  assign n16435 = ~n6198 & n9684;
  assign n16436 = ~n16434 & ~n16435;
  assign n16437 = ~n16431 & n16436;
  assign n16438 = pi232 & ~n16437;
  assign n16439 = ~n16430 & ~n16438;
  assign n16440 = pi39 & ~n16439;
  assign n16441 = ~n9686 & n13809;
  assign n16442 = ~pi39 & ~n16441;
  assign n16443 = n10146 & ~n16442;
  assign n16444 = ~n16440 & n16443;
  assign n16445 = ~pi138 & n16444;
  assign n16446 = ~pi118 & n13757;
  assign n16447 = ~pi139 & n16446;
  assign n16448 = ~n16445 & ~n16447;
  assign n16449 = ~n16429 & n16448;
  assign n16450 = ~pi138 & ~n8933;
  assign n16451 = n16428 & n16450;
  assign n16452 = n16444 & ~n16450;
  assign n16453 = n16447 & ~n16452;
  assign n16454 = ~n16451 & n16453;
  assign po295 = ~n16449 & ~n16454;
  assign n16456 = ~n9358 & ~n15634;
  assign n16457 = pi169 & n13630;
  assign n16458 = ~n16456 & ~n16457;
  assign n16459 = pi299 & ~n16458;
  assign n16460 = pi191 & n16387;
  assign n16461 = ~pi191 & n16375;
  assign n16462 = pi232 & ~n16461;
  assign n16463 = ~n16460 & n16462;
  assign n16464 = ~n16459 & n16463;
  assign n16465 = n16379 & ~n16464;
  assign n16466 = pi191 & n16410;
  assign n16467 = ~pi169 & n9033;
  assign n16468 = ~n16403 & ~n16467;
  assign n16469 = n9028 & ~n16468;
  assign n16470 = n9030 & ~n16469;
  assign n16471 = ~pi191 & n16396;
  assign n16472 = ~n16470 & ~n16471;
  assign n16473 = ~n16466 & n16472;
  assign n16474 = pi232 & ~n16473;
  assign n16475 = ~n16402 & ~n16474;
  assign n16476 = pi39 & ~n16475;
  assign n16477 = n3206 & ~n16476;
  assign n16478 = ~n16465 & n16477;
  assign n16479 = ~pi87 & ~n16478;
  assign n16480 = n16374 & ~n16479;
  assign n16481 = ~pi92 & ~n16480;
  assign n16482 = n16373 & ~n16481;
  assign n16483 = ~pi55 & ~n16482;
  assign n16484 = ~n16425 & ~n16483;
  assign n16485 = n3293 & ~n16484;
  assign n16486 = n9666 & ~n16485;
  assign n16487 = pi139 & n16486;
  assign n16488 = ~n6198 & n8970;
  assign n16489 = ~n11413 & ~n16488;
  assign n16490 = ~n11410 & n15645;
  assign n16491 = n8969 & ~n16433;
  assign n16492 = ~n16490 & ~n16491;
  assign n16493 = n16489 & n16492;
  assign n16494 = pi232 & ~n16493;
  assign n16495 = ~n16430 & ~n16494;
  assign n16496 = pi39 & ~n16495;
  assign n16497 = n13809 & ~n15658;
  assign n16498 = ~pi39 & ~n16497;
  assign n16499 = n10146 & ~n16498;
  assign n16500 = ~n16496 & n16499;
  assign n16501 = ~pi139 & n16500;
  assign n16502 = ~n16446 & ~n16501;
  assign n16503 = ~n16487 & n16502;
  assign n16504 = ~pi139 & ~n8934;
  assign n16505 = n16486 & n16504;
  assign n16506 = n16500 & ~n16504;
  assign n16507 = n16446 & ~n16506;
  assign n16508 = ~n16505 & n16507;
  assign po296 = ~n16503 & ~n16508;
  assign n16510 = pi140 & ~n3267;
  assign n16511 = ~pi661 & ~pi681;
  assign n16512 = ~pi662 & n16511;
  assign n16513 = pi680 & ~n16512;
  assign n16514 = ~n6166 & n6435;
  assign n16515 = ~pi120 & ~n16514;
  assign n16516 = pi120 & ~n3095;
  assign n16517 = ~n16515 & ~n16516;
  assign n16518 = n2754 & n16517;
  assign n16519 = pi665 & pi1091;
  assign n16520 = pi621 & pi1091;
  assign n16521 = pi603 & ~n16520;
  assign n16522 = ~n16519 & ~n16521;
  assign n16523 = n16518 & ~n16522;
  assign n16524 = pi616 & ~n16523;
  assign n16525 = pi614 & ~n16523;
  assign n16526 = pi642 & ~n16523;
  assign n16527 = n2754 & n16514;
  assign n16528 = ~pi120 & ~n16527;
  assign n16529 = n2754 & n3095;
  assign n16530 = n6169 & n14187;
  assign n16531 = n16529 & ~n16530;
  assign n16532 = pi120 & ~n16531;
  assign n16533 = pi1091 & ~n16532;
  assign n16534 = ~n16528 & n16533;
  assign n16535 = pi665 & n16534;
  assign n16536 = pi120 & ~n16529;
  assign n16537 = ~pi1091 & ~n16536;
  assign n16538 = pi120 & pi824;
  assign n16539 = n6169 & n16538;
  assign n16540 = n16537 & ~n16539;
  assign n16541 = ~n16528 & n16540;
  assign n16542 = ~n16534 & ~n16541;
  assign n16543 = n16518 & n16521;
  assign n16544 = ~n16542 & n16543;
  assign n16545 = ~n16535 & ~n16544;
  assign n16546 = ~n6162 & n16518;
  assign n16547 = n16519 & n16546;
  assign n16548 = ~pi603 & n16547;
  assign n16549 = n16545 & ~n16548;
  assign n16550 = ~n6162 & n16542;
  assign n16551 = n16543 & ~n16550;
  assign n16552 = n16518 & n16519;
  assign n16553 = n6162 & ~n16552;
  assign n16554 = ~n6162 & ~n16535;
  assign n16555 = ~n16553 & ~n16554;
  assign n16556 = ~pi642 & ~n16555;
  assign n16557 = ~n16551 & n16556;
  assign n16558 = n16549 & n16557;
  assign n16559 = ~n16526 & ~n16558;
  assign n16560 = ~pi614 & ~n16559;
  assign n16561 = ~n16525 & ~n16560;
  assign n16562 = ~pi616 & ~n16561;
  assign n16563 = ~n16524 & ~n16562;
  assign n16564 = n16513 & ~n16563;
  assign n16565 = pi616 & ~n16518;
  assign n16566 = pi614 & ~n16518;
  assign n16567 = ~n6155 & ~n16518;
  assign n16568 = n6162 & ~n16518;
  assign n16569 = ~n16550 & ~n16568;
  assign n16570 = n6155 & ~n16569;
  assign n16571 = ~n16567 & ~n16570;
  assign n16572 = ~pi614 & ~n16571;
  assign n16573 = ~n16566 & ~n16572;
  assign n16574 = ~pi616 & ~n16573;
  assign n16575 = ~n16565 & ~n16574;
  assign n16576 = ~pi680 & ~n16575;
  assign n16577 = n6160 & ~n16555;
  assign n16578 = ~n16551 & n16577;
  assign n16579 = ~n16576 & ~n16578;
  assign n16580 = ~n16564 & n16579;
  assign n16581 = n6215 & ~n16580;
  assign n16582 = n6162 & ~n16542;
  assign n16583 = ~n16546 & ~n16582;
  assign n16584 = ~n6157 & ~n16583;
  assign n16585 = n16542 & ~n16584;
  assign n16586 = ~pi680 & n16585;
  assign n16587 = n6160 & n16545;
  assign n16588 = n16543 & ~n16583;
  assign n16589 = ~n16535 & ~n16547;
  assign n16590 = ~n16588 & n16589;
  assign n16591 = ~pi614 & ~pi642;
  assign n16592 = ~pi616 & n16591;
  assign n16593 = n16549 & n16592;
  assign n16594 = ~n16590 & ~n16593;
  assign n16595 = n16513 & ~n16594;
  assign n16596 = ~n16587 & ~n16595;
  assign n16597 = ~n16586 & n16596;
  assign n16598 = ~n6215 & ~n16597;
  assign n16599 = pi223 & ~n16598;
  assign n16600 = ~n16581 & n16599;
  assign n16601 = ~pi603 & ~n16518;
  assign n16602 = ~pi824 & ~n16514;
  assign n16603 = n6435 & ~n10149;
  assign n16604 = pi1092 & n16603;
  assign n16605 = ~n10972 & ~n16604;
  assign n16606 = ~n16602 & ~n16605;
  assign n16607 = pi1093 & n16606;
  assign n16608 = ~pi120 & ~n16607;
  assign n16609 = n16537 & ~n16608;
  assign n16610 = n2733 & n16527;
  assign n16611 = ~pi829 & ~n16606;
  assign n16612 = pi829 & ~n16604;
  assign n16613 = n7473 & ~n16612;
  assign n16614 = ~n16611 & n16613;
  assign n16615 = ~n16610 & ~n16614;
  assign n16616 = pi1091 & ~n16615;
  assign n16617 = ~pi120 & ~n16616;
  assign n16618 = ~n16536 & ~n16617;
  assign n16619 = ~n16609 & ~n16618;
  assign n16620 = ~n6162 & n16619;
  assign n16621 = ~n16568 & ~n16620;
  assign n16622 = pi603 & ~n16621;
  assign n16623 = ~n16601 & ~n16622;
  assign n16624 = ~n16522 & n16623;
  assign n16625 = ~pi642 & ~n16624;
  assign n16626 = ~n16526 & ~n16625;
  assign n16627 = ~pi614 & ~n16626;
  assign n16628 = ~n16525 & ~n16627;
  assign n16629 = ~pi616 & ~n16628;
  assign n16630 = ~n16524 & ~n16629;
  assign n16631 = n16513 & ~n16630;
  assign n16632 = ~pi642 & ~n16623;
  assign n16633 = ~n16567 & ~n16632;
  assign n16634 = ~pi614 & ~n16633;
  assign n16635 = ~n16566 & ~n16634;
  assign n16636 = ~pi616 & ~n16635;
  assign n16637 = ~n16565 & ~n16636;
  assign n16638 = ~pi680 & ~n16637;
  assign n16639 = n16519 & n16618;
  assign n16640 = ~n6162 & ~n16639;
  assign n16641 = ~n16553 & ~n16640;
  assign n16642 = n16521 & n16621;
  assign n16643 = ~n16641 & ~n16642;
  assign n16644 = n6160 & n16643;
  assign n16645 = ~n16638 & ~n16644;
  assign n16646 = ~n16631 & n16645;
  assign n16647 = n6215 & n16646;
  assign n16648 = n6162 & ~n16619;
  assign n16649 = ~n16546 & ~n16648;
  assign n16650 = ~n6157 & n16649;
  assign n16651 = n6157 & n16619;
  assign n16652 = ~n16650 & ~n16651;
  assign n16653 = ~n16522 & n16652;
  assign n16654 = n16513 & ~n16653;
  assign n16655 = ~pi680 & ~n16652;
  assign n16656 = ~n16520 & ~n16619;
  assign n16657 = pi603 & n16656;
  assign n16658 = pi603 & ~pi621;
  assign n16659 = n16639 & ~n16658;
  assign n16660 = n6160 & ~n16659;
  assign n16661 = ~n16657 & n16660;
  assign n16662 = ~n16655 & ~n16661;
  assign n16663 = ~n16654 & n16662;
  assign n16664 = ~n6215 & n16663;
  assign n16665 = ~n3052 & ~n16664;
  assign n16666 = ~n16647 & n16665;
  assign n16667 = pi680 & n16522;
  assign n16668 = n16518 & ~n16667;
  assign n16669 = n3052 & ~n16668;
  assign n16670 = ~pi223 & ~n16669;
  assign n16671 = ~n16666 & n16670;
  assign n16672 = ~n16600 & ~n16671;
  assign n16673 = ~pi299 & ~n16672;
  assign n16674 = ~n6189 & ~n16663;
  assign n16675 = n6189 & ~n16646;
  assign n16676 = ~n16674 & ~n16675;
  assign n16677 = ~n3329 & ~n16676;
  assign n16678 = n3329 & ~n16668;
  assign n16679 = ~pi215 & ~n16678;
  assign n16680 = ~n16677 & n16679;
  assign n16681 = n6189 & ~n16580;
  assign n16682 = ~n6189 & ~n16597;
  assign n16683 = pi215 & ~n16682;
  assign n16684 = ~n16681 & n16683;
  assign n16685 = ~n16680 & ~n16684;
  assign n16686 = pi299 & ~n16685;
  assign n16687 = ~n16673 & ~n16686;
  assign n16688 = ~pi140 & n16687;
  assign n16689 = n16518 & ~n16519;
  assign n16690 = ~n16519 & ~n16619;
  assign n16691 = ~n16689 & ~n16690;
  assign n16692 = ~n16521 & ~n16649;
  assign n16693 = ~n16691 & n16692;
  assign n16694 = pi616 & ~n16693;
  assign n16695 = n16520 & n16618;
  assign n16696 = ~pi665 & n16695;
  assign n16697 = pi603 & ~n16696;
  assign n16698 = ~n16649 & ~n16691;
  assign n16699 = ~pi603 & ~n16698;
  assign n16700 = ~n16697 & ~n16699;
  assign n16701 = n16592 & ~n16700;
  assign n16702 = n16693 & ~n16701;
  assign n16703 = n16591 & n16700;
  assign n16704 = ~pi616 & ~n16703;
  assign n16705 = ~n16702 & n16704;
  assign n16706 = ~n16694 & ~n16705;
  assign n16707 = ~n16512 & ~n16706;
  assign n16708 = n6160 & n16690;
  assign n16709 = ~n16697 & n16708;
  assign n16710 = ~n16513 & ~n16709;
  assign n16711 = ~n16707 & ~n16710;
  assign n16712 = ~n6189 & ~n16711;
  assign n16713 = n16518 & ~n16521;
  assign n16714 = ~n16519 & n16713;
  assign n16715 = pi616 & ~n16714;
  assign n16716 = n16513 & ~n16715;
  assign n16717 = n16518 & n16520;
  assign n16718 = n6162 & ~n16717;
  assign n16719 = ~n6162 & ~n16695;
  assign n16720 = ~n16718 & ~n16719;
  assign n16721 = pi603 & ~n16720;
  assign n16722 = pi603 & pi665;
  assign n16723 = ~pi603 & ~n16689;
  assign n16724 = ~n16722 & ~n16723;
  assign n16725 = ~n16721 & n16724;
  assign n16726 = n16591 & n16725;
  assign n16727 = ~n16591 & n16714;
  assign n16728 = ~pi616 & ~n16727;
  assign n16729 = ~n16726 & n16728;
  assign n16730 = n16716 & ~n16729;
  assign n16731 = n16621 & n16644;
  assign n16732 = ~n16730 & ~n16731;
  assign n16733 = n6189 & n16732;
  assign n16734 = ~n3329 & ~n16733;
  assign n16735 = ~n16712 & n16734;
  assign n16736 = n3329 & n16518;
  assign n16737 = ~pi215 & ~n16736;
  assign n16738 = ~n16679 & ~n16737;
  assign n16739 = ~n16735 & ~n16738;
  assign n16740 = n2754 & ~n16521;
  assign n16741 = ~n16583 & n16740;
  assign n16742 = n16724 & n16741;
  assign n16743 = pi616 & ~n16742;
  assign n16744 = pi614 & ~pi616;
  assign n16745 = ~n16742 & n16744;
  assign n16746 = pi621 & n16534;
  assign n16747 = ~n6162 & ~n16746;
  assign n16748 = ~n16718 & ~n16747;
  assign n16749 = pi603 & ~n16748;
  assign n16750 = n16724 & ~n16749;
  assign n16751 = ~pi642 & ~n16750;
  assign n16752 = n16742 & ~n16751;
  assign n16753 = n6156 & ~n16752;
  assign n16754 = ~n16745 & ~n16753;
  assign n16755 = ~n16743 & n16754;
  assign n16756 = ~n16512 & ~n16755;
  assign n16757 = ~n16542 & n16667;
  assign n16758 = ~n16513 & ~n16757;
  assign n16759 = ~n16756 & ~n16758;
  assign n16760 = ~n6189 & n16759;
  assign n16761 = ~n16592 & n16713;
  assign n16762 = n16592 & ~n16601;
  assign n16763 = ~n16749 & n16762;
  assign n16764 = ~n16761 & ~n16763;
  assign n16765 = ~n16519 & ~n16764;
  assign n16766 = ~pi616 & ~n16765;
  assign n16767 = n16716 & ~n16766;
  assign n16768 = n6160 & n16569;
  assign n16769 = ~n16749 & n16768;
  assign n16770 = n16724 & n16769;
  assign n16771 = ~n16767 & ~n16770;
  assign n16772 = n6189 & ~n16771;
  assign n16773 = pi215 & ~n16772;
  assign n16774 = ~n16760 & n16773;
  assign n16775 = ~n16739 & ~n16774;
  assign n16776 = pi299 & ~n16775;
  assign n16777 = ~n6215 & n16711;
  assign n16778 = n6215 & ~n16732;
  assign n16779 = ~n3052 & ~n16778;
  assign n16780 = ~n16777 & n16779;
  assign n16781 = n3052 & n16518;
  assign n16782 = n16521 & n16781;
  assign n16783 = ~pi223 & ~n16782;
  assign n16784 = n2754 & n16521;
  assign n16785 = pi680 & ~n16519;
  assign n16786 = n2754 & n16785;
  assign n16787 = ~n16521 & n16786;
  assign n16788 = ~n16784 & ~n16787;
  assign n16789 = n16518 & ~n16788;
  assign n16790 = n3052 & ~n16789;
  assign n16791 = n16783 & ~n16790;
  assign n16792 = ~n16780 & n16791;
  assign n16793 = ~n6215 & ~n16759;
  assign n16794 = n6215 & n16771;
  assign n16795 = pi223 & ~n16794;
  assign n16796 = ~n16793 & n16795;
  assign n16797 = ~pi299 & ~n16796;
  assign n16798 = ~n16792 & n16797;
  assign n16799 = ~n16776 & ~n16798;
  assign n16800 = pi140 & n16799;
  assign n16801 = pi761 & ~n16800;
  assign n16802 = ~n16688 & n16801;
  assign n16803 = ~n16657 & ~n16700;
  assign n16804 = n16592 & ~n16803;
  assign n16805 = n16521 & ~n16649;
  assign n16806 = ~n16698 & ~n16805;
  assign n16807 = ~n16592 & ~n16806;
  assign n16808 = n16513 & ~n16807;
  assign n16809 = ~n16804 & n16808;
  assign n16810 = ~n6160 & ~n16652;
  assign n16811 = n6160 & n16619;
  assign n16812 = ~n16810 & ~n16811;
  assign n16813 = n16521 & n16812;
  assign n16814 = ~n16513 & ~n16708;
  assign n16815 = ~n16813 & n16814;
  assign n16816 = ~n16809 & ~n16815;
  assign n16817 = ~n6215 & n16816;
  assign n16818 = n16519 & ~n16658;
  assign n16819 = n16518 & ~n16818;
  assign n16820 = ~n16592 & n16819;
  assign n16821 = n16513 & ~n16820;
  assign n16822 = ~n16721 & n16762;
  assign n16823 = n16519 & n16822;
  assign n16824 = n16592 & n16623;
  assign n16825 = ~n16823 & n16824;
  assign n16826 = n16821 & ~n16825;
  assign n16827 = n16543 & ~n16592;
  assign n16828 = n16592 & n16642;
  assign n16829 = ~n16827 & ~n16828;
  assign n16830 = ~pi680 & n16829;
  assign n16831 = n16621 & ~n16691;
  assign n16832 = n6160 & ~n16831;
  assign n16833 = ~n16642 & n16832;
  assign n16834 = ~n16830 & ~n16833;
  assign n16835 = ~n16826 & n16834;
  assign n16836 = n6215 & n16835;
  assign n16837 = ~n3052 & ~n16836;
  assign n16838 = ~n16817 & n16837;
  assign n16839 = ~pi223 & ~n16790;
  assign n16840 = ~n16838 & n16839;
  assign n16841 = ~n6157 & n16689;
  assign n16842 = ~n16550 & n16689;
  assign n16843 = ~n16841 & ~n16842;
  assign n16844 = ~n16551 & n16843;
  assign n16845 = n16592 & ~n16844;
  assign n16846 = n16821 & ~n16845;
  assign n16847 = n16550 & n16592;
  assign n16848 = n16588 & ~n16847;
  assign n16849 = ~n6160 & n16848;
  assign n16850 = ~n16551 & ~n16849;
  assign n16851 = n16512 & ~n16842;
  assign n16852 = pi680 & ~n16851;
  assign n16853 = n16850 & ~n16852;
  assign n16854 = ~n16846 & ~n16853;
  assign n16855 = n6215 & ~n16854;
  assign n16856 = ~n16544 & ~n16849;
  assign n16857 = ~n16583 & n16689;
  assign n16858 = ~n16843 & n16852;
  assign n16859 = n16857 & n16858;
  assign n16860 = n16856 & ~n16859;
  assign n16861 = ~n6215 & n16860;
  assign n16862 = pi223 & ~n16861;
  assign n16863 = ~n16855 & n16862;
  assign n16864 = ~pi299 & ~n16863;
  assign n16865 = ~n16840 & n16864;
  assign n16866 = ~n6189 & n16816;
  assign n16867 = n6189 & n16835;
  assign n16868 = ~n16866 & ~n16867;
  assign n16869 = ~n3329 & ~n16868;
  assign n16870 = n3329 & n16789;
  assign n16871 = ~pi215 & ~n16870;
  assign n16872 = ~n16869 & n16871;
  assign n16873 = n6189 & n16854;
  assign n16874 = ~n6189 & ~n16860;
  assign n16875 = pi215 & ~n16874;
  assign n16876 = ~n16873 & n16875;
  assign n16877 = ~n16872 & ~n16876;
  assign n16878 = pi299 & ~n16877;
  assign n16879 = ~n16865 & ~n16878;
  assign n16880 = pi140 & n16879;
  assign n16881 = ~n16521 & n16652;
  assign n16882 = ~pi680 & ~n16881;
  assign n16883 = ~n6191 & n16639;
  assign n16884 = ~n6157 & n16547;
  assign n16885 = ~n16883 & ~n16884;
  assign n16886 = n16818 & ~n16885;
  assign n16887 = n16513 & ~n16886;
  assign n16888 = ~n16660 & ~n16887;
  assign n16889 = ~n16882 & n16888;
  assign n16890 = ~n6215 & n16889;
  assign n16891 = n16552 & ~n16658;
  assign n16892 = ~n16592 & n16891;
  assign n16893 = n16513 & ~n16892;
  assign n16894 = ~n16823 & n16893;
  assign n16895 = ~n16761 & ~n16822;
  assign n16896 = ~pi680 & n16895;
  assign n16897 = n16641 & n16818;
  assign n16898 = n6160 & ~n16897;
  assign n16899 = ~n16896 & ~n16898;
  assign n16900 = ~n16894 & n16899;
  assign n16901 = n6215 & n16900;
  assign n16902 = ~n16890 & ~n16901;
  assign n16903 = ~n3052 & ~n16902;
  assign n16904 = ~n16521 & ~n16785;
  assign n16905 = n16529 & n16904;
  assign n16906 = ~n16515 & n16905;
  assign n16907 = n3052 & n16906;
  assign n16908 = ~pi223 & ~n16907;
  assign n16909 = ~n16903 & n16908;
  assign n16910 = ~n16589 & ~n16764;
  assign n16911 = n16513 & ~n16910;
  assign n16912 = n6157 & ~n16534;
  assign n16913 = n16741 & ~n16912;
  assign n16914 = ~pi680 & ~n16913;
  assign n16915 = pi680 & ~n16535;
  assign n16916 = ~n16658 & ~n16915;
  assign n16917 = n6160 & ~n16916;
  assign n16918 = ~n16914 & ~n16917;
  assign n16919 = ~n16911 & n16918;
  assign n16920 = ~n6215 & n16919;
  assign n16921 = ~n6160 & ~n16764;
  assign n16922 = ~n16785 & n16921;
  assign n16923 = n6160 & ~n16658;
  assign n16924 = n16555 & n16923;
  assign n16925 = ~n16922 & ~n16924;
  assign n16926 = n6215 & ~n16925;
  assign n16927 = pi223 & ~n16926;
  assign n16928 = ~n16920 & n16927;
  assign n16929 = ~n16909 & ~n16928;
  assign n16930 = ~pi299 & ~n16929;
  assign n16931 = ~n6189 & n16889;
  assign n16932 = n6189 & n16900;
  assign n16933 = ~n16931 & ~n16932;
  assign n16934 = ~n3329 & ~n16933;
  assign n16935 = n3329 & n16906;
  assign n16936 = ~pi215 & ~n16935;
  assign n16937 = ~n16934 & n16936;
  assign n16938 = ~n6189 & n16919;
  assign n16939 = n6189 & ~n16925;
  assign n16940 = pi215 & ~n16939;
  assign n16941 = ~n16938 & n16940;
  assign n16942 = ~n16937 & ~n16941;
  assign n16943 = pi299 & ~n16942;
  assign n16944 = ~n16930 & ~n16943;
  assign n16945 = ~pi140 & ~n16944;
  assign n16946 = ~pi761 & ~n16945;
  assign n16947 = ~n16880 & n16946;
  assign n16948 = ~n16802 & ~n16947;
  assign n16949 = pi39 & ~n16948;
  assign n16950 = ~pi102 & ~n11239;
  assign n16951 = ~pi98 & ~n2596;
  assign n16952 = ~n16950 & n16951;
  assign n16953 = n7429 & n12123;
  assign n16954 = n16952 & n16953;
  assign n16955 = n8859 & n9127;
  assign n16956 = n16954 & n16955;
  assign n16957 = ~pi40 & ~n16956;
  assign n16958 = n10227 & ~n16957;
  assign n16959 = ~pi252 & ~n16958;
  assign n16960 = n2536 & n2572;
  assign n16961 = n8858 & n16954;
  assign n16962 = ~pi47 & ~n16961;
  assign n16963 = pi314 & n10202;
  assign n16964 = n16962 & ~n16963;
  assign n16965 = n16960 & ~n16964;
  assign n16966 = ~pi35 & ~n16965;
  assign n16967 = ~pi40 & n10220;
  assign n16968 = ~n16966 & n16967;
  assign n16969 = pi252 & ~n2553;
  assign n16970 = ~n16968 & n16969;
  assign n16971 = ~n16959 & ~n16970;
  assign n16972 = n3092 & n16971;
  assign n16973 = pi1092 & ~n12135;
  assign n16974 = n16972 & n16973;
  assign n16975 = ~pi88 & ~n16952;
  assign n16976 = n10946 & ~n16975;
  assign n16977 = n2519 & n16976;
  assign n16978 = ~pi47 & ~n16963;
  assign n16979 = ~n16977 & n16978;
  assign n16980 = n16960 & ~n16979;
  assign n16981 = ~pi35 & ~n16980;
  assign n16982 = pi252 & n10220;
  assign n16983 = ~n16981 & n16982;
  assign n16984 = ~pi252 & n9269;
  assign n16985 = n16976 & n16984;
  assign n16986 = ~pi40 & ~n16985;
  assign n16987 = ~n16983 & n16986;
  assign n16988 = n7474 & n10227;
  assign n16989 = ~n16987 & n16988;
  assign n16990 = ~n16974 & ~n16989;
  assign n16991 = pi1093 & ~n16990;
  assign n16992 = ~n2733 & ~n16991;
  assign n16993 = pi1092 & n10018;
  assign po1106 = n2733 & n16993;
  assign n16995 = n16972 & po1106;
  assign n16996 = ~n2734 & ~n16995;
  assign n16997 = ~n16992 & ~n16996;
  assign n16998 = pi621 & n16997;
  assign n16999 = ~pi210 & ~n16998;
  assign n17000 = ~n3359 & ~n16987;
  assign n17001 = ~pi32 & ~n17000;
  assign n17002 = pi32 & ~n6366;
  assign n17003 = ~pi95 & n6257;
  assign n17004 = ~n17002 & n17003;
  assign n17005 = ~n17001 & n17004;
  assign n17006 = pi824 & n17005;
  assign n17007 = ~n16974 & ~n17006;
  assign n17008 = ~pi32 & ~n16971;
  assign n17009 = n17004 & ~n17008;
  assign n17010 = ~pi824 & pi829;
  assign n17011 = n17009 & n17010;
  assign n17012 = n17007 & ~n17011;
  assign n17013 = pi1093 & ~n17012;
  assign n17014 = ~n2733 & ~n17013;
  assign n17015 = ~n16996 & ~n17014;
  assign n17016 = pi621 & n17015;
  assign n17017 = pi210 & ~n17016;
  assign n17018 = ~n16999 & ~n17017;
  assign n17019 = pi603 & ~n17018;
  assign n17020 = ~pi1091 & n16991;
  assign n17021 = ~n16997 & ~n17020;
  assign n17022 = ~pi210 & n17021;
  assign n17023 = n7536 & ~n17007;
  assign n17024 = ~n17015 & ~n17023;
  assign n17025 = pi210 & n17024;
  assign n17026 = ~n17022 & ~n17025;
  assign n17027 = ~n17019 & n17026;
  assign n17028 = pi299 & ~n17027;
  assign n17029 = ~pi198 & ~n16998;
  assign n17030 = pi198 & ~n17016;
  assign n17031 = ~n17029 & ~n17030;
  assign n17032 = pi621 & ~n17020;
  assign n17033 = ~n17021 & ~n17032;
  assign n17034 = ~pi198 & n17033;
  assign n17035 = pi621 & ~n17023;
  assign n17036 = ~n17024 & ~n17035;
  assign n17037 = pi198 & n17036;
  assign n17038 = ~n17034 & ~n17037;
  assign n17039 = ~pi603 & ~n17038;
  assign n17040 = ~n17031 & ~n17039;
  assign n17041 = ~pi299 & n17040;
  assign n17042 = ~n17028 & ~n17041;
  assign n17043 = pi665 & ~n17020;
  assign n17044 = ~n17021 & ~n17043;
  assign n17045 = ~pi198 & ~n17044;
  assign n17046 = pi665 & ~n17023;
  assign n17047 = ~n17024 & ~n17046;
  assign n17048 = pi198 & ~n17047;
  assign n17049 = ~n17045 & ~n17048;
  assign n17050 = pi680 & n17049;
  assign n17051 = ~pi299 & ~n17050;
  assign n17052 = pi210 & ~n17047;
  assign n17053 = ~pi210 & ~n17044;
  assign n17054 = ~n17052 & ~n17053;
  assign n17055 = pi680 & n17054;
  assign n17056 = pi299 & ~n17055;
  assign n17057 = ~n17051 & ~n17056;
  assign n17058 = ~n16722 & n17057;
  assign n17059 = n17042 & n17058;
  assign n17060 = pi140 & ~n17059;
  assign n17061 = ~pi198 & n17021;
  assign n17062 = pi198 & n17024;
  assign n17063 = ~n17061 & ~n17062;
  assign n17064 = pi665 & n17015;
  assign n17065 = pi198 & ~n17064;
  assign n17066 = pi665 & n16997;
  assign n17067 = ~pi198 & ~n17066;
  assign n17068 = ~n17065 & ~n17067;
  assign n17069 = pi680 & ~n17068;
  assign n17070 = n17063 & ~n17069;
  assign n17071 = ~pi299 & ~n17070;
  assign n17072 = ~pi210 & ~n17066;
  assign n17073 = pi210 & ~n17064;
  assign n17074 = ~n17072 & ~n17073;
  assign n17075 = pi680 & ~n17074;
  assign n17076 = n17026 & ~n17075;
  assign n17077 = pi299 & ~n17076;
  assign n17078 = ~n17071 & ~n17077;
  assign n17079 = pi603 & ~n17038;
  assign n17080 = ~pi299 & ~n17079;
  assign n17081 = ~pi210 & ~n17033;
  assign n17082 = pi210 & ~n17036;
  assign n17083 = ~n17081 & ~n17082;
  assign n17084 = pi603 & n17083;
  assign n17085 = pi299 & ~n17084;
  assign n17086 = ~n17080 & ~n17085;
  assign n17087 = pi680 & n17086;
  assign n17088 = ~n17078 & ~n17087;
  assign n17089 = ~pi140 & ~n17088;
  assign n17090 = pi761 & ~n17089;
  assign n17091 = ~n17060 & n17090;
  assign n17092 = n17042 & n17078;
  assign n17093 = ~pi140 & n17092;
  assign n17094 = ~n17057 & ~n17086;
  assign n17095 = pi140 & n17094;
  assign n17096 = ~pi761 & ~n17095;
  assign n17097 = ~n17093 & n17096;
  assign n17098 = ~pi39 & ~n17097;
  assign n17099 = ~n17091 & n17098;
  assign n17100 = ~pi38 & ~n17099;
  assign n17101 = ~n16949 & n17100;
  assign n17102 = ~pi140 & ~n16905;
  assign n17103 = pi140 & ~n16788;
  assign n17104 = n3095 & n17103;
  assign n17105 = ~pi761 & ~n17104;
  assign n17106 = ~n17102 & n17105;
  assign n17107 = n16529 & n16667;
  assign n17108 = ~pi140 & ~n16529;
  assign n17109 = pi761 & ~n17108;
  assign n17110 = ~n17107 & n17109;
  assign n17111 = ~n17106 & ~n17110;
  assign n17112 = ~pi39 & ~n17111;
  assign n17113 = pi39 & pi140;
  assign n17114 = pi38 & ~n17113;
  assign n17115 = ~n17112 & n17114;
  assign n17116 = ~n17101 & ~n17115;
  assign n17117 = ~pi738 & ~n17116;
  assign n17118 = pi299 & ~n17026;
  assign n17119 = ~pi299 & ~n17063;
  assign n17120 = ~n17118 & ~n17119;
  assign n17121 = ~pi39 & ~n17120;
  assign n17122 = pi681 & n16585;
  assign n17123 = ~n6158 & ~n16575;
  assign n17124 = n6158 & n16542;
  assign n17125 = ~n6162 & ~n17124;
  assign n17126 = ~n17123 & n17125;
  assign n17127 = ~n16582 & ~n17126;
  assign n17128 = ~pi661 & ~n17127;
  assign n17129 = pi661 & ~n16585;
  assign n17130 = ~pi681 & ~n17129;
  assign n17131 = ~n17128 & n17130;
  assign n17132 = ~n17122 & ~n17131;
  assign n17133 = ~n6215 & ~n17132;
  assign n17134 = pi681 & ~n16575;
  assign n17135 = ~pi616 & ~n16512;
  assign n17136 = n16573 & n17135;
  assign n17137 = pi680 & ~n16569;
  assign n17138 = ~pi616 & n16512;
  assign n17139 = ~n17137 & n17138;
  assign n17140 = ~n16576 & n17139;
  assign n17141 = ~n17136 & ~n17140;
  assign n17142 = ~pi680 & ~n16518;
  assign n17143 = pi616 & n16512;
  assign n17144 = ~n17142 & n17143;
  assign n17145 = ~n17137 & n17144;
  assign n17146 = pi616 & n16518;
  assign n17147 = ~n16512 & n17146;
  assign n17148 = ~n17145 & ~n17147;
  assign n17149 = ~pi681 & n17148;
  assign n17150 = n17141 & n17149;
  assign n17151 = ~n17134 & ~n17150;
  assign n17152 = n6215 & ~n17151;
  assign n17153 = ~n17133 & ~n17152;
  assign n17154 = pi223 & ~n17153;
  assign n17155 = pi681 & ~n16637;
  assign n17156 = ~pi616 & ~n16633;
  assign n17157 = ~pi614 & ~n6160;
  assign n17158 = ~n16565 & n17157;
  assign n17159 = ~n17156 & n17158;
  assign n17160 = ~pi614 & n6160;
  assign n17161 = n16621 & n17160;
  assign n17162 = ~n17159 & ~n17161;
  assign n17163 = pi680 & ~n16621;
  assign n17164 = pi614 & n16512;
  assign n17165 = ~n17142 & n17164;
  assign n17166 = ~n17163 & n17165;
  assign n17167 = pi614 & n16518;
  assign n17168 = ~n16512 & n17167;
  assign n17169 = ~n17166 & ~n17168;
  assign n17170 = ~pi681 & n17169;
  assign n17171 = n17162 & n17170;
  assign n17172 = ~n17155 & ~n17171;
  assign n17173 = n6215 & ~n17172;
  assign n17174 = ~n6215 & ~n16812;
  assign n17175 = ~n17173 & ~n17174;
  assign n17176 = ~n3052 & n17175;
  assign n17177 = ~n16781 & ~n17176;
  assign n17178 = ~pi223 & n17177;
  assign n17179 = ~n17154 & ~n17178;
  assign n17180 = ~pi299 & ~n17179;
  assign n17181 = n6188 & ~n17172;
  assign n17182 = ~n6188 & ~n16812;
  assign n17183 = n6183 & ~n17182;
  assign n17184 = ~n17181 & n17183;
  assign n17185 = ~n3329 & n17184;
  assign n17186 = ~n6183 & n16812;
  assign n17187 = ~n3329 & n17186;
  assign n17188 = n16737 & ~n17187;
  assign n17189 = ~n17185 & n17188;
  assign n17190 = ~n6183 & n17132;
  assign n17191 = ~n6188 & ~n17132;
  assign n17192 = n6188 & ~n17151;
  assign n17193 = n6183 & ~n17192;
  assign n17194 = ~n17191 & n17193;
  assign n17195 = ~n17190 & ~n17194;
  assign n17196 = pi215 & n17195;
  assign n17197 = ~n17189 & ~n17196;
  assign n17198 = pi299 & ~n17197;
  assign n17199 = ~n17180 & ~n17198;
  assign n17200 = pi39 & ~n17199;
  assign n17201 = ~n17121 & ~n17200;
  assign n17202 = pi761 & n17201;
  assign n17203 = ~pi39 & ~n17042;
  assign n17204 = n16621 & ~n16721;
  assign n17205 = n6160 & ~n17204;
  assign n17206 = ~n6160 & n16895;
  assign n17207 = ~n17205 & ~n17206;
  assign n17208 = n6189 & ~n17207;
  assign n17209 = ~n16521 & n16812;
  assign n17210 = ~n6189 & ~n17209;
  assign n17211 = ~n3329 & ~n17210;
  assign n17212 = ~n17208 & n17211;
  assign n17213 = n3329 & n16713;
  assign n17214 = ~n17212 & ~n17213;
  assign n17215 = ~pi215 & ~n17214;
  assign n17216 = ~n16769 & ~n16921;
  assign n17217 = n6189 & n17216;
  assign n17218 = ~n6160 & ~n16913;
  assign n17219 = ~n16542 & n16740;
  assign n17220 = n6160 & ~n17219;
  assign n17221 = ~n17218 & ~n17220;
  assign n17222 = ~n6189 & ~n17221;
  assign n17223 = pi215 & ~n17222;
  assign n17224 = ~n17217 & n17223;
  assign n17225 = ~n17215 & ~n17224;
  assign n17226 = pi299 & ~n17225;
  assign n17227 = n6215 & ~n17207;
  assign n17228 = ~n6215 & ~n17209;
  assign n17229 = ~n3052 & ~n17228;
  assign n17230 = ~n17227 & n17229;
  assign n17231 = n3052 & n16713;
  assign n17232 = ~n17230 & ~n17231;
  assign n17233 = ~pi223 & ~n17232;
  assign n17234 = n6215 & n17216;
  assign n17235 = ~n6215 & ~n17221;
  assign n17236 = pi223 & ~n17235;
  assign n17237 = ~n17234 & n17236;
  assign n17238 = ~n17233 & ~n17237;
  assign n17239 = ~pi299 & ~n17238;
  assign n17240 = ~n17226 & ~n17239;
  assign n17241 = pi39 & n17240;
  assign n17242 = ~n17203 & ~n17241;
  assign n17243 = ~pi761 & n17242;
  assign n17244 = ~pi140 & ~n17243;
  assign n17245 = ~n17202 & n17244;
  assign n17246 = ~pi39 & ~n17086;
  assign n17247 = ~n6189 & ~n16813;
  assign n17248 = n6160 & n16642;
  assign n17249 = ~n6160 & ~n16829;
  assign n17250 = ~n17248 & ~n17249;
  assign n17251 = n6189 & n17250;
  assign n17252 = ~n3329 & ~n17251;
  assign n17253 = ~n17247 & n17252;
  assign n17254 = n3329 & n16517;
  assign n17255 = n16784 & n17254;
  assign n17256 = ~pi215 & ~n17255;
  assign n17257 = ~n17253 & n17256;
  assign n17258 = ~n6189 & n16583;
  assign n17259 = ~n16850 & ~n17258;
  assign n17260 = pi215 & ~n17259;
  assign n17261 = pi299 & ~n17260;
  assign n17262 = ~n17257 & n17261;
  assign n17263 = ~n6215 & ~n16813;
  assign n17264 = n6215 & n17250;
  assign n17265 = ~n3052 & ~n17264;
  assign n17266 = ~n17263 & n17265;
  assign n17267 = n16783 & ~n17266;
  assign n17268 = ~n6215 & n16583;
  assign n17269 = ~n16850 & ~n17268;
  assign n17270 = pi223 & ~n17269;
  assign n17271 = ~pi299 & ~n17270;
  assign n17272 = ~n17267 & n17271;
  assign n17273 = ~n17262 & ~n17272;
  assign n17274 = pi39 & n17273;
  assign n17275 = ~n17246 & ~n17274;
  assign n17276 = pi140 & ~pi761;
  assign n17277 = n17275 & n17276;
  assign n17278 = ~n17245 & ~n17277;
  assign n17279 = ~pi38 & ~n17278;
  assign n17280 = n2754 & n6234;
  assign n17281 = ~pi140 & ~n17280;
  assign n17282 = n6234 & n16784;
  assign n17283 = ~pi761 & n17282;
  assign n17284 = ~n17281 & ~n17283;
  assign n17285 = pi38 & ~n17284;
  assign n17286 = ~n17279 & ~n17285;
  assign n17287 = pi738 & ~n17286;
  assign n17288 = n3267 & ~n17287;
  assign n17289 = ~n17117 & n17288;
  assign n17290 = ~n16510 & ~n17289;
  assign n17291 = ~pi625 & n17290;
  assign n17292 = n3267 & n17286;
  assign n17293 = ~n16510 & ~n17292;
  assign n17294 = pi625 & n17293;
  assign n17295 = ~pi1153 & ~n17294;
  assign n17296 = ~n17291 & n17295;
  assign n17297 = n16781 & n16785;
  assign n17298 = n16652 & n16785;
  assign n17299 = ~n16512 & n17298;
  assign n17300 = ~n16708 & ~n17299;
  assign n17301 = ~n6215 & n17300;
  assign n17302 = n6157 & n16831;
  assign n17303 = ~n16841 & ~n17302;
  assign n17304 = ~n16512 & n17303;
  assign n17305 = n16512 & ~n16831;
  assign n17306 = pi680 & ~n17305;
  assign n17307 = ~n17304 & n17306;
  assign n17308 = n6215 & ~n17307;
  assign n17309 = ~n3052 & ~n17308;
  assign n17310 = ~n17301 & n17309;
  assign n17311 = ~n17297 & ~n17310;
  assign n17312 = ~pi223 & ~n17311;
  assign n17313 = pi680 & ~n16843;
  assign n17314 = ~n17268 & n17313;
  assign n17315 = pi223 & ~n16851;
  assign n17316 = n17314 & n17315;
  assign n17317 = ~n17312 & ~n17316;
  assign n17318 = ~pi299 & ~n17317;
  assign n17319 = n6189 & ~n17307;
  assign n17320 = ~n6189 & n17300;
  assign n17321 = ~n3329 & ~n17320;
  assign n17322 = ~n17319 & n17321;
  assign n17323 = n16518 & n16785;
  assign n17324 = n3329 & n17323;
  assign n17325 = ~n17322 & ~n17324;
  assign n17326 = ~pi215 & ~n17325;
  assign n17327 = ~n17258 & n17313;
  assign n17328 = pi215 & ~n16851;
  assign n17329 = n17327 & n17328;
  assign n17330 = ~n17326 & ~n17329;
  assign n17331 = pi299 & ~n17330;
  assign n17332 = ~n17318 & ~n17331;
  assign n17333 = pi140 & ~n17332;
  assign n17334 = n6157 & n16641;
  assign n17335 = ~n6157 & n16552;
  assign n17336 = pi680 & ~n17335;
  assign n17337 = ~n17334 & n17336;
  assign n17338 = ~n16638 & ~n17337;
  assign n17339 = ~n16512 & n17338;
  assign n17340 = pi680 & ~n16641;
  assign n17341 = n16512 & ~n17340;
  assign n17342 = ~n16638 & n17341;
  assign n17343 = ~n17339 & ~n17342;
  assign n17344 = n6215 & n17343;
  assign n17345 = ~n16512 & ~n16885;
  assign n17346 = n16512 & n16639;
  assign n17347 = pi680 & ~n17346;
  assign n17348 = ~n17345 & n17347;
  assign n17349 = ~n16655 & ~n17348;
  assign n17350 = ~n6215 & ~n17349;
  assign n17351 = ~n3052 & ~n17350;
  assign n17352 = ~n17344 & n17351;
  assign n17353 = n16781 & ~n16785;
  assign n17354 = ~pi223 & ~n17353;
  assign n17355 = ~n17352 & n17354;
  assign n17356 = ~n16555 & n17336;
  assign n17357 = ~n16577 & ~n17356;
  assign n17358 = ~n16585 & ~n16785;
  assign n17359 = n17357 & n17358;
  assign n17360 = ~n6215 & n17359;
  assign n17361 = ~n16576 & n17357;
  assign n17362 = n6215 & n17361;
  assign n17363 = pi223 & ~n17362;
  assign n17364 = ~n17360 & n17363;
  assign n17365 = ~n17355 & ~n17364;
  assign n17366 = ~pi299 & ~n17365;
  assign n17367 = n6189 & n17343;
  assign n17368 = ~n6189 & ~n17349;
  assign n17369 = ~n3329 & ~n17368;
  assign n17370 = ~n17367 & n17369;
  assign n17371 = n2754 & ~n16785;
  assign n17372 = n17254 & n17371;
  assign n17373 = ~pi215 & ~n17372;
  assign n17374 = ~n17370 & n17373;
  assign n17375 = ~n6189 & n17359;
  assign n17376 = n6189 & n17361;
  assign n17377 = pi215 & ~n17376;
  assign n17378 = ~n17375 & n17377;
  assign n17379 = ~n17374 & ~n17378;
  assign n17380 = pi299 & ~n17379;
  assign n17381 = ~n17366 & ~n17380;
  assign n17382 = pi39 & n17381;
  assign n17383 = ~n17113 & ~n17382;
  assign n17384 = ~n17333 & ~n17383;
  assign n17385 = ~pi140 & ~n17078;
  assign n17386 = pi140 & n17057;
  assign n17387 = ~pi39 & ~n17386;
  assign n17388 = ~n17385 & n17387;
  assign n17389 = ~n17384 & ~n17388;
  assign n17390 = ~pi38 & ~n17389;
  assign n17391 = n6234 & n16786;
  assign n17392 = pi38 & ~n17391;
  assign n17393 = ~n17281 & n17392;
  assign n17394 = ~pi738 & ~n17393;
  assign n17395 = ~n17390 & n17394;
  assign n17396 = ~pi38 & ~n17201;
  assign n17397 = n2754 & n6109;
  assign n17398 = pi38 & ~n17397;
  assign n17399 = ~n17396 & ~n17398;
  assign n17400 = ~pi140 & pi738;
  assign n17401 = ~n17399 & n17400;
  assign n17402 = n3267 & ~n17401;
  assign n17403 = ~n17395 & n17402;
  assign n17404 = ~n16510 & ~n17403;
  assign n17405 = pi625 & n17404;
  assign n17406 = n3267 & n17399;
  assign n17407 = ~pi140 & ~n17406;
  assign n17408 = ~pi625 & n17407;
  assign n17409 = pi1153 & ~n17408;
  assign n17410 = ~n17405 & n17409;
  assign n17411 = ~pi608 & ~n17410;
  assign n17412 = ~n17296 & n17411;
  assign n17413 = pi625 & n17290;
  assign n17414 = ~pi625 & n17293;
  assign n17415 = pi1153 & ~n17414;
  assign n17416 = ~n17413 & n17415;
  assign n17417 = ~pi625 & n17404;
  assign n17418 = pi625 & n17407;
  assign n17419 = ~pi1153 & ~n17418;
  assign n17420 = ~n17417 & n17419;
  assign n17421 = pi608 & ~n17420;
  assign n17422 = ~n17416 & n17421;
  assign n17423 = ~n17412 & ~n17422;
  assign n17424 = pi778 & ~n17423;
  assign n17425 = ~pi778 & n17290;
  assign n17426 = ~n17424 & ~n17425;
  assign n17427 = ~pi609 & ~n17426;
  assign n17428 = ~pi778 & ~n17404;
  assign n17429 = ~n17410 & ~n17420;
  assign n17430 = pi778 & ~n17429;
  assign n17431 = ~n17428 & ~n17430;
  assign n17432 = pi609 & n17431;
  assign n17433 = ~pi1155 & ~n17432;
  assign n17434 = ~n17427 & n17433;
  assign n17435 = ~pi608 & pi1153;
  assign n17436 = pi608 & ~pi1153;
  assign n17437 = ~n17435 & ~n17436;
  assign n17438 = pi778 & ~n17437;
  assign n17439 = pi609 & ~n17438;
  assign n17440 = ~n17407 & ~n17439;
  assign n17441 = ~n17293 & ~n17438;
  assign n17442 = pi609 & n17441;
  assign n17443 = ~n17440 & ~n17442;
  assign n17444 = pi1155 & ~n17443;
  assign n17445 = ~pi660 & ~n17444;
  assign n17446 = ~n17434 & n17445;
  assign n17447 = pi609 & ~n17426;
  assign n17448 = ~pi609 & n17431;
  assign n17449 = pi1155 & ~n17448;
  assign n17450 = ~n17447 & n17449;
  assign n17451 = ~pi609 & ~n17438;
  assign n17452 = ~n17407 & ~n17451;
  assign n17453 = ~pi609 & n17441;
  assign n17454 = ~n17452 & ~n17453;
  assign n17455 = ~pi1155 & ~n17454;
  assign n17456 = pi660 & ~n17455;
  assign n17457 = ~n17450 & n17456;
  assign n17458 = ~n17446 & ~n17457;
  assign n17459 = pi785 & ~n17458;
  assign n17460 = ~pi785 & ~n17426;
  assign n17461 = ~n17459 & ~n17460;
  assign n17462 = ~pi618 & ~n17461;
  assign n17463 = ~pi660 & ~pi1155;
  assign n17464 = pi660 & pi1155;
  assign n17465 = pi785 & ~n17464;
  assign n17466 = ~n17463 & n17465;
  assign n17467 = ~n17431 & ~n17466;
  assign n17468 = ~n17407 & n17466;
  assign n17469 = ~n17467 & ~n17468;
  assign n17470 = pi618 & n17469;
  assign n17471 = ~pi1154 & ~n17470;
  assign n17472 = ~n17462 & n17471;
  assign n17473 = ~n17407 & n17438;
  assign n17474 = ~n17441 & ~n17473;
  assign n17475 = ~pi785 & ~n17474;
  assign n17476 = ~n17444 & ~n17455;
  assign n17477 = pi785 & ~n17476;
  assign n17478 = ~n17475 & ~n17477;
  assign n17479 = pi618 & n17478;
  assign n17480 = ~pi618 & n17407;
  assign n17481 = pi1154 & ~n17480;
  assign n17482 = ~n17479 & n17481;
  assign n17483 = ~pi627 & ~n17482;
  assign n17484 = ~n17472 & n17483;
  assign n17485 = pi618 & ~n17461;
  assign n17486 = ~pi618 & n17469;
  assign n17487 = pi1154 & ~n17486;
  assign n17488 = ~n17485 & n17487;
  assign n17489 = ~pi618 & n17478;
  assign n17490 = pi618 & n17407;
  assign n17491 = ~pi1154 & ~n17490;
  assign n17492 = ~n17489 & n17491;
  assign n17493 = pi627 & ~n17492;
  assign n17494 = ~n17488 & n17493;
  assign n17495 = ~n17484 & ~n17494;
  assign n17496 = pi781 & ~n17495;
  assign n17497 = ~pi781 & ~n17461;
  assign n17498 = ~n17496 & ~n17497;
  assign n17499 = ~pi619 & ~n17498;
  assign n17500 = ~pi627 & ~pi1154;
  assign n17501 = pi627 & pi1154;
  assign n17502 = pi781 & ~n17501;
  assign n17503 = ~n17500 & n17502;
  assign n17504 = n17469 & ~n17503;
  assign n17505 = n17407 & n17503;
  assign n17506 = ~n17504 & ~n17505;
  assign n17507 = pi619 & ~n17506;
  assign n17508 = ~pi1159 & ~n17507;
  assign n17509 = ~n17499 & n17508;
  assign n17510 = ~pi781 & ~n17478;
  assign n17511 = ~n17482 & ~n17492;
  assign n17512 = pi781 & ~n17511;
  assign n17513 = ~n17510 & ~n17512;
  assign n17514 = pi619 & n17513;
  assign n17515 = ~pi619 & n17407;
  assign n17516 = pi1159 & ~n17515;
  assign n17517 = ~n17514 & n17516;
  assign n17518 = ~pi648 & ~n17517;
  assign n17519 = ~n17509 & n17518;
  assign n17520 = pi619 & ~n17498;
  assign n17521 = ~pi619 & ~n17506;
  assign n17522 = pi1159 & ~n17521;
  assign n17523 = ~n17520 & n17522;
  assign n17524 = ~pi619 & n17513;
  assign n17525 = pi619 & n17407;
  assign n17526 = ~pi1159 & ~n17525;
  assign n17527 = ~n17524 & n17526;
  assign n17528 = pi648 & ~n17527;
  assign n17529 = ~n17523 & n17528;
  assign n17530 = ~n17519 & ~n17529;
  assign n17531 = pi789 & ~n17530;
  assign n17532 = ~pi789 & ~n17498;
  assign n17533 = ~n17531 & ~n17532;
  assign n17534 = ~pi788 & n17533;
  assign n17535 = ~pi626 & n17533;
  assign n17536 = ~pi648 & pi1159;
  assign n17537 = pi648 & ~pi1159;
  assign n17538 = ~n17536 & ~n17537;
  assign n17539 = pi789 & ~n17538;
  assign n17540 = n17506 & ~n17539;
  assign n17541 = ~n17407 & n17539;
  assign n17542 = ~n17540 & ~n17541;
  assign n17543 = pi626 & ~n17542;
  assign n17544 = ~pi641 & ~n17543;
  assign n17545 = ~n17535 & n17544;
  assign n17546 = ~pi641 & ~pi1158;
  assign n17547 = ~pi789 & ~n17513;
  assign n17548 = ~n17517 & ~n17527;
  assign n17549 = pi789 & ~n17548;
  assign n17550 = ~n17547 & ~n17549;
  assign n17551 = ~pi626 & n17550;
  assign n17552 = pi626 & n17407;
  assign n17553 = ~pi1158 & ~n17552;
  assign n17554 = ~n17551 & n17553;
  assign n17555 = ~n17546 & ~n17554;
  assign n17556 = ~n17545 & ~n17555;
  assign n17557 = pi626 & n17533;
  assign n17558 = ~pi626 & ~n17542;
  assign n17559 = pi641 & ~n17558;
  assign n17560 = ~n17557 & n17559;
  assign n17561 = pi641 & pi1158;
  assign n17562 = pi626 & n17550;
  assign n17563 = ~pi626 & n17407;
  assign n17564 = pi1158 & ~n17563;
  assign n17565 = ~n17562 & n17564;
  assign n17566 = ~n17561 & ~n17565;
  assign n17567 = ~n17560 & ~n17566;
  assign n17568 = ~n17556 & ~n17567;
  assign n17569 = pi788 & ~n17568;
  assign n17570 = ~n17534 & ~n17569;
  assign n17571 = ~pi628 & n17570;
  assign n17572 = ~n17554 & ~n17565;
  assign n17573 = pi788 & ~n17572;
  assign n17574 = ~pi788 & ~n17550;
  assign n17575 = ~n17573 & ~n17574;
  assign n17576 = pi628 & n17575;
  assign n17577 = ~pi1156 & ~n17576;
  assign n17578 = ~n17571 & n17577;
  assign n17579 = ~pi641 & pi1158;
  assign n17580 = pi641 & ~pi1158;
  assign n17581 = ~n17579 & ~n17580;
  assign n17582 = pi788 & ~n17581;
  assign n17583 = n17542 & ~n17582;
  assign n17584 = n17407 & n17582;
  assign n17585 = ~n17583 & ~n17584;
  assign n17586 = pi628 & ~n17585;
  assign n17587 = ~pi628 & n17407;
  assign n17588 = pi1156 & ~n17587;
  assign n17589 = ~n17586 & n17588;
  assign n17590 = ~pi629 & ~n17589;
  assign n17591 = ~n17578 & n17590;
  assign n17592 = pi628 & n17570;
  assign n17593 = ~pi628 & n17575;
  assign n17594 = pi1156 & ~n17593;
  assign n17595 = ~n17592 & n17594;
  assign n17596 = ~pi628 & ~n17585;
  assign n17597 = pi628 & n17407;
  assign n17598 = ~pi1156 & ~n17597;
  assign n17599 = ~n17596 & n17598;
  assign n17600 = pi629 & ~n17599;
  assign n17601 = ~n17595 & n17600;
  assign n17602 = ~n17591 & ~n17601;
  assign n17603 = pi792 & ~n17602;
  assign n17604 = ~pi792 & n17570;
  assign n17605 = ~n17603 & ~n17604;
  assign n17606 = ~pi647 & ~n17605;
  assign n17607 = ~pi629 & pi1156;
  assign n17608 = pi629 & ~pi1156;
  assign n17609 = ~n17607 & ~n17608;
  assign n17610 = pi792 & ~n17609;
  assign n17611 = n17575 & ~n17610;
  assign n17612 = n17407 & n17610;
  assign n17613 = ~n17611 & ~n17612;
  assign n17614 = pi647 & ~n17613;
  assign n17615 = ~pi1157 & ~n17614;
  assign n17616 = ~n17606 & n17615;
  assign n17617 = ~pi792 & n17585;
  assign n17618 = ~n17589 & ~n17599;
  assign n17619 = pi792 & ~n17618;
  assign n17620 = ~n17617 & ~n17619;
  assign n17621 = pi647 & n17620;
  assign n17622 = ~pi647 & n17407;
  assign n17623 = pi1157 & ~n17622;
  assign n17624 = ~n17621 & n17623;
  assign n17625 = ~pi630 & ~n17624;
  assign n17626 = ~n17616 & n17625;
  assign n17627 = pi647 & ~n17605;
  assign n17628 = ~pi647 & ~n17613;
  assign n17629 = pi1157 & ~n17628;
  assign n17630 = ~n17627 & n17629;
  assign n17631 = ~pi647 & n17620;
  assign n17632 = pi647 & n17407;
  assign n17633 = ~pi1157 & ~n17632;
  assign n17634 = ~n17631 & n17633;
  assign n17635 = pi630 & ~n17634;
  assign n17636 = ~n17630 & n17635;
  assign n17637 = ~n17626 & ~n17636;
  assign n17638 = pi787 & ~n17637;
  assign n17639 = ~pi787 & ~n17605;
  assign n17640 = ~n17638 & ~n17639;
  assign n17641 = ~pi644 & ~n17640;
  assign n17642 = ~pi787 & ~n17620;
  assign n17643 = ~n17624 & ~n17634;
  assign n17644 = pi787 & ~n17643;
  assign n17645 = ~n17642 & ~n17644;
  assign n17646 = pi644 & n17645;
  assign n17647 = ~pi715 & ~n17646;
  assign n17648 = ~n17641 & n17647;
  assign n17649 = ~pi630 & pi1157;
  assign n17650 = pi630 & ~pi1157;
  assign n17651 = ~n17649 & ~n17650;
  assign n17652 = pi787 & ~n17651;
  assign n17653 = n17613 & ~n17652;
  assign n17654 = ~n17407 & n17652;
  assign n17655 = ~n17653 & ~n17654;
  assign n17656 = ~pi644 & n17655;
  assign n17657 = pi644 & n17407;
  assign n17658 = pi715 & ~n17657;
  assign n17659 = ~n17656 & n17658;
  assign n17660 = ~pi1160 & ~n17659;
  assign n17661 = ~n17648 & n17660;
  assign n17662 = pi644 & ~n17640;
  assign n17663 = ~pi644 & n17645;
  assign n17664 = pi715 & ~n17663;
  assign n17665 = ~n17662 & n17664;
  assign n17666 = pi644 & n17655;
  assign n17667 = ~pi644 & n17407;
  assign n17668 = ~pi715 & ~n17667;
  assign n17669 = ~n17666 & n17668;
  assign n17670 = pi1160 & ~n17669;
  assign n17671 = ~n17665 & n17670;
  assign n17672 = pi790 & ~n17671;
  assign n17673 = ~n17661 & n17672;
  assign n17674 = ~pi790 & n17640;
  assign n17675 = ~po1038 & ~n17674;
  assign n17676 = ~n17673 & n17675;
  assign n17677 = ~pi140 & po1038;
  assign n17678 = ~pi832 & ~n17677;
  assign n17679 = ~n17676 & n17678;
  assign n17680 = ~pi140 & ~n2754;
  assign n17681 = ~pi738 & n16786;
  assign n17682 = ~n17680 & ~n17681;
  assign n17683 = ~pi778 & n17682;
  assign n17684 = ~pi625 & n17681;
  assign n17685 = ~n17682 & ~n17684;
  assign n17686 = pi1153 & ~n17685;
  assign n17687 = ~pi1153 & ~n17680;
  assign n17688 = ~n17684 & n17687;
  assign n17689 = ~n17686 & ~n17688;
  assign n17690 = pi778 & ~n17689;
  assign n17691 = ~n17683 & ~n17690;
  assign n17692 = n2754 & n17466;
  assign n17693 = n17691 & ~n17692;
  assign n17694 = n2754 & n17503;
  assign n17695 = n17693 & ~n17694;
  assign n17696 = n2754 & n17539;
  assign n17697 = n17695 & ~n17696;
  assign n17698 = ~pi626 & pi1158;
  assign n17699 = pi626 & ~pi1158;
  assign n17700 = ~n17698 & ~n17699;
  assign n17701 = ~pi626 & pi641;
  assign n17702 = pi626 & ~pi641;
  assign n17703 = ~n17701 & ~n17702;
  assign n17704 = ~n17700 & ~n17703;
  assign n17705 = n17697 & n17704;
  assign n17706 = n2754 & n17438;
  assign n17707 = ~pi761 & n16784;
  assign n17708 = ~n17680 & ~n17707;
  assign n17709 = ~n17706 & ~n17708;
  assign n17710 = ~pi785 & ~n17709;
  assign n17711 = n2754 & ~n17439;
  assign n17712 = ~n17708 & ~n17711;
  assign n17713 = pi1155 & ~n17712;
  assign n17714 = pi609 & n2754;
  assign n17715 = n17709 & ~n17714;
  assign n17716 = ~pi1155 & ~n17715;
  assign n17717 = ~n17713 & ~n17716;
  assign n17718 = pi785 & ~n17717;
  assign n17719 = ~n17710 & ~n17718;
  assign n17720 = ~pi781 & ~n17719;
  assign n17721 = ~pi618 & n2754;
  assign n17722 = n17719 & ~n17721;
  assign n17723 = pi1154 & ~n17722;
  assign n17724 = pi618 & n2754;
  assign n17725 = n17719 & ~n17724;
  assign n17726 = ~pi1154 & ~n17725;
  assign n17727 = ~n17723 & ~n17726;
  assign n17728 = pi781 & ~n17727;
  assign n17729 = ~n17720 & ~n17728;
  assign n17730 = ~pi789 & ~n17729;
  assign n17731 = pi619 & n17729;
  assign n17732 = ~pi619 & n17680;
  assign n17733 = pi1159 & ~n17732;
  assign n17734 = ~n17731 & n17733;
  assign n17735 = ~pi619 & n17729;
  assign n17736 = pi619 & n17680;
  assign n17737 = ~pi1159 & ~n17736;
  assign n17738 = ~n17735 & n17737;
  assign n17739 = ~n17734 & ~n17738;
  assign n17740 = pi789 & ~n17739;
  assign n17741 = ~n17730 & ~n17740;
  assign n17742 = pi626 & n17741;
  assign n17743 = ~pi626 & n17680;
  assign n17744 = pi1158 & ~n17743;
  assign n17745 = ~n17742 & n17744;
  assign n17746 = ~pi626 & n17741;
  assign n17747 = pi626 & n17680;
  assign n17748 = ~pi1158 & ~n17747;
  assign n17749 = ~n17746 & n17748;
  assign n17750 = ~n17745 & ~n17749;
  assign n17751 = ~n17581 & n17750;
  assign n17752 = ~n17705 & ~n17751;
  assign n17753 = pi788 & ~n17752;
  assign n17754 = ~n16521 & ~n17682;
  assign n17755 = pi625 & n17754;
  assign n17756 = n17708 & ~n17754;
  assign n17757 = ~n17755 & ~n17756;
  assign n17758 = n17687 & ~n17757;
  assign n17759 = ~pi608 & ~n17686;
  assign n17760 = ~n17758 & n17759;
  assign n17761 = pi1153 & n17708;
  assign n17762 = ~n17755 & n17761;
  assign n17763 = pi608 & ~n17688;
  assign n17764 = ~n17762 & n17763;
  assign n17765 = ~n17760 & ~n17764;
  assign n17766 = pi778 & ~n17765;
  assign n17767 = ~pi778 & ~n17756;
  assign n17768 = ~n17766 & ~n17767;
  assign n17769 = ~pi609 & ~n17768;
  assign n17770 = pi609 & n17691;
  assign n17771 = ~pi1155 & ~n17770;
  assign n17772 = ~n17769 & n17771;
  assign n17773 = ~pi660 & ~n17713;
  assign n17774 = ~n17772 & n17773;
  assign n17775 = pi609 & ~n17768;
  assign n17776 = ~pi609 & n17691;
  assign n17777 = pi1155 & ~n17776;
  assign n17778 = ~n17775 & n17777;
  assign n17779 = pi660 & ~n17716;
  assign n17780 = ~n17778 & n17779;
  assign n17781 = ~n17774 & ~n17780;
  assign n17782 = pi785 & ~n17781;
  assign n17783 = ~pi785 & ~n17768;
  assign n17784 = ~n17782 & ~n17783;
  assign n17785 = ~pi618 & ~n17784;
  assign n17786 = pi618 & n17693;
  assign n17787 = ~pi1154 & ~n17786;
  assign n17788 = ~n17785 & n17787;
  assign n17789 = ~pi627 & ~n17723;
  assign n17790 = ~n17788 & n17789;
  assign n17791 = pi618 & ~n17784;
  assign n17792 = ~pi618 & n17693;
  assign n17793 = pi1154 & ~n17792;
  assign n17794 = ~n17791 & n17793;
  assign n17795 = pi627 & ~n17726;
  assign n17796 = ~n17794 & n17795;
  assign n17797 = ~n17790 & ~n17796;
  assign n17798 = pi781 & ~n17797;
  assign n17799 = ~pi781 & ~n17784;
  assign n17800 = ~n17798 & ~n17799;
  assign n17801 = pi619 & ~n17800;
  assign n17802 = ~pi619 & n17695;
  assign n17803 = pi1159 & ~n17802;
  assign n17804 = ~n17801 & n17803;
  assign n17805 = pi648 & ~n17738;
  assign n17806 = ~n17804 & n17805;
  assign n17807 = ~pi619 & ~n17800;
  assign n17808 = pi619 & n17695;
  assign n17809 = ~pi1159 & ~n17808;
  assign n17810 = ~n17807 & n17809;
  assign n17811 = ~pi648 & ~n17734;
  assign n17812 = ~n17810 & n17811;
  assign n17813 = pi789 & ~n17812;
  assign n17814 = ~n17806 & n17813;
  assign n17815 = ~pi789 & n17800;
  assign n17816 = pi788 & ~n17700;
  assign n17817 = ~n17582 & ~n17816;
  assign n17818 = ~n17815 & n17817;
  assign n17819 = ~n17814 & n17818;
  assign n17820 = ~n17753 & ~n17819;
  assign n17821 = ~pi628 & ~n17820;
  assign n17822 = ~pi788 & ~n17741;
  assign n17823 = pi788 & ~n17750;
  assign n17824 = ~n17822 & ~n17823;
  assign n17825 = pi628 & n17824;
  assign n17826 = ~pi1156 & ~n17825;
  assign n17827 = ~n17821 & n17826;
  assign n17828 = n2754 & n17582;
  assign n17829 = n17697 & ~n17828;
  assign n17830 = ~pi628 & n2754;
  assign n17831 = n17829 & ~n17830;
  assign n17832 = pi1156 & ~n17831;
  assign n17833 = ~pi629 & ~n17832;
  assign n17834 = ~n17827 & n17833;
  assign n17835 = pi628 & ~n17820;
  assign n17836 = ~pi628 & n17824;
  assign n17837 = pi1156 & ~n17836;
  assign n17838 = ~n17835 & n17837;
  assign n17839 = pi628 & n2754;
  assign n17840 = n17829 & ~n17839;
  assign n17841 = ~pi1156 & ~n17840;
  assign n17842 = pi629 & ~n17841;
  assign n17843 = ~n17838 & n17842;
  assign n17844 = ~n17834 & ~n17843;
  assign n17845 = pi792 & ~n17844;
  assign n17846 = ~pi792 & ~n17820;
  assign n17847 = ~n17845 & ~n17846;
  assign n17848 = ~pi647 & ~n17847;
  assign n17849 = ~n17610 & n17824;
  assign n17850 = n17610 & n17680;
  assign n17851 = ~n17849 & ~n17850;
  assign n17852 = pi647 & ~n17851;
  assign n17853 = ~pi1157 & ~n17852;
  assign n17854 = ~n17848 & n17853;
  assign n17855 = ~pi628 & pi1156;
  assign n17856 = pi628 & ~pi1156;
  assign n17857 = ~n17855 & ~n17856;
  assign n17858 = pi792 & ~n17857;
  assign n17859 = n2754 & n17858;
  assign n17860 = n17829 & ~n17859;
  assign n17861 = pi647 & n17860;
  assign n17862 = ~pi647 & n17680;
  assign n17863 = pi1157 & ~n17862;
  assign n17864 = ~n17861 & n17863;
  assign n17865 = ~pi630 & ~n17864;
  assign n17866 = ~n17854 & n17865;
  assign n17867 = pi647 & ~n17847;
  assign n17868 = ~pi647 & ~n17851;
  assign n17869 = pi1157 & ~n17868;
  assign n17870 = ~n17867 & n17869;
  assign n17871 = ~pi647 & n17860;
  assign n17872 = pi647 & n17680;
  assign n17873 = ~pi1157 & ~n17872;
  assign n17874 = ~n17871 & n17873;
  assign n17875 = pi630 & ~n17874;
  assign n17876 = ~n17870 & n17875;
  assign n17877 = ~n17866 & ~n17876;
  assign n17878 = pi787 & ~n17877;
  assign n17879 = ~pi787 & ~n17847;
  assign n17880 = ~n17878 & ~n17879;
  assign n17881 = pi644 & ~n17880;
  assign n17882 = ~pi787 & ~n17860;
  assign n17883 = ~n17864 & ~n17874;
  assign n17884 = pi787 & ~n17883;
  assign n17885 = ~n17882 & ~n17884;
  assign n17886 = ~pi644 & n17885;
  assign n17887 = pi715 & ~n17886;
  assign n17888 = ~n17881 & n17887;
  assign n17889 = n17652 & ~n17680;
  assign n17890 = ~n17652 & n17851;
  assign n17891 = ~n17889 & ~n17890;
  assign n17892 = pi644 & n17891;
  assign n17893 = ~pi644 & n17680;
  assign n17894 = ~pi715 & ~n17893;
  assign n17895 = ~n17892 & n17894;
  assign n17896 = pi1160 & ~n17895;
  assign n17897 = ~n17888 & n17896;
  assign n17898 = ~pi644 & ~n17880;
  assign n17899 = pi644 & n17885;
  assign n17900 = ~pi715 & ~n17899;
  assign n17901 = ~n17898 & n17900;
  assign n17902 = ~pi644 & n17891;
  assign n17903 = pi644 & n17680;
  assign n17904 = pi715 & ~n17903;
  assign n17905 = ~n17902 & n17904;
  assign n17906 = ~pi1160 & ~n17905;
  assign n17907 = ~n17901 & n17906;
  assign n17908 = ~n17897 & ~n17907;
  assign n17909 = pi790 & ~n17908;
  assign n17910 = ~pi790 & ~n17880;
  assign n17911 = pi832 & ~n17910;
  assign n17912 = ~n17909 & n17911;
  assign po297 = ~n17679 & ~n17912;
  assign n17914 = pi141 & ~n3267;
  assign n17915 = ~pi141 & n16687;
  assign n17916 = pi141 & n16799;
  assign n17917 = ~pi749 & ~n17916;
  assign n17918 = ~n17915 & n17917;
  assign n17919 = pi141 & n16879;
  assign n17920 = ~pi141 & ~n16944;
  assign n17921 = pi749 & ~n17920;
  assign n17922 = ~n17919 & n17921;
  assign n17923 = pi39 & ~n17922;
  assign n17924 = ~n17918 & n17923;
  assign n17925 = pi141 & n17059;
  assign n17926 = ~pi141 & n17088;
  assign n17927 = ~pi749 & ~n17926;
  assign n17928 = ~n17925 & n17927;
  assign n17929 = ~pi141 & ~n17092;
  assign n17930 = pi141 & ~n17094;
  assign n17931 = pi749 & ~n17930;
  assign n17932 = ~n17929 & n17931;
  assign n17933 = ~pi39 & ~n17932;
  assign n17934 = ~n17928 & n17933;
  assign n17935 = ~pi38 & ~n17934;
  assign n17936 = ~n17924 & n17935;
  assign n17937 = ~pi141 & ~n17280;
  assign n17938 = pi749 & n17282;
  assign n17939 = ~n17937 & ~n17938;
  assign n17940 = ~pi39 & n17107;
  assign n17941 = pi38 & ~n17940;
  assign n17942 = n17939 & n17941;
  assign n17943 = pi706 & ~n17942;
  assign n17944 = ~n17936 & n17943;
  assign n17945 = pi38 & ~n17939;
  assign n17946 = ~pi749 & n17199;
  assign n17947 = pi141 & n17273;
  assign n17948 = ~n17946 & ~n17947;
  assign n17949 = pi39 & ~n17948;
  assign n17950 = ~pi141 & n17242;
  assign n17951 = pi141 & n17246;
  assign n17952 = pi749 & ~n17951;
  assign n17953 = ~n17950 & n17952;
  assign n17954 = ~pi39 & n17120;
  assign n17955 = ~pi141 & ~pi749;
  assign n17956 = ~n17954 & n17955;
  assign n17957 = ~n17953 & ~n17956;
  assign n17958 = ~pi38 & ~n17957;
  assign n17959 = ~n17949 & n17958;
  assign n17960 = ~n17945 & ~n17959;
  assign n17961 = ~pi706 & ~n17960;
  assign n17962 = n3267 & ~n17961;
  assign n17963 = ~n17944 & n17962;
  assign n17964 = ~n17914 & ~n17963;
  assign n17965 = ~pi625 & n17964;
  assign n17966 = n3267 & n17960;
  assign n17967 = ~n17914 & ~n17966;
  assign n17968 = pi625 & n17967;
  assign n17969 = ~pi1153 & ~n17968;
  assign n17970 = ~n17965 & n17969;
  assign n17971 = ~pi39 & n17078;
  assign n17972 = ~n17382 & ~n17971;
  assign n17973 = ~pi141 & n17972;
  assign n17974 = pi39 & ~n17332;
  assign n17975 = ~pi39 & n17057;
  assign n17976 = ~n17974 & ~n17975;
  assign n17977 = pi141 & ~n17976;
  assign n17978 = ~pi38 & ~n17977;
  assign n17979 = ~n17973 & n17978;
  assign n17980 = n17392 & ~n17937;
  assign n17981 = pi706 & ~n17980;
  assign n17982 = ~n17979 & n17981;
  assign n17983 = ~pi141 & ~pi706;
  assign n17984 = ~n17399 & n17983;
  assign n17985 = n3267 & ~n17984;
  assign n17986 = ~n17982 & n17985;
  assign n17987 = ~n17914 & ~n17986;
  assign n17988 = pi625 & n17987;
  assign n17989 = ~pi141 & ~n17406;
  assign n17990 = ~pi625 & n17989;
  assign n17991 = pi1153 & ~n17990;
  assign n17992 = ~n17988 & n17991;
  assign n17993 = ~pi608 & ~n17992;
  assign n17994 = ~n17970 & n17993;
  assign n17995 = pi625 & n17964;
  assign n17996 = ~pi625 & n17967;
  assign n17997 = pi1153 & ~n17996;
  assign n17998 = ~n17995 & n17997;
  assign n17999 = ~pi625 & n17987;
  assign n18000 = pi625 & n17989;
  assign n18001 = ~pi1153 & ~n18000;
  assign n18002 = ~n17999 & n18001;
  assign n18003 = pi608 & ~n18002;
  assign n18004 = ~n17998 & n18003;
  assign n18005 = ~n17994 & ~n18004;
  assign n18006 = pi778 & ~n18005;
  assign n18007 = ~pi778 & n17964;
  assign n18008 = ~n18006 & ~n18007;
  assign n18009 = ~pi609 & ~n18008;
  assign n18010 = ~pi778 & ~n17987;
  assign n18011 = ~n17992 & ~n18002;
  assign n18012 = pi778 & ~n18011;
  assign n18013 = ~n18010 & ~n18012;
  assign n18014 = pi609 & n18013;
  assign n18015 = ~pi1155 & ~n18014;
  assign n18016 = ~n18009 & n18015;
  assign n18017 = ~n17439 & ~n17989;
  assign n18018 = ~n17438 & ~n17967;
  assign n18019 = pi609 & n18018;
  assign n18020 = ~n18017 & ~n18019;
  assign n18021 = pi1155 & ~n18020;
  assign n18022 = ~pi660 & ~n18021;
  assign n18023 = ~n18016 & n18022;
  assign n18024 = pi609 & ~n18008;
  assign n18025 = ~pi609 & n18013;
  assign n18026 = pi1155 & ~n18025;
  assign n18027 = ~n18024 & n18026;
  assign n18028 = ~n17451 & ~n17989;
  assign n18029 = ~pi609 & n18018;
  assign n18030 = ~n18028 & ~n18029;
  assign n18031 = ~pi1155 & ~n18030;
  assign n18032 = pi660 & ~n18031;
  assign n18033 = ~n18027 & n18032;
  assign n18034 = ~n18023 & ~n18033;
  assign n18035 = pi785 & ~n18034;
  assign n18036 = ~pi785 & ~n18008;
  assign n18037 = ~n18035 & ~n18036;
  assign n18038 = ~pi618 & ~n18037;
  assign n18039 = ~n17466 & ~n18013;
  assign n18040 = n17466 & ~n17989;
  assign n18041 = ~n18039 & ~n18040;
  assign n18042 = pi618 & n18041;
  assign n18043 = ~pi1154 & ~n18042;
  assign n18044 = ~n18038 & n18043;
  assign n18045 = n17438 & ~n17989;
  assign n18046 = ~n18018 & ~n18045;
  assign n18047 = ~pi785 & ~n18046;
  assign n18048 = ~n18021 & ~n18031;
  assign n18049 = pi785 & ~n18048;
  assign n18050 = ~n18047 & ~n18049;
  assign n18051 = pi618 & n18050;
  assign n18052 = ~pi618 & n17989;
  assign n18053 = pi1154 & ~n18052;
  assign n18054 = ~n18051 & n18053;
  assign n18055 = ~pi627 & ~n18054;
  assign n18056 = ~n18044 & n18055;
  assign n18057 = pi618 & ~n18037;
  assign n18058 = ~pi618 & n18041;
  assign n18059 = pi1154 & ~n18058;
  assign n18060 = ~n18057 & n18059;
  assign n18061 = ~pi618 & n18050;
  assign n18062 = pi618 & n17989;
  assign n18063 = ~pi1154 & ~n18062;
  assign n18064 = ~n18061 & n18063;
  assign n18065 = pi627 & ~n18064;
  assign n18066 = ~n18060 & n18065;
  assign n18067 = ~n18056 & ~n18066;
  assign n18068 = pi781 & ~n18067;
  assign n18069 = ~pi781 & ~n18037;
  assign n18070 = ~n18068 & ~n18069;
  assign n18071 = ~pi619 & ~n18070;
  assign n18072 = ~n17503 & n18041;
  assign n18073 = n17503 & n17989;
  assign n18074 = ~n18072 & ~n18073;
  assign n18075 = pi619 & ~n18074;
  assign n18076 = ~pi1159 & ~n18075;
  assign n18077 = ~n18071 & n18076;
  assign n18078 = ~pi781 & ~n18050;
  assign n18079 = ~n18054 & ~n18064;
  assign n18080 = pi781 & ~n18079;
  assign n18081 = ~n18078 & ~n18080;
  assign n18082 = pi619 & n18081;
  assign n18083 = ~pi619 & n17989;
  assign n18084 = pi1159 & ~n18083;
  assign n18085 = ~n18082 & n18084;
  assign n18086 = ~pi648 & ~n18085;
  assign n18087 = ~n18077 & n18086;
  assign n18088 = pi619 & ~n18070;
  assign n18089 = ~pi619 & ~n18074;
  assign n18090 = pi1159 & ~n18089;
  assign n18091 = ~n18088 & n18090;
  assign n18092 = ~pi619 & n18081;
  assign n18093 = pi619 & n17989;
  assign n18094 = ~pi1159 & ~n18093;
  assign n18095 = ~n18092 & n18094;
  assign n18096 = pi648 & ~n18095;
  assign n18097 = ~n18091 & n18096;
  assign n18098 = ~n18087 & ~n18097;
  assign n18099 = pi789 & ~n18098;
  assign n18100 = ~pi789 & ~n18070;
  assign n18101 = ~n18099 & ~n18100;
  assign n18102 = ~pi788 & n18101;
  assign n18103 = ~pi626 & n18101;
  assign n18104 = n17539 & ~n17989;
  assign n18105 = ~n17539 & n18074;
  assign n18106 = ~n18104 & ~n18105;
  assign n18107 = pi626 & ~n18106;
  assign n18108 = ~pi641 & ~n18107;
  assign n18109 = ~n18103 & n18108;
  assign n18110 = ~pi789 & ~n18081;
  assign n18111 = ~n18085 & ~n18095;
  assign n18112 = pi789 & ~n18111;
  assign n18113 = ~n18110 & ~n18112;
  assign n18114 = ~pi626 & n18113;
  assign n18115 = pi626 & n17989;
  assign n18116 = ~pi1158 & ~n18115;
  assign n18117 = ~n18114 & n18116;
  assign n18118 = ~n17546 & ~n18117;
  assign n18119 = ~n18109 & ~n18118;
  assign n18120 = pi626 & n18101;
  assign n18121 = ~pi626 & ~n18106;
  assign n18122 = pi641 & ~n18121;
  assign n18123 = ~n18120 & n18122;
  assign n18124 = pi626 & n18113;
  assign n18125 = ~pi626 & n17989;
  assign n18126 = pi1158 & ~n18125;
  assign n18127 = ~n18124 & n18126;
  assign n18128 = ~n17561 & ~n18127;
  assign n18129 = ~n18123 & ~n18128;
  assign n18130 = ~n18119 & ~n18129;
  assign n18131 = pi788 & ~n18130;
  assign n18132 = ~n18102 & ~n18131;
  assign n18133 = ~pi628 & n18132;
  assign n18134 = ~n18117 & ~n18127;
  assign n18135 = pi788 & ~n18134;
  assign n18136 = ~pi788 & ~n18113;
  assign n18137 = ~n18135 & ~n18136;
  assign n18138 = pi628 & n18137;
  assign n18139 = ~pi1156 & ~n18138;
  assign n18140 = ~n18133 & n18139;
  assign n18141 = ~n17582 & n18106;
  assign n18142 = n17582 & n17989;
  assign n18143 = ~n18141 & ~n18142;
  assign n18144 = pi628 & ~n18143;
  assign n18145 = ~pi628 & n17989;
  assign n18146 = pi1156 & ~n18145;
  assign n18147 = ~n18144 & n18146;
  assign n18148 = ~pi629 & ~n18147;
  assign n18149 = ~n18140 & n18148;
  assign n18150 = pi628 & n18132;
  assign n18151 = ~pi628 & n18137;
  assign n18152 = pi1156 & ~n18151;
  assign n18153 = ~n18150 & n18152;
  assign n18154 = ~pi628 & ~n18143;
  assign n18155 = pi628 & n17989;
  assign n18156 = ~pi1156 & ~n18155;
  assign n18157 = ~n18154 & n18156;
  assign n18158 = pi629 & ~n18157;
  assign n18159 = ~n18153 & n18158;
  assign n18160 = ~n18149 & ~n18159;
  assign n18161 = pi792 & ~n18160;
  assign n18162 = ~pi792 & n18132;
  assign n18163 = ~n18161 & ~n18162;
  assign n18164 = ~pi647 & ~n18163;
  assign n18165 = ~n17610 & n18137;
  assign n18166 = n17610 & n17989;
  assign n18167 = ~n18165 & ~n18166;
  assign n18168 = pi647 & ~n18167;
  assign n18169 = ~pi1157 & ~n18168;
  assign n18170 = ~n18164 & n18169;
  assign n18171 = ~pi792 & n18143;
  assign n18172 = ~n18147 & ~n18157;
  assign n18173 = pi792 & ~n18172;
  assign n18174 = ~n18171 & ~n18173;
  assign n18175 = pi647 & n18174;
  assign n18176 = ~pi647 & n17989;
  assign n18177 = pi1157 & ~n18176;
  assign n18178 = ~n18175 & n18177;
  assign n18179 = ~pi630 & ~n18178;
  assign n18180 = ~n18170 & n18179;
  assign n18181 = pi647 & ~n18163;
  assign n18182 = ~pi647 & ~n18167;
  assign n18183 = pi1157 & ~n18182;
  assign n18184 = ~n18181 & n18183;
  assign n18185 = ~pi647 & n18174;
  assign n18186 = pi647 & n17989;
  assign n18187 = ~pi1157 & ~n18186;
  assign n18188 = ~n18185 & n18187;
  assign n18189 = pi630 & ~n18188;
  assign n18190 = ~n18184 & n18189;
  assign n18191 = ~n18180 & ~n18190;
  assign n18192 = pi787 & ~n18191;
  assign n18193 = ~pi787 & ~n18163;
  assign n18194 = ~n18192 & ~n18193;
  assign n18195 = ~pi644 & ~n18194;
  assign n18196 = ~pi787 & ~n18174;
  assign n18197 = ~n18178 & ~n18188;
  assign n18198 = pi787 & ~n18197;
  assign n18199 = ~n18196 & ~n18198;
  assign n18200 = pi644 & n18199;
  assign n18201 = ~pi715 & ~n18200;
  assign n18202 = ~n18195 & n18201;
  assign n18203 = n17652 & ~n17989;
  assign n18204 = ~n17652 & n18167;
  assign n18205 = ~n18203 & ~n18204;
  assign n18206 = ~pi644 & n18205;
  assign n18207 = pi644 & n17989;
  assign n18208 = pi715 & ~n18207;
  assign n18209 = ~n18206 & n18208;
  assign n18210 = ~pi1160 & ~n18209;
  assign n18211 = ~n18202 & n18210;
  assign n18212 = pi644 & ~n18194;
  assign n18213 = ~pi644 & n18199;
  assign n18214 = pi715 & ~n18213;
  assign n18215 = ~n18212 & n18214;
  assign n18216 = pi644 & n18205;
  assign n18217 = ~pi644 & n17989;
  assign n18218 = ~pi715 & ~n18217;
  assign n18219 = ~n18216 & n18218;
  assign n18220 = pi1160 & ~n18219;
  assign n18221 = ~n18215 & n18220;
  assign n18222 = pi790 & ~n18221;
  assign n18223 = ~n18211 & n18222;
  assign n18224 = ~pi790 & n18194;
  assign n18225 = ~po1038 & ~n18224;
  assign n18226 = ~n18223 & n18225;
  assign n18227 = ~pi141 & po1038;
  assign n18228 = ~pi832 & ~n18227;
  assign n18229 = ~n18226 & n18228;
  assign n18230 = ~pi141 & ~n2754;
  assign n18231 = pi706 & n16786;
  assign n18232 = ~n18230 & ~n18231;
  assign n18233 = ~pi778 & n18232;
  assign n18234 = ~pi625 & n18231;
  assign n18235 = ~n18232 & ~n18234;
  assign n18236 = pi1153 & ~n18235;
  assign n18237 = ~pi1153 & ~n18230;
  assign n18238 = ~n18234 & n18237;
  assign n18239 = ~n18236 & ~n18238;
  assign n18240 = pi778 & ~n18239;
  assign n18241 = ~n18233 & ~n18240;
  assign n18242 = ~n17692 & n18241;
  assign n18243 = ~n17694 & n18242;
  assign n18244 = ~n17696 & n18243;
  assign n18245 = n17704 & n18244;
  assign n18246 = pi749 & n16784;
  assign n18247 = ~n18230 & ~n18246;
  assign n18248 = ~n17706 & ~n18247;
  assign n18249 = ~pi785 & ~n18248;
  assign n18250 = ~n17711 & ~n18247;
  assign n18251 = pi1155 & ~n18250;
  assign n18252 = ~n17714 & n18248;
  assign n18253 = ~pi1155 & ~n18252;
  assign n18254 = ~n18251 & ~n18253;
  assign n18255 = pi785 & ~n18254;
  assign n18256 = ~n18249 & ~n18255;
  assign n18257 = ~pi781 & ~n18256;
  assign n18258 = ~n17721 & n18256;
  assign n18259 = pi1154 & ~n18258;
  assign n18260 = ~n17724 & n18256;
  assign n18261 = ~pi1154 & ~n18260;
  assign n18262 = ~n18259 & ~n18261;
  assign n18263 = pi781 & ~n18262;
  assign n18264 = ~n18257 & ~n18263;
  assign n18265 = ~pi789 & ~n18264;
  assign n18266 = pi619 & n18264;
  assign n18267 = ~pi619 & n18230;
  assign n18268 = pi1159 & ~n18267;
  assign n18269 = ~n18266 & n18268;
  assign n18270 = ~pi619 & n18264;
  assign n18271 = pi619 & n18230;
  assign n18272 = ~pi1159 & ~n18271;
  assign n18273 = ~n18270 & n18272;
  assign n18274 = ~n18269 & ~n18273;
  assign n18275 = pi789 & ~n18274;
  assign n18276 = ~n18265 & ~n18275;
  assign n18277 = pi626 & n18276;
  assign n18278 = ~pi626 & n18230;
  assign n18279 = pi1158 & ~n18278;
  assign n18280 = ~n18277 & n18279;
  assign n18281 = ~pi626 & n18276;
  assign n18282 = pi626 & n18230;
  assign n18283 = ~pi1158 & ~n18282;
  assign n18284 = ~n18281 & n18283;
  assign n18285 = ~n18280 & ~n18284;
  assign n18286 = ~n17581 & n18285;
  assign n18287 = ~n18245 & ~n18286;
  assign n18288 = pi788 & ~n18287;
  assign n18289 = ~n16521 & ~n18232;
  assign n18290 = pi625 & n18289;
  assign n18291 = n18247 & ~n18289;
  assign n18292 = ~n18290 & ~n18291;
  assign n18293 = n18237 & ~n18292;
  assign n18294 = ~pi608 & ~n18236;
  assign n18295 = ~n18293 & n18294;
  assign n18296 = pi1153 & n18247;
  assign n18297 = ~n18290 & n18296;
  assign n18298 = pi608 & ~n18238;
  assign n18299 = ~n18297 & n18298;
  assign n18300 = ~n18295 & ~n18299;
  assign n18301 = pi778 & ~n18300;
  assign n18302 = ~pi778 & ~n18291;
  assign n18303 = ~n18301 & ~n18302;
  assign n18304 = ~pi609 & ~n18303;
  assign n18305 = pi609 & n18241;
  assign n18306 = ~pi1155 & ~n18305;
  assign n18307 = ~n18304 & n18306;
  assign n18308 = ~pi660 & ~n18251;
  assign n18309 = ~n18307 & n18308;
  assign n18310 = pi609 & ~n18303;
  assign n18311 = ~pi609 & n18241;
  assign n18312 = pi1155 & ~n18311;
  assign n18313 = ~n18310 & n18312;
  assign n18314 = pi660 & ~n18253;
  assign n18315 = ~n18313 & n18314;
  assign n18316 = ~n18309 & ~n18315;
  assign n18317 = pi785 & ~n18316;
  assign n18318 = ~pi785 & ~n18303;
  assign n18319 = ~n18317 & ~n18318;
  assign n18320 = ~pi618 & ~n18319;
  assign n18321 = pi618 & n18242;
  assign n18322 = ~pi1154 & ~n18321;
  assign n18323 = ~n18320 & n18322;
  assign n18324 = ~pi627 & ~n18259;
  assign n18325 = ~n18323 & n18324;
  assign n18326 = pi618 & ~n18319;
  assign n18327 = ~pi618 & n18242;
  assign n18328 = pi1154 & ~n18327;
  assign n18329 = ~n18326 & n18328;
  assign n18330 = pi627 & ~n18261;
  assign n18331 = ~n18329 & n18330;
  assign n18332 = ~n18325 & ~n18331;
  assign n18333 = pi781 & ~n18332;
  assign n18334 = ~pi781 & ~n18319;
  assign n18335 = ~n18333 & ~n18334;
  assign n18336 = pi619 & ~n18335;
  assign n18337 = ~pi619 & n18243;
  assign n18338 = pi1159 & ~n18337;
  assign n18339 = ~n18336 & n18338;
  assign n18340 = pi648 & ~n18273;
  assign n18341 = ~n18339 & n18340;
  assign n18342 = ~pi619 & ~n18335;
  assign n18343 = pi619 & n18243;
  assign n18344 = ~pi1159 & ~n18343;
  assign n18345 = ~n18342 & n18344;
  assign n18346 = ~pi648 & ~n18269;
  assign n18347 = ~n18345 & n18346;
  assign n18348 = pi789 & ~n18347;
  assign n18349 = ~n18341 & n18348;
  assign n18350 = ~pi789 & n18335;
  assign n18351 = n17817 & ~n18350;
  assign n18352 = ~n18349 & n18351;
  assign n18353 = ~n18288 & ~n18352;
  assign n18354 = ~pi628 & ~n18353;
  assign n18355 = ~pi788 & ~n18276;
  assign n18356 = pi788 & ~n18285;
  assign n18357 = ~n18355 & ~n18356;
  assign n18358 = pi628 & n18357;
  assign n18359 = ~pi1156 & ~n18358;
  assign n18360 = ~n18354 & n18359;
  assign n18361 = ~n17828 & n18244;
  assign n18362 = ~n17830 & n18361;
  assign n18363 = pi1156 & ~n18362;
  assign n18364 = ~pi629 & ~n18363;
  assign n18365 = ~n18360 & n18364;
  assign n18366 = pi628 & ~n18353;
  assign n18367 = ~pi628 & n18357;
  assign n18368 = pi1156 & ~n18367;
  assign n18369 = ~n18366 & n18368;
  assign n18370 = ~n17839 & n18361;
  assign n18371 = ~pi1156 & ~n18370;
  assign n18372 = pi629 & ~n18371;
  assign n18373 = ~n18369 & n18372;
  assign n18374 = ~n18365 & ~n18373;
  assign n18375 = pi792 & ~n18374;
  assign n18376 = ~pi792 & ~n18353;
  assign n18377 = ~n18375 & ~n18376;
  assign n18378 = ~pi647 & ~n18377;
  assign n18379 = ~n17610 & n18357;
  assign n18380 = n17610 & n18230;
  assign n18381 = ~n18379 & ~n18380;
  assign n18382 = pi647 & ~n18381;
  assign n18383 = ~pi1157 & ~n18382;
  assign n18384 = ~n18378 & n18383;
  assign n18385 = ~n17859 & n18361;
  assign n18386 = pi647 & n18385;
  assign n18387 = ~pi647 & n18230;
  assign n18388 = pi1157 & ~n18387;
  assign n18389 = ~n18386 & n18388;
  assign n18390 = ~pi630 & ~n18389;
  assign n18391 = ~n18384 & n18390;
  assign n18392 = pi647 & ~n18377;
  assign n18393 = ~pi647 & ~n18381;
  assign n18394 = pi1157 & ~n18393;
  assign n18395 = ~n18392 & n18394;
  assign n18396 = ~pi647 & n18385;
  assign n18397 = pi647 & n18230;
  assign n18398 = ~pi1157 & ~n18397;
  assign n18399 = ~n18396 & n18398;
  assign n18400 = pi630 & ~n18399;
  assign n18401 = ~n18395 & n18400;
  assign n18402 = ~n18391 & ~n18401;
  assign n18403 = pi787 & ~n18402;
  assign n18404 = ~pi787 & ~n18377;
  assign n18405 = ~n18403 & ~n18404;
  assign n18406 = pi644 & ~n18405;
  assign n18407 = ~pi787 & ~n18385;
  assign n18408 = ~n18389 & ~n18399;
  assign n18409 = pi787 & ~n18408;
  assign n18410 = ~n18407 & ~n18409;
  assign n18411 = ~pi644 & n18410;
  assign n18412 = pi715 & ~n18411;
  assign n18413 = ~n18406 & n18412;
  assign n18414 = n17652 & ~n18230;
  assign n18415 = ~n17652 & n18381;
  assign n18416 = ~n18414 & ~n18415;
  assign n18417 = pi644 & n18416;
  assign n18418 = ~pi644 & n18230;
  assign n18419 = ~pi715 & ~n18418;
  assign n18420 = ~n18417 & n18419;
  assign n18421 = pi1160 & ~n18420;
  assign n18422 = ~n18413 & n18421;
  assign n18423 = ~pi644 & ~n18405;
  assign n18424 = pi644 & n18410;
  assign n18425 = ~pi715 & ~n18424;
  assign n18426 = ~n18423 & n18425;
  assign n18427 = ~pi644 & n18416;
  assign n18428 = pi644 & n18230;
  assign n18429 = pi715 & ~n18428;
  assign n18430 = ~n18427 & n18429;
  assign n18431 = ~pi1160 & ~n18430;
  assign n18432 = ~n18426 & n18431;
  assign n18433 = ~n18422 & ~n18432;
  assign n18434 = pi790 & ~n18433;
  assign n18435 = ~pi790 & ~n18405;
  assign n18436 = pi832 & ~n18435;
  assign n18437 = ~n18434 & n18436;
  assign po298 = ~n18229 & ~n18437;
  assign n18439 = pi142 & ~n3267;
  assign n18440 = pi142 & ~n17040;
  assign n18441 = n17070 & n18440;
  assign n18442 = ~pi142 & ~n17079;
  assign n18443 = ~n17050 & n18442;
  assign n18444 = ~n18441 & ~n18443;
  assign n18445 = pi743 & ~n18444;
  assign n18446 = ~n16722 & n17049;
  assign n18447 = ~n17040 & n18446;
  assign n18448 = pi680 & n18447;
  assign n18449 = ~pi142 & n18448;
  assign n18450 = pi142 & ~n17070;
  assign n18451 = ~n17079 & n18450;
  assign n18452 = ~pi743 & ~n18451;
  assign n18453 = ~n18449 & n18452;
  assign n18454 = ~pi299 & ~n18453;
  assign n18455 = ~n18445 & n18454;
  assign n18456 = ~n16722 & n17054;
  assign n18457 = n17027 & n18456;
  assign n18458 = pi680 & n18457;
  assign n18459 = ~pi142 & n18458;
  assign n18460 = pi142 & ~n17076;
  assign n18461 = ~n17084 & n18460;
  assign n18462 = ~pi743 & ~n18461;
  assign n18463 = ~n18459 & n18462;
  assign n18464 = ~pi142 & ~n17084;
  assign n18465 = ~n17055 & n18464;
  assign n18466 = pi142 & n17027;
  assign n18467 = ~n17075 & n18466;
  assign n18468 = ~n18465 & ~n18467;
  assign n18469 = pi743 & ~n18468;
  assign n18470 = pi299 & ~n18469;
  assign n18471 = ~n18463 & n18470;
  assign n18472 = ~n18455 & ~n18471;
  assign n18473 = pi735 & ~n18472;
  assign n18474 = pi743 & ~n18442;
  assign n18475 = ~n18440 & n18474;
  assign n18476 = pi142 & ~pi743;
  assign n18477 = ~n17063 & n18476;
  assign n18478 = ~pi299 & ~n18477;
  assign n18479 = ~n18475 & n18478;
  assign n18480 = pi142 & ~n17026;
  assign n18481 = ~pi743 & ~n18480;
  assign n18482 = ~n18464 & ~n18481;
  assign n18483 = ~n18466 & n18482;
  assign n18484 = pi299 & ~n18483;
  assign n18485 = ~n18479 & ~n18484;
  assign n18486 = ~pi735 & n18485;
  assign n18487 = ~pi39 & ~n18486;
  assign n18488 = ~n18473 & n18487;
  assign n18489 = pi142 & n16919;
  assign n18490 = ~pi142 & n16860;
  assign n18491 = pi743 & ~n18490;
  assign n18492 = ~n18489 & n18491;
  assign n18493 = ~pi142 & ~n16759;
  assign n18494 = pi142 & n16597;
  assign n18495 = ~pi743 & ~n18494;
  assign n18496 = ~n18493 & n18495;
  assign n18497 = ~n18492 & ~n18496;
  assign n18498 = pi735 & ~n18497;
  assign n18499 = pi142 & ~n17132;
  assign n18500 = ~pi743 & ~n18499;
  assign n18501 = pi142 & ~n17221;
  assign n18502 = pi743 & n16856;
  assign n18503 = ~n18501 & n18502;
  assign n18504 = ~n18500 & ~n18503;
  assign n18505 = ~pi735 & n18504;
  assign n18506 = ~n18498 & ~n18505;
  assign n18507 = ~n6189 & n18506;
  assign n18508 = pi142 & ~n16925;
  assign n18509 = ~pi142 & ~n16854;
  assign n18510 = pi743 & ~n18509;
  assign n18511 = ~n18508 & n18510;
  assign n18512 = pi142 & n16580;
  assign n18513 = ~pi142 & n16771;
  assign n18514 = ~pi743 & ~n18513;
  assign n18515 = ~n18512 & n18514;
  assign n18516 = ~n18511 & ~n18515;
  assign n18517 = pi735 & ~n18516;
  assign n18518 = pi142 & ~n17151;
  assign n18519 = ~pi743 & ~n18518;
  assign n18520 = pi142 & n17216;
  assign n18521 = pi743 & n16850;
  assign n18522 = ~n18520 & n18521;
  assign n18523 = ~n18519 & ~n18522;
  assign n18524 = ~pi735 & n18523;
  assign n18525 = ~n18517 & ~n18524;
  assign n18526 = n6189 & n18525;
  assign n18527 = pi215 & ~n18526;
  assign n18528 = ~n18507 & n18527;
  assign n18529 = ~pi142 & ~n16835;
  assign n18530 = pi142 & n16900;
  assign n18531 = pi743 & ~n18530;
  assign n18532 = ~n18529 & n18531;
  assign n18533 = pi142 & n16646;
  assign n18534 = ~pi142 & n16732;
  assign n18535 = ~pi743 & ~n18534;
  assign n18536 = ~n18533 & n18535;
  assign n18537 = ~n18532 & ~n18536;
  assign n18538 = pi735 & ~n18537;
  assign n18539 = ~pi142 & n17250;
  assign n18540 = pi142 & n17207;
  assign n18541 = ~n18539 & ~n18540;
  assign n18542 = pi743 & ~n18541;
  assign n18543 = pi142 & ~n17172;
  assign n18544 = ~pi743 & ~n18543;
  assign n18545 = ~n18542 & ~n18544;
  assign n18546 = ~pi735 & n18545;
  assign n18547 = ~n18538 & ~n18546;
  assign n18548 = n6189 & ~n18547;
  assign n18549 = ~pi142 & ~n16816;
  assign n18550 = pi142 & n16889;
  assign n18551 = pi743 & ~n18550;
  assign n18552 = ~n18549 & n18551;
  assign n18553 = ~pi142 & ~n16711;
  assign n18554 = pi142 & n16663;
  assign n18555 = ~pi743 & ~n18554;
  assign n18556 = ~n18553 & n18555;
  assign n18557 = ~n18552 & ~n18556;
  assign n18558 = pi735 & ~n18557;
  assign n18559 = pi142 & ~n16812;
  assign n18560 = pi743 & n16813;
  assign n18561 = ~n18559 & ~n18560;
  assign n18562 = ~pi735 & ~n18561;
  assign n18563 = ~n18558 & ~n18562;
  assign n18564 = ~n6189 & ~n18563;
  assign n18565 = ~n3329 & ~n18564;
  assign n18566 = ~n18548 & n18565;
  assign n18567 = pi142 & ~n16518;
  assign n18568 = pi743 & n16543;
  assign n18569 = ~n18567 & ~n18568;
  assign n18570 = ~pi735 & n18569;
  assign n18571 = pi142 & ~n16529;
  assign n18572 = pi743 & n16784;
  assign n18573 = n3095 & n18572;
  assign n18574 = ~n18571 & ~n18573;
  assign n18575 = ~n17107 & n18574;
  assign n18576 = ~n16515 & ~n18575;
  assign n18577 = pi735 & ~n18576;
  assign n18578 = ~n18567 & n18577;
  assign n18579 = ~n18570 & ~n18578;
  assign n18580 = n3329 & ~n18579;
  assign n18581 = ~pi215 & ~n18580;
  assign n18582 = ~n18566 & n18581;
  assign n18583 = ~n18528 & ~n18582;
  assign n18584 = pi299 & ~n18583;
  assign n18585 = ~n6215 & n18506;
  assign n18586 = n6215 & n18525;
  assign n18587 = pi223 & ~n18586;
  assign n18588 = ~n18585 & n18587;
  assign n18589 = n6215 & ~n18547;
  assign n18590 = ~n6215 & ~n18563;
  assign n18591 = ~n3052 & ~n18590;
  assign n18592 = ~n18589 & n18591;
  assign n18593 = n3052 & ~n18579;
  assign n18594 = ~pi223 & ~n18593;
  assign n18595 = ~n18592 & n18594;
  assign n18596 = ~n18588 & ~n18595;
  assign n18597 = ~pi299 & ~n18596;
  assign n18598 = pi39 & ~n18597;
  assign n18599 = ~n18584 & n18598;
  assign n18600 = ~n18488 & ~n18599;
  assign n18601 = ~pi38 & ~n18600;
  assign n18602 = pi39 & pi142;
  assign n18603 = pi38 & ~n18602;
  assign n18604 = ~pi39 & ~n18574;
  assign n18605 = pi735 & n17940;
  assign n18606 = ~n18604 & ~n18605;
  assign n18607 = n18603 & n18606;
  assign n18608 = n3267 & ~n18607;
  assign n18609 = ~n18601 & n18608;
  assign n18610 = ~n18439 & ~n18609;
  assign n18611 = pi625 & n18610;
  assign n18612 = ~n6189 & ~n18561;
  assign n18613 = n6189 & n18545;
  assign n18614 = ~n18612 & ~n18613;
  assign n18615 = ~n3329 & ~n18614;
  assign n18616 = n3329 & ~n18569;
  assign n18617 = ~pi215 & ~n18616;
  assign n18618 = ~n18615 & n18617;
  assign n18619 = ~n6189 & n18504;
  assign n18620 = n6189 & n18523;
  assign n18621 = pi215 & ~n18620;
  assign n18622 = ~n18619 & n18621;
  assign n18623 = ~n18618 & ~n18622;
  assign n18624 = pi299 & ~n18623;
  assign n18625 = n6215 & n18545;
  assign n18626 = ~n6215 & ~n18561;
  assign n18627 = ~n3052 & ~n18626;
  assign n18628 = ~n18625 & n18627;
  assign n18629 = n3052 & n18569;
  assign n18630 = ~pi223 & ~n18629;
  assign n18631 = ~n18628 & n18630;
  assign n18632 = ~n6215 & ~n18504;
  assign n18633 = n6215 & ~n18523;
  assign n18634 = pi223 & ~n18633;
  assign n18635 = ~n18632 & n18634;
  assign n18636 = ~pi299 & ~n18635;
  assign n18637 = ~n18631 & n18636;
  assign n18638 = pi39 & ~n18637;
  assign n18639 = ~n18624 & n18638;
  assign n18640 = ~pi39 & n18485;
  assign n18641 = ~pi38 & ~n18640;
  assign n18642 = ~n18639 & n18641;
  assign n18643 = n18603 & ~n18604;
  assign n18644 = n3267 & ~n18643;
  assign n18645 = ~n18642 & n18644;
  assign n18646 = ~n18439 & ~n18645;
  assign n18647 = ~pi625 & n18646;
  assign n18648 = pi1153 & ~n18647;
  assign n18649 = ~n18611 & n18648;
  assign n18650 = ~pi142 & ~n17307;
  assign n18651 = pi142 & ~n17343;
  assign n18652 = ~n18650 & ~n18651;
  assign n18653 = pi735 & ~n18652;
  assign n18654 = ~pi735 & ~n18543;
  assign n18655 = ~n18653 & ~n18654;
  assign n18656 = n6215 & n18655;
  assign n18657 = ~pi142 & n17300;
  assign n18658 = pi142 & n17349;
  assign n18659 = ~n18657 & ~n18658;
  assign n18660 = pi735 & ~n18659;
  assign n18661 = ~pi735 & ~n18559;
  assign n18662 = ~n18660 & ~n18661;
  assign n18663 = ~n6215 & n18662;
  assign n18664 = ~n3052 & ~n18663;
  assign n18665 = ~n18656 & n18664;
  assign n18666 = pi735 & n16786;
  assign n18667 = n16517 & n18666;
  assign n18668 = ~n18567 & ~n18667;
  assign n18669 = n3052 & n18668;
  assign n18670 = ~pi223 & ~n18669;
  assign n18671 = ~n18665 & n18670;
  assign n18672 = ~pi735 & ~n18499;
  assign n18673 = pi142 & ~n17359;
  assign n18674 = ~pi142 & n16858;
  assign n18675 = n16857 & n18674;
  assign n18676 = pi735 & ~n18675;
  assign n18677 = ~n18673 & n18676;
  assign n18678 = ~n18672 & ~n18677;
  assign n18679 = ~n6215 & ~n18678;
  assign n18680 = ~pi735 & ~n18518;
  assign n18681 = pi142 & ~n17361;
  assign n18682 = pi735 & ~n18674;
  assign n18683 = ~n18681 & n18682;
  assign n18684 = ~n18680 & ~n18683;
  assign n18685 = n6215 & ~n18684;
  assign n18686 = pi223 & ~n18685;
  assign n18687 = ~n18679 & n18686;
  assign n18688 = ~pi299 & ~n18687;
  assign n18689 = ~n18671 & n18688;
  assign n18690 = n6189 & n18655;
  assign n18691 = ~n6189 & n18662;
  assign n18692 = ~n3329 & ~n18691;
  assign n18693 = ~n18690 & n18692;
  assign n18694 = n3329 & n18668;
  assign n18695 = ~pi215 & ~n18694;
  assign n18696 = ~n18693 & n18695;
  assign n18697 = ~n6189 & ~n18678;
  assign n18698 = n6189 & ~n18684;
  assign n18699 = pi215 & ~n18698;
  assign n18700 = ~n18697 & n18699;
  assign n18701 = pi299 & ~n18700;
  assign n18702 = ~n18696 & n18701;
  assign n18703 = pi39 & ~n18702;
  assign n18704 = ~n18689 & n18703;
  assign n18705 = pi142 & n17078;
  assign n18706 = ~pi142 & ~n17057;
  assign n18707 = pi735 & ~n18706;
  assign n18708 = ~n18705 & n18707;
  assign n18709 = pi142 & ~pi735;
  assign n18710 = ~n17120 & n18709;
  assign n18711 = ~n18708 & ~n18710;
  assign n18712 = ~pi39 & ~n18711;
  assign n18713 = ~pi38 & ~n18712;
  assign n18714 = ~n18704 & n18713;
  assign n18715 = n3095 & n18666;
  assign n18716 = ~n18571 & ~n18715;
  assign n18717 = ~pi39 & ~n18716;
  assign n18718 = n18603 & ~n18717;
  assign n18719 = n3267 & ~n18718;
  assign n18720 = ~n18714 & n18719;
  assign n18721 = ~n18439 & ~n18720;
  assign n18722 = ~pi625 & n18721;
  assign n18723 = n3267 & ~n17398;
  assign n18724 = pi142 & ~n18723;
  assign n18725 = pi39 & ~n17180;
  assign n18726 = pi142 & ~n17954;
  assign n18727 = ~n18725 & n18726;
  assign n18728 = ~n6189 & ~n18499;
  assign n18729 = n6189 & ~n18518;
  assign n18730 = pi215 & ~n18729;
  assign n18731 = ~n18728 & n18730;
  assign n18732 = ~n6189 & ~n18559;
  assign n18733 = n6189 & ~n18543;
  assign n18734 = ~n18732 & ~n18733;
  assign n18735 = ~n3329 & ~n18734;
  assign n18736 = n3329 & ~n18567;
  assign n18737 = ~pi215 & ~n18736;
  assign n18738 = ~n18735 & n18737;
  assign n18739 = ~n18731 & ~n18738;
  assign n18740 = pi39 & pi299;
  assign n18741 = ~n18739 & n18740;
  assign n18742 = ~n18727 & ~n18741;
  assign n18743 = n14755 & ~n18742;
  assign n18744 = ~n18724 & ~n18743;
  assign n18745 = pi625 & n18744;
  assign n18746 = ~pi1153 & ~n18745;
  assign n18747 = ~n18722 & n18746;
  assign n18748 = pi608 & ~n18747;
  assign n18749 = ~n18649 & n18748;
  assign n18750 = ~pi625 & n18610;
  assign n18751 = pi625 & n18646;
  assign n18752 = ~pi1153 & ~n18751;
  assign n18753 = ~n18750 & n18752;
  assign n18754 = pi625 & n18721;
  assign n18755 = ~pi625 & n18744;
  assign n18756 = pi1153 & ~n18755;
  assign n18757 = ~n18754 & n18756;
  assign n18758 = ~pi608 & ~n18757;
  assign n18759 = ~n18753 & n18758;
  assign n18760 = ~n18749 & ~n18759;
  assign n18761 = pi778 & ~n18760;
  assign n18762 = ~pi778 & n18610;
  assign n18763 = ~n18761 & ~n18762;
  assign n18764 = ~pi609 & ~n18763;
  assign n18765 = ~pi778 & ~n18721;
  assign n18766 = ~n18747 & ~n18757;
  assign n18767 = pi778 & ~n18766;
  assign n18768 = ~n18765 & ~n18767;
  assign n18769 = pi609 & n18768;
  assign n18770 = ~pi1155 & ~n18769;
  assign n18771 = ~n18764 & n18770;
  assign n18772 = ~n17439 & ~n18744;
  assign n18773 = ~n17438 & ~n18646;
  assign n18774 = pi609 & n18773;
  assign n18775 = ~n18772 & ~n18774;
  assign n18776 = pi1155 & ~n18775;
  assign n18777 = ~pi660 & ~n18776;
  assign n18778 = ~n18771 & n18777;
  assign n18779 = pi609 & ~n18763;
  assign n18780 = ~pi609 & n18768;
  assign n18781 = pi1155 & ~n18780;
  assign n18782 = ~n18779 & n18781;
  assign n18783 = ~n17451 & ~n18744;
  assign n18784 = ~pi609 & n18773;
  assign n18785 = ~n18783 & ~n18784;
  assign n18786 = ~pi1155 & ~n18785;
  assign n18787 = pi660 & ~n18786;
  assign n18788 = ~n18782 & n18787;
  assign n18789 = ~n18778 & ~n18788;
  assign n18790 = pi785 & ~n18789;
  assign n18791 = ~pi785 & ~n18763;
  assign n18792 = ~n18790 & ~n18791;
  assign n18793 = ~pi618 & ~n18792;
  assign n18794 = ~n17466 & n18768;
  assign n18795 = n17466 & n18744;
  assign n18796 = ~n18794 & ~n18795;
  assign n18797 = pi618 & ~n18796;
  assign n18798 = ~pi1154 & ~n18797;
  assign n18799 = ~n18793 & n18798;
  assign n18800 = n17438 & ~n18744;
  assign n18801 = ~n18773 & ~n18800;
  assign n18802 = ~pi785 & ~n18801;
  assign n18803 = ~n18776 & ~n18786;
  assign n18804 = pi785 & ~n18803;
  assign n18805 = ~n18802 & ~n18804;
  assign n18806 = pi618 & n18805;
  assign n18807 = ~pi618 & n18744;
  assign n18808 = pi1154 & ~n18807;
  assign n18809 = ~n18806 & n18808;
  assign n18810 = ~pi627 & ~n18809;
  assign n18811 = ~n18799 & n18810;
  assign n18812 = pi618 & ~n18792;
  assign n18813 = ~pi618 & ~n18796;
  assign n18814 = pi1154 & ~n18813;
  assign n18815 = ~n18812 & n18814;
  assign n18816 = ~pi618 & n18805;
  assign n18817 = pi618 & n18744;
  assign n18818 = ~pi1154 & ~n18817;
  assign n18819 = ~n18816 & n18818;
  assign n18820 = pi627 & ~n18819;
  assign n18821 = ~n18815 & n18820;
  assign n18822 = ~n18811 & ~n18821;
  assign n18823 = pi781 & ~n18822;
  assign n18824 = ~pi781 & ~n18792;
  assign n18825 = ~n18823 & ~n18824;
  assign n18826 = ~pi619 & ~n18825;
  assign n18827 = n17503 & ~n18744;
  assign n18828 = ~n17503 & n18796;
  assign n18829 = ~n18827 & ~n18828;
  assign n18830 = pi619 & n18829;
  assign n18831 = ~pi1159 & ~n18830;
  assign n18832 = ~n18826 & n18831;
  assign n18833 = ~pi781 & ~n18805;
  assign n18834 = ~n18809 & ~n18819;
  assign n18835 = pi781 & ~n18834;
  assign n18836 = ~n18833 & ~n18835;
  assign n18837 = pi619 & n18836;
  assign n18838 = ~pi619 & n18744;
  assign n18839 = pi1159 & ~n18838;
  assign n18840 = ~n18837 & n18839;
  assign n18841 = ~pi648 & ~n18840;
  assign n18842 = ~n18832 & n18841;
  assign n18843 = pi619 & ~n18825;
  assign n18844 = ~pi619 & n18829;
  assign n18845 = pi1159 & ~n18844;
  assign n18846 = ~n18843 & n18845;
  assign n18847 = ~pi619 & n18836;
  assign n18848 = pi619 & n18744;
  assign n18849 = ~pi1159 & ~n18848;
  assign n18850 = ~n18847 & n18849;
  assign n18851 = pi648 & ~n18850;
  assign n18852 = ~n18846 & n18851;
  assign n18853 = ~n18842 & ~n18852;
  assign n18854 = pi789 & ~n18853;
  assign n18855 = ~pi789 & ~n18825;
  assign n18856 = ~n18854 & ~n18855;
  assign n18857 = ~pi788 & n18856;
  assign n18858 = ~pi626 & n18856;
  assign n18859 = ~n17539 & n18829;
  assign n18860 = n17539 & n18744;
  assign n18861 = ~n18859 & ~n18860;
  assign n18862 = pi626 & n18861;
  assign n18863 = ~pi641 & ~n18862;
  assign n18864 = ~n18858 & n18863;
  assign n18865 = ~pi789 & ~n18836;
  assign n18866 = ~n18840 & ~n18850;
  assign n18867 = pi789 & ~n18866;
  assign n18868 = ~n18865 & ~n18867;
  assign n18869 = ~pi626 & n18868;
  assign n18870 = pi626 & n18744;
  assign n18871 = ~pi1158 & ~n18870;
  assign n18872 = ~n18869 & n18871;
  assign n18873 = ~n17546 & ~n18872;
  assign n18874 = ~n18864 & ~n18873;
  assign n18875 = pi626 & n18856;
  assign n18876 = ~pi626 & n18861;
  assign n18877 = pi641 & ~n18876;
  assign n18878 = ~n18875 & n18877;
  assign n18879 = pi626 & n18868;
  assign n18880 = ~pi626 & n18744;
  assign n18881 = pi1158 & ~n18880;
  assign n18882 = ~n18879 & n18881;
  assign n18883 = ~n17561 & ~n18882;
  assign n18884 = ~n18878 & ~n18883;
  assign n18885 = ~n18874 & ~n18884;
  assign n18886 = pi788 & ~n18885;
  assign n18887 = ~n18857 & ~n18886;
  assign n18888 = ~pi628 & n18887;
  assign n18889 = ~n18872 & ~n18882;
  assign n18890 = pi788 & ~n18889;
  assign n18891 = ~pi788 & ~n18868;
  assign n18892 = ~n18890 & ~n18891;
  assign n18893 = pi628 & n18892;
  assign n18894 = ~pi1156 & ~n18893;
  assign n18895 = ~n18888 & n18894;
  assign n18896 = ~n17582 & ~n18861;
  assign n18897 = n17582 & n18744;
  assign n18898 = ~n18896 & ~n18897;
  assign n18899 = pi628 & ~n18898;
  assign n18900 = ~pi628 & n18744;
  assign n18901 = pi1156 & ~n18900;
  assign n18902 = ~n18899 & n18901;
  assign n18903 = ~pi629 & ~n18902;
  assign n18904 = ~n18895 & n18903;
  assign n18905 = pi628 & n18887;
  assign n18906 = ~pi628 & n18892;
  assign n18907 = pi1156 & ~n18906;
  assign n18908 = ~n18905 & n18907;
  assign n18909 = ~pi628 & ~n18898;
  assign n18910 = pi628 & n18744;
  assign n18911 = ~pi1156 & ~n18910;
  assign n18912 = ~n18909 & n18911;
  assign n18913 = pi629 & ~n18912;
  assign n18914 = ~n18908 & n18913;
  assign n18915 = ~n18904 & ~n18914;
  assign n18916 = pi792 & ~n18915;
  assign n18917 = ~pi792 & n18887;
  assign n18918 = ~n18916 & ~n18917;
  assign n18919 = ~pi647 & ~n18918;
  assign n18920 = ~n17610 & n18892;
  assign n18921 = n17610 & n18744;
  assign n18922 = ~n18920 & ~n18921;
  assign n18923 = pi647 & ~n18922;
  assign n18924 = ~pi1157 & ~n18923;
  assign n18925 = ~n18919 & n18924;
  assign n18926 = ~pi792 & n18898;
  assign n18927 = ~n18902 & ~n18912;
  assign n18928 = pi792 & ~n18927;
  assign n18929 = ~n18926 & ~n18928;
  assign n18930 = pi647 & n18929;
  assign n18931 = ~pi647 & n18744;
  assign n18932 = pi1157 & ~n18931;
  assign n18933 = ~n18930 & n18932;
  assign n18934 = ~pi630 & ~n18933;
  assign n18935 = ~n18925 & n18934;
  assign n18936 = pi647 & ~n18918;
  assign n18937 = ~pi647 & ~n18922;
  assign n18938 = pi1157 & ~n18937;
  assign n18939 = ~n18936 & n18938;
  assign n18940 = ~pi647 & n18929;
  assign n18941 = pi647 & n18744;
  assign n18942 = ~pi1157 & ~n18941;
  assign n18943 = ~n18940 & n18942;
  assign n18944 = pi630 & ~n18943;
  assign n18945 = ~n18939 & n18944;
  assign n18946 = ~n18935 & ~n18945;
  assign n18947 = pi787 & ~n18946;
  assign n18948 = ~pi787 & ~n18918;
  assign n18949 = ~n18947 & ~n18948;
  assign n18950 = ~pi644 & ~n18949;
  assign n18951 = ~pi787 & ~n18929;
  assign n18952 = ~n18933 & ~n18943;
  assign n18953 = pi787 & ~n18952;
  assign n18954 = ~n18951 & ~n18953;
  assign n18955 = pi644 & n18954;
  assign n18956 = ~pi715 & ~n18955;
  assign n18957 = ~n18950 & n18956;
  assign n18958 = n17652 & ~n18744;
  assign n18959 = ~n17652 & n18922;
  assign n18960 = ~n18958 & ~n18959;
  assign n18961 = ~pi644 & n18960;
  assign n18962 = pi644 & n18744;
  assign n18963 = pi715 & ~n18962;
  assign n18964 = ~n18961 & n18963;
  assign n18965 = ~pi1160 & ~n18964;
  assign n18966 = ~n18957 & n18965;
  assign n18967 = pi644 & ~n18949;
  assign n18968 = ~pi644 & n18954;
  assign n18969 = pi715 & ~n18968;
  assign n18970 = ~n18967 & n18969;
  assign n18971 = pi644 & n18960;
  assign n18972 = ~pi644 & n18744;
  assign n18973 = ~pi715 & ~n18972;
  assign n18974 = ~n18971 & n18973;
  assign n18975 = pi1160 & ~n18974;
  assign n18976 = ~n18970 & n18975;
  assign n18977 = pi790 & ~n18976;
  assign n18978 = ~n18966 & n18977;
  assign n18979 = ~pi790 & n18949;
  assign n18980 = n6286 & ~n18979;
  assign n18981 = ~n18978 & n18980;
  assign n18982 = ~pi142 & ~n6286;
  assign n18983 = ~pi57 & ~n18982;
  assign n18984 = ~n18981 & n18983;
  assign n18985 = pi57 & pi142;
  assign n18986 = ~pi832 & ~n18985;
  assign n18987 = ~n18984 & n18986;
  assign n18988 = ~n17438 & n18572;
  assign n18989 = pi609 & n18988;
  assign n18990 = pi142 & ~n2754;
  assign n18991 = pi1155 & ~n18990;
  assign n18992 = ~n18989 & n18991;
  assign n18993 = ~pi609 & n18988;
  assign n18994 = ~pi1155 & ~n18990;
  assign n18995 = ~n18993 & n18994;
  assign n18996 = ~n18992 & ~n18995;
  assign n18997 = pi785 & ~n18996;
  assign n18998 = ~pi785 & ~n18990;
  assign n18999 = ~n18988 & n18998;
  assign n19000 = ~n18997 & ~n18999;
  assign n19001 = ~pi781 & ~n19000;
  assign n19002 = pi618 & n19000;
  assign n19003 = ~pi618 & n18990;
  assign n19004 = pi1154 & ~n19003;
  assign n19005 = ~n19002 & n19004;
  assign n19006 = ~pi618 & n19000;
  assign n19007 = pi618 & n18990;
  assign n19008 = ~pi1154 & ~n19007;
  assign n19009 = ~n19006 & n19008;
  assign n19010 = ~n19005 & ~n19009;
  assign n19011 = pi781 & ~n19010;
  assign n19012 = ~n19001 & ~n19011;
  assign n19013 = ~pi789 & ~n19012;
  assign n19014 = pi619 & n19012;
  assign n19015 = ~pi619 & n18990;
  assign n19016 = pi1159 & ~n19015;
  assign n19017 = ~n19014 & n19016;
  assign n19018 = ~pi619 & n19012;
  assign n19019 = pi619 & n18990;
  assign n19020 = ~pi1159 & ~n19019;
  assign n19021 = ~n19018 & n19020;
  assign n19022 = ~n19017 & ~n19021;
  assign n19023 = pi789 & ~n19022;
  assign n19024 = ~n19013 & ~n19023;
  assign n19025 = pi626 & n19024;
  assign n19026 = ~pi626 & n18990;
  assign n19027 = pi1158 & ~n19026;
  assign n19028 = ~n19025 & n19027;
  assign n19029 = ~pi626 & n19024;
  assign n19030 = pi626 & n18990;
  assign n19031 = ~pi1158 & ~n19030;
  assign n19032 = ~n19029 & n19031;
  assign n19033 = ~n19028 & ~n19032;
  assign n19034 = ~n17581 & n19033;
  assign n19035 = ~pi625 & pi1153;
  assign n19036 = pi625 & ~pi1153;
  assign n19037 = ~n19035 & ~n19036;
  assign n19038 = pi778 & ~n19037;
  assign n19039 = n18666 & ~n19038;
  assign n19040 = ~n18990 & ~n19039;
  assign n19041 = ~n17692 & ~n19040;
  assign n19042 = ~n17694 & n19041;
  assign n19043 = ~n17696 & n17704;
  assign n19044 = n19042 & n19043;
  assign n19045 = ~n19034 & ~n19044;
  assign n19046 = pi788 & ~n19045;
  assign n19047 = pi735 & n16787;
  assign n19048 = pi625 & n19047;
  assign n19049 = ~n18572 & ~n18990;
  assign n19050 = ~n19047 & n19049;
  assign n19051 = ~n19048 & ~n19050;
  assign n19052 = ~pi1153 & ~n19051;
  assign n19053 = pi625 & n18666;
  assign n19054 = pi1153 & ~n18990;
  assign n19055 = ~n19053 & n19054;
  assign n19056 = ~pi608 & ~n19055;
  assign n19057 = ~n19052 & n19056;
  assign n19058 = ~n18572 & ~n19048;
  assign n19059 = pi1153 & ~n19058;
  assign n19060 = ~pi625 & ~pi1153;
  assign n19061 = n18666 & n19060;
  assign n19062 = ~n18990 & ~n19061;
  assign n19063 = ~n19059 & n19062;
  assign n19064 = pi608 & ~n19063;
  assign n19065 = ~n19057 & ~n19064;
  assign n19066 = pi778 & ~n19065;
  assign n19067 = ~pi778 & ~n19050;
  assign n19068 = ~n19066 & ~n19067;
  assign n19069 = ~pi609 & ~n19068;
  assign n19070 = pi609 & ~n19040;
  assign n19071 = ~pi1155 & ~n19070;
  assign n19072 = ~n19069 & n19071;
  assign n19073 = ~pi660 & ~n18992;
  assign n19074 = ~n19072 & n19073;
  assign n19075 = pi609 & ~n19068;
  assign n19076 = ~pi609 & ~n19040;
  assign n19077 = pi1155 & ~n19076;
  assign n19078 = ~n19075 & n19077;
  assign n19079 = pi660 & ~n18995;
  assign n19080 = ~n19078 & n19079;
  assign n19081 = ~n19074 & ~n19080;
  assign n19082 = pi785 & ~n19081;
  assign n19083 = ~pi785 & ~n19068;
  assign n19084 = ~n19082 & ~n19083;
  assign n19085 = ~pi618 & ~n19084;
  assign n19086 = pi618 & n19041;
  assign n19087 = ~pi1154 & ~n19086;
  assign n19088 = ~n19085 & n19087;
  assign n19089 = ~pi627 & ~n19005;
  assign n19090 = ~n19088 & n19089;
  assign n19091 = pi618 & ~n19084;
  assign n19092 = ~pi618 & n19041;
  assign n19093 = pi1154 & ~n19092;
  assign n19094 = ~n19091 & n19093;
  assign n19095 = pi627 & ~n19009;
  assign n19096 = ~n19094 & n19095;
  assign n19097 = ~n19090 & ~n19096;
  assign n19098 = pi781 & ~n19097;
  assign n19099 = ~pi781 & ~n19084;
  assign n19100 = ~n19098 & ~n19099;
  assign n19101 = pi619 & ~n19100;
  assign n19102 = ~pi619 & n19042;
  assign n19103 = pi1159 & ~n19102;
  assign n19104 = ~n19101 & n19103;
  assign n19105 = pi648 & ~n19021;
  assign n19106 = ~n19104 & n19105;
  assign n19107 = ~pi619 & ~n19100;
  assign n19108 = pi619 & n19042;
  assign n19109 = ~pi1159 & ~n19108;
  assign n19110 = ~n19107 & n19109;
  assign n19111 = ~pi648 & ~n19017;
  assign n19112 = ~n19110 & n19111;
  assign n19113 = pi789 & ~n19112;
  assign n19114 = ~n19106 & n19113;
  assign n19115 = ~pi789 & n19100;
  assign n19116 = n17817 & ~n19115;
  assign n19117 = ~n19114 & n19116;
  assign n19118 = ~n19046 & ~n19117;
  assign n19119 = ~pi628 & n19118;
  assign n19120 = ~pi788 & ~n19024;
  assign n19121 = pi788 & ~n19033;
  assign n19122 = ~n19120 & ~n19121;
  assign n19123 = pi628 & ~n19122;
  assign n19124 = ~pi1156 & ~n19123;
  assign n19125 = ~n19119 & n19124;
  assign n19126 = ~n17539 & ~n17582;
  assign n19127 = ~n17466 & ~n17503;
  assign n19128 = n19126 & n19127;
  assign n19129 = ~n19040 & n19128;
  assign n19130 = pi628 & n19129;
  assign n19131 = ~n18990 & ~n19130;
  assign n19132 = pi1156 & ~n19131;
  assign n19133 = ~pi629 & ~n19132;
  assign n19134 = ~n19125 & n19133;
  assign n19135 = pi628 & n19118;
  assign n19136 = ~pi628 & ~n19122;
  assign n19137 = pi1156 & ~n19136;
  assign n19138 = ~n19135 & n19137;
  assign n19139 = ~pi628 & n19129;
  assign n19140 = ~n18990 & ~n19139;
  assign n19141 = ~pi1156 & ~n19140;
  assign n19142 = pi629 & ~n19141;
  assign n19143 = ~n19138 & n19142;
  assign n19144 = ~n19134 & ~n19143;
  assign n19145 = pi792 & ~n19144;
  assign n19146 = ~pi792 & n19118;
  assign n19147 = ~n19145 & ~n19146;
  assign n19148 = ~pi647 & n19147;
  assign n19149 = ~n17610 & n19122;
  assign n19150 = n17610 & n18990;
  assign n19151 = ~n19149 & ~n19150;
  assign n19152 = pi647 & ~n19151;
  assign n19153 = ~pi1157 & ~n19152;
  assign n19154 = ~n19148 & n19153;
  assign n19155 = ~pi628 & ~pi1156;
  assign n19156 = pi628 & pi1156;
  assign n19157 = pi792 & ~n19156;
  assign n19158 = ~n19155 & n19157;
  assign n19159 = n19129 & ~n19158;
  assign n19160 = pi647 & n19159;
  assign n19161 = pi1157 & ~n18990;
  assign n19162 = ~n19160 & n19161;
  assign n19163 = ~pi630 & ~n19162;
  assign n19164 = ~n19154 & n19163;
  assign n19165 = pi647 & n19147;
  assign n19166 = ~pi647 & ~n19151;
  assign n19167 = pi1157 & ~n19166;
  assign n19168 = ~n19165 & n19167;
  assign n19169 = ~pi647 & n19159;
  assign n19170 = ~pi1157 & ~n18990;
  assign n19171 = ~n19169 & n19170;
  assign n19172 = pi630 & ~n19171;
  assign n19173 = ~n19168 & n19172;
  assign n19174 = ~n19164 & ~n19173;
  assign n19175 = pi787 & ~n19174;
  assign n19176 = ~pi787 & n19147;
  assign n19177 = ~n19175 & ~n19176;
  assign n19178 = pi644 & ~n19177;
  assign n19179 = ~pi647 & pi1157;
  assign n19180 = pi647 & ~pi1157;
  assign n19181 = ~n19179 & ~n19180;
  assign n19182 = pi787 & ~n19181;
  assign n19183 = n19159 & ~n19182;
  assign n19184 = ~n18990 & ~n19183;
  assign n19185 = ~pi644 & ~n19184;
  assign n19186 = pi715 & ~n19185;
  assign n19187 = ~n19178 & n19186;
  assign n19188 = n17652 & ~n18990;
  assign n19189 = ~n17652 & n19151;
  assign n19190 = ~n19188 & ~n19189;
  assign n19191 = pi644 & n19190;
  assign n19192 = ~pi644 & n18990;
  assign n19193 = ~pi715 & ~n19192;
  assign n19194 = ~n19191 & n19193;
  assign n19195 = pi1160 & ~n19194;
  assign n19196 = ~n19187 & n19195;
  assign n19197 = ~pi644 & ~n19177;
  assign n19198 = pi644 & ~n19184;
  assign n19199 = ~pi715 & ~n19198;
  assign n19200 = ~n19197 & n19199;
  assign n19201 = ~pi644 & n19190;
  assign n19202 = pi644 & n18990;
  assign n19203 = pi715 & ~n19202;
  assign n19204 = ~n19201 & n19203;
  assign n19205 = ~pi1160 & ~n19204;
  assign n19206 = ~n19200 & n19205;
  assign n19207 = ~n19196 & ~n19206;
  assign n19208 = pi790 & ~n19207;
  assign n19209 = ~pi790 & ~n19177;
  assign n19210 = pi832 & ~n19209;
  assign n19211 = ~n19208 & n19210;
  assign po299 = ~n18987 & ~n19211;
  assign n19213 = pi143 & ~n3267;
  assign n19214 = ~pi143 & ~n17399;
  assign n19215 = pi774 & ~n19214;
  assign n19216 = n6109 & n16784;
  assign n19217 = pi38 & n19216;
  assign n19218 = ~pi38 & n17275;
  assign n19219 = pi143 & ~n19218;
  assign n19220 = ~pi38 & ~n17242;
  assign n19221 = n6234 & n16740;
  assign n19222 = pi38 & ~n19221;
  assign n19223 = ~n19220 & ~n19222;
  assign n19224 = ~pi143 & ~pi774;
  assign n19225 = n19223 & n19224;
  assign n19226 = ~n19219 & ~n19225;
  assign n19227 = ~n19217 & ~n19226;
  assign n19228 = ~n19215 & ~n19227;
  assign n19229 = ~pi687 & n19228;
  assign n19230 = ~n16667 & n17280;
  assign n19231 = pi38 & n19230;
  assign n19232 = pi39 & ~n16687;
  assign n19233 = ~pi39 & ~n17088;
  assign n19234 = ~n19232 & ~n19233;
  assign n19235 = ~pi38 & ~n19234;
  assign n19236 = ~n19231 & ~n19235;
  assign n19237 = ~pi143 & n19236;
  assign n19238 = ~pi39 & ~n17059;
  assign n19239 = pi39 & ~n16799;
  assign n19240 = ~n19238 & ~n19239;
  assign n19241 = ~pi38 & n19240;
  assign n19242 = pi143 & n19241;
  assign n19243 = pi38 & n17940;
  assign n19244 = pi774 & ~n19243;
  assign n19245 = ~n19242 & n19244;
  assign n19246 = ~n19237 & n19245;
  assign n19247 = n6234 & ~n16788;
  assign n19248 = pi38 & ~n19247;
  assign n19249 = pi39 & ~n16879;
  assign n19250 = ~n17057 & n17246;
  assign n19251 = ~n19249 & ~n19250;
  assign n19252 = ~pi38 & ~n19251;
  assign n19253 = ~n19248 & ~n19252;
  assign n19254 = pi143 & n19253;
  assign n19255 = pi39 & ~n16944;
  assign n19256 = ~pi39 & ~n17092;
  assign n19257 = ~pi38 & n19256;
  assign n19258 = ~pi39 & n16905;
  assign n19259 = pi38 & ~n19258;
  assign n19260 = ~n19257 & ~n19259;
  assign n19261 = ~n19255 & n19260;
  assign n19262 = ~pi143 & ~n19261;
  assign n19263 = ~pi774 & ~n19262;
  assign n19264 = ~n19254 & n19263;
  assign n19265 = pi687 & ~n19264;
  assign n19266 = ~n19246 & n19265;
  assign n19267 = n3267 & ~n19266;
  assign n19268 = ~n19229 & n19267;
  assign n19269 = ~n19213 & ~n19268;
  assign n19270 = ~pi625 & n19269;
  assign n19271 = n3267 & ~n19228;
  assign n19272 = ~n19213 & ~n19271;
  assign n19273 = pi625 & n19272;
  assign n19274 = ~pi1153 & ~n19273;
  assign n19275 = ~n19270 & n19274;
  assign n19276 = ~pi143 & n17972;
  assign n19277 = pi143 & ~n17976;
  assign n19278 = ~pi38 & ~n19277;
  assign n19279 = ~n19276 & n19278;
  assign n19280 = ~pi143 & ~n17280;
  assign n19281 = n17392 & ~n19280;
  assign n19282 = pi687 & ~n19281;
  assign n19283 = ~n19279 & n19282;
  assign n19284 = ~pi687 & n19214;
  assign n19285 = n3267 & ~n19284;
  assign n19286 = ~n19283 & n19285;
  assign n19287 = ~n19213 & ~n19286;
  assign n19288 = pi625 & n19287;
  assign n19289 = ~pi143 & ~n17406;
  assign n19290 = ~pi625 & n19289;
  assign n19291 = pi1153 & ~n19290;
  assign n19292 = ~n19288 & n19291;
  assign n19293 = ~pi608 & ~n19292;
  assign n19294 = ~n19275 & n19293;
  assign n19295 = pi625 & n19269;
  assign n19296 = ~pi625 & n19272;
  assign n19297 = pi1153 & ~n19296;
  assign n19298 = ~n19295 & n19297;
  assign n19299 = ~pi625 & n19287;
  assign n19300 = pi625 & n19289;
  assign n19301 = ~pi1153 & ~n19300;
  assign n19302 = ~n19299 & n19301;
  assign n19303 = pi608 & ~n19302;
  assign n19304 = ~n19298 & n19303;
  assign n19305 = ~n19294 & ~n19304;
  assign n19306 = pi778 & ~n19305;
  assign n19307 = ~pi778 & n19269;
  assign n19308 = ~n19306 & ~n19307;
  assign n19309 = ~pi609 & ~n19308;
  assign n19310 = ~pi778 & ~n19287;
  assign n19311 = ~n19292 & ~n19302;
  assign n19312 = pi778 & ~n19311;
  assign n19313 = ~n19310 & ~n19312;
  assign n19314 = pi609 & n19313;
  assign n19315 = ~pi1155 & ~n19314;
  assign n19316 = ~n19309 & n19315;
  assign n19317 = ~n17439 & ~n19289;
  assign n19318 = ~n17438 & ~n19272;
  assign n19319 = pi609 & n19318;
  assign n19320 = ~n19317 & ~n19319;
  assign n19321 = pi1155 & ~n19320;
  assign n19322 = ~pi660 & ~n19321;
  assign n19323 = ~n19316 & n19322;
  assign n19324 = pi609 & ~n19308;
  assign n19325 = ~pi609 & n19313;
  assign n19326 = pi1155 & ~n19325;
  assign n19327 = ~n19324 & n19326;
  assign n19328 = ~n17451 & ~n19289;
  assign n19329 = ~pi609 & n19318;
  assign n19330 = ~n19328 & ~n19329;
  assign n19331 = ~pi1155 & ~n19330;
  assign n19332 = pi660 & ~n19331;
  assign n19333 = ~n19327 & n19332;
  assign n19334 = ~n19323 & ~n19333;
  assign n19335 = pi785 & ~n19334;
  assign n19336 = ~pi785 & ~n19308;
  assign n19337 = ~n19335 & ~n19336;
  assign n19338 = ~pi618 & ~n19337;
  assign n19339 = ~n17466 & ~n19313;
  assign n19340 = n17466 & ~n19289;
  assign n19341 = ~n19339 & ~n19340;
  assign n19342 = pi618 & n19341;
  assign n19343 = ~pi1154 & ~n19342;
  assign n19344 = ~n19338 & n19343;
  assign n19345 = n17438 & ~n19289;
  assign n19346 = ~n19318 & ~n19345;
  assign n19347 = ~pi785 & ~n19346;
  assign n19348 = ~n19321 & ~n19331;
  assign n19349 = pi785 & ~n19348;
  assign n19350 = ~n19347 & ~n19349;
  assign n19351 = pi618 & n19350;
  assign n19352 = ~pi618 & n19289;
  assign n19353 = pi1154 & ~n19352;
  assign n19354 = ~n19351 & n19353;
  assign n19355 = ~pi627 & ~n19354;
  assign n19356 = ~n19344 & n19355;
  assign n19357 = pi618 & ~n19337;
  assign n19358 = ~pi618 & n19341;
  assign n19359 = pi1154 & ~n19358;
  assign n19360 = ~n19357 & n19359;
  assign n19361 = ~pi618 & n19350;
  assign n19362 = pi618 & n19289;
  assign n19363 = ~pi1154 & ~n19362;
  assign n19364 = ~n19361 & n19363;
  assign n19365 = pi627 & ~n19364;
  assign n19366 = ~n19360 & n19365;
  assign n19367 = ~n19356 & ~n19366;
  assign n19368 = pi781 & ~n19367;
  assign n19369 = ~pi781 & ~n19337;
  assign n19370 = ~n19368 & ~n19369;
  assign n19371 = ~pi619 & ~n19370;
  assign n19372 = ~n17503 & n19341;
  assign n19373 = n17503 & n19289;
  assign n19374 = ~n19372 & ~n19373;
  assign n19375 = pi619 & ~n19374;
  assign n19376 = ~pi1159 & ~n19375;
  assign n19377 = ~n19371 & n19376;
  assign n19378 = ~pi781 & ~n19350;
  assign n19379 = ~n19354 & ~n19364;
  assign n19380 = pi781 & ~n19379;
  assign n19381 = ~n19378 & ~n19380;
  assign n19382 = pi619 & n19381;
  assign n19383 = ~pi619 & n19289;
  assign n19384 = pi1159 & ~n19383;
  assign n19385 = ~n19382 & n19384;
  assign n19386 = ~pi648 & ~n19385;
  assign n19387 = ~n19377 & n19386;
  assign n19388 = pi619 & ~n19370;
  assign n19389 = ~pi619 & ~n19374;
  assign n19390 = pi1159 & ~n19389;
  assign n19391 = ~n19388 & n19390;
  assign n19392 = ~pi619 & n19381;
  assign n19393 = pi619 & n19289;
  assign n19394 = ~pi1159 & ~n19393;
  assign n19395 = ~n19392 & n19394;
  assign n19396 = pi648 & ~n19395;
  assign n19397 = ~n19391 & n19396;
  assign n19398 = ~n19387 & ~n19397;
  assign n19399 = pi789 & ~n19398;
  assign n19400 = ~pi789 & ~n19370;
  assign n19401 = ~n19399 & ~n19400;
  assign n19402 = ~pi788 & n19401;
  assign n19403 = ~pi626 & n19401;
  assign n19404 = n17539 & ~n19289;
  assign n19405 = ~n17539 & n19374;
  assign n19406 = ~n19404 & ~n19405;
  assign n19407 = pi626 & ~n19406;
  assign n19408 = ~pi641 & ~n19407;
  assign n19409 = ~n19403 & n19408;
  assign n19410 = ~pi789 & ~n19381;
  assign n19411 = ~n19385 & ~n19395;
  assign n19412 = pi789 & ~n19411;
  assign n19413 = ~n19410 & ~n19412;
  assign n19414 = ~pi626 & n19413;
  assign n19415 = pi626 & n19289;
  assign n19416 = ~pi1158 & ~n19415;
  assign n19417 = ~n19414 & n19416;
  assign n19418 = ~n17546 & ~n19417;
  assign n19419 = ~n19409 & ~n19418;
  assign n19420 = pi626 & n19401;
  assign n19421 = ~pi626 & ~n19406;
  assign n19422 = pi641 & ~n19421;
  assign n19423 = ~n19420 & n19422;
  assign n19424 = pi626 & n19413;
  assign n19425 = ~pi626 & n19289;
  assign n19426 = pi1158 & ~n19425;
  assign n19427 = ~n19424 & n19426;
  assign n19428 = ~n17561 & ~n19427;
  assign n19429 = ~n19423 & ~n19428;
  assign n19430 = ~n19419 & ~n19429;
  assign n19431 = pi788 & ~n19430;
  assign n19432 = ~n19402 & ~n19431;
  assign n19433 = ~pi628 & n19432;
  assign n19434 = ~n19417 & ~n19427;
  assign n19435 = pi788 & ~n19434;
  assign n19436 = ~pi788 & ~n19413;
  assign n19437 = ~n19435 & ~n19436;
  assign n19438 = pi628 & n19437;
  assign n19439 = ~pi1156 & ~n19438;
  assign n19440 = ~n19433 & n19439;
  assign n19441 = ~n17582 & n19406;
  assign n19442 = n17582 & n19289;
  assign n19443 = ~n19441 & ~n19442;
  assign n19444 = pi628 & ~n19443;
  assign n19445 = ~pi628 & n19289;
  assign n19446 = pi1156 & ~n19445;
  assign n19447 = ~n19444 & n19446;
  assign n19448 = ~pi629 & ~n19447;
  assign n19449 = ~n19440 & n19448;
  assign n19450 = pi628 & n19432;
  assign n19451 = ~pi628 & n19437;
  assign n19452 = pi1156 & ~n19451;
  assign n19453 = ~n19450 & n19452;
  assign n19454 = ~pi628 & ~n19443;
  assign n19455 = pi628 & n19289;
  assign n19456 = ~pi1156 & ~n19455;
  assign n19457 = ~n19454 & n19456;
  assign n19458 = pi629 & ~n19457;
  assign n19459 = ~n19453 & n19458;
  assign n19460 = ~n19449 & ~n19459;
  assign n19461 = pi792 & ~n19460;
  assign n19462 = ~pi792 & n19432;
  assign n19463 = ~n19461 & ~n19462;
  assign n19464 = ~pi647 & ~n19463;
  assign n19465 = ~n17610 & n19437;
  assign n19466 = n17610 & n19289;
  assign n19467 = ~n19465 & ~n19466;
  assign n19468 = pi647 & ~n19467;
  assign n19469 = ~pi1157 & ~n19468;
  assign n19470 = ~n19464 & n19469;
  assign n19471 = ~pi792 & n19443;
  assign n19472 = ~n19447 & ~n19457;
  assign n19473 = pi792 & ~n19472;
  assign n19474 = ~n19471 & ~n19473;
  assign n19475 = pi647 & n19474;
  assign n19476 = ~pi647 & n19289;
  assign n19477 = pi1157 & ~n19476;
  assign n19478 = ~n19475 & n19477;
  assign n19479 = ~pi630 & ~n19478;
  assign n19480 = ~n19470 & n19479;
  assign n19481 = pi647 & ~n19463;
  assign n19482 = ~pi647 & ~n19467;
  assign n19483 = pi1157 & ~n19482;
  assign n19484 = ~n19481 & n19483;
  assign n19485 = ~pi647 & n19474;
  assign n19486 = pi647 & n19289;
  assign n19487 = ~pi1157 & ~n19486;
  assign n19488 = ~n19485 & n19487;
  assign n19489 = pi630 & ~n19488;
  assign n19490 = ~n19484 & n19489;
  assign n19491 = ~n19480 & ~n19490;
  assign n19492 = pi787 & ~n19491;
  assign n19493 = ~pi787 & ~n19463;
  assign n19494 = ~n19492 & ~n19493;
  assign n19495 = ~pi644 & ~n19494;
  assign n19496 = ~pi787 & ~n19474;
  assign n19497 = ~n19478 & ~n19488;
  assign n19498 = pi787 & ~n19497;
  assign n19499 = ~n19496 & ~n19498;
  assign n19500 = pi644 & n19499;
  assign n19501 = ~pi715 & ~n19500;
  assign n19502 = ~n19495 & n19501;
  assign n19503 = n17652 & ~n19289;
  assign n19504 = ~n17652 & n19467;
  assign n19505 = ~n19503 & ~n19504;
  assign n19506 = ~pi644 & n19505;
  assign n19507 = pi644 & n19289;
  assign n19508 = pi715 & ~n19507;
  assign n19509 = ~n19506 & n19508;
  assign n19510 = ~pi1160 & ~n19509;
  assign n19511 = ~n19502 & n19510;
  assign n19512 = pi644 & ~n19494;
  assign n19513 = ~pi644 & n19499;
  assign n19514 = pi715 & ~n19513;
  assign n19515 = ~n19512 & n19514;
  assign n19516 = pi644 & n19505;
  assign n19517 = ~pi644 & n19289;
  assign n19518 = ~pi715 & ~n19517;
  assign n19519 = ~n19516 & n19518;
  assign n19520 = pi1160 & ~n19519;
  assign n19521 = ~n19515 & n19520;
  assign n19522 = pi790 & ~n19521;
  assign n19523 = ~n19511 & n19522;
  assign n19524 = ~pi790 & n19494;
  assign n19525 = ~po1038 & ~n19524;
  assign n19526 = ~n19523 & n19525;
  assign n19527 = ~pi143 & po1038;
  assign n19528 = ~pi832 & ~n19527;
  assign n19529 = ~n19526 & n19528;
  assign n19530 = ~pi143 & ~n2754;
  assign n19531 = pi687 & n16786;
  assign n19532 = ~n19530 & ~n19531;
  assign n19533 = ~pi778 & n19532;
  assign n19534 = ~pi625 & n19531;
  assign n19535 = ~n19532 & ~n19534;
  assign n19536 = pi1153 & ~n19535;
  assign n19537 = ~pi1153 & ~n19530;
  assign n19538 = ~n19534 & n19537;
  assign n19539 = ~n19536 & ~n19538;
  assign n19540 = pi778 & ~n19539;
  assign n19541 = ~n19533 & ~n19540;
  assign n19542 = ~n17692 & n19541;
  assign n19543 = ~n17694 & n19542;
  assign n19544 = ~n17696 & n19543;
  assign n19545 = n17704 & n19544;
  assign n19546 = ~pi774 & n16784;
  assign n19547 = ~n19530 & ~n19546;
  assign n19548 = ~n17706 & ~n19547;
  assign n19549 = ~pi785 & ~n19548;
  assign n19550 = ~n17711 & ~n19547;
  assign n19551 = pi1155 & ~n19550;
  assign n19552 = ~n17714 & n19548;
  assign n19553 = ~pi1155 & ~n19552;
  assign n19554 = ~n19551 & ~n19553;
  assign n19555 = pi785 & ~n19554;
  assign n19556 = ~n19549 & ~n19555;
  assign n19557 = ~pi781 & ~n19556;
  assign n19558 = ~n17721 & n19556;
  assign n19559 = pi1154 & ~n19558;
  assign n19560 = ~n17724 & n19556;
  assign n19561 = ~pi1154 & ~n19560;
  assign n19562 = ~n19559 & ~n19561;
  assign n19563 = pi781 & ~n19562;
  assign n19564 = ~n19557 & ~n19563;
  assign n19565 = ~pi789 & ~n19564;
  assign n19566 = pi619 & n19564;
  assign n19567 = ~pi619 & n19530;
  assign n19568 = pi1159 & ~n19567;
  assign n19569 = ~n19566 & n19568;
  assign n19570 = ~pi619 & n19564;
  assign n19571 = pi619 & n19530;
  assign n19572 = ~pi1159 & ~n19571;
  assign n19573 = ~n19570 & n19572;
  assign n19574 = ~n19569 & ~n19573;
  assign n19575 = pi789 & ~n19574;
  assign n19576 = ~n19565 & ~n19575;
  assign n19577 = pi626 & n19576;
  assign n19578 = ~pi626 & n19530;
  assign n19579 = pi1158 & ~n19578;
  assign n19580 = ~n19577 & n19579;
  assign n19581 = ~pi626 & n19576;
  assign n19582 = pi626 & n19530;
  assign n19583 = ~pi1158 & ~n19582;
  assign n19584 = ~n19581 & n19583;
  assign n19585 = ~n19580 & ~n19584;
  assign n19586 = ~n17581 & n19585;
  assign n19587 = ~n19545 & ~n19586;
  assign n19588 = pi788 & ~n19587;
  assign n19589 = ~n16521 & ~n19532;
  assign n19590 = pi625 & n19589;
  assign n19591 = n19547 & ~n19589;
  assign n19592 = ~n19590 & ~n19591;
  assign n19593 = n19537 & ~n19592;
  assign n19594 = ~pi608 & ~n19536;
  assign n19595 = ~n19593 & n19594;
  assign n19596 = pi1153 & n19547;
  assign n19597 = ~n19590 & n19596;
  assign n19598 = pi608 & ~n19538;
  assign n19599 = ~n19597 & n19598;
  assign n19600 = ~n19595 & ~n19599;
  assign n19601 = pi778 & ~n19600;
  assign n19602 = ~pi778 & ~n19591;
  assign n19603 = ~n19601 & ~n19602;
  assign n19604 = ~pi609 & ~n19603;
  assign n19605 = pi609 & n19541;
  assign n19606 = ~pi1155 & ~n19605;
  assign n19607 = ~n19604 & n19606;
  assign n19608 = ~pi660 & ~n19551;
  assign n19609 = ~n19607 & n19608;
  assign n19610 = pi609 & ~n19603;
  assign n19611 = ~pi609 & n19541;
  assign n19612 = pi1155 & ~n19611;
  assign n19613 = ~n19610 & n19612;
  assign n19614 = pi660 & ~n19553;
  assign n19615 = ~n19613 & n19614;
  assign n19616 = ~n19609 & ~n19615;
  assign n19617 = pi785 & ~n19616;
  assign n19618 = ~pi785 & ~n19603;
  assign n19619 = ~n19617 & ~n19618;
  assign n19620 = ~pi618 & ~n19619;
  assign n19621 = pi618 & n19542;
  assign n19622 = ~pi1154 & ~n19621;
  assign n19623 = ~n19620 & n19622;
  assign n19624 = ~pi627 & ~n19559;
  assign n19625 = ~n19623 & n19624;
  assign n19626 = pi618 & ~n19619;
  assign n19627 = ~pi618 & n19542;
  assign n19628 = pi1154 & ~n19627;
  assign n19629 = ~n19626 & n19628;
  assign n19630 = pi627 & ~n19561;
  assign n19631 = ~n19629 & n19630;
  assign n19632 = ~n19625 & ~n19631;
  assign n19633 = pi781 & ~n19632;
  assign n19634 = ~pi781 & ~n19619;
  assign n19635 = ~n19633 & ~n19634;
  assign n19636 = pi619 & ~n19635;
  assign n19637 = ~pi619 & n19543;
  assign n19638 = pi1159 & ~n19637;
  assign n19639 = ~n19636 & n19638;
  assign n19640 = pi648 & ~n19573;
  assign n19641 = ~n19639 & n19640;
  assign n19642 = ~pi619 & ~n19635;
  assign n19643 = pi619 & n19543;
  assign n19644 = ~pi1159 & ~n19643;
  assign n19645 = ~n19642 & n19644;
  assign n19646 = ~pi648 & ~n19569;
  assign n19647 = ~n19645 & n19646;
  assign n19648 = pi789 & ~n19647;
  assign n19649 = ~n19641 & n19648;
  assign n19650 = ~pi789 & n19635;
  assign n19651 = n17817 & ~n19650;
  assign n19652 = ~n19649 & n19651;
  assign n19653 = ~n19588 & ~n19652;
  assign n19654 = ~pi628 & ~n19653;
  assign n19655 = ~pi788 & ~n19576;
  assign n19656 = pi788 & ~n19585;
  assign n19657 = ~n19655 & ~n19656;
  assign n19658 = pi628 & n19657;
  assign n19659 = ~pi1156 & ~n19658;
  assign n19660 = ~n19654 & n19659;
  assign n19661 = ~n17828 & n19544;
  assign n19662 = ~n17830 & n19661;
  assign n19663 = pi1156 & ~n19662;
  assign n19664 = ~pi629 & ~n19663;
  assign n19665 = ~n19660 & n19664;
  assign n19666 = pi628 & ~n19653;
  assign n19667 = ~pi628 & n19657;
  assign n19668 = pi1156 & ~n19667;
  assign n19669 = ~n19666 & n19668;
  assign n19670 = ~n17839 & n19661;
  assign n19671 = ~pi1156 & ~n19670;
  assign n19672 = pi629 & ~n19671;
  assign n19673 = ~n19669 & n19672;
  assign n19674 = ~n19665 & ~n19673;
  assign n19675 = pi792 & ~n19674;
  assign n19676 = ~pi792 & ~n19653;
  assign n19677 = ~n19675 & ~n19676;
  assign n19678 = ~pi647 & ~n19677;
  assign n19679 = ~n17610 & n19657;
  assign n19680 = n17610 & n19530;
  assign n19681 = ~n19679 & ~n19680;
  assign n19682 = pi647 & ~n19681;
  assign n19683 = ~pi1157 & ~n19682;
  assign n19684 = ~n19678 & n19683;
  assign n19685 = ~n17859 & n19661;
  assign n19686 = pi647 & n19685;
  assign n19687 = ~pi647 & n19530;
  assign n19688 = pi1157 & ~n19687;
  assign n19689 = ~n19686 & n19688;
  assign n19690 = ~pi630 & ~n19689;
  assign n19691 = ~n19684 & n19690;
  assign n19692 = pi647 & ~n19677;
  assign n19693 = ~pi647 & ~n19681;
  assign n19694 = pi1157 & ~n19693;
  assign n19695 = ~n19692 & n19694;
  assign n19696 = ~pi647 & n19685;
  assign n19697 = pi647 & n19530;
  assign n19698 = ~pi1157 & ~n19697;
  assign n19699 = ~n19696 & n19698;
  assign n19700 = pi630 & ~n19699;
  assign n19701 = ~n19695 & n19700;
  assign n19702 = ~n19691 & ~n19701;
  assign n19703 = pi787 & ~n19702;
  assign n19704 = ~pi787 & ~n19677;
  assign n19705 = ~n19703 & ~n19704;
  assign n19706 = pi644 & ~n19705;
  assign n19707 = ~pi787 & ~n19685;
  assign n19708 = ~n19689 & ~n19699;
  assign n19709 = pi787 & ~n19708;
  assign n19710 = ~n19707 & ~n19709;
  assign n19711 = ~pi644 & n19710;
  assign n19712 = pi715 & ~n19711;
  assign n19713 = ~n19706 & n19712;
  assign n19714 = n17652 & ~n19530;
  assign n19715 = ~n17652 & n19681;
  assign n19716 = ~n19714 & ~n19715;
  assign n19717 = pi644 & n19716;
  assign n19718 = ~pi644 & n19530;
  assign n19719 = ~pi715 & ~n19718;
  assign n19720 = ~n19717 & n19719;
  assign n19721 = pi1160 & ~n19720;
  assign n19722 = ~n19713 & n19721;
  assign n19723 = ~pi644 & ~n19705;
  assign n19724 = pi644 & n19710;
  assign n19725 = ~pi715 & ~n19724;
  assign n19726 = ~n19723 & n19725;
  assign n19727 = ~pi644 & n19716;
  assign n19728 = pi644 & n19530;
  assign n19729 = pi715 & ~n19728;
  assign n19730 = ~n19727 & n19729;
  assign n19731 = ~pi1160 & ~n19730;
  assign n19732 = ~n19726 & n19731;
  assign n19733 = ~n19722 & ~n19732;
  assign n19734 = pi790 & ~n19733;
  assign n19735 = ~pi790 & ~n19705;
  assign n19736 = pi832 & ~n19735;
  assign n19737 = ~n19734 & n19736;
  assign po300 = ~n19529 & ~n19737;
  assign n19739 = pi144 & ~n3267;
  assign n19740 = pi144 & ~n16687;
  assign n19741 = ~pi144 & ~n16799;
  assign n19742 = ~pi758 & ~n19741;
  assign n19743 = ~n19740 & n19742;
  assign n19744 = ~pi144 & ~n16879;
  assign n19745 = pi144 & n16944;
  assign n19746 = pi758 & ~n19745;
  assign n19747 = ~n19744 & n19746;
  assign n19748 = pi39 & ~n19747;
  assign n19749 = ~n19743 & n19748;
  assign n19750 = pi144 & ~n17088;
  assign n19751 = ~pi144 & ~n17059;
  assign n19752 = ~pi758 & ~n19751;
  assign n19753 = ~n19750 & n19752;
  assign n19754 = pi144 & n17092;
  assign n19755 = ~pi144 & n17094;
  assign n19756 = pi758 & ~n19755;
  assign n19757 = ~n19754 & n19756;
  assign n19758 = ~pi39 & ~n19757;
  assign n19759 = ~n19753 & n19758;
  assign n19760 = ~pi38 & ~n19759;
  assign n19761 = ~n19749 & n19760;
  assign n19762 = pi758 & n16521;
  assign n19763 = n17280 & ~n19762;
  assign n19764 = ~pi144 & ~n17280;
  assign n19765 = pi38 & ~n19764;
  assign n19766 = ~n19763 & n19765;
  assign n19767 = pi736 & ~n19243;
  assign n19768 = ~n19766 & n19767;
  assign n19769 = ~n19761 & n19768;
  assign n19770 = ~pi758 & ~n17199;
  assign n19771 = pi758 & n17240;
  assign n19772 = ~n19770 & ~n19771;
  assign n19773 = pi39 & ~n19772;
  assign n19774 = pi758 & n17042;
  assign n19775 = ~pi758 & n17120;
  assign n19776 = ~pi39 & ~n19775;
  assign n19777 = ~n19774 & n19776;
  assign n19778 = ~n19773 & ~n19777;
  assign n19779 = pi144 & ~n19778;
  assign n19780 = ~pi144 & pi758;
  assign n19781 = n17275 & n19780;
  assign n19782 = ~n19779 & ~n19781;
  assign n19783 = ~pi38 & ~n19782;
  assign n19784 = ~n19766 & ~n19783;
  assign n19785 = n3267 & ~n19784;
  assign n19786 = pi736 & n3267;
  assign n19787 = ~n19785 & ~n19786;
  assign n19788 = ~n19769 & ~n19787;
  assign n19789 = ~n19739 & ~n19788;
  assign n19790 = ~pi625 & n19789;
  assign n19791 = ~n19739 & ~n19785;
  assign n19792 = pi625 & n19791;
  assign n19793 = ~pi1153 & ~n19792;
  assign n19794 = ~n19790 & n19793;
  assign n19795 = pi144 & ~n17406;
  assign n19796 = ~n19786 & ~n19795;
  assign n19797 = pi144 & ~n17972;
  assign n19798 = ~pi144 & n17976;
  assign n19799 = ~pi38 & ~n19798;
  assign n19800 = ~n19797 & n19799;
  assign n19801 = ~n16785 & n17280;
  assign n19802 = pi38 & ~n19801;
  assign n19803 = ~n19764 & n19802;
  assign n19804 = n19786 & ~n19803;
  assign n19805 = ~n19800 & n19804;
  assign n19806 = ~n19796 & ~n19805;
  assign n19807 = pi625 & ~n19806;
  assign n19808 = ~pi625 & ~n19795;
  assign n19809 = pi1153 & ~n19808;
  assign n19810 = ~n19807 & n19809;
  assign n19811 = ~pi608 & ~n19810;
  assign n19812 = ~n19794 & n19811;
  assign n19813 = pi625 & n19789;
  assign n19814 = ~pi625 & n19791;
  assign n19815 = pi1153 & ~n19814;
  assign n19816 = ~n19813 & n19815;
  assign n19817 = ~pi625 & ~n19806;
  assign n19818 = pi625 & ~n19795;
  assign n19819 = ~pi1153 & ~n19818;
  assign n19820 = ~n19817 & n19819;
  assign n19821 = pi608 & ~n19820;
  assign n19822 = ~n19816 & n19821;
  assign n19823 = ~n19812 & ~n19822;
  assign n19824 = pi778 & ~n19823;
  assign n19825 = ~pi778 & n19789;
  assign n19826 = ~n19824 & ~n19825;
  assign n19827 = ~pi609 & ~n19826;
  assign n19828 = ~pi778 & n19806;
  assign n19829 = ~n19810 & ~n19820;
  assign n19830 = pi778 & ~n19829;
  assign n19831 = ~n19828 & ~n19830;
  assign n19832 = pi609 & n19831;
  assign n19833 = ~pi1155 & ~n19832;
  assign n19834 = ~n19827 & n19833;
  assign n19835 = n17438 & ~n19795;
  assign n19836 = ~n17438 & n19791;
  assign n19837 = ~n19835 & ~n19836;
  assign n19838 = pi609 & ~n19837;
  assign n19839 = ~pi609 & ~n19795;
  assign n19840 = pi1155 & ~n19839;
  assign n19841 = ~n19838 & n19840;
  assign n19842 = ~pi660 & ~n19841;
  assign n19843 = ~n19834 & n19842;
  assign n19844 = pi609 & ~n19826;
  assign n19845 = ~pi609 & n19831;
  assign n19846 = pi1155 & ~n19845;
  assign n19847 = ~n19844 & n19846;
  assign n19848 = ~pi609 & ~n19837;
  assign n19849 = pi609 & ~n19795;
  assign n19850 = ~pi1155 & ~n19849;
  assign n19851 = ~n19848 & n19850;
  assign n19852 = pi660 & ~n19851;
  assign n19853 = ~n19847 & n19852;
  assign n19854 = ~n19843 & ~n19853;
  assign n19855 = pi785 & ~n19854;
  assign n19856 = ~pi785 & ~n19826;
  assign n19857 = ~n19855 & ~n19856;
  assign n19858 = ~pi618 & ~n19857;
  assign n19859 = n17466 & ~n19795;
  assign n19860 = ~n17466 & n19831;
  assign n19861 = ~n19859 & ~n19860;
  assign n19862 = pi618 & ~n19861;
  assign n19863 = ~pi1154 & ~n19862;
  assign n19864 = ~n19858 & n19863;
  assign n19865 = ~pi785 & n19837;
  assign n19866 = ~n19841 & ~n19851;
  assign n19867 = pi785 & ~n19866;
  assign n19868 = ~n19865 & ~n19867;
  assign n19869 = pi618 & n19868;
  assign n19870 = ~pi618 & ~n19795;
  assign n19871 = pi1154 & ~n19870;
  assign n19872 = ~n19869 & n19871;
  assign n19873 = ~pi627 & ~n19872;
  assign n19874 = ~n19864 & n19873;
  assign n19875 = pi618 & ~n19857;
  assign n19876 = ~pi618 & ~n19861;
  assign n19877 = pi1154 & ~n19876;
  assign n19878 = ~n19875 & n19877;
  assign n19879 = ~pi618 & n19868;
  assign n19880 = pi618 & ~n19795;
  assign n19881 = ~pi1154 & ~n19880;
  assign n19882 = ~n19879 & n19881;
  assign n19883 = pi627 & ~n19882;
  assign n19884 = ~n19878 & n19883;
  assign n19885 = ~n19874 & ~n19884;
  assign n19886 = pi781 & ~n19885;
  assign n19887 = ~pi781 & ~n19857;
  assign n19888 = ~n19886 & ~n19887;
  assign n19889 = ~pi619 & ~n19888;
  assign n19890 = ~n17503 & n19861;
  assign n19891 = n17503 & n19795;
  assign n19892 = ~n19890 & ~n19891;
  assign n19893 = pi619 & n19892;
  assign n19894 = ~pi1159 & ~n19893;
  assign n19895 = ~n19889 & n19894;
  assign n19896 = ~pi781 & ~n19868;
  assign n19897 = ~n19872 & ~n19882;
  assign n19898 = pi781 & ~n19897;
  assign n19899 = ~n19896 & ~n19898;
  assign n19900 = pi619 & n19899;
  assign n19901 = ~pi619 & ~n19795;
  assign n19902 = pi1159 & ~n19901;
  assign n19903 = ~n19900 & n19902;
  assign n19904 = ~pi648 & ~n19903;
  assign n19905 = ~n19895 & n19904;
  assign n19906 = pi619 & ~n19888;
  assign n19907 = ~pi619 & n19892;
  assign n19908 = pi1159 & ~n19907;
  assign n19909 = ~n19906 & n19908;
  assign n19910 = ~pi619 & n19899;
  assign n19911 = pi619 & ~n19795;
  assign n19912 = ~pi1159 & ~n19911;
  assign n19913 = ~n19910 & n19912;
  assign n19914 = pi648 & ~n19913;
  assign n19915 = ~n19909 & n19914;
  assign n19916 = ~n19905 & ~n19915;
  assign n19917 = pi789 & ~n19916;
  assign n19918 = ~pi789 & ~n19888;
  assign n19919 = ~n19917 & ~n19918;
  assign n19920 = ~pi788 & n19919;
  assign n19921 = ~pi626 & n19919;
  assign n19922 = n17539 & ~n19795;
  assign n19923 = ~n17539 & n19892;
  assign n19924 = ~n19922 & ~n19923;
  assign n19925 = pi626 & n19924;
  assign n19926 = ~pi641 & ~n19925;
  assign n19927 = ~n19921 & n19926;
  assign n19928 = ~pi789 & ~n19899;
  assign n19929 = ~n19903 & ~n19913;
  assign n19930 = pi789 & ~n19929;
  assign n19931 = ~n19928 & ~n19930;
  assign n19932 = ~pi626 & n19931;
  assign n19933 = pi626 & ~n19795;
  assign n19934 = ~pi1158 & ~n19933;
  assign n19935 = ~n19932 & n19934;
  assign n19936 = ~n17546 & ~n19935;
  assign n19937 = ~n19927 & ~n19936;
  assign n19938 = pi626 & n19919;
  assign n19939 = ~pi626 & n19924;
  assign n19940 = pi641 & ~n19939;
  assign n19941 = ~n19938 & n19940;
  assign n19942 = pi626 & n19931;
  assign n19943 = ~pi626 & ~n19795;
  assign n19944 = pi1158 & ~n19943;
  assign n19945 = ~n19942 & n19944;
  assign n19946 = ~n17561 & ~n19945;
  assign n19947 = ~n19941 & ~n19946;
  assign n19948 = ~n19937 & ~n19947;
  assign n19949 = pi788 & ~n19948;
  assign n19950 = ~n19920 & ~n19949;
  assign n19951 = ~pi628 & n19950;
  assign n19952 = ~n19935 & ~n19945;
  assign n19953 = pi788 & ~n19952;
  assign n19954 = ~pi788 & ~n19931;
  assign n19955 = ~n19953 & ~n19954;
  assign n19956 = pi628 & n19955;
  assign n19957 = ~pi1156 & ~n19956;
  assign n19958 = ~n19951 & n19957;
  assign n19959 = ~n17582 & n19924;
  assign n19960 = n17582 & n19795;
  assign n19961 = ~n19959 & ~n19960;
  assign n19962 = pi628 & n19961;
  assign n19963 = ~pi628 & ~n19795;
  assign n19964 = pi1156 & ~n19963;
  assign n19965 = ~n19962 & n19964;
  assign n19966 = ~pi629 & ~n19965;
  assign n19967 = ~n19958 & n19966;
  assign n19968 = pi628 & n19950;
  assign n19969 = ~pi628 & n19955;
  assign n19970 = pi1156 & ~n19969;
  assign n19971 = ~n19968 & n19970;
  assign n19972 = ~pi628 & n19961;
  assign n19973 = pi628 & ~n19795;
  assign n19974 = ~pi1156 & ~n19973;
  assign n19975 = ~n19972 & n19974;
  assign n19976 = pi629 & ~n19975;
  assign n19977 = ~n19971 & n19976;
  assign n19978 = ~n19967 & ~n19977;
  assign n19979 = pi792 & ~n19978;
  assign n19980 = ~pi792 & n19950;
  assign n19981 = ~n19979 & ~n19980;
  assign n19982 = ~pi647 & ~n19981;
  assign n19983 = ~n17610 & ~n19955;
  assign n19984 = n17610 & n19795;
  assign n19985 = ~n19983 & ~n19984;
  assign n19986 = pi647 & n19985;
  assign n19987 = ~pi1157 & ~n19986;
  assign n19988 = ~n19982 & n19987;
  assign n19989 = ~pi792 & ~n19961;
  assign n19990 = ~n19965 & ~n19975;
  assign n19991 = pi792 & ~n19990;
  assign n19992 = ~n19989 & ~n19991;
  assign n19993 = pi647 & n19992;
  assign n19994 = ~pi647 & ~n19795;
  assign n19995 = pi1157 & ~n19994;
  assign n19996 = ~n19993 & n19995;
  assign n19997 = ~pi630 & ~n19996;
  assign n19998 = ~n19988 & n19997;
  assign n19999 = pi647 & ~n19981;
  assign n20000 = ~pi647 & n19985;
  assign n20001 = pi1157 & ~n20000;
  assign n20002 = ~n19999 & n20001;
  assign n20003 = ~pi647 & n19992;
  assign n20004 = pi647 & ~n19795;
  assign n20005 = ~pi1157 & ~n20004;
  assign n20006 = ~n20003 & n20005;
  assign n20007 = pi630 & ~n20006;
  assign n20008 = ~n20002 & n20007;
  assign n20009 = ~n19998 & ~n20008;
  assign n20010 = pi787 & ~n20009;
  assign n20011 = ~pi787 & ~n19981;
  assign n20012 = ~n20010 & ~n20011;
  assign n20013 = ~pi644 & ~n20012;
  assign n20014 = ~pi787 & ~n19992;
  assign n20015 = ~n19996 & ~n20006;
  assign n20016 = pi787 & ~n20015;
  assign n20017 = ~n20014 & ~n20016;
  assign n20018 = pi644 & n20017;
  assign n20019 = ~pi715 & ~n20018;
  assign n20020 = ~n20013 & n20019;
  assign n20021 = n17652 & ~n19795;
  assign n20022 = ~n17652 & n19985;
  assign n20023 = ~n20021 & ~n20022;
  assign n20024 = ~pi644 & ~n20023;
  assign n20025 = pi644 & ~n19795;
  assign n20026 = pi715 & ~n20025;
  assign n20027 = ~n20024 & n20026;
  assign n20028 = ~pi1160 & ~n20027;
  assign n20029 = ~n20020 & n20028;
  assign n20030 = pi644 & ~n20012;
  assign n20031 = ~pi644 & n20017;
  assign n20032 = pi715 & ~n20031;
  assign n20033 = ~n20030 & n20032;
  assign n20034 = pi644 & ~n20023;
  assign n20035 = ~pi644 & ~n19795;
  assign n20036 = ~pi715 & ~n20035;
  assign n20037 = ~n20034 & n20036;
  assign n20038 = pi1160 & ~n20037;
  assign n20039 = ~n20033 & n20038;
  assign n20040 = pi790 & ~n20039;
  assign n20041 = ~n20029 & n20040;
  assign n20042 = ~pi790 & n20012;
  assign n20043 = n6286 & ~n20042;
  assign n20044 = ~n20041 & n20043;
  assign n20045 = ~pi144 & ~n6286;
  assign n20046 = ~pi57 & ~n20045;
  assign n20047 = ~n20044 & n20046;
  assign n20048 = pi57 & pi144;
  assign n20049 = ~pi832 & ~n20048;
  assign n20050 = ~n20047 & n20049;
  assign n20051 = pi144 & ~n2754;
  assign n20052 = pi736 & n16786;
  assign n20053 = ~n20051 & ~n20052;
  assign n20054 = ~pi778 & n20053;
  assign n20055 = pi625 & n20052;
  assign n20056 = ~n20053 & ~n20055;
  assign n20057 = ~pi1153 & ~n20056;
  assign n20058 = pi1153 & ~n20051;
  assign n20059 = ~n20055 & n20058;
  assign n20060 = ~n20057 & ~n20059;
  assign n20061 = pi778 & ~n20060;
  assign n20062 = ~n20054 & ~n20061;
  assign n20063 = n19128 & n20062;
  assign n20064 = ~pi628 & n20063;
  assign n20065 = pi629 & ~n20064;
  assign n20066 = pi609 & pi1155;
  assign n20067 = ~pi609 & ~pi1155;
  assign n20068 = pi785 & ~n20067;
  assign n20069 = ~n20066 & n20068;
  assign n20070 = pi758 & n16784;
  assign n20071 = ~n20069 & n20070;
  assign n20072 = pi618 & pi1154;
  assign n20073 = ~pi618 & ~pi1154;
  assign n20074 = pi781 & ~n20073;
  assign n20075 = ~n20072 & n20074;
  assign n20076 = ~pi619 & pi1159;
  assign n20077 = pi619 & ~pi1159;
  assign n20078 = ~n20076 & ~n20077;
  assign n20079 = pi789 & ~n20078;
  assign n20080 = ~n17438 & ~n20079;
  assign n20081 = ~n20075 & n20080;
  assign n20082 = n20071 & n20081;
  assign n20083 = ~n17816 & n20082;
  assign n20084 = pi628 & ~n20083;
  assign n20085 = ~n20065 & ~n20084;
  assign n20086 = ~pi1156 & ~n20085;
  assign n20087 = pi628 & n20063;
  assign n20088 = ~pi628 & ~n20083;
  assign n20089 = pi629 & ~n20088;
  assign n20090 = pi1156 & ~n20089;
  assign n20091 = ~n20087 & n20090;
  assign n20092 = ~n20086 & ~n20091;
  assign n20093 = ~n20051 & ~n20092;
  assign n20094 = pi792 & n20093;
  assign n20095 = ~n17692 & n20062;
  assign n20096 = ~n17694 & n20095;
  assign n20097 = ~n17696 & n20096;
  assign n20098 = n17699 & n20097;
  assign n20099 = pi626 & n20082;
  assign n20100 = ~n20051 & ~n20099;
  assign n20101 = pi1158 & ~n20100;
  assign n20102 = ~pi641 & ~n20101;
  assign n20103 = ~n20098 & n20102;
  assign n20104 = n17698 & n20097;
  assign n20105 = ~pi626 & n20082;
  assign n20106 = ~n20051 & ~n20105;
  assign n20107 = ~pi1158 & ~n20106;
  assign n20108 = pi641 & ~n20107;
  assign n20109 = ~n20104 & n20108;
  assign n20110 = pi788 & ~n20109;
  assign n20111 = ~n20103 & n20110;
  assign n20112 = ~n20051 & ~n20070;
  assign n20113 = pi736 & n16787;
  assign n20114 = n20112 & ~n20113;
  assign n20115 = pi625 & n20113;
  assign n20116 = ~n20114 & ~n20115;
  assign n20117 = ~pi1153 & ~n20116;
  assign n20118 = ~pi608 & ~n20059;
  assign n20119 = ~n20117 & n20118;
  assign n20120 = pi1153 & n20112;
  assign n20121 = ~n20115 & n20120;
  assign n20122 = pi608 & ~n20057;
  assign n20123 = ~n20121 & n20122;
  assign n20124 = ~n20119 & ~n20123;
  assign n20125 = pi778 & ~n20124;
  assign n20126 = ~pi778 & ~n20114;
  assign n20127 = ~n20125 & ~n20126;
  assign n20128 = ~pi609 & ~n20127;
  assign n20129 = pi609 & n20062;
  assign n20130 = ~pi1155 & ~n20129;
  assign n20131 = ~n20128 & n20130;
  assign n20132 = n17439 & n20070;
  assign n20133 = pi1155 & ~n20051;
  assign n20134 = ~n20132 & n20133;
  assign n20135 = ~pi660 & ~n20134;
  assign n20136 = ~n20131 & n20135;
  assign n20137 = pi609 & ~n20127;
  assign n20138 = ~pi609 & n20062;
  assign n20139 = pi1155 & ~n20138;
  assign n20140 = ~n20137 & n20139;
  assign n20141 = n17451 & n20070;
  assign n20142 = ~pi1155 & ~n20051;
  assign n20143 = ~n20141 & n20142;
  assign n20144 = pi660 & ~n20143;
  assign n20145 = ~n20140 & n20144;
  assign n20146 = ~n20136 & ~n20145;
  assign n20147 = pi785 & ~n20146;
  assign n20148 = ~pi785 & ~n20127;
  assign n20149 = ~n20147 & ~n20148;
  assign n20150 = ~pi618 & ~n20149;
  assign n20151 = pi618 & n20095;
  assign n20152 = ~pi1154 & ~n20151;
  assign n20153 = ~n20150 & n20152;
  assign n20154 = pi618 & ~n17438;
  assign n20155 = n20071 & n20154;
  assign n20156 = pi1154 & ~n20051;
  assign n20157 = ~n20155 & n20156;
  assign n20158 = ~pi627 & ~n20157;
  assign n20159 = ~n20153 & n20158;
  assign n20160 = pi618 & ~n20149;
  assign n20161 = ~pi618 & n20095;
  assign n20162 = pi1154 & ~n20161;
  assign n20163 = ~n20160 & n20162;
  assign n20164 = ~pi618 & ~n17438;
  assign n20165 = n20071 & n20164;
  assign n20166 = ~pi1154 & ~n20051;
  assign n20167 = ~n20165 & n20166;
  assign n20168 = pi627 & ~n20167;
  assign n20169 = ~n20163 & n20168;
  assign n20170 = ~n20159 & ~n20169;
  assign n20171 = pi781 & ~n20170;
  assign n20172 = ~pi781 & ~n20149;
  assign n20173 = ~n20171 & ~n20172;
  assign n20174 = pi619 & ~n20173;
  assign n20175 = ~pi619 & n20096;
  assign n20176 = pi1159 & ~n20175;
  assign n20177 = ~n20174 & n20176;
  assign n20178 = n20071 & ~n20075;
  assign n20179 = ~pi619 & ~n17438;
  assign n20180 = n20178 & n20179;
  assign n20181 = ~pi1159 & ~n20051;
  assign n20182 = ~n20180 & n20181;
  assign n20183 = pi648 & ~n20182;
  assign n20184 = ~n20177 & n20183;
  assign n20185 = ~pi619 & ~n20173;
  assign n20186 = pi619 & n20096;
  assign n20187 = ~pi1159 & ~n20186;
  assign n20188 = ~n20185 & n20187;
  assign n20189 = pi619 & ~n17438;
  assign n20190 = n20178 & n20189;
  assign n20191 = pi1159 & ~n20051;
  assign n20192 = ~n20190 & n20191;
  assign n20193 = ~pi648 & ~n20192;
  assign n20194 = ~n20188 & n20193;
  assign n20195 = pi789 & ~n20194;
  assign n20196 = ~n20184 & n20195;
  assign n20197 = ~pi789 & n20173;
  assign n20198 = n17817 & ~n20197;
  assign n20199 = ~n20196 & n20198;
  assign n20200 = ~n20111 & ~n20199;
  assign n20201 = ~n20094 & ~n20200;
  assign n20202 = ~pi629 & n19155;
  assign n20203 = pi629 & n19156;
  assign n20204 = pi792 & ~n20203;
  assign n20205 = ~n20202 & n20204;
  assign n20206 = ~n20093 & n20205;
  assign n20207 = ~n17652 & ~n19182;
  assign n20208 = ~n20206 & n20207;
  assign n20209 = ~n20201 & n20208;
  assign n20210 = ~n17610 & n20083;
  assign n20211 = ~pi630 & n20210;
  assign n20212 = pi647 & ~n20211;
  assign n20213 = ~n19158 & n20063;
  assign n20214 = pi630 & ~n20213;
  assign n20215 = ~n20212 & ~n20214;
  assign n20216 = ~pi1157 & ~n20215;
  assign n20217 = ~pi630 & ~n20213;
  assign n20218 = pi647 & ~n20217;
  assign n20219 = pi630 & n20210;
  assign n20220 = pi1157 & ~n20219;
  assign n20221 = ~n20218 & n20220;
  assign n20222 = ~n20216 & ~n20221;
  assign n20223 = pi787 & ~n20051;
  assign n20224 = ~n20222 & n20223;
  assign n20225 = ~n20209 & ~n20224;
  assign n20226 = pi644 & n20225;
  assign n20227 = ~n19182 & n20213;
  assign n20228 = ~n20051 & ~n20227;
  assign n20229 = ~pi644 & ~n20228;
  assign n20230 = pi715 & ~n20229;
  assign n20231 = ~n20226 & n20230;
  assign n20232 = ~n17652 & n20210;
  assign n20233 = pi644 & n20232;
  assign n20234 = ~pi715 & ~n20051;
  assign n20235 = ~n20233 & n20234;
  assign n20236 = pi1160 & ~n20235;
  assign n20237 = ~n20231 & n20236;
  assign n20238 = ~pi644 & n20225;
  assign n20239 = pi644 & ~n20228;
  assign n20240 = ~pi715 & ~n20239;
  assign n20241 = ~n20238 & n20240;
  assign n20242 = ~pi644 & n20232;
  assign n20243 = pi715 & ~n20051;
  assign n20244 = ~n20242 & n20243;
  assign n20245 = ~pi1160 & ~n20244;
  assign n20246 = ~n20241 & n20245;
  assign n20247 = ~n20237 & ~n20246;
  assign n20248 = pi790 & ~n20247;
  assign n20249 = ~pi790 & n20225;
  assign n20250 = pi832 & ~n20249;
  assign n20251 = ~n20248 & n20250;
  assign po301 = ~n20050 & ~n20251;
  assign n20253 = ~pi145 & ~n17406;
  assign n20254 = n17539 & ~n20253;
  assign n20255 = ~pi698 & n3267;
  assign n20256 = n20253 & ~n20255;
  assign n20257 = pi145 & ~n17976;
  assign n20258 = ~pi38 & ~n20257;
  assign n20259 = n3267 & ~n20258;
  assign n20260 = ~pi145 & n17972;
  assign n20261 = ~n20259 & ~n20260;
  assign n20262 = ~pi145 & ~n17280;
  assign n20263 = n17392 & ~n20262;
  assign n20264 = ~pi698 & ~n20263;
  assign n20265 = ~n20261 & n20264;
  assign n20266 = ~n20256 & ~n20265;
  assign n20267 = ~pi778 & n20266;
  assign n20268 = pi625 & ~n20266;
  assign n20269 = ~pi625 & n20253;
  assign n20270 = pi1153 & ~n20269;
  assign n20271 = ~n20268 & n20270;
  assign n20272 = ~pi625 & ~n20266;
  assign n20273 = pi625 & n20253;
  assign n20274 = ~pi1153 & ~n20273;
  assign n20275 = ~n20272 & n20274;
  assign n20276 = ~n20271 & ~n20275;
  assign n20277 = pi778 & ~n20276;
  assign n20278 = ~n20267 & ~n20277;
  assign n20279 = ~n17466 & ~n20278;
  assign n20280 = n17466 & ~n20253;
  assign n20281 = ~n20279 & ~n20280;
  assign n20282 = ~n17503 & n20281;
  assign n20283 = n17503 & n20253;
  assign n20284 = ~n20282 & ~n20283;
  assign n20285 = ~n17539 & n20284;
  assign n20286 = ~n20254 & ~n20285;
  assign n20287 = ~n17582 & n20286;
  assign n20288 = n17582 & n20253;
  assign n20289 = ~n20287 & ~n20288;
  assign n20290 = ~pi792 & n20289;
  assign n20291 = pi628 & ~n20289;
  assign n20292 = ~pi628 & n20253;
  assign n20293 = pi1156 & ~n20292;
  assign n20294 = ~n20291 & n20293;
  assign n20295 = ~pi628 & ~n20289;
  assign n20296 = pi628 & n20253;
  assign n20297 = ~pi1156 & ~n20296;
  assign n20298 = ~n20295 & n20297;
  assign n20299 = ~n20294 & ~n20298;
  assign n20300 = pi792 & ~n20299;
  assign n20301 = ~n20290 & ~n20300;
  assign n20302 = ~pi647 & ~n20301;
  assign n20303 = pi647 & ~n20253;
  assign n20304 = ~n20302 & ~n20303;
  assign n20305 = ~pi1157 & n20304;
  assign n20306 = pi647 & ~n20301;
  assign n20307 = ~pi647 & ~n20253;
  assign n20308 = ~n20306 & ~n20307;
  assign n20309 = pi1157 & n20308;
  assign n20310 = ~n20305 & ~n20309;
  assign n20311 = pi787 & ~n20310;
  assign n20312 = ~pi787 & n20301;
  assign n20313 = ~n20311 & ~n20312;
  assign n20314 = ~pi644 & ~n20313;
  assign n20315 = pi715 & ~n20314;
  assign n20316 = pi145 & ~n3267;
  assign n20317 = ~pi145 & ~n17201;
  assign n20318 = pi767 & ~n20317;
  assign n20319 = pi145 & ~n17275;
  assign n20320 = ~pi145 & ~pi767;
  assign n20321 = n17242 & n20320;
  assign n20322 = ~n20319 & ~n20321;
  assign n20323 = ~n20318 & n20322;
  assign n20324 = ~pi38 & ~n20323;
  assign n20325 = ~pi767 & n17282;
  assign n20326 = pi38 & ~n20262;
  assign n20327 = ~n20325 & n20326;
  assign n20328 = ~n20324 & ~n20327;
  assign n20329 = n3267 & ~n20328;
  assign n20330 = ~n20316 & ~n20329;
  assign n20331 = ~n17438 & ~n20330;
  assign n20332 = n17438 & ~n20253;
  assign n20333 = ~n20331 & ~n20332;
  assign n20334 = ~pi785 & ~n20333;
  assign n20335 = ~n17439 & ~n20253;
  assign n20336 = pi609 & n20331;
  assign n20337 = ~n20335 & ~n20336;
  assign n20338 = pi1155 & ~n20337;
  assign n20339 = ~n17451 & ~n20253;
  assign n20340 = ~pi609 & n20331;
  assign n20341 = ~n20339 & ~n20340;
  assign n20342 = ~pi1155 & ~n20341;
  assign n20343 = ~n20338 & ~n20342;
  assign n20344 = pi785 & ~n20343;
  assign n20345 = ~n20334 & ~n20344;
  assign n20346 = ~pi781 & ~n20345;
  assign n20347 = pi618 & n20345;
  assign n20348 = ~pi618 & n20253;
  assign n20349 = pi1154 & ~n20348;
  assign n20350 = ~n20347 & n20349;
  assign n20351 = ~pi618 & n20345;
  assign n20352 = pi618 & n20253;
  assign n20353 = ~pi1154 & ~n20352;
  assign n20354 = ~n20351 & n20353;
  assign n20355 = ~n20350 & ~n20354;
  assign n20356 = pi781 & ~n20355;
  assign n20357 = ~n20346 & ~n20356;
  assign n20358 = ~pi789 & ~n20357;
  assign n20359 = pi619 & n20357;
  assign n20360 = ~pi619 & n20253;
  assign n20361 = pi1159 & ~n20360;
  assign n20362 = ~n20359 & n20361;
  assign n20363 = ~pi619 & n20357;
  assign n20364 = pi619 & n20253;
  assign n20365 = ~pi1159 & ~n20364;
  assign n20366 = ~n20363 & n20365;
  assign n20367 = ~n20362 & ~n20366;
  assign n20368 = pi789 & ~n20367;
  assign n20369 = ~n20358 & ~n20368;
  assign n20370 = ~pi788 & ~n20369;
  assign n20371 = pi626 & n20369;
  assign n20372 = ~pi626 & n20253;
  assign n20373 = pi1158 & ~n20372;
  assign n20374 = ~n20371 & n20373;
  assign n20375 = ~pi626 & n20369;
  assign n20376 = pi626 & n20253;
  assign n20377 = ~pi1158 & ~n20376;
  assign n20378 = ~n20375 & n20377;
  assign n20379 = ~n20374 & ~n20378;
  assign n20380 = pi788 & ~n20379;
  assign n20381 = ~n20370 & ~n20380;
  assign n20382 = ~n17610 & n20381;
  assign n20383 = n17610 & n20253;
  assign n20384 = ~n20382 & ~n20383;
  assign n20385 = ~n17652 & ~n20384;
  assign n20386 = n17652 & n20253;
  assign n20387 = ~n20385 & ~n20386;
  assign n20388 = pi644 & ~n20387;
  assign n20389 = ~pi644 & n20253;
  assign n20390 = ~pi715 & ~n20389;
  assign n20391 = ~n20388 & n20390;
  assign n20392 = pi1160 & ~n20391;
  assign n20393 = ~n20315 & n20392;
  assign n20394 = pi630 & ~pi647;
  assign n20395 = pi1157 & n20394;
  assign n20396 = ~pi630 & pi647;
  assign n20397 = ~pi1157 & n20396;
  assign n20398 = ~n20395 & ~n20397;
  assign n20399 = n20384 & ~n20398;
  assign n20400 = n17650 & ~n20304;
  assign n20401 = n17649 & ~n20308;
  assign n20402 = ~n20400 & ~n20401;
  assign n20403 = ~n20399 & n20402;
  assign n20404 = pi787 & ~n20403;
  assign n20405 = ~pi628 & pi629;
  assign n20406 = pi1156 & n20405;
  assign n20407 = pi628 & ~pi629;
  assign n20408 = ~pi1156 & n20407;
  assign n20409 = ~n20406 & ~n20408;
  assign n20410 = ~n20381 & ~n20409;
  assign n20411 = ~pi629 & n20294;
  assign n20412 = pi629 & n20298;
  assign n20413 = ~n20411 & ~n20412;
  assign n20414 = ~n20410 & n20413;
  assign n20415 = pi792 & ~n20414;
  assign n20416 = pi698 & n20328;
  assign n20417 = ~pi145 & n16687;
  assign n20418 = pi145 & n16799;
  assign n20419 = pi767 & ~n20418;
  assign n20420 = ~n20417 & n20419;
  assign n20421 = pi145 & n16879;
  assign n20422 = ~pi145 & ~n16944;
  assign n20423 = ~pi767 & ~n20422;
  assign n20424 = ~n20421 & n20423;
  assign n20425 = pi39 & ~n20424;
  assign n20426 = ~n20420 & n20425;
  assign n20427 = ~pi145 & ~n17088;
  assign n20428 = pi145 & ~n17059;
  assign n20429 = pi767 & ~n20428;
  assign n20430 = ~n20427 & n20429;
  assign n20431 = ~pi145 & n17092;
  assign n20432 = pi145 & n17094;
  assign n20433 = ~pi767 & ~n20432;
  assign n20434 = ~n20431 & n20433;
  assign n20435 = ~n20430 & ~n20434;
  assign n20436 = ~pi39 & ~n20435;
  assign n20437 = ~pi38 & ~n20436;
  assign n20438 = ~n20426 & n20437;
  assign n20439 = ~pi767 & ~n16905;
  assign n20440 = n19230 & ~n20439;
  assign n20441 = ~pi145 & ~n20440;
  assign n20442 = ~pi767 & n16784;
  assign n20443 = ~n16787 & ~n20442;
  assign n20444 = pi145 & ~n20443;
  assign n20445 = n6234 & n20444;
  assign n20446 = pi38 & ~n20445;
  assign n20447 = ~n20441 & n20446;
  assign n20448 = ~pi698 & ~n20447;
  assign n20449 = ~n20438 & n20448;
  assign n20450 = n3267 & ~n20449;
  assign n20451 = ~n20416 & n20450;
  assign n20452 = ~n20316 & ~n20451;
  assign n20453 = ~pi625 & n20452;
  assign n20454 = pi625 & n20330;
  assign n20455 = ~pi1153 & ~n20454;
  assign n20456 = ~n20453 & n20455;
  assign n20457 = ~pi608 & ~n20271;
  assign n20458 = ~n20456 & n20457;
  assign n20459 = pi625 & n20452;
  assign n20460 = ~pi625 & n20330;
  assign n20461 = pi1153 & ~n20460;
  assign n20462 = ~n20459 & n20461;
  assign n20463 = pi608 & ~n20275;
  assign n20464 = ~n20462 & n20463;
  assign n20465 = ~n20458 & ~n20464;
  assign n20466 = pi778 & ~n20465;
  assign n20467 = ~pi778 & n20452;
  assign n20468 = ~n20466 & ~n20467;
  assign n20469 = ~pi609 & ~n20468;
  assign n20470 = pi609 & n20278;
  assign n20471 = ~pi1155 & ~n20470;
  assign n20472 = ~n20469 & n20471;
  assign n20473 = ~pi660 & ~n20338;
  assign n20474 = ~n20472 & n20473;
  assign n20475 = pi609 & ~n20468;
  assign n20476 = ~pi609 & n20278;
  assign n20477 = pi1155 & ~n20476;
  assign n20478 = ~n20475 & n20477;
  assign n20479 = pi660 & ~n20342;
  assign n20480 = ~n20478 & n20479;
  assign n20481 = ~n20474 & ~n20480;
  assign n20482 = pi785 & ~n20481;
  assign n20483 = ~pi785 & ~n20468;
  assign n20484 = ~n20482 & ~n20483;
  assign n20485 = ~pi618 & ~n20484;
  assign n20486 = pi618 & n20281;
  assign n20487 = ~pi1154 & ~n20486;
  assign n20488 = ~n20485 & n20487;
  assign n20489 = ~pi627 & ~n20350;
  assign n20490 = ~n20488 & n20489;
  assign n20491 = pi618 & ~n20484;
  assign n20492 = ~pi618 & n20281;
  assign n20493 = pi1154 & ~n20492;
  assign n20494 = ~n20491 & n20493;
  assign n20495 = pi627 & ~n20354;
  assign n20496 = ~n20494 & n20495;
  assign n20497 = ~n20490 & ~n20496;
  assign n20498 = pi781 & ~n20497;
  assign n20499 = ~pi781 & ~n20484;
  assign n20500 = ~n20498 & ~n20499;
  assign n20501 = pi619 & ~n20500;
  assign n20502 = ~pi619 & ~n20284;
  assign n20503 = pi1159 & ~n20502;
  assign n20504 = ~n20501 & n20503;
  assign n20505 = pi648 & ~n20366;
  assign n20506 = ~n20504 & n20505;
  assign n20507 = ~pi619 & ~n20500;
  assign n20508 = pi619 & ~n20284;
  assign n20509 = ~pi1159 & ~n20508;
  assign n20510 = ~n20507 & n20509;
  assign n20511 = ~pi648 & ~n20362;
  assign n20512 = ~n20510 & n20511;
  assign n20513 = pi789 & ~n20512;
  assign n20514 = ~n20506 & n20513;
  assign n20515 = ~pi789 & n20500;
  assign n20516 = n17817 & ~n20515;
  assign n20517 = ~n20514 & n20516;
  assign n20518 = n17704 & n20286;
  assign n20519 = ~n17581 & n20379;
  assign n20520 = ~n20518 & ~n20519;
  assign n20521 = pi788 & ~n20520;
  assign n20522 = ~n20205 & ~n20521;
  assign n20523 = ~n20517 & n20522;
  assign n20524 = ~n20415 & ~n20523;
  assign n20525 = n20207 & ~n20524;
  assign n20526 = ~n20404 & ~n20525;
  assign n20527 = ~pi644 & n20526;
  assign n20528 = pi644 & ~n20313;
  assign n20529 = ~pi715 & ~n20528;
  assign n20530 = ~n20527 & n20529;
  assign n20531 = ~pi644 & ~n20387;
  assign n20532 = pi644 & n20253;
  assign n20533 = pi715 & ~n20532;
  assign n20534 = ~n20531 & n20533;
  assign n20535 = ~pi1160 & ~n20534;
  assign n20536 = ~n20530 & n20535;
  assign n20537 = ~n20393 & ~n20536;
  assign n20538 = pi790 & ~n20537;
  assign n20539 = pi644 & n20392;
  assign n20540 = pi790 & ~n20539;
  assign n20541 = n20526 & ~n20540;
  assign n20542 = ~n20538 & ~n20541;
  assign n20543 = ~po1038 & ~n20542;
  assign n20544 = ~pi145 & po1038;
  assign n20545 = ~pi832 & ~n20544;
  assign n20546 = ~n20543 & n20545;
  assign n20547 = ~pi145 & ~n2754;
  assign n20548 = ~n20442 & ~n20547;
  assign n20549 = ~n17706 & ~n20548;
  assign n20550 = ~pi785 & ~n20549;
  assign n20551 = ~n17711 & ~n20548;
  assign n20552 = pi1155 & ~n20551;
  assign n20553 = ~n17714 & n20549;
  assign n20554 = ~pi1155 & ~n20553;
  assign n20555 = ~n20552 & ~n20554;
  assign n20556 = pi785 & ~n20555;
  assign n20557 = ~n20550 & ~n20556;
  assign n20558 = ~pi781 & ~n20557;
  assign n20559 = ~n17721 & n20557;
  assign n20560 = pi1154 & ~n20559;
  assign n20561 = ~n17724 & n20557;
  assign n20562 = ~pi1154 & ~n20561;
  assign n20563 = ~n20560 & ~n20562;
  assign n20564 = pi781 & ~n20563;
  assign n20565 = ~n20558 & ~n20564;
  assign n20566 = ~pi789 & ~n20565;
  assign n20567 = pi619 & n20565;
  assign n20568 = ~pi619 & n20547;
  assign n20569 = pi1159 & ~n20568;
  assign n20570 = ~n20567 & n20569;
  assign n20571 = ~pi619 & n20565;
  assign n20572 = pi619 & n20547;
  assign n20573 = ~pi1159 & ~n20572;
  assign n20574 = ~n20571 & n20573;
  assign n20575 = ~n20570 & ~n20574;
  assign n20576 = pi789 & ~n20575;
  assign n20577 = ~n20566 & ~n20576;
  assign n20578 = ~pi788 & ~n20577;
  assign n20579 = pi626 & n20577;
  assign n20580 = ~pi626 & n20547;
  assign n20581 = pi1158 & ~n20580;
  assign n20582 = ~n20579 & n20581;
  assign n20583 = ~pi626 & n20577;
  assign n20584 = pi626 & n20547;
  assign n20585 = ~pi1158 & ~n20584;
  assign n20586 = ~n20583 & n20585;
  assign n20587 = ~n20582 & ~n20586;
  assign n20588 = pi788 & ~n20587;
  assign n20589 = ~n20578 & ~n20588;
  assign n20590 = ~n17610 & n20589;
  assign n20591 = n17610 & n20547;
  assign n20592 = ~n20590 & ~n20591;
  assign n20593 = ~n20398 & n20592;
  assign n20594 = ~pi698 & n16786;
  assign n20595 = ~n20547 & ~n20594;
  assign n20596 = ~pi778 & n20595;
  assign n20597 = ~pi625 & n20594;
  assign n20598 = ~n20595 & ~n20597;
  assign n20599 = pi1153 & ~n20598;
  assign n20600 = ~pi1153 & ~n20547;
  assign n20601 = ~n20597 & n20600;
  assign n20602 = ~n20599 & ~n20601;
  assign n20603 = pi778 & ~n20602;
  assign n20604 = ~n20596 & ~n20603;
  assign n20605 = ~n17692 & n20604;
  assign n20606 = ~n17694 & n20605;
  assign n20607 = ~n17696 & n20606;
  assign n20608 = ~n17828 & n20607;
  assign n20609 = ~n17859 & n20608;
  assign n20610 = ~pi647 & n20609;
  assign n20611 = pi647 & n20547;
  assign n20612 = ~pi1157 & ~n20611;
  assign n20613 = ~n20610 & n20612;
  assign n20614 = pi647 & ~n20609;
  assign n20615 = ~pi647 & ~n20547;
  assign n20616 = ~n20614 & ~n20615;
  assign n20617 = pi1157 & ~n20616;
  assign n20618 = ~n20613 & ~n20617;
  assign n20619 = ~n17651 & ~n20618;
  assign n20620 = ~n20593 & ~n20619;
  assign n20621 = pi787 & ~n20620;
  assign n20622 = n17704 & n20607;
  assign n20623 = ~n17581 & n20587;
  assign n20624 = ~n20622 & ~n20623;
  assign n20625 = pi788 & ~n20624;
  assign n20626 = ~n16521 & ~n20595;
  assign n20627 = pi625 & n20626;
  assign n20628 = n20548 & ~n20626;
  assign n20629 = ~n20627 & ~n20628;
  assign n20630 = n20600 & ~n20629;
  assign n20631 = ~pi608 & ~n20599;
  assign n20632 = ~n20630 & n20631;
  assign n20633 = pi1153 & n20548;
  assign n20634 = ~n20627 & n20633;
  assign n20635 = pi608 & ~n20601;
  assign n20636 = ~n20634 & n20635;
  assign n20637 = ~n20632 & ~n20636;
  assign n20638 = pi778 & ~n20637;
  assign n20639 = ~pi778 & ~n20628;
  assign n20640 = ~n20638 & ~n20639;
  assign n20641 = ~pi609 & ~n20640;
  assign n20642 = pi609 & n20604;
  assign n20643 = ~pi1155 & ~n20642;
  assign n20644 = ~n20641 & n20643;
  assign n20645 = ~pi660 & ~n20552;
  assign n20646 = ~n20644 & n20645;
  assign n20647 = pi609 & ~n20640;
  assign n20648 = ~pi609 & n20604;
  assign n20649 = pi1155 & ~n20648;
  assign n20650 = ~n20647 & n20649;
  assign n20651 = pi660 & ~n20554;
  assign n20652 = ~n20650 & n20651;
  assign n20653 = ~n20646 & ~n20652;
  assign n20654 = pi785 & ~n20653;
  assign n20655 = ~pi785 & ~n20640;
  assign n20656 = ~n20654 & ~n20655;
  assign n20657 = ~pi618 & ~n20656;
  assign n20658 = pi618 & n20605;
  assign n20659 = ~pi1154 & ~n20658;
  assign n20660 = ~n20657 & n20659;
  assign n20661 = ~pi627 & ~n20560;
  assign n20662 = ~n20660 & n20661;
  assign n20663 = pi618 & ~n20656;
  assign n20664 = ~pi618 & n20605;
  assign n20665 = pi1154 & ~n20664;
  assign n20666 = ~n20663 & n20665;
  assign n20667 = pi627 & ~n20562;
  assign n20668 = ~n20666 & n20667;
  assign n20669 = ~n20662 & ~n20668;
  assign n20670 = pi781 & ~n20669;
  assign n20671 = ~pi781 & ~n20656;
  assign n20672 = ~n20670 & ~n20671;
  assign n20673 = pi619 & ~n20672;
  assign n20674 = ~pi619 & n20606;
  assign n20675 = pi1159 & ~n20674;
  assign n20676 = ~n20673 & n20675;
  assign n20677 = pi648 & ~n20574;
  assign n20678 = ~n20676 & n20677;
  assign n20679 = ~pi619 & ~n20672;
  assign n20680 = pi619 & n20606;
  assign n20681 = ~pi1159 & ~n20680;
  assign n20682 = ~n20679 & n20681;
  assign n20683 = ~pi648 & ~n20570;
  assign n20684 = ~n20682 & n20683;
  assign n20685 = pi789 & ~n20684;
  assign n20686 = ~n20678 & n20685;
  assign n20687 = ~pi789 & n20672;
  assign n20688 = n17817 & ~n20687;
  assign n20689 = ~n20686 & n20688;
  assign n20690 = ~n20625 & ~n20689;
  assign n20691 = ~n20205 & ~n20690;
  assign n20692 = n17856 & n20589;
  assign n20693 = pi1156 & ~n17830;
  assign n20694 = n20608 & n20693;
  assign n20695 = ~n20692 & ~n20694;
  assign n20696 = ~pi629 & ~n20695;
  assign n20697 = ~pi1156 & ~n17839;
  assign n20698 = n20608 & n20697;
  assign n20699 = n17855 & n20589;
  assign n20700 = ~n20698 & ~n20699;
  assign n20701 = pi629 & ~n20700;
  assign n20702 = ~n20696 & ~n20701;
  assign n20703 = pi792 & ~n20702;
  assign n20704 = n20207 & ~n20703;
  assign n20705 = ~n20691 & n20704;
  assign n20706 = ~n20621 & ~n20705;
  assign n20707 = pi644 & n20706;
  assign n20708 = ~pi787 & ~n20609;
  assign n20709 = pi787 & ~n20618;
  assign n20710 = ~n20708 & ~n20709;
  assign n20711 = ~pi644 & n20710;
  assign n20712 = pi715 & ~n20711;
  assign n20713 = ~n20707 & n20712;
  assign n20714 = ~n17652 & ~n20592;
  assign n20715 = n17652 & n20547;
  assign n20716 = ~n20714 & ~n20715;
  assign n20717 = pi644 & ~n20716;
  assign n20718 = ~pi644 & n20547;
  assign n20719 = ~pi715 & ~n20718;
  assign n20720 = ~n20717 & n20719;
  assign n20721 = pi1160 & ~n20720;
  assign n20722 = ~n20713 & n20721;
  assign n20723 = ~pi644 & n20706;
  assign n20724 = pi644 & n20710;
  assign n20725 = ~pi715 & ~n20724;
  assign n20726 = ~n20723 & n20725;
  assign n20727 = ~pi644 & ~n20716;
  assign n20728 = pi644 & n20547;
  assign n20729 = pi715 & ~n20728;
  assign n20730 = ~n20727 & n20729;
  assign n20731 = ~pi1160 & ~n20730;
  assign n20732 = ~n20726 & n20731;
  assign n20733 = ~n20722 & ~n20732;
  assign n20734 = pi790 & ~n20733;
  assign n20735 = ~pi790 & n20706;
  assign n20736 = pi832 & ~n20735;
  assign n20737 = ~n20734 & n20736;
  assign po302 = ~n20546 & ~n20737;
  assign n20739 = ~pi907 & n6188;
  assign n20740 = pi146 & ~n16812;
  assign n20741 = ~n20739 & n20740;
  assign n20742 = pi146 & ~n17172;
  assign n20743 = n20739 & n20742;
  assign n20744 = pi735 & pi907;
  assign n20745 = n16812 & n20744;
  assign n20746 = ~pi947 & ~n20745;
  assign n20747 = ~n20743 & n20746;
  assign n20748 = pi743 & n16812;
  assign n20749 = pi947 & ~n20740;
  assign n20750 = ~n20748 & n20749;
  assign n20751 = ~n20747 & ~n20750;
  assign n20752 = ~n20741 & ~n20751;
  assign n20753 = ~n3329 & ~n20752;
  assign n20754 = pi743 & pi947;
  assign n20755 = pi907 & ~pi947;
  assign n20756 = pi735 & n20755;
  assign n20757 = ~n20754 & ~n20756;
  assign n20758 = n16518 & ~n20757;
  assign n20759 = pi146 & ~n16518;
  assign n20760 = ~n20758 & ~n20759;
  assign n20761 = n3329 & ~n20760;
  assign n20762 = ~pi215 & ~n20761;
  assign n20763 = ~n20753 & n20762;
  assign n20764 = pi146 & n17195;
  assign n20765 = n17132 & ~n20757;
  assign n20766 = pi215 & ~n20765;
  assign n20767 = ~n20764 & n20766;
  assign n20768 = ~n20763 & ~n20767;
  assign n20769 = pi299 & ~n20768;
  assign n20770 = n16812 & ~n20757;
  assign n20771 = ~n6215 & ~n20740;
  assign n20772 = ~n20770 & n20771;
  assign n20773 = n17172 & ~n20757;
  assign n20774 = n6215 & ~n20742;
  assign n20775 = ~n20773 & n20774;
  assign n20776 = ~n20772 & ~n20775;
  assign n20777 = ~n3052 & ~n20776;
  assign n20778 = n3052 & n20760;
  assign n20779 = ~pi223 & ~n20778;
  assign n20780 = ~n20777 & n20779;
  assign n20781 = pi146 & ~n17132;
  assign n20782 = ~n20765 & ~n20781;
  assign n20783 = ~n6215 & ~n20782;
  assign n20784 = n17151 & n20757;
  assign n20785 = ~pi146 & ~n17151;
  assign n20786 = n6215 & ~n20785;
  assign n20787 = ~n20784 & n20786;
  assign n20788 = ~n20783 & ~n20787;
  assign n20789 = pi223 & ~n20788;
  assign n20790 = ~pi299 & ~n20789;
  assign n20791 = ~n20780 & n20790;
  assign n20792 = ~n20769 & ~n20791;
  assign n20793 = pi39 & ~n20792;
  assign n20794 = n17063 & n20757;
  assign n20795 = ~pi146 & ~n17063;
  assign n20796 = ~pi299 & ~n20795;
  assign n20797 = ~n20794 & n20796;
  assign n20798 = n17026 & n20757;
  assign n20799 = ~pi146 & ~n17026;
  assign n20800 = pi299 & ~n20799;
  assign n20801 = ~n20798 & n20800;
  assign n20802 = ~pi39 & ~n20801;
  assign n20803 = ~n20797 & n20802;
  assign n20804 = ~pi38 & ~n20803;
  assign n20805 = ~n20793 & n20804;
  assign n20806 = ~pi146 & ~n17280;
  assign n20807 = n2754 & n20757;
  assign n20808 = n6234 & n20807;
  assign n20809 = pi38 & ~n20808;
  assign n20810 = ~n20806 & n20809;
  assign n20811 = n10143 & ~n20810;
  assign n20812 = ~n20805 & n20811;
  assign n20813 = ~pi146 & ~n10143;
  assign n20814 = ~pi832 & ~n20813;
  assign n20815 = ~n20812 & n20814;
  assign n20816 = ~pi146 & ~n2754;
  assign n20817 = pi832 & ~n20816;
  assign n20818 = ~n20807 & n20817;
  assign po303 = n20815 | n20818;
  assign n20820 = ~pi770 & pi947;
  assign n20821 = pi726 & n20755;
  assign n20822 = ~n20820 & ~n20821;
  assign n20823 = n2754 & ~n20822;
  assign n20824 = ~pi147 & ~n2754;
  assign n20825 = pi832 & ~n20824;
  assign n20826 = ~n20823 & n20825;
  assign n20827 = ~pi947 & n17120;
  assign n20828 = ~pi39 & ~n20827;
  assign n20829 = ~pi299 & n17179;
  assign n20830 = pi947 & n20829;
  assign n20831 = ~pi947 & n16736;
  assign n20832 = n16812 & n20755;
  assign n20833 = ~n17184 & ~n20832;
  assign n20834 = ~n3329 & ~n20833;
  assign n20835 = ~pi215 & ~n20834;
  assign n20836 = ~n20831 & n20835;
  assign n20837 = pi215 & ~n17194;
  assign n20838 = n17132 & n20755;
  assign n20839 = n20837 & ~n20838;
  assign n20840 = ~n20836 & ~n20839;
  assign n20841 = pi299 & ~n20840;
  assign n20842 = ~n17180 & ~n20841;
  assign n20843 = ~n20830 & n20842;
  assign n20844 = pi39 & ~n20843;
  assign n20845 = ~n20828 & ~n20844;
  assign n20846 = ~pi38 & n20845;
  assign n20847 = pi38 & ~pi947;
  assign n20848 = n17397 & n20847;
  assign n20849 = ~n20846 & ~n20848;
  assign n20850 = ~pi770 & n20849;
  assign n20851 = pi770 & ~n17399;
  assign n20852 = ~n20850 & ~n20851;
  assign n20853 = ~pi147 & ~n20852;
  assign n20854 = ~n17398 & ~n20848;
  assign n20855 = pi947 & n17120;
  assign n20856 = ~pi39 & ~n20855;
  assign n20857 = pi947 & n17179;
  assign n20858 = ~pi299 & ~n20857;
  assign n20859 = pi215 & pi947;
  assign n20860 = n17132 & n20859;
  assign n20861 = pi299 & ~n20860;
  assign n20862 = pi947 & n16812;
  assign n20863 = ~n3329 & ~n20862;
  assign n20864 = pi947 & n16518;
  assign n20865 = n3329 & ~n20864;
  assign n20866 = ~pi215 & ~n20865;
  assign n20867 = ~n20863 & n20866;
  assign n20868 = n20861 & ~n20867;
  assign n20869 = ~n20858 & ~n20868;
  assign n20870 = pi39 & ~n20869;
  assign n20871 = ~n20856 & ~n20870;
  assign n20872 = ~pi38 & ~n20871;
  assign n20873 = n20854 & ~n20872;
  assign n20874 = pi147 & ~pi770;
  assign n20875 = n20873 & n20874;
  assign n20876 = ~pi726 & ~n20875;
  assign n20877 = ~n20853 & n20876;
  assign n20878 = n16736 & ~n20755;
  assign n20879 = ~n17184 & ~n20862;
  assign n20880 = ~n3329 & ~n20879;
  assign n20881 = ~pi215 & ~n20880;
  assign n20882 = ~n20878 & n20881;
  assign n20883 = ~n20837 & ~n20882;
  assign n20884 = ~n20860 & ~n20883;
  assign n20885 = pi299 & ~n20884;
  assign n20886 = ~n20755 & n20829;
  assign n20887 = ~n20885 & ~n20886;
  assign n20888 = pi39 & ~n20887;
  assign n20889 = n17120 & ~n20755;
  assign n20890 = ~pi39 & n20889;
  assign n20891 = ~n20888 & ~n20890;
  assign n20892 = ~pi147 & n20891;
  assign n20893 = pi215 & ~n20838;
  assign n20894 = ~n3329 & ~n20832;
  assign n20895 = pi907 & n16518;
  assign n20896 = ~pi947 & n20895;
  assign n20897 = n3329 & ~n20896;
  assign n20898 = ~n20894 & ~n20897;
  assign n20899 = ~pi215 & ~n20898;
  assign n20900 = ~n20893 & ~n20899;
  assign n20901 = pi299 & ~n20900;
  assign n20902 = n17179 & n20755;
  assign n20903 = ~pi299 & ~n20902;
  assign n20904 = ~n20901 & ~n20903;
  assign n20905 = pi39 & ~n20904;
  assign n20906 = n17120 & n20755;
  assign n20907 = ~pi39 & ~n20906;
  assign n20908 = ~n20905 & ~n20907;
  assign n20909 = pi147 & n20908;
  assign n20910 = ~pi38 & ~n20909;
  assign n20911 = ~n20892 & n20910;
  assign n20912 = ~pi147 & ~n17280;
  assign n20913 = n17280 & n20755;
  assign n20914 = pi38 & ~n20913;
  assign n20915 = ~n20912 & n20914;
  assign n20916 = pi770 & ~n20915;
  assign n20917 = ~n20911 & n20916;
  assign n20918 = pi299 & pi947;
  assign n20919 = pi299 & ~n20883;
  assign n20920 = ~n20918 & ~n20919;
  assign n20921 = ~n6183 & n17179;
  assign n20922 = ~pi299 & n20921;
  assign n20923 = ~n17180 & ~n20922;
  assign n20924 = n20920 & n20923;
  assign n20925 = pi39 & n20924;
  assign n20926 = ~n6183 & n17120;
  assign n20927 = ~pi39 & ~n20926;
  assign n20928 = n17120 & n20927;
  assign n20929 = ~n20925 & ~n20928;
  assign n20930 = ~pi147 & n20929;
  assign n20931 = ~n6183 & n16518;
  assign n20932 = n3329 & n20931;
  assign n20933 = ~pi215 & ~n20932;
  assign n20934 = ~n17187 & n20933;
  assign n20935 = pi215 & ~n17190;
  assign n20936 = pi299 & ~n20935;
  assign n20937 = ~n20934 & n20936;
  assign n20938 = ~n20922 & ~n20937;
  assign n20939 = pi39 & n20938;
  assign n20940 = ~n20927 & ~n20939;
  assign n20941 = pi147 & n20940;
  assign n20942 = ~pi38 & ~n20941;
  assign n20943 = ~n20930 & n20942;
  assign n20944 = n6183 & n17397;
  assign n20945 = ~pi147 & ~n20944;
  assign n20946 = ~n6183 & n17280;
  assign n20947 = pi38 & ~n20946;
  assign n20948 = ~n20945 & n20947;
  assign n20949 = ~pi770 & ~n20948;
  assign n20950 = ~n20943 & n20949;
  assign n20951 = pi726 & ~n20950;
  assign n20952 = ~n20917 & n20951;
  assign n20953 = n10143 & ~n20952;
  assign n20954 = ~n20877 & n20953;
  assign n20955 = ~pi147 & ~n10143;
  assign n20956 = ~pi832 & ~n20955;
  assign n20957 = ~n20954 & n20956;
  assign po304 = ~n20826 & ~n20957;
  assign n20959 = ~pi148 & n20924;
  assign n20960 = pi148 & n20938;
  assign n20961 = pi749 & ~n20960;
  assign n20962 = ~n20959 & n20961;
  assign n20963 = ~n9684 & ~n20887;
  assign n20964 = ~n17180 & ~n20901;
  assign n20965 = pi148 & ~n20964;
  assign n20966 = ~pi749 & ~n20965;
  assign n20967 = ~n20963 & n20966;
  assign n20968 = pi39 & ~n20967;
  assign n20969 = ~n20962 & n20968;
  assign n20970 = ~pi148 & ~n17120;
  assign n20971 = ~pi39 & ~n20970;
  assign n20972 = ~pi749 & pi947;
  assign n20973 = n20926 & ~n20972;
  assign n20974 = n20971 & ~n20973;
  assign n20975 = ~pi38 & ~n20974;
  assign n20976 = ~n20969 & n20975;
  assign n20977 = n20946 & ~n20972;
  assign n20978 = ~pi148 & ~n17280;
  assign n20979 = ~n20977 & ~n20978;
  assign n20980 = pi38 & ~n20979;
  assign n20981 = pi706 & ~n20980;
  assign n20982 = ~n20976 & n20981;
  assign n20983 = n3267 & n6286;
  assign n20984 = ~pi148 & ~n20840;
  assign n20985 = ~n20860 & ~n20867;
  assign n20986 = pi148 & ~n20985;
  assign n20987 = pi299 & ~n20986;
  assign n20988 = ~n20984 & n20987;
  assign n20989 = ~pi148 & ~n17179;
  assign n20990 = n20858 & ~n20989;
  assign n20991 = pi749 & ~n20990;
  assign n20992 = ~n20988 & n20991;
  assign n20993 = ~pi148 & ~pi749;
  assign n20994 = ~n17199 & n20993;
  assign n20995 = pi39 & ~n20994;
  assign n20996 = ~n20992 & n20995;
  assign n20997 = pi749 & pi947;
  assign n20998 = n17120 & n20997;
  assign n20999 = n20971 & ~n20998;
  assign n21000 = ~pi38 & ~n20999;
  assign n21001 = ~n20996 & n21000;
  assign n21002 = pi148 & ~n17397;
  assign n21003 = n17280 & ~n20997;
  assign n21004 = pi38 & ~n21003;
  assign n21005 = ~n21002 & n21004;
  assign n21006 = ~pi706 & ~n21005;
  assign n21007 = ~n21001 & n21006;
  assign n21008 = n20983 & ~n21007;
  assign n21009 = ~n20982 & n21008;
  assign n21010 = ~pi148 & ~n20983;
  assign n21011 = ~pi57 & ~n21010;
  assign n21012 = ~n21009 & n21011;
  assign n21013 = pi57 & pi148;
  assign n21014 = ~pi832 & ~n21013;
  assign n21015 = ~n21012 & n21014;
  assign n21016 = pi706 & n20755;
  assign n21017 = n2754 & ~n20997;
  assign n21018 = ~n21016 & n21017;
  assign n21019 = pi148 & ~n2754;
  assign n21020 = pi832 & ~n21019;
  assign n21021 = ~n21018 & n21020;
  assign po305 = n21015 | n21021;
  assign n21023 = ~pi755 & pi947;
  assign n21024 = ~pi725 & n20755;
  assign n21025 = ~n21023 & ~n21024;
  assign n21026 = n2754 & ~n21025;
  assign n21027 = ~pi149 & ~n2754;
  assign n21028 = pi832 & ~n21027;
  assign n21029 = ~n21026 & n21028;
  assign n21030 = pi149 & ~n17397;
  assign n21031 = n17280 & ~n21023;
  assign n21032 = pi38 & ~n21031;
  assign n21033 = ~n21030 & n21032;
  assign n21034 = ~pi149 & ~n20840;
  assign n21035 = ~n16029 & ~n20868;
  assign n21036 = ~n21034 & ~n21035;
  assign n21037 = ~pi149 & ~n17179;
  assign n21038 = n20858 & ~n21037;
  assign n21039 = ~pi755 & ~n21038;
  assign n21040 = ~n21036 & n21039;
  assign n21041 = ~pi149 & pi755;
  assign n21042 = ~n17199 & n21041;
  assign n21043 = pi39 & ~n21042;
  assign n21044 = ~n21040 & n21043;
  assign n21045 = n17120 & n21023;
  assign n21046 = ~pi149 & ~n17120;
  assign n21047 = ~pi39 & ~n21046;
  assign n21048 = ~n21045 & n21047;
  assign n21049 = ~pi38 & ~n21048;
  assign n21050 = ~n21044 & n21049;
  assign n21051 = ~n21033 & ~n21050;
  assign n21052 = pi725 & ~n21051;
  assign n21053 = ~n20906 & n21048;
  assign n21054 = ~pi149 & n20924;
  assign n21055 = pi149 & n20938;
  assign n21056 = ~pi755 & ~n21055;
  assign n21057 = ~n21054 & n21056;
  assign n21058 = ~pi149 & n20885;
  assign n21059 = pi149 & ~n20964;
  assign n21060 = pi755 & ~n20886;
  assign n21061 = ~n21059 & n21060;
  assign n21062 = ~n21058 & n21061;
  assign n21063 = pi39 & ~n21062;
  assign n21064 = ~n21057 & n21063;
  assign n21065 = ~n21053 & ~n21064;
  assign n21066 = ~pi38 & ~n21065;
  assign n21067 = ~n6183 & n16529;
  assign n21068 = pi755 & pi947;
  assign n21069 = ~pi39 & ~n21068;
  assign n21070 = n21067 & n21069;
  assign n21071 = ~pi149 & ~n17280;
  assign n21072 = pi38 & ~n21071;
  assign n21073 = ~n21070 & n21072;
  assign n21074 = ~pi725 & ~n21073;
  assign n21075 = ~n21066 & n21074;
  assign n21076 = ~n21052 & ~n21075;
  assign n21077 = n10143 & ~n21076;
  assign n21078 = ~pi149 & ~n10143;
  assign n21079 = ~pi832 & ~n21078;
  assign n21080 = ~n21077 & n21079;
  assign po306 = ~n21029 & ~n21080;
  assign n21082 = ~pi150 & n20843;
  assign n21083 = pi150 & ~n20869;
  assign n21084 = ~pi751 & ~n21083;
  assign n21085 = ~n21082 & n21084;
  assign n21086 = ~pi150 & pi751;
  assign n21087 = ~n17199 & n21086;
  assign n21088 = ~n21085 & ~n21087;
  assign n21089 = pi39 & ~n21088;
  assign n21090 = pi150 & ~n17120;
  assign n21091 = pi751 & n17120;
  assign n21092 = ~n21090 & ~n21091;
  assign n21093 = n20828 & n21092;
  assign n21094 = ~pi38 & ~n21093;
  assign n21095 = ~n21089 & n21094;
  assign n21096 = pi150 & ~n17397;
  assign n21097 = ~pi751 & pi947;
  assign n21098 = n17280 & ~n21097;
  assign n21099 = ~n21096 & ~n21098;
  assign n21100 = pi38 & ~n21099;
  assign n21101 = pi701 & ~n21100;
  assign n21102 = ~n21095 & n21101;
  assign n21103 = ~pi150 & ~n20887;
  assign n21104 = pi150 & ~n20904;
  assign n21105 = pi751 & ~n21104;
  assign n21106 = ~n21103 & n21105;
  assign n21107 = ~pi150 & n20924;
  assign n21108 = pi150 & n20938;
  assign n21109 = ~pi751 & ~n21108;
  assign n21110 = ~n21107 & n21109;
  assign n21111 = ~n21106 & ~n21110;
  assign n21112 = pi39 & ~n21111;
  assign n21113 = n20889 & ~n21097;
  assign n21114 = ~pi39 & ~n21090;
  assign n21115 = ~n21113 & n21114;
  assign n21116 = ~pi38 & ~n21115;
  assign n21117 = ~n21112 & n21116;
  assign n21118 = pi751 & pi947;
  assign n21119 = ~pi39 & ~n21118;
  assign n21120 = n21067 & n21119;
  assign n21121 = ~pi150 & ~n17280;
  assign n21122 = pi38 & ~n21121;
  assign n21123 = ~n21120 & n21122;
  assign n21124 = ~pi701 & ~n21123;
  assign n21125 = ~n21117 & n21124;
  assign n21126 = ~n21102 & ~n21125;
  assign n21127 = n10143 & ~n21126;
  assign n21128 = ~pi150 & ~n10143;
  assign n21129 = ~pi832 & ~n21128;
  assign n21130 = ~n21127 & n21129;
  assign n21131 = ~pi701 & n20755;
  assign n21132 = ~n21097 & ~n21131;
  assign n21133 = n2754 & ~n21132;
  assign n21134 = ~pi150 & ~n2754;
  assign n21135 = pi832 & ~n21134;
  assign n21136 = ~n21133 & n21135;
  assign po307 = ~n21130 & ~n21136;
  assign n21138 = ~pi745 & pi947;
  assign n21139 = ~pi723 & n20755;
  assign n21140 = ~n21138 & ~n21139;
  assign n21141 = n2754 & ~n21140;
  assign n21142 = ~pi151 & ~n2754;
  assign n21143 = pi832 & ~n21142;
  assign n21144 = ~n21141 & n21143;
  assign n21145 = ~pi151 & ~n17120;
  assign n21146 = ~pi745 & n20855;
  assign n21147 = ~n21145 & ~n21146;
  assign n21148 = n20907 & n21147;
  assign n21149 = ~n17194 & ~n20838;
  assign n21150 = ~pi151 & n21149;
  assign n21151 = ~n17190 & ~n21150;
  assign n21152 = pi215 & ~n21151;
  assign n21153 = pi151 & ~n3329;
  assign n21154 = ~n17186 & n21153;
  assign n21155 = ~n17185 & ~n21154;
  assign n21156 = ~pi151 & ~n16518;
  assign n21157 = n20897 & ~n21156;
  assign n21158 = ~n20931 & n21157;
  assign n21159 = ~pi215 & ~n21158;
  assign n21160 = n21155 & n21159;
  assign n21161 = ~n21152 & ~n21160;
  assign n21162 = pi299 & ~n21161;
  assign n21163 = pi151 & ~n20921;
  assign n21164 = ~n20923 & ~n21163;
  assign n21165 = ~n21162 & ~n21164;
  assign n21166 = ~pi745 & ~n21165;
  assign n21167 = n21155 & ~n21157;
  assign n21168 = n20881 & n21167;
  assign n21169 = ~n21152 & ~n21168;
  assign n21170 = ~n20860 & ~n21169;
  assign n21171 = pi299 & ~n21170;
  assign n21172 = ~pi151 & ~n17179;
  assign n21173 = n20903 & ~n21172;
  assign n21174 = pi745 & ~n21173;
  assign n21175 = ~n21171 & n21174;
  assign n21176 = pi39 & ~n21175;
  assign n21177 = ~n21166 & n21176;
  assign n21178 = ~n21148 & ~n21177;
  assign n21179 = ~pi38 & ~n21178;
  assign n21180 = pi745 & pi947;
  assign n21181 = ~pi39 & ~n21180;
  assign n21182 = n21067 & n21181;
  assign n21183 = ~pi151 & ~n17280;
  assign n21184 = pi38 & ~n21183;
  assign n21185 = ~n21182 & n21184;
  assign n21186 = ~pi723 & ~n21185;
  assign n21187 = ~n21179 & n21186;
  assign n21188 = ~pi745 & ~n17180;
  assign n21189 = ~pi151 & ~n17199;
  assign n21190 = ~n21188 & n21189;
  assign n21191 = n20865 & ~n21156;
  assign n21192 = n21155 & ~n21191;
  assign n21193 = n20835 & n21192;
  assign n21194 = n20893 & ~n21151;
  assign n21195 = pi299 & ~n21194;
  assign n21196 = ~n21193 & n21195;
  assign n21197 = ~pi745 & ~n20858;
  assign n21198 = ~n21196 & n21197;
  assign n21199 = ~n21190 & ~n21198;
  assign n21200 = pi39 & ~n21199;
  assign n21201 = ~pi39 & ~n21147;
  assign n21202 = ~pi38 & ~n21201;
  assign n21203 = ~n21200 & n21202;
  assign n21204 = pi151 & ~n17397;
  assign n21205 = n17280 & ~n21138;
  assign n21206 = ~n21204 & ~n21205;
  assign n21207 = pi38 & ~n21206;
  assign n21208 = pi723 & ~n21207;
  assign n21209 = ~n21203 & n21208;
  assign n21210 = ~n21187 & ~n21209;
  assign n21211 = n10143 & ~n21210;
  assign n21212 = ~pi151 & ~n10143;
  assign n21213 = ~pi832 & ~n21212;
  assign n21214 = ~n21211 & n21213;
  assign po308 = ~n21144 & ~n21214;
  assign n21216 = ~pi152 & ~n17175;
  assign n21217 = ~pi947 & n17175;
  assign n21218 = ~n3052 & ~n21217;
  assign n21219 = ~n21216 & n21218;
  assign n21220 = ~n6183 & n17175;
  assign n21221 = ~n3052 & ~n21220;
  assign n21222 = ~n21219 & n21221;
  assign n21223 = pi152 & ~n16518;
  assign n21224 = ~n20931 & ~n21223;
  assign n21225 = n3052 & n21224;
  assign n21226 = ~pi223 & ~n21225;
  assign n21227 = ~n21222 & n21226;
  assign n21228 = n17153 & ~n20755;
  assign n21229 = pi223 & ~n21228;
  assign n21230 = ~pi152 & ~n17153;
  assign n21231 = n21229 & ~n21230;
  assign n21232 = ~pi947 & n17153;
  assign n21233 = pi223 & ~n21232;
  assign n21234 = ~n21230 & n21233;
  assign n21235 = ~pi299 & ~n21234;
  assign n21236 = ~n21231 & n21235;
  assign n21237 = ~n21227 & n21236;
  assign n21238 = n3329 & n21224;
  assign n21239 = ~pi215 & ~n21238;
  assign n21240 = pi152 & n20879;
  assign n21241 = n20894 & ~n21240;
  assign n21242 = ~n17186 & n21241;
  assign n21243 = n21239 & ~n21242;
  assign n21244 = ~pi152 & ~n17190;
  assign n21245 = n20837 & ~n21244;
  assign n21246 = pi299 & ~n21245;
  assign n21247 = ~n21243 & n21246;
  assign n21248 = pi759 & ~n21247;
  assign n21249 = ~n21237 & n21248;
  assign n21250 = ~n20896 & ~n21223;
  assign n21251 = n3052 & ~n21250;
  assign n21252 = n17175 & ~n20755;
  assign n21253 = ~n3052 & ~n21252;
  assign n21254 = ~n21216 & n21253;
  assign n21255 = ~n21251 & ~n21254;
  assign n21256 = ~pi223 & ~n21255;
  assign n21257 = ~pi299 & ~n21231;
  assign n21258 = ~n21256 & n21257;
  assign n21259 = ~n20878 & n21239;
  assign n21260 = ~n21241 & n21259;
  assign n21261 = ~n20755 & ~n20935;
  assign n21262 = n21245 & ~n21261;
  assign n21263 = pi299 & ~n21262;
  assign n21264 = ~n21260 & n21263;
  assign n21265 = ~pi759 & ~n21264;
  assign n21266 = ~n21258 & n21265;
  assign n21267 = pi39 & ~n21266;
  assign n21268 = ~n21249 & n21267;
  assign n21269 = pi152 & ~n17120;
  assign n21270 = pi759 & pi947;
  assign n21271 = ~pi39 & ~n21270;
  assign n21272 = ~n17121 & ~n21271;
  assign n21273 = ~n21269 & ~n21272;
  assign n21274 = ~n20906 & n21273;
  assign n21275 = ~pi38 & ~n21274;
  assign n21276 = ~n21268 & n21275;
  assign n21277 = n16529 & ~n20755;
  assign n21278 = n21271 & n21277;
  assign n21279 = ~pi152 & ~n17280;
  assign n21280 = pi38 & ~n21279;
  assign n21281 = ~n21278 & n21280;
  assign n21282 = pi696 & ~n21281;
  assign n21283 = ~n21276 & n21282;
  assign n21284 = ~n20834 & ~n21241;
  assign n21285 = ~n20862 & ~n21284;
  assign n21286 = ~n20864 & ~n21223;
  assign n21287 = n3329 & n21286;
  assign n21288 = ~pi215 & ~n21287;
  assign n21289 = ~n21285 & n21288;
  assign n21290 = pi152 & n20839;
  assign n21291 = n20861 & ~n21290;
  assign n21292 = ~n21289 & n21291;
  assign n21293 = n3052 & ~n21286;
  assign n21294 = ~n21219 & ~n21293;
  assign n21295 = ~pi223 & ~n21294;
  assign n21296 = n21235 & ~n21295;
  assign n21297 = pi759 & ~n21296;
  assign n21298 = ~n21292 & n21297;
  assign n21299 = ~pi759 & ~n17199;
  assign n21300 = pi152 & n21299;
  assign n21301 = pi39 & ~n21300;
  assign n21302 = ~n21298 & n21301;
  assign n21303 = ~pi38 & ~n21273;
  assign n21304 = ~n21302 & n21303;
  assign n21305 = ~pi152 & ~n17397;
  assign n21306 = n17280 & ~n21270;
  assign n21307 = pi38 & ~n21306;
  assign n21308 = ~n21305 & n21307;
  assign n21309 = ~pi696 & ~n21308;
  assign n21310 = ~n21304 & n21309;
  assign n21311 = ~n21283 & ~n21310;
  assign n21312 = n10143 & ~n21311;
  assign n21313 = ~pi152 & ~n10143;
  assign n21314 = ~pi832 & ~n21313;
  assign n21315 = ~n21312 & n21314;
  assign n21316 = pi696 & n20755;
  assign n21317 = n2754 & ~n21270;
  assign n21318 = ~n21316 & n21317;
  assign n21319 = ~pi152 & ~n2754;
  assign n21320 = pi832 & ~n21319;
  assign n21321 = ~n21318 & n21320;
  assign po309 = n21315 | n21321;
  assign n21323 = pi766 & pi947;
  assign n21324 = n2754 & ~n21323;
  assign n21325 = pi700 & n20755;
  assign n21326 = n21324 & ~n21325;
  assign n21327 = pi153 & ~n2754;
  assign n21328 = pi832 & ~n21327;
  assign n21329 = ~n21326 & n21328;
  assign n21330 = ~pi153 & ~n17120;
  assign n21331 = ~pi766 & n17954;
  assign n21332 = ~n20856 & ~n21331;
  assign n21333 = ~n21330 & ~n21332;
  assign n21334 = ~n20906 & n21333;
  assign n21335 = pi153 & ~n17190;
  assign n21336 = n20837 & ~n21335;
  assign n21337 = pi153 & ~n3329;
  assign n21338 = ~n17186 & n21337;
  assign n21339 = ~n17185 & ~n21338;
  assign n21340 = ~pi153 & ~n16518;
  assign n21341 = n20865 & ~n21340;
  assign n21342 = ~n20895 & n21341;
  assign n21343 = ~pi215 & ~n21342;
  assign n21344 = n21339 & n21343;
  assign n21345 = ~n21336 & ~n21344;
  assign n21346 = pi299 & ~n21345;
  assign n21347 = pi153 & ~n20921;
  assign n21348 = ~n20923 & ~n21347;
  assign n21349 = ~n21346 & ~n21348;
  assign n21350 = pi766 & ~n21349;
  assign n21351 = n20897 & ~n21340;
  assign n21352 = ~n20880 & ~n21351;
  assign n21353 = n21339 & n21352;
  assign n21354 = ~pi215 & ~n21353;
  assign n21355 = n20935 & ~n21336;
  assign n21356 = ~n20860 & ~n21355;
  assign n21357 = ~n21354 & n21356;
  assign n21358 = pi299 & ~n21357;
  assign n21359 = ~pi153 & ~n17179;
  assign n21360 = n20903 & ~n21359;
  assign n21361 = ~pi766 & ~n21360;
  assign n21362 = ~n21358 & n21361;
  assign n21363 = pi39 & ~n21362;
  assign n21364 = ~n21350 & n21363;
  assign n21365 = ~n21334 & ~n21364;
  assign n21366 = ~pi38 & ~n21365;
  assign n21367 = ~pi766 & pi947;
  assign n21368 = ~pi39 & ~n21367;
  assign n21369 = n21067 & n21368;
  assign n21370 = ~pi153 & ~n17280;
  assign n21371 = pi38 & ~n21370;
  assign n21372 = ~n21369 & n21371;
  assign n21373 = ~n21366 & ~n21372;
  assign n21374 = pi700 & ~n21373;
  assign n21375 = n20858 & ~n21359;
  assign n21376 = n21339 & ~n21341;
  assign n21377 = n20835 & n21376;
  assign n21378 = n20839 & ~n21335;
  assign n21379 = pi299 & ~n21378;
  assign n21380 = ~n21377 & n21379;
  assign n21381 = pi766 & ~n21380;
  assign n21382 = ~n21375 & n21381;
  assign n21383 = ~pi153 & ~pi766;
  assign n21384 = ~n17199 & n21383;
  assign n21385 = pi39 & ~n21384;
  assign n21386 = ~n21382 & n21385;
  assign n21387 = ~pi38 & ~n21333;
  assign n21388 = ~n21386 & n21387;
  assign n21389 = pi153 & ~n17397;
  assign n21390 = n6234 & n21324;
  assign n21391 = pi38 & ~n21390;
  assign n21392 = ~n21389 & n21391;
  assign n21393 = ~pi700 & ~n21392;
  assign n21394 = ~n21388 & n21393;
  assign n21395 = n20983 & ~n21394;
  assign n21396 = ~n21374 & n21395;
  assign n21397 = ~pi153 & ~n20983;
  assign n21398 = ~pi57 & ~n21397;
  assign n21399 = ~n21396 & n21398;
  assign n21400 = pi57 & pi153;
  assign n21401 = ~pi832 & ~n21400;
  assign n21402 = ~n21399 & n21401;
  assign po310 = n21329 | n21402;
  assign n21404 = ~pi742 & pi947;
  assign n21405 = ~pi704 & n20755;
  assign n21406 = ~n21404 & ~n21405;
  assign n21407 = n2754 & ~n21406;
  assign n21408 = ~pi154 & ~n2754;
  assign n21409 = pi832 & ~n21408;
  assign n21410 = ~n21407 & n21409;
  assign n21411 = ~pi154 & ~n17120;
  assign n21412 = n20907 & ~n21411;
  assign n21413 = ~n20926 & n21412;
  assign n21414 = ~pi154 & ~n20924;
  assign n21415 = pi154 & ~n20938;
  assign n21416 = pi39 & ~n21415;
  assign n21417 = ~n21414 & n21416;
  assign n21418 = ~n21413 & ~n21417;
  assign n21419 = ~pi38 & ~n21418;
  assign n21420 = ~pi154 & ~n17280;
  assign n21421 = n20947 & ~n21420;
  assign n21422 = ~pi742 & ~n21421;
  assign n21423 = ~n21419 & n21422;
  assign n21424 = ~pi154 & n20887;
  assign n21425 = pi154 & n20904;
  assign n21426 = pi39 & ~n21425;
  assign n21427 = ~n21424 & n21426;
  assign n21428 = ~n21412 & ~n21427;
  assign n21429 = ~pi38 & ~n21428;
  assign n21430 = n20914 & ~n21420;
  assign n21431 = pi742 & ~n21430;
  assign n21432 = ~n21429 & n21431;
  assign n21433 = ~pi704 & ~n21432;
  assign n21434 = ~n21423 & n21433;
  assign n21435 = n20856 & ~n21411;
  assign n21436 = ~pi154 & ~n20843;
  assign n21437 = pi154 & n20869;
  assign n21438 = pi39 & ~n21437;
  assign n21439 = ~n21436 & n21438;
  assign n21440 = ~n21435 & ~n21439;
  assign n21441 = ~pi38 & ~n21440;
  assign n21442 = ~pi154 & ~n17397;
  assign n21443 = ~n20854 & ~n21442;
  assign n21444 = ~pi742 & ~n21443;
  assign n21445 = ~n21441 & n21444;
  assign n21446 = ~pi154 & pi742;
  assign n21447 = ~n17399 & n21446;
  assign n21448 = pi704 & ~n21447;
  assign n21449 = ~n21445 & n21448;
  assign n21450 = n10143 & ~n21449;
  assign n21451 = ~n21434 & n21450;
  assign n21452 = ~pi154 & ~n10143;
  assign n21453 = ~pi832 & ~n21452;
  assign n21454 = ~n21451 & n21453;
  assign po311 = ~n21410 & ~n21454;
  assign n21456 = ~pi38 & ~n20908;
  assign n21457 = ~n20914 & ~n21456;
  assign n21458 = pi757 & n21457;
  assign n21459 = ~pi38 & ~n20940;
  assign n21460 = ~n20947 & ~n21459;
  assign n21461 = ~pi757 & n21460;
  assign n21462 = ~pi686 & ~n21461;
  assign n21463 = ~n21458 & n21462;
  assign n21464 = ~pi757 & n20873;
  assign n21465 = pi686 & ~n21464;
  assign n21466 = n10143 & ~n21465;
  assign n21467 = ~n21463 & n21466;
  assign n21468 = pi155 & ~n21467;
  assign n21469 = ~pi38 & ~n20891;
  assign n21470 = n17280 & n20914;
  assign n21471 = ~n21469 & ~n21470;
  assign n21472 = pi757 & n21471;
  assign n21473 = ~pi38 & ~n20929;
  assign n21474 = pi38 & n20944;
  assign n21475 = ~n21473 & ~n21474;
  assign n21476 = ~pi757 & n21475;
  assign n21477 = ~pi686 & ~n21476;
  assign n21478 = ~n21472 & n21477;
  assign n21479 = ~pi757 & n20849;
  assign n21480 = pi757 & ~n17399;
  assign n21481 = pi686 & ~n21480;
  assign n21482 = ~n21479 & n21481;
  assign n21483 = ~n21478 & ~n21482;
  assign n21484 = ~pi155 & n10143;
  assign n21485 = ~n21483 & n21484;
  assign n21486 = ~n21468 & ~n21485;
  assign n21487 = ~pi832 & ~n21486;
  assign n21488 = ~pi757 & pi947;
  assign n21489 = ~pi686 & n20755;
  assign n21490 = ~n21488 & ~n21489;
  assign n21491 = n2754 & ~n21490;
  assign n21492 = ~pi155 & ~n2754;
  assign n21493 = pi832 & ~n21492;
  assign n21494 = ~n21491 & n21493;
  assign po312 = ~n21487 & ~n21494;
  assign n21496 = ~pi741 & pi947;
  assign n21497 = ~pi724 & n20755;
  assign n21498 = ~n21496 & ~n21497;
  assign n21499 = n2754 & ~n21498;
  assign n21500 = ~pi156 & ~n2754;
  assign n21501 = pi832 & ~n21500;
  assign n21502 = ~n21499 & n21501;
  assign n21503 = pi741 & ~n21471;
  assign n21504 = ~pi741 & ~n21475;
  assign n21505 = ~pi724 & ~n21504;
  assign n21506 = ~n21503 & n21505;
  assign n21507 = ~pi741 & ~n20849;
  assign n21508 = pi741 & n17399;
  assign n21509 = pi724 & ~n21508;
  assign n21510 = ~n21507 & n21509;
  assign n21511 = n10143 & ~n21510;
  assign n21512 = ~n21506 & n21511;
  assign n21513 = ~pi156 & ~n21512;
  assign n21514 = pi741 & ~n21457;
  assign n21515 = ~pi741 & ~n21460;
  assign n21516 = ~pi724 & ~n21515;
  assign n21517 = ~n21514 & n21516;
  assign n21518 = pi724 & ~pi741;
  assign n21519 = n20873 & n21518;
  assign n21520 = ~n21517 & ~n21519;
  assign n21521 = pi156 & n10143;
  assign n21522 = ~n21520 & n21521;
  assign n21523 = ~pi832 & ~n21522;
  assign n21524 = ~n21513 & n21523;
  assign po313 = ~n21502 & ~n21524;
  assign n21526 = ~pi760 & pi947;
  assign n21527 = ~pi688 & n20755;
  assign n21528 = ~n21526 & ~n21527;
  assign n21529 = n2754 & ~n21528;
  assign n21530 = ~pi157 & ~n2754;
  assign n21531 = pi832 & ~n21530;
  assign n21532 = ~n21529 & n21531;
  assign n21533 = pi157 & ~n17397;
  assign n21534 = n17280 & ~n21526;
  assign n21535 = pi38 & ~n21534;
  assign n21536 = ~n21533 & n21535;
  assign n21537 = ~pi157 & ~n20840;
  assign n21538 = ~n13723 & ~n20868;
  assign n21539 = ~n21537 & ~n21538;
  assign n21540 = ~pi157 & ~n17179;
  assign n21541 = n20858 & ~n21540;
  assign n21542 = ~pi760 & ~n21541;
  assign n21543 = ~n21539 & n21542;
  assign n21544 = ~pi157 & pi760;
  assign n21545 = ~n17199 & n21544;
  assign n21546 = pi39 & ~n21545;
  assign n21547 = ~n21543 & n21546;
  assign n21548 = n17120 & n21526;
  assign n21549 = ~pi157 & ~n17120;
  assign n21550 = ~pi39 & ~n21549;
  assign n21551 = ~n21548 & n21550;
  assign n21552 = ~pi38 & ~n21551;
  assign n21553 = ~n21547 & n21552;
  assign n21554 = ~n21536 & ~n21553;
  assign n21555 = pi688 & ~n21554;
  assign n21556 = ~n20906 & n21551;
  assign n21557 = ~pi760 & n20924;
  assign n21558 = pi760 & ~n20887;
  assign n21559 = ~pi157 & ~n21558;
  assign n21560 = ~n21557 & n21559;
  assign n21561 = pi760 & ~n20904;
  assign n21562 = ~pi760 & n20938;
  assign n21563 = pi157 & ~n21562;
  assign n21564 = ~n21561 & n21563;
  assign n21565 = pi39 & ~n21564;
  assign n21566 = ~n21560 & n21565;
  assign n21567 = ~n21556 & ~n21566;
  assign n21568 = ~pi38 & ~n21567;
  assign n21569 = pi760 & pi947;
  assign n21570 = ~pi39 & ~n21569;
  assign n21571 = n21067 & n21570;
  assign n21572 = ~pi157 & ~n17280;
  assign n21573 = pi38 & ~n21572;
  assign n21574 = ~n21571 & n21573;
  assign n21575 = ~pi688 & ~n21574;
  assign n21576 = ~n21568 & n21575;
  assign n21577 = ~n21555 & ~n21576;
  assign n21578 = n10143 & ~n21577;
  assign n21579 = ~pi157 & ~n10143;
  assign n21580 = ~pi832 & ~n21579;
  assign n21581 = ~n21578 & n21580;
  assign po314 = ~n21532 & ~n21581;
  assign n21583 = ~pi158 & n20843;
  assign n21584 = pi158 & ~n20869;
  assign n21585 = ~pi753 & ~n21584;
  assign n21586 = ~n21583 & n21585;
  assign n21587 = ~pi158 & pi753;
  assign n21588 = ~n17199 & n21587;
  assign n21589 = ~n21586 & ~n21588;
  assign n21590 = pi39 & ~n21589;
  assign n21591 = pi158 & ~n17120;
  assign n21592 = pi753 & n17120;
  assign n21593 = ~n21591 & ~n21592;
  assign n21594 = n20828 & n21593;
  assign n21595 = ~pi38 & ~n21594;
  assign n21596 = ~n21590 & n21595;
  assign n21597 = pi158 & ~n17397;
  assign n21598 = ~pi753 & pi947;
  assign n21599 = n17280 & ~n21598;
  assign n21600 = ~n21597 & ~n21599;
  assign n21601 = pi38 & ~n21600;
  assign n21602 = pi702 & ~n21601;
  assign n21603 = ~n21596 & n21602;
  assign n21604 = ~pi158 & ~n20887;
  assign n21605 = pi158 & ~n20904;
  assign n21606 = pi753 & ~n21605;
  assign n21607 = ~n21604 & n21606;
  assign n21608 = ~pi158 & n20924;
  assign n21609 = pi158 & n20938;
  assign n21610 = ~pi753 & ~n21609;
  assign n21611 = ~n21608 & n21610;
  assign n21612 = ~n21607 & ~n21611;
  assign n21613 = pi39 & ~n21612;
  assign n21614 = n20889 & ~n21598;
  assign n21615 = ~pi39 & ~n21591;
  assign n21616 = ~n21614 & n21615;
  assign n21617 = ~pi38 & ~n21616;
  assign n21618 = ~n21613 & n21617;
  assign n21619 = pi753 & pi947;
  assign n21620 = ~pi39 & ~n21619;
  assign n21621 = n21067 & n21620;
  assign n21622 = ~pi158 & ~n17280;
  assign n21623 = pi38 & ~n21622;
  assign n21624 = ~n21621 & n21623;
  assign n21625 = ~pi702 & ~n21624;
  assign n21626 = ~n21618 & n21625;
  assign n21627 = ~n21603 & ~n21626;
  assign n21628 = n10143 & ~n21627;
  assign n21629 = ~pi158 & ~n10143;
  assign n21630 = ~pi832 & ~n21629;
  assign n21631 = ~n21628 & n21630;
  assign n21632 = ~pi702 & n20755;
  assign n21633 = ~n21598 & ~n21632;
  assign n21634 = n2754 & ~n21633;
  assign n21635 = ~pi158 & ~n2754;
  assign n21636 = pi832 & ~n21635;
  assign n21637 = ~n21634 & n21636;
  assign po315 = ~n21631 & ~n21637;
  assign n21639 = ~pi159 & n20843;
  assign n21640 = pi159 & ~n20869;
  assign n21641 = ~pi754 & ~n21640;
  assign n21642 = ~n21639 & n21641;
  assign n21643 = ~pi159 & pi754;
  assign n21644 = ~n17199 & n21643;
  assign n21645 = ~n21642 & ~n21644;
  assign n21646 = pi39 & ~n21645;
  assign n21647 = pi159 & ~n17120;
  assign n21648 = pi754 & n17120;
  assign n21649 = ~n21647 & ~n21648;
  assign n21650 = n20828 & n21649;
  assign n21651 = ~pi38 & ~n21650;
  assign n21652 = ~n21646 & n21651;
  assign n21653 = pi159 & ~n17397;
  assign n21654 = ~pi754 & pi947;
  assign n21655 = n17280 & ~n21654;
  assign n21656 = ~n21653 & ~n21655;
  assign n21657 = pi38 & ~n21656;
  assign n21658 = pi709 & ~n21657;
  assign n21659 = ~n21652 & n21658;
  assign n21660 = ~pi159 & ~n20887;
  assign n21661 = pi159 & ~n20904;
  assign n21662 = pi754 & ~n21661;
  assign n21663 = ~n21660 & n21662;
  assign n21664 = ~pi159 & n20924;
  assign n21665 = pi159 & n20938;
  assign n21666 = ~pi754 & ~n21665;
  assign n21667 = ~n21664 & n21666;
  assign n21668 = ~n21663 & ~n21667;
  assign n21669 = pi39 & ~n21668;
  assign n21670 = n20889 & ~n21654;
  assign n21671 = ~pi39 & ~n21647;
  assign n21672 = ~n21670 & n21671;
  assign n21673 = ~pi38 & ~n21672;
  assign n21674 = ~n21669 & n21673;
  assign n21675 = pi754 & pi947;
  assign n21676 = ~pi39 & ~n21675;
  assign n21677 = n21067 & n21676;
  assign n21678 = ~pi159 & ~n17280;
  assign n21679 = pi38 & ~n21678;
  assign n21680 = ~n21677 & n21679;
  assign n21681 = ~pi709 & ~n21680;
  assign n21682 = ~n21674 & n21681;
  assign n21683 = ~n21659 & ~n21682;
  assign n21684 = n10143 & ~n21683;
  assign n21685 = ~pi159 & ~n10143;
  assign n21686 = ~pi832 & ~n21685;
  assign n21687 = ~n21684 & n21686;
  assign n21688 = ~pi709 & n20755;
  assign n21689 = ~n21654 & ~n21688;
  assign n21690 = n2754 & ~n21689;
  assign n21691 = ~pi159 & ~n2754;
  assign n21692 = pi832 & ~n21691;
  assign n21693 = ~n21690 & n21692;
  assign po316 = ~n21687 & ~n21693;
  assign n21695 = ~pi756 & pi947;
  assign n21696 = ~pi734 & n20755;
  assign n21697 = ~n21695 & ~n21696;
  assign n21698 = n2754 & ~n21697;
  assign n21699 = ~pi160 & ~n2754;
  assign n21700 = pi832 & ~n21699;
  assign n21701 = ~n21698 & n21700;
  assign n21702 = pi160 & ~n17397;
  assign n21703 = n17280 & ~n21695;
  assign n21704 = pi38 & ~n21703;
  assign n21705 = ~n21702 & n21704;
  assign n21706 = ~pi160 & ~n20840;
  assign n21707 = pi160 & ~n20985;
  assign n21708 = pi299 & ~n21707;
  assign n21709 = ~n21706 & n21708;
  assign n21710 = ~pi160 & ~n17179;
  assign n21711 = n20858 & ~n21710;
  assign n21712 = ~pi756 & ~n21711;
  assign n21713 = ~n21709 & n21712;
  assign n21714 = ~pi160 & pi756;
  assign n21715 = ~n17199 & n21714;
  assign n21716 = pi39 & ~n21715;
  assign n21717 = ~n21713 & n21716;
  assign n21718 = n17120 & n21695;
  assign n21719 = ~pi160 & ~n17120;
  assign n21720 = ~pi39 & ~n21719;
  assign n21721 = ~n21718 & n21720;
  assign n21722 = ~pi38 & ~n21721;
  assign n21723 = ~n21717 & n21722;
  assign n21724 = ~n21705 & ~n21723;
  assign n21725 = pi734 & ~n21724;
  assign n21726 = ~n20906 & n21721;
  assign n21727 = ~pi160 & n20924;
  assign n21728 = pi160 & n20938;
  assign n21729 = ~pi756 & ~n21728;
  assign n21730 = ~n21727 & n21729;
  assign n21731 = ~pi160 & n20885;
  assign n21732 = pi160 & ~n20964;
  assign n21733 = pi756 & ~n20886;
  assign n21734 = ~n21732 & n21733;
  assign n21735 = ~n21731 & n21734;
  assign n21736 = pi39 & ~n21735;
  assign n21737 = ~n21730 & n21736;
  assign n21738 = ~n21726 & ~n21737;
  assign n21739 = ~pi38 & ~n21738;
  assign n21740 = pi756 & pi947;
  assign n21741 = ~pi39 & ~n21740;
  assign n21742 = n21067 & n21741;
  assign n21743 = ~pi160 & ~n17280;
  assign n21744 = pi38 & ~n21743;
  assign n21745 = ~n21742 & n21744;
  assign n21746 = ~pi734 & ~n21745;
  assign n21747 = ~n21739 & n21746;
  assign n21748 = ~n21725 & ~n21747;
  assign n21749 = n10143 & ~n21748;
  assign n21750 = ~pi160 & ~n10143;
  assign n21751 = ~pi832 & ~n21750;
  assign n21752 = ~n21749 & n21751;
  assign po317 = ~n21701 & ~n21752;
  assign n21754 = ~pi161 & ~n17175;
  assign n21755 = n21218 & ~n21754;
  assign n21756 = n21221 & ~n21755;
  assign n21757 = pi161 & ~n16518;
  assign n21758 = ~n20931 & ~n21757;
  assign n21759 = n3052 & n21758;
  assign n21760 = ~pi223 & ~n21759;
  assign n21761 = ~n21756 & n21760;
  assign n21762 = ~pi161 & ~n17153;
  assign n21763 = n21229 & ~n21762;
  assign n21764 = n21233 & ~n21762;
  assign n21765 = ~pi299 & ~n21764;
  assign n21766 = ~n21763 & n21765;
  assign n21767 = ~n21761 & n21766;
  assign n21768 = n3329 & n21758;
  assign n21769 = ~pi215 & ~n21768;
  assign n21770 = pi161 & n20879;
  assign n21771 = n20894 & ~n21770;
  assign n21772 = ~n17186 & n21771;
  assign n21773 = n21769 & ~n21772;
  assign n21774 = ~pi161 & ~n17190;
  assign n21775 = n20837 & ~n21774;
  assign n21776 = pi299 & ~n21775;
  assign n21777 = ~n21773 & n21776;
  assign n21778 = pi758 & ~n21777;
  assign n21779 = ~n21767 & n21778;
  assign n21780 = ~n20896 & ~n21757;
  assign n21781 = n3052 & ~n21780;
  assign n21782 = n21253 & ~n21754;
  assign n21783 = ~n21781 & ~n21782;
  assign n21784 = ~pi223 & ~n21783;
  assign n21785 = ~pi299 & ~n21763;
  assign n21786 = ~n21784 & n21785;
  assign n21787 = ~n20878 & n21769;
  assign n21788 = ~n21771 & n21787;
  assign n21789 = ~n21261 & n21775;
  assign n21790 = pi299 & ~n21789;
  assign n21791 = ~n21788 & n21790;
  assign n21792 = ~pi758 & ~n21791;
  assign n21793 = ~n21786 & n21792;
  assign n21794 = pi39 & ~n21793;
  assign n21795 = ~n21779 & n21794;
  assign n21796 = pi161 & ~n17120;
  assign n21797 = pi758 & pi947;
  assign n21798 = ~pi39 & ~n21797;
  assign n21799 = ~n17121 & ~n21798;
  assign n21800 = ~n21796 & ~n21799;
  assign n21801 = ~n20906 & n21800;
  assign n21802 = ~pi38 & ~n21801;
  assign n21803 = ~n21795 & n21802;
  assign n21804 = n21277 & n21798;
  assign n21805 = ~pi161 & ~n17280;
  assign n21806 = pi38 & ~n21805;
  assign n21807 = ~n21804 & n21806;
  assign n21808 = pi736 & ~n21807;
  assign n21809 = ~n21803 & n21808;
  assign n21810 = ~n20834 & ~n21771;
  assign n21811 = ~n20862 & ~n21810;
  assign n21812 = ~n20864 & ~n21757;
  assign n21813 = n3329 & n21812;
  assign n21814 = ~pi215 & ~n21813;
  assign n21815 = ~n21811 & n21814;
  assign n21816 = pi161 & n20839;
  assign n21817 = n20861 & ~n21816;
  assign n21818 = ~n21815 & n21817;
  assign n21819 = n3052 & ~n21812;
  assign n21820 = ~n21755 & ~n21819;
  assign n21821 = ~pi223 & ~n21820;
  assign n21822 = n21765 & ~n21821;
  assign n21823 = pi758 & ~n21822;
  assign n21824 = ~n21818 & n21823;
  assign n21825 = pi161 & n19770;
  assign n21826 = pi39 & ~n21825;
  assign n21827 = ~n21824 & n21826;
  assign n21828 = ~pi38 & ~n21800;
  assign n21829 = ~n21827 & n21828;
  assign n21830 = ~pi161 & ~n17397;
  assign n21831 = n17280 & ~n21797;
  assign n21832 = pi38 & ~n21831;
  assign n21833 = ~n21830 & n21832;
  assign n21834 = ~pi736 & ~n21833;
  assign n21835 = ~n21829 & n21834;
  assign n21836 = ~n21809 & ~n21835;
  assign n21837 = n10143 & ~n21836;
  assign n21838 = ~pi161 & ~n10143;
  assign n21839 = ~pi832 & ~n21838;
  assign n21840 = ~n21837 & n21839;
  assign n21841 = pi736 & n20755;
  assign n21842 = n2754 & ~n21797;
  assign n21843 = ~n21841 & n21842;
  assign n21844 = ~pi161 & ~n2754;
  assign n21845 = pi832 & ~n21844;
  assign n21846 = ~n21843 & n21845;
  assign po318 = n21840 | n21846;
  assign n21848 = pi162 & ~n17397;
  assign n21849 = ~pi761 & pi947;
  assign n21850 = n17280 & ~n21849;
  assign n21851 = pi38 & ~n21850;
  assign n21852 = ~n21848 & n21851;
  assign n21853 = ~pi761 & n20842;
  assign n21854 = pi761 & n17199;
  assign n21855 = ~pi162 & ~n21854;
  assign n21856 = ~n21853 & n21855;
  assign n21857 = n15018 & ~n20985;
  assign n21858 = ~n20830 & ~n21857;
  assign n21859 = ~pi761 & ~n21858;
  assign n21860 = pi39 & ~n21859;
  assign n21861 = ~n21856 & n21860;
  assign n21862 = n17120 & n21849;
  assign n21863 = ~pi162 & ~n17120;
  assign n21864 = ~pi39 & ~n21863;
  assign n21865 = ~n21862 & n21864;
  assign n21866 = ~pi38 & ~n21865;
  assign n21867 = ~n21861 & n21866;
  assign n21868 = ~n21852 & ~n21867;
  assign n21869 = pi738 & ~n21868;
  assign n21870 = ~n20906 & n21865;
  assign n21871 = ~pi162 & n20924;
  assign n21872 = pi162 & n20938;
  assign n21873 = ~pi761 & ~n21872;
  assign n21874 = ~n21871 & n21873;
  assign n21875 = ~n15018 & ~n20887;
  assign n21876 = pi162 & ~n20964;
  assign n21877 = pi761 & ~n21876;
  assign n21878 = ~n21875 & n21877;
  assign n21879 = pi39 & ~n21878;
  assign n21880 = ~n21874 & n21879;
  assign n21881 = ~n21870 & ~n21880;
  assign n21882 = ~pi38 & ~n21881;
  assign n21883 = pi761 & pi947;
  assign n21884 = ~pi39 & ~n21883;
  assign n21885 = n21067 & n21884;
  assign n21886 = ~pi162 & ~n17280;
  assign n21887 = pi38 & ~n21886;
  assign n21888 = ~n21885 & n21887;
  assign n21889 = ~pi738 & ~n21888;
  assign n21890 = ~n21882 & n21889;
  assign n21891 = ~n21869 & ~n21890;
  assign n21892 = n10143 & ~n21891;
  assign n21893 = ~pi162 & ~n10143;
  assign n21894 = ~pi832 & ~n21893;
  assign n21895 = ~n21892 & n21894;
  assign n21896 = ~pi738 & n20755;
  assign n21897 = ~n21849 & ~n21896;
  assign n21898 = n2754 & ~n21897;
  assign n21899 = ~pi162 & ~n2754;
  assign n21900 = pi832 & ~n21899;
  assign n21901 = ~n21898 & n21900;
  assign po319 = ~n21895 & ~n21901;
  assign n21903 = ~pi777 & pi947;
  assign n21904 = ~pi737 & n20755;
  assign n21905 = ~n21903 & ~n21904;
  assign n21906 = n2754 & ~n21905;
  assign n21907 = ~pi163 & ~n2754;
  assign n21908 = pi832 & ~n21907;
  assign n21909 = ~n21906 & n21908;
  assign n21910 = pi163 & ~n17397;
  assign n21911 = n17280 & ~n21903;
  assign n21912 = pi38 & ~n21911;
  assign n21913 = ~n21910 & n21912;
  assign n21914 = ~pi163 & ~n20840;
  assign n21915 = ~n14625 & ~n20868;
  assign n21916 = ~n21914 & ~n21915;
  assign n21917 = ~pi163 & ~n17179;
  assign n21918 = n20858 & ~n21917;
  assign n21919 = ~pi777 & ~n21918;
  assign n21920 = ~n21916 & n21919;
  assign n21921 = ~pi163 & pi777;
  assign n21922 = ~n17199 & n21921;
  assign n21923 = pi39 & ~n21922;
  assign n21924 = ~n21920 & n21923;
  assign n21925 = n17120 & n21903;
  assign n21926 = ~pi163 & ~n17120;
  assign n21927 = ~pi39 & ~n21926;
  assign n21928 = ~n21925 & n21927;
  assign n21929 = ~pi38 & ~n21928;
  assign n21930 = ~n21924 & n21929;
  assign n21931 = ~n21913 & ~n21930;
  assign n21932 = pi737 & ~n21931;
  assign n21933 = ~n20906 & n21928;
  assign n21934 = ~pi163 & n20924;
  assign n21935 = pi163 & n20938;
  assign n21936 = ~pi777 & ~n21935;
  assign n21937 = ~n21934 & n21936;
  assign n21938 = ~pi163 & n20885;
  assign n21939 = pi163 & ~n20964;
  assign n21940 = pi777 & ~n20886;
  assign n21941 = ~n21939 & n21940;
  assign n21942 = ~n21938 & n21941;
  assign n21943 = pi39 & ~n21942;
  assign n21944 = ~n21937 & n21943;
  assign n21945 = ~n21933 & ~n21944;
  assign n21946 = ~pi38 & ~n21945;
  assign n21947 = pi777 & pi947;
  assign n21948 = ~pi39 & ~n21947;
  assign n21949 = n21067 & n21948;
  assign n21950 = ~pi163 & ~n17280;
  assign n21951 = pi38 & ~n21950;
  assign n21952 = ~n21949 & n21951;
  assign n21953 = ~pi737 & ~n21952;
  assign n21954 = ~n21946 & n21953;
  assign n21955 = ~n21932 & ~n21954;
  assign n21956 = n10143 & ~n21955;
  assign n21957 = ~pi163 & ~n10143;
  assign n21958 = ~pi832 & ~n21957;
  assign n21959 = ~n21956 & n21958;
  assign po320 = ~n21909 & ~n21959;
  assign n21961 = ~pi752 & pi947;
  assign n21962 = pi703 & n20755;
  assign n21963 = ~n21961 & ~n21962;
  assign n21964 = n2754 & ~n21963;
  assign n21965 = ~pi164 & ~n2754;
  assign n21966 = pi832 & ~n21965;
  assign n21967 = ~n21964 & n21966;
  assign n21968 = ~pi164 & n20929;
  assign n21969 = pi164 & n20940;
  assign n21970 = ~pi38 & ~n21969;
  assign n21971 = ~n21968 & n21970;
  assign n21972 = ~pi164 & ~n20944;
  assign n21973 = n20947 & ~n21972;
  assign n21974 = ~pi752 & ~n21973;
  assign n21975 = ~n21971 & n21974;
  assign n21976 = ~pi164 & n20891;
  assign n21977 = pi164 & n20908;
  assign n21978 = ~pi38 & ~n21977;
  assign n21979 = ~n21976 & n21978;
  assign n21980 = ~pi164 & ~n17280;
  assign n21981 = n20914 & ~n21980;
  assign n21982 = pi752 & ~n21981;
  assign n21983 = ~n21979 & n21982;
  assign n21984 = ~n21975 & ~n21983;
  assign n21985 = pi703 & ~n21984;
  assign n21986 = pi164 & ~n20848;
  assign n21987 = ~pi752 & ~n21986;
  assign n21988 = ~n20849 & n21987;
  assign n21989 = ~pi752 & n20873;
  assign n21990 = pi164 & ~n21989;
  assign n21991 = pi752 & n17399;
  assign n21992 = ~pi703 & ~n21991;
  assign n21993 = ~n21990 & n21992;
  assign n21994 = ~n21988 & n21993;
  assign n21995 = ~n21985 & ~n21994;
  assign n21996 = n10143 & ~n21995;
  assign n21997 = ~pi164 & ~n10143;
  assign n21998 = ~pi832 & ~n21997;
  assign n21999 = ~n21996 & n21998;
  assign po321 = ~n21967 & ~n21999;
  assign n22001 = ~pi774 & pi947;
  assign n22002 = pi687 & n20755;
  assign n22003 = ~n22001 & ~n22002;
  assign n22004 = n2754 & ~n22003;
  assign n22005 = ~pi165 & ~n2754;
  assign n22006 = pi832 & ~n22005;
  assign n22007 = ~n22004 & n22006;
  assign n22008 = ~pi165 & n20929;
  assign n22009 = pi165 & n20940;
  assign n22010 = ~pi38 & ~n22009;
  assign n22011 = ~n22008 & n22010;
  assign n22012 = ~pi165 & ~n20944;
  assign n22013 = n20947 & ~n22012;
  assign n22014 = ~pi774 & ~n22013;
  assign n22015 = ~n22011 & n22014;
  assign n22016 = ~pi165 & n20891;
  assign n22017 = pi165 & n20908;
  assign n22018 = ~pi38 & ~n22017;
  assign n22019 = ~n22016 & n22018;
  assign n22020 = ~pi165 & ~n17280;
  assign n22021 = n20914 & ~n22020;
  assign n22022 = pi774 & ~n22021;
  assign n22023 = ~n22019 & n22022;
  assign n22024 = ~n22015 & ~n22023;
  assign n22025 = pi687 & ~n22024;
  assign n22026 = pi165 & ~n20848;
  assign n22027 = ~pi774 & ~n22026;
  assign n22028 = ~n20849 & n22027;
  assign n22029 = ~pi774 & n20873;
  assign n22030 = pi165 & ~n22029;
  assign n22031 = pi774 & n17399;
  assign n22032 = ~pi687 & ~n22031;
  assign n22033 = ~n22030 & n22032;
  assign n22034 = ~n22028 & n22033;
  assign n22035 = ~n22025 & ~n22034;
  assign n22036 = n10143 & ~n22035;
  assign n22037 = ~pi165 & ~n10143;
  assign n22038 = ~pi832 & ~n22037;
  assign n22039 = ~n22036 & n22038;
  assign po322 = ~n22007 & ~n22039;
  assign n22041 = pi166 & n20879;
  assign n22042 = n20894 & ~n22041;
  assign n22043 = ~n20834 & ~n22042;
  assign n22044 = ~n20862 & ~n22043;
  assign n22045 = pi166 & ~n16518;
  assign n22046 = ~n20864 & ~n22045;
  assign n22047 = n3329 & n22046;
  assign n22048 = ~pi215 & ~n22047;
  assign n22049 = ~n22044 & n22048;
  assign n22050 = pi166 & n20839;
  assign n22051 = n20861 & ~n22050;
  assign n22052 = ~n22049 & n22051;
  assign n22053 = ~pi166 & ~n17153;
  assign n22054 = n21233 & ~n22053;
  assign n22055 = ~pi299 & ~n22054;
  assign n22056 = n3052 & ~n22046;
  assign n22057 = ~pi166 & ~n17175;
  assign n22058 = n21218 & ~n22057;
  assign n22059 = ~n22056 & ~n22058;
  assign n22060 = ~pi223 & ~n22059;
  assign n22061 = n22055 & ~n22060;
  assign n22062 = pi772 & ~n22061;
  assign n22063 = ~n22052 & n22062;
  assign n22064 = ~pi772 & ~n17199;
  assign n22065 = pi166 & n22064;
  assign n22066 = pi39 & ~n22065;
  assign n22067 = ~n22063 & n22066;
  assign n22068 = pi166 & ~n17120;
  assign n22069 = pi772 & pi947;
  assign n22070 = ~pi39 & ~n22069;
  assign n22071 = ~n17121 & ~n22070;
  assign n22072 = ~n22068 & ~n22071;
  assign n22073 = ~pi38 & ~n22072;
  assign n22074 = ~n22067 & n22073;
  assign n22075 = ~pi166 & ~n17397;
  assign n22076 = n17280 & ~n22069;
  assign n22077 = pi38 & ~n22076;
  assign n22078 = ~n22075 & n22077;
  assign n22079 = ~pi727 & ~n22078;
  assign n22080 = ~n22074 & n22079;
  assign n22081 = ~n20931 & ~n22045;
  assign n22082 = n3329 & n22081;
  assign n22083 = ~pi215 & ~n22082;
  assign n22084 = ~n20878 & n22083;
  assign n22085 = ~n22042 & n22084;
  assign n22086 = ~pi166 & ~n17190;
  assign n22087 = n20837 & ~n22086;
  assign n22088 = ~n21261 & n22087;
  assign n22089 = pi299 & ~n22088;
  assign n22090 = ~n22085 & n22089;
  assign n22091 = ~n21252 & ~n22057;
  assign n22092 = ~n3052 & ~n22091;
  assign n22093 = n3052 & n22081;
  assign n22094 = ~pi223 & ~n22093;
  assign n22095 = n3052 & n20864;
  assign n22096 = n22094 & ~n22095;
  assign n22097 = ~n22092 & n22096;
  assign n22098 = ~n6183 & n17153;
  assign n22099 = ~pi166 & ~n22098;
  assign n22100 = n21229 & ~n22099;
  assign n22101 = ~pi299 & ~n22100;
  assign n22102 = ~n22097 & n22101;
  assign n22103 = ~pi772 & ~n22102;
  assign n22104 = ~n22090 & n22103;
  assign n22105 = ~n17186 & n22042;
  assign n22106 = n22083 & ~n22105;
  assign n22107 = pi299 & ~n22087;
  assign n22108 = ~n22106 & n22107;
  assign n22109 = n21221 & ~n22091;
  assign n22110 = n22094 & ~n22109;
  assign n22111 = n22055 & ~n22100;
  assign n22112 = ~n22110 & n22111;
  assign n22113 = pi772 & ~n22112;
  assign n22114 = ~n22108 & n22113;
  assign n22115 = pi39 & ~n22114;
  assign n22116 = ~n22104 & n22115;
  assign n22117 = ~n20906 & n22072;
  assign n22118 = ~pi38 & ~n22117;
  assign n22119 = ~n22116 & n22118;
  assign n22120 = ~pi166 & ~n17280;
  assign n22121 = n21277 & n22070;
  assign n22122 = pi38 & ~n22121;
  assign n22123 = ~n22120 & n22122;
  assign n22124 = pi727 & ~n22123;
  assign n22125 = ~n22119 & n22124;
  assign n22126 = ~n22080 & ~n22125;
  assign n22127 = n10143 & ~n22126;
  assign n22128 = ~pi166 & ~n10143;
  assign n22129 = ~pi832 & ~n22128;
  assign n22130 = ~n22127 & n22129;
  assign n22131 = pi727 & n20755;
  assign n22132 = n2754 & ~n22069;
  assign n22133 = ~n22131 & n22132;
  assign n22134 = ~pi166 & ~n2754;
  assign n22135 = pi832 & ~n22134;
  assign n22136 = ~n22133 & n22135;
  assign po323 = n22130 | n22136;
  assign n22138 = ~pi768 & pi947;
  assign n22139 = pi705 & n20755;
  assign n22140 = ~n22138 & ~n22139;
  assign n22141 = n2754 & ~n22140;
  assign n22142 = ~pi167 & ~n2754;
  assign n22143 = pi832 & ~n22142;
  assign n22144 = ~n22141 & n22143;
  assign n22145 = ~pi167 & n20929;
  assign n22146 = pi167 & n20940;
  assign n22147 = ~pi38 & ~n22146;
  assign n22148 = ~n22145 & n22147;
  assign n22149 = ~pi167 & ~n20944;
  assign n22150 = n20947 & ~n22149;
  assign n22151 = ~pi768 & ~n22150;
  assign n22152 = ~n22148 & n22151;
  assign n22153 = ~pi167 & n20891;
  assign n22154 = pi167 & n20908;
  assign n22155 = ~pi38 & ~n22154;
  assign n22156 = ~n22153 & n22155;
  assign n22157 = ~pi167 & ~n17280;
  assign n22158 = n20914 & ~n22157;
  assign n22159 = pi768 & ~n22158;
  assign n22160 = ~n22156 & n22159;
  assign n22161 = pi705 & ~n22160;
  assign n22162 = ~n22152 & n22161;
  assign n22163 = ~pi167 & ~n20845;
  assign n22164 = pi167 & n20871;
  assign n22165 = ~pi38 & ~n22164;
  assign n22166 = ~n22163 & n22165;
  assign n22167 = ~pi167 & ~n17397;
  assign n22168 = ~n20854 & ~n22167;
  assign n22169 = ~pi768 & ~n22168;
  assign n22170 = ~n22166 & n22169;
  assign n22171 = pi768 & ~n17399;
  assign n22172 = ~pi167 & n22171;
  assign n22173 = ~pi705 & ~n22172;
  assign n22174 = ~n22170 & n22173;
  assign n22175 = n10143 & ~n22174;
  assign n22176 = ~n22162 & n22175;
  assign n22177 = ~pi167 & ~n10143;
  assign n22178 = ~pi832 & ~n22177;
  assign n22179 = ~n22176 & n22178;
  assign po324 = ~n22144 & ~n22179;
  assign n22181 = pi763 & pi947;
  assign n22182 = n2754 & ~n22181;
  assign n22183 = pi699 & n20755;
  assign n22184 = n22182 & ~n22183;
  assign n22185 = pi168 & ~n2754;
  assign n22186 = pi832 & ~n22185;
  assign n22187 = ~n22184 & n22186;
  assign n22188 = ~pi168 & ~n17120;
  assign n22189 = ~pi763 & n17954;
  assign n22190 = ~n20856 & ~n22189;
  assign n22191 = ~n22188 & ~n22190;
  assign n22192 = ~n20906 & n22191;
  assign n22193 = pi168 & ~n17190;
  assign n22194 = n20837 & ~n22193;
  assign n22195 = pi168 & ~n3329;
  assign n22196 = ~n17186 & n22195;
  assign n22197 = ~n17185 & ~n22196;
  assign n22198 = ~pi168 & ~n16518;
  assign n22199 = n20865 & ~n22198;
  assign n22200 = ~n20895 & n22199;
  assign n22201 = ~pi215 & ~n22200;
  assign n22202 = n22197 & n22201;
  assign n22203 = ~n22194 & ~n22202;
  assign n22204 = pi299 & ~n22203;
  assign n22205 = pi168 & ~n20921;
  assign n22206 = ~n20923 & ~n22205;
  assign n22207 = ~n22204 & ~n22206;
  assign n22208 = pi763 & ~n22207;
  assign n22209 = n20897 & ~n22198;
  assign n22210 = ~n20880 & ~n22209;
  assign n22211 = n22197 & n22210;
  assign n22212 = ~pi215 & ~n22211;
  assign n22213 = n20935 & ~n22194;
  assign n22214 = ~n20860 & ~n22213;
  assign n22215 = ~n22212 & n22214;
  assign n22216 = pi299 & ~n22215;
  assign n22217 = ~pi168 & ~n17179;
  assign n22218 = n20903 & ~n22217;
  assign n22219 = ~pi763 & ~n22218;
  assign n22220 = ~n22216 & n22219;
  assign n22221 = pi39 & ~n22220;
  assign n22222 = ~n22208 & n22221;
  assign n22223 = ~n22192 & ~n22222;
  assign n22224 = ~pi38 & ~n22223;
  assign n22225 = ~pi763 & pi947;
  assign n22226 = ~pi39 & ~n22225;
  assign n22227 = n21067 & n22226;
  assign n22228 = ~pi168 & ~n17280;
  assign n22229 = pi38 & ~n22228;
  assign n22230 = ~n22227 & n22229;
  assign n22231 = ~n22224 & ~n22230;
  assign n22232 = pi699 & ~n22231;
  assign n22233 = n20858 & ~n22217;
  assign n22234 = n22197 & ~n22199;
  assign n22235 = n20835 & n22234;
  assign n22236 = n20839 & ~n22193;
  assign n22237 = pi299 & ~n22236;
  assign n22238 = ~n22235 & n22237;
  assign n22239 = pi763 & ~n22238;
  assign n22240 = ~n22233 & n22239;
  assign n22241 = ~pi168 & ~pi763;
  assign n22242 = ~n17199 & n22241;
  assign n22243 = pi39 & ~n22242;
  assign n22244 = ~n22240 & n22243;
  assign n22245 = ~pi38 & ~n22191;
  assign n22246 = ~n22244 & n22245;
  assign n22247 = pi168 & ~n17397;
  assign n22248 = n6234 & n22182;
  assign n22249 = pi38 & ~n22248;
  assign n22250 = ~n22247 & n22249;
  assign n22251 = ~pi699 & ~n22250;
  assign n22252 = ~n22246 & n22251;
  assign n22253 = n20983 & ~n22252;
  assign n22254 = ~n22232 & n22253;
  assign n22255 = ~pi168 & ~n20983;
  assign n22256 = ~pi57 & ~n22255;
  assign n22257 = ~n22254 & n22256;
  assign n22258 = pi57 & pi168;
  assign n22259 = ~pi832 & ~n22258;
  assign n22260 = ~n22257 & n22259;
  assign po325 = n22187 | n22260;
  assign n22262 = pi746 & pi947;
  assign n22263 = n2754 & ~n22262;
  assign n22264 = pi729 & n20755;
  assign n22265 = n22263 & ~n22264;
  assign n22266 = pi169 & ~n2754;
  assign n22267 = pi832 & ~n22266;
  assign n22268 = ~n22265 & n22267;
  assign n22269 = ~pi169 & ~n17120;
  assign n22270 = ~pi746 & n17954;
  assign n22271 = ~n20856 & ~n22270;
  assign n22272 = ~n22269 & ~n22271;
  assign n22273 = ~n20906 & n22272;
  assign n22274 = pi169 & ~n17190;
  assign n22275 = n20837 & ~n22274;
  assign n22276 = pi169 & ~n3329;
  assign n22277 = ~n17186 & n22276;
  assign n22278 = ~n17185 & ~n22277;
  assign n22279 = ~pi169 & ~n16518;
  assign n22280 = n20865 & ~n22279;
  assign n22281 = ~n20895 & n22280;
  assign n22282 = ~pi215 & ~n22281;
  assign n22283 = n22278 & n22282;
  assign n22284 = ~n22275 & ~n22283;
  assign n22285 = pi299 & ~n22284;
  assign n22286 = pi169 & ~n20921;
  assign n22287 = ~n20923 & ~n22286;
  assign n22288 = ~n22285 & ~n22287;
  assign n22289 = pi746 & ~n22288;
  assign n22290 = n20897 & ~n22279;
  assign n22291 = ~n20880 & ~n22290;
  assign n22292 = n22278 & n22291;
  assign n22293 = ~pi215 & ~n22292;
  assign n22294 = n20935 & ~n22275;
  assign n22295 = ~n20860 & ~n22294;
  assign n22296 = ~n22293 & n22295;
  assign n22297 = pi299 & ~n22296;
  assign n22298 = ~pi169 & ~n17179;
  assign n22299 = n20903 & ~n22298;
  assign n22300 = ~pi746 & ~n22299;
  assign n22301 = ~n22297 & n22300;
  assign n22302 = pi39 & ~n22301;
  assign n22303 = ~n22289 & n22302;
  assign n22304 = ~n22273 & ~n22303;
  assign n22305 = ~pi38 & ~n22304;
  assign n22306 = ~pi746 & pi947;
  assign n22307 = ~pi39 & ~n22306;
  assign n22308 = n21067 & n22307;
  assign n22309 = ~pi169 & ~n17280;
  assign n22310 = pi38 & ~n22309;
  assign n22311 = ~n22308 & n22310;
  assign n22312 = ~n22305 & ~n22311;
  assign n22313 = pi729 & ~n22312;
  assign n22314 = n20858 & ~n22298;
  assign n22315 = n22278 & ~n22280;
  assign n22316 = n20835 & n22315;
  assign n22317 = n20839 & ~n22274;
  assign n22318 = pi299 & ~n22317;
  assign n22319 = ~n22316 & n22318;
  assign n22320 = pi746 & ~n22319;
  assign n22321 = ~n22314 & n22320;
  assign n22322 = ~pi169 & ~pi746;
  assign n22323 = ~n17199 & n22322;
  assign n22324 = pi39 & ~n22323;
  assign n22325 = ~n22321 & n22324;
  assign n22326 = ~pi38 & ~n22272;
  assign n22327 = ~n22325 & n22326;
  assign n22328 = pi169 & ~n17397;
  assign n22329 = n6234 & n22263;
  assign n22330 = pi38 & ~n22329;
  assign n22331 = ~n22328 & n22330;
  assign n22332 = ~pi729 & ~n22331;
  assign n22333 = ~n22327 & n22332;
  assign n22334 = n20983 & ~n22333;
  assign n22335 = ~n22313 & n22334;
  assign n22336 = ~pi169 & ~n20983;
  assign n22337 = ~pi57 & ~n22336;
  assign n22338 = ~n22335 & n22337;
  assign n22339 = pi57 & pi169;
  assign n22340 = ~pi832 & ~n22339;
  assign n22341 = ~n22338 & n22340;
  assign po326 = n22268 | n22341;
  assign n22343 = pi730 & n20755;
  assign n22344 = pi748 & pi947;
  assign n22345 = n2754 & ~n22344;
  assign n22346 = ~n22343 & n22345;
  assign n22347 = pi170 & ~n2754;
  assign n22348 = pi832 & ~n22347;
  assign n22349 = ~n22346 & n22348;
  assign n22350 = pi170 & ~n3329;
  assign n22351 = ~n17186 & n22350;
  assign n22352 = ~n17185 & ~n22351;
  assign n22353 = ~pi170 & ~n16518;
  assign n22354 = n20897 & ~n22353;
  assign n22355 = ~n20880 & ~n22354;
  assign n22356 = n22352 & n22355;
  assign n22357 = ~pi215 & ~n22356;
  assign n22358 = pi170 & ~n17190;
  assign n22359 = n20837 & ~n22358;
  assign n22360 = n20935 & ~n22359;
  assign n22361 = ~n20860 & ~n22360;
  assign n22362 = ~n22357 & n22361;
  assign n22363 = pi299 & ~n22362;
  assign n22364 = ~pi170 & ~n17179;
  assign n22365 = ~pi299 & ~n22364;
  assign n22366 = ~n20902 & n22365;
  assign n22367 = ~n22363 & ~n22366;
  assign n22368 = pi39 & ~n22367;
  assign n22369 = ~pi170 & ~n17120;
  assign n22370 = n20907 & ~n22369;
  assign n22371 = ~n22368 & ~n22370;
  assign n22372 = ~pi38 & ~n22371;
  assign n22373 = ~pi170 & ~n17280;
  assign n22374 = n20914 & ~n22373;
  assign n22375 = ~pi748 & ~n22374;
  assign n22376 = ~n22372 & n22375;
  assign n22377 = n20927 & ~n22369;
  assign n22378 = pi170 & ~n20921;
  assign n22379 = ~n20923 & ~n22378;
  assign n22380 = n20865 & ~n22353;
  assign n22381 = ~n20895 & n22380;
  assign n22382 = ~pi215 & ~n22381;
  assign n22383 = n22352 & n22382;
  assign n22384 = ~n22359 & ~n22383;
  assign n22385 = pi299 & ~n22384;
  assign n22386 = pi39 & ~n22385;
  assign n22387 = ~n22379 & n22386;
  assign n22388 = ~n22377 & ~n22387;
  assign n22389 = ~pi38 & ~n22388;
  assign n22390 = n20947 & ~n22373;
  assign n22391 = pi748 & ~n22390;
  assign n22392 = ~n22389 & n22391;
  assign n22393 = pi730 & ~n22392;
  assign n22394 = ~n22376 & n22393;
  assign n22395 = n20856 & ~n22369;
  assign n22396 = n22352 & ~n22380;
  assign n22397 = n20835 & n22396;
  assign n22398 = n20839 & ~n22358;
  assign n22399 = pi299 & ~n22398;
  assign n22400 = ~n22397 & n22399;
  assign n22401 = ~n20857 & n22365;
  assign n22402 = ~n22400 & ~n22401;
  assign n22403 = pi39 & ~n22402;
  assign n22404 = ~n22395 & ~n22403;
  assign n22405 = ~pi38 & ~n22404;
  assign n22406 = ~pi170 & ~n17397;
  assign n22407 = ~n20854 & ~n22406;
  assign n22408 = pi748 & ~n22407;
  assign n22409 = ~n22405 & n22408;
  assign n22410 = ~pi170 & ~pi748;
  assign n22411 = ~n17399 & n22410;
  assign n22412 = ~pi730 & ~n22411;
  assign n22413 = ~n22409 & n22412;
  assign n22414 = n20983 & ~n22413;
  assign n22415 = ~n22394 & n22414;
  assign n22416 = ~pi170 & ~n20983;
  assign n22417 = ~pi57 & ~n22416;
  assign n22418 = ~n22415 & n22417;
  assign n22419 = pi57 & pi170;
  assign n22420 = ~pi832 & ~n22419;
  assign n22421 = ~n22418 & n22420;
  assign po327 = n22349 | n22421;
  assign n22423 = pi764 & pi947;
  assign n22424 = n2754 & ~n22423;
  assign n22425 = pi691 & n20755;
  assign n22426 = n22424 & ~n22425;
  assign n22427 = pi171 & ~n2754;
  assign n22428 = pi832 & ~n22427;
  assign n22429 = ~n22426 & n22428;
  assign n22430 = ~pi171 & ~n17120;
  assign n22431 = ~pi764 & n17954;
  assign n22432 = ~n20856 & ~n22431;
  assign n22433 = ~n22430 & ~n22432;
  assign n22434 = ~n20906 & n22433;
  assign n22435 = pi171 & ~n17190;
  assign n22436 = n20837 & ~n22435;
  assign n22437 = pi171 & ~n3329;
  assign n22438 = ~n17186 & n22437;
  assign n22439 = ~n17185 & ~n22438;
  assign n22440 = ~pi171 & ~n16518;
  assign n22441 = n20865 & ~n22440;
  assign n22442 = ~n20895 & n22441;
  assign n22443 = ~pi215 & ~n22442;
  assign n22444 = n22439 & n22443;
  assign n22445 = ~n22436 & ~n22444;
  assign n22446 = pi299 & ~n22445;
  assign n22447 = pi171 & ~n20921;
  assign n22448 = ~n20923 & ~n22447;
  assign n22449 = ~n22446 & ~n22448;
  assign n22450 = pi764 & ~n22449;
  assign n22451 = n20897 & ~n22440;
  assign n22452 = ~n20880 & ~n22451;
  assign n22453 = n22439 & n22452;
  assign n22454 = ~pi215 & ~n22453;
  assign n22455 = n20935 & ~n22436;
  assign n22456 = ~n20860 & ~n22455;
  assign n22457 = ~n22454 & n22456;
  assign n22458 = pi299 & ~n22457;
  assign n22459 = ~pi171 & ~n17179;
  assign n22460 = n20903 & ~n22459;
  assign n22461 = ~pi764 & ~n22460;
  assign n22462 = ~n22458 & n22461;
  assign n22463 = pi39 & ~n22462;
  assign n22464 = ~n22450 & n22463;
  assign n22465 = ~n22434 & ~n22464;
  assign n22466 = ~pi38 & ~n22465;
  assign n22467 = ~pi764 & pi947;
  assign n22468 = ~pi39 & ~n22467;
  assign n22469 = n21067 & n22468;
  assign n22470 = ~pi171 & ~n17280;
  assign n22471 = pi38 & ~n22470;
  assign n22472 = ~n22469 & n22471;
  assign n22473 = ~n22466 & ~n22472;
  assign n22474 = pi691 & ~n22473;
  assign n22475 = n20858 & ~n22459;
  assign n22476 = n22439 & ~n22441;
  assign n22477 = n20835 & n22476;
  assign n22478 = n20839 & ~n22435;
  assign n22479 = pi299 & ~n22478;
  assign n22480 = ~n22477 & n22479;
  assign n22481 = pi764 & ~n22480;
  assign n22482 = ~n22475 & n22481;
  assign n22483 = ~pi171 & ~pi764;
  assign n22484 = ~n17199 & n22483;
  assign n22485 = pi39 & ~n22484;
  assign n22486 = ~n22482 & n22485;
  assign n22487 = ~pi38 & ~n22433;
  assign n22488 = ~n22486 & n22487;
  assign n22489 = pi171 & ~n17397;
  assign n22490 = n6234 & n22424;
  assign n22491 = pi38 & ~n22490;
  assign n22492 = ~n22489 & n22491;
  assign n22493 = ~pi691 & ~n22492;
  assign n22494 = ~n22488 & n22493;
  assign n22495 = n20983 & ~n22494;
  assign n22496 = ~n22474 & n22495;
  assign n22497 = ~pi171 & ~n20983;
  assign n22498 = ~pi57 & ~n22497;
  assign n22499 = ~n22496 & n22498;
  assign n22500 = pi57 & pi171;
  assign n22501 = ~pi832 & ~n22500;
  assign n22502 = ~n22499 & n22501;
  assign po328 = n22429 | n22502;
  assign n22504 = pi739 & pi947;
  assign n22505 = n2754 & ~n22504;
  assign n22506 = pi690 & n20755;
  assign n22507 = n22505 & ~n22506;
  assign n22508 = pi172 & ~n2754;
  assign n22509 = pi832 & ~n22508;
  assign n22510 = ~n22507 & n22509;
  assign n22511 = n17120 & n22504;
  assign n22512 = ~pi172 & ~n17120;
  assign n22513 = ~pi39 & ~n22512;
  assign n22514 = ~n22511 & n22513;
  assign n22515 = ~n20906 & n22514;
  assign n22516 = pi172 & ~n17190;
  assign n22517 = n20837 & ~n22516;
  assign n22518 = pi172 & ~n3329;
  assign n22519 = ~n17186 & n22518;
  assign n22520 = ~n17185 & ~n22519;
  assign n22521 = ~pi172 & ~n16518;
  assign n22522 = n20865 & ~n22521;
  assign n22523 = ~n20895 & n22522;
  assign n22524 = ~pi215 & ~n22523;
  assign n22525 = n22520 & n22524;
  assign n22526 = ~n22517 & ~n22525;
  assign n22527 = pi299 & ~n22526;
  assign n22528 = pi172 & ~n20921;
  assign n22529 = ~n20923 & ~n22528;
  assign n22530 = ~n22527 & ~n22529;
  assign n22531 = pi739 & ~n22530;
  assign n22532 = n20897 & ~n22521;
  assign n22533 = ~n20880 & ~n22532;
  assign n22534 = n22520 & n22533;
  assign n22535 = ~pi215 & ~n22534;
  assign n22536 = n20935 & ~n22517;
  assign n22537 = ~n20860 & ~n22536;
  assign n22538 = ~n22535 & n22537;
  assign n22539 = pi299 & ~n22538;
  assign n22540 = ~pi172 & ~n17179;
  assign n22541 = n20903 & ~n22540;
  assign n22542 = ~pi739 & ~n22541;
  assign n22543 = ~n22539 & n22542;
  assign n22544 = pi39 & ~n22543;
  assign n22545 = ~n22531 & n22544;
  assign n22546 = ~n22515 & ~n22545;
  assign n22547 = ~pi38 & ~n22546;
  assign n22548 = ~pi739 & pi947;
  assign n22549 = ~pi39 & ~n22548;
  assign n22550 = n21067 & n22549;
  assign n22551 = ~pi172 & ~n17280;
  assign n22552 = pi38 & ~n22551;
  assign n22553 = ~n22550 & n22552;
  assign n22554 = ~n22547 & ~n22553;
  assign n22555 = pi690 & ~n22554;
  assign n22556 = n20858 & ~n22540;
  assign n22557 = n22520 & ~n22522;
  assign n22558 = n20835 & n22557;
  assign n22559 = n20839 & ~n22516;
  assign n22560 = pi299 & ~n22559;
  assign n22561 = ~n22558 & n22560;
  assign n22562 = pi739 & ~n22561;
  assign n22563 = ~n22556 & n22562;
  assign n22564 = ~pi172 & ~pi739;
  assign n22565 = ~n17199 & n22564;
  assign n22566 = pi39 & ~n22565;
  assign n22567 = ~n22563 & n22566;
  assign n22568 = ~pi38 & ~n22514;
  assign n22569 = ~n22567 & n22568;
  assign n22570 = pi172 & ~n17397;
  assign n22571 = n6234 & n22505;
  assign n22572 = pi38 & ~n22571;
  assign n22573 = ~n22570 & n22572;
  assign n22574 = ~pi690 & ~n22573;
  assign n22575 = ~n22569 & n22574;
  assign n22576 = n20983 & ~n22575;
  assign n22577 = ~n22555 & n22576;
  assign n22578 = ~pi172 & ~n20983;
  assign n22579 = ~pi57 & ~n22578;
  assign n22580 = ~n22577 & n22579;
  assign n22581 = pi57 & pi172;
  assign n22582 = ~pi832 & ~n22581;
  assign n22583 = ~n22580 & n22582;
  assign po329 = n22510 | n22583;
  assign n22585 = ~pi173 & ~n17406;
  assign n22586 = n17539 & ~n22585;
  assign n22587 = ~pi723 & n3267;
  assign n22588 = n22585 & ~n22587;
  assign n22589 = pi173 & ~n17976;
  assign n22590 = ~pi38 & ~n22589;
  assign n22591 = n3267 & ~n22590;
  assign n22592 = ~pi173 & n17972;
  assign n22593 = ~n22591 & ~n22592;
  assign n22594 = ~pi173 & ~n17280;
  assign n22595 = n17392 & ~n22594;
  assign n22596 = ~pi723 & ~n22595;
  assign n22597 = ~n22593 & n22596;
  assign n22598 = ~n22588 & ~n22597;
  assign n22599 = ~pi778 & n22598;
  assign n22600 = pi625 & ~n22598;
  assign n22601 = ~pi625 & n22585;
  assign n22602 = pi1153 & ~n22601;
  assign n22603 = ~n22600 & n22602;
  assign n22604 = ~pi625 & ~n22598;
  assign n22605 = pi625 & n22585;
  assign n22606 = ~pi1153 & ~n22605;
  assign n22607 = ~n22604 & n22606;
  assign n22608 = ~n22603 & ~n22607;
  assign n22609 = pi778 & ~n22608;
  assign n22610 = ~n22599 & ~n22609;
  assign n22611 = ~n17466 & ~n22610;
  assign n22612 = n17466 & ~n22585;
  assign n22613 = ~n22611 & ~n22612;
  assign n22614 = ~n17503 & n22613;
  assign n22615 = n17503 & n22585;
  assign n22616 = ~n22614 & ~n22615;
  assign n22617 = ~n17539 & n22616;
  assign n22618 = ~n22586 & ~n22617;
  assign n22619 = ~n17582 & n22618;
  assign n22620 = n17582 & n22585;
  assign n22621 = ~n22619 & ~n22620;
  assign n22622 = ~pi792 & n22621;
  assign n22623 = pi628 & ~n22621;
  assign n22624 = ~pi628 & n22585;
  assign n22625 = pi1156 & ~n22624;
  assign n22626 = ~n22623 & n22625;
  assign n22627 = ~pi628 & ~n22621;
  assign n22628 = pi628 & n22585;
  assign n22629 = ~pi1156 & ~n22628;
  assign n22630 = ~n22627 & n22629;
  assign n22631 = ~n22626 & ~n22630;
  assign n22632 = pi792 & ~n22631;
  assign n22633 = ~n22622 & ~n22632;
  assign n22634 = ~pi647 & ~n22633;
  assign n22635 = pi647 & ~n22585;
  assign n22636 = ~n22634 & ~n22635;
  assign n22637 = ~pi1157 & n22636;
  assign n22638 = pi647 & ~n22633;
  assign n22639 = ~pi647 & ~n22585;
  assign n22640 = ~n22638 & ~n22639;
  assign n22641 = pi1157 & n22640;
  assign n22642 = ~n22637 & ~n22641;
  assign n22643 = pi787 & ~n22642;
  assign n22644 = ~pi787 & n22633;
  assign n22645 = ~n22643 & ~n22644;
  assign n22646 = ~pi644 & ~n22645;
  assign n22647 = pi715 & ~n22646;
  assign n22648 = pi173 & ~n3267;
  assign n22649 = ~pi173 & ~n17201;
  assign n22650 = pi745 & ~n22649;
  assign n22651 = pi173 & ~n17275;
  assign n22652 = ~pi173 & ~pi745;
  assign n22653 = n17242 & n22652;
  assign n22654 = ~n22651 & ~n22653;
  assign n22655 = ~n22650 & n22654;
  assign n22656 = ~pi38 & ~n22655;
  assign n22657 = ~pi745 & n17282;
  assign n22658 = pi38 & ~n22594;
  assign n22659 = ~n22657 & n22658;
  assign n22660 = ~n22656 & ~n22659;
  assign n22661 = n3267 & ~n22660;
  assign n22662 = ~n22648 & ~n22661;
  assign n22663 = ~n17438 & ~n22662;
  assign n22664 = n17438 & ~n22585;
  assign n22665 = ~n22663 & ~n22664;
  assign n22666 = ~pi785 & ~n22665;
  assign n22667 = ~n17439 & ~n22585;
  assign n22668 = pi609 & n22663;
  assign n22669 = ~n22667 & ~n22668;
  assign n22670 = pi1155 & ~n22669;
  assign n22671 = ~n17451 & ~n22585;
  assign n22672 = ~pi609 & n22663;
  assign n22673 = ~n22671 & ~n22672;
  assign n22674 = ~pi1155 & ~n22673;
  assign n22675 = ~n22670 & ~n22674;
  assign n22676 = pi785 & ~n22675;
  assign n22677 = ~n22666 & ~n22676;
  assign n22678 = ~pi781 & ~n22677;
  assign n22679 = pi618 & n22677;
  assign n22680 = ~pi618 & n22585;
  assign n22681 = pi1154 & ~n22680;
  assign n22682 = ~n22679 & n22681;
  assign n22683 = ~pi618 & n22677;
  assign n22684 = pi618 & n22585;
  assign n22685 = ~pi1154 & ~n22684;
  assign n22686 = ~n22683 & n22685;
  assign n22687 = ~n22682 & ~n22686;
  assign n22688 = pi781 & ~n22687;
  assign n22689 = ~n22678 & ~n22688;
  assign n22690 = ~pi789 & ~n22689;
  assign n22691 = pi619 & n22689;
  assign n22692 = ~pi619 & n22585;
  assign n22693 = pi1159 & ~n22692;
  assign n22694 = ~n22691 & n22693;
  assign n22695 = ~pi619 & n22689;
  assign n22696 = pi619 & n22585;
  assign n22697 = ~pi1159 & ~n22696;
  assign n22698 = ~n22695 & n22697;
  assign n22699 = ~n22694 & ~n22698;
  assign n22700 = pi789 & ~n22699;
  assign n22701 = ~n22690 & ~n22700;
  assign n22702 = ~pi788 & ~n22701;
  assign n22703 = pi626 & n22701;
  assign n22704 = ~pi626 & n22585;
  assign n22705 = pi1158 & ~n22704;
  assign n22706 = ~n22703 & n22705;
  assign n22707 = ~pi626 & n22701;
  assign n22708 = pi626 & n22585;
  assign n22709 = ~pi1158 & ~n22708;
  assign n22710 = ~n22707 & n22709;
  assign n22711 = ~n22706 & ~n22710;
  assign n22712 = pi788 & ~n22711;
  assign n22713 = ~n22702 & ~n22712;
  assign n22714 = ~n17610 & n22713;
  assign n22715 = n17610 & n22585;
  assign n22716 = ~n22714 & ~n22715;
  assign n22717 = ~n17652 & ~n22716;
  assign n22718 = n17652 & n22585;
  assign n22719 = ~n22717 & ~n22718;
  assign n22720 = pi644 & ~n22719;
  assign n22721 = ~pi644 & n22585;
  assign n22722 = ~pi715 & ~n22721;
  assign n22723 = ~n22720 & n22722;
  assign n22724 = pi1160 & ~n22723;
  assign n22725 = ~n22647 & n22724;
  assign n22726 = ~n20398 & n22716;
  assign n22727 = n17650 & ~n22636;
  assign n22728 = n17649 & ~n22640;
  assign n22729 = ~n22727 & ~n22728;
  assign n22730 = ~n22726 & n22729;
  assign n22731 = pi787 & ~n22730;
  assign n22732 = ~n20409 & ~n22713;
  assign n22733 = ~pi629 & n22626;
  assign n22734 = pi629 & n22630;
  assign n22735 = ~n22733 & ~n22734;
  assign n22736 = ~n22732 & n22735;
  assign n22737 = pi792 & ~n22736;
  assign n22738 = pi723 & n22660;
  assign n22739 = ~pi173 & n16687;
  assign n22740 = pi173 & n16799;
  assign n22741 = pi745 & ~n22740;
  assign n22742 = ~n22739 & n22741;
  assign n22743 = pi173 & n16879;
  assign n22744 = ~pi173 & ~n16944;
  assign n22745 = ~pi745 & ~n22744;
  assign n22746 = ~n22743 & n22745;
  assign n22747 = pi39 & ~n22746;
  assign n22748 = ~n22742 & n22747;
  assign n22749 = ~pi173 & ~n17088;
  assign n22750 = pi173 & ~n17059;
  assign n22751 = pi745 & ~n22750;
  assign n22752 = ~n22749 & n22751;
  assign n22753 = ~pi173 & n17092;
  assign n22754 = pi173 & n17094;
  assign n22755 = ~pi745 & ~n22754;
  assign n22756 = ~n22753 & n22755;
  assign n22757 = ~n22752 & ~n22756;
  assign n22758 = ~pi39 & ~n22757;
  assign n22759 = ~pi38 & ~n22758;
  assign n22760 = ~n22748 & n22759;
  assign n22761 = ~pi745 & ~n16905;
  assign n22762 = n19230 & ~n22761;
  assign n22763 = ~pi173 & ~n22762;
  assign n22764 = ~pi745 & n16784;
  assign n22765 = ~n16787 & ~n22764;
  assign n22766 = pi173 & ~n22765;
  assign n22767 = n6234 & n22766;
  assign n22768 = pi38 & ~n22767;
  assign n22769 = ~n22763 & n22768;
  assign n22770 = ~pi723 & ~n22769;
  assign n22771 = ~n22760 & n22770;
  assign n22772 = n3267 & ~n22771;
  assign n22773 = ~n22738 & n22772;
  assign n22774 = ~n22648 & ~n22773;
  assign n22775 = ~pi625 & n22774;
  assign n22776 = pi625 & n22662;
  assign n22777 = ~pi1153 & ~n22776;
  assign n22778 = ~n22775 & n22777;
  assign n22779 = ~pi608 & ~n22603;
  assign n22780 = ~n22778 & n22779;
  assign n22781 = pi625 & n22774;
  assign n22782 = ~pi625 & n22662;
  assign n22783 = pi1153 & ~n22782;
  assign n22784 = ~n22781 & n22783;
  assign n22785 = pi608 & ~n22607;
  assign n22786 = ~n22784 & n22785;
  assign n22787 = ~n22780 & ~n22786;
  assign n22788 = pi778 & ~n22787;
  assign n22789 = ~pi778 & n22774;
  assign n22790 = ~n22788 & ~n22789;
  assign n22791 = ~pi609 & ~n22790;
  assign n22792 = pi609 & n22610;
  assign n22793 = ~pi1155 & ~n22792;
  assign n22794 = ~n22791 & n22793;
  assign n22795 = ~pi660 & ~n22670;
  assign n22796 = ~n22794 & n22795;
  assign n22797 = pi609 & ~n22790;
  assign n22798 = ~pi609 & n22610;
  assign n22799 = pi1155 & ~n22798;
  assign n22800 = ~n22797 & n22799;
  assign n22801 = pi660 & ~n22674;
  assign n22802 = ~n22800 & n22801;
  assign n22803 = ~n22796 & ~n22802;
  assign n22804 = pi785 & ~n22803;
  assign n22805 = ~pi785 & ~n22790;
  assign n22806 = ~n22804 & ~n22805;
  assign n22807 = ~pi618 & ~n22806;
  assign n22808 = pi618 & n22613;
  assign n22809 = ~pi1154 & ~n22808;
  assign n22810 = ~n22807 & n22809;
  assign n22811 = ~pi627 & ~n22682;
  assign n22812 = ~n22810 & n22811;
  assign n22813 = pi618 & ~n22806;
  assign n22814 = ~pi618 & n22613;
  assign n22815 = pi1154 & ~n22814;
  assign n22816 = ~n22813 & n22815;
  assign n22817 = pi627 & ~n22686;
  assign n22818 = ~n22816 & n22817;
  assign n22819 = ~n22812 & ~n22818;
  assign n22820 = pi781 & ~n22819;
  assign n22821 = ~pi781 & ~n22806;
  assign n22822 = ~n22820 & ~n22821;
  assign n22823 = pi619 & ~n22822;
  assign n22824 = ~pi619 & ~n22616;
  assign n22825 = pi1159 & ~n22824;
  assign n22826 = ~n22823 & n22825;
  assign n22827 = pi648 & ~n22698;
  assign n22828 = ~n22826 & n22827;
  assign n22829 = ~pi619 & ~n22822;
  assign n22830 = pi619 & ~n22616;
  assign n22831 = ~pi1159 & ~n22830;
  assign n22832 = ~n22829 & n22831;
  assign n22833 = ~pi648 & ~n22694;
  assign n22834 = ~n22832 & n22833;
  assign n22835 = pi789 & ~n22834;
  assign n22836 = ~n22828 & n22835;
  assign n22837 = ~pi789 & n22822;
  assign n22838 = n17817 & ~n22837;
  assign n22839 = ~n22836 & n22838;
  assign n22840 = n17704 & n22618;
  assign n22841 = ~n17581 & n22711;
  assign n22842 = ~n22840 & ~n22841;
  assign n22843 = pi788 & ~n22842;
  assign n22844 = ~n20205 & ~n22843;
  assign n22845 = ~n22839 & n22844;
  assign n22846 = ~n22737 & ~n22845;
  assign n22847 = n20207 & ~n22846;
  assign n22848 = ~n22731 & ~n22847;
  assign n22849 = ~pi644 & n22848;
  assign n22850 = pi644 & ~n22645;
  assign n22851 = ~pi715 & ~n22850;
  assign n22852 = ~n22849 & n22851;
  assign n22853 = ~pi644 & ~n22719;
  assign n22854 = pi644 & n22585;
  assign n22855 = pi715 & ~n22854;
  assign n22856 = ~n22853 & n22855;
  assign n22857 = ~pi1160 & ~n22856;
  assign n22858 = ~n22852 & n22857;
  assign n22859 = ~n22725 & ~n22858;
  assign n22860 = pi790 & ~n22859;
  assign n22861 = pi644 & n22724;
  assign n22862 = pi790 & ~n22861;
  assign n22863 = n22848 & ~n22862;
  assign n22864 = ~n22860 & ~n22863;
  assign n22865 = ~po1038 & ~n22864;
  assign n22866 = ~pi173 & po1038;
  assign n22867 = ~pi832 & ~n22866;
  assign n22868 = ~n22865 & n22867;
  assign n22869 = ~pi173 & ~n2754;
  assign n22870 = ~n22764 & ~n22869;
  assign n22871 = ~n17706 & ~n22870;
  assign n22872 = ~pi785 & ~n22871;
  assign n22873 = n17451 & n22764;
  assign n22874 = n22871 & ~n22873;
  assign n22875 = pi1155 & ~n22874;
  assign n22876 = ~pi1155 & ~n22869;
  assign n22877 = ~n22873 & n22876;
  assign n22878 = ~n22875 & ~n22877;
  assign n22879 = pi785 & ~n22878;
  assign n22880 = ~n22872 & ~n22879;
  assign n22881 = ~pi781 & ~n22880;
  assign n22882 = ~n17721 & n22880;
  assign n22883 = pi1154 & ~n22882;
  assign n22884 = ~n17724 & n22880;
  assign n22885 = ~pi1154 & ~n22884;
  assign n22886 = ~n22883 & ~n22885;
  assign n22887 = pi781 & ~n22886;
  assign n22888 = ~n22881 & ~n22887;
  assign n22889 = ~pi789 & ~n22888;
  assign n22890 = ~pi619 & n2754;
  assign n22891 = n22888 & ~n22890;
  assign n22892 = pi1159 & ~n22891;
  assign n22893 = pi619 & n2754;
  assign n22894 = n22888 & ~n22893;
  assign n22895 = ~pi1159 & ~n22894;
  assign n22896 = ~n22892 & ~n22895;
  assign n22897 = pi789 & ~n22896;
  assign n22898 = ~n22889 & ~n22897;
  assign n22899 = ~pi788 & ~n22898;
  assign n22900 = pi626 & n22898;
  assign n22901 = ~pi626 & n22869;
  assign n22902 = pi1158 & ~n22901;
  assign n22903 = ~n22900 & n22902;
  assign n22904 = ~pi626 & n22898;
  assign n22905 = pi626 & n22869;
  assign n22906 = ~pi1158 & ~n22905;
  assign n22907 = ~n22904 & n22906;
  assign n22908 = ~n22903 & ~n22907;
  assign n22909 = pi788 & ~n22908;
  assign n22910 = ~n22899 & ~n22909;
  assign n22911 = ~n17610 & n22910;
  assign n22912 = n17610 & n22869;
  assign n22913 = ~n22911 & ~n22912;
  assign n22914 = ~n20398 & n22913;
  assign n22915 = ~pi723 & n16786;
  assign n22916 = ~n22869 & ~n22915;
  assign n22917 = ~pi778 & ~n22916;
  assign n22918 = ~pi625 & n22915;
  assign n22919 = ~n22916 & ~n22918;
  assign n22920 = pi1153 & ~n22919;
  assign n22921 = ~pi1153 & ~n22869;
  assign n22922 = ~n22918 & n22921;
  assign n22923 = pi778 & ~n22922;
  assign n22924 = ~n22920 & n22923;
  assign n22925 = ~n22917 & ~n22924;
  assign n22926 = ~n17692 & ~n22925;
  assign n22927 = ~n17694 & n22926;
  assign n22928 = ~n17696 & n22927;
  assign n22929 = ~n17828 & n22928;
  assign n22930 = ~n17859 & n22929;
  assign n22931 = ~pi647 & n22930;
  assign n22932 = pi647 & n22869;
  assign n22933 = ~pi1157 & ~n22932;
  assign n22934 = ~n22931 & n22933;
  assign n22935 = pi647 & ~n22930;
  assign n22936 = ~pi647 & ~n22869;
  assign n22937 = ~n22935 & ~n22936;
  assign n22938 = pi1157 & ~n22937;
  assign n22939 = ~n22934 & ~n22938;
  assign n22940 = ~n17651 & ~n22939;
  assign n22941 = ~n22914 & ~n22940;
  assign n22942 = pi787 & ~n22941;
  assign n22943 = n17704 & n22928;
  assign n22944 = ~n17581 & n22908;
  assign n22945 = ~n22943 & ~n22944;
  assign n22946 = pi788 & ~n22945;
  assign n22947 = ~n16521 & ~n22916;
  assign n22948 = pi625 & n22947;
  assign n22949 = n22870 & ~n22947;
  assign n22950 = ~n22948 & ~n22949;
  assign n22951 = n22921 & ~n22950;
  assign n22952 = ~pi608 & ~n22920;
  assign n22953 = ~n22951 & n22952;
  assign n22954 = pi1153 & n22870;
  assign n22955 = ~n22948 & n22954;
  assign n22956 = pi608 & ~n22922;
  assign n22957 = ~n22955 & n22956;
  assign n22958 = ~n22953 & ~n22957;
  assign n22959 = pi778 & ~n22958;
  assign n22960 = ~pi778 & ~n22949;
  assign n22961 = ~n22959 & ~n22960;
  assign n22962 = ~pi609 & ~n22961;
  assign n22963 = pi609 & ~n22925;
  assign n22964 = ~pi1155 & ~n22963;
  assign n22965 = ~n22962 & n22964;
  assign n22966 = ~pi660 & ~n22875;
  assign n22967 = ~n22965 & n22966;
  assign n22968 = pi609 & ~n22961;
  assign n22969 = ~pi609 & ~n22925;
  assign n22970 = pi1155 & ~n22969;
  assign n22971 = ~n22968 & n22970;
  assign n22972 = pi660 & ~n22877;
  assign n22973 = ~n22971 & n22972;
  assign n22974 = ~n22967 & ~n22973;
  assign n22975 = pi785 & ~n22974;
  assign n22976 = ~pi785 & ~n22961;
  assign n22977 = ~n22975 & ~n22976;
  assign n22978 = ~pi618 & ~n22977;
  assign n22979 = pi618 & n22926;
  assign n22980 = ~pi1154 & ~n22979;
  assign n22981 = ~n22978 & n22980;
  assign n22982 = ~pi627 & ~n22883;
  assign n22983 = ~n22981 & n22982;
  assign n22984 = pi618 & ~n22977;
  assign n22985 = ~pi618 & n22926;
  assign n22986 = pi1154 & ~n22985;
  assign n22987 = ~n22984 & n22986;
  assign n22988 = pi627 & ~n22885;
  assign n22989 = ~n22987 & n22988;
  assign n22990 = ~n22983 & ~n22989;
  assign n22991 = pi781 & ~n22990;
  assign n22992 = ~pi781 & ~n22977;
  assign n22993 = ~n22991 & ~n22992;
  assign n22994 = pi619 & ~n22993;
  assign n22995 = ~pi619 & n22927;
  assign n22996 = pi1159 & ~n22995;
  assign n22997 = ~n22994 & n22996;
  assign n22998 = pi648 & ~n22895;
  assign n22999 = ~n22997 & n22998;
  assign n23000 = ~pi619 & ~n22993;
  assign n23001 = pi619 & n22927;
  assign n23002 = ~pi1159 & ~n23001;
  assign n23003 = ~n23000 & n23002;
  assign n23004 = ~pi648 & ~n22892;
  assign n23005 = ~n23003 & n23004;
  assign n23006 = pi789 & ~n23005;
  assign n23007 = ~n22999 & n23006;
  assign n23008 = ~pi789 & n22993;
  assign n23009 = n17817 & ~n23008;
  assign n23010 = ~n23007 & n23009;
  assign n23011 = ~n22946 & ~n23010;
  assign n23012 = ~n20205 & ~n23011;
  assign n23013 = n17856 & n22910;
  assign n23014 = n20693 & n22929;
  assign n23015 = ~n23013 & ~n23014;
  assign n23016 = ~pi629 & ~n23015;
  assign n23017 = n20697 & n22929;
  assign n23018 = n17855 & n22910;
  assign n23019 = ~n23017 & ~n23018;
  assign n23020 = pi629 & ~n23019;
  assign n23021 = ~n23016 & ~n23020;
  assign n23022 = pi792 & ~n23021;
  assign n23023 = n20207 & ~n23022;
  assign n23024 = ~n23012 & n23023;
  assign n23025 = ~n22942 & ~n23024;
  assign n23026 = pi644 & n23025;
  assign n23027 = ~pi787 & ~n22930;
  assign n23028 = pi787 & ~n22939;
  assign n23029 = ~n23027 & ~n23028;
  assign n23030 = ~pi644 & n23029;
  assign n23031 = pi715 & ~n23030;
  assign n23032 = ~n23026 & n23031;
  assign n23033 = ~n17652 & ~n22913;
  assign n23034 = n17652 & n22869;
  assign n23035 = ~n23033 & ~n23034;
  assign n23036 = pi644 & ~n23035;
  assign n23037 = ~pi644 & n22869;
  assign n23038 = ~pi715 & ~n23037;
  assign n23039 = ~n23036 & n23038;
  assign n23040 = pi1160 & ~n23039;
  assign n23041 = ~n23032 & n23040;
  assign n23042 = ~pi644 & n23025;
  assign n23043 = pi644 & n23029;
  assign n23044 = ~pi715 & ~n23043;
  assign n23045 = ~n23042 & n23044;
  assign n23046 = ~pi644 & ~n23035;
  assign n23047 = pi644 & n22869;
  assign n23048 = pi715 & ~n23047;
  assign n23049 = ~n23046 & n23048;
  assign n23050 = ~pi1160 & ~n23049;
  assign n23051 = ~n23045 & n23050;
  assign n23052 = ~n23041 & ~n23051;
  assign n23053 = pi790 & ~n23052;
  assign n23054 = ~pi790 & n23025;
  assign n23055 = pi832 & ~n23054;
  assign n23056 = ~n23053 & n23055;
  assign po330 = ~n22868 & ~n23056;
  assign n23058 = pi174 & ~n3267;
  assign n23059 = pi174 & ~n16687;
  assign n23060 = ~pi174 & ~n16799;
  assign n23061 = ~pi759 & ~n23060;
  assign n23062 = ~n23059 & n23061;
  assign n23063 = ~pi174 & ~n16879;
  assign n23064 = pi174 & n16944;
  assign n23065 = pi759 & ~n23064;
  assign n23066 = ~n23063 & n23065;
  assign n23067 = pi39 & ~n23066;
  assign n23068 = ~n23062 & n23067;
  assign n23069 = pi174 & ~n17088;
  assign n23070 = ~pi174 & ~n17059;
  assign n23071 = ~pi759 & ~n23070;
  assign n23072 = ~n23069 & n23071;
  assign n23073 = pi174 & n17092;
  assign n23074 = ~pi174 & n17094;
  assign n23075 = pi759 & ~n23074;
  assign n23076 = ~n23073 & n23075;
  assign n23077 = ~pi39 & ~n23076;
  assign n23078 = ~n23072 & n23077;
  assign n23079 = ~pi38 & ~n23078;
  assign n23080 = ~n23068 & n23079;
  assign n23081 = pi759 & n16521;
  assign n23082 = n17280 & ~n23081;
  assign n23083 = ~pi174 & ~n17280;
  assign n23084 = pi38 & ~n23083;
  assign n23085 = ~n23082 & n23084;
  assign n23086 = pi696 & ~n19243;
  assign n23087 = ~n23085 & n23086;
  assign n23088 = ~n23080 & n23087;
  assign n23089 = pi759 & n17240;
  assign n23090 = ~n21299 & ~n23089;
  assign n23091 = pi39 & ~n23090;
  assign n23092 = pi759 & n17042;
  assign n23093 = ~pi759 & n17120;
  assign n23094 = ~pi39 & ~n23093;
  assign n23095 = ~n23092 & n23094;
  assign n23096 = ~n23091 & ~n23095;
  assign n23097 = pi174 & ~n23096;
  assign n23098 = ~pi174 & pi759;
  assign n23099 = n17275 & n23098;
  assign n23100 = ~n23097 & ~n23099;
  assign n23101 = ~pi38 & ~n23100;
  assign n23102 = ~n23085 & ~n23101;
  assign n23103 = n3267 & ~n23102;
  assign n23104 = pi696 & n3267;
  assign n23105 = ~n23103 & ~n23104;
  assign n23106 = ~n23088 & ~n23105;
  assign n23107 = ~n23058 & ~n23106;
  assign n23108 = ~pi625 & n23107;
  assign n23109 = ~n23058 & ~n23103;
  assign n23110 = pi625 & n23109;
  assign n23111 = ~pi1153 & ~n23110;
  assign n23112 = ~n23108 & n23111;
  assign n23113 = pi174 & ~n17406;
  assign n23114 = ~n23104 & ~n23113;
  assign n23115 = pi174 & ~n17972;
  assign n23116 = ~pi174 & n17976;
  assign n23117 = ~pi38 & ~n23116;
  assign n23118 = ~n23115 & n23117;
  assign n23119 = n19802 & ~n23083;
  assign n23120 = n23104 & ~n23119;
  assign n23121 = ~n23118 & n23120;
  assign n23122 = ~n23114 & ~n23121;
  assign n23123 = pi625 & ~n23122;
  assign n23124 = ~pi625 & ~n23113;
  assign n23125 = pi1153 & ~n23124;
  assign n23126 = ~n23123 & n23125;
  assign n23127 = ~pi608 & ~n23126;
  assign n23128 = ~n23112 & n23127;
  assign n23129 = pi625 & n23107;
  assign n23130 = ~pi625 & n23109;
  assign n23131 = pi1153 & ~n23130;
  assign n23132 = ~n23129 & n23131;
  assign n23133 = ~pi625 & ~n23122;
  assign n23134 = pi625 & ~n23113;
  assign n23135 = ~pi1153 & ~n23134;
  assign n23136 = ~n23133 & n23135;
  assign n23137 = pi608 & ~n23136;
  assign n23138 = ~n23132 & n23137;
  assign n23139 = ~n23128 & ~n23138;
  assign n23140 = pi778 & ~n23139;
  assign n23141 = ~pi778 & n23107;
  assign n23142 = ~n23140 & ~n23141;
  assign n23143 = ~pi609 & ~n23142;
  assign n23144 = ~pi778 & n23122;
  assign n23145 = ~n23126 & ~n23136;
  assign n23146 = pi778 & ~n23145;
  assign n23147 = ~n23144 & ~n23146;
  assign n23148 = pi609 & n23147;
  assign n23149 = ~pi1155 & ~n23148;
  assign n23150 = ~n23143 & n23149;
  assign n23151 = n17438 & ~n23113;
  assign n23152 = ~n17438 & n23109;
  assign n23153 = ~n23151 & ~n23152;
  assign n23154 = pi609 & ~n23153;
  assign n23155 = ~pi609 & ~n23113;
  assign n23156 = pi1155 & ~n23155;
  assign n23157 = ~n23154 & n23156;
  assign n23158 = ~pi660 & ~n23157;
  assign n23159 = ~n23150 & n23158;
  assign n23160 = pi609 & ~n23142;
  assign n23161 = ~pi609 & n23147;
  assign n23162 = pi1155 & ~n23161;
  assign n23163 = ~n23160 & n23162;
  assign n23164 = ~pi609 & ~n23153;
  assign n23165 = pi609 & ~n23113;
  assign n23166 = ~pi1155 & ~n23165;
  assign n23167 = ~n23164 & n23166;
  assign n23168 = pi660 & ~n23167;
  assign n23169 = ~n23163 & n23168;
  assign n23170 = ~n23159 & ~n23169;
  assign n23171 = pi785 & ~n23170;
  assign n23172 = ~pi785 & ~n23142;
  assign n23173 = ~n23171 & ~n23172;
  assign n23174 = ~pi618 & ~n23173;
  assign n23175 = n17466 & ~n23113;
  assign n23176 = ~n17466 & n23147;
  assign n23177 = ~n23175 & ~n23176;
  assign n23178 = pi618 & ~n23177;
  assign n23179 = ~pi1154 & ~n23178;
  assign n23180 = ~n23174 & n23179;
  assign n23181 = ~pi785 & n23153;
  assign n23182 = ~n23157 & ~n23167;
  assign n23183 = pi785 & ~n23182;
  assign n23184 = ~n23181 & ~n23183;
  assign n23185 = pi618 & n23184;
  assign n23186 = ~pi618 & ~n23113;
  assign n23187 = pi1154 & ~n23186;
  assign n23188 = ~n23185 & n23187;
  assign n23189 = ~pi627 & ~n23188;
  assign n23190 = ~n23180 & n23189;
  assign n23191 = pi618 & ~n23173;
  assign n23192 = ~pi618 & ~n23177;
  assign n23193 = pi1154 & ~n23192;
  assign n23194 = ~n23191 & n23193;
  assign n23195 = ~pi618 & n23184;
  assign n23196 = pi618 & ~n23113;
  assign n23197 = ~pi1154 & ~n23196;
  assign n23198 = ~n23195 & n23197;
  assign n23199 = pi627 & ~n23198;
  assign n23200 = ~n23194 & n23199;
  assign n23201 = ~n23190 & ~n23200;
  assign n23202 = pi781 & ~n23201;
  assign n23203 = ~pi781 & ~n23173;
  assign n23204 = ~n23202 & ~n23203;
  assign n23205 = ~pi619 & ~n23204;
  assign n23206 = ~n17503 & n23177;
  assign n23207 = n17503 & n23113;
  assign n23208 = ~n23206 & ~n23207;
  assign n23209 = pi619 & n23208;
  assign n23210 = ~pi1159 & ~n23209;
  assign n23211 = ~n23205 & n23210;
  assign n23212 = ~pi781 & ~n23184;
  assign n23213 = ~n23188 & ~n23198;
  assign n23214 = pi781 & ~n23213;
  assign n23215 = ~n23212 & ~n23214;
  assign n23216 = pi619 & n23215;
  assign n23217 = ~pi619 & ~n23113;
  assign n23218 = pi1159 & ~n23217;
  assign n23219 = ~n23216 & n23218;
  assign n23220 = ~pi648 & ~n23219;
  assign n23221 = ~n23211 & n23220;
  assign n23222 = pi619 & ~n23204;
  assign n23223 = ~pi619 & n23208;
  assign n23224 = pi1159 & ~n23223;
  assign n23225 = ~n23222 & n23224;
  assign n23226 = ~pi619 & n23215;
  assign n23227 = pi619 & ~n23113;
  assign n23228 = ~pi1159 & ~n23227;
  assign n23229 = ~n23226 & n23228;
  assign n23230 = pi648 & ~n23229;
  assign n23231 = ~n23225 & n23230;
  assign n23232 = ~n23221 & ~n23231;
  assign n23233 = pi789 & ~n23232;
  assign n23234 = ~pi789 & ~n23204;
  assign n23235 = ~n23233 & ~n23234;
  assign n23236 = ~pi788 & n23235;
  assign n23237 = ~pi626 & n23235;
  assign n23238 = n17539 & ~n23113;
  assign n23239 = ~n17539 & n23208;
  assign n23240 = ~n23238 & ~n23239;
  assign n23241 = pi626 & n23240;
  assign n23242 = ~pi641 & ~n23241;
  assign n23243 = ~n23237 & n23242;
  assign n23244 = ~pi789 & ~n23215;
  assign n23245 = ~n23219 & ~n23229;
  assign n23246 = pi789 & ~n23245;
  assign n23247 = ~n23244 & ~n23246;
  assign n23248 = ~pi626 & ~n23247;
  assign n23249 = pi626 & n23113;
  assign n23250 = pi641 & ~n23249;
  assign n23251 = ~n23248 & n23250;
  assign n23252 = ~pi1158 & ~n23251;
  assign n23253 = ~n23243 & n23252;
  assign n23254 = pi626 & n23235;
  assign n23255 = ~pi626 & n23240;
  assign n23256 = pi641 & ~n23255;
  assign n23257 = ~n23254 & n23256;
  assign n23258 = pi626 & ~n23247;
  assign n23259 = ~pi626 & n23113;
  assign n23260 = ~pi641 & ~n23259;
  assign n23261 = ~n23258 & n23260;
  assign n23262 = pi1158 & ~n23261;
  assign n23263 = ~n23257 & n23262;
  assign n23264 = ~n23253 & ~n23263;
  assign n23265 = pi788 & ~n23264;
  assign n23266 = ~n23236 & ~n23265;
  assign n23267 = ~pi628 & n23266;
  assign n23268 = ~n17816 & ~n23247;
  assign n23269 = n17816 & n23113;
  assign n23270 = ~n23268 & ~n23269;
  assign n23271 = pi628 & n23270;
  assign n23272 = ~pi1156 & ~n23271;
  assign n23273 = ~n23267 & n23272;
  assign n23274 = ~n17582 & n23240;
  assign n23275 = n17582 & n23113;
  assign n23276 = ~n23274 & ~n23275;
  assign n23277 = pi628 & n23276;
  assign n23278 = ~pi628 & ~n23113;
  assign n23279 = pi1156 & ~n23278;
  assign n23280 = ~n23277 & n23279;
  assign n23281 = ~pi629 & ~n23280;
  assign n23282 = ~n23273 & n23281;
  assign n23283 = pi628 & n23266;
  assign n23284 = ~pi628 & n23270;
  assign n23285 = pi1156 & ~n23284;
  assign n23286 = ~n23283 & n23285;
  assign n23287 = ~pi628 & n23276;
  assign n23288 = pi628 & ~n23113;
  assign n23289 = ~pi1156 & ~n23288;
  assign n23290 = ~n23287 & n23289;
  assign n23291 = pi629 & ~n23290;
  assign n23292 = ~n23286 & n23291;
  assign n23293 = ~n23282 & ~n23292;
  assign n23294 = pi792 & ~n23293;
  assign n23295 = ~pi792 & n23266;
  assign n23296 = ~n23294 & ~n23295;
  assign n23297 = ~pi647 & ~n23296;
  assign n23298 = ~n17610 & ~n23270;
  assign n23299 = n17610 & n23113;
  assign n23300 = ~n23298 & ~n23299;
  assign n23301 = pi647 & n23300;
  assign n23302 = ~pi1157 & ~n23301;
  assign n23303 = ~n23297 & n23302;
  assign n23304 = ~pi792 & ~n23276;
  assign n23305 = ~n23280 & ~n23290;
  assign n23306 = pi792 & ~n23305;
  assign n23307 = ~n23304 & ~n23306;
  assign n23308 = pi647 & n23307;
  assign n23309 = ~pi647 & ~n23113;
  assign n23310 = pi1157 & ~n23309;
  assign n23311 = ~n23308 & n23310;
  assign n23312 = ~pi630 & ~n23311;
  assign n23313 = ~n23303 & n23312;
  assign n23314 = pi647 & ~n23296;
  assign n23315 = ~pi647 & n23300;
  assign n23316 = pi1157 & ~n23315;
  assign n23317 = ~n23314 & n23316;
  assign n23318 = ~pi647 & n23307;
  assign n23319 = pi647 & ~n23113;
  assign n23320 = ~pi1157 & ~n23319;
  assign n23321 = ~n23318 & n23320;
  assign n23322 = pi630 & ~n23321;
  assign n23323 = ~n23317 & n23322;
  assign n23324 = ~n23313 & ~n23323;
  assign n23325 = pi787 & ~n23324;
  assign n23326 = ~pi787 & ~n23296;
  assign n23327 = ~n23325 & ~n23326;
  assign n23328 = ~pi644 & ~n23327;
  assign n23329 = ~pi787 & ~n23307;
  assign n23330 = ~n23311 & ~n23321;
  assign n23331 = pi787 & ~n23330;
  assign n23332 = ~n23329 & ~n23331;
  assign n23333 = pi644 & n23332;
  assign n23334 = ~pi715 & ~n23333;
  assign n23335 = ~n23328 & n23334;
  assign n23336 = n17652 & ~n23113;
  assign n23337 = ~n17652 & n23300;
  assign n23338 = ~n23336 & ~n23337;
  assign n23339 = ~pi644 & ~n23338;
  assign n23340 = pi644 & ~n23113;
  assign n23341 = pi715 & ~n23340;
  assign n23342 = ~n23339 & n23341;
  assign n23343 = ~pi1160 & ~n23342;
  assign n23344 = ~n23335 & n23343;
  assign n23345 = pi644 & ~n23327;
  assign n23346 = ~pi644 & n23332;
  assign n23347 = pi715 & ~n23346;
  assign n23348 = ~n23345 & n23347;
  assign n23349 = pi644 & ~n23338;
  assign n23350 = ~pi644 & ~n23113;
  assign n23351 = ~pi715 & ~n23350;
  assign n23352 = ~n23349 & n23351;
  assign n23353 = pi1160 & ~n23352;
  assign n23354 = ~n23348 & n23353;
  assign n23355 = pi790 & ~n23354;
  assign n23356 = ~n23344 & n23355;
  assign n23357 = ~pi790 & n23327;
  assign n23358 = n6286 & ~n23357;
  assign n23359 = ~n23356 & n23358;
  assign n23360 = ~pi174 & ~n6286;
  assign n23361 = ~pi57 & ~n23360;
  assign n23362 = ~n23359 & n23361;
  assign n23363 = pi57 & pi174;
  assign n23364 = ~pi832 & ~n23363;
  assign n23365 = ~n23362 & n23364;
  assign n23366 = pi174 & ~n2754;
  assign n23367 = pi759 & n16784;
  assign n23368 = ~n23366 & ~n23367;
  assign n23369 = pi696 & n16787;
  assign n23370 = n23368 & ~n23369;
  assign n23371 = pi625 & n23369;
  assign n23372 = ~n23370 & ~n23371;
  assign n23373 = ~pi1153 & ~n23372;
  assign n23374 = pi696 & n16786;
  assign n23375 = pi625 & n23374;
  assign n23376 = pi1153 & ~n23366;
  assign n23377 = ~n23375 & n23376;
  assign n23378 = ~pi608 & ~n23377;
  assign n23379 = ~n23373 & n23378;
  assign n23380 = pi1153 & n23368;
  assign n23381 = ~n23371 & n23380;
  assign n23382 = ~n23366 & ~n23374;
  assign n23383 = ~n23375 & ~n23382;
  assign n23384 = ~pi1153 & ~n23383;
  assign n23385 = pi608 & ~n23384;
  assign n23386 = ~n23381 & n23385;
  assign n23387 = ~n23379 & ~n23386;
  assign n23388 = pi778 & ~n23387;
  assign n23389 = ~pi778 & ~n23370;
  assign n23390 = ~n23388 & ~n23389;
  assign n23391 = ~pi609 & ~n23390;
  assign n23392 = ~pi778 & n23382;
  assign n23393 = ~n23377 & ~n23384;
  assign n23394 = pi778 & ~n23393;
  assign n23395 = ~n23392 & ~n23394;
  assign n23396 = pi609 & n23395;
  assign n23397 = ~pi1155 & ~n23396;
  assign n23398 = ~n23391 & n23397;
  assign n23399 = n17439 & n23367;
  assign n23400 = pi1155 & ~n23366;
  assign n23401 = ~n23399 & n23400;
  assign n23402 = ~pi660 & ~n23401;
  assign n23403 = ~n23398 & n23402;
  assign n23404 = pi609 & ~n23390;
  assign n23405 = ~pi609 & n23395;
  assign n23406 = pi1155 & ~n23405;
  assign n23407 = ~n23404 & n23406;
  assign n23408 = n17451 & n23367;
  assign n23409 = ~pi1155 & ~n23366;
  assign n23410 = ~n23408 & n23409;
  assign n23411 = pi660 & ~n23410;
  assign n23412 = ~n23407 & n23411;
  assign n23413 = ~n23403 & ~n23412;
  assign n23414 = pi785 & ~n23413;
  assign n23415 = ~pi785 & ~n23390;
  assign n23416 = ~n23414 & ~n23415;
  assign n23417 = ~pi618 & ~n23416;
  assign n23418 = ~n17692 & n23395;
  assign n23419 = pi618 & n23418;
  assign n23420 = ~pi1154 & ~n23419;
  assign n23421 = ~n23417 & n23420;
  assign n23422 = ~n20069 & n23367;
  assign n23423 = n20154 & n23422;
  assign n23424 = pi1154 & ~n23366;
  assign n23425 = ~n23423 & n23424;
  assign n23426 = ~pi627 & ~n23425;
  assign n23427 = ~n23421 & n23426;
  assign n23428 = pi618 & ~n23416;
  assign n23429 = ~pi618 & n23418;
  assign n23430 = pi1154 & ~n23429;
  assign n23431 = ~n23428 & n23430;
  assign n23432 = n20164 & n23422;
  assign n23433 = ~pi1154 & ~n23366;
  assign n23434 = ~n23432 & n23433;
  assign n23435 = pi627 & ~n23434;
  assign n23436 = ~n23431 & n23435;
  assign n23437 = ~n23427 & ~n23436;
  assign n23438 = pi781 & ~n23437;
  assign n23439 = ~pi781 & ~n23416;
  assign n23440 = pi648 & n20076;
  assign n23441 = ~pi648 & n20077;
  assign n23442 = ~n23440 & ~n23441;
  assign n23443 = n17538 & n23442;
  assign n23444 = pi789 & ~n23443;
  assign n23445 = ~n23439 & ~n23444;
  assign n23446 = ~n23438 & n23445;
  assign n23447 = n19127 & n23395;
  assign n23448 = ~n23442 & ~n23447;
  assign n23449 = ~n20075 & n23422;
  assign n23450 = n20179 & n23449;
  assign n23451 = n17537 & ~n23450;
  assign n23452 = n20189 & n23449;
  assign n23453 = n17536 & ~n23452;
  assign n23454 = ~n23451 & ~n23453;
  assign n23455 = ~n23448 & n23454;
  assign n23456 = pi789 & ~n23366;
  assign n23457 = ~n23455 & n23456;
  assign n23458 = n17817 & ~n23457;
  assign n23459 = ~n23446 & n23458;
  assign n23460 = ~n17539 & n23447;
  assign n23461 = ~n23366 & ~n23460;
  assign n23462 = n17699 & ~n23461;
  assign n23463 = n20081 & n23422;
  assign n23464 = pi626 & n23463;
  assign n23465 = ~n23366 & ~n23464;
  assign n23466 = pi1158 & ~n23465;
  assign n23467 = ~pi641 & ~n23466;
  assign n23468 = ~n23462 & n23467;
  assign n23469 = n17698 & ~n23461;
  assign n23470 = ~pi626 & n23463;
  assign n23471 = ~n23366 & ~n23470;
  assign n23472 = ~pi1158 & ~n23471;
  assign n23473 = pi641 & ~n23472;
  assign n23474 = ~n23469 & n23473;
  assign n23475 = pi788 & ~n23474;
  assign n23476 = ~n23468 & n23475;
  assign n23477 = ~n20205 & ~n23476;
  assign n23478 = ~n23459 & n23477;
  assign n23479 = ~n17816 & n23463;
  assign n23480 = ~pi629 & n23479;
  assign n23481 = pi628 & ~n23480;
  assign n23482 = n19128 & n23395;
  assign n23483 = pi629 & ~n23482;
  assign n23484 = ~n23481 & ~n23483;
  assign n23485 = ~pi1156 & ~n23484;
  assign n23486 = pi628 & n23482;
  assign n23487 = ~pi628 & ~n23479;
  assign n23488 = pi629 & ~n23487;
  assign n23489 = pi1156 & ~n23488;
  assign n23490 = ~n23486 & n23489;
  assign n23491 = ~n23485 & ~n23490;
  assign n23492 = pi792 & ~n23366;
  assign n23493 = ~n23491 & n23492;
  assign n23494 = ~n23478 & ~n23493;
  assign n23495 = n20207 & ~n23494;
  assign n23496 = ~n17610 & n23479;
  assign n23497 = ~pi630 & n23496;
  assign n23498 = pi647 & ~n23497;
  assign n23499 = ~n19158 & n23482;
  assign n23500 = pi630 & ~n23499;
  assign n23501 = ~n23498 & ~n23500;
  assign n23502 = ~pi1157 & ~n23501;
  assign n23503 = ~pi630 & ~n23499;
  assign n23504 = pi647 & ~n23503;
  assign n23505 = pi630 & n23496;
  assign n23506 = pi1157 & ~n23505;
  assign n23507 = ~n23504 & n23506;
  assign n23508 = ~n23502 & ~n23507;
  assign n23509 = pi787 & ~n23366;
  assign n23510 = ~n23508 & n23509;
  assign n23511 = ~n23495 & ~n23510;
  assign n23512 = pi644 & n23511;
  assign n23513 = ~n19182 & n23499;
  assign n23514 = ~n23366 & ~n23513;
  assign n23515 = ~pi644 & ~n23514;
  assign n23516 = pi715 & ~n23515;
  assign n23517 = ~n23512 & n23516;
  assign n23518 = ~n17610 & ~n17652;
  assign n23519 = n23479 & n23518;
  assign n23520 = pi644 & n23519;
  assign n23521 = ~pi715 & ~n23366;
  assign n23522 = ~n23520 & n23521;
  assign n23523 = pi1160 & ~n23522;
  assign n23524 = ~n23517 & n23523;
  assign n23525 = ~pi644 & n23511;
  assign n23526 = pi644 & ~n23514;
  assign n23527 = ~pi715 & ~n23526;
  assign n23528 = ~n23525 & n23527;
  assign n23529 = ~pi644 & n23519;
  assign n23530 = pi715 & ~n23366;
  assign n23531 = ~n23529 & n23530;
  assign n23532 = ~pi1160 & ~n23531;
  assign n23533 = ~n23528 & n23532;
  assign n23534 = ~n23524 & ~n23533;
  assign n23535 = pi790 & ~n23534;
  assign n23536 = ~pi790 & n23511;
  assign n23537 = pi832 & ~n23536;
  assign n23538 = ~n23535 & n23537;
  assign po331 = ~n23365 & ~n23538;
  assign n23540 = ~pi175 & ~n2754;
  assign n23541 = pi766 & n16784;
  assign n23542 = ~n23540 & ~n23541;
  assign n23543 = ~n17706 & ~n23542;
  assign n23544 = ~pi785 & ~n23543;
  assign n23545 = n17451 & n23541;
  assign n23546 = n23543 & ~n23545;
  assign n23547 = pi1155 & ~n23546;
  assign n23548 = ~pi1155 & ~n23540;
  assign n23549 = ~n23545 & n23548;
  assign n23550 = ~n23547 & ~n23549;
  assign n23551 = pi785 & ~n23550;
  assign n23552 = ~n23544 & ~n23551;
  assign n23553 = ~pi781 & ~n23552;
  assign n23554 = ~n17721 & n23552;
  assign n23555 = pi1154 & ~n23554;
  assign n23556 = ~n17724 & n23552;
  assign n23557 = ~pi1154 & ~n23556;
  assign n23558 = ~n23555 & ~n23557;
  assign n23559 = pi781 & ~n23558;
  assign n23560 = ~n23553 & ~n23559;
  assign n23561 = ~pi789 & ~n23560;
  assign n23562 = ~n22890 & n23560;
  assign n23563 = pi1159 & ~n23562;
  assign n23564 = ~n22893 & n23560;
  assign n23565 = ~pi1159 & ~n23564;
  assign n23566 = ~n23563 & ~n23565;
  assign n23567 = pi789 & ~n23566;
  assign n23568 = ~n23561 & ~n23567;
  assign n23569 = ~n17816 & n23568;
  assign n23570 = n17816 & n23540;
  assign n23571 = ~n23569 & ~n23570;
  assign n23572 = ~n17610 & ~n23571;
  assign n23573 = n17610 & n23540;
  assign n23574 = ~n23572 & ~n23573;
  assign n23575 = ~n20398 & n23574;
  assign n23576 = pi700 & n16786;
  assign n23577 = ~n23540 & ~n23576;
  assign n23578 = ~pi778 & ~n23577;
  assign n23579 = ~pi625 & n23576;
  assign n23580 = ~n23577 & ~n23579;
  assign n23581 = pi1153 & ~n23580;
  assign n23582 = ~pi1153 & ~n23540;
  assign n23583 = ~n23579 & n23582;
  assign n23584 = pi778 & ~n23583;
  assign n23585 = ~n23581 & n23584;
  assign n23586 = ~n23578 & ~n23585;
  assign n23587 = ~n17692 & ~n23586;
  assign n23588 = ~n17694 & n23587;
  assign n23589 = ~n17696 & n23588;
  assign n23590 = ~n17828 & n23589;
  assign n23591 = ~n17859 & n23590;
  assign n23592 = ~pi647 & n23591;
  assign n23593 = pi647 & n23540;
  assign n23594 = ~pi1157 & ~n23593;
  assign n23595 = ~n23592 & n23594;
  assign n23596 = pi647 & ~n23591;
  assign n23597 = ~pi647 & ~n23540;
  assign n23598 = ~n23596 & ~n23597;
  assign n23599 = pi1157 & ~n23598;
  assign n23600 = ~n23595 & ~n23599;
  assign n23601 = ~n17651 & ~n23600;
  assign n23602 = ~n23575 & ~n23601;
  assign n23603 = pi787 & ~n23602;
  assign n23604 = pi626 & ~n23568;
  assign n23605 = ~pi626 & ~n23540;
  assign n23606 = n17579 & ~n23605;
  assign n23607 = ~n23604 & n23606;
  assign n23608 = n17704 & n23589;
  assign n23609 = ~pi626 & ~n23568;
  assign n23610 = pi626 & ~n23540;
  assign n23611 = n17580 & ~n23610;
  assign n23612 = ~n23609 & n23611;
  assign n23613 = ~n23608 & ~n23612;
  assign n23614 = ~n23607 & n23613;
  assign n23615 = pi788 & ~n23614;
  assign n23616 = ~n16521 & ~n23577;
  assign n23617 = pi625 & n23616;
  assign n23618 = n23542 & ~n23616;
  assign n23619 = ~n23617 & ~n23618;
  assign n23620 = n23582 & ~n23619;
  assign n23621 = ~pi608 & ~n23581;
  assign n23622 = ~n23620 & n23621;
  assign n23623 = pi1153 & n23542;
  assign n23624 = ~n23617 & n23623;
  assign n23625 = pi608 & ~n23583;
  assign n23626 = ~n23624 & n23625;
  assign n23627 = ~n23622 & ~n23626;
  assign n23628 = pi778 & ~n23627;
  assign n23629 = ~pi778 & ~n23618;
  assign n23630 = ~n23628 & ~n23629;
  assign n23631 = ~pi609 & ~n23630;
  assign n23632 = pi609 & ~n23586;
  assign n23633 = ~pi1155 & ~n23632;
  assign n23634 = ~n23631 & n23633;
  assign n23635 = ~pi660 & ~n23547;
  assign n23636 = ~n23634 & n23635;
  assign n23637 = pi609 & ~n23630;
  assign n23638 = ~pi609 & ~n23586;
  assign n23639 = pi1155 & ~n23638;
  assign n23640 = ~n23637 & n23639;
  assign n23641 = pi660 & ~n23549;
  assign n23642 = ~n23640 & n23641;
  assign n23643 = ~n23636 & ~n23642;
  assign n23644 = pi785 & ~n23643;
  assign n23645 = ~pi785 & ~n23630;
  assign n23646 = ~n23644 & ~n23645;
  assign n23647 = ~pi618 & ~n23646;
  assign n23648 = pi618 & n23587;
  assign n23649 = ~pi1154 & ~n23648;
  assign n23650 = ~n23647 & n23649;
  assign n23651 = ~pi627 & ~n23555;
  assign n23652 = ~n23650 & n23651;
  assign n23653 = pi618 & ~n23646;
  assign n23654 = ~pi618 & n23587;
  assign n23655 = pi1154 & ~n23654;
  assign n23656 = ~n23653 & n23655;
  assign n23657 = pi627 & ~n23557;
  assign n23658 = ~n23656 & n23657;
  assign n23659 = ~n23652 & ~n23658;
  assign n23660 = pi781 & ~n23659;
  assign n23661 = ~pi781 & ~n23646;
  assign n23662 = ~n23660 & ~n23661;
  assign n23663 = pi619 & ~n23662;
  assign n23664 = ~pi619 & n23588;
  assign n23665 = pi1159 & ~n23664;
  assign n23666 = ~n23663 & n23665;
  assign n23667 = pi648 & ~n23565;
  assign n23668 = ~n23666 & n23667;
  assign n23669 = ~pi619 & ~n23662;
  assign n23670 = pi619 & n23588;
  assign n23671 = ~pi1159 & ~n23670;
  assign n23672 = ~n23669 & n23671;
  assign n23673 = ~pi648 & ~n23563;
  assign n23674 = ~n23672 & n23673;
  assign n23675 = pi789 & ~n23674;
  assign n23676 = ~n23668 & n23675;
  assign n23677 = ~pi789 & n23662;
  assign n23678 = n17817 & ~n23677;
  assign n23679 = ~n23676 & n23678;
  assign n23680 = ~n23615 & ~n23679;
  assign n23681 = ~n20205 & ~n23680;
  assign n23682 = n17856 & ~n23571;
  assign n23683 = n20693 & n23590;
  assign n23684 = ~n23682 & ~n23683;
  assign n23685 = ~pi629 & ~n23684;
  assign n23686 = n20697 & n23590;
  assign n23687 = n17855 & ~n23571;
  assign n23688 = ~n23686 & ~n23687;
  assign n23689 = pi629 & ~n23688;
  assign n23690 = ~n23685 & ~n23689;
  assign n23691 = pi792 & ~n23690;
  assign n23692 = n20207 & ~n23691;
  assign n23693 = ~n23681 & n23692;
  assign n23694 = ~n23603 & ~n23693;
  assign n23695 = pi644 & n23694;
  assign n23696 = ~pi787 & ~n23591;
  assign n23697 = pi787 & ~n23600;
  assign n23698 = ~n23696 & ~n23697;
  assign n23699 = ~pi644 & n23698;
  assign n23700 = pi715 & ~n23699;
  assign n23701 = ~n23695 & n23700;
  assign n23702 = ~n17652 & ~n23574;
  assign n23703 = n17652 & n23540;
  assign n23704 = ~n23702 & ~n23703;
  assign n23705 = pi644 & ~n23704;
  assign n23706 = ~pi644 & n23540;
  assign n23707 = ~pi715 & ~n23706;
  assign n23708 = ~n23705 & n23707;
  assign n23709 = pi1160 & ~n23708;
  assign n23710 = ~n23701 & n23709;
  assign n23711 = ~pi644 & n23694;
  assign n23712 = pi644 & n23698;
  assign n23713 = ~pi715 & ~n23712;
  assign n23714 = ~n23711 & n23713;
  assign n23715 = ~pi644 & ~n23704;
  assign n23716 = pi644 & n23540;
  assign n23717 = pi715 & ~n23716;
  assign n23718 = ~n23715 & n23717;
  assign n23719 = ~pi1160 & ~n23718;
  assign n23720 = ~n23714 & n23719;
  assign n23721 = ~n23710 & ~n23720;
  assign n23722 = pi790 & ~n23721;
  assign n23723 = ~pi790 & n23694;
  assign n23724 = pi832 & ~n23723;
  assign n23725 = ~n23722 & n23724;
  assign n23726 = ~pi175 & ~n17406;
  assign n23727 = n17539 & ~n23726;
  assign n23728 = pi175 & ~n3267;
  assign n23729 = ~pi175 & n17972;
  assign n23730 = pi175 & ~n17976;
  assign n23731 = ~pi38 & ~n23730;
  assign n23732 = ~n23729 & n23731;
  assign n23733 = ~pi175 & ~n17280;
  assign n23734 = n17392 & ~n23733;
  assign n23735 = pi700 & ~n23734;
  assign n23736 = ~n23732 & n23735;
  assign n23737 = ~pi175 & ~pi700;
  assign n23738 = ~n17399 & n23737;
  assign n23739 = n3267 & ~n23738;
  assign n23740 = ~n23736 & n23739;
  assign n23741 = ~n23728 & ~n23740;
  assign n23742 = ~pi778 & ~n23741;
  assign n23743 = pi625 & n23741;
  assign n23744 = ~pi625 & n23726;
  assign n23745 = pi1153 & ~n23744;
  assign n23746 = ~n23743 & n23745;
  assign n23747 = ~pi625 & n23741;
  assign n23748 = pi625 & n23726;
  assign n23749 = ~pi1153 & ~n23748;
  assign n23750 = ~n23747 & n23749;
  assign n23751 = ~n23746 & ~n23750;
  assign n23752 = pi778 & ~n23751;
  assign n23753 = ~n23742 & ~n23752;
  assign n23754 = ~n17466 & ~n23753;
  assign n23755 = n17466 & ~n23726;
  assign n23756 = ~n23754 & ~n23755;
  assign n23757 = ~n17503 & n23756;
  assign n23758 = n17503 & n23726;
  assign n23759 = ~n23757 & ~n23758;
  assign n23760 = ~n17539 & n23759;
  assign n23761 = ~n23727 & ~n23760;
  assign n23762 = ~n17582 & n23761;
  assign n23763 = n17582 & n23726;
  assign n23764 = ~n23762 & ~n23763;
  assign n23765 = ~pi628 & ~n23764;
  assign n23766 = pi628 & n23726;
  assign n23767 = ~n23765 & ~n23766;
  assign n23768 = ~pi1156 & ~n23767;
  assign n23769 = pi628 & ~n23764;
  assign n23770 = ~pi628 & n23726;
  assign n23771 = ~n23769 & ~n23770;
  assign n23772 = pi1156 & ~n23771;
  assign n23773 = ~n23768 & ~n23772;
  assign n23774 = pi792 & ~n23773;
  assign n23775 = ~pi792 & ~n23764;
  assign n23776 = ~n23774 & ~n23775;
  assign n23777 = ~pi647 & ~n23776;
  assign n23778 = pi647 & n23726;
  assign n23779 = ~n23777 & ~n23778;
  assign n23780 = ~pi1157 & ~n23779;
  assign n23781 = pi647 & ~n23776;
  assign n23782 = ~pi647 & n23726;
  assign n23783 = ~n23781 & ~n23782;
  assign n23784 = pi1157 & ~n23783;
  assign n23785 = ~n23780 & ~n23784;
  assign n23786 = pi787 & ~n23785;
  assign n23787 = ~pi787 & ~n23776;
  assign n23788 = ~n23786 & ~n23787;
  assign n23789 = ~pi644 & ~n23788;
  assign n23790 = pi715 & ~n23789;
  assign n23791 = ~pi766 & n17199;
  assign n23792 = pi175 & n17273;
  assign n23793 = ~n23791 & ~n23792;
  assign n23794 = pi39 & ~n23793;
  assign n23795 = ~pi175 & pi766;
  assign n23796 = n17242 & n23795;
  assign n23797 = pi766 & ~n17246;
  assign n23798 = pi175 & ~n23797;
  assign n23799 = ~n21331 & ~n23798;
  assign n23800 = ~n23796 & n23799;
  assign n23801 = ~n23794 & n23800;
  assign n23802 = ~pi38 & ~n23801;
  assign n23803 = pi766 & n17282;
  assign n23804 = pi38 & ~n23733;
  assign n23805 = ~n23803 & n23804;
  assign n23806 = ~n23802 & ~n23805;
  assign n23807 = n3267 & ~n23806;
  assign n23808 = ~n23728 & ~n23807;
  assign n23809 = ~n17438 & ~n23808;
  assign n23810 = n17438 & ~n23726;
  assign n23811 = ~n23809 & ~n23810;
  assign n23812 = ~pi785 & ~n23811;
  assign n23813 = ~n17439 & ~n23726;
  assign n23814 = pi609 & n23809;
  assign n23815 = ~n23813 & ~n23814;
  assign n23816 = pi1155 & ~n23815;
  assign n23817 = ~n17451 & ~n23726;
  assign n23818 = ~pi609 & n23809;
  assign n23819 = ~n23817 & ~n23818;
  assign n23820 = ~pi1155 & ~n23819;
  assign n23821 = ~n23816 & ~n23820;
  assign n23822 = pi785 & ~n23821;
  assign n23823 = ~n23812 & ~n23822;
  assign n23824 = ~pi781 & ~n23823;
  assign n23825 = pi618 & n23823;
  assign n23826 = ~pi618 & n23726;
  assign n23827 = pi1154 & ~n23826;
  assign n23828 = ~n23825 & n23827;
  assign n23829 = ~pi618 & n23823;
  assign n23830 = pi618 & n23726;
  assign n23831 = ~pi1154 & ~n23830;
  assign n23832 = ~n23829 & n23831;
  assign n23833 = ~n23828 & ~n23832;
  assign n23834 = pi781 & ~n23833;
  assign n23835 = ~n23824 & ~n23834;
  assign n23836 = ~pi789 & ~n23835;
  assign n23837 = pi619 & n23835;
  assign n23838 = ~pi619 & n23726;
  assign n23839 = pi1159 & ~n23838;
  assign n23840 = ~n23837 & n23839;
  assign n23841 = ~pi619 & n23835;
  assign n23842 = pi619 & n23726;
  assign n23843 = ~pi1159 & ~n23842;
  assign n23844 = ~n23841 & n23843;
  assign n23845 = ~n23840 & ~n23844;
  assign n23846 = pi789 & ~n23845;
  assign n23847 = ~n23836 & ~n23846;
  assign n23848 = ~n17816 & n23847;
  assign n23849 = n17816 & n23726;
  assign n23850 = ~n23848 & ~n23849;
  assign n23851 = ~n17610 & ~n23850;
  assign n23852 = n17610 & n23726;
  assign n23853 = ~n23851 & ~n23852;
  assign n23854 = ~n17652 & ~n23853;
  assign n23855 = n17652 & n23726;
  assign n23856 = ~n23854 & ~n23855;
  assign n23857 = pi644 & ~n23856;
  assign n23858 = ~pi644 & n23726;
  assign n23859 = ~pi715 & ~n23858;
  assign n23860 = ~n23857 & n23859;
  assign n23861 = pi1160 & ~n23860;
  assign n23862 = ~n23790 & n23861;
  assign n23863 = pi644 & ~n23788;
  assign n23864 = ~pi715 & ~n23863;
  assign n23865 = ~pi644 & ~n23856;
  assign n23866 = pi644 & n23726;
  assign n23867 = pi715 & ~n23866;
  assign n23868 = ~n23865 & n23867;
  assign n23869 = ~pi1160 & ~n23868;
  assign n23870 = ~n23864 & n23869;
  assign n23871 = ~n23862 & ~n23870;
  assign n23872 = pi790 & ~n23871;
  assign n23873 = pi644 & n23861;
  assign n23874 = ~pi644 & n23869;
  assign n23875 = pi790 & ~n23874;
  assign n23876 = ~n23873 & n23875;
  assign n23877 = ~n20409 & n23850;
  assign n23878 = n17608 & n23767;
  assign n23879 = n17607 & n23771;
  assign n23880 = ~n23878 & ~n23879;
  assign n23881 = ~n23877 & n23880;
  assign n23882 = pi792 & ~n23881;
  assign n23883 = ~pi700 & n23806;
  assign n23884 = ~pi175 & n16687;
  assign n23885 = pi175 & n16799;
  assign n23886 = ~pi766 & ~n23885;
  assign n23887 = ~n23884 & n23886;
  assign n23888 = pi175 & n16879;
  assign n23889 = ~pi175 & ~n16944;
  assign n23890 = pi766 & ~n23889;
  assign n23891 = ~n23888 & n23890;
  assign n23892 = pi39 & ~n23891;
  assign n23893 = ~n23887 & n23892;
  assign n23894 = pi175 & n17059;
  assign n23895 = ~pi175 & n17088;
  assign n23896 = ~pi766 & ~n23895;
  assign n23897 = ~n23894 & n23896;
  assign n23898 = ~pi175 & ~n17092;
  assign n23899 = pi175 & ~n17094;
  assign n23900 = pi766 & ~n23899;
  assign n23901 = ~n23898 & n23900;
  assign n23902 = ~pi39 & ~n23901;
  assign n23903 = ~n23897 & n23902;
  assign n23904 = ~pi38 & ~n23903;
  assign n23905 = ~n23893 & n23904;
  assign n23906 = ~n16522 & n16529;
  assign n23907 = ~pi766 & n23906;
  assign n23908 = ~n16905 & ~n23907;
  assign n23909 = ~pi39 & ~n23908;
  assign n23910 = ~pi175 & ~n23909;
  assign n23911 = ~n16787 & ~n23541;
  assign n23912 = pi175 & ~n23911;
  assign n23913 = n6234 & n23912;
  assign n23914 = pi38 & ~n23913;
  assign n23915 = ~n23910 & n23914;
  assign n23916 = pi700 & ~n23915;
  assign n23917 = ~n23905 & n23916;
  assign n23918 = n3267 & ~n23917;
  assign n23919 = ~n23883 & n23918;
  assign n23920 = ~n23728 & ~n23919;
  assign n23921 = ~pi625 & n23920;
  assign n23922 = pi625 & n23808;
  assign n23923 = ~pi1153 & ~n23922;
  assign n23924 = ~n23921 & n23923;
  assign n23925 = ~pi608 & ~n23746;
  assign n23926 = ~n23924 & n23925;
  assign n23927 = pi625 & n23920;
  assign n23928 = ~pi625 & n23808;
  assign n23929 = pi1153 & ~n23928;
  assign n23930 = ~n23927 & n23929;
  assign n23931 = pi608 & ~n23750;
  assign n23932 = ~n23930 & n23931;
  assign n23933 = ~n23926 & ~n23932;
  assign n23934 = pi778 & ~n23933;
  assign n23935 = ~pi778 & n23920;
  assign n23936 = ~n23934 & ~n23935;
  assign n23937 = ~pi609 & ~n23936;
  assign n23938 = pi609 & n23753;
  assign n23939 = ~pi1155 & ~n23938;
  assign n23940 = ~n23937 & n23939;
  assign n23941 = ~pi660 & ~n23816;
  assign n23942 = ~n23940 & n23941;
  assign n23943 = pi609 & ~n23936;
  assign n23944 = ~pi609 & n23753;
  assign n23945 = pi1155 & ~n23944;
  assign n23946 = ~n23943 & n23945;
  assign n23947 = pi660 & ~n23820;
  assign n23948 = ~n23946 & n23947;
  assign n23949 = ~n23942 & ~n23948;
  assign n23950 = pi785 & ~n23949;
  assign n23951 = ~pi785 & ~n23936;
  assign n23952 = ~n23950 & ~n23951;
  assign n23953 = ~pi618 & ~n23952;
  assign n23954 = pi618 & n23756;
  assign n23955 = ~pi1154 & ~n23954;
  assign n23956 = ~n23953 & n23955;
  assign n23957 = ~pi627 & ~n23828;
  assign n23958 = ~n23956 & n23957;
  assign n23959 = pi618 & ~n23952;
  assign n23960 = ~pi618 & n23756;
  assign n23961 = pi1154 & ~n23960;
  assign n23962 = ~n23959 & n23961;
  assign n23963 = pi627 & ~n23832;
  assign n23964 = ~n23962 & n23963;
  assign n23965 = ~n23958 & ~n23964;
  assign n23966 = pi781 & ~n23965;
  assign n23967 = ~pi781 & ~n23952;
  assign n23968 = ~n23966 & ~n23967;
  assign n23969 = pi619 & ~n23968;
  assign n23970 = ~pi619 & ~n23759;
  assign n23971 = pi1159 & ~n23970;
  assign n23972 = ~n23969 & n23971;
  assign n23973 = pi648 & ~n23844;
  assign n23974 = ~n23972 & n23973;
  assign n23975 = ~pi619 & ~n23968;
  assign n23976 = pi619 & ~n23759;
  assign n23977 = ~pi1159 & ~n23976;
  assign n23978 = ~n23975 & n23977;
  assign n23979 = ~pi648 & ~n23840;
  assign n23980 = ~n23978 & n23979;
  assign n23981 = pi789 & ~n23980;
  assign n23982 = ~n23974 & n23981;
  assign n23983 = ~pi789 & n23968;
  assign n23984 = n17817 & ~n23983;
  assign n23985 = ~n23982 & n23984;
  assign n23986 = pi626 & ~n23847;
  assign n23987 = ~pi626 & ~n23726;
  assign n23988 = n17579 & ~n23987;
  assign n23989 = ~n23986 & n23988;
  assign n23990 = n17704 & n23761;
  assign n23991 = ~pi626 & ~n23847;
  assign n23992 = pi626 & ~n23726;
  assign n23993 = n17580 & ~n23992;
  assign n23994 = ~n23991 & n23993;
  assign n23995 = ~n23990 & ~n23994;
  assign n23996 = ~n23989 & n23995;
  assign n23997 = pi788 & ~n23996;
  assign n23998 = ~n20205 & ~n23997;
  assign n23999 = ~n23985 & n23998;
  assign n24000 = ~n23882 & ~n23999;
  assign n24001 = n20207 & ~n24000;
  assign n24002 = n17649 & n23783;
  assign n24003 = n17650 & n23779;
  assign n24004 = ~n20398 & n23853;
  assign n24005 = ~n24003 & ~n24004;
  assign n24006 = ~n24002 & n24005;
  assign n24007 = pi787 & ~n24006;
  assign n24008 = ~n24001 & ~n24007;
  assign n24009 = ~n23876 & n24008;
  assign n24010 = ~n23872 & ~n24009;
  assign n24011 = ~po1038 & ~n24010;
  assign n24012 = ~pi175 & po1038;
  assign n24013 = ~pi832 & ~n24012;
  assign n24014 = ~n24011 & n24013;
  assign po332 = ~n23725 & ~n24014;
  assign n24016 = ~pi176 & ~n2754;
  assign n24017 = ~pi742 & n16784;
  assign n24018 = ~n24016 & ~n24017;
  assign n24019 = ~n17706 & ~n24018;
  assign n24020 = ~pi785 & ~n24019;
  assign n24021 = ~n17711 & ~n24018;
  assign n24022 = pi1155 & ~n24021;
  assign n24023 = ~n17714 & n24019;
  assign n24024 = ~pi1155 & ~n24023;
  assign n24025 = ~n24022 & ~n24024;
  assign n24026 = pi785 & ~n24025;
  assign n24027 = ~n24020 & ~n24026;
  assign n24028 = ~pi781 & ~n24027;
  assign n24029 = ~n17721 & n24027;
  assign n24030 = pi1154 & ~n24029;
  assign n24031 = ~n17724 & n24027;
  assign n24032 = ~pi1154 & ~n24031;
  assign n24033 = ~n24030 & ~n24032;
  assign n24034 = pi781 & ~n24033;
  assign n24035 = ~n24028 & ~n24034;
  assign n24036 = ~pi789 & ~n24035;
  assign n24037 = pi619 & n24035;
  assign n24038 = ~pi619 & n24016;
  assign n24039 = pi1159 & ~n24038;
  assign n24040 = ~n24037 & n24039;
  assign n24041 = ~pi619 & n24035;
  assign n24042 = pi619 & n24016;
  assign n24043 = ~pi1159 & ~n24042;
  assign n24044 = ~n24041 & n24043;
  assign n24045 = ~n24040 & ~n24044;
  assign n24046 = pi789 & ~n24045;
  assign n24047 = ~n24036 & ~n24046;
  assign n24048 = ~n17816 & n24047;
  assign n24049 = n17816 & n24016;
  assign n24050 = ~n24048 & ~n24049;
  assign n24051 = ~n17610 & ~n24050;
  assign n24052 = n17610 & n24016;
  assign n24053 = ~n24051 & ~n24052;
  assign n24054 = ~n20398 & n24053;
  assign n24055 = ~pi704 & n16786;
  assign n24056 = ~n24016 & ~n24055;
  assign n24057 = ~pi778 & n24056;
  assign n24058 = ~pi625 & n24055;
  assign n24059 = ~n24056 & ~n24058;
  assign n24060 = pi1153 & ~n24059;
  assign n24061 = ~pi1153 & ~n24016;
  assign n24062 = ~n24058 & n24061;
  assign n24063 = ~n24060 & ~n24062;
  assign n24064 = pi778 & ~n24063;
  assign n24065 = ~n24057 & ~n24064;
  assign n24066 = ~n17692 & n24065;
  assign n24067 = ~n17694 & n24066;
  assign n24068 = ~n17696 & n24067;
  assign n24069 = ~n17828 & n24068;
  assign n24070 = ~n17859 & n24069;
  assign n24071 = ~pi647 & n24070;
  assign n24072 = pi647 & n24016;
  assign n24073 = ~pi1157 & ~n24072;
  assign n24074 = ~n24071 & n24073;
  assign n24075 = pi647 & ~n24070;
  assign n24076 = ~pi647 & ~n24016;
  assign n24077 = ~n24075 & ~n24076;
  assign n24078 = pi1157 & ~n24077;
  assign n24079 = ~n24074 & ~n24078;
  assign n24080 = ~n17651 & ~n24079;
  assign n24081 = ~n24054 & ~n24080;
  assign n24082 = pi787 & ~n24081;
  assign n24083 = pi626 & ~n24047;
  assign n24084 = ~pi626 & ~n24016;
  assign n24085 = n17579 & ~n24084;
  assign n24086 = ~n24083 & n24085;
  assign n24087 = n17704 & n24068;
  assign n24088 = ~pi626 & ~n24047;
  assign n24089 = pi626 & ~n24016;
  assign n24090 = n17580 & ~n24089;
  assign n24091 = ~n24088 & n24090;
  assign n24092 = ~n24087 & ~n24091;
  assign n24093 = ~n24086 & n24092;
  assign n24094 = pi788 & ~n24093;
  assign n24095 = ~n16521 & ~n24056;
  assign n24096 = pi625 & n24095;
  assign n24097 = n24018 & ~n24095;
  assign n24098 = ~n24096 & ~n24097;
  assign n24099 = n24061 & ~n24098;
  assign n24100 = ~pi608 & ~n24060;
  assign n24101 = ~n24099 & n24100;
  assign n24102 = pi1153 & n24018;
  assign n24103 = ~n24096 & n24102;
  assign n24104 = pi608 & ~n24062;
  assign n24105 = ~n24103 & n24104;
  assign n24106 = ~n24101 & ~n24105;
  assign n24107 = pi778 & ~n24106;
  assign n24108 = ~pi778 & ~n24097;
  assign n24109 = ~n24107 & ~n24108;
  assign n24110 = ~pi609 & ~n24109;
  assign n24111 = pi609 & n24065;
  assign n24112 = ~pi1155 & ~n24111;
  assign n24113 = ~n24110 & n24112;
  assign n24114 = ~pi660 & ~n24022;
  assign n24115 = ~n24113 & n24114;
  assign n24116 = pi609 & ~n24109;
  assign n24117 = ~pi609 & n24065;
  assign n24118 = pi1155 & ~n24117;
  assign n24119 = ~n24116 & n24118;
  assign n24120 = pi660 & ~n24024;
  assign n24121 = ~n24119 & n24120;
  assign n24122 = ~n24115 & ~n24121;
  assign n24123 = pi785 & ~n24122;
  assign n24124 = ~pi785 & ~n24109;
  assign n24125 = ~n24123 & ~n24124;
  assign n24126 = ~pi618 & ~n24125;
  assign n24127 = pi618 & n24066;
  assign n24128 = ~pi1154 & ~n24127;
  assign n24129 = ~n24126 & n24128;
  assign n24130 = ~pi627 & ~n24030;
  assign n24131 = ~n24129 & n24130;
  assign n24132 = pi618 & ~n24125;
  assign n24133 = ~pi618 & n24066;
  assign n24134 = pi1154 & ~n24133;
  assign n24135 = ~n24132 & n24134;
  assign n24136 = pi627 & ~n24032;
  assign n24137 = ~n24135 & n24136;
  assign n24138 = ~n24131 & ~n24137;
  assign n24139 = pi781 & ~n24138;
  assign n24140 = ~pi781 & ~n24125;
  assign n24141 = ~n24139 & ~n24140;
  assign n24142 = pi619 & ~n24141;
  assign n24143 = ~pi619 & n24067;
  assign n24144 = pi1159 & ~n24143;
  assign n24145 = ~n24142 & n24144;
  assign n24146 = pi648 & ~n24044;
  assign n24147 = ~n24145 & n24146;
  assign n24148 = ~pi619 & ~n24141;
  assign n24149 = pi619 & n24067;
  assign n24150 = ~pi1159 & ~n24149;
  assign n24151 = ~n24148 & n24150;
  assign n24152 = ~pi648 & ~n24040;
  assign n24153 = ~n24151 & n24152;
  assign n24154 = pi789 & ~n24153;
  assign n24155 = ~n24147 & n24154;
  assign n24156 = ~pi789 & n24141;
  assign n24157 = n17817 & ~n24156;
  assign n24158 = ~n24155 & n24157;
  assign n24159 = ~n24094 & ~n24158;
  assign n24160 = ~n20205 & ~n24159;
  assign n24161 = n17856 & ~n24050;
  assign n24162 = n20693 & n24069;
  assign n24163 = ~n24161 & ~n24162;
  assign n24164 = ~pi629 & ~n24163;
  assign n24165 = n20697 & n24069;
  assign n24166 = n17855 & ~n24050;
  assign n24167 = ~n24165 & ~n24166;
  assign n24168 = pi629 & ~n24167;
  assign n24169 = ~n24164 & ~n24168;
  assign n24170 = pi792 & ~n24169;
  assign n24171 = n20207 & ~n24170;
  assign n24172 = ~n24160 & n24171;
  assign n24173 = ~n24082 & ~n24172;
  assign n24174 = pi644 & n24173;
  assign n24175 = ~pi787 & ~n24070;
  assign n24176 = pi787 & ~n24079;
  assign n24177 = ~n24175 & ~n24176;
  assign n24178 = ~pi644 & n24177;
  assign n24179 = pi715 & ~n24178;
  assign n24180 = ~n24174 & n24179;
  assign n24181 = ~n17652 & ~n24053;
  assign n24182 = n17652 & n24016;
  assign n24183 = ~n24181 & ~n24182;
  assign n24184 = pi644 & ~n24183;
  assign n24185 = ~pi644 & n24016;
  assign n24186 = ~pi715 & ~n24185;
  assign n24187 = ~n24184 & n24186;
  assign n24188 = pi1160 & ~n24187;
  assign n24189 = ~n24180 & n24188;
  assign n24190 = ~pi644 & n24173;
  assign n24191 = pi644 & n24177;
  assign n24192 = ~pi715 & ~n24191;
  assign n24193 = ~n24190 & n24192;
  assign n24194 = ~pi644 & ~n24183;
  assign n24195 = pi644 & n24016;
  assign n24196 = pi715 & ~n24195;
  assign n24197 = ~n24194 & n24196;
  assign n24198 = ~pi1160 & ~n24197;
  assign n24199 = ~n24193 & n24198;
  assign n24200 = ~n24189 & ~n24199;
  assign n24201 = pi790 & ~n24200;
  assign n24202 = ~pi790 & n24173;
  assign n24203 = pi832 & ~n24202;
  assign n24204 = ~n24201 & n24203;
  assign n24205 = ~pi176 & ~n17406;
  assign n24206 = n17539 & ~n24205;
  assign n24207 = ~pi38 & n17976;
  assign n24208 = n3267 & ~n17392;
  assign n24209 = ~n24207 & n24208;
  assign n24210 = pi176 & ~n24209;
  assign n24211 = ~pi38 & n17972;
  assign n24212 = ~n19802 & ~n24211;
  assign n24213 = ~pi176 & n24212;
  assign n24214 = ~pi704 & ~n24213;
  assign n24215 = ~pi176 & ~n17399;
  assign n24216 = pi704 & n24215;
  assign n24217 = n3267 & ~n24216;
  assign n24218 = ~n24214 & n24217;
  assign n24219 = ~n24210 & ~n24218;
  assign n24220 = ~pi778 & ~n24219;
  assign n24221 = pi625 & n24219;
  assign n24222 = ~pi625 & n24205;
  assign n24223 = pi1153 & ~n24222;
  assign n24224 = ~n24221 & n24223;
  assign n24225 = ~pi625 & n24219;
  assign n24226 = pi625 & n24205;
  assign n24227 = ~pi1153 & ~n24226;
  assign n24228 = ~n24225 & n24227;
  assign n24229 = ~n24224 & ~n24228;
  assign n24230 = pi778 & ~n24229;
  assign n24231 = ~n24220 & ~n24230;
  assign n24232 = ~n17466 & ~n24231;
  assign n24233 = n17466 & ~n24205;
  assign n24234 = ~n24232 & ~n24233;
  assign n24235 = ~n17503 & n24234;
  assign n24236 = n17503 & n24205;
  assign n24237 = ~n24235 & ~n24236;
  assign n24238 = ~n17539 & n24237;
  assign n24239 = ~n24206 & ~n24238;
  assign n24240 = ~n17582 & n24239;
  assign n24241 = n17582 & n24205;
  assign n24242 = ~n24240 & ~n24241;
  assign n24243 = ~pi628 & ~n24242;
  assign n24244 = pi628 & n24205;
  assign n24245 = ~n24243 & ~n24244;
  assign n24246 = ~pi1156 & ~n24245;
  assign n24247 = pi628 & ~n24242;
  assign n24248 = ~pi628 & n24205;
  assign n24249 = ~n24247 & ~n24248;
  assign n24250 = pi1156 & ~n24249;
  assign n24251 = ~n24246 & ~n24250;
  assign n24252 = pi792 & ~n24251;
  assign n24253 = ~pi792 & ~n24242;
  assign n24254 = ~n24252 & ~n24253;
  assign n24255 = ~pi647 & ~n24254;
  assign n24256 = pi647 & n24205;
  assign n24257 = ~n24255 & ~n24256;
  assign n24258 = ~pi1157 & ~n24257;
  assign n24259 = pi647 & ~n24254;
  assign n24260 = ~pi647 & n24205;
  assign n24261 = ~n24259 & ~n24260;
  assign n24262 = pi1157 & ~n24261;
  assign n24263 = ~n24258 & ~n24262;
  assign n24264 = pi787 & ~n24263;
  assign n24265 = ~pi787 & ~n24254;
  assign n24266 = ~n24264 & ~n24265;
  assign n24267 = ~pi644 & ~n24266;
  assign n24268 = pi715 & ~n24267;
  assign n24269 = pi176 & ~n3267;
  assign n24270 = ~pi176 & n19223;
  assign n24271 = ~n19217 & ~n19218;
  assign n24272 = pi176 & n24271;
  assign n24273 = ~n24270 & ~n24272;
  assign n24274 = ~pi742 & ~n24273;
  assign n24275 = pi742 & ~n24215;
  assign n24276 = ~n24274 & ~n24275;
  assign n24277 = n3267 & ~n24276;
  assign n24278 = ~n24269 & ~n24277;
  assign n24279 = ~n17438 & ~n24278;
  assign n24280 = n17438 & ~n24205;
  assign n24281 = ~n24279 & ~n24280;
  assign n24282 = ~pi785 & ~n24281;
  assign n24283 = ~n17439 & ~n24205;
  assign n24284 = pi609 & n24279;
  assign n24285 = ~n24283 & ~n24284;
  assign n24286 = pi1155 & ~n24285;
  assign n24287 = ~n17451 & ~n24205;
  assign n24288 = ~pi609 & n24279;
  assign n24289 = ~n24287 & ~n24288;
  assign n24290 = ~pi1155 & ~n24289;
  assign n24291 = ~n24286 & ~n24290;
  assign n24292 = pi785 & ~n24291;
  assign n24293 = ~n24282 & ~n24292;
  assign n24294 = ~pi781 & ~n24293;
  assign n24295 = pi618 & n24293;
  assign n24296 = ~pi618 & n24205;
  assign n24297 = pi1154 & ~n24296;
  assign n24298 = ~n24295 & n24297;
  assign n24299 = ~pi618 & n24293;
  assign n24300 = pi618 & n24205;
  assign n24301 = ~pi1154 & ~n24300;
  assign n24302 = ~n24299 & n24301;
  assign n24303 = ~n24298 & ~n24302;
  assign n24304 = pi781 & ~n24303;
  assign n24305 = ~n24294 & ~n24304;
  assign n24306 = ~pi789 & ~n24305;
  assign n24307 = pi619 & n24305;
  assign n24308 = ~pi619 & n24205;
  assign n24309 = pi1159 & ~n24308;
  assign n24310 = ~n24307 & n24309;
  assign n24311 = ~pi619 & n24305;
  assign n24312 = pi619 & n24205;
  assign n24313 = ~pi1159 & ~n24312;
  assign n24314 = ~n24311 & n24313;
  assign n24315 = ~n24310 & ~n24314;
  assign n24316 = pi789 & ~n24315;
  assign n24317 = ~n24306 & ~n24316;
  assign n24318 = ~n17816 & n24317;
  assign n24319 = n17816 & n24205;
  assign n24320 = ~n24318 & ~n24319;
  assign n24321 = ~n17610 & ~n24320;
  assign n24322 = n17610 & n24205;
  assign n24323 = ~n24321 & ~n24322;
  assign n24324 = ~n17652 & ~n24323;
  assign n24325 = n17652 & n24205;
  assign n24326 = ~n24324 & ~n24325;
  assign n24327 = pi644 & ~n24326;
  assign n24328 = ~pi644 & n24205;
  assign n24329 = ~pi715 & ~n24328;
  assign n24330 = ~n24327 & n24329;
  assign n24331 = pi1160 & ~n24330;
  assign n24332 = ~n24268 & n24331;
  assign n24333 = pi644 & ~n24266;
  assign n24334 = ~pi715 & ~n24333;
  assign n24335 = ~pi644 & ~n24326;
  assign n24336 = pi644 & n24205;
  assign n24337 = pi715 & ~n24336;
  assign n24338 = ~n24335 & n24337;
  assign n24339 = ~pi1160 & ~n24338;
  assign n24340 = ~n24334 & n24339;
  assign n24341 = ~n24332 & ~n24340;
  assign n24342 = pi790 & ~n24341;
  assign n24343 = pi644 & n24331;
  assign n24344 = ~pi644 & n24339;
  assign n24345 = pi790 & ~n24344;
  assign n24346 = ~n24343 & n24345;
  assign n24347 = n17649 & n24261;
  assign n24348 = n17650 & n24257;
  assign n24349 = ~n20398 & n24323;
  assign n24350 = ~n24348 & ~n24349;
  assign n24351 = ~n24347 & n24350;
  assign n24352 = pi787 & ~n24351;
  assign n24353 = ~n20409 & n24320;
  assign n24354 = n17608 & n24245;
  assign n24355 = n17607 & n24249;
  assign n24356 = ~n24354 & ~n24355;
  assign n24357 = ~n24353 & n24356;
  assign n24358 = pi792 & ~n24357;
  assign n24359 = pi626 & ~n24317;
  assign n24360 = ~pi626 & ~n24205;
  assign n24361 = n17579 & ~n24360;
  assign n24362 = ~n24359 & n24361;
  assign n24363 = n17704 & n24239;
  assign n24364 = ~pi626 & ~n24317;
  assign n24365 = pi626 & ~n24205;
  assign n24366 = n17580 & ~n24365;
  assign n24367 = ~n24364 & n24366;
  assign n24368 = ~n24363 & ~n24367;
  assign n24369 = ~n24362 & n24368;
  assign n24370 = pi788 & ~n24369;
  assign n24371 = pi704 & n24276;
  assign n24372 = ~pi176 & n19236;
  assign n24373 = ~n19241 & ~n19243;
  assign n24374 = pi176 & ~n24373;
  assign n24375 = pi742 & ~n24374;
  assign n24376 = ~n24372 & n24375;
  assign n24377 = pi176 & n19253;
  assign n24378 = ~pi176 & ~n19261;
  assign n24379 = ~pi742 & ~n24378;
  assign n24380 = ~n24377 & n24379;
  assign n24381 = ~pi704 & ~n24380;
  assign n24382 = ~n24376 & n24381;
  assign n24383 = n3267 & ~n24382;
  assign n24384 = ~n24371 & n24383;
  assign n24385 = ~n24269 & ~n24384;
  assign n24386 = ~pi625 & n24385;
  assign n24387 = pi625 & n24278;
  assign n24388 = ~pi1153 & ~n24387;
  assign n24389 = ~n24386 & n24388;
  assign n24390 = ~pi608 & ~n24224;
  assign n24391 = ~n24389 & n24390;
  assign n24392 = pi625 & n24385;
  assign n24393 = ~pi625 & n24278;
  assign n24394 = pi1153 & ~n24393;
  assign n24395 = ~n24392 & n24394;
  assign n24396 = pi608 & ~n24228;
  assign n24397 = ~n24395 & n24396;
  assign n24398 = ~n24391 & ~n24397;
  assign n24399 = pi778 & ~n24398;
  assign n24400 = ~pi778 & n24385;
  assign n24401 = ~n24399 & ~n24400;
  assign n24402 = ~pi609 & ~n24401;
  assign n24403 = pi609 & n24231;
  assign n24404 = ~pi1155 & ~n24403;
  assign n24405 = ~n24402 & n24404;
  assign n24406 = ~pi660 & ~n24286;
  assign n24407 = ~n24405 & n24406;
  assign n24408 = pi609 & ~n24401;
  assign n24409 = ~pi609 & n24231;
  assign n24410 = pi1155 & ~n24409;
  assign n24411 = ~n24408 & n24410;
  assign n24412 = pi660 & ~n24290;
  assign n24413 = ~n24411 & n24412;
  assign n24414 = ~n24407 & ~n24413;
  assign n24415 = pi785 & ~n24414;
  assign n24416 = ~pi785 & ~n24401;
  assign n24417 = ~n24415 & ~n24416;
  assign n24418 = ~pi618 & ~n24417;
  assign n24419 = pi618 & n24234;
  assign n24420 = ~pi1154 & ~n24419;
  assign n24421 = ~n24418 & n24420;
  assign n24422 = ~pi627 & ~n24298;
  assign n24423 = ~n24421 & n24422;
  assign n24424 = pi618 & ~n24417;
  assign n24425 = ~pi618 & n24234;
  assign n24426 = pi1154 & ~n24425;
  assign n24427 = ~n24424 & n24426;
  assign n24428 = pi627 & ~n24302;
  assign n24429 = ~n24427 & n24428;
  assign n24430 = ~n24423 & ~n24429;
  assign n24431 = pi781 & ~n24430;
  assign n24432 = ~pi781 & ~n24417;
  assign n24433 = ~n24431 & ~n24432;
  assign n24434 = pi619 & ~n24433;
  assign n24435 = ~pi619 & ~n24237;
  assign n24436 = pi1159 & ~n24435;
  assign n24437 = ~n24434 & n24436;
  assign n24438 = pi648 & ~n24314;
  assign n24439 = ~n24437 & n24438;
  assign n24440 = ~pi619 & ~n24433;
  assign n24441 = pi619 & ~n24237;
  assign n24442 = ~pi1159 & ~n24441;
  assign n24443 = ~n24440 & n24442;
  assign n24444 = ~pi648 & ~n24310;
  assign n24445 = ~n24443 & n24444;
  assign n24446 = pi789 & ~n24445;
  assign n24447 = ~n24439 & n24446;
  assign n24448 = ~pi789 & n24433;
  assign n24449 = n17817 & ~n24448;
  assign n24450 = ~n24447 & n24449;
  assign n24451 = ~n24370 & ~n24450;
  assign n24452 = ~n24358 & ~n24451;
  assign n24453 = n20205 & n24357;
  assign n24454 = n20207 & ~n24453;
  assign n24455 = ~n24452 & n24454;
  assign n24456 = ~n24352 & ~n24455;
  assign n24457 = ~n24346 & n24456;
  assign n24458 = ~n24342 & ~n24457;
  assign n24459 = ~po1038 & ~n24458;
  assign n24460 = ~pi176 & po1038;
  assign n24461 = ~pi832 & ~n24460;
  assign n24462 = ~n24459 & n24461;
  assign po333 = ~n24204 & ~n24462;
  assign n24464 = pi177 & ~n3267;
  assign n24465 = ~pi757 & ~n19223;
  assign n24466 = ~n21480 & ~n24465;
  assign n24467 = ~pi177 & ~n24466;
  assign n24468 = ~pi177 & ~n19217;
  assign n24469 = ~pi757 & ~n24468;
  assign n24470 = ~n24271 & n24469;
  assign n24471 = ~n24467 & ~n24470;
  assign n24472 = pi686 & ~n24471;
  assign n24473 = ~pi177 & n19234;
  assign n24474 = pi177 & n19240;
  assign n24475 = ~pi38 & ~n24474;
  assign n24476 = ~n24473 & n24475;
  assign n24477 = ~pi177 & ~n17280;
  assign n24478 = n17941 & ~n24477;
  assign n24479 = pi757 & ~n24478;
  assign n24480 = ~n24476 & n24479;
  assign n24481 = pi177 & n19251;
  assign n24482 = ~n19255 & ~n19256;
  assign n24483 = ~pi177 & ~n24482;
  assign n24484 = ~pi38 & ~n24483;
  assign n24485 = ~n24481 & n24484;
  assign n24486 = ~pi177 & ~n19258;
  assign n24487 = pi177 & n19247;
  assign n24488 = pi38 & ~n24487;
  assign n24489 = ~n24486 & n24488;
  assign n24490 = ~pi757 & ~n24489;
  assign n24491 = ~n24485 & n24490;
  assign n24492 = ~n24480 & ~n24491;
  assign n24493 = ~pi686 & ~n24492;
  assign n24494 = n3267 & ~n24493;
  assign n24495 = ~n24472 & n24494;
  assign n24496 = ~n24464 & ~n24495;
  assign n24497 = ~pi625 & n24496;
  assign n24498 = n3267 & n24471;
  assign n24499 = ~n24464 & ~n24498;
  assign n24500 = pi625 & n24499;
  assign n24501 = ~pi1153 & ~n24500;
  assign n24502 = ~n24497 & n24501;
  assign n24503 = ~pi177 & n17972;
  assign n24504 = pi177 & ~n17976;
  assign n24505 = ~pi38 & ~n24504;
  assign n24506 = ~n24503 & n24505;
  assign n24507 = n17392 & ~n24477;
  assign n24508 = ~pi686 & ~n24507;
  assign n24509 = ~n24506 & n24508;
  assign n24510 = ~pi177 & pi686;
  assign n24511 = ~n17399 & n24510;
  assign n24512 = n3267 & ~n24511;
  assign n24513 = ~n24509 & n24512;
  assign n24514 = ~n24464 & ~n24513;
  assign n24515 = pi625 & n24514;
  assign n24516 = ~pi177 & ~n17406;
  assign n24517 = ~pi625 & n24516;
  assign n24518 = pi1153 & ~n24517;
  assign n24519 = ~n24515 & n24518;
  assign n24520 = ~pi608 & ~n24519;
  assign n24521 = ~n24502 & n24520;
  assign n24522 = pi625 & n24496;
  assign n24523 = ~pi625 & n24499;
  assign n24524 = pi1153 & ~n24523;
  assign n24525 = ~n24522 & n24524;
  assign n24526 = ~pi625 & n24514;
  assign n24527 = pi625 & n24516;
  assign n24528 = ~pi1153 & ~n24527;
  assign n24529 = ~n24526 & n24528;
  assign n24530 = pi608 & ~n24529;
  assign n24531 = ~n24525 & n24530;
  assign n24532 = ~n24521 & ~n24531;
  assign n24533 = pi778 & ~n24532;
  assign n24534 = ~pi778 & n24496;
  assign n24535 = ~n24533 & ~n24534;
  assign n24536 = ~pi609 & ~n24535;
  assign n24537 = ~pi778 & ~n24514;
  assign n24538 = ~n24519 & ~n24529;
  assign n24539 = pi778 & ~n24538;
  assign n24540 = ~n24537 & ~n24539;
  assign n24541 = pi609 & n24540;
  assign n24542 = ~pi1155 & ~n24541;
  assign n24543 = ~n24536 & n24542;
  assign n24544 = ~n17439 & ~n24516;
  assign n24545 = ~n17438 & ~n24499;
  assign n24546 = pi609 & n24545;
  assign n24547 = ~n24544 & ~n24546;
  assign n24548 = pi1155 & ~n24547;
  assign n24549 = ~pi660 & ~n24548;
  assign n24550 = ~n24543 & n24549;
  assign n24551 = pi609 & ~n24535;
  assign n24552 = ~pi609 & n24540;
  assign n24553 = pi1155 & ~n24552;
  assign n24554 = ~n24551 & n24553;
  assign n24555 = ~n17451 & ~n24516;
  assign n24556 = ~pi609 & n24545;
  assign n24557 = ~n24555 & ~n24556;
  assign n24558 = ~pi1155 & ~n24557;
  assign n24559 = pi660 & ~n24558;
  assign n24560 = ~n24554 & n24559;
  assign n24561 = ~n24550 & ~n24560;
  assign n24562 = pi785 & ~n24561;
  assign n24563 = ~pi785 & ~n24535;
  assign n24564 = ~n24562 & ~n24563;
  assign n24565 = ~pi618 & ~n24564;
  assign n24566 = ~n17466 & ~n24540;
  assign n24567 = n17466 & ~n24516;
  assign n24568 = ~n24566 & ~n24567;
  assign n24569 = pi618 & n24568;
  assign n24570 = ~pi1154 & ~n24569;
  assign n24571 = ~n24565 & n24570;
  assign n24572 = n17438 & ~n24516;
  assign n24573 = ~n24545 & ~n24572;
  assign n24574 = ~pi785 & ~n24573;
  assign n24575 = ~n24548 & ~n24558;
  assign n24576 = pi785 & ~n24575;
  assign n24577 = ~n24574 & ~n24576;
  assign n24578 = pi618 & n24577;
  assign n24579 = ~pi618 & n24516;
  assign n24580 = pi1154 & ~n24579;
  assign n24581 = ~n24578 & n24580;
  assign n24582 = ~pi627 & ~n24581;
  assign n24583 = ~n24571 & n24582;
  assign n24584 = pi618 & ~n24564;
  assign n24585 = ~pi618 & n24568;
  assign n24586 = pi1154 & ~n24585;
  assign n24587 = ~n24584 & n24586;
  assign n24588 = ~pi618 & n24577;
  assign n24589 = pi618 & n24516;
  assign n24590 = ~pi1154 & ~n24589;
  assign n24591 = ~n24588 & n24590;
  assign n24592 = pi627 & ~n24591;
  assign n24593 = ~n24587 & n24592;
  assign n24594 = ~n24583 & ~n24593;
  assign n24595 = pi781 & ~n24594;
  assign n24596 = ~pi781 & ~n24564;
  assign n24597 = ~n24595 & ~n24596;
  assign n24598 = ~pi619 & ~n24597;
  assign n24599 = ~n17503 & n24568;
  assign n24600 = n17503 & n24516;
  assign n24601 = ~n24599 & ~n24600;
  assign n24602 = pi619 & ~n24601;
  assign n24603 = ~pi1159 & ~n24602;
  assign n24604 = ~n24598 & n24603;
  assign n24605 = ~pi781 & ~n24577;
  assign n24606 = ~n24581 & ~n24591;
  assign n24607 = pi781 & ~n24606;
  assign n24608 = ~n24605 & ~n24607;
  assign n24609 = pi619 & n24608;
  assign n24610 = ~pi619 & n24516;
  assign n24611 = pi1159 & ~n24610;
  assign n24612 = ~n24609 & n24611;
  assign n24613 = ~pi648 & ~n24612;
  assign n24614 = ~n24604 & n24613;
  assign n24615 = pi619 & ~n24597;
  assign n24616 = ~pi619 & ~n24601;
  assign n24617 = pi1159 & ~n24616;
  assign n24618 = ~n24615 & n24617;
  assign n24619 = ~pi619 & n24608;
  assign n24620 = pi619 & n24516;
  assign n24621 = ~pi1159 & ~n24620;
  assign n24622 = ~n24619 & n24621;
  assign n24623 = pi648 & ~n24622;
  assign n24624 = ~n24618 & n24623;
  assign n24625 = ~n24614 & ~n24624;
  assign n24626 = pi789 & ~n24625;
  assign n24627 = ~pi789 & ~n24597;
  assign n24628 = ~n24626 & ~n24627;
  assign n24629 = ~pi788 & n24628;
  assign n24630 = ~pi626 & n24628;
  assign n24631 = n17539 & ~n24516;
  assign n24632 = ~n17539 & n24601;
  assign n24633 = ~n24631 & ~n24632;
  assign n24634 = pi626 & ~n24633;
  assign n24635 = ~pi641 & ~n24634;
  assign n24636 = ~n24630 & n24635;
  assign n24637 = ~pi789 & ~n24608;
  assign n24638 = ~n24612 & ~n24622;
  assign n24639 = pi789 & ~n24638;
  assign n24640 = ~n24637 & ~n24639;
  assign n24641 = ~pi626 & ~n24640;
  assign n24642 = pi626 & ~n24516;
  assign n24643 = pi641 & ~n24642;
  assign n24644 = ~n24641 & n24643;
  assign n24645 = ~pi1158 & ~n24644;
  assign n24646 = ~n24636 & n24645;
  assign n24647 = pi626 & n24628;
  assign n24648 = ~pi626 & ~n24633;
  assign n24649 = pi641 & ~n24648;
  assign n24650 = ~n24647 & n24649;
  assign n24651 = pi626 & ~n24640;
  assign n24652 = ~pi626 & ~n24516;
  assign n24653 = ~pi641 & ~n24652;
  assign n24654 = ~n24651 & n24653;
  assign n24655 = pi1158 & ~n24654;
  assign n24656 = ~n24650 & n24655;
  assign n24657 = ~n24646 & ~n24656;
  assign n24658 = pi788 & ~n24657;
  assign n24659 = ~n24629 & ~n24658;
  assign n24660 = ~pi628 & n24659;
  assign n24661 = ~n17816 & n24640;
  assign n24662 = n17816 & n24516;
  assign n24663 = ~n24661 & ~n24662;
  assign n24664 = pi628 & ~n24663;
  assign n24665 = ~pi1156 & ~n24664;
  assign n24666 = ~n24660 & n24665;
  assign n24667 = ~n17582 & n24633;
  assign n24668 = n17582 & n24516;
  assign n24669 = ~n24667 & ~n24668;
  assign n24670 = pi628 & ~n24669;
  assign n24671 = ~pi628 & n24516;
  assign n24672 = pi1156 & ~n24671;
  assign n24673 = ~n24670 & n24672;
  assign n24674 = ~pi629 & ~n24673;
  assign n24675 = ~n24666 & n24674;
  assign n24676 = pi628 & n24659;
  assign n24677 = ~pi628 & ~n24663;
  assign n24678 = pi1156 & ~n24677;
  assign n24679 = ~n24676 & n24678;
  assign n24680 = ~pi628 & ~n24669;
  assign n24681 = pi628 & n24516;
  assign n24682 = ~pi1156 & ~n24681;
  assign n24683 = ~n24680 & n24682;
  assign n24684 = pi629 & ~n24683;
  assign n24685 = ~n24679 & n24684;
  assign n24686 = ~n24675 & ~n24685;
  assign n24687 = pi792 & ~n24686;
  assign n24688 = ~pi792 & n24659;
  assign n24689 = ~n24687 & ~n24688;
  assign n24690 = ~pi647 & ~n24689;
  assign n24691 = ~n17610 & ~n24663;
  assign n24692 = n17610 & n24516;
  assign n24693 = ~n24691 & ~n24692;
  assign n24694 = pi647 & ~n24693;
  assign n24695 = ~pi1157 & ~n24694;
  assign n24696 = ~n24690 & n24695;
  assign n24697 = ~pi792 & n24669;
  assign n24698 = ~n24673 & ~n24683;
  assign n24699 = pi792 & ~n24698;
  assign n24700 = ~n24697 & ~n24699;
  assign n24701 = pi647 & n24700;
  assign n24702 = ~pi647 & n24516;
  assign n24703 = pi1157 & ~n24702;
  assign n24704 = ~n24701 & n24703;
  assign n24705 = ~pi630 & ~n24704;
  assign n24706 = ~n24696 & n24705;
  assign n24707 = pi647 & ~n24689;
  assign n24708 = ~pi647 & ~n24693;
  assign n24709 = pi1157 & ~n24708;
  assign n24710 = ~n24707 & n24709;
  assign n24711 = ~pi647 & n24700;
  assign n24712 = pi647 & n24516;
  assign n24713 = ~pi1157 & ~n24712;
  assign n24714 = ~n24711 & n24713;
  assign n24715 = pi630 & ~n24714;
  assign n24716 = ~n24710 & n24715;
  assign n24717 = ~n24706 & ~n24716;
  assign n24718 = pi787 & ~n24717;
  assign n24719 = ~pi787 & ~n24689;
  assign n24720 = ~n24718 & ~n24719;
  assign n24721 = ~pi644 & ~n24720;
  assign n24722 = ~pi787 & ~n24700;
  assign n24723 = ~n24704 & ~n24714;
  assign n24724 = pi787 & ~n24723;
  assign n24725 = ~n24722 & ~n24724;
  assign n24726 = pi644 & n24725;
  assign n24727 = ~pi715 & ~n24726;
  assign n24728 = ~n24721 & n24727;
  assign n24729 = n17652 & ~n24516;
  assign n24730 = ~n17652 & n24693;
  assign n24731 = ~n24729 & ~n24730;
  assign n24732 = ~pi644 & n24731;
  assign n24733 = pi644 & n24516;
  assign n24734 = pi715 & ~n24733;
  assign n24735 = ~n24732 & n24734;
  assign n24736 = ~pi1160 & ~n24735;
  assign n24737 = ~n24728 & n24736;
  assign n24738 = pi644 & ~n24720;
  assign n24739 = ~pi644 & n24725;
  assign n24740 = pi715 & ~n24739;
  assign n24741 = ~n24738 & n24740;
  assign n24742 = pi644 & n24731;
  assign n24743 = ~pi644 & n24516;
  assign n24744 = ~pi715 & ~n24743;
  assign n24745 = ~n24742 & n24744;
  assign n24746 = pi1160 & ~n24745;
  assign n24747 = ~n24741 & n24746;
  assign n24748 = pi790 & ~n24747;
  assign n24749 = ~n24737 & n24748;
  assign n24750 = ~pi790 & n24720;
  assign n24751 = ~po1038 & ~n24750;
  assign n24752 = ~n24749 & n24751;
  assign n24753 = ~pi177 & po1038;
  assign n24754 = ~pi832 & ~n24753;
  assign n24755 = ~n24752 & n24754;
  assign n24756 = ~pi177 & ~n2754;
  assign n24757 = ~pi757 & n16784;
  assign n24758 = ~n24756 & ~n24757;
  assign n24759 = ~n17706 & ~n24758;
  assign n24760 = ~pi785 & ~n24759;
  assign n24761 = ~n17711 & ~n24758;
  assign n24762 = pi1155 & ~n24761;
  assign n24763 = ~n17714 & n24759;
  assign n24764 = ~pi1155 & ~n24763;
  assign n24765 = ~n24762 & ~n24764;
  assign n24766 = pi785 & ~n24765;
  assign n24767 = ~n24760 & ~n24766;
  assign n24768 = ~pi781 & ~n24767;
  assign n24769 = ~n17721 & n24767;
  assign n24770 = pi1154 & ~n24769;
  assign n24771 = ~n17724 & n24767;
  assign n24772 = ~pi1154 & ~n24771;
  assign n24773 = ~n24770 & ~n24772;
  assign n24774 = pi781 & ~n24773;
  assign n24775 = ~n24768 & ~n24774;
  assign n24776 = ~pi789 & ~n24775;
  assign n24777 = pi619 & n24775;
  assign n24778 = ~pi619 & n24756;
  assign n24779 = pi1159 & ~n24778;
  assign n24780 = ~n24777 & n24779;
  assign n24781 = ~pi619 & n24775;
  assign n24782 = pi619 & n24756;
  assign n24783 = ~pi1159 & ~n24782;
  assign n24784 = ~n24781 & n24783;
  assign n24785 = ~n24780 & ~n24784;
  assign n24786 = pi789 & ~n24785;
  assign n24787 = ~n24776 & ~n24786;
  assign n24788 = ~n17816 & n24787;
  assign n24789 = n17816 & n24756;
  assign n24790 = ~n24788 & ~n24789;
  assign n24791 = ~n17610 & ~n24790;
  assign n24792 = n17610 & n24756;
  assign n24793 = ~n24791 & ~n24792;
  assign n24794 = ~n20398 & n24793;
  assign n24795 = ~pi686 & n16786;
  assign n24796 = ~n24756 & ~n24795;
  assign n24797 = ~pi778 & n24796;
  assign n24798 = ~pi625 & n24795;
  assign n24799 = ~n24796 & ~n24798;
  assign n24800 = pi1153 & ~n24799;
  assign n24801 = ~pi1153 & ~n24756;
  assign n24802 = ~n24798 & n24801;
  assign n24803 = ~n24800 & ~n24802;
  assign n24804 = pi778 & ~n24803;
  assign n24805 = ~n24797 & ~n24804;
  assign n24806 = ~n17692 & n24805;
  assign n24807 = ~n17694 & n24806;
  assign n24808 = ~n17696 & n24807;
  assign n24809 = ~n17828 & n24808;
  assign n24810 = ~n17859 & n24809;
  assign n24811 = ~pi647 & n24810;
  assign n24812 = pi647 & n24756;
  assign n24813 = ~pi1157 & ~n24812;
  assign n24814 = ~n24811 & n24813;
  assign n24815 = pi647 & ~n24810;
  assign n24816 = ~pi647 & ~n24756;
  assign n24817 = ~n24815 & ~n24816;
  assign n24818 = pi1157 & ~n24817;
  assign n24819 = ~n24814 & ~n24818;
  assign n24820 = ~n17651 & ~n24819;
  assign n24821 = ~n24794 & ~n24820;
  assign n24822 = pi787 & ~n24821;
  assign n24823 = pi626 & ~n24787;
  assign n24824 = ~pi626 & ~n24756;
  assign n24825 = n17579 & ~n24824;
  assign n24826 = ~n24823 & n24825;
  assign n24827 = n17704 & n24808;
  assign n24828 = ~pi626 & ~n24787;
  assign n24829 = pi626 & ~n24756;
  assign n24830 = n17580 & ~n24829;
  assign n24831 = ~n24828 & n24830;
  assign n24832 = ~n24827 & ~n24831;
  assign n24833 = ~n24826 & n24832;
  assign n24834 = pi788 & ~n24833;
  assign n24835 = ~n16521 & ~n24796;
  assign n24836 = pi625 & n24835;
  assign n24837 = n24758 & ~n24835;
  assign n24838 = ~n24836 & ~n24837;
  assign n24839 = n24801 & ~n24838;
  assign n24840 = ~pi608 & ~n24800;
  assign n24841 = ~n24839 & n24840;
  assign n24842 = pi1153 & n24758;
  assign n24843 = ~n24836 & n24842;
  assign n24844 = pi608 & ~n24802;
  assign n24845 = ~n24843 & n24844;
  assign n24846 = ~n24841 & ~n24845;
  assign n24847 = pi778 & ~n24846;
  assign n24848 = ~pi778 & ~n24837;
  assign n24849 = ~n24847 & ~n24848;
  assign n24850 = ~pi609 & ~n24849;
  assign n24851 = pi609 & n24805;
  assign n24852 = ~pi1155 & ~n24851;
  assign n24853 = ~n24850 & n24852;
  assign n24854 = ~pi660 & ~n24762;
  assign n24855 = ~n24853 & n24854;
  assign n24856 = pi609 & ~n24849;
  assign n24857 = ~pi609 & n24805;
  assign n24858 = pi1155 & ~n24857;
  assign n24859 = ~n24856 & n24858;
  assign n24860 = pi660 & ~n24764;
  assign n24861 = ~n24859 & n24860;
  assign n24862 = ~n24855 & ~n24861;
  assign n24863 = pi785 & ~n24862;
  assign n24864 = ~pi785 & ~n24849;
  assign n24865 = ~n24863 & ~n24864;
  assign n24866 = ~pi618 & ~n24865;
  assign n24867 = pi618 & n24806;
  assign n24868 = ~pi1154 & ~n24867;
  assign n24869 = ~n24866 & n24868;
  assign n24870 = ~pi627 & ~n24770;
  assign n24871 = ~n24869 & n24870;
  assign n24872 = pi618 & ~n24865;
  assign n24873 = ~pi618 & n24806;
  assign n24874 = pi1154 & ~n24873;
  assign n24875 = ~n24872 & n24874;
  assign n24876 = pi627 & ~n24772;
  assign n24877 = ~n24875 & n24876;
  assign n24878 = ~n24871 & ~n24877;
  assign n24879 = pi781 & ~n24878;
  assign n24880 = ~pi781 & ~n24865;
  assign n24881 = ~n24879 & ~n24880;
  assign n24882 = pi619 & ~n24881;
  assign n24883 = ~pi619 & n24807;
  assign n24884 = pi1159 & ~n24883;
  assign n24885 = ~n24882 & n24884;
  assign n24886 = pi648 & ~n24784;
  assign n24887 = ~n24885 & n24886;
  assign n24888 = ~pi619 & ~n24881;
  assign n24889 = pi619 & n24807;
  assign n24890 = ~pi1159 & ~n24889;
  assign n24891 = ~n24888 & n24890;
  assign n24892 = ~pi648 & ~n24780;
  assign n24893 = ~n24891 & n24892;
  assign n24894 = pi789 & ~n24893;
  assign n24895 = ~n24887 & n24894;
  assign n24896 = ~pi789 & n24881;
  assign n24897 = n17817 & ~n24896;
  assign n24898 = ~n24895 & n24897;
  assign n24899 = ~n24834 & ~n24898;
  assign n24900 = ~n20205 & ~n24899;
  assign n24901 = n17856 & ~n24790;
  assign n24902 = n20693 & n24809;
  assign n24903 = ~n24901 & ~n24902;
  assign n24904 = ~pi629 & ~n24903;
  assign n24905 = n20697 & n24809;
  assign n24906 = n17855 & ~n24790;
  assign n24907 = ~n24905 & ~n24906;
  assign n24908 = pi629 & ~n24907;
  assign n24909 = ~n24904 & ~n24908;
  assign n24910 = pi792 & ~n24909;
  assign n24911 = n20207 & ~n24910;
  assign n24912 = ~n24900 & n24911;
  assign n24913 = ~n24822 & ~n24912;
  assign n24914 = pi644 & n24913;
  assign n24915 = ~pi787 & ~n24810;
  assign n24916 = pi787 & ~n24819;
  assign n24917 = ~n24915 & ~n24916;
  assign n24918 = ~pi644 & n24917;
  assign n24919 = pi715 & ~n24918;
  assign n24920 = ~n24914 & n24919;
  assign n24921 = ~n17652 & ~n24793;
  assign n24922 = n17652 & n24756;
  assign n24923 = ~n24921 & ~n24922;
  assign n24924 = pi644 & ~n24923;
  assign n24925 = ~pi644 & n24756;
  assign n24926 = ~pi715 & ~n24925;
  assign n24927 = ~n24924 & n24926;
  assign n24928 = pi1160 & ~n24927;
  assign n24929 = ~n24920 & n24928;
  assign n24930 = ~pi644 & n24913;
  assign n24931 = pi644 & n24917;
  assign n24932 = ~pi715 & ~n24931;
  assign n24933 = ~n24930 & n24932;
  assign n24934 = ~pi644 & ~n24923;
  assign n24935 = pi644 & n24756;
  assign n24936 = pi715 & ~n24935;
  assign n24937 = ~n24934 & n24936;
  assign n24938 = ~pi1160 & ~n24937;
  assign n24939 = ~n24933 & n24938;
  assign n24940 = ~n24929 & ~n24939;
  assign n24941 = pi790 & ~n24940;
  assign n24942 = ~pi790 & n24913;
  assign n24943 = pi832 & ~n24942;
  assign n24944 = ~n24941 & n24943;
  assign po334 = ~n24755 & ~n24944;
  assign n24946 = ~pi178 & ~n2754;
  assign n24947 = ~pi760 & n16784;
  assign n24948 = ~n24946 & ~n24947;
  assign n24949 = ~n17706 & ~n24948;
  assign n24950 = ~pi785 & ~n24949;
  assign n24951 = n17451 & n24947;
  assign n24952 = n24949 & ~n24951;
  assign n24953 = pi1155 & ~n24952;
  assign n24954 = ~pi1155 & ~n24946;
  assign n24955 = ~n24951 & n24954;
  assign n24956 = ~n24953 & ~n24955;
  assign n24957 = pi785 & ~n24956;
  assign n24958 = ~n24950 & ~n24957;
  assign n24959 = ~pi781 & ~n24958;
  assign n24960 = ~n17721 & n24958;
  assign n24961 = pi1154 & ~n24960;
  assign n24962 = ~n17724 & n24958;
  assign n24963 = ~pi1154 & ~n24962;
  assign n24964 = ~n24961 & ~n24963;
  assign n24965 = pi781 & ~n24964;
  assign n24966 = ~n24959 & ~n24965;
  assign n24967 = ~pi789 & ~n24966;
  assign n24968 = ~n22890 & n24966;
  assign n24969 = pi1159 & ~n24968;
  assign n24970 = ~n22893 & n24966;
  assign n24971 = ~pi1159 & ~n24970;
  assign n24972 = ~n24969 & ~n24971;
  assign n24973 = pi789 & ~n24972;
  assign n24974 = ~n24967 & ~n24973;
  assign n24975 = ~n17816 & n24974;
  assign n24976 = n17816 & n24946;
  assign n24977 = ~n24975 & ~n24976;
  assign n24978 = ~n17610 & ~n24977;
  assign n24979 = n17610 & n24946;
  assign n24980 = ~n24978 & ~n24979;
  assign n24981 = ~n20398 & n24980;
  assign n24982 = ~pi688 & n16786;
  assign n24983 = ~n24946 & ~n24982;
  assign n24984 = ~pi778 & ~n24983;
  assign n24985 = ~pi625 & n24982;
  assign n24986 = ~n24983 & ~n24985;
  assign n24987 = pi1153 & ~n24986;
  assign n24988 = ~pi1153 & ~n24946;
  assign n24989 = ~n24985 & n24988;
  assign n24990 = pi778 & ~n24989;
  assign n24991 = ~n24987 & n24990;
  assign n24992 = ~n24984 & ~n24991;
  assign n24993 = ~n17692 & ~n24992;
  assign n24994 = ~n17694 & n24993;
  assign n24995 = ~n17696 & n24994;
  assign n24996 = ~n17828 & n24995;
  assign n24997 = ~n17859 & n24996;
  assign n24998 = ~pi647 & n24997;
  assign n24999 = pi647 & n24946;
  assign n25000 = ~pi1157 & ~n24999;
  assign n25001 = ~n24998 & n25000;
  assign n25002 = pi647 & ~n24997;
  assign n25003 = ~pi647 & ~n24946;
  assign n25004 = ~n25002 & ~n25003;
  assign n25005 = pi1157 & ~n25004;
  assign n25006 = ~n25001 & ~n25005;
  assign n25007 = ~n17651 & ~n25006;
  assign n25008 = ~n24981 & ~n25007;
  assign n25009 = pi787 & ~n25008;
  assign n25010 = pi626 & ~n24974;
  assign n25011 = ~pi626 & ~n24946;
  assign n25012 = n17579 & ~n25011;
  assign n25013 = ~n25010 & n25012;
  assign n25014 = n17704 & n24995;
  assign n25015 = ~pi626 & ~n24974;
  assign n25016 = pi626 & ~n24946;
  assign n25017 = n17580 & ~n25016;
  assign n25018 = ~n25015 & n25017;
  assign n25019 = ~n25014 & ~n25018;
  assign n25020 = ~n25013 & n25019;
  assign n25021 = pi788 & ~n25020;
  assign n25022 = ~n16521 & ~n24983;
  assign n25023 = pi625 & n25022;
  assign n25024 = n24948 & ~n25022;
  assign n25025 = ~n25023 & ~n25024;
  assign n25026 = n24988 & ~n25025;
  assign n25027 = ~pi608 & ~n24987;
  assign n25028 = ~n25026 & n25027;
  assign n25029 = pi1153 & n24948;
  assign n25030 = ~n25023 & n25029;
  assign n25031 = pi608 & ~n24989;
  assign n25032 = ~n25030 & n25031;
  assign n25033 = ~n25028 & ~n25032;
  assign n25034 = pi778 & ~n25033;
  assign n25035 = ~pi778 & ~n25024;
  assign n25036 = ~n25034 & ~n25035;
  assign n25037 = ~pi609 & ~n25036;
  assign n25038 = pi609 & ~n24992;
  assign n25039 = ~pi1155 & ~n25038;
  assign n25040 = ~n25037 & n25039;
  assign n25041 = ~pi660 & ~n24953;
  assign n25042 = ~n25040 & n25041;
  assign n25043 = pi609 & ~n25036;
  assign n25044 = ~pi609 & ~n24992;
  assign n25045 = pi1155 & ~n25044;
  assign n25046 = ~n25043 & n25045;
  assign n25047 = pi660 & ~n24955;
  assign n25048 = ~n25046 & n25047;
  assign n25049 = ~n25042 & ~n25048;
  assign n25050 = pi785 & ~n25049;
  assign n25051 = ~pi785 & ~n25036;
  assign n25052 = ~n25050 & ~n25051;
  assign n25053 = ~pi618 & ~n25052;
  assign n25054 = pi618 & n24993;
  assign n25055 = ~pi1154 & ~n25054;
  assign n25056 = ~n25053 & n25055;
  assign n25057 = ~pi627 & ~n24961;
  assign n25058 = ~n25056 & n25057;
  assign n25059 = pi618 & ~n25052;
  assign n25060 = ~pi618 & n24993;
  assign n25061 = pi1154 & ~n25060;
  assign n25062 = ~n25059 & n25061;
  assign n25063 = pi627 & ~n24963;
  assign n25064 = ~n25062 & n25063;
  assign n25065 = ~n25058 & ~n25064;
  assign n25066 = pi781 & ~n25065;
  assign n25067 = ~pi781 & ~n25052;
  assign n25068 = ~n25066 & ~n25067;
  assign n25069 = pi619 & ~n25068;
  assign n25070 = ~pi619 & n24994;
  assign n25071 = pi1159 & ~n25070;
  assign n25072 = ~n25069 & n25071;
  assign n25073 = pi648 & ~n24971;
  assign n25074 = ~n25072 & n25073;
  assign n25075 = ~pi619 & ~n25068;
  assign n25076 = pi619 & n24994;
  assign n25077 = ~pi1159 & ~n25076;
  assign n25078 = ~n25075 & n25077;
  assign n25079 = ~pi648 & ~n24969;
  assign n25080 = ~n25078 & n25079;
  assign n25081 = pi789 & ~n25080;
  assign n25082 = ~n25074 & n25081;
  assign n25083 = ~pi789 & n25068;
  assign n25084 = n17817 & ~n25083;
  assign n25085 = ~n25082 & n25084;
  assign n25086 = ~n25021 & ~n25085;
  assign n25087 = ~n20205 & ~n25086;
  assign n25088 = n17856 & ~n24977;
  assign n25089 = n20693 & n24996;
  assign n25090 = ~n25088 & ~n25089;
  assign n25091 = ~pi629 & ~n25090;
  assign n25092 = n20697 & n24996;
  assign n25093 = n17855 & ~n24977;
  assign n25094 = ~n25092 & ~n25093;
  assign n25095 = pi629 & ~n25094;
  assign n25096 = ~n25091 & ~n25095;
  assign n25097 = pi792 & ~n25096;
  assign n25098 = n20207 & ~n25097;
  assign n25099 = ~n25087 & n25098;
  assign n25100 = ~n25009 & ~n25099;
  assign n25101 = pi644 & n25100;
  assign n25102 = ~pi787 & ~n24997;
  assign n25103 = pi787 & ~n25006;
  assign n25104 = ~n25102 & ~n25103;
  assign n25105 = ~pi644 & n25104;
  assign n25106 = pi715 & ~n25105;
  assign n25107 = ~n25101 & n25106;
  assign n25108 = ~n17652 & ~n24980;
  assign n25109 = n17652 & n24946;
  assign n25110 = ~n25108 & ~n25109;
  assign n25111 = pi644 & ~n25110;
  assign n25112 = ~pi644 & n24946;
  assign n25113 = ~pi715 & ~n25112;
  assign n25114 = ~n25111 & n25113;
  assign n25115 = pi1160 & ~n25114;
  assign n25116 = ~n25107 & n25115;
  assign n25117 = ~pi644 & n25100;
  assign n25118 = pi644 & n25104;
  assign n25119 = ~pi715 & ~n25118;
  assign n25120 = ~n25117 & n25119;
  assign n25121 = ~pi644 & ~n25110;
  assign n25122 = pi644 & n24946;
  assign n25123 = pi715 & ~n25122;
  assign n25124 = ~n25121 & n25123;
  assign n25125 = ~pi1160 & ~n25124;
  assign n25126 = ~n25120 & n25125;
  assign n25127 = ~n25116 & ~n25126;
  assign n25128 = pi790 & ~n25127;
  assign n25129 = ~pi790 & n25100;
  assign n25130 = pi832 & ~n25129;
  assign n25131 = ~n25128 & n25130;
  assign n25132 = ~pi178 & ~n17406;
  assign n25133 = n17539 & ~n25132;
  assign n25134 = ~pi688 & n3267;
  assign n25135 = n25132 & ~n25134;
  assign n25136 = pi178 & ~n17976;
  assign n25137 = ~pi38 & ~n25136;
  assign n25138 = n3267 & ~n25137;
  assign n25139 = ~pi178 & n17972;
  assign n25140 = ~n25138 & ~n25139;
  assign n25141 = ~pi178 & ~n17280;
  assign n25142 = n17392 & ~n25141;
  assign n25143 = ~pi688 & ~n25142;
  assign n25144 = ~n25140 & n25143;
  assign n25145 = ~n25135 & ~n25144;
  assign n25146 = ~pi778 & n25145;
  assign n25147 = pi625 & ~n25145;
  assign n25148 = ~pi625 & n25132;
  assign n25149 = pi1153 & ~n25148;
  assign n25150 = ~n25147 & n25149;
  assign n25151 = ~pi625 & ~n25145;
  assign n25152 = pi625 & n25132;
  assign n25153 = ~pi1153 & ~n25152;
  assign n25154 = ~n25151 & n25153;
  assign n25155 = ~n25150 & ~n25154;
  assign n25156 = pi778 & ~n25155;
  assign n25157 = ~n25146 & ~n25156;
  assign n25158 = ~n17466 & ~n25157;
  assign n25159 = n17466 & ~n25132;
  assign n25160 = ~n25158 & ~n25159;
  assign n25161 = ~n17503 & n25160;
  assign n25162 = n17503 & n25132;
  assign n25163 = ~n25161 & ~n25162;
  assign n25164 = ~n17539 & n25163;
  assign n25165 = ~n25133 & ~n25164;
  assign n25166 = ~n17582 & n25165;
  assign n25167 = n17582 & n25132;
  assign n25168 = ~n25166 & ~n25167;
  assign n25169 = ~pi792 & n25168;
  assign n25170 = pi628 & ~n25168;
  assign n25171 = ~pi628 & n25132;
  assign n25172 = pi1156 & ~n25171;
  assign n25173 = ~n25170 & n25172;
  assign n25174 = ~pi628 & ~n25168;
  assign n25175 = pi628 & n25132;
  assign n25176 = ~pi1156 & ~n25175;
  assign n25177 = ~n25174 & n25176;
  assign n25178 = ~n25173 & ~n25177;
  assign n25179 = pi792 & ~n25178;
  assign n25180 = ~n25169 & ~n25179;
  assign n25181 = ~pi647 & ~n25180;
  assign n25182 = pi647 & ~n25132;
  assign n25183 = ~n25181 & ~n25182;
  assign n25184 = ~pi1157 & n25183;
  assign n25185 = pi647 & ~n25180;
  assign n25186 = ~pi647 & ~n25132;
  assign n25187 = ~n25185 & ~n25186;
  assign n25188 = pi1157 & n25187;
  assign n25189 = ~n25184 & ~n25188;
  assign n25190 = pi787 & ~n25189;
  assign n25191 = ~pi787 & n25180;
  assign n25192 = ~n25190 & ~n25191;
  assign n25193 = ~pi644 & ~n25192;
  assign n25194 = pi715 & ~n25193;
  assign n25195 = pi178 & ~n3267;
  assign n25196 = ~pi760 & n17282;
  assign n25197 = ~n25141 & ~n25196;
  assign n25198 = pi38 & ~n25197;
  assign n25199 = ~pi178 & n17242;
  assign n25200 = pi178 & ~n17275;
  assign n25201 = ~pi760 & ~n25200;
  assign n25202 = ~n25199 & n25201;
  assign n25203 = ~pi178 & pi760;
  assign n25204 = ~n17201 & n25203;
  assign n25205 = ~n25202 & ~n25204;
  assign n25206 = ~pi38 & ~n25205;
  assign n25207 = ~n25198 & ~n25206;
  assign n25208 = n3267 & n25207;
  assign n25209 = ~n25195 & ~n25208;
  assign n25210 = ~n17438 & ~n25209;
  assign n25211 = n17438 & ~n25132;
  assign n25212 = ~n25210 & ~n25211;
  assign n25213 = ~pi785 & ~n25212;
  assign n25214 = ~n17439 & ~n25132;
  assign n25215 = pi609 & n25210;
  assign n25216 = ~n25214 & ~n25215;
  assign n25217 = pi1155 & ~n25216;
  assign n25218 = ~n17451 & ~n25132;
  assign n25219 = ~pi609 & n25210;
  assign n25220 = ~n25218 & ~n25219;
  assign n25221 = ~pi1155 & ~n25220;
  assign n25222 = ~n25217 & ~n25221;
  assign n25223 = pi785 & ~n25222;
  assign n25224 = ~n25213 & ~n25223;
  assign n25225 = ~pi781 & ~n25224;
  assign n25226 = pi618 & n25224;
  assign n25227 = ~pi618 & n25132;
  assign n25228 = pi1154 & ~n25227;
  assign n25229 = ~n25226 & n25228;
  assign n25230 = ~pi618 & n25224;
  assign n25231 = pi618 & n25132;
  assign n25232 = ~pi1154 & ~n25231;
  assign n25233 = ~n25230 & n25232;
  assign n25234 = ~n25229 & ~n25233;
  assign n25235 = pi781 & ~n25234;
  assign n25236 = ~n25225 & ~n25235;
  assign n25237 = ~pi789 & ~n25236;
  assign n25238 = pi619 & n25236;
  assign n25239 = ~pi619 & n25132;
  assign n25240 = pi1159 & ~n25239;
  assign n25241 = ~n25238 & n25240;
  assign n25242 = ~pi619 & n25236;
  assign n25243 = pi619 & n25132;
  assign n25244 = ~pi1159 & ~n25243;
  assign n25245 = ~n25242 & n25244;
  assign n25246 = ~n25241 & ~n25245;
  assign n25247 = pi789 & ~n25246;
  assign n25248 = ~n25237 & ~n25247;
  assign n25249 = ~n17816 & n25248;
  assign n25250 = n17816 & n25132;
  assign n25251 = ~n25249 & ~n25250;
  assign n25252 = ~n17610 & ~n25251;
  assign n25253 = n17610 & n25132;
  assign n25254 = ~n25252 & ~n25253;
  assign n25255 = ~n17652 & ~n25254;
  assign n25256 = n17652 & n25132;
  assign n25257 = ~n25255 & ~n25256;
  assign n25258 = pi644 & ~n25257;
  assign n25259 = ~pi644 & n25132;
  assign n25260 = ~pi715 & ~n25259;
  assign n25261 = ~n25258 & n25260;
  assign n25262 = pi1160 & ~n25261;
  assign n25263 = ~n25194 & n25262;
  assign n25264 = pi644 & ~n25192;
  assign n25265 = ~pi715 & ~n25264;
  assign n25266 = ~pi644 & ~n25257;
  assign n25267 = pi644 & n25132;
  assign n25268 = pi715 & ~n25267;
  assign n25269 = ~n25266 & n25268;
  assign n25270 = ~pi1160 & ~n25269;
  assign n25271 = ~n25265 & n25270;
  assign n25272 = ~n25263 & ~n25271;
  assign n25273 = pi790 & ~n25272;
  assign n25274 = pi644 & n25262;
  assign n25275 = ~pi644 & n25270;
  assign n25276 = pi790 & ~n25275;
  assign n25277 = ~n25274 & n25276;
  assign n25278 = ~n20409 & n25251;
  assign n25279 = ~pi629 & n25173;
  assign n25280 = pi629 & n25177;
  assign n25281 = ~n25279 & ~n25280;
  assign n25282 = ~n25278 & n25281;
  assign n25283 = pi792 & ~n25282;
  assign n25284 = pi688 & ~n25207;
  assign n25285 = ~pi178 & n16687;
  assign n25286 = pi178 & n16799;
  assign n25287 = pi760 & ~n25286;
  assign n25288 = ~n25285 & n25287;
  assign n25289 = pi178 & n16879;
  assign n25290 = ~pi178 & ~n16944;
  assign n25291 = ~pi760 & ~n25290;
  assign n25292 = ~n25289 & n25291;
  assign n25293 = pi39 & ~n25292;
  assign n25294 = ~n25288 & n25293;
  assign n25295 = ~pi178 & ~n17088;
  assign n25296 = pi178 & ~n17059;
  assign n25297 = pi760 & ~n25296;
  assign n25298 = ~n25295 & n25297;
  assign n25299 = ~pi178 & n17092;
  assign n25300 = pi178 & n17094;
  assign n25301 = ~pi760 & ~n25300;
  assign n25302 = ~n25299 & n25301;
  assign n25303 = ~n25298 & ~n25302;
  assign n25304 = ~pi39 & ~n25303;
  assign n25305 = ~pi38 & ~n25304;
  assign n25306 = ~n25294 & n25305;
  assign n25307 = ~pi760 & ~n16905;
  assign n25308 = n19230 & ~n25307;
  assign n25309 = ~pi178 & ~n25308;
  assign n25310 = ~n16787 & ~n24947;
  assign n25311 = pi178 & ~n25310;
  assign n25312 = n6234 & n25311;
  assign n25313 = pi38 & ~n25312;
  assign n25314 = ~n25309 & n25313;
  assign n25315 = ~pi688 & ~n25314;
  assign n25316 = ~n25306 & n25315;
  assign n25317 = n3267 & ~n25316;
  assign n25318 = ~n25284 & n25317;
  assign n25319 = ~n25195 & ~n25318;
  assign n25320 = ~pi625 & n25319;
  assign n25321 = pi625 & n25209;
  assign n25322 = ~pi1153 & ~n25321;
  assign n25323 = ~n25320 & n25322;
  assign n25324 = ~pi608 & ~n25150;
  assign n25325 = ~n25323 & n25324;
  assign n25326 = pi625 & n25319;
  assign n25327 = ~pi625 & n25209;
  assign n25328 = pi1153 & ~n25327;
  assign n25329 = ~n25326 & n25328;
  assign n25330 = pi608 & ~n25154;
  assign n25331 = ~n25329 & n25330;
  assign n25332 = ~n25325 & ~n25331;
  assign n25333 = pi778 & ~n25332;
  assign n25334 = ~pi778 & n25319;
  assign n25335 = ~n25333 & ~n25334;
  assign n25336 = ~pi609 & ~n25335;
  assign n25337 = pi609 & n25157;
  assign n25338 = ~pi1155 & ~n25337;
  assign n25339 = ~n25336 & n25338;
  assign n25340 = ~pi660 & ~n25217;
  assign n25341 = ~n25339 & n25340;
  assign n25342 = pi609 & ~n25335;
  assign n25343 = ~pi609 & n25157;
  assign n25344 = pi1155 & ~n25343;
  assign n25345 = ~n25342 & n25344;
  assign n25346 = pi660 & ~n25221;
  assign n25347 = ~n25345 & n25346;
  assign n25348 = ~n25341 & ~n25347;
  assign n25349 = pi785 & ~n25348;
  assign n25350 = ~pi785 & ~n25335;
  assign n25351 = ~n25349 & ~n25350;
  assign n25352 = ~pi618 & ~n25351;
  assign n25353 = pi618 & n25160;
  assign n25354 = ~pi1154 & ~n25353;
  assign n25355 = ~n25352 & n25354;
  assign n25356 = ~pi627 & ~n25229;
  assign n25357 = ~n25355 & n25356;
  assign n25358 = pi618 & ~n25351;
  assign n25359 = ~pi618 & n25160;
  assign n25360 = pi1154 & ~n25359;
  assign n25361 = ~n25358 & n25360;
  assign n25362 = pi627 & ~n25233;
  assign n25363 = ~n25361 & n25362;
  assign n25364 = ~n25357 & ~n25363;
  assign n25365 = pi781 & ~n25364;
  assign n25366 = ~pi781 & ~n25351;
  assign n25367 = ~n25365 & ~n25366;
  assign n25368 = pi619 & ~n25367;
  assign n25369 = ~pi619 & ~n25163;
  assign n25370 = pi1159 & ~n25369;
  assign n25371 = ~n25368 & n25370;
  assign n25372 = pi648 & ~n25245;
  assign n25373 = ~n25371 & n25372;
  assign n25374 = ~pi619 & ~n25367;
  assign n25375 = pi619 & ~n25163;
  assign n25376 = ~pi1159 & ~n25375;
  assign n25377 = ~n25374 & n25376;
  assign n25378 = ~pi648 & ~n25241;
  assign n25379 = ~n25377 & n25378;
  assign n25380 = pi789 & ~n25379;
  assign n25381 = ~n25373 & n25380;
  assign n25382 = ~pi789 & n25367;
  assign n25383 = n17817 & ~n25382;
  assign n25384 = ~n25381 & n25383;
  assign n25385 = pi626 & ~n25248;
  assign n25386 = ~pi626 & ~n25132;
  assign n25387 = n17579 & ~n25386;
  assign n25388 = ~n25385 & n25387;
  assign n25389 = n17704 & n25165;
  assign n25390 = ~pi626 & ~n25248;
  assign n25391 = pi626 & ~n25132;
  assign n25392 = n17580 & ~n25391;
  assign n25393 = ~n25390 & n25392;
  assign n25394 = ~n25389 & ~n25393;
  assign n25395 = ~n25388 & n25394;
  assign n25396 = pi788 & ~n25395;
  assign n25397 = ~n20205 & ~n25396;
  assign n25398 = ~n25384 & n25397;
  assign n25399 = ~n25283 & ~n25398;
  assign n25400 = n20207 & ~n25399;
  assign n25401 = ~n20398 & n25254;
  assign n25402 = n17650 & ~n25183;
  assign n25403 = n17649 & ~n25187;
  assign n25404 = ~n25402 & ~n25403;
  assign n25405 = ~n25401 & n25404;
  assign n25406 = pi787 & ~n25405;
  assign n25407 = ~n25400 & ~n25406;
  assign n25408 = ~n25277 & n25407;
  assign n25409 = ~n25273 & ~n25408;
  assign n25410 = ~po1038 & ~n25409;
  assign n25411 = ~pi178 & po1038;
  assign n25412 = ~pi832 & ~n25411;
  assign n25413 = ~n25410 & n25412;
  assign po335 = ~n25131 & ~n25413;
  assign n25415 = pi179 & ~n3267;
  assign n25416 = ~pi179 & ~n17280;
  assign n25417 = n17941 & ~n25416;
  assign n25418 = ~pi179 & n16687;
  assign n25419 = pi179 & n16799;
  assign n25420 = pi39 & ~n25419;
  assign n25421 = ~n25418 & n25420;
  assign n25422 = pi179 & n17059;
  assign n25423 = ~pi179 & n17088;
  assign n25424 = ~pi39 & ~n25423;
  assign n25425 = ~n25422 & n25424;
  assign n25426 = ~n25421 & ~n25425;
  assign n25427 = ~pi38 & ~n25426;
  assign n25428 = ~n25417 & ~n25427;
  assign n25429 = pi741 & ~n25428;
  assign n25430 = pi179 & n19253;
  assign n25431 = ~pi179 & ~n19261;
  assign n25432 = ~pi741 & ~n25431;
  assign n25433 = ~n25430 & n25432;
  assign n25434 = ~pi724 & ~n25433;
  assign n25435 = ~n25429 & n25434;
  assign n25436 = ~pi741 & ~n24271;
  assign n25437 = pi179 & ~n25436;
  assign n25438 = ~pi179 & ~pi741;
  assign n25439 = ~n19217 & n25438;
  assign n25440 = n19223 & n25439;
  assign n25441 = ~n25437 & ~n25440;
  assign n25442 = ~n21508 & n25441;
  assign n25443 = n3267 & ~n25442;
  assign n25444 = ~pi724 & n3267;
  assign n25445 = ~n25443 & ~n25444;
  assign n25446 = ~n25435 & ~n25445;
  assign n25447 = ~n25415 & ~n25446;
  assign n25448 = ~pi625 & n25447;
  assign n25449 = ~n25415 & ~n25443;
  assign n25450 = pi625 & n25449;
  assign n25451 = ~pi1153 & ~n25450;
  assign n25452 = ~n25448 & n25451;
  assign n25453 = ~pi179 & ~n17406;
  assign n25454 = ~n25444 & n25453;
  assign n25455 = ~pi179 & n17972;
  assign n25456 = pi179 & ~n17976;
  assign n25457 = ~pi38 & ~n25456;
  assign n25458 = n3267 & ~n25457;
  assign n25459 = ~n25455 & ~n25458;
  assign n25460 = n17392 & ~n25416;
  assign n25461 = ~pi724 & ~n25460;
  assign n25462 = ~n25459 & n25461;
  assign n25463 = ~n25454 & ~n25462;
  assign n25464 = pi625 & ~n25463;
  assign n25465 = ~pi625 & n25453;
  assign n25466 = pi1153 & ~n25465;
  assign n25467 = ~n25464 & n25466;
  assign n25468 = ~pi608 & ~n25467;
  assign n25469 = ~n25452 & n25468;
  assign n25470 = pi625 & n25447;
  assign n25471 = ~pi625 & n25449;
  assign n25472 = pi1153 & ~n25471;
  assign n25473 = ~n25470 & n25472;
  assign n25474 = ~pi625 & ~n25463;
  assign n25475 = pi625 & n25453;
  assign n25476 = ~pi1153 & ~n25475;
  assign n25477 = ~n25474 & n25476;
  assign n25478 = pi608 & ~n25477;
  assign n25479 = ~n25473 & n25478;
  assign n25480 = ~n25469 & ~n25479;
  assign n25481 = pi778 & ~n25480;
  assign n25482 = ~pi778 & n25447;
  assign n25483 = ~n25481 & ~n25482;
  assign n25484 = ~pi609 & ~n25483;
  assign n25485 = ~pi778 & n25463;
  assign n25486 = ~n25467 & ~n25477;
  assign n25487 = pi778 & ~n25486;
  assign n25488 = ~n25485 & ~n25487;
  assign n25489 = pi609 & n25488;
  assign n25490 = ~pi1155 & ~n25489;
  assign n25491 = ~n25484 & n25490;
  assign n25492 = ~n17439 & ~n25453;
  assign n25493 = ~n17438 & ~n25449;
  assign n25494 = pi609 & n25493;
  assign n25495 = ~n25492 & ~n25494;
  assign n25496 = pi1155 & ~n25495;
  assign n25497 = ~pi660 & ~n25496;
  assign n25498 = ~n25491 & n25497;
  assign n25499 = pi609 & ~n25483;
  assign n25500 = ~pi609 & n25488;
  assign n25501 = pi1155 & ~n25500;
  assign n25502 = ~n25499 & n25501;
  assign n25503 = ~n17451 & ~n25453;
  assign n25504 = ~pi609 & n25493;
  assign n25505 = ~n25503 & ~n25504;
  assign n25506 = ~pi1155 & ~n25505;
  assign n25507 = pi660 & ~n25506;
  assign n25508 = ~n25502 & n25507;
  assign n25509 = ~n25498 & ~n25508;
  assign n25510 = pi785 & ~n25509;
  assign n25511 = ~pi785 & ~n25483;
  assign n25512 = ~n25510 & ~n25511;
  assign n25513 = ~pi618 & ~n25512;
  assign n25514 = ~n17466 & ~n25488;
  assign n25515 = n17466 & ~n25453;
  assign n25516 = ~n25514 & ~n25515;
  assign n25517 = pi618 & n25516;
  assign n25518 = ~pi1154 & ~n25517;
  assign n25519 = ~n25513 & n25518;
  assign n25520 = n17438 & ~n25453;
  assign n25521 = ~n25493 & ~n25520;
  assign n25522 = ~pi785 & ~n25521;
  assign n25523 = ~n25496 & ~n25506;
  assign n25524 = pi785 & ~n25523;
  assign n25525 = ~n25522 & ~n25524;
  assign n25526 = pi618 & n25525;
  assign n25527 = ~pi618 & n25453;
  assign n25528 = pi1154 & ~n25527;
  assign n25529 = ~n25526 & n25528;
  assign n25530 = ~pi627 & ~n25529;
  assign n25531 = ~n25519 & n25530;
  assign n25532 = pi618 & ~n25512;
  assign n25533 = ~pi618 & n25516;
  assign n25534 = pi1154 & ~n25533;
  assign n25535 = ~n25532 & n25534;
  assign n25536 = ~pi618 & n25525;
  assign n25537 = pi618 & n25453;
  assign n25538 = ~pi1154 & ~n25537;
  assign n25539 = ~n25536 & n25538;
  assign n25540 = pi627 & ~n25539;
  assign n25541 = ~n25535 & n25540;
  assign n25542 = ~n25531 & ~n25541;
  assign n25543 = pi781 & ~n25542;
  assign n25544 = ~pi781 & ~n25512;
  assign n25545 = ~n25543 & ~n25544;
  assign n25546 = ~pi619 & ~n25545;
  assign n25547 = ~n17503 & n25516;
  assign n25548 = n17503 & n25453;
  assign n25549 = ~n25547 & ~n25548;
  assign n25550 = pi619 & ~n25549;
  assign n25551 = ~pi1159 & ~n25550;
  assign n25552 = ~n25546 & n25551;
  assign n25553 = ~pi781 & ~n25525;
  assign n25554 = ~n25529 & ~n25539;
  assign n25555 = pi781 & ~n25554;
  assign n25556 = ~n25553 & ~n25555;
  assign n25557 = pi619 & n25556;
  assign n25558 = ~pi619 & n25453;
  assign n25559 = pi1159 & ~n25558;
  assign n25560 = ~n25557 & n25559;
  assign n25561 = ~pi648 & ~n25560;
  assign n25562 = ~n25552 & n25561;
  assign n25563 = pi619 & ~n25545;
  assign n25564 = ~pi619 & ~n25549;
  assign n25565 = pi1159 & ~n25564;
  assign n25566 = ~n25563 & n25565;
  assign n25567 = ~pi619 & n25556;
  assign n25568 = pi619 & n25453;
  assign n25569 = ~pi1159 & ~n25568;
  assign n25570 = ~n25567 & n25569;
  assign n25571 = pi648 & ~n25570;
  assign n25572 = ~n25566 & n25571;
  assign n25573 = ~n25562 & ~n25572;
  assign n25574 = pi789 & ~n25573;
  assign n25575 = ~pi789 & ~n25545;
  assign n25576 = ~n25574 & ~n25575;
  assign n25577 = ~pi788 & n25576;
  assign n25578 = ~pi626 & n25576;
  assign n25579 = n17539 & ~n25453;
  assign n25580 = ~n17539 & n25549;
  assign n25581 = ~n25579 & ~n25580;
  assign n25582 = pi626 & ~n25581;
  assign n25583 = ~pi641 & ~n25582;
  assign n25584 = ~n25578 & n25583;
  assign n25585 = ~pi789 & ~n25556;
  assign n25586 = ~n25560 & ~n25570;
  assign n25587 = pi789 & ~n25586;
  assign n25588 = ~n25585 & ~n25587;
  assign n25589 = ~pi626 & ~n25588;
  assign n25590 = pi626 & ~n25453;
  assign n25591 = pi641 & ~n25590;
  assign n25592 = ~n25589 & n25591;
  assign n25593 = ~pi1158 & ~n25592;
  assign n25594 = ~n25584 & n25593;
  assign n25595 = pi626 & n25576;
  assign n25596 = ~pi626 & ~n25581;
  assign n25597 = pi641 & ~n25596;
  assign n25598 = ~n25595 & n25597;
  assign n25599 = pi626 & ~n25588;
  assign n25600 = ~pi626 & ~n25453;
  assign n25601 = ~pi641 & ~n25600;
  assign n25602 = ~n25599 & n25601;
  assign n25603 = pi1158 & ~n25602;
  assign n25604 = ~n25598 & n25603;
  assign n25605 = ~n25594 & ~n25604;
  assign n25606 = pi788 & ~n25605;
  assign n25607 = ~n25577 & ~n25606;
  assign n25608 = ~pi628 & n25607;
  assign n25609 = ~n17816 & n25588;
  assign n25610 = n17816 & n25453;
  assign n25611 = ~n25609 & ~n25610;
  assign n25612 = pi628 & ~n25611;
  assign n25613 = ~pi1156 & ~n25612;
  assign n25614 = ~n25608 & n25613;
  assign n25615 = ~n17582 & n25581;
  assign n25616 = n17582 & n25453;
  assign n25617 = ~n25615 & ~n25616;
  assign n25618 = pi628 & ~n25617;
  assign n25619 = ~pi628 & n25453;
  assign n25620 = pi1156 & ~n25619;
  assign n25621 = ~n25618 & n25620;
  assign n25622 = ~pi629 & ~n25621;
  assign n25623 = ~n25614 & n25622;
  assign n25624 = pi628 & n25607;
  assign n25625 = ~pi628 & ~n25611;
  assign n25626 = pi1156 & ~n25625;
  assign n25627 = ~n25624 & n25626;
  assign n25628 = ~pi628 & ~n25617;
  assign n25629 = pi628 & n25453;
  assign n25630 = ~pi1156 & ~n25629;
  assign n25631 = ~n25628 & n25630;
  assign n25632 = pi629 & ~n25631;
  assign n25633 = ~n25627 & n25632;
  assign n25634 = ~n25623 & ~n25633;
  assign n25635 = pi792 & ~n25634;
  assign n25636 = ~pi792 & n25607;
  assign n25637 = ~n25635 & ~n25636;
  assign n25638 = ~pi647 & ~n25637;
  assign n25639 = ~n17610 & ~n25611;
  assign n25640 = n17610 & n25453;
  assign n25641 = ~n25639 & ~n25640;
  assign n25642 = pi647 & ~n25641;
  assign n25643 = ~pi1157 & ~n25642;
  assign n25644 = ~n25638 & n25643;
  assign n25645 = ~pi792 & n25617;
  assign n25646 = ~n25621 & ~n25631;
  assign n25647 = pi792 & ~n25646;
  assign n25648 = ~n25645 & ~n25647;
  assign n25649 = pi647 & n25648;
  assign n25650 = ~pi647 & n25453;
  assign n25651 = pi1157 & ~n25650;
  assign n25652 = ~n25649 & n25651;
  assign n25653 = ~pi630 & ~n25652;
  assign n25654 = ~n25644 & n25653;
  assign n25655 = pi647 & ~n25637;
  assign n25656 = ~pi647 & ~n25641;
  assign n25657 = pi1157 & ~n25656;
  assign n25658 = ~n25655 & n25657;
  assign n25659 = ~pi647 & n25648;
  assign n25660 = pi647 & n25453;
  assign n25661 = ~pi1157 & ~n25660;
  assign n25662 = ~n25659 & n25661;
  assign n25663 = pi630 & ~n25662;
  assign n25664 = ~n25658 & n25663;
  assign n25665 = ~n25654 & ~n25664;
  assign n25666 = pi787 & ~n25665;
  assign n25667 = ~pi787 & ~n25637;
  assign n25668 = ~n25666 & ~n25667;
  assign n25669 = ~pi644 & ~n25668;
  assign n25670 = ~pi787 & ~n25648;
  assign n25671 = ~n25652 & ~n25662;
  assign n25672 = pi787 & ~n25671;
  assign n25673 = ~n25670 & ~n25672;
  assign n25674 = pi644 & n25673;
  assign n25675 = ~pi715 & ~n25674;
  assign n25676 = ~n25669 & n25675;
  assign n25677 = n17652 & ~n25453;
  assign n25678 = ~n17652 & n25641;
  assign n25679 = ~n25677 & ~n25678;
  assign n25680 = ~pi644 & n25679;
  assign n25681 = pi644 & n25453;
  assign n25682 = pi715 & ~n25681;
  assign n25683 = ~n25680 & n25682;
  assign n25684 = ~pi1160 & ~n25683;
  assign n25685 = ~n25676 & n25684;
  assign n25686 = pi644 & ~n25668;
  assign n25687 = ~pi644 & n25673;
  assign n25688 = pi715 & ~n25687;
  assign n25689 = ~n25686 & n25688;
  assign n25690 = pi644 & n25679;
  assign n25691 = ~pi644 & n25453;
  assign n25692 = ~pi715 & ~n25691;
  assign n25693 = ~n25690 & n25692;
  assign n25694 = pi1160 & ~n25693;
  assign n25695 = ~n25689 & n25694;
  assign n25696 = pi790 & ~n25695;
  assign n25697 = ~n25685 & n25696;
  assign n25698 = ~pi790 & n25668;
  assign n25699 = ~po1038 & ~n25698;
  assign n25700 = ~n25697 & n25699;
  assign n25701 = ~pi179 & po1038;
  assign n25702 = ~pi832 & ~n25701;
  assign n25703 = ~n25700 & n25702;
  assign n25704 = ~pi179 & ~n2754;
  assign n25705 = ~pi741 & n16784;
  assign n25706 = ~n25704 & ~n25705;
  assign n25707 = ~n17706 & ~n25706;
  assign n25708 = ~pi785 & ~n25707;
  assign n25709 = ~n17711 & ~n25706;
  assign n25710 = pi1155 & ~n25709;
  assign n25711 = ~n17714 & n25707;
  assign n25712 = ~pi1155 & ~n25711;
  assign n25713 = ~n25710 & ~n25712;
  assign n25714 = pi785 & ~n25713;
  assign n25715 = ~n25708 & ~n25714;
  assign n25716 = ~pi781 & ~n25715;
  assign n25717 = ~n17721 & n25715;
  assign n25718 = pi1154 & ~n25717;
  assign n25719 = ~n17724 & n25715;
  assign n25720 = ~pi1154 & ~n25719;
  assign n25721 = ~n25718 & ~n25720;
  assign n25722 = pi781 & ~n25721;
  assign n25723 = ~n25716 & ~n25722;
  assign n25724 = ~pi789 & ~n25723;
  assign n25725 = pi619 & n25723;
  assign n25726 = ~pi619 & n25704;
  assign n25727 = pi1159 & ~n25726;
  assign n25728 = ~n25725 & n25727;
  assign n25729 = ~pi619 & n25723;
  assign n25730 = pi619 & n25704;
  assign n25731 = ~pi1159 & ~n25730;
  assign n25732 = ~n25729 & n25731;
  assign n25733 = ~n25728 & ~n25732;
  assign n25734 = pi789 & ~n25733;
  assign n25735 = ~n25724 & ~n25734;
  assign n25736 = ~n17816 & n25735;
  assign n25737 = n17816 & n25704;
  assign n25738 = ~n25736 & ~n25737;
  assign n25739 = ~n17610 & ~n25738;
  assign n25740 = n17610 & n25704;
  assign n25741 = ~n25739 & ~n25740;
  assign n25742 = ~n20398 & n25741;
  assign n25743 = ~pi724 & n16786;
  assign n25744 = ~n25704 & ~n25743;
  assign n25745 = ~pi778 & n25744;
  assign n25746 = ~pi625 & n25743;
  assign n25747 = ~n25744 & ~n25746;
  assign n25748 = pi1153 & ~n25747;
  assign n25749 = ~pi1153 & ~n25704;
  assign n25750 = ~n25746 & n25749;
  assign n25751 = ~n25748 & ~n25750;
  assign n25752 = pi778 & ~n25751;
  assign n25753 = ~n25745 & ~n25752;
  assign n25754 = ~n17692 & n25753;
  assign n25755 = ~n17694 & n25754;
  assign n25756 = ~n17696 & n25755;
  assign n25757 = ~n17828 & n25756;
  assign n25758 = ~n17859 & n25757;
  assign n25759 = ~pi647 & n25758;
  assign n25760 = pi647 & n25704;
  assign n25761 = ~pi1157 & ~n25760;
  assign n25762 = ~n25759 & n25761;
  assign n25763 = pi647 & ~n25758;
  assign n25764 = ~pi647 & ~n25704;
  assign n25765 = ~n25763 & ~n25764;
  assign n25766 = pi1157 & ~n25765;
  assign n25767 = ~n25762 & ~n25766;
  assign n25768 = ~n17651 & ~n25767;
  assign n25769 = ~n25742 & ~n25768;
  assign n25770 = pi787 & ~n25769;
  assign n25771 = pi626 & ~n25735;
  assign n25772 = ~pi626 & ~n25704;
  assign n25773 = n17579 & ~n25772;
  assign n25774 = ~n25771 & n25773;
  assign n25775 = n17704 & n25756;
  assign n25776 = ~pi626 & ~n25735;
  assign n25777 = pi626 & ~n25704;
  assign n25778 = n17580 & ~n25777;
  assign n25779 = ~n25776 & n25778;
  assign n25780 = ~n25775 & ~n25779;
  assign n25781 = ~n25774 & n25780;
  assign n25782 = pi788 & ~n25781;
  assign n25783 = ~n16521 & ~n25744;
  assign n25784 = pi625 & n25783;
  assign n25785 = n25706 & ~n25783;
  assign n25786 = ~n25784 & ~n25785;
  assign n25787 = n25749 & ~n25786;
  assign n25788 = ~pi608 & ~n25748;
  assign n25789 = ~n25787 & n25788;
  assign n25790 = pi1153 & n25706;
  assign n25791 = ~n25784 & n25790;
  assign n25792 = pi608 & ~n25750;
  assign n25793 = ~n25791 & n25792;
  assign n25794 = ~n25789 & ~n25793;
  assign n25795 = pi778 & ~n25794;
  assign n25796 = ~pi778 & ~n25785;
  assign n25797 = ~n25795 & ~n25796;
  assign n25798 = ~pi609 & ~n25797;
  assign n25799 = pi609 & n25753;
  assign n25800 = ~pi1155 & ~n25799;
  assign n25801 = ~n25798 & n25800;
  assign n25802 = ~pi660 & ~n25710;
  assign n25803 = ~n25801 & n25802;
  assign n25804 = pi609 & ~n25797;
  assign n25805 = ~pi609 & n25753;
  assign n25806 = pi1155 & ~n25805;
  assign n25807 = ~n25804 & n25806;
  assign n25808 = pi660 & ~n25712;
  assign n25809 = ~n25807 & n25808;
  assign n25810 = ~n25803 & ~n25809;
  assign n25811 = pi785 & ~n25810;
  assign n25812 = ~pi785 & ~n25797;
  assign n25813 = ~n25811 & ~n25812;
  assign n25814 = ~pi618 & ~n25813;
  assign n25815 = pi618 & n25754;
  assign n25816 = ~pi1154 & ~n25815;
  assign n25817 = ~n25814 & n25816;
  assign n25818 = ~pi627 & ~n25718;
  assign n25819 = ~n25817 & n25818;
  assign n25820 = pi618 & ~n25813;
  assign n25821 = ~pi618 & n25754;
  assign n25822 = pi1154 & ~n25821;
  assign n25823 = ~n25820 & n25822;
  assign n25824 = pi627 & ~n25720;
  assign n25825 = ~n25823 & n25824;
  assign n25826 = ~n25819 & ~n25825;
  assign n25827 = pi781 & ~n25826;
  assign n25828 = ~pi781 & ~n25813;
  assign n25829 = ~n25827 & ~n25828;
  assign n25830 = pi619 & ~n25829;
  assign n25831 = ~pi619 & n25755;
  assign n25832 = pi1159 & ~n25831;
  assign n25833 = ~n25830 & n25832;
  assign n25834 = pi648 & ~n25732;
  assign n25835 = ~n25833 & n25834;
  assign n25836 = ~pi619 & ~n25829;
  assign n25837 = pi619 & n25755;
  assign n25838 = ~pi1159 & ~n25837;
  assign n25839 = ~n25836 & n25838;
  assign n25840 = ~pi648 & ~n25728;
  assign n25841 = ~n25839 & n25840;
  assign n25842 = pi789 & ~n25841;
  assign n25843 = ~n25835 & n25842;
  assign n25844 = ~pi789 & n25829;
  assign n25845 = n17817 & ~n25844;
  assign n25846 = ~n25843 & n25845;
  assign n25847 = ~n25782 & ~n25846;
  assign n25848 = ~n20205 & ~n25847;
  assign n25849 = n17856 & ~n25738;
  assign n25850 = n20693 & n25757;
  assign n25851 = ~n25849 & ~n25850;
  assign n25852 = ~pi629 & ~n25851;
  assign n25853 = n20697 & n25757;
  assign n25854 = n17855 & ~n25738;
  assign n25855 = ~n25853 & ~n25854;
  assign n25856 = pi629 & ~n25855;
  assign n25857 = ~n25852 & ~n25856;
  assign n25858 = pi792 & ~n25857;
  assign n25859 = n20207 & ~n25858;
  assign n25860 = ~n25848 & n25859;
  assign n25861 = ~n25770 & ~n25860;
  assign n25862 = pi644 & n25861;
  assign n25863 = ~pi787 & ~n25758;
  assign n25864 = pi787 & ~n25767;
  assign n25865 = ~n25863 & ~n25864;
  assign n25866 = ~pi644 & n25865;
  assign n25867 = pi715 & ~n25866;
  assign n25868 = ~n25862 & n25867;
  assign n25869 = ~n17652 & ~n25741;
  assign n25870 = n17652 & n25704;
  assign n25871 = ~n25869 & ~n25870;
  assign n25872 = pi644 & ~n25871;
  assign n25873 = ~pi644 & n25704;
  assign n25874 = ~pi715 & ~n25873;
  assign n25875 = ~n25872 & n25874;
  assign n25876 = pi1160 & ~n25875;
  assign n25877 = ~n25868 & n25876;
  assign n25878 = ~pi644 & n25861;
  assign n25879 = pi644 & n25865;
  assign n25880 = ~pi715 & ~n25879;
  assign n25881 = ~n25878 & n25880;
  assign n25882 = ~pi644 & ~n25871;
  assign n25883 = pi644 & n25704;
  assign n25884 = pi715 & ~n25883;
  assign n25885 = ~n25882 & n25884;
  assign n25886 = ~pi1160 & ~n25885;
  assign n25887 = ~n25881 & n25886;
  assign n25888 = ~n25877 & ~n25887;
  assign n25889 = pi790 & ~n25888;
  assign n25890 = ~pi790 & n25861;
  assign n25891 = pi832 & ~n25890;
  assign n25892 = ~n25889 & n25891;
  assign po336 = ~n25703 & ~n25892;
  assign n25894 = ~pi180 & ~n2754;
  assign n25895 = ~pi753 & n16784;
  assign n25896 = ~n25894 & ~n25895;
  assign n25897 = ~n17706 & ~n25896;
  assign n25898 = ~pi785 & ~n25897;
  assign n25899 = n17451 & n25895;
  assign n25900 = n25897 & ~n25899;
  assign n25901 = pi1155 & ~n25900;
  assign n25902 = ~pi1155 & ~n25894;
  assign n25903 = ~n25899 & n25902;
  assign n25904 = ~n25901 & ~n25903;
  assign n25905 = pi785 & ~n25904;
  assign n25906 = ~n25898 & ~n25905;
  assign n25907 = ~pi781 & ~n25906;
  assign n25908 = ~n17721 & n25906;
  assign n25909 = pi1154 & ~n25908;
  assign n25910 = ~n17724 & n25906;
  assign n25911 = ~pi1154 & ~n25910;
  assign n25912 = ~n25909 & ~n25911;
  assign n25913 = pi781 & ~n25912;
  assign n25914 = ~n25907 & ~n25913;
  assign n25915 = ~pi789 & ~n25914;
  assign n25916 = ~n22890 & n25914;
  assign n25917 = pi1159 & ~n25916;
  assign n25918 = ~n22893 & n25914;
  assign n25919 = ~pi1159 & ~n25918;
  assign n25920 = ~n25917 & ~n25919;
  assign n25921 = pi789 & ~n25920;
  assign n25922 = ~n25915 & ~n25921;
  assign n25923 = ~n17816 & n25922;
  assign n25924 = n17816 & n25894;
  assign n25925 = ~n25923 & ~n25924;
  assign n25926 = ~n17610 & ~n25925;
  assign n25927 = n17610 & n25894;
  assign n25928 = ~n25926 & ~n25927;
  assign n25929 = ~n20398 & n25928;
  assign n25930 = ~pi702 & n16786;
  assign n25931 = ~n25894 & ~n25930;
  assign n25932 = ~pi778 & ~n25931;
  assign n25933 = ~pi625 & n25930;
  assign n25934 = ~n25931 & ~n25933;
  assign n25935 = pi1153 & ~n25934;
  assign n25936 = ~pi1153 & ~n25894;
  assign n25937 = ~n25933 & n25936;
  assign n25938 = pi778 & ~n25937;
  assign n25939 = ~n25935 & n25938;
  assign n25940 = ~n25932 & ~n25939;
  assign n25941 = ~n17692 & ~n25940;
  assign n25942 = ~n17694 & n25941;
  assign n25943 = ~n17696 & n25942;
  assign n25944 = ~n17828 & n25943;
  assign n25945 = ~n17859 & n25944;
  assign n25946 = ~pi647 & n25945;
  assign n25947 = pi647 & n25894;
  assign n25948 = ~pi1157 & ~n25947;
  assign n25949 = ~n25946 & n25948;
  assign n25950 = pi647 & ~n25945;
  assign n25951 = ~pi647 & ~n25894;
  assign n25952 = ~n25950 & ~n25951;
  assign n25953 = pi1157 & ~n25952;
  assign n25954 = ~n25949 & ~n25953;
  assign n25955 = ~n17651 & ~n25954;
  assign n25956 = ~n25929 & ~n25955;
  assign n25957 = pi787 & ~n25956;
  assign n25958 = pi626 & ~n25922;
  assign n25959 = ~pi626 & ~n25894;
  assign n25960 = n17579 & ~n25959;
  assign n25961 = ~n25958 & n25960;
  assign n25962 = n17704 & n25943;
  assign n25963 = ~pi626 & ~n25922;
  assign n25964 = pi626 & ~n25894;
  assign n25965 = n17580 & ~n25964;
  assign n25966 = ~n25963 & n25965;
  assign n25967 = ~n25962 & ~n25966;
  assign n25968 = ~n25961 & n25967;
  assign n25969 = pi788 & ~n25968;
  assign n25970 = ~n16521 & ~n25931;
  assign n25971 = pi625 & n25970;
  assign n25972 = n25896 & ~n25970;
  assign n25973 = ~n25971 & ~n25972;
  assign n25974 = n25936 & ~n25973;
  assign n25975 = ~pi608 & ~n25935;
  assign n25976 = ~n25974 & n25975;
  assign n25977 = pi1153 & n25896;
  assign n25978 = ~n25971 & n25977;
  assign n25979 = pi608 & ~n25937;
  assign n25980 = ~n25978 & n25979;
  assign n25981 = ~n25976 & ~n25980;
  assign n25982 = pi778 & ~n25981;
  assign n25983 = ~pi778 & ~n25972;
  assign n25984 = ~n25982 & ~n25983;
  assign n25985 = ~pi609 & ~n25984;
  assign n25986 = pi609 & ~n25940;
  assign n25987 = ~pi1155 & ~n25986;
  assign n25988 = ~n25985 & n25987;
  assign n25989 = ~pi660 & ~n25901;
  assign n25990 = ~n25988 & n25989;
  assign n25991 = pi609 & ~n25984;
  assign n25992 = ~pi609 & ~n25940;
  assign n25993 = pi1155 & ~n25992;
  assign n25994 = ~n25991 & n25993;
  assign n25995 = pi660 & ~n25903;
  assign n25996 = ~n25994 & n25995;
  assign n25997 = ~n25990 & ~n25996;
  assign n25998 = pi785 & ~n25997;
  assign n25999 = ~pi785 & ~n25984;
  assign n26000 = ~n25998 & ~n25999;
  assign n26001 = ~pi618 & ~n26000;
  assign n26002 = pi618 & n25941;
  assign n26003 = ~pi1154 & ~n26002;
  assign n26004 = ~n26001 & n26003;
  assign n26005 = ~pi627 & ~n25909;
  assign n26006 = ~n26004 & n26005;
  assign n26007 = pi618 & ~n26000;
  assign n26008 = ~pi618 & n25941;
  assign n26009 = pi1154 & ~n26008;
  assign n26010 = ~n26007 & n26009;
  assign n26011 = pi627 & ~n25911;
  assign n26012 = ~n26010 & n26011;
  assign n26013 = ~n26006 & ~n26012;
  assign n26014 = pi781 & ~n26013;
  assign n26015 = ~pi781 & ~n26000;
  assign n26016 = ~n26014 & ~n26015;
  assign n26017 = pi619 & ~n26016;
  assign n26018 = ~pi619 & n25942;
  assign n26019 = pi1159 & ~n26018;
  assign n26020 = ~n26017 & n26019;
  assign n26021 = pi648 & ~n25919;
  assign n26022 = ~n26020 & n26021;
  assign n26023 = ~pi619 & ~n26016;
  assign n26024 = pi619 & n25942;
  assign n26025 = ~pi1159 & ~n26024;
  assign n26026 = ~n26023 & n26025;
  assign n26027 = ~pi648 & ~n25917;
  assign n26028 = ~n26026 & n26027;
  assign n26029 = pi789 & ~n26028;
  assign n26030 = ~n26022 & n26029;
  assign n26031 = ~pi789 & n26016;
  assign n26032 = n17817 & ~n26031;
  assign n26033 = ~n26030 & n26032;
  assign n26034 = ~n25969 & ~n26033;
  assign n26035 = ~n20205 & ~n26034;
  assign n26036 = n17856 & ~n25925;
  assign n26037 = n20693 & n25944;
  assign n26038 = ~n26036 & ~n26037;
  assign n26039 = ~pi629 & ~n26038;
  assign n26040 = n20697 & n25944;
  assign n26041 = n17855 & ~n25925;
  assign n26042 = ~n26040 & ~n26041;
  assign n26043 = pi629 & ~n26042;
  assign n26044 = ~n26039 & ~n26043;
  assign n26045 = pi792 & ~n26044;
  assign n26046 = n20207 & ~n26045;
  assign n26047 = ~n26035 & n26046;
  assign n26048 = ~n25957 & ~n26047;
  assign n26049 = pi644 & n26048;
  assign n26050 = ~pi787 & ~n25945;
  assign n26051 = pi787 & ~n25954;
  assign n26052 = ~n26050 & ~n26051;
  assign n26053 = ~pi644 & n26052;
  assign n26054 = pi715 & ~n26053;
  assign n26055 = ~n26049 & n26054;
  assign n26056 = ~n17652 & ~n25928;
  assign n26057 = n17652 & n25894;
  assign n26058 = ~n26056 & ~n26057;
  assign n26059 = pi644 & ~n26058;
  assign n26060 = ~pi644 & n25894;
  assign n26061 = ~pi715 & ~n26060;
  assign n26062 = ~n26059 & n26061;
  assign n26063 = pi1160 & ~n26062;
  assign n26064 = ~n26055 & n26063;
  assign n26065 = ~pi644 & n26048;
  assign n26066 = pi644 & n26052;
  assign n26067 = ~pi715 & ~n26066;
  assign n26068 = ~n26065 & n26067;
  assign n26069 = ~pi644 & ~n26058;
  assign n26070 = pi644 & n25894;
  assign n26071 = pi715 & ~n26070;
  assign n26072 = ~n26069 & n26071;
  assign n26073 = ~pi1160 & ~n26072;
  assign n26074 = ~n26068 & n26073;
  assign n26075 = ~n26064 & ~n26074;
  assign n26076 = pi790 & ~n26075;
  assign n26077 = ~pi790 & n26048;
  assign n26078 = pi832 & ~n26077;
  assign n26079 = ~n26076 & n26078;
  assign n26080 = ~pi180 & ~n17406;
  assign n26081 = n17539 & ~n26080;
  assign n26082 = ~pi702 & n3267;
  assign n26083 = n26080 & ~n26082;
  assign n26084 = pi180 & ~n17976;
  assign n26085 = ~pi38 & ~n26084;
  assign n26086 = n3267 & ~n26085;
  assign n26087 = ~pi180 & n17972;
  assign n26088 = ~n26086 & ~n26087;
  assign n26089 = ~pi180 & ~n17280;
  assign n26090 = n17392 & ~n26089;
  assign n26091 = ~pi702 & ~n26090;
  assign n26092 = ~n26088 & n26091;
  assign n26093 = ~n26083 & ~n26092;
  assign n26094 = ~pi778 & n26093;
  assign n26095 = pi625 & ~n26093;
  assign n26096 = ~pi625 & n26080;
  assign n26097 = pi1153 & ~n26096;
  assign n26098 = ~n26095 & n26097;
  assign n26099 = ~pi625 & ~n26093;
  assign n26100 = pi625 & n26080;
  assign n26101 = ~pi1153 & ~n26100;
  assign n26102 = ~n26099 & n26101;
  assign n26103 = ~n26098 & ~n26102;
  assign n26104 = pi778 & ~n26103;
  assign n26105 = ~n26094 & ~n26104;
  assign n26106 = ~n17466 & ~n26105;
  assign n26107 = n17466 & ~n26080;
  assign n26108 = ~n26106 & ~n26107;
  assign n26109 = ~n17503 & n26108;
  assign n26110 = n17503 & n26080;
  assign n26111 = ~n26109 & ~n26110;
  assign n26112 = ~n17539 & n26111;
  assign n26113 = ~n26081 & ~n26112;
  assign n26114 = ~n17582 & n26113;
  assign n26115 = n17582 & n26080;
  assign n26116 = ~n26114 & ~n26115;
  assign n26117 = ~pi792 & n26116;
  assign n26118 = pi628 & ~n26116;
  assign n26119 = ~pi628 & n26080;
  assign n26120 = pi1156 & ~n26119;
  assign n26121 = ~n26118 & n26120;
  assign n26122 = ~pi628 & ~n26116;
  assign n26123 = pi628 & n26080;
  assign n26124 = ~pi1156 & ~n26123;
  assign n26125 = ~n26122 & n26124;
  assign n26126 = ~n26121 & ~n26125;
  assign n26127 = pi792 & ~n26126;
  assign n26128 = ~n26117 & ~n26127;
  assign n26129 = ~pi647 & ~n26128;
  assign n26130 = pi647 & ~n26080;
  assign n26131 = ~n26129 & ~n26130;
  assign n26132 = ~pi1157 & n26131;
  assign n26133 = pi647 & ~n26128;
  assign n26134 = ~pi647 & ~n26080;
  assign n26135 = ~n26133 & ~n26134;
  assign n26136 = pi1157 & n26135;
  assign n26137 = ~n26132 & ~n26136;
  assign n26138 = pi787 & ~n26137;
  assign n26139 = ~pi787 & n26128;
  assign n26140 = ~n26138 & ~n26139;
  assign n26141 = ~pi644 & ~n26140;
  assign n26142 = pi715 & ~n26141;
  assign n26143 = pi180 & ~n3267;
  assign n26144 = pi753 & n17199;
  assign n26145 = pi180 & n17273;
  assign n26146 = ~n26144 & ~n26145;
  assign n26147 = pi39 & ~n26146;
  assign n26148 = ~pi180 & ~pi753;
  assign n26149 = n17242 & n26148;
  assign n26150 = pi180 & pi753;
  assign n26151 = pi180 & ~n17086;
  assign n26152 = ~n21592 & ~n26151;
  assign n26153 = ~pi39 & ~n26152;
  assign n26154 = ~n26150 & ~n26153;
  assign n26155 = ~n26149 & n26154;
  assign n26156 = ~n26147 & n26155;
  assign n26157 = ~pi38 & ~n26156;
  assign n26158 = ~pi753 & n17282;
  assign n26159 = pi38 & ~n26089;
  assign n26160 = ~n26158 & n26159;
  assign n26161 = ~n26157 & ~n26160;
  assign n26162 = n3267 & ~n26161;
  assign n26163 = ~n26143 & ~n26162;
  assign n26164 = ~n17438 & ~n26163;
  assign n26165 = n17438 & ~n26080;
  assign n26166 = ~n26164 & ~n26165;
  assign n26167 = ~pi785 & ~n26166;
  assign n26168 = ~n17439 & ~n26080;
  assign n26169 = pi609 & n26164;
  assign n26170 = ~n26168 & ~n26169;
  assign n26171 = pi1155 & ~n26170;
  assign n26172 = ~n17451 & ~n26080;
  assign n26173 = ~pi609 & n26164;
  assign n26174 = ~n26172 & ~n26173;
  assign n26175 = ~pi1155 & ~n26174;
  assign n26176 = ~n26171 & ~n26175;
  assign n26177 = pi785 & ~n26176;
  assign n26178 = ~n26167 & ~n26177;
  assign n26179 = ~pi781 & ~n26178;
  assign n26180 = pi618 & n26178;
  assign n26181 = ~pi618 & n26080;
  assign n26182 = pi1154 & ~n26181;
  assign n26183 = ~n26180 & n26182;
  assign n26184 = ~pi618 & n26178;
  assign n26185 = pi618 & n26080;
  assign n26186 = ~pi1154 & ~n26185;
  assign n26187 = ~n26184 & n26186;
  assign n26188 = ~n26183 & ~n26187;
  assign n26189 = pi781 & ~n26188;
  assign n26190 = ~n26179 & ~n26189;
  assign n26191 = ~pi789 & ~n26190;
  assign n26192 = pi619 & n26190;
  assign n26193 = ~pi619 & n26080;
  assign n26194 = pi1159 & ~n26193;
  assign n26195 = ~n26192 & n26194;
  assign n26196 = ~pi619 & n26190;
  assign n26197 = pi619 & n26080;
  assign n26198 = ~pi1159 & ~n26197;
  assign n26199 = ~n26196 & n26198;
  assign n26200 = ~n26195 & ~n26199;
  assign n26201 = pi789 & ~n26200;
  assign n26202 = ~n26191 & ~n26201;
  assign n26203 = ~n17816 & n26202;
  assign n26204 = n17816 & n26080;
  assign n26205 = ~n26203 & ~n26204;
  assign n26206 = ~n17610 & ~n26205;
  assign n26207 = n17610 & n26080;
  assign n26208 = ~n26206 & ~n26207;
  assign n26209 = ~n17652 & ~n26208;
  assign n26210 = n17652 & n26080;
  assign n26211 = ~n26209 & ~n26210;
  assign n26212 = pi644 & ~n26211;
  assign n26213 = ~pi644 & n26080;
  assign n26214 = ~pi715 & ~n26213;
  assign n26215 = ~n26212 & n26214;
  assign n26216 = pi1160 & ~n26215;
  assign n26217 = ~n26142 & n26216;
  assign n26218 = pi644 & ~n26140;
  assign n26219 = ~pi715 & ~n26218;
  assign n26220 = ~pi644 & ~n26211;
  assign n26221 = pi644 & n26080;
  assign n26222 = pi715 & ~n26221;
  assign n26223 = ~n26220 & n26222;
  assign n26224 = ~pi1160 & ~n26223;
  assign n26225 = ~n26219 & n26224;
  assign n26226 = ~n26217 & ~n26225;
  assign n26227 = pi790 & ~n26226;
  assign n26228 = pi644 & n26216;
  assign n26229 = ~pi644 & n26224;
  assign n26230 = pi790 & ~n26229;
  assign n26231 = ~n26228 & n26230;
  assign n26232 = ~n20409 & n26205;
  assign n26233 = ~pi629 & n26121;
  assign n26234 = pi629 & n26125;
  assign n26235 = ~n26233 & ~n26234;
  assign n26236 = ~n26232 & n26235;
  assign n26237 = pi792 & ~n26236;
  assign n26238 = pi702 & n26161;
  assign n26239 = ~pi180 & n16687;
  assign n26240 = pi180 & n16799;
  assign n26241 = pi753 & ~n26240;
  assign n26242 = ~n26239 & n26241;
  assign n26243 = pi180 & n16879;
  assign n26244 = ~pi180 & ~n16944;
  assign n26245 = ~pi753 & ~n26244;
  assign n26246 = ~n26243 & n26245;
  assign n26247 = pi39 & ~n26246;
  assign n26248 = ~n26242 & n26247;
  assign n26249 = ~pi180 & ~n17088;
  assign n26250 = pi180 & ~n17059;
  assign n26251 = pi753 & ~n26250;
  assign n26252 = ~n26249 & n26251;
  assign n26253 = ~pi180 & n17092;
  assign n26254 = pi180 & n17094;
  assign n26255 = ~pi753 & ~n26254;
  assign n26256 = ~n26253 & n26255;
  assign n26257 = ~n26252 & ~n26256;
  assign n26258 = ~pi39 & ~n26257;
  assign n26259 = ~pi38 & ~n26258;
  assign n26260 = ~n26248 & n26259;
  assign n26261 = ~pi753 & ~n16905;
  assign n26262 = n19230 & ~n26261;
  assign n26263 = ~pi180 & ~n26262;
  assign n26264 = ~n16787 & ~n25895;
  assign n26265 = pi180 & ~n26264;
  assign n26266 = n6234 & n26265;
  assign n26267 = pi38 & ~n26266;
  assign n26268 = ~n26263 & n26267;
  assign n26269 = ~pi702 & ~n26268;
  assign n26270 = ~n26260 & n26269;
  assign n26271 = n3267 & ~n26270;
  assign n26272 = ~n26238 & n26271;
  assign n26273 = ~n26143 & ~n26272;
  assign n26274 = ~pi625 & n26273;
  assign n26275 = pi625 & n26163;
  assign n26276 = ~pi1153 & ~n26275;
  assign n26277 = ~n26274 & n26276;
  assign n26278 = ~pi608 & ~n26098;
  assign n26279 = ~n26277 & n26278;
  assign n26280 = pi625 & n26273;
  assign n26281 = ~pi625 & n26163;
  assign n26282 = pi1153 & ~n26281;
  assign n26283 = ~n26280 & n26282;
  assign n26284 = pi608 & ~n26102;
  assign n26285 = ~n26283 & n26284;
  assign n26286 = ~n26279 & ~n26285;
  assign n26287 = pi778 & ~n26286;
  assign n26288 = ~pi778 & n26273;
  assign n26289 = ~n26287 & ~n26288;
  assign n26290 = ~pi609 & ~n26289;
  assign n26291 = pi609 & n26105;
  assign n26292 = ~pi1155 & ~n26291;
  assign n26293 = ~n26290 & n26292;
  assign n26294 = ~pi660 & ~n26171;
  assign n26295 = ~n26293 & n26294;
  assign n26296 = pi609 & ~n26289;
  assign n26297 = ~pi609 & n26105;
  assign n26298 = pi1155 & ~n26297;
  assign n26299 = ~n26296 & n26298;
  assign n26300 = pi660 & ~n26175;
  assign n26301 = ~n26299 & n26300;
  assign n26302 = ~n26295 & ~n26301;
  assign n26303 = pi785 & ~n26302;
  assign n26304 = ~pi785 & ~n26289;
  assign n26305 = ~n26303 & ~n26304;
  assign n26306 = ~pi618 & ~n26305;
  assign n26307 = pi618 & n26108;
  assign n26308 = ~pi1154 & ~n26307;
  assign n26309 = ~n26306 & n26308;
  assign n26310 = ~pi627 & ~n26183;
  assign n26311 = ~n26309 & n26310;
  assign n26312 = pi618 & ~n26305;
  assign n26313 = ~pi618 & n26108;
  assign n26314 = pi1154 & ~n26313;
  assign n26315 = ~n26312 & n26314;
  assign n26316 = pi627 & ~n26187;
  assign n26317 = ~n26315 & n26316;
  assign n26318 = ~n26311 & ~n26317;
  assign n26319 = pi781 & ~n26318;
  assign n26320 = ~pi781 & ~n26305;
  assign n26321 = ~n26319 & ~n26320;
  assign n26322 = pi619 & ~n26321;
  assign n26323 = ~pi619 & ~n26111;
  assign n26324 = pi1159 & ~n26323;
  assign n26325 = ~n26322 & n26324;
  assign n26326 = pi648 & ~n26199;
  assign n26327 = ~n26325 & n26326;
  assign n26328 = ~pi619 & ~n26321;
  assign n26329 = pi619 & ~n26111;
  assign n26330 = ~pi1159 & ~n26329;
  assign n26331 = ~n26328 & n26330;
  assign n26332 = ~pi648 & ~n26195;
  assign n26333 = ~n26331 & n26332;
  assign n26334 = pi789 & ~n26333;
  assign n26335 = ~n26327 & n26334;
  assign n26336 = ~pi789 & n26321;
  assign n26337 = n17817 & ~n26336;
  assign n26338 = ~n26335 & n26337;
  assign n26339 = pi626 & ~n26202;
  assign n26340 = ~pi626 & ~n26080;
  assign n26341 = n17579 & ~n26340;
  assign n26342 = ~n26339 & n26341;
  assign n26343 = n17704 & n26113;
  assign n26344 = ~pi626 & ~n26202;
  assign n26345 = pi626 & ~n26080;
  assign n26346 = n17580 & ~n26345;
  assign n26347 = ~n26344 & n26346;
  assign n26348 = ~n26343 & ~n26347;
  assign n26349 = ~n26342 & n26348;
  assign n26350 = pi788 & ~n26349;
  assign n26351 = ~n20205 & ~n26350;
  assign n26352 = ~n26338 & n26351;
  assign n26353 = ~n26237 & ~n26352;
  assign n26354 = n20207 & ~n26353;
  assign n26355 = ~n20398 & n26208;
  assign n26356 = n17650 & ~n26131;
  assign n26357 = n17649 & ~n26135;
  assign n26358 = ~n26356 & ~n26357;
  assign n26359 = ~n26355 & n26358;
  assign n26360 = pi787 & ~n26359;
  assign n26361 = ~n26354 & ~n26360;
  assign n26362 = ~n26231 & n26361;
  assign n26363 = ~n26227 & ~n26362;
  assign n26364 = ~po1038 & ~n26363;
  assign n26365 = ~pi180 & po1038;
  assign n26366 = ~pi832 & ~n26365;
  assign n26367 = ~n26364 & n26366;
  assign po337 = ~n26079 & ~n26367;
  assign n26369 = ~pi181 & ~n2754;
  assign n26370 = ~pi754 & n16784;
  assign n26371 = ~n26369 & ~n26370;
  assign n26372 = ~n17706 & ~n26371;
  assign n26373 = ~pi785 & ~n26372;
  assign n26374 = n17451 & n26370;
  assign n26375 = n26372 & ~n26374;
  assign n26376 = pi1155 & ~n26375;
  assign n26377 = ~pi1155 & ~n26369;
  assign n26378 = ~n26374 & n26377;
  assign n26379 = ~n26376 & ~n26378;
  assign n26380 = pi785 & ~n26379;
  assign n26381 = ~n26373 & ~n26380;
  assign n26382 = ~pi781 & ~n26381;
  assign n26383 = ~n17721 & n26381;
  assign n26384 = pi1154 & ~n26383;
  assign n26385 = ~n17724 & n26381;
  assign n26386 = ~pi1154 & ~n26385;
  assign n26387 = ~n26384 & ~n26386;
  assign n26388 = pi781 & ~n26387;
  assign n26389 = ~n26382 & ~n26388;
  assign n26390 = ~pi789 & ~n26389;
  assign n26391 = ~n22890 & n26389;
  assign n26392 = pi1159 & ~n26391;
  assign n26393 = ~n22893 & n26389;
  assign n26394 = ~pi1159 & ~n26393;
  assign n26395 = ~n26392 & ~n26394;
  assign n26396 = pi789 & ~n26395;
  assign n26397 = ~n26390 & ~n26396;
  assign n26398 = ~n17816 & n26397;
  assign n26399 = n17816 & n26369;
  assign n26400 = ~n26398 & ~n26399;
  assign n26401 = ~n17610 & ~n26400;
  assign n26402 = n17610 & n26369;
  assign n26403 = ~n26401 & ~n26402;
  assign n26404 = ~n20398 & n26403;
  assign n26405 = ~pi709 & n16786;
  assign n26406 = ~n26369 & ~n26405;
  assign n26407 = ~pi778 & ~n26406;
  assign n26408 = ~pi625 & n26405;
  assign n26409 = ~n26406 & ~n26408;
  assign n26410 = pi1153 & ~n26409;
  assign n26411 = ~pi1153 & ~n26369;
  assign n26412 = ~n26408 & n26411;
  assign n26413 = pi778 & ~n26412;
  assign n26414 = ~n26410 & n26413;
  assign n26415 = ~n26407 & ~n26414;
  assign n26416 = ~n17692 & ~n26415;
  assign n26417 = ~n17694 & n26416;
  assign n26418 = ~n17696 & n26417;
  assign n26419 = ~n17828 & n26418;
  assign n26420 = ~n17859 & n26419;
  assign n26421 = ~pi647 & n26420;
  assign n26422 = pi647 & n26369;
  assign n26423 = ~pi1157 & ~n26422;
  assign n26424 = ~n26421 & n26423;
  assign n26425 = pi647 & ~n26420;
  assign n26426 = ~pi647 & ~n26369;
  assign n26427 = ~n26425 & ~n26426;
  assign n26428 = pi1157 & ~n26427;
  assign n26429 = ~n26424 & ~n26428;
  assign n26430 = ~n17651 & ~n26429;
  assign n26431 = ~n26404 & ~n26430;
  assign n26432 = pi787 & ~n26431;
  assign n26433 = pi626 & ~n26397;
  assign n26434 = ~pi626 & ~n26369;
  assign n26435 = n17579 & ~n26434;
  assign n26436 = ~n26433 & n26435;
  assign n26437 = n17704 & n26418;
  assign n26438 = ~pi626 & ~n26397;
  assign n26439 = pi626 & ~n26369;
  assign n26440 = n17580 & ~n26439;
  assign n26441 = ~n26438 & n26440;
  assign n26442 = ~n26437 & ~n26441;
  assign n26443 = ~n26436 & n26442;
  assign n26444 = pi788 & ~n26443;
  assign n26445 = ~n16521 & ~n26406;
  assign n26446 = pi625 & n26445;
  assign n26447 = n26371 & ~n26445;
  assign n26448 = ~n26446 & ~n26447;
  assign n26449 = n26411 & ~n26448;
  assign n26450 = ~pi608 & ~n26410;
  assign n26451 = ~n26449 & n26450;
  assign n26452 = pi1153 & n26371;
  assign n26453 = ~n26446 & n26452;
  assign n26454 = pi608 & ~n26412;
  assign n26455 = ~n26453 & n26454;
  assign n26456 = ~n26451 & ~n26455;
  assign n26457 = pi778 & ~n26456;
  assign n26458 = ~pi778 & ~n26447;
  assign n26459 = ~n26457 & ~n26458;
  assign n26460 = ~pi609 & ~n26459;
  assign n26461 = pi609 & ~n26415;
  assign n26462 = ~pi1155 & ~n26461;
  assign n26463 = ~n26460 & n26462;
  assign n26464 = ~pi660 & ~n26376;
  assign n26465 = ~n26463 & n26464;
  assign n26466 = pi609 & ~n26459;
  assign n26467 = ~pi609 & ~n26415;
  assign n26468 = pi1155 & ~n26467;
  assign n26469 = ~n26466 & n26468;
  assign n26470 = pi660 & ~n26378;
  assign n26471 = ~n26469 & n26470;
  assign n26472 = ~n26465 & ~n26471;
  assign n26473 = pi785 & ~n26472;
  assign n26474 = ~pi785 & ~n26459;
  assign n26475 = ~n26473 & ~n26474;
  assign n26476 = ~pi618 & ~n26475;
  assign n26477 = pi618 & n26416;
  assign n26478 = ~pi1154 & ~n26477;
  assign n26479 = ~n26476 & n26478;
  assign n26480 = ~pi627 & ~n26384;
  assign n26481 = ~n26479 & n26480;
  assign n26482 = pi618 & ~n26475;
  assign n26483 = ~pi618 & n26416;
  assign n26484 = pi1154 & ~n26483;
  assign n26485 = ~n26482 & n26484;
  assign n26486 = pi627 & ~n26386;
  assign n26487 = ~n26485 & n26486;
  assign n26488 = ~n26481 & ~n26487;
  assign n26489 = pi781 & ~n26488;
  assign n26490 = ~pi781 & ~n26475;
  assign n26491 = ~n26489 & ~n26490;
  assign n26492 = pi619 & ~n26491;
  assign n26493 = ~pi619 & n26417;
  assign n26494 = pi1159 & ~n26493;
  assign n26495 = ~n26492 & n26494;
  assign n26496 = pi648 & ~n26394;
  assign n26497 = ~n26495 & n26496;
  assign n26498 = ~pi619 & ~n26491;
  assign n26499 = pi619 & n26417;
  assign n26500 = ~pi1159 & ~n26499;
  assign n26501 = ~n26498 & n26500;
  assign n26502 = ~pi648 & ~n26392;
  assign n26503 = ~n26501 & n26502;
  assign n26504 = pi789 & ~n26503;
  assign n26505 = ~n26497 & n26504;
  assign n26506 = ~pi789 & n26491;
  assign n26507 = n17817 & ~n26506;
  assign n26508 = ~n26505 & n26507;
  assign n26509 = ~n26444 & ~n26508;
  assign n26510 = ~n20205 & ~n26509;
  assign n26511 = n17856 & ~n26400;
  assign n26512 = n20693 & n26419;
  assign n26513 = ~n26511 & ~n26512;
  assign n26514 = ~pi629 & ~n26513;
  assign n26515 = n20697 & n26419;
  assign n26516 = n17855 & ~n26400;
  assign n26517 = ~n26515 & ~n26516;
  assign n26518 = pi629 & ~n26517;
  assign n26519 = ~n26514 & ~n26518;
  assign n26520 = pi792 & ~n26519;
  assign n26521 = n20207 & ~n26520;
  assign n26522 = ~n26510 & n26521;
  assign n26523 = ~n26432 & ~n26522;
  assign n26524 = pi644 & n26523;
  assign n26525 = ~pi787 & ~n26420;
  assign n26526 = pi787 & ~n26429;
  assign n26527 = ~n26525 & ~n26526;
  assign n26528 = ~pi644 & n26527;
  assign n26529 = pi715 & ~n26528;
  assign n26530 = ~n26524 & n26529;
  assign n26531 = ~n17652 & ~n26403;
  assign n26532 = n17652 & n26369;
  assign n26533 = ~n26531 & ~n26532;
  assign n26534 = pi644 & ~n26533;
  assign n26535 = ~pi644 & n26369;
  assign n26536 = ~pi715 & ~n26535;
  assign n26537 = ~n26534 & n26536;
  assign n26538 = pi1160 & ~n26537;
  assign n26539 = ~n26530 & n26538;
  assign n26540 = ~pi644 & n26523;
  assign n26541 = pi644 & n26527;
  assign n26542 = ~pi715 & ~n26541;
  assign n26543 = ~n26540 & n26542;
  assign n26544 = ~pi644 & ~n26533;
  assign n26545 = pi644 & n26369;
  assign n26546 = pi715 & ~n26545;
  assign n26547 = ~n26544 & n26546;
  assign n26548 = ~pi1160 & ~n26547;
  assign n26549 = ~n26543 & n26548;
  assign n26550 = ~n26539 & ~n26549;
  assign n26551 = pi790 & ~n26550;
  assign n26552 = ~pi790 & n26523;
  assign n26553 = pi832 & ~n26552;
  assign n26554 = ~n26551 & n26553;
  assign n26555 = ~pi181 & ~n17406;
  assign n26556 = n17539 & ~n26555;
  assign n26557 = ~pi709 & n3267;
  assign n26558 = n26555 & ~n26557;
  assign n26559 = pi181 & ~n17976;
  assign n26560 = ~pi38 & ~n26559;
  assign n26561 = n3267 & ~n26560;
  assign n26562 = ~pi181 & n17972;
  assign n26563 = ~n26561 & ~n26562;
  assign n26564 = ~pi181 & ~n17280;
  assign n26565 = n17392 & ~n26564;
  assign n26566 = ~pi709 & ~n26565;
  assign n26567 = ~n26563 & n26566;
  assign n26568 = ~n26558 & ~n26567;
  assign n26569 = ~pi778 & n26568;
  assign n26570 = pi625 & ~n26568;
  assign n26571 = ~pi625 & n26555;
  assign n26572 = pi1153 & ~n26571;
  assign n26573 = ~n26570 & n26572;
  assign n26574 = ~pi625 & ~n26568;
  assign n26575 = pi625 & n26555;
  assign n26576 = ~pi1153 & ~n26575;
  assign n26577 = ~n26574 & n26576;
  assign n26578 = ~n26573 & ~n26577;
  assign n26579 = pi778 & ~n26578;
  assign n26580 = ~n26569 & ~n26579;
  assign n26581 = ~n17466 & ~n26580;
  assign n26582 = n17466 & ~n26555;
  assign n26583 = ~n26581 & ~n26582;
  assign n26584 = ~n17503 & n26583;
  assign n26585 = n17503 & n26555;
  assign n26586 = ~n26584 & ~n26585;
  assign n26587 = ~n17539 & n26586;
  assign n26588 = ~n26556 & ~n26587;
  assign n26589 = ~n17582 & n26588;
  assign n26590 = n17582 & n26555;
  assign n26591 = ~n26589 & ~n26590;
  assign n26592 = ~pi792 & n26591;
  assign n26593 = pi628 & ~n26591;
  assign n26594 = ~pi628 & n26555;
  assign n26595 = pi1156 & ~n26594;
  assign n26596 = ~n26593 & n26595;
  assign n26597 = ~pi628 & ~n26591;
  assign n26598 = pi628 & n26555;
  assign n26599 = ~pi1156 & ~n26598;
  assign n26600 = ~n26597 & n26599;
  assign n26601 = ~n26596 & ~n26600;
  assign n26602 = pi792 & ~n26601;
  assign n26603 = ~n26592 & ~n26602;
  assign n26604 = ~pi647 & ~n26603;
  assign n26605 = pi647 & ~n26555;
  assign n26606 = ~n26604 & ~n26605;
  assign n26607 = ~pi1157 & n26606;
  assign n26608 = pi647 & ~n26603;
  assign n26609 = ~pi647 & ~n26555;
  assign n26610 = ~n26608 & ~n26609;
  assign n26611 = pi1157 & n26610;
  assign n26612 = ~n26607 & ~n26611;
  assign n26613 = pi787 & ~n26612;
  assign n26614 = ~pi787 & n26603;
  assign n26615 = ~n26613 & ~n26614;
  assign n26616 = ~pi644 & ~n26615;
  assign n26617 = pi715 & ~n26616;
  assign n26618 = pi181 & ~n3267;
  assign n26619 = pi754 & n17199;
  assign n26620 = pi181 & n17273;
  assign n26621 = ~n26619 & ~n26620;
  assign n26622 = pi39 & ~n26621;
  assign n26623 = ~pi181 & ~pi754;
  assign n26624 = n17242 & n26623;
  assign n26625 = pi181 & pi754;
  assign n26626 = pi181 & ~n17086;
  assign n26627 = ~n21648 & ~n26626;
  assign n26628 = ~pi39 & ~n26627;
  assign n26629 = ~n26625 & ~n26628;
  assign n26630 = ~n26624 & n26629;
  assign n26631 = ~n26622 & n26630;
  assign n26632 = ~pi38 & ~n26631;
  assign n26633 = ~pi754 & n17282;
  assign n26634 = pi38 & ~n26564;
  assign n26635 = ~n26633 & n26634;
  assign n26636 = ~n26632 & ~n26635;
  assign n26637 = n3267 & ~n26636;
  assign n26638 = ~n26618 & ~n26637;
  assign n26639 = ~n17438 & ~n26638;
  assign n26640 = n17438 & ~n26555;
  assign n26641 = ~n26639 & ~n26640;
  assign n26642 = ~pi785 & ~n26641;
  assign n26643 = ~n17439 & ~n26555;
  assign n26644 = pi609 & n26639;
  assign n26645 = ~n26643 & ~n26644;
  assign n26646 = pi1155 & ~n26645;
  assign n26647 = ~n17451 & ~n26555;
  assign n26648 = ~pi609 & n26639;
  assign n26649 = ~n26647 & ~n26648;
  assign n26650 = ~pi1155 & ~n26649;
  assign n26651 = ~n26646 & ~n26650;
  assign n26652 = pi785 & ~n26651;
  assign n26653 = ~n26642 & ~n26652;
  assign n26654 = ~pi781 & ~n26653;
  assign n26655 = pi618 & n26653;
  assign n26656 = ~pi618 & n26555;
  assign n26657 = pi1154 & ~n26656;
  assign n26658 = ~n26655 & n26657;
  assign n26659 = ~pi618 & n26653;
  assign n26660 = pi618 & n26555;
  assign n26661 = ~pi1154 & ~n26660;
  assign n26662 = ~n26659 & n26661;
  assign n26663 = ~n26658 & ~n26662;
  assign n26664 = pi781 & ~n26663;
  assign n26665 = ~n26654 & ~n26664;
  assign n26666 = ~pi789 & ~n26665;
  assign n26667 = pi619 & n26665;
  assign n26668 = ~pi619 & n26555;
  assign n26669 = pi1159 & ~n26668;
  assign n26670 = ~n26667 & n26669;
  assign n26671 = ~pi619 & n26665;
  assign n26672 = pi619 & n26555;
  assign n26673 = ~pi1159 & ~n26672;
  assign n26674 = ~n26671 & n26673;
  assign n26675 = ~n26670 & ~n26674;
  assign n26676 = pi789 & ~n26675;
  assign n26677 = ~n26666 & ~n26676;
  assign n26678 = ~n17816 & n26677;
  assign n26679 = n17816 & n26555;
  assign n26680 = ~n26678 & ~n26679;
  assign n26681 = ~n17610 & ~n26680;
  assign n26682 = n17610 & n26555;
  assign n26683 = ~n26681 & ~n26682;
  assign n26684 = ~n17652 & ~n26683;
  assign n26685 = n17652 & n26555;
  assign n26686 = ~n26684 & ~n26685;
  assign n26687 = pi644 & ~n26686;
  assign n26688 = ~pi644 & n26555;
  assign n26689 = ~pi715 & ~n26688;
  assign n26690 = ~n26687 & n26689;
  assign n26691 = pi1160 & ~n26690;
  assign n26692 = ~n26617 & n26691;
  assign n26693 = pi644 & ~n26615;
  assign n26694 = ~pi715 & ~n26693;
  assign n26695 = ~pi644 & ~n26686;
  assign n26696 = pi644 & n26555;
  assign n26697 = pi715 & ~n26696;
  assign n26698 = ~n26695 & n26697;
  assign n26699 = ~pi1160 & ~n26698;
  assign n26700 = ~n26694 & n26699;
  assign n26701 = ~n26692 & ~n26700;
  assign n26702 = pi790 & ~n26701;
  assign n26703 = pi644 & n26691;
  assign n26704 = ~pi644 & n26699;
  assign n26705 = pi790 & ~n26704;
  assign n26706 = ~n26703 & n26705;
  assign n26707 = ~n20409 & n26680;
  assign n26708 = ~pi629 & n26596;
  assign n26709 = pi629 & n26600;
  assign n26710 = ~n26708 & ~n26709;
  assign n26711 = ~n26707 & n26710;
  assign n26712 = pi792 & ~n26711;
  assign n26713 = pi709 & n26636;
  assign n26714 = ~pi181 & n16687;
  assign n26715 = pi181 & n16799;
  assign n26716 = pi754 & ~n26715;
  assign n26717 = ~n26714 & n26716;
  assign n26718 = pi181 & n16879;
  assign n26719 = ~pi181 & ~n16944;
  assign n26720 = ~pi754 & ~n26719;
  assign n26721 = ~n26718 & n26720;
  assign n26722 = pi39 & ~n26721;
  assign n26723 = ~n26717 & n26722;
  assign n26724 = ~pi181 & ~n17088;
  assign n26725 = pi181 & ~n17059;
  assign n26726 = pi754 & ~n26725;
  assign n26727 = ~n26724 & n26726;
  assign n26728 = ~pi181 & n17092;
  assign n26729 = pi181 & n17094;
  assign n26730 = ~pi754 & ~n26729;
  assign n26731 = ~n26728 & n26730;
  assign n26732 = ~n26727 & ~n26731;
  assign n26733 = ~pi39 & ~n26732;
  assign n26734 = ~pi38 & ~n26733;
  assign n26735 = ~n26723 & n26734;
  assign n26736 = ~pi754 & ~n16905;
  assign n26737 = n19230 & ~n26736;
  assign n26738 = ~pi181 & ~n26737;
  assign n26739 = ~n16787 & ~n26370;
  assign n26740 = pi181 & ~n26739;
  assign n26741 = n6234 & n26740;
  assign n26742 = pi38 & ~n26741;
  assign n26743 = ~n26738 & n26742;
  assign n26744 = ~pi709 & ~n26743;
  assign n26745 = ~n26735 & n26744;
  assign n26746 = n3267 & ~n26745;
  assign n26747 = ~n26713 & n26746;
  assign n26748 = ~n26618 & ~n26747;
  assign n26749 = ~pi625 & n26748;
  assign n26750 = pi625 & n26638;
  assign n26751 = ~pi1153 & ~n26750;
  assign n26752 = ~n26749 & n26751;
  assign n26753 = ~pi608 & ~n26573;
  assign n26754 = ~n26752 & n26753;
  assign n26755 = pi625 & n26748;
  assign n26756 = ~pi625 & n26638;
  assign n26757 = pi1153 & ~n26756;
  assign n26758 = ~n26755 & n26757;
  assign n26759 = pi608 & ~n26577;
  assign n26760 = ~n26758 & n26759;
  assign n26761 = ~n26754 & ~n26760;
  assign n26762 = pi778 & ~n26761;
  assign n26763 = ~pi778 & n26748;
  assign n26764 = ~n26762 & ~n26763;
  assign n26765 = ~pi609 & ~n26764;
  assign n26766 = pi609 & n26580;
  assign n26767 = ~pi1155 & ~n26766;
  assign n26768 = ~n26765 & n26767;
  assign n26769 = ~pi660 & ~n26646;
  assign n26770 = ~n26768 & n26769;
  assign n26771 = pi609 & ~n26764;
  assign n26772 = ~pi609 & n26580;
  assign n26773 = pi1155 & ~n26772;
  assign n26774 = ~n26771 & n26773;
  assign n26775 = pi660 & ~n26650;
  assign n26776 = ~n26774 & n26775;
  assign n26777 = ~n26770 & ~n26776;
  assign n26778 = pi785 & ~n26777;
  assign n26779 = ~pi785 & ~n26764;
  assign n26780 = ~n26778 & ~n26779;
  assign n26781 = ~pi618 & ~n26780;
  assign n26782 = pi618 & n26583;
  assign n26783 = ~pi1154 & ~n26782;
  assign n26784 = ~n26781 & n26783;
  assign n26785 = ~pi627 & ~n26658;
  assign n26786 = ~n26784 & n26785;
  assign n26787 = pi618 & ~n26780;
  assign n26788 = ~pi618 & n26583;
  assign n26789 = pi1154 & ~n26788;
  assign n26790 = ~n26787 & n26789;
  assign n26791 = pi627 & ~n26662;
  assign n26792 = ~n26790 & n26791;
  assign n26793 = ~n26786 & ~n26792;
  assign n26794 = pi781 & ~n26793;
  assign n26795 = ~pi781 & ~n26780;
  assign n26796 = ~n26794 & ~n26795;
  assign n26797 = pi619 & ~n26796;
  assign n26798 = ~pi619 & ~n26586;
  assign n26799 = pi1159 & ~n26798;
  assign n26800 = ~n26797 & n26799;
  assign n26801 = pi648 & ~n26674;
  assign n26802 = ~n26800 & n26801;
  assign n26803 = ~pi619 & ~n26796;
  assign n26804 = pi619 & ~n26586;
  assign n26805 = ~pi1159 & ~n26804;
  assign n26806 = ~n26803 & n26805;
  assign n26807 = ~pi648 & ~n26670;
  assign n26808 = ~n26806 & n26807;
  assign n26809 = pi789 & ~n26808;
  assign n26810 = ~n26802 & n26809;
  assign n26811 = ~pi789 & n26796;
  assign n26812 = n17817 & ~n26811;
  assign n26813 = ~n26810 & n26812;
  assign n26814 = pi626 & ~n26677;
  assign n26815 = ~pi626 & ~n26555;
  assign n26816 = n17579 & ~n26815;
  assign n26817 = ~n26814 & n26816;
  assign n26818 = n17704 & n26588;
  assign n26819 = ~pi626 & ~n26677;
  assign n26820 = pi626 & ~n26555;
  assign n26821 = n17580 & ~n26820;
  assign n26822 = ~n26819 & n26821;
  assign n26823 = ~n26818 & ~n26822;
  assign n26824 = ~n26817 & n26823;
  assign n26825 = pi788 & ~n26824;
  assign n26826 = ~n20205 & ~n26825;
  assign n26827 = ~n26813 & n26826;
  assign n26828 = ~n26712 & ~n26827;
  assign n26829 = n20207 & ~n26828;
  assign n26830 = ~n20398 & n26683;
  assign n26831 = n17650 & ~n26606;
  assign n26832 = n17649 & ~n26610;
  assign n26833 = ~n26831 & ~n26832;
  assign n26834 = ~n26830 & n26833;
  assign n26835 = pi787 & ~n26834;
  assign n26836 = ~n26829 & ~n26835;
  assign n26837 = ~n26706 & n26836;
  assign n26838 = ~n26702 & ~n26837;
  assign n26839 = ~po1038 & ~n26838;
  assign n26840 = ~pi181 & po1038;
  assign n26841 = ~pi832 & ~n26840;
  assign n26842 = ~n26839 & n26841;
  assign po338 = ~n26554 & ~n26842;
  assign n26844 = ~pi182 & ~n2754;
  assign n26845 = ~pi756 & n16784;
  assign n26846 = ~n26844 & ~n26845;
  assign n26847 = ~n17706 & ~n26846;
  assign n26848 = ~pi785 & ~n26847;
  assign n26849 = n17451 & n26845;
  assign n26850 = n26847 & ~n26849;
  assign n26851 = pi1155 & ~n26850;
  assign n26852 = ~pi1155 & ~n26844;
  assign n26853 = ~n26849 & n26852;
  assign n26854 = ~n26851 & ~n26853;
  assign n26855 = pi785 & ~n26854;
  assign n26856 = ~n26848 & ~n26855;
  assign n26857 = ~pi781 & ~n26856;
  assign n26858 = ~n17721 & n26856;
  assign n26859 = pi1154 & ~n26858;
  assign n26860 = ~n17724 & n26856;
  assign n26861 = ~pi1154 & ~n26860;
  assign n26862 = ~n26859 & ~n26861;
  assign n26863 = pi781 & ~n26862;
  assign n26864 = ~n26857 & ~n26863;
  assign n26865 = ~pi789 & ~n26864;
  assign n26866 = ~n22890 & n26864;
  assign n26867 = pi1159 & ~n26866;
  assign n26868 = ~n22893 & n26864;
  assign n26869 = ~pi1159 & ~n26868;
  assign n26870 = ~n26867 & ~n26869;
  assign n26871 = pi789 & ~n26870;
  assign n26872 = ~n26865 & ~n26871;
  assign n26873 = ~n17816 & n26872;
  assign n26874 = n17816 & n26844;
  assign n26875 = ~n26873 & ~n26874;
  assign n26876 = ~n17610 & ~n26875;
  assign n26877 = n17610 & n26844;
  assign n26878 = ~n26876 & ~n26877;
  assign n26879 = ~n20398 & n26878;
  assign n26880 = ~pi734 & n16786;
  assign n26881 = ~n26844 & ~n26880;
  assign n26882 = ~pi778 & ~n26881;
  assign n26883 = ~pi625 & n26880;
  assign n26884 = ~n26881 & ~n26883;
  assign n26885 = pi1153 & ~n26884;
  assign n26886 = ~pi1153 & ~n26844;
  assign n26887 = ~n26883 & n26886;
  assign n26888 = pi778 & ~n26887;
  assign n26889 = ~n26885 & n26888;
  assign n26890 = ~n26882 & ~n26889;
  assign n26891 = ~n17692 & ~n26890;
  assign n26892 = ~n17694 & n26891;
  assign n26893 = ~n17696 & n26892;
  assign n26894 = ~n17828 & n26893;
  assign n26895 = ~n17859 & n26894;
  assign n26896 = ~pi647 & n26895;
  assign n26897 = pi647 & n26844;
  assign n26898 = ~pi1157 & ~n26897;
  assign n26899 = ~n26896 & n26898;
  assign n26900 = pi647 & ~n26895;
  assign n26901 = ~pi647 & ~n26844;
  assign n26902 = ~n26900 & ~n26901;
  assign n26903 = pi1157 & ~n26902;
  assign n26904 = ~n26899 & ~n26903;
  assign n26905 = ~n17651 & ~n26904;
  assign n26906 = ~n26879 & ~n26905;
  assign n26907 = pi787 & ~n26906;
  assign n26908 = pi626 & ~n26872;
  assign n26909 = ~pi626 & ~n26844;
  assign n26910 = n17579 & ~n26909;
  assign n26911 = ~n26908 & n26910;
  assign n26912 = n17704 & n26893;
  assign n26913 = ~pi626 & ~n26872;
  assign n26914 = pi626 & ~n26844;
  assign n26915 = n17580 & ~n26914;
  assign n26916 = ~n26913 & n26915;
  assign n26917 = ~n26912 & ~n26916;
  assign n26918 = ~n26911 & n26917;
  assign n26919 = pi788 & ~n26918;
  assign n26920 = ~n16521 & ~n26881;
  assign n26921 = pi625 & n26920;
  assign n26922 = n26846 & ~n26920;
  assign n26923 = ~n26921 & ~n26922;
  assign n26924 = n26886 & ~n26923;
  assign n26925 = ~pi608 & ~n26885;
  assign n26926 = ~n26924 & n26925;
  assign n26927 = pi1153 & n26846;
  assign n26928 = ~n26921 & n26927;
  assign n26929 = pi608 & ~n26887;
  assign n26930 = ~n26928 & n26929;
  assign n26931 = ~n26926 & ~n26930;
  assign n26932 = pi778 & ~n26931;
  assign n26933 = ~pi778 & ~n26922;
  assign n26934 = ~n26932 & ~n26933;
  assign n26935 = ~pi609 & ~n26934;
  assign n26936 = pi609 & ~n26890;
  assign n26937 = ~pi1155 & ~n26936;
  assign n26938 = ~n26935 & n26937;
  assign n26939 = ~pi660 & ~n26851;
  assign n26940 = ~n26938 & n26939;
  assign n26941 = pi609 & ~n26934;
  assign n26942 = ~pi609 & ~n26890;
  assign n26943 = pi1155 & ~n26942;
  assign n26944 = ~n26941 & n26943;
  assign n26945 = pi660 & ~n26853;
  assign n26946 = ~n26944 & n26945;
  assign n26947 = ~n26940 & ~n26946;
  assign n26948 = pi785 & ~n26947;
  assign n26949 = ~pi785 & ~n26934;
  assign n26950 = ~n26948 & ~n26949;
  assign n26951 = ~pi618 & ~n26950;
  assign n26952 = pi618 & n26891;
  assign n26953 = ~pi1154 & ~n26952;
  assign n26954 = ~n26951 & n26953;
  assign n26955 = ~pi627 & ~n26859;
  assign n26956 = ~n26954 & n26955;
  assign n26957 = pi618 & ~n26950;
  assign n26958 = ~pi618 & n26891;
  assign n26959 = pi1154 & ~n26958;
  assign n26960 = ~n26957 & n26959;
  assign n26961 = pi627 & ~n26861;
  assign n26962 = ~n26960 & n26961;
  assign n26963 = ~n26956 & ~n26962;
  assign n26964 = pi781 & ~n26963;
  assign n26965 = ~pi781 & ~n26950;
  assign n26966 = ~n26964 & ~n26965;
  assign n26967 = pi619 & ~n26966;
  assign n26968 = ~pi619 & n26892;
  assign n26969 = pi1159 & ~n26968;
  assign n26970 = ~n26967 & n26969;
  assign n26971 = pi648 & ~n26869;
  assign n26972 = ~n26970 & n26971;
  assign n26973 = ~pi619 & ~n26966;
  assign n26974 = pi619 & n26892;
  assign n26975 = ~pi1159 & ~n26974;
  assign n26976 = ~n26973 & n26975;
  assign n26977 = ~pi648 & ~n26867;
  assign n26978 = ~n26976 & n26977;
  assign n26979 = pi789 & ~n26978;
  assign n26980 = ~n26972 & n26979;
  assign n26981 = ~pi789 & n26966;
  assign n26982 = n17817 & ~n26981;
  assign n26983 = ~n26980 & n26982;
  assign n26984 = ~n26919 & ~n26983;
  assign n26985 = ~n20205 & ~n26984;
  assign n26986 = n17856 & ~n26875;
  assign n26987 = n20693 & n26894;
  assign n26988 = ~n26986 & ~n26987;
  assign n26989 = ~pi629 & ~n26988;
  assign n26990 = n20697 & n26894;
  assign n26991 = n17855 & ~n26875;
  assign n26992 = ~n26990 & ~n26991;
  assign n26993 = pi629 & ~n26992;
  assign n26994 = ~n26989 & ~n26993;
  assign n26995 = pi792 & ~n26994;
  assign n26996 = n20207 & ~n26995;
  assign n26997 = ~n26985 & n26996;
  assign n26998 = ~n26907 & ~n26997;
  assign n26999 = pi644 & n26998;
  assign n27000 = ~pi787 & ~n26895;
  assign n27001 = pi787 & ~n26904;
  assign n27002 = ~n27000 & ~n27001;
  assign n27003 = ~pi644 & n27002;
  assign n27004 = pi715 & ~n27003;
  assign n27005 = ~n26999 & n27004;
  assign n27006 = ~n17652 & ~n26878;
  assign n27007 = n17652 & n26844;
  assign n27008 = ~n27006 & ~n27007;
  assign n27009 = pi644 & ~n27008;
  assign n27010 = ~pi644 & n26844;
  assign n27011 = ~pi715 & ~n27010;
  assign n27012 = ~n27009 & n27011;
  assign n27013 = pi1160 & ~n27012;
  assign n27014 = ~n27005 & n27013;
  assign n27015 = ~pi644 & n26998;
  assign n27016 = pi644 & n27002;
  assign n27017 = ~pi715 & ~n27016;
  assign n27018 = ~n27015 & n27017;
  assign n27019 = ~pi644 & ~n27008;
  assign n27020 = pi644 & n26844;
  assign n27021 = pi715 & ~n27020;
  assign n27022 = ~n27019 & n27021;
  assign n27023 = ~pi1160 & ~n27022;
  assign n27024 = ~n27018 & n27023;
  assign n27025 = ~n27014 & ~n27024;
  assign n27026 = pi790 & ~n27025;
  assign n27027 = ~pi790 & n26998;
  assign n27028 = pi832 & ~n27027;
  assign n27029 = ~n27026 & n27028;
  assign n27030 = ~pi182 & ~n17406;
  assign n27031 = n17539 & ~n27030;
  assign n27032 = ~pi734 & n3267;
  assign n27033 = n27030 & ~n27032;
  assign n27034 = pi182 & ~n17976;
  assign n27035 = ~pi38 & ~n27034;
  assign n27036 = n3267 & ~n27035;
  assign n27037 = ~pi182 & n17972;
  assign n27038 = ~n27036 & ~n27037;
  assign n27039 = ~pi182 & ~n17280;
  assign n27040 = n17392 & ~n27039;
  assign n27041 = ~pi734 & ~n27040;
  assign n27042 = ~n27038 & n27041;
  assign n27043 = ~n27033 & ~n27042;
  assign n27044 = ~pi778 & n27043;
  assign n27045 = pi625 & ~n27043;
  assign n27046 = ~pi625 & n27030;
  assign n27047 = pi1153 & ~n27046;
  assign n27048 = ~n27045 & n27047;
  assign n27049 = ~pi625 & ~n27043;
  assign n27050 = pi625 & n27030;
  assign n27051 = ~pi1153 & ~n27050;
  assign n27052 = ~n27049 & n27051;
  assign n27053 = ~n27048 & ~n27052;
  assign n27054 = pi778 & ~n27053;
  assign n27055 = ~n27044 & ~n27054;
  assign n27056 = ~n17466 & ~n27055;
  assign n27057 = n17466 & ~n27030;
  assign n27058 = ~n27056 & ~n27057;
  assign n27059 = ~n17503 & n27058;
  assign n27060 = n17503 & n27030;
  assign n27061 = ~n27059 & ~n27060;
  assign n27062 = ~n17539 & n27061;
  assign n27063 = ~n27031 & ~n27062;
  assign n27064 = ~n17582 & n27063;
  assign n27065 = n17582 & n27030;
  assign n27066 = ~n27064 & ~n27065;
  assign n27067 = ~pi792 & n27066;
  assign n27068 = pi628 & ~n27066;
  assign n27069 = ~pi628 & n27030;
  assign n27070 = pi1156 & ~n27069;
  assign n27071 = ~n27068 & n27070;
  assign n27072 = ~pi628 & ~n27066;
  assign n27073 = pi628 & n27030;
  assign n27074 = ~pi1156 & ~n27073;
  assign n27075 = ~n27072 & n27074;
  assign n27076 = ~n27071 & ~n27075;
  assign n27077 = pi792 & ~n27076;
  assign n27078 = ~n27067 & ~n27077;
  assign n27079 = ~pi647 & ~n27078;
  assign n27080 = pi647 & ~n27030;
  assign n27081 = ~n27079 & ~n27080;
  assign n27082 = ~pi1157 & n27081;
  assign n27083 = pi647 & ~n27078;
  assign n27084 = ~pi647 & ~n27030;
  assign n27085 = ~n27083 & ~n27084;
  assign n27086 = pi1157 & n27085;
  assign n27087 = ~n27082 & ~n27086;
  assign n27088 = pi787 & ~n27087;
  assign n27089 = ~pi787 & n27078;
  assign n27090 = ~n27088 & ~n27089;
  assign n27091 = ~pi644 & ~n27090;
  assign n27092 = pi715 & ~n27091;
  assign n27093 = pi182 & ~n3267;
  assign n27094 = ~pi756 & n17282;
  assign n27095 = ~n27039 & ~n27094;
  assign n27096 = pi38 & ~n27095;
  assign n27097 = ~pi182 & n17242;
  assign n27098 = pi182 & ~n17275;
  assign n27099 = ~pi756 & ~n27098;
  assign n27100 = ~n27097 & n27099;
  assign n27101 = ~pi182 & pi756;
  assign n27102 = ~n17201 & n27101;
  assign n27103 = ~n27100 & ~n27102;
  assign n27104 = ~pi38 & ~n27103;
  assign n27105 = ~n27096 & ~n27104;
  assign n27106 = n3267 & n27105;
  assign n27107 = ~n27093 & ~n27106;
  assign n27108 = ~n17438 & ~n27107;
  assign n27109 = n17438 & ~n27030;
  assign n27110 = ~n27108 & ~n27109;
  assign n27111 = ~pi785 & ~n27110;
  assign n27112 = ~n17439 & ~n27030;
  assign n27113 = pi609 & n27108;
  assign n27114 = ~n27112 & ~n27113;
  assign n27115 = pi1155 & ~n27114;
  assign n27116 = ~n17451 & ~n27030;
  assign n27117 = ~pi609 & n27108;
  assign n27118 = ~n27116 & ~n27117;
  assign n27119 = ~pi1155 & ~n27118;
  assign n27120 = ~n27115 & ~n27119;
  assign n27121 = pi785 & ~n27120;
  assign n27122 = ~n27111 & ~n27121;
  assign n27123 = ~pi781 & ~n27122;
  assign n27124 = pi618 & n27122;
  assign n27125 = ~pi618 & n27030;
  assign n27126 = pi1154 & ~n27125;
  assign n27127 = ~n27124 & n27126;
  assign n27128 = ~pi618 & n27122;
  assign n27129 = pi618 & n27030;
  assign n27130 = ~pi1154 & ~n27129;
  assign n27131 = ~n27128 & n27130;
  assign n27132 = ~n27127 & ~n27131;
  assign n27133 = pi781 & ~n27132;
  assign n27134 = ~n27123 & ~n27133;
  assign n27135 = ~pi789 & ~n27134;
  assign n27136 = pi619 & n27134;
  assign n27137 = ~pi619 & n27030;
  assign n27138 = pi1159 & ~n27137;
  assign n27139 = ~n27136 & n27138;
  assign n27140 = ~pi619 & n27134;
  assign n27141 = pi619 & n27030;
  assign n27142 = ~pi1159 & ~n27141;
  assign n27143 = ~n27140 & n27142;
  assign n27144 = ~n27139 & ~n27143;
  assign n27145 = pi789 & ~n27144;
  assign n27146 = ~n27135 & ~n27145;
  assign n27147 = ~n17816 & n27146;
  assign n27148 = n17816 & n27030;
  assign n27149 = ~n27147 & ~n27148;
  assign n27150 = ~n17610 & ~n27149;
  assign n27151 = n17610 & n27030;
  assign n27152 = ~n27150 & ~n27151;
  assign n27153 = ~n17652 & ~n27152;
  assign n27154 = n17652 & n27030;
  assign n27155 = ~n27153 & ~n27154;
  assign n27156 = pi644 & ~n27155;
  assign n27157 = ~pi644 & n27030;
  assign n27158 = ~pi715 & ~n27157;
  assign n27159 = ~n27156 & n27158;
  assign n27160 = pi1160 & ~n27159;
  assign n27161 = ~n27092 & n27160;
  assign n27162 = pi644 & ~n27090;
  assign n27163 = ~pi715 & ~n27162;
  assign n27164 = ~pi644 & ~n27155;
  assign n27165 = pi644 & n27030;
  assign n27166 = pi715 & ~n27165;
  assign n27167 = ~n27164 & n27166;
  assign n27168 = ~pi1160 & ~n27167;
  assign n27169 = ~n27163 & n27168;
  assign n27170 = ~n27161 & ~n27169;
  assign n27171 = pi790 & ~n27170;
  assign n27172 = pi644 & n27160;
  assign n27173 = ~pi644 & n27168;
  assign n27174 = pi790 & ~n27173;
  assign n27175 = ~n27172 & n27174;
  assign n27176 = ~n20409 & n27149;
  assign n27177 = ~pi629 & n27071;
  assign n27178 = pi629 & n27075;
  assign n27179 = ~n27177 & ~n27178;
  assign n27180 = ~n27176 & n27179;
  assign n27181 = pi792 & ~n27180;
  assign n27182 = pi734 & ~n27105;
  assign n27183 = ~pi182 & n16687;
  assign n27184 = pi182 & n16799;
  assign n27185 = pi756 & ~n27184;
  assign n27186 = ~n27183 & n27185;
  assign n27187 = pi182 & n16879;
  assign n27188 = ~pi182 & ~n16944;
  assign n27189 = ~pi756 & ~n27188;
  assign n27190 = ~n27187 & n27189;
  assign n27191 = pi39 & ~n27190;
  assign n27192 = ~n27186 & n27191;
  assign n27193 = ~pi182 & ~n17088;
  assign n27194 = pi182 & ~n17059;
  assign n27195 = pi756 & ~n27194;
  assign n27196 = ~n27193 & n27195;
  assign n27197 = ~pi182 & n17092;
  assign n27198 = pi182 & n17094;
  assign n27199 = ~pi756 & ~n27198;
  assign n27200 = ~n27197 & n27199;
  assign n27201 = ~n27196 & ~n27200;
  assign n27202 = ~pi39 & ~n27201;
  assign n27203 = ~pi38 & ~n27202;
  assign n27204 = ~n27192 & n27203;
  assign n27205 = ~pi756 & ~n16905;
  assign n27206 = n19230 & ~n27205;
  assign n27207 = ~pi182 & ~n27206;
  assign n27208 = ~n16787 & ~n26845;
  assign n27209 = pi182 & ~n27208;
  assign n27210 = n6234 & n27209;
  assign n27211 = pi38 & ~n27210;
  assign n27212 = ~n27207 & n27211;
  assign n27213 = ~pi734 & ~n27212;
  assign n27214 = ~n27204 & n27213;
  assign n27215 = n3267 & ~n27214;
  assign n27216 = ~n27182 & n27215;
  assign n27217 = ~n27093 & ~n27216;
  assign n27218 = ~pi625 & n27217;
  assign n27219 = pi625 & n27107;
  assign n27220 = ~pi1153 & ~n27219;
  assign n27221 = ~n27218 & n27220;
  assign n27222 = ~pi608 & ~n27048;
  assign n27223 = ~n27221 & n27222;
  assign n27224 = pi625 & n27217;
  assign n27225 = ~pi625 & n27107;
  assign n27226 = pi1153 & ~n27225;
  assign n27227 = ~n27224 & n27226;
  assign n27228 = pi608 & ~n27052;
  assign n27229 = ~n27227 & n27228;
  assign n27230 = ~n27223 & ~n27229;
  assign n27231 = pi778 & ~n27230;
  assign n27232 = ~pi778 & n27217;
  assign n27233 = ~n27231 & ~n27232;
  assign n27234 = ~pi609 & ~n27233;
  assign n27235 = pi609 & n27055;
  assign n27236 = ~pi1155 & ~n27235;
  assign n27237 = ~n27234 & n27236;
  assign n27238 = ~pi660 & ~n27115;
  assign n27239 = ~n27237 & n27238;
  assign n27240 = pi609 & ~n27233;
  assign n27241 = ~pi609 & n27055;
  assign n27242 = pi1155 & ~n27241;
  assign n27243 = ~n27240 & n27242;
  assign n27244 = pi660 & ~n27119;
  assign n27245 = ~n27243 & n27244;
  assign n27246 = ~n27239 & ~n27245;
  assign n27247 = pi785 & ~n27246;
  assign n27248 = ~pi785 & ~n27233;
  assign n27249 = ~n27247 & ~n27248;
  assign n27250 = ~pi618 & ~n27249;
  assign n27251 = pi618 & n27058;
  assign n27252 = ~pi1154 & ~n27251;
  assign n27253 = ~n27250 & n27252;
  assign n27254 = ~pi627 & ~n27127;
  assign n27255 = ~n27253 & n27254;
  assign n27256 = pi618 & ~n27249;
  assign n27257 = ~pi618 & n27058;
  assign n27258 = pi1154 & ~n27257;
  assign n27259 = ~n27256 & n27258;
  assign n27260 = pi627 & ~n27131;
  assign n27261 = ~n27259 & n27260;
  assign n27262 = ~n27255 & ~n27261;
  assign n27263 = pi781 & ~n27262;
  assign n27264 = ~pi781 & ~n27249;
  assign n27265 = ~n27263 & ~n27264;
  assign n27266 = pi619 & ~n27265;
  assign n27267 = ~pi619 & ~n27061;
  assign n27268 = pi1159 & ~n27267;
  assign n27269 = ~n27266 & n27268;
  assign n27270 = pi648 & ~n27143;
  assign n27271 = ~n27269 & n27270;
  assign n27272 = ~pi619 & ~n27265;
  assign n27273 = pi619 & ~n27061;
  assign n27274 = ~pi1159 & ~n27273;
  assign n27275 = ~n27272 & n27274;
  assign n27276 = ~pi648 & ~n27139;
  assign n27277 = ~n27275 & n27276;
  assign n27278 = pi789 & ~n27277;
  assign n27279 = ~n27271 & n27278;
  assign n27280 = ~pi789 & n27265;
  assign n27281 = n17817 & ~n27280;
  assign n27282 = ~n27279 & n27281;
  assign n27283 = pi626 & ~n27146;
  assign n27284 = ~pi626 & ~n27030;
  assign n27285 = n17579 & ~n27284;
  assign n27286 = ~n27283 & n27285;
  assign n27287 = n17704 & n27063;
  assign n27288 = ~pi626 & ~n27146;
  assign n27289 = pi626 & ~n27030;
  assign n27290 = n17580 & ~n27289;
  assign n27291 = ~n27288 & n27290;
  assign n27292 = ~n27287 & ~n27291;
  assign n27293 = ~n27286 & n27292;
  assign n27294 = pi788 & ~n27293;
  assign n27295 = ~n20205 & ~n27294;
  assign n27296 = ~n27282 & n27295;
  assign n27297 = ~n27181 & ~n27296;
  assign n27298 = n20207 & ~n27297;
  assign n27299 = ~n20398 & n27152;
  assign n27300 = n17650 & ~n27081;
  assign n27301 = n17649 & ~n27085;
  assign n27302 = ~n27300 & ~n27301;
  assign n27303 = ~n27299 & n27302;
  assign n27304 = pi787 & ~n27303;
  assign n27305 = ~n27298 & ~n27304;
  assign n27306 = ~n27175 & n27305;
  assign n27307 = ~n27171 & ~n27306;
  assign n27308 = ~po1038 & ~n27307;
  assign n27309 = ~pi182 & po1038;
  assign n27310 = ~pi832 & ~n27309;
  assign n27311 = ~n27308 & n27310;
  assign po339 = ~n27029 & ~n27311;
  assign n27313 = ~pi183 & ~n2754;
  assign n27314 = ~pi755 & n16784;
  assign n27315 = ~n27313 & ~n27314;
  assign n27316 = ~n17706 & ~n27315;
  assign n27317 = ~pi785 & ~n27316;
  assign n27318 = n17451 & n27314;
  assign n27319 = n27316 & ~n27318;
  assign n27320 = pi1155 & ~n27319;
  assign n27321 = ~pi1155 & ~n27313;
  assign n27322 = ~n27318 & n27321;
  assign n27323 = ~n27320 & ~n27322;
  assign n27324 = pi785 & ~n27323;
  assign n27325 = ~n27317 & ~n27324;
  assign n27326 = ~pi781 & ~n27325;
  assign n27327 = ~n17721 & n27325;
  assign n27328 = pi1154 & ~n27327;
  assign n27329 = ~n17724 & n27325;
  assign n27330 = ~pi1154 & ~n27329;
  assign n27331 = ~n27328 & ~n27330;
  assign n27332 = pi781 & ~n27331;
  assign n27333 = ~n27326 & ~n27332;
  assign n27334 = ~pi789 & ~n27333;
  assign n27335 = ~n22890 & n27333;
  assign n27336 = pi1159 & ~n27335;
  assign n27337 = ~n22893 & n27333;
  assign n27338 = ~pi1159 & ~n27337;
  assign n27339 = ~n27336 & ~n27338;
  assign n27340 = pi789 & ~n27339;
  assign n27341 = ~n27334 & ~n27340;
  assign n27342 = ~n17816 & n27341;
  assign n27343 = n17816 & n27313;
  assign n27344 = ~n27342 & ~n27343;
  assign n27345 = ~n17610 & ~n27344;
  assign n27346 = n17610 & n27313;
  assign n27347 = ~n27345 & ~n27346;
  assign n27348 = ~n20398 & n27347;
  assign n27349 = ~pi725 & n16786;
  assign n27350 = ~n27313 & ~n27349;
  assign n27351 = ~pi778 & ~n27350;
  assign n27352 = ~pi625 & n27349;
  assign n27353 = ~n27350 & ~n27352;
  assign n27354 = pi1153 & ~n27353;
  assign n27355 = ~pi1153 & ~n27313;
  assign n27356 = ~n27352 & n27355;
  assign n27357 = pi778 & ~n27356;
  assign n27358 = ~n27354 & n27357;
  assign n27359 = ~n27351 & ~n27358;
  assign n27360 = ~n17692 & ~n27359;
  assign n27361 = ~n17694 & n27360;
  assign n27362 = ~n17696 & n27361;
  assign n27363 = ~n17828 & n27362;
  assign n27364 = ~n17859 & n27363;
  assign n27365 = ~pi647 & n27364;
  assign n27366 = pi647 & n27313;
  assign n27367 = ~pi1157 & ~n27366;
  assign n27368 = ~n27365 & n27367;
  assign n27369 = pi647 & ~n27364;
  assign n27370 = ~pi647 & ~n27313;
  assign n27371 = ~n27369 & ~n27370;
  assign n27372 = pi1157 & ~n27371;
  assign n27373 = ~n27368 & ~n27372;
  assign n27374 = ~n17651 & ~n27373;
  assign n27375 = ~n27348 & ~n27374;
  assign n27376 = pi787 & ~n27375;
  assign n27377 = pi626 & ~n27341;
  assign n27378 = ~pi626 & ~n27313;
  assign n27379 = n17579 & ~n27378;
  assign n27380 = ~n27377 & n27379;
  assign n27381 = n17704 & n27362;
  assign n27382 = ~pi626 & ~n27341;
  assign n27383 = pi626 & ~n27313;
  assign n27384 = n17580 & ~n27383;
  assign n27385 = ~n27382 & n27384;
  assign n27386 = ~n27381 & ~n27385;
  assign n27387 = ~n27380 & n27386;
  assign n27388 = pi788 & ~n27387;
  assign n27389 = ~n16521 & ~n27350;
  assign n27390 = pi625 & n27389;
  assign n27391 = n27315 & ~n27389;
  assign n27392 = ~n27390 & ~n27391;
  assign n27393 = n27355 & ~n27392;
  assign n27394 = ~pi608 & ~n27354;
  assign n27395 = ~n27393 & n27394;
  assign n27396 = pi1153 & n27315;
  assign n27397 = ~n27390 & n27396;
  assign n27398 = pi608 & ~n27356;
  assign n27399 = ~n27397 & n27398;
  assign n27400 = ~n27395 & ~n27399;
  assign n27401 = pi778 & ~n27400;
  assign n27402 = ~pi778 & ~n27391;
  assign n27403 = ~n27401 & ~n27402;
  assign n27404 = ~pi609 & ~n27403;
  assign n27405 = pi609 & ~n27359;
  assign n27406 = ~pi1155 & ~n27405;
  assign n27407 = ~n27404 & n27406;
  assign n27408 = ~pi660 & ~n27320;
  assign n27409 = ~n27407 & n27408;
  assign n27410 = pi609 & ~n27403;
  assign n27411 = ~pi609 & ~n27359;
  assign n27412 = pi1155 & ~n27411;
  assign n27413 = ~n27410 & n27412;
  assign n27414 = pi660 & ~n27322;
  assign n27415 = ~n27413 & n27414;
  assign n27416 = ~n27409 & ~n27415;
  assign n27417 = pi785 & ~n27416;
  assign n27418 = ~pi785 & ~n27403;
  assign n27419 = ~n27417 & ~n27418;
  assign n27420 = ~pi618 & ~n27419;
  assign n27421 = pi618 & n27360;
  assign n27422 = ~pi1154 & ~n27421;
  assign n27423 = ~n27420 & n27422;
  assign n27424 = ~pi627 & ~n27328;
  assign n27425 = ~n27423 & n27424;
  assign n27426 = pi618 & ~n27419;
  assign n27427 = ~pi618 & n27360;
  assign n27428 = pi1154 & ~n27427;
  assign n27429 = ~n27426 & n27428;
  assign n27430 = pi627 & ~n27330;
  assign n27431 = ~n27429 & n27430;
  assign n27432 = ~n27425 & ~n27431;
  assign n27433 = pi781 & ~n27432;
  assign n27434 = ~pi781 & ~n27419;
  assign n27435 = ~n27433 & ~n27434;
  assign n27436 = pi619 & ~n27435;
  assign n27437 = ~pi619 & n27361;
  assign n27438 = pi1159 & ~n27437;
  assign n27439 = ~n27436 & n27438;
  assign n27440 = pi648 & ~n27338;
  assign n27441 = ~n27439 & n27440;
  assign n27442 = ~pi619 & ~n27435;
  assign n27443 = pi619 & n27361;
  assign n27444 = ~pi1159 & ~n27443;
  assign n27445 = ~n27442 & n27444;
  assign n27446 = ~pi648 & ~n27336;
  assign n27447 = ~n27445 & n27446;
  assign n27448 = pi789 & ~n27447;
  assign n27449 = ~n27441 & n27448;
  assign n27450 = ~pi789 & n27435;
  assign n27451 = n17817 & ~n27450;
  assign n27452 = ~n27449 & n27451;
  assign n27453 = ~n27388 & ~n27452;
  assign n27454 = ~n20205 & ~n27453;
  assign n27455 = n17856 & ~n27344;
  assign n27456 = n20693 & n27363;
  assign n27457 = ~n27455 & ~n27456;
  assign n27458 = ~pi629 & ~n27457;
  assign n27459 = n20697 & n27363;
  assign n27460 = n17855 & ~n27344;
  assign n27461 = ~n27459 & ~n27460;
  assign n27462 = pi629 & ~n27461;
  assign n27463 = ~n27458 & ~n27462;
  assign n27464 = pi792 & ~n27463;
  assign n27465 = n20207 & ~n27464;
  assign n27466 = ~n27454 & n27465;
  assign n27467 = ~n27376 & ~n27466;
  assign n27468 = pi644 & n27467;
  assign n27469 = ~pi787 & ~n27364;
  assign n27470 = pi787 & ~n27373;
  assign n27471 = ~n27469 & ~n27470;
  assign n27472 = ~pi644 & n27471;
  assign n27473 = pi715 & ~n27472;
  assign n27474 = ~n27468 & n27473;
  assign n27475 = ~n17652 & ~n27347;
  assign n27476 = n17652 & n27313;
  assign n27477 = ~n27475 & ~n27476;
  assign n27478 = pi644 & ~n27477;
  assign n27479 = ~pi644 & n27313;
  assign n27480 = ~pi715 & ~n27479;
  assign n27481 = ~n27478 & n27480;
  assign n27482 = pi1160 & ~n27481;
  assign n27483 = ~n27474 & n27482;
  assign n27484 = ~pi644 & n27467;
  assign n27485 = pi644 & n27471;
  assign n27486 = ~pi715 & ~n27485;
  assign n27487 = ~n27484 & n27486;
  assign n27488 = ~pi644 & ~n27477;
  assign n27489 = pi644 & n27313;
  assign n27490 = pi715 & ~n27489;
  assign n27491 = ~n27488 & n27490;
  assign n27492 = ~pi1160 & ~n27491;
  assign n27493 = ~n27487 & n27492;
  assign n27494 = ~n27483 & ~n27493;
  assign n27495 = pi790 & ~n27494;
  assign n27496 = ~pi790 & n27467;
  assign n27497 = pi832 & ~n27496;
  assign n27498 = ~n27495 & n27497;
  assign n27499 = ~pi183 & ~n17406;
  assign n27500 = n17539 & ~n27499;
  assign n27501 = ~pi725 & n3267;
  assign n27502 = n27499 & ~n27501;
  assign n27503 = pi183 & ~n17976;
  assign n27504 = ~pi38 & ~n27503;
  assign n27505 = n3267 & ~n27504;
  assign n27506 = ~pi183 & n17972;
  assign n27507 = ~n27505 & ~n27506;
  assign n27508 = ~pi183 & ~n17280;
  assign n27509 = n17392 & ~n27508;
  assign n27510 = ~pi725 & ~n27509;
  assign n27511 = ~n27507 & n27510;
  assign n27512 = ~n27502 & ~n27511;
  assign n27513 = ~pi778 & n27512;
  assign n27514 = pi625 & ~n27512;
  assign n27515 = ~pi625 & n27499;
  assign n27516 = pi1153 & ~n27515;
  assign n27517 = ~n27514 & n27516;
  assign n27518 = ~pi625 & ~n27512;
  assign n27519 = pi625 & n27499;
  assign n27520 = ~pi1153 & ~n27519;
  assign n27521 = ~n27518 & n27520;
  assign n27522 = ~n27517 & ~n27521;
  assign n27523 = pi778 & ~n27522;
  assign n27524 = ~n27513 & ~n27523;
  assign n27525 = ~n17466 & ~n27524;
  assign n27526 = n17466 & ~n27499;
  assign n27527 = ~n27525 & ~n27526;
  assign n27528 = ~n17503 & n27527;
  assign n27529 = n17503 & n27499;
  assign n27530 = ~n27528 & ~n27529;
  assign n27531 = ~n17539 & n27530;
  assign n27532 = ~n27500 & ~n27531;
  assign n27533 = ~n17582 & n27532;
  assign n27534 = n17582 & n27499;
  assign n27535 = ~n27533 & ~n27534;
  assign n27536 = ~pi792 & n27535;
  assign n27537 = pi628 & ~n27535;
  assign n27538 = ~pi628 & n27499;
  assign n27539 = pi1156 & ~n27538;
  assign n27540 = ~n27537 & n27539;
  assign n27541 = ~pi628 & ~n27535;
  assign n27542 = pi628 & n27499;
  assign n27543 = ~pi1156 & ~n27542;
  assign n27544 = ~n27541 & n27543;
  assign n27545 = ~n27540 & ~n27544;
  assign n27546 = pi792 & ~n27545;
  assign n27547 = ~n27536 & ~n27546;
  assign n27548 = ~pi647 & ~n27547;
  assign n27549 = pi647 & ~n27499;
  assign n27550 = ~n27548 & ~n27549;
  assign n27551 = ~pi1157 & n27550;
  assign n27552 = pi647 & ~n27547;
  assign n27553 = ~pi647 & ~n27499;
  assign n27554 = ~n27552 & ~n27553;
  assign n27555 = pi1157 & n27554;
  assign n27556 = ~n27551 & ~n27555;
  assign n27557 = pi787 & ~n27556;
  assign n27558 = ~pi787 & n27547;
  assign n27559 = ~n27557 & ~n27558;
  assign n27560 = ~pi644 & ~n27559;
  assign n27561 = pi715 & ~n27560;
  assign n27562 = pi183 & ~n3267;
  assign n27563 = ~pi755 & n17282;
  assign n27564 = ~n27508 & ~n27563;
  assign n27565 = pi38 & ~n27564;
  assign n27566 = ~pi183 & n17242;
  assign n27567 = pi183 & ~n17275;
  assign n27568 = ~pi755 & ~n27567;
  assign n27569 = ~n27566 & n27568;
  assign n27570 = ~pi183 & pi755;
  assign n27571 = ~n17201 & n27570;
  assign n27572 = ~n27569 & ~n27571;
  assign n27573 = ~pi38 & ~n27572;
  assign n27574 = ~n27565 & ~n27573;
  assign n27575 = n3267 & n27574;
  assign n27576 = ~n27562 & ~n27575;
  assign n27577 = ~n17438 & ~n27576;
  assign n27578 = n17438 & ~n27499;
  assign n27579 = ~n27577 & ~n27578;
  assign n27580 = ~pi785 & ~n27579;
  assign n27581 = ~n17439 & ~n27499;
  assign n27582 = pi609 & n27577;
  assign n27583 = ~n27581 & ~n27582;
  assign n27584 = pi1155 & ~n27583;
  assign n27585 = ~n17451 & ~n27499;
  assign n27586 = ~pi609 & n27577;
  assign n27587 = ~n27585 & ~n27586;
  assign n27588 = ~pi1155 & ~n27587;
  assign n27589 = ~n27584 & ~n27588;
  assign n27590 = pi785 & ~n27589;
  assign n27591 = ~n27580 & ~n27590;
  assign n27592 = ~pi781 & ~n27591;
  assign n27593 = pi618 & n27591;
  assign n27594 = ~pi618 & n27499;
  assign n27595 = pi1154 & ~n27594;
  assign n27596 = ~n27593 & n27595;
  assign n27597 = ~pi618 & n27591;
  assign n27598 = pi618 & n27499;
  assign n27599 = ~pi1154 & ~n27598;
  assign n27600 = ~n27597 & n27599;
  assign n27601 = ~n27596 & ~n27600;
  assign n27602 = pi781 & ~n27601;
  assign n27603 = ~n27592 & ~n27602;
  assign n27604 = ~pi789 & ~n27603;
  assign n27605 = pi619 & n27603;
  assign n27606 = ~pi619 & n27499;
  assign n27607 = pi1159 & ~n27606;
  assign n27608 = ~n27605 & n27607;
  assign n27609 = ~pi619 & n27603;
  assign n27610 = pi619 & n27499;
  assign n27611 = ~pi1159 & ~n27610;
  assign n27612 = ~n27609 & n27611;
  assign n27613 = ~n27608 & ~n27612;
  assign n27614 = pi789 & ~n27613;
  assign n27615 = ~n27604 & ~n27614;
  assign n27616 = ~n17816 & n27615;
  assign n27617 = n17816 & n27499;
  assign n27618 = ~n27616 & ~n27617;
  assign n27619 = ~n17610 & ~n27618;
  assign n27620 = n17610 & n27499;
  assign n27621 = ~n27619 & ~n27620;
  assign n27622 = ~n17652 & ~n27621;
  assign n27623 = n17652 & n27499;
  assign n27624 = ~n27622 & ~n27623;
  assign n27625 = pi644 & ~n27624;
  assign n27626 = ~pi644 & n27499;
  assign n27627 = ~pi715 & ~n27626;
  assign n27628 = ~n27625 & n27627;
  assign n27629 = pi1160 & ~n27628;
  assign n27630 = ~n27561 & n27629;
  assign n27631 = pi644 & ~n27559;
  assign n27632 = ~pi715 & ~n27631;
  assign n27633 = ~pi644 & ~n27624;
  assign n27634 = pi644 & n27499;
  assign n27635 = pi715 & ~n27634;
  assign n27636 = ~n27633 & n27635;
  assign n27637 = ~pi1160 & ~n27636;
  assign n27638 = ~n27632 & n27637;
  assign n27639 = ~n27630 & ~n27638;
  assign n27640 = pi790 & ~n27639;
  assign n27641 = pi644 & n27629;
  assign n27642 = ~pi644 & n27637;
  assign n27643 = pi790 & ~n27642;
  assign n27644 = ~n27641 & n27643;
  assign n27645 = ~n20409 & n27618;
  assign n27646 = ~pi629 & n27540;
  assign n27647 = pi629 & n27544;
  assign n27648 = ~n27646 & ~n27647;
  assign n27649 = ~n27645 & n27648;
  assign n27650 = pi792 & ~n27649;
  assign n27651 = pi725 & ~n27574;
  assign n27652 = ~pi183 & n16687;
  assign n27653 = pi183 & n16799;
  assign n27654 = pi755 & ~n27653;
  assign n27655 = ~n27652 & n27654;
  assign n27656 = pi183 & n16879;
  assign n27657 = ~pi183 & ~n16944;
  assign n27658 = ~pi755 & ~n27657;
  assign n27659 = ~n27656 & n27658;
  assign n27660 = pi39 & ~n27659;
  assign n27661 = ~n27655 & n27660;
  assign n27662 = ~pi183 & ~n17088;
  assign n27663 = pi183 & ~n17059;
  assign n27664 = pi755 & ~n27663;
  assign n27665 = ~n27662 & n27664;
  assign n27666 = ~pi183 & n17092;
  assign n27667 = pi183 & n17094;
  assign n27668 = ~pi755 & ~n27667;
  assign n27669 = ~n27666 & n27668;
  assign n27670 = ~n27665 & ~n27669;
  assign n27671 = ~pi39 & ~n27670;
  assign n27672 = ~pi38 & ~n27671;
  assign n27673 = ~n27661 & n27672;
  assign n27674 = ~pi755 & ~n16905;
  assign n27675 = n19230 & ~n27674;
  assign n27676 = ~pi183 & ~n27675;
  assign n27677 = ~n16787 & ~n27314;
  assign n27678 = pi183 & ~n27677;
  assign n27679 = n6234 & n27678;
  assign n27680 = pi38 & ~n27679;
  assign n27681 = ~n27676 & n27680;
  assign n27682 = ~pi725 & ~n27681;
  assign n27683 = ~n27673 & n27682;
  assign n27684 = n3267 & ~n27683;
  assign n27685 = ~n27651 & n27684;
  assign n27686 = ~n27562 & ~n27685;
  assign n27687 = ~pi625 & n27686;
  assign n27688 = pi625 & n27576;
  assign n27689 = ~pi1153 & ~n27688;
  assign n27690 = ~n27687 & n27689;
  assign n27691 = ~pi608 & ~n27517;
  assign n27692 = ~n27690 & n27691;
  assign n27693 = pi625 & n27686;
  assign n27694 = ~pi625 & n27576;
  assign n27695 = pi1153 & ~n27694;
  assign n27696 = ~n27693 & n27695;
  assign n27697 = pi608 & ~n27521;
  assign n27698 = ~n27696 & n27697;
  assign n27699 = ~n27692 & ~n27698;
  assign n27700 = pi778 & ~n27699;
  assign n27701 = ~pi778 & n27686;
  assign n27702 = ~n27700 & ~n27701;
  assign n27703 = ~pi609 & ~n27702;
  assign n27704 = pi609 & n27524;
  assign n27705 = ~pi1155 & ~n27704;
  assign n27706 = ~n27703 & n27705;
  assign n27707 = ~pi660 & ~n27584;
  assign n27708 = ~n27706 & n27707;
  assign n27709 = pi609 & ~n27702;
  assign n27710 = ~pi609 & n27524;
  assign n27711 = pi1155 & ~n27710;
  assign n27712 = ~n27709 & n27711;
  assign n27713 = pi660 & ~n27588;
  assign n27714 = ~n27712 & n27713;
  assign n27715 = ~n27708 & ~n27714;
  assign n27716 = pi785 & ~n27715;
  assign n27717 = ~pi785 & ~n27702;
  assign n27718 = ~n27716 & ~n27717;
  assign n27719 = ~pi618 & ~n27718;
  assign n27720 = pi618 & n27527;
  assign n27721 = ~pi1154 & ~n27720;
  assign n27722 = ~n27719 & n27721;
  assign n27723 = ~pi627 & ~n27596;
  assign n27724 = ~n27722 & n27723;
  assign n27725 = pi618 & ~n27718;
  assign n27726 = ~pi618 & n27527;
  assign n27727 = pi1154 & ~n27726;
  assign n27728 = ~n27725 & n27727;
  assign n27729 = pi627 & ~n27600;
  assign n27730 = ~n27728 & n27729;
  assign n27731 = ~n27724 & ~n27730;
  assign n27732 = pi781 & ~n27731;
  assign n27733 = ~pi781 & ~n27718;
  assign n27734 = ~n27732 & ~n27733;
  assign n27735 = pi619 & ~n27734;
  assign n27736 = ~pi619 & ~n27530;
  assign n27737 = pi1159 & ~n27736;
  assign n27738 = ~n27735 & n27737;
  assign n27739 = pi648 & ~n27612;
  assign n27740 = ~n27738 & n27739;
  assign n27741 = ~pi619 & ~n27734;
  assign n27742 = pi619 & ~n27530;
  assign n27743 = ~pi1159 & ~n27742;
  assign n27744 = ~n27741 & n27743;
  assign n27745 = ~pi648 & ~n27608;
  assign n27746 = ~n27744 & n27745;
  assign n27747 = pi789 & ~n27746;
  assign n27748 = ~n27740 & n27747;
  assign n27749 = ~pi789 & n27734;
  assign n27750 = n17817 & ~n27749;
  assign n27751 = ~n27748 & n27750;
  assign n27752 = pi626 & ~n27615;
  assign n27753 = ~pi626 & ~n27499;
  assign n27754 = n17579 & ~n27753;
  assign n27755 = ~n27752 & n27754;
  assign n27756 = n17704 & n27532;
  assign n27757 = ~pi626 & ~n27615;
  assign n27758 = pi626 & ~n27499;
  assign n27759 = n17580 & ~n27758;
  assign n27760 = ~n27757 & n27759;
  assign n27761 = ~n27756 & ~n27760;
  assign n27762 = ~n27755 & n27761;
  assign n27763 = pi788 & ~n27762;
  assign n27764 = ~n20205 & ~n27763;
  assign n27765 = ~n27751 & n27764;
  assign n27766 = ~n27650 & ~n27765;
  assign n27767 = n20207 & ~n27766;
  assign n27768 = ~n20398 & n27621;
  assign n27769 = n17650 & ~n27550;
  assign n27770 = n17649 & ~n27554;
  assign n27771 = ~n27769 & ~n27770;
  assign n27772 = ~n27768 & n27771;
  assign n27773 = pi787 & ~n27772;
  assign n27774 = ~n27767 & ~n27773;
  assign n27775 = ~n27644 & n27774;
  assign n27776 = ~n27640 & ~n27775;
  assign n27777 = ~po1038 & ~n27776;
  assign n27778 = ~pi183 & po1038;
  assign n27779 = ~pi832 & ~n27778;
  assign n27780 = ~n27777 & n27779;
  assign po340 = ~n27498 & ~n27780;
  assign n27782 = ~pi184 & ~n2754;
  assign n27783 = ~pi777 & n16784;
  assign n27784 = ~n27782 & ~n27783;
  assign n27785 = ~n17706 & ~n27784;
  assign n27786 = ~pi785 & ~n27785;
  assign n27787 = n17451 & n27783;
  assign n27788 = n27785 & ~n27787;
  assign n27789 = pi1155 & ~n27788;
  assign n27790 = ~pi1155 & ~n27782;
  assign n27791 = ~n27787 & n27790;
  assign n27792 = ~n27789 & ~n27791;
  assign n27793 = pi785 & ~n27792;
  assign n27794 = ~n27786 & ~n27793;
  assign n27795 = ~pi781 & ~n27794;
  assign n27796 = ~n17721 & n27794;
  assign n27797 = pi1154 & ~n27796;
  assign n27798 = ~n17724 & n27794;
  assign n27799 = ~pi1154 & ~n27798;
  assign n27800 = ~n27797 & ~n27799;
  assign n27801 = pi781 & ~n27800;
  assign n27802 = ~n27795 & ~n27801;
  assign n27803 = ~pi789 & ~n27802;
  assign n27804 = ~n22890 & n27802;
  assign n27805 = pi1159 & ~n27804;
  assign n27806 = ~n22893 & n27802;
  assign n27807 = ~pi1159 & ~n27806;
  assign n27808 = ~n27805 & ~n27807;
  assign n27809 = pi789 & ~n27808;
  assign n27810 = ~n27803 & ~n27809;
  assign n27811 = ~n17816 & n27810;
  assign n27812 = n17816 & n27782;
  assign n27813 = ~n27811 & ~n27812;
  assign n27814 = ~n17610 & ~n27813;
  assign n27815 = n17610 & n27782;
  assign n27816 = ~n27814 & ~n27815;
  assign n27817 = ~n20398 & n27816;
  assign n27818 = ~pi737 & n16786;
  assign n27819 = ~n27782 & ~n27818;
  assign n27820 = ~pi778 & ~n27819;
  assign n27821 = ~pi625 & n27818;
  assign n27822 = ~n27819 & ~n27821;
  assign n27823 = pi1153 & ~n27822;
  assign n27824 = ~pi1153 & ~n27782;
  assign n27825 = ~n27821 & n27824;
  assign n27826 = pi778 & ~n27825;
  assign n27827 = ~n27823 & n27826;
  assign n27828 = ~n27820 & ~n27827;
  assign n27829 = ~n17692 & ~n27828;
  assign n27830 = ~n17694 & n27829;
  assign n27831 = ~n17696 & n27830;
  assign n27832 = ~n17828 & n27831;
  assign n27833 = ~n17859 & n27832;
  assign n27834 = ~pi647 & n27833;
  assign n27835 = pi647 & n27782;
  assign n27836 = ~pi1157 & ~n27835;
  assign n27837 = ~n27834 & n27836;
  assign n27838 = pi647 & ~n27833;
  assign n27839 = ~pi647 & ~n27782;
  assign n27840 = ~n27838 & ~n27839;
  assign n27841 = pi1157 & ~n27840;
  assign n27842 = ~n27837 & ~n27841;
  assign n27843 = ~n17651 & ~n27842;
  assign n27844 = ~n27817 & ~n27843;
  assign n27845 = pi787 & ~n27844;
  assign n27846 = pi626 & ~n27810;
  assign n27847 = ~pi626 & ~n27782;
  assign n27848 = n17579 & ~n27847;
  assign n27849 = ~n27846 & n27848;
  assign n27850 = n17704 & n27831;
  assign n27851 = ~pi626 & ~n27810;
  assign n27852 = pi626 & ~n27782;
  assign n27853 = n17580 & ~n27852;
  assign n27854 = ~n27851 & n27853;
  assign n27855 = ~n27850 & ~n27854;
  assign n27856 = ~n27849 & n27855;
  assign n27857 = pi788 & ~n27856;
  assign n27858 = ~n16521 & ~n27819;
  assign n27859 = pi625 & n27858;
  assign n27860 = n27784 & ~n27858;
  assign n27861 = ~n27859 & ~n27860;
  assign n27862 = n27824 & ~n27861;
  assign n27863 = ~pi608 & ~n27823;
  assign n27864 = ~n27862 & n27863;
  assign n27865 = pi1153 & n27784;
  assign n27866 = ~n27859 & n27865;
  assign n27867 = pi608 & ~n27825;
  assign n27868 = ~n27866 & n27867;
  assign n27869 = ~n27864 & ~n27868;
  assign n27870 = pi778 & ~n27869;
  assign n27871 = ~pi778 & ~n27860;
  assign n27872 = ~n27870 & ~n27871;
  assign n27873 = ~pi609 & ~n27872;
  assign n27874 = pi609 & ~n27828;
  assign n27875 = ~pi1155 & ~n27874;
  assign n27876 = ~n27873 & n27875;
  assign n27877 = ~pi660 & ~n27789;
  assign n27878 = ~n27876 & n27877;
  assign n27879 = pi609 & ~n27872;
  assign n27880 = ~pi609 & ~n27828;
  assign n27881 = pi1155 & ~n27880;
  assign n27882 = ~n27879 & n27881;
  assign n27883 = pi660 & ~n27791;
  assign n27884 = ~n27882 & n27883;
  assign n27885 = ~n27878 & ~n27884;
  assign n27886 = pi785 & ~n27885;
  assign n27887 = ~pi785 & ~n27872;
  assign n27888 = ~n27886 & ~n27887;
  assign n27889 = ~pi618 & ~n27888;
  assign n27890 = pi618 & n27829;
  assign n27891 = ~pi1154 & ~n27890;
  assign n27892 = ~n27889 & n27891;
  assign n27893 = ~pi627 & ~n27797;
  assign n27894 = ~n27892 & n27893;
  assign n27895 = pi618 & ~n27888;
  assign n27896 = ~pi618 & n27829;
  assign n27897 = pi1154 & ~n27896;
  assign n27898 = ~n27895 & n27897;
  assign n27899 = pi627 & ~n27799;
  assign n27900 = ~n27898 & n27899;
  assign n27901 = ~n27894 & ~n27900;
  assign n27902 = pi781 & ~n27901;
  assign n27903 = ~pi781 & ~n27888;
  assign n27904 = ~n27902 & ~n27903;
  assign n27905 = pi619 & ~n27904;
  assign n27906 = ~pi619 & n27830;
  assign n27907 = pi1159 & ~n27906;
  assign n27908 = ~n27905 & n27907;
  assign n27909 = pi648 & ~n27807;
  assign n27910 = ~n27908 & n27909;
  assign n27911 = ~pi619 & ~n27904;
  assign n27912 = pi619 & n27830;
  assign n27913 = ~pi1159 & ~n27912;
  assign n27914 = ~n27911 & n27913;
  assign n27915 = ~pi648 & ~n27805;
  assign n27916 = ~n27914 & n27915;
  assign n27917 = pi789 & ~n27916;
  assign n27918 = ~n27910 & n27917;
  assign n27919 = ~pi789 & n27904;
  assign n27920 = n17817 & ~n27919;
  assign n27921 = ~n27918 & n27920;
  assign n27922 = ~n27857 & ~n27921;
  assign n27923 = ~n20205 & ~n27922;
  assign n27924 = n17856 & ~n27813;
  assign n27925 = n20693 & n27832;
  assign n27926 = ~n27924 & ~n27925;
  assign n27927 = ~pi629 & ~n27926;
  assign n27928 = n20697 & n27832;
  assign n27929 = n17855 & ~n27813;
  assign n27930 = ~n27928 & ~n27929;
  assign n27931 = pi629 & ~n27930;
  assign n27932 = ~n27927 & ~n27931;
  assign n27933 = pi792 & ~n27932;
  assign n27934 = n20207 & ~n27933;
  assign n27935 = ~n27923 & n27934;
  assign n27936 = ~n27845 & ~n27935;
  assign n27937 = pi644 & n27936;
  assign n27938 = ~pi787 & ~n27833;
  assign n27939 = pi787 & ~n27842;
  assign n27940 = ~n27938 & ~n27939;
  assign n27941 = ~pi644 & n27940;
  assign n27942 = pi715 & ~n27941;
  assign n27943 = ~n27937 & n27942;
  assign n27944 = ~n17652 & ~n27816;
  assign n27945 = n17652 & n27782;
  assign n27946 = ~n27944 & ~n27945;
  assign n27947 = pi644 & ~n27946;
  assign n27948 = ~pi644 & n27782;
  assign n27949 = ~pi715 & ~n27948;
  assign n27950 = ~n27947 & n27949;
  assign n27951 = pi1160 & ~n27950;
  assign n27952 = ~n27943 & n27951;
  assign n27953 = ~pi644 & n27936;
  assign n27954 = pi644 & n27940;
  assign n27955 = ~pi715 & ~n27954;
  assign n27956 = ~n27953 & n27955;
  assign n27957 = ~pi644 & ~n27946;
  assign n27958 = pi644 & n27782;
  assign n27959 = pi715 & ~n27958;
  assign n27960 = ~n27957 & n27959;
  assign n27961 = ~pi1160 & ~n27960;
  assign n27962 = ~n27956 & n27961;
  assign n27963 = ~n27952 & ~n27962;
  assign n27964 = pi790 & ~n27963;
  assign n27965 = ~pi790 & n27936;
  assign n27966 = pi832 & ~n27965;
  assign n27967 = ~n27964 & n27966;
  assign n27968 = ~pi184 & ~n17406;
  assign n27969 = n17539 & ~n27968;
  assign n27970 = ~pi737 & n3267;
  assign n27971 = n27968 & ~n27970;
  assign n27972 = pi184 & ~n17976;
  assign n27973 = ~pi38 & ~n27972;
  assign n27974 = n3267 & ~n27973;
  assign n27975 = ~pi184 & n17972;
  assign n27976 = ~n27974 & ~n27975;
  assign n27977 = ~pi184 & ~n17280;
  assign n27978 = n17392 & ~n27977;
  assign n27979 = ~pi737 & ~n27978;
  assign n27980 = ~n27976 & n27979;
  assign n27981 = ~n27971 & ~n27980;
  assign n27982 = ~pi778 & n27981;
  assign n27983 = pi625 & ~n27981;
  assign n27984 = ~pi625 & n27968;
  assign n27985 = pi1153 & ~n27984;
  assign n27986 = ~n27983 & n27985;
  assign n27987 = ~pi625 & ~n27981;
  assign n27988 = pi625 & n27968;
  assign n27989 = ~pi1153 & ~n27988;
  assign n27990 = ~n27987 & n27989;
  assign n27991 = ~n27986 & ~n27990;
  assign n27992 = pi778 & ~n27991;
  assign n27993 = ~n27982 & ~n27992;
  assign n27994 = ~n17466 & ~n27993;
  assign n27995 = n17466 & ~n27968;
  assign n27996 = ~n27994 & ~n27995;
  assign n27997 = ~n17503 & n27996;
  assign n27998 = n17503 & n27968;
  assign n27999 = ~n27997 & ~n27998;
  assign n28000 = ~n17539 & n27999;
  assign n28001 = ~n27969 & ~n28000;
  assign n28002 = ~n17582 & n28001;
  assign n28003 = n17582 & n27968;
  assign n28004 = ~n28002 & ~n28003;
  assign n28005 = ~pi792 & n28004;
  assign n28006 = pi628 & ~n28004;
  assign n28007 = ~pi628 & n27968;
  assign n28008 = pi1156 & ~n28007;
  assign n28009 = ~n28006 & n28008;
  assign n28010 = ~pi628 & ~n28004;
  assign n28011 = pi628 & n27968;
  assign n28012 = ~pi1156 & ~n28011;
  assign n28013 = ~n28010 & n28012;
  assign n28014 = ~n28009 & ~n28013;
  assign n28015 = pi792 & ~n28014;
  assign n28016 = ~n28005 & ~n28015;
  assign n28017 = ~pi647 & ~n28016;
  assign n28018 = pi647 & ~n27968;
  assign n28019 = ~n28017 & ~n28018;
  assign n28020 = ~pi1157 & n28019;
  assign n28021 = pi647 & ~n28016;
  assign n28022 = ~pi647 & ~n27968;
  assign n28023 = ~n28021 & ~n28022;
  assign n28024 = pi1157 & n28023;
  assign n28025 = ~n28020 & ~n28024;
  assign n28026 = pi787 & ~n28025;
  assign n28027 = ~pi787 & n28016;
  assign n28028 = ~n28026 & ~n28027;
  assign n28029 = ~pi644 & ~n28028;
  assign n28030 = pi715 & ~n28029;
  assign n28031 = pi184 & ~n3267;
  assign n28032 = ~pi777 & n17282;
  assign n28033 = ~n27977 & ~n28032;
  assign n28034 = pi38 & ~n28033;
  assign n28035 = ~pi184 & n17242;
  assign n28036 = pi184 & ~n17275;
  assign n28037 = ~pi777 & ~n28036;
  assign n28038 = ~n28035 & n28037;
  assign n28039 = ~pi184 & pi777;
  assign n28040 = ~n17201 & n28039;
  assign n28041 = ~n28038 & ~n28040;
  assign n28042 = ~pi38 & ~n28041;
  assign n28043 = ~n28034 & ~n28042;
  assign n28044 = n3267 & n28043;
  assign n28045 = ~n28031 & ~n28044;
  assign n28046 = ~n17438 & ~n28045;
  assign n28047 = n17438 & ~n27968;
  assign n28048 = ~n28046 & ~n28047;
  assign n28049 = ~pi785 & ~n28048;
  assign n28050 = ~n17439 & ~n27968;
  assign n28051 = pi609 & n28046;
  assign n28052 = ~n28050 & ~n28051;
  assign n28053 = pi1155 & ~n28052;
  assign n28054 = ~n17451 & ~n27968;
  assign n28055 = ~pi609 & n28046;
  assign n28056 = ~n28054 & ~n28055;
  assign n28057 = ~pi1155 & ~n28056;
  assign n28058 = ~n28053 & ~n28057;
  assign n28059 = pi785 & ~n28058;
  assign n28060 = ~n28049 & ~n28059;
  assign n28061 = ~pi781 & ~n28060;
  assign n28062 = pi618 & n28060;
  assign n28063 = ~pi618 & n27968;
  assign n28064 = pi1154 & ~n28063;
  assign n28065 = ~n28062 & n28064;
  assign n28066 = ~pi618 & n28060;
  assign n28067 = pi618 & n27968;
  assign n28068 = ~pi1154 & ~n28067;
  assign n28069 = ~n28066 & n28068;
  assign n28070 = ~n28065 & ~n28069;
  assign n28071 = pi781 & ~n28070;
  assign n28072 = ~n28061 & ~n28071;
  assign n28073 = ~pi789 & ~n28072;
  assign n28074 = pi619 & n28072;
  assign n28075 = ~pi619 & n27968;
  assign n28076 = pi1159 & ~n28075;
  assign n28077 = ~n28074 & n28076;
  assign n28078 = ~pi619 & n28072;
  assign n28079 = pi619 & n27968;
  assign n28080 = ~pi1159 & ~n28079;
  assign n28081 = ~n28078 & n28080;
  assign n28082 = ~n28077 & ~n28081;
  assign n28083 = pi789 & ~n28082;
  assign n28084 = ~n28073 & ~n28083;
  assign n28085 = ~n17816 & n28084;
  assign n28086 = n17816 & n27968;
  assign n28087 = ~n28085 & ~n28086;
  assign n28088 = ~n17610 & ~n28087;
  assign n28089 = n17610 & n27968;
  assign n28090 = ~n28088 & ~n28089;
  assign n28091 = ~n17652 & ~n28090;
  assign n28092 = n17652 & n27968;
  assign n28093 = ~n28091 & ~n28092;
  assign n28094 = pi644 & ~n28093;
  assign n28095 = ~pi644 & n27968;
  assign n28096 = ~pi715 & ~n28095;
  assign n28097 = ~n28094 & n28096;
  assign n28098 = pi1160 & ~n28097;
  assign n28099 = ~n28030 & n28098;
  assign n28100 = pi644 & ~n28028;
  assign n28101 = ~pi715 & ~n28100;
  assign n28102 = ~pi644 & ~n28093;
  assign n28103 = pi644 & n27968;
  assign n28104 = pi715 & ~n28103;
  assign n28105 = ~n28102 & n28104;
  assign n28106 = ~pi1160 & ~n28105;
  assign n28107 = ~n28101 & n28106;
  assign n28108 = ~n28099 & ~n28107;
  assign n28109 = pi790 & ~n28108;
  assign n28110 = pi644 & n28098;
  assign n28111 = ~pi644 & n28106;
  assign n28112 = pi790 & ~n28111;
  assign n28113 = ~n28110 & n28112;
  assign n28114 = ~n20409 & n28087;
  assign n28115 = ~pi629 & n28009;
  assign n28116 = pi629 & n28013;
  assign n28117 = ~n28115 & ~n28116;
  assign n28118 = ~n28114 & n28117;
  assign n28119 = pi792 & ~n28118;
  assign n28120 = pi737 & ~n28043;
  assign n28121 = ~pi184 & n16687;
  assign n28122 = pi184 & n16799;
  assign n28123 = pi777 & ~n28122;
  assign n28124 = ~n28121 & n28123;
  assign n28125 = pi184 & n16879;
  assign n28126 = ~pi184 & ~n16944;
  assign n28127 = ~pi777 & ~n28126;
  assign n28128 = ~n28125 & n28127;
  assign n28129 = pi39 & ~n28128;
  assign n28130 = ~n28124 & n28129;
  assign n28131 = ~pi184 & ~n17088;
  assign n28132 = pi184 & ~n17059;
  assign n28133 = pi777 & ~n28132;
  assign n28134 = ~n28131 & n28133;
  assign n28135 = ~pi184 & n17092;
  assign n28136 = pi184 & n17094;
  assign n28137 = ~pi777 & ~n28136;
  assign n28138 = ~n28135 & n28137;
  assign n28139 = ~n28134 & ~n28138;
  assign n28140 = ~pi39 & ~n28139;
  assign n28141 = ~pi38 & ~n28140;
  assign n28142 = ~n28130 & n28141;
  assign n28143 = ~pi777 & ~n16905;
  assign n28144 = n19230 & ~n28143;
  assign n28145 = ~pi184 & ~n28144;
  assign n28146 = ~n16787 & ~n27783;
  assign n28147 = pi184 & ~n28146;
  assign n28148 = n6234 & n28147;
  assign n28149 = pi38 & ~n28148;
  assign n28150 = ~n28145 & n28149;
  assign n28151 = ~pi737 & ~n28150;
  assign n28152 = ~n28142 & n28151;
  assign n28153 = n3267 & ~n28152;
  assign n28154 = ~n28120 & n28153;
  assign n28155 = ~n28031 & ~n28154;
  assign n28156 = ~pi625 & n28155;
  assign n28157 = pi625 & n28045;
  assign n28158 = ~pi1153 & ~n28157;
  assign n28159 = ~n28156 & n28158;
  assign n28160 = ~pi608 & ~n27986;
  assign n28161 = ~n28159 & n28160;
  assign n28162 = pi625 & n28155;
  assign n28163 = ~pi625 & n28045;
  assign n28164 = pi1153 & ~n28163;
  assign n28165 = ~n28162 & n28164;
  assign n28166 = pi608 & ~n27990;
  assign n28167 = ~n28165 & n28166;
  assign n28168 = ~n28161 & ~n28167;
  assign n28169 = pi778 & ~n28168;
  assign n28170 = ~pi778 & n28155;
  assign n28171 = ~n28169 & ~n28170;
  assign n28172 = ~pi609 & ~n28171;
  assign n28173 = pi609 & n27993;
  assign n28174 = ~pi1155 & ~n28173;
  assign n28175 = ~n28172 & n28174;
  assign n28176 = ~pi660 & ~n28053;
  assign n28177 = ~n28175 & n28176;
  assign n28178 = pi609 & ~n28171;
  assign n28179 = ~pi609 & n27993;
  assign n28180 = pi1155 & ~n28179;
  assign n28181 = ~n28178 & n28180;
  assign n28182 = pi660 & ~n28057;
  assign n28183 = ~n28181 & n28182;
  assign n28184 = ~n28177 & ~n28183;
  assign n28185 = pi785 & ~n28184;
  assign n28186 = ~pi785 & ~n28171;
  assign n28187 = ~n28185 & ~n28186;
  assign n28188 = ~pi618 & ~n28187;
  assign n28189 = pi618 & n27996;
  assign n28190 = ~pi1154 & ~n28189;
  assign n28191 = ~n28188 & n28190;
  assign n28192 = ~pi627 & ~n28065;
  assign n28193 = ~n28191 & n28192;
  assign n28194 = pi618 & ~n28187;
  assign n28195 = ~pi618 & n27996;
  assign n28196 = pi1154 & ~n28195;
  assign n28197 = ~n28194 & n28196;
  assign n28198 = pi627 & ~n28069;
  assign n28199 = ~n28197 & n28198;
  assign n28200 = ~n28193 & ~n28199;
  assign n28201 = pi781 & ~n28200;
  assign n28202 = ~pi781 & ~n28187;
  assign n28203 = ~n28201 & ~n28202;
  assign n28204 = pi619 & ~n28203;
  assign n28205 = ~pi619 & ~n27999;
  assign n28206 = pi1159 & ~n28205;
  assign n28207 = ~n28204 & n28206;
  assign n28208 = pi648 & ~n28081;
  assign n28209 = ~n28207 & n28208;
  assign n28210 = ~pi619 & ~n28203;
  assign n28211 = pi619 & ~n27999;
  assign n28212 = ~pi1159 & ~n28211;
  assign n28213 = ~n28210 & n28212;
  assign n28214 = ~pi648 & ~n28077;
  assign n28215 = ~n28213 & n28214;
  assign n28216 = pi789 & ~n28215;
  assign n28217 = ~n28209 & n28216;
  assign n28218 = ~pi789 & n28203;
  assign n28219 = n17817 & ~n28218;
  assign n28220 = ~n28217 & n28219;
  assign n28221 = pi626 & ~n28084;
  assign n28222 = ~pi626 & ~n27968;
  assign n28223 = n17579 & ~n28222;
  assign n28224 = ~n28221 & n28223;
  assign n28225 = n17704 & n28001;
  assign n28226 = ~pi626 & ~n28084;
  assign n28227 = pi626 & ~n27968;
  assign n28228 = n17580 & ~n28227;
  assign n28229 = ~n28226 & n28228;
  assign n28230 = ~n28225 & ~n28229;
  assign n28231 = ~n28224 & n28230;
  assign n28232 = pi788 & ~n28231;
  assign n28233 = ~n20205 & ~n28232;
  assign n28234 = ~n28220 & n28233;
  assign n28235 = ~n28119 & ~n28234;
  assign n28236 = n20207 & ~n28235;
  assign n28237 = ~n20398 & n28090;
  assign n28238 = n17650 & ~n28019;
  assign n28239 = n17649 & ~n28023;
  assign n28240 = ~n28238 & ~n28239;
  assign n28241 = ~n28237 & n28240;
  assign n28242 = pi787 & ~n28241;
  assign n28243 = ~n28236 & ~n28242;
  assign n28244 = ~n28113 & n28243;
  assign n28245 = ~n28109 & ~n28244;
  assign n28246 = ~po1038 & ~n28245;
  assign n28247 = ~pi184 & po1038;
  assign n28248 = ~pi832 & ~n28247;
  assign n28249 = ~n28246 & n28248;
  assign po341 = ~n27967 & ~n28249;
  assign n28251 = ~pi185 & ~n2754;
  assign n28252 = ~pi751 & n16784;
  assign n28253 = ~n28251 & ~n28252;
  assign n28254 = ~n17706 & ~n28253;
  assign n28255 = ~pi785 & ~n28254;
  assign n28256 = n17451 & n28252;
  assign n28257 = n28254 & ~n28256;
  assign n28258 = pi1155 & ~n28257;
  assign n28259 = ~pi1155 & ~n28251;
  assign n28260 = ~n28256 & n28259;
  assign n28261 = ~n28258 & ~n28260;
  assign n28262 = pi785 & ~n28261;
  assign n28263 = ~n28255 & ~n28262;
  assign n28264 = ~pi781 & ~n28263;
  assign n28265 = ~n17721 & n28263;
  assign n28266 = pi1154 & ~n28265;
  assign n28267 = ~n17724 & n28263;
  assign n28268 = ~pi1154 & ~n28267;
  assign n28269 = ~n28266 & ~n28268;
  assign n28270 = pi781 & ~n28269;
  assign n28271 = ~n28264 & ~n28270;
  assign n28272 = ~pi789 & ~n28271;
  assign n28273 = ~n22890 & n28271;
  assign n28274 = pi1159 & ~n28273;
  assign n28275 = ~n22893 & n28271;
  assign n28276 = ~pi1159 & ~n28275;
  assign n28277 = ~n28274 & ~n28276;
  assign n28278 = pi789 & ~n28277;
  assign n28279 = ~n28272 & ~n28278;
  assign n28280 = ~n17816 & n28279;
  assign n28281 = n17816 & n28251;
  assign n28282 = ~n28280 & ~n28281;
  assign n28283 = ~n17610 & ~n28282;
  assign n28284 = n17610 & n28251;
  assign n28285 = ~n28283 & ~n28284;
  assign n28286 = ~n20398 & n28285;
  assign n28287 = ~pi701 & n16786;
  assign n28288 = ~n28251 & ~n28287;
  assign n28289 = ~pi778 & ~n28288;
  assign n28290 = ~pi625 & n28287;
  assign n28291 = ~n28288 & ~n28290;
  assign n28292 = pi1153 & ~n28291;
  assign n28293 = ~pi1153 & ~n28251;
  assign n28294 = ~n28290 & n28293;
  assign n28295 = pi778 & ~n28294;
  assign n28296 = ~n28292 & n28295;
  assign n28297 = ~n28289 & ~n28296;
  assign n28298 = ~n17692 & ~n28297;
  assign n28299 = ~n17694 & n28298;
  assign n28300 = ~n17696 & n28299;
  assign n28301 = ~n17828 & n28300;
  assign n28302 = ~n17859 & n28301;
  assign n28303 = ~pi647 & n28302;
  assign n28304 = pi647 & n28251;
  assign n28305 = ~pi1157 & ~n28304;
  assign n28306 = ~n28303 & n28305;
  assign n28307 = pi647 & ~n28302;
  assign n28308 = ~pi647 & ~n28251;
  assign n28309 = ~n28307 & ~n28308;
  assign n28310 = pi1157 & ~n28309;
  assign n28311 = ~n28306 & ~n28310;
  assign n28312 = ~n17651 & ~n28311;
  assign n28313 = ~n28286 & ~n28312;
  assign n28314 = pi787 & ~n28313;
  assign n28315 = pi626 & ~n28279;
  assign n28316 = ~pi626 & ~n28251;
  assign n28317 = n17579 & ~n28316;
  assign n28318 = ~n28315 & n28317;
  assign n28319 = n17704 & n28300;
  assign n28320 = ~pi626 & ~n28279;
  assign n28321 = pi626 & ~n28251;
  assign n28322 = n17580 & ~n28321;
  assign n28323 = ~n28320 & n28322;
  assign n28324 = ~n28319 & ~n28323;
  assign n28325 = ~n28318 & n28324;
  assign n28326 = pi788 & ~n28325;
  assign n28327 = ~n16521 & ~n28288;
  assign n28328 = pi625 & n28327;
  assign n28329 = n28253 & ~n28327;
  assign n28330 = ~n28328 & ~n28329;
  assign n28331 = n28293 & ~n28330;
  assign n28332 = ~pi608 & ~n28292;
  assign n28333 = ~n28331 & n28332;
  assign n28334 = pi1153 & n28253;
  assign n28335 = ~n28328 & n28334;
  assign n28336 = pi608 & ~n28294;
  assign n28337 = ~n28335 & n28336;
  assign n28338 = ~n28333 & ~n28337;
  assign n28339 = pi778 & ~n28338;
  assign n28340 = ~pi778 & ~n28329;
  assign n28341 = ~n28339 & ~n28340;
  assign n28342 = ~pi609 & ~n28341;
  assign n28343 = pi609 & ~n28297;
  assign n28344 = ~pi1155 & ~n28343;
  assign n28345 = ~n28342 & n28344;
  assign n28346 = ~pi660 & ~n28258;
  assign n28347 = ~n28345 & n28346;
  assign n28348 = pi609 & ~n28341;
  assign n28349 = ~pi609 & ~n28297;
  assign n28350 = pi1155 & ~n28349;
  assign n28351 = ~n28348 & n28350;
  assign n28352 = pi660 & ~n28260;
  assign n28353 = ~n28351 & n28352;
  assign n28354 = ~n28347 & ~n28353;
  assign n28355 = pi785 & ~n28354;
  assign n28356 = ~pi785 & ~n28341;
  assign n28357 = ~n28355 & ~n28356;
  assign n28358 = ~pi618 & ~n28357;
  assign n28359 = pi618 & n28298;
  assign n28360 = ~pi1154 & ~n28359;
  assign n28361 = ~n28358 & n28360;
  assign n28362 = ~pi627 & ~n28266;
  assign n28363 = ~n28361 & n28362;
  assign n28364 = pi618 & ~n28357;
  assign n28365 = ~pi618 & n28298;
  assign n28366 = pi1154 & ~n28365;
  assign n28367 = ~n28364 & n28366;
  assign n28368 = pi627 & ~n28268;
  assign n28369 = ~n28367 & n28368;
  assign n28370 = ~n28363 & ~n28369;
  assign n28371 = pi781 & ~n28370;
  assign n28372 = ~pi781 & ~n28357;
  assign n28373 = ~n28371 & ~n28372;
  assign n28374 = pi619 & ~n28373;
  assign n28375 = ~pi619 & n28299;
  assign n28376 = pi1159 & ~n28375;
  assign n28377 = ~n28374 & n28376;
  assign n28378 = pi648 & ~n28276;
  assign n28379 = ~n28377 & n28378;
  assign n28380 = ~pi619 & ~n28373;
  assign n28381 = pi619 & n28299;
  assign n28382 = ~pi1159 & ~n28381;
  assign n28383 = ~n28380 & n28382;
  assign n28384 = ~pi648 & ~n28274;
  assign n28385 = ~n28383 & n28384;
  assign n28386 = pi789 & ~n28385;
  assign n28387 = ~n28379 & n28386;
  assign n28388 = ~pi789 & n28373;
  assign n28389 = n17817 & ~n28388;
  assign n28390 = ~n28387 & n28389;
  assign n28391 = ~n28326 & ~n28390;
  assign n28392 = ~n20205 & ~n28391;
  assign n28393 = n17856 & ~n28282;
  assign n28394 = n20693 & n28301;
  assign n28395 = ~n28393 & ~n28394;
  assign n28396 = ~pi629 & ~n28395;
  assign n28397 = n20697 & n28301;
  assign n28398 = n17855 & ~n28282;
  assign n28399 = ~n28397 & ~n28398;
  assign n28400 = pi629 & ~n28399;
  assign n28401 = ~n28396 & ~n28400;
  assign n28402 = pi792 & ~n28401;
  assign n28403 = n20207 & ~n28402;
  assign n28404 = ~n28392 & n28403;
  assign n28405 = ~n28314 & ~n28404;
  assign n28406 = pi644 & n28405;
  assign n28407 = ~pi787 & ~n28302;
  assign n28408 = pi787 & ~n28311;
  assign n28409 = ~n28407 & ~n28408;
  assign n28410 = ~pi644 & n28409;
  assign n28411 = pi715 & ~n28410;
  assign n28412 = ~n28406 & n28411;
  assign n28413 = ~n17652 & ~n28285;
  assign n28414 = n17652 & n28251;
  assign n28415 = ~n28413 & ~n28414;
  assign n28416 = pi644 & ~n28415;
  assign n28417 = ~pi644 & n28251;
  assign n28418 = ~pi715 & ~n28417;
  assign n28419 = ~n28416 & n28418;
  assign n28420 = pi1160 & ~n28419;
  assign n28421 = ~n28412 & n28420;
  assign n28422 = ~pi644 & n28405;
  assign n28423 = pi644 & n28409;
  assign n28424 = ~pi715 & ~n28423;
  assign n28425 = ~n28422 & n28424;
  assign n28426 = ~pi644 & ~n28415;
  assign n28427 = pi644 & n28251;
  assign n28428 = pi715 & ~n28427;
  assign n28429 = ~n28426 & n28428;
  assign n28430 = ~pi1160 & ~n28429;
  assign n28431 = ~n28425 & n28430;
  assign n28432 = ~n28421 & ~n28431;
  assign n28433 = pi790 & ~n28432;
  assign n28434 = ~pi790 & n28405;
  assign n28435 = pi832 & ~n28434;
  assign n28436 = ~n28433 & n28435;
  assign n28437 = ~pi185 & ~n17406;
  assign n28438 = n17539 & ~n28437;
  assign n28439 = ~pi701 & n3267;
  assign n28440 = n28437 & ~n28439;
  assign n28441 = pi185 & ~n17976;
  assign n28442 = ~pi38 & ~n28441;
  assign n28443 = n3267 & ~n28442;
  assign n28444 = ~pi185 & n17972;
  assign n28445 = ~n28443 & ~n28444;
  assign n28446 = ~pi185 & ~n17280;
  assign n28447 = n17392 & ~n28446;
  assign n28448 = ~pi701 & ~n28447;
  assign n28449 = ~n28445 & n28448;
  assign n28450 = ~n28440 & ~n28449;
  assign n28451 = ~pi778 & n28450;
  assign n28452 = pi625 & ~n28450;
  assign n28453 = ~pi625 & n28437;
  assign n28454 = pi1153 & ~n28453;
  assign n28455 = ~n28452 & n28454;
  assign n28456 = ~pi625 & ~n28450;
  assign n28457 = pi625 & n28437;
  assign n28458 = ~pi1153 & ~n28457;
  assign n28459 = ~n28456 & n28458;
  assign n28460 = ~n28455 & ~n28459;
  assign n28461 = pi778 & ~n28460;
  assign n28462 = ~n28451 & ~n28461;
  assign n28463 = ~n17466 & ~n28462;
  assign n28464 = n17466 & ~n28437;
  assign n28465 = ~n28463 & ~n28464;
  assign n28466 = ~n17503 & n28465;
  assign n28467 = n17503 & n28437;
  assign n28468 = ~n28466 & ~n28467;
  assign n28469 = ~n17539 & n28468;
  assign n28470 = ~n28438 & ~n28469;
  assign n28471 = ~n17582 & n28470;
  assign n28472 = n17582 & n28437;
  assign n28473 = ~n28471 & ~n28472;
  assign n28474 = ~pi792 & n28473;
  assign n28475 = pi628 & ~n28473;
  assign n28476 = ~pi628 & n28437;
  assign n28477 = pi1156 & ~n28476;
  assign n28478 = ~n28475 & n28477;
  assign n28479 = ~pi628 & ~n28473;
  assign n28480 = pi628 & n28437;
  assign n28481 = ~pi1156 & ~n28480;
  assign n28482 = ~n28479 & n28481;
  assign n28483 = ~n28478 & ~n28482;
  assign n28484 = pi792 & ~n28483;
  assign n28485 = ~n28474 & ~n28484;
  assign n28486 = ~pi647 & ~n28485;
  assign n28487 = pi647 & ~n28437;
  assign n28488 = ~n28486 & ~n28487;
  assign n28489 = ~pi1157 & n28488;
  assign n28490 = pi647 & ~n28485;
  assign n28491 = ~pi647 & ~n28437;
  assign n28492 = ~n28490 & ~n28491;
  assign n28493 = pi1157 & n28492;
  assign n28494 = ~n28489 & ~n28493;
  assign n28495 = pi787 & ~n28494;
  assign n28496 = ~pi787 & n28485;
  assign n28497 = ~n28495 & ~n28496;
  assign n28498 = ~pi644 & ~n28497;
  assign n28499 = pi715 & ~n28498;
  assign n28500 = pi185 & ~n3267;
  assign n28501 = pi751 & n17199;
  assign n28502 = pi185 & n17273;
  assign n28503 = ~n28501 & ~n28502;
  assign n28504 = pi39 & ~n28503;
  assign n28505 = ~pi185 & ~pi751;
  assign n28506 = n17242 & n28505;
  assign n28507 = pi185 & pi751;
  assign n28508 = pi185 & ~n17086;
  assign n28509 = ~n21091 & ~n28508;
  assign n28510 = ~pi39 & ~n28509;
  assign n28511 = ~n28507 & ~n28510;
  assign n28512 = ~n28506 & n28511;
  assign n28513 = ~n28504 & n28512;
  assign n28514 = ~pi38 & ~n28513;
  assign n28515 = ~pi751 & n17282;
  assign n28516 = pi38 & ~n28446;
  assign n28517 = ~n28515 & n28516;
  assign n28518 = ~n28514 & ~n28517;
  assign n28519 = n3267 & ~n28518;
  assign n28520 = ~n28500 & ~n28519;
  assign n28521 = ~n17438 & ~n28520;
  assign n28522 = n17438 & ~n28437;
  assign n28523 = ~n28521 & ~n28522;
  assign n28524 = ~pi785 & ~n28523;
  assign n28525 = ~n17439 & ~n28437;
  assign n28526 = pi609 & n28521;
  assign n28527 = ~n28525 & ~n28526;
  assign n28528 = pi1155 & ~n28527;
  assign n28529 = ~n17451 & ~n28437;
  assign n28530 = ~pi609 & n28521;
  assign n28531 = ~n28529 & ~n28530;
  assign n28532 = ~pi1155 & ~n28531;
  assign n28533 = ~n28528 & ~n28532;
  assign n28534 = pi785 & ~n28533;
  assign n28535 = ~n28524 & ~n28534;
  assign n28536 = ~pi781 & ~n28535;
  assign n28537 = pi618 & n28535;
  assign n28538 = ~pi618 & n28437;
  assign n28539 = pi1154 & ~n28538;
  assign n28540 = ~n28537 & n28539;
  assign n28541 = ~pi618 & n28535;
  assign n28542 = pi618 & n28437;
  assign n28543 = ~pi1154 & ~n28542;
  assign n28544 = ~n28541 & n28543;
  assign n28545 = ~n28540 & ~n28544;
  assign n28546 = pi781 & ~n28545;
  assign n28547 = ~n28536 & ~n28546;
  assign n28548 = ~pi789 & ~n28547;
  assign n28549 = pi619 & n28547;
  assign n28550 = ~pi619 & n28437;
  assign n28551 = pi1159 & ~n28550;
  assign n28552 = ~n28549 & n28551;
  assign n28553 = ~pi619 & n28547;
  assign n28554 = pi619 & n28437;
  assign n28555 = ~pi1159 & ~n28554;
  assign n28556 = ~n28553 & n28555;
  assign n28557 = ~n28552 & ~n28556;
  assign n28558 = pi789 & ~n28557;
  assign n28559 = ~n28548 & ~n28558;
  assign n28560 = ~n17816 & n28559;
  assign n28561 = n17816 & n28437;
  assign n28562 = ~n28560 & ~n28561;
  assign n28563 = ~n17610 & ~n28562;
  assign n28564 = n17610 & n28437;
  assign n28565 = ~n28563 & ~n28564;
  assign n28566 = ~n17652 & ~n28565;
  assign n28567 = n17652 & n28437;
  assign n28568 = ~n28566 & ~n28567;
  assign n28569 = pi644 & ~n28568;
  assign n28570 = ~pi644 & n28437;
  assign n28571 = ~pi715 & ~n28570;
  assign n28572 = ~n28569 & n28571;
  assign n28573 = pi1160 & ~n28572;
  assign n28574 = ~n28499 & n28573;
  assign n28575 = pi644 & ~n28497;
  assign n28576 = ~pi715 & ~n28575;
  assign n28577 = ~pi644 & ~n28568;
  assign n28578 = pi644 & n28437;
  assign n28579 = pi715 & ~n28578;
  assign n28580 = ~n28577 & n28579;
  assign n28581 = ~pi1160 & ~n28580;
  assign n28582 = ~n28576 & n28581;
  assign n28583 = ~n28574 & ~n28582;
  assign n28584 = pi790 & ~n28583;
  assign n28585 = pi644 & n28573;
  assign n28586 = ~pi644 & n28581;
  assign n28587 = pi790 & ~n28586;
  assign n28588 = ~n28585 & n28587;
  assign n28589 = ~n20409 & n28562;
  assign n28590 = ~pi629 & n28478;
  assign n28591 = pi629 & n28482;
  assign n28592 = ~n28590 & ~n28591;
  assign n28593 = ~n28589 & n28592;
  assign n28594 = pi792 & ~n28593;
  assign n28595 = pi701 & n28518;
  assign n28596 = ~pi185 & n16687;
  assign n28597 = pi185 & n16799;
  assign n28598 = pi751 & ~n28597;
  assign n28599 = ~n28596 & n28598;
  assign n28600 = pi185 & n16879;
  assign n28601 = ~pi185 & ~n16944;
  assign n28602 = ~pi751 & ~n28601;
  assign n28603 = ~n28600 & n28602;
  assign n28604 = pi39 & ~n28603;
  assign n28605 = ~n28599 & n28604;
  assign n28606 = ~pi185 & ~n17088;
  assign n28607 = pi185 & ~n17059;
  assign n28608 = pi751 & ~n28607;
  assign n28609 = ~n28606 & n28608;
  assign n28610 = ~pi185 & n17092;
  assign n28611 = pi185 & n17094;
  assign n28612 = ~pi751 & ~n28611;
  assign n28613 = ~n28610 & n28612;
  assign n28614 = ~n28609 & ~n28613;
  assign n28615 = ~pi39 & ~n28614;
  assign n28616 = ~pi38 & ~n28615;
  assign n28617 = ~n28605 & n28616;
  assign n28618 = ~pi751 & ~n16905;
  assign n28619 = n19230 & ~n28618;
  assign n28620 = ~pi185 & ~n28619;
  assign n28621 = ~n16787 & ~n28252;
  assign n28622 = pi185 & ~n28621;
  assign n28623 = n6234 & n28622;
  assign n28624 = pi38 & ~n28623;
  assign n28625 = ~n28620 & n28624;
  assign n28626 = ~pi701 & ~n28625;
  assign n28627 = ~n28617 & n28626;
  assign n28628 = n3267 & ~n28627;
  assign n28629 = ~n28595 & n28628;
  assign n28630 = ~n28500 & ~n28629;
  assign n28631 = ~pi625 & n28630;
  assign n28632 = pi625 & n28520;
  assign n28633 = ~pi1153 & ~n28632;
  assign n28634 = ~n28631 & n28633;
  assign n28635 = ~pi608 & ~n28455;
  assign n28636 = ~n28634 & n28635;
  assign n28637 = pi625 & n28630;
  assign n28638 = ~pi625 & n28520;
  assign n28639 = pi1153 & ~n28638;
  assign n28640 = ~n28637 & n28639;
  assign n28641 = pi608 & ~n28459;
  assign n28642 = ~n28640 & n28641;
  assign n28643 = ~n28636 & ~n28642;
  assign n28644 = pi778 & ~n28643;
  assign n28645 = ~pi778 & n28630;
  assign n28646 = ~n28644 & ~n28645;
  assign n28647 = ~pi609 & ~n28646;
  assign n28648 = pi609 & n28462;
  assign n28649 = ~pi1155 & ~n28648;
  assign n28650 = ~n28647 & n28649;
  assign n28651 = ~pi660 & ~n28528;
  assign n28652 = ~n28650 & n28651;
  assign n28653 = pi609 & ~n28646;
  assign n28654 = ~pi609 & n28462;
  assign n28655 = pi1155 & ~n28654;
  assign n28656 = ~n28653 & n28655;
  assign n28657 = pi660 & ~n28532;
  assign n28658 = ~n28656 & n28657;
  assign n28659 = ~n28652 & ~n28658;
  assign n28660 = pi785 & ~n28659;
  assign n28661 = ~pi785 & ~n28646;
  assign n28662 = ~n28660 & ~n28661;
  assign n28663 = ~pi618 & ~n28662;
  assign n28664 = pi618 & n28465;
  assign n28665 = ~pi1154 & ~n28664;
  assign n28666 = ~n28663 & n28665;
  assign n28667 = ~pi627 & ~n28540;
  assign n28668 = ~n28666 & n28667;
  assign n28669 = pi618 & ~n28662;
  assign n28670 = ~pi618 & n28465;
  assign n28671 = pi1154 & ~n28670;
  assign n28672 = ~n28669 & n28671;
  assign n28673 = pi627 & ~n28544;
  assign n28674 = ~n28672 & n28673;
  assign n28675 = ~n28668 & ~n28674;
  assign n28676 = pi781 & ~n28675;
  assign n28677 = ~pi781 & ~n28662;
  assign n28678 = ~n28676 & ~n28677;
  assign n28679 = pi619 & ~n28678;
  assign n28680 = ~pi619 & ~n28468;
  assign n28681 = pi1159 & ~n28680;
  assign n28682 = ~n28679 & n28681;
  assign n28683 = pi648 & ~n28556;
  assign n28684 = ~n28682 & n28683;
  assign n28685 = ~pi619 & ~n28678;
  assign n28686 = pi619 & ~n28468;
  assign n28687 = ~pi1159 & ~n28686;
  assign n28688 = ~n28685 & n28687;
  assign n28689 = ~pi648 & ~n28552;
  assign n28690 = ~n28688 & n28689;
  assign n28691 = pi789 & ~n28690;
  assign n28692 = ~n28684 & n28691;
  assign n28693 = ~pi789 & n28678;
  assign n28694 = n17817 & ~n28693;
  assign n28695 = ~n28692 & n28694;
  assign n28696 = pi626 & ~n28559;
  assign n28697 = ~pi626 & ~n28437;
  assign n28698 = n17579 & ~n28697;
  assign n28699 = ~n28696 & n28698;
  assign n28700 = n17704 & n28470;
  assign n28701 = ~pi626 & ~n28559;
  assign n28702 = pi626 & ~n28437;
  assign n28703 = n17580 & ~n28702;
  assign n28704 = ~n28701 & n28703;
  assign n28705 = ~n28700 & ~n28704;
  assign n28706 = ~n28699 & n28705;
  assign n28707 = pi788 & ~n28706;
  assign n28708 = ~n20205 & ~n28707;
  assign n28709 = ~n28695 & n28708;
  assign n28710 = ~n28594 & ~n28709;
  assign n28711 = n20207 & ~n28710;
  assign n28712 = ~n20398 & n28565;
  assign n28713 = n17650 & ~n28488;
  assign n28714 = n17649 & ~n28492;
  assign n28715 = ~n28713 & ~n28714;
  assign n28716 = ~n28712 & n28715;
  assign n28717 = pi787 & ~n28716;
  assign n28718 = ~n28711 & ~n28717;
  assign n28719 = ~n28588 & n28718;
  assign n28720 = ~n28584 & ~n28719;
  assign n28721 = ~po1038 & ~n28720;
  assign n28722 = ~pi185 & po1038;
  assign n28723 = ~pi832 & ~n28722;
  assign n28724 = ~n28721 & n28723;
  assign po342 = ~n28436 & ~n28724;
  assign n28726 = pi186 & ~n3267;
  assign n28727 = ~pi186 & ~n17399;
  assign n28728 = pi752 & ~n28727;
  assign n28729 = pi186 & ~n19218;
  assign n28730 = ~pi186 & ~pi752;
  assign n28731 = n19223 & n28730;
  assign n28732 = ~n28729 & ~n28731;
  assign n28733 = ~n19217 & ~n28732;
  assign n28734 = ~n28728 & ~n28733;
  assign n28735 = ~pi703 & n28734;
  assign n28736 = ~pi186 & n19236;
  assign n28737 = pi186 & n19241;
  assign n28738 = pi752 & ~n19243;
  assign n28739 = ~n28737 & n28738;
  assign n28740 = ~n28736 & n28739;
  assign n28741 = pi186 & n19253;
  assign n28742 = ~pi186 & ~n19261;
  assign n28743 = ~pi752 & ~n28742;
  assign n28744 = ~n28741 & n28743;
  assign n28745 = pi703 & ~n28744;
  assign n28746 = ~n28740 & n28745;
  assign n28747 = n3267 & ~n28746;
  assign n28748 = ~n28735 & n28747;
  assign n28749 = ~n28726 & ~n28748;
  assign n28750 = ~pi625 & n28749;
  assign n28751 = n3267 & ~n28734;
  assign n28752 = ~n28726 & ~n28751;
  assign n28753 = pi625 & n28752;
  assign n28754 = ~pi1153 & ~n28753;
  assign n28755 = ~n28750 & n28754;
  assign n28756 = ~pi186 & n17972;
  assign n28757 = pi186 & ~n17976;
  assign n28758 = ~pi38 & ~n28757;
  assign n28759 = ~n28756 & n28758;
  assign n28760 = ~pi186 & ~n17280;
  assign n28761 = n17392 & ~n28760;
  assign n28762 = pi703 & ~n28761;
  assign n28763 = ~n28759 & n28762;
  assign n28764 = ~pi703 & n28727;
  assign n28765 = n3267 & ~n28764;
  assign n28766 = ~n28763 & n28765;
  assign n28767 = ~n28726 & ~n28766;
  assign n28768 = pi625 & n28767;
  assign n28769 = ~pi186 & ~n17406;
  assign n28770 = ~pi625 & n28769;
  assign n28771 = pi1153 & ~n28770;
  assign n28772 = ~n28768 & n28771;
  assign n28773 = ~pi608 & ~n28772;
  assign n28774 = ~n28755 & n28773;
  assign n28775 = pi625 & n28749;
  assign n28776 = ~pi625 & n28752;
  assign n28777 = pi1153 & ~n28776;
  assign n28778 = ~n28775 & n28777;
  assign n28779 = ~pi625 & n28767;
  assign n28780 = pi625 & n28769;
  assign n28781 = ~pi1153 & ~n28780;
  assign n28782 = ~n28779 & n28781;
  assign n28783 = pi608 & ~n28782;
  assign n28784 = ~n28778 & n28783;
  assign n28785 = ~n28774 & ~n28784;
  assign n28786 = pi778 & ~n28785;
  assign n28787 = ~pi778 & n28749;
  assign n28788 = ~n28786 & ~n28787;
  assign n28789 = ~pi609 & ~n28788;
  assign n28790 = ~pi778 & ~n28767;
  assign n28791 = ~n28772 & ~n28782;
  assign n28792 = pi778 & ~n28791;
  assign n28793 = ~n28790 & ~n28792;
  assign n28794 = pi609 & n28793;
  assign n28795 = ~pi1155 & ~n28794;
  assign n28796 = ~n28789 & n28795;
  assign n28797 = ~n17439 & ~n28769;
  assign n28798 = ~n17438 & ~n28752;
  assign n28799 = pi609 & n28798;
  assign n28800 = ~n28797 & ~n28799;
  assign n28801 = pi1155 & ~n28800;
  assign n28802 = ~pi660 & ~n28801;
  assign n28803 = ~n28796 & n28802;
  assign n28804 = pi609 & ~n28788;
  assign n28805 = ~pi609 & n28793;
  assign n28806 = pi1155 & ~n28805;
  assign n28807 = ~n28804 & n28806;
  assign n28808 = ~n17451 & ~n28769;
  assign n28809 = ~pi609 & n28798;
  assign n28810 = ~n28808 & ~n28809;
  assign n28811 = ~pi1155 & ~n28810;
  assign n28812 = pi660 & ~n28811;
  assign n28813 = ~n28807 & n28812;
  assign n28814 = ~n28803 & ~n28813;
  assign n28815 = pi785 & ~n28814;
  assign n28816 = ~pi785 & ~n28788;
  assign n28817 = ~n28815 & ~n28816;
  assign n28818 = ~pi618 & ~n28817;
  assign n28819 = ~n17466 & ~n28793;
  assign n28820 = n17466 & ~n28769;
  assign n28821 = ~n28819 & ~n28820;
  assign n28822 = pi618 & n28821;
  assign n28823 = ~pi1154 & ~n28822;
  assign n28824 = ~n28818 & n28823;
  assign n28825 = n17438 & ~n28769;
  assign n28826 = ~n28798 & ~n28825;
  assign n28827 = ~pi785 & ~n28826;
  assign n28828 = ~n28801 & ~n28811;
  assign n28829 = pi785 & ~n28828;
  assign n28830 = ~n28827 & ~n28829;
  assign n28831 = pi618 & n28830;
  assign n28832 = ~pi618 & n28769;
  assign n28833 = pi1154 & ~n28832;
  assign n28834 = ~n28831 & n28833;
  assign n28835 = ~pi627 & ~n28834;
  assign n28836 = ~n28824 & n28835;
  assign n28837 = pi618 & ~n28817;
  assign n28838 = ~pi618 & n28821;
  assign n28839 = pi1154 & ~n28838;
  assign n28840 = ~n28837 & n28839;
  assign n28841 = ~pi618 & n28830;
  assign n28842 = pi618 & n28769;
  assign n28843 = ~pi1154 & ~n28842;
  assign n28844 = ~n28841 & n28843;
  assign n28845 = pi627 & ~n28844;
  assign n28846 = ~n28840 & n28845;
  assign n28847 = ~n28836 & ~n28846;
  assign n28848 = pi781 & ~n28847;
  assign n28849 = ~pi781 & ~n28817;
  assign n28850 = ~n28848 & ~n28849;
  assign n28851 = ~pi619 & ~n28850;
  assign n28852 = ~n17503 & n28821;
  assign n28853 = n17503 & n28769;
  assign n28854 = ~n28852 & ~n28853;
  assign n28855 = pi619 & ~n28854;
  assign n28856 = ~pi1159 & ~n28855;
  assign n28857 = ~n28851 & n28856;
  assign n28858 = ~pi781 & ~n28830;
  assign n28859 = ~n28834 & ~n28844;
  assign n28860 = pi781 & ~n28859;
  assign n28861 = ~n28858 & ~n28860;
  assign n28862 = pi619 & n28861;
  assign n28863 = ~pi619 & n28769;
  assign n28864 = pi1159 & ~n28863;
  assign n28865 = ~n28862 & n28864;
  assign n28866 = ~pi648 & ~n28865;
  assign n28867 = ~n28857 & n28866;
  assign n28868 = pi619 & ~n28850;
  assign n28869 = ~pi619 & ~n28854;
  assign n28870 = pi1159 & ~n28869;
  assign n28871 = ~n28868 & n28870;
  assign n28872 = ~pi619 & n28861;
  assign n28873 = pi619 & n28769;
  assign n28874 = ~pi1159 & ~n28873;
  assign n28875 = ~n28872 & n28874;
  assign n28876 = pi648 & ~n28875;
  assign n28877 = ~n28871 & n28876;
  assign n28878 = ~n28867 & ~n28877;
  assign n28879 = pi789 & ~n28878;
  assign n28880 = ~pi789 & ~n28850;
  assign n28881 = ~n28879 & ~n28880;
  assign n28882 = ~pi788 & n28881;
  assign n28883 = ~pi626 & n28881;
  assign n28884 = n17539 & ~n28769;
  assign n28885 = ~n17539 & n28854;
  assign n28886 = ~n28884 & ~n28885;
  assign n28887 = pi626 & ~n28886;
  assign n28888 = ~pi641 & ~n28887;
  assign n28889 = ~n28883 & n28888;
  assign n28890 = ~pi789 & ~n28861;
  assign n28891 = ~n28865 & ~n28875;
  assign n28892 = pi789 & ~n28891;
  assign n28893 = ~n28890 & ~n28892;
  assign n28894 = ~pi626 & ~n28893;
  assign n28895 = pi626 & ~n28769;
  assign n28896 = pi641 & ~n28895;
  assign n28897 = ~n28894 & n28896;
  assign n28898 = ~pi1158 & ~n28897;
  assign n28899 = ~n28889 & n28898;
  assign n28900 = pi626 & n28881;
  assign n28901 = ~pi626 & ~n28886;
  assign n28902 = pi641 & ~n28901;
  assign n28903 = ~n28900 & n28902;
  assign n28904 = pi626 & ~n28893;
  assign n28905 = ~pi626 & ~n28769;
  assign n28906 = ~pi641 & ~n28905;
  assign n28907 = ~n28904 & n28906;
  assign n28908 = pi1158 & ~n28907;
  assign n28909 = ~n28903 & n28908;
  assign n28910 = ~n28899 & ~n28909;
  assign n28911 = pi788 & ~n28910;
  assign n28912 = ~n28882 & ~n28911;
  assign n28913 = ~pi628 & n28912;
  assign n28914 = ~n17816 & n28893;
  assign n28915 = n17816 & n28769;
  assign n28916 = ~n28914 & ~n28915;
  assign n28917 = pi628 & ~n28916;
  assign n28918 = ~pi1156 & ~n28917;
  assign n28919 = ~n28913 & n28918;
  assign n28920 = ~n17582 & n28886;
  assign n28921 = n17582 & n28769;
  assign n28922 = ~n28920 & ~n28921;
  assign n28923 = pi628 & ~n28922;
  assign n28924 = ~pi628 & n28769;
  assign n28925 = pi1156 & ~n28924;
  assign n28926 = ~n28923 & n28925;
  assign n28927 = ~pi629 & ~n28926;
  assign n28928 = ~n28919 & n28927;
  assign n28929 = pi628 & n28912;
  assign n28930 = ~pi628 & ~n28916;
  assign n28931 = pi1156 & ~n28930;
  assign n28932 = ~n28929 & n28931;
  assign n28933 = ~pi628 & ~n28922;
  assign n28934 = pi628 & n28769;
  assign n28935 = ~pi1156 & ~n28934;
  assign n28936 = ~n28933 & n28935;
  assign n28937 = pi629 & ~n28936;
  assign n28938 = ~n28932 & n28937;
  assign n28939 = ~n28928 & ~n28938;
  assign n28940 = pi792 & ~n28939;
  assign n28941 = ~pi792 & n28912;
  assign n28942 = ~n28940 & ~n28941;
  assign n28943 = ~pi647 & ~n28942;
  assign n28944 = ~n17610 & ~n28916;
  assign n28945 = n17610 & n28769;
  assign n28946 = ~n28944 & ~n28945;
  assign n28947 = pi647 & ~n28946;
  assign n28948 = ~pi1157 & ~n28947;
  assign n28949 = ~n28943 & n28948;
  assign n28950 = ~pi792 & n28922;
  assign n28951 = ~n28926 & ~n28936;
  assign n28952 = pi792 & ~n28951;
  assign n28953 = ~n28950 & ~n28952;
  assign n28954 = pi647 & n28953;
  assign n28955 = ~pi647 & n28769;
  assign n28956 = pi1157 & ~n28955;
  assign n28957 = ~n28954 & n28956;
  assign n28958 = ~pi630 & ~n28957;
  assign n28959 = ~n28949 & n28958;
  assign n28960 = pi647 & ~n28942;
  assign n28961 = ~pi647 & ~n28946;
  assign n28962 = pi1157 & ~n28961;
  assign n28963 = ~n28960 & n28962;
  assign n28964 = ~pi647 & n28953;
  assign n28965 = pi647 & n28769;
  assign n28966 = ~pi1157 & ~n28965;
  assign n28967 = ~n28964 & n28966;
  assign n28968 = pi630 & ~n28967;
  assign n28969 = ~n28963 & n28968;
  assign n28970 = ~n28959 & ~n28969;
  assign n28971 = pi787 & ~n28970;
  assign n28972 = ~pi787 & ~n28942;
  assign n28973 = ~n28971 & ~n28972;
  assign n28974 = ~pi644 & ~n28973;
  assign n28975 = ~pi787 & ~n28953;
  assign n28976 = ~n28957 & ~n28967;
  assign n28977 = pi787 & ~n28976;
  assign n28978 = ~n28975 & ~n28977;
  assign n28979 = pi644 & n28978;
  assign n28980 = ~pi715 & ~n28979;
  assign n28981 = ~n28974 & n28980;
  assign n28982 = n17652 & ~n28769;
  assign n28983 = ~n17652 & n28946;
  assign n28984 = ~n28982 & ~n28983;
  assign n28985 = ~pi644 & n28984;
  assign n28986 = pi644 & n28769;
  assign n28987 = pi715 & ~n28986;
  assign n28988 = ~n28985 & n28987;
  assign n28989 = ~pi1160 & ~n28988;
  assign n28990 = ~n28981 & n28989;
  assign n28991 = pi644 & ~n28973;
  assign n28992 = ~pi644 & n28978;
  assign n28993 = pi715 & ~n28992;
  assign n28994 = ~n28991 & n28993;
  assign n28995 = pi644 & n28984;
  assign n28996 = ~pi644 & n28769;
  assign n28997 = ~pi715 & ~n28996;
  assign n28998 = ~n28995 & n28997;
  assign n28999 = pi1160 & ~n28998;
  assign n29000 = ~n28994 & n28999;
  assign n29001 = pi790 & ~n29000;
  assign n29002 = ~n28990 & n29001;
  assign n29003 = ~pi790 & n28973;
  assign n29004 = ~po1038 & ~n29003;
  assign n29005 = ~n29002 & n29004;
  assign n29006 = ~pi186 & po1038;
  assign n29007 = ~pi832 & ~n29006;
  assign n29008 = ~n29005 & n29007;
  assign n29009 = ~pi186 & ~n2754;
  assign n29010 = ~pi752 & n16784;
  assign n29011 = ~n29009 & ~n29010;
  assign n29012 = ~n17706 & ~n29011;
  assign n29013 = ~pi785 & ~n29012;
  assign n29014 = ~n17711 & ~n29011;
  assign n29015 = pi1155 & ~n29014;
  assign n29016 = ~n17714 & n29012;
  assign n29017 = ~pi1155 & ~n29016;
  assign n29018 = ~n29015 & ~n29017;
  assign n29019 = pi785 & ~n29018;
  assign n29020 = ~n29013 & ~n29019;
  assign n29021 = ~pi781 & ~n29020;
  assign n29022 = ~n17721 & n29020;
  assign n29023 = pi1154 & ~n29022;
  assign n29024 = ~n17724 & n29020;
  assign n29025 = ~pi1154 & ~n29024;
  assign n29026 = ~n29023 & ~n29025;
  assign n29027 = pi781 & ~n29026;
  assign n29028 = ~n29021 & ~n29027;
  assign n29029 = ~pi789 & ~n29028;
  assign n29030 = pi619 & n29028;
  assign n29031 = ~pi619 & n29009;
  assign n29032 = pi1159 & ~n29031;
  assign n29033 = ~n29030 & n29032;
  assign n29034 = ~pi619 & n29028;
  assign n29035 = pi619 & n29009;
  assign n29036 = ~pi1159 & ~n29035;
  assign n29037 = ~n29034 & n29036;
  assign n29038 = ~n29033 & ~n29037;
  assign n29039 = pi789 & ~n29038;
  assign n29040 = ~n29029 & ~n29039;
  assign n29041 = ~n17816 & n29040;
  assign n29042 = n17816 & n29009;
  assign n29043 = ~n29041 & ~n29042;
  assign n29044 = ~n17610 & ~n29043;
  assign n29045 = n17610 & n29009;
  assign n29046 = ~n29044 & ~n29045;
  assign n29047 = ~n20398 & n29046;
  assign n29048 = pi703 & n16786;
  assign n29049 = ~n29009 & ~n29048;
  assign n29050 = ~pi778 & n29049;
  assign n29051 = ~pi625 & n29048;
  assign n29052 = ~n29049 & ~n29051;
  assign n29053 = pi1153 & ~n29052;
  assign n29054 = ~pi1153 & ~n29009;
  assign n29055 = ~n29051 & n29054;
  assign n29056 = ~n29053 & ~n29055;
  assign n29057 = pi778 & ~n29056;
  assign n29058 = ~n29050 & ~n29057;
  assign n29059 = ~n17692 & n29058;
  assign n29060 = ~n17694 & n29059;
  assign n29061 = ~n17696 & n29060;
  assign n29062 = ~n17828 & n29061;
  assign n29063 = ~n17859 & n29062;
  assign n29064 = ~pi647 & n29063;
  assign n29065 = pi647 & n29009;
  assign n29066 = ~pi1157 & ~n29065;
  assign n29067 = ~n29064 & n29066;
  assign n29068 = pi647 & ~n29063;
  assign n29069 = ~pi647 & ~n29009;
  assign n29070 = ~n29068 & ~n29069;
  assign n29071 = pi1157 & ~n29070;
  assign n29072 = ~n29067 & ~n29071;
  assign n29073 = ~n17651 & ~n29072;
  assign n29074 = ~n29047 & ~n29073;
  assign n29075 = pi787 & ~n29074;
  assign n29076 = pi626 & ~n29040;
  assign n29077 = ~pi626 & ~n29009;
  assign n29078 = n17579 & ~n29077;
  assign n29079 = ~n29076 & n29078;
  assign n29080 = n17704 & n29061;
  assign n29081 = ~pi626 & ~n29040;
  assign n29082 = pi626 & ~n29009;
  assign n29083 = n17580 & ~n29082;
  assign n29084 = ~n29081 & n29083;
  assign n29085 = ~n29080 & ~n29084;
  assign n29086 = ~n29079 & n29085;
  assign n29087 = pi788 & ~n29086;
  assign n29088 = ~n16521 & ~n29049;
  assign n29089 = pi625 & n29088;
  assign n29090 = n29011 & ~n29088;
  assign n29091 = ~n29089 & ~n29090;
  assign n29092 = n29054 & ~n29091;
  assign n29093 = ~pi608 & ~n29053;
  assign n29094 = ~n29092 & n29093;
  assign n29095 = pi1153 & n29011;
  assign n29096 = ~n29089 & n29095;
  assign n29097 = pi608 & ~n29055;
  assign n29098 = ~n29096 & n29097;
  assign n29099 = ~n29094 & ~n29098;
  assign n29100 = pi778 & ~n29099;
  assign n29101 = ~pi778 & ~n29090;
  assign n29102 = ~n29100 & ~n29101;
  assign n29103 = ~pi609 & ~n29102;
  assign n29104 = pi609 & n29058;
  assign n29105 = ~pi1155 & ~n29104;
  assign n29106 = ~n29103 & n29105;
  assign n29107 = ~pi660 & ~n29015;
  assign n29108 = ~n29106 & n29107;
  assign n29109 = pi609 & ~n29102;
  assign n29110 = ~pi609 & n29058;
  assign n29111 = pi1155 & ~n29110;
  assign n29112 = ~n29109 & n29111;
  assign n29113 = pi660 & ~n29017;
  assign n29114 = ~n29112 & n29113;
  assign n29115 = ~n29108 & ~n29114;
  assign n29116 = pi785 & ~n29115;
  assign n29117 = ~pi785 & ~n29102;
  assign n29118 = ~n29116 & ~n29117;
  assign n29119 = ~pi618 & ~n29118;
  assign n29120 = pi618 & n29059;
  assign n29121 = ~pi1154 & ~n29120;
  assign n29122 = ~n29119 & n29121;
  assign n29123 = ~pi627 & ~n29023;
  assign n29124 = ~n29122 & n29123;
  assign n29125 = pi618 & ~n29118;
  assign n29126 = ~pi618 & n29059;
  assign n29127 = pi1154 & ~n29126;
  assign n29128 = ~n29125 & n29127;
  assign n29129 = pi627 & ~n29025;
  assign n29130 = ~n29128 & n29129;
  assign n29131 = ~n29124 & ~n29130;
  assign n29132 = pi781 & ~n29131;
  assign n29133 = ~pi781 & ~n29118;
  assign n29134 = ~n29132 & ~n29133;
  assign n29135 = pi619 & ~n29134;
  assign n29136 = ~pi619 & n29060;
  assign n29137 = pi1159 & ~n29136;
  assign n29138 = ~n29135 & n29137;
  assign n29139 = pi648 & ~n29037;
  assign n29140 = ~n29138 & n29139;
  assign n29141 = ~pi619 & ~n29134;
  assign n29142 = pi619 & n29060;
  assign n29143 = ~pi1159 & ~n29142;
  assign n29144 = ~n29141 & n29143;
  assign n29145 = ~pi648 & ~n29033;
  assign n29146 = ~n29144 & n29145;
  assign n29147 = pi789 & ~n29146;
  assign n29148 = ~n29140 & n29147;
  assign n29149 = ~pi789 & n29134;
  assign n29150 = n17817 & ~n29149;
  assign n29151 = ~n29148 & n29150;
  assign n29152 = ~n29087 & ~n29151;
  assign n29153 = ~n20205 & ~n29152;
  assign n29154 = n17856 & ~n29043;
  assign n29155 = n20693 & n29062;
  assign n29156 = ~n29154 & ~n29155;
  assign n29157 = ~pi629 & ~n29156;
  assign n29158 = n20697 & n29062;
  assign n29159 = n17855 & ~n29043;
  assign n29160 = ~n29158 & ~n29159;
  assign n29161 = pi629 & ~n29160;
  assign n29162 = ~n29157 & ~n29161;
  assign n29163 = pi792 & ~n29162;
  assign n29164 = n20207 & ~n29163;
  assign n29165 = ~n29153 & n29164;
  assign n29166 = ~n29075 & ~n29165;
  assign n29167 = pi644 & n29166;
  assign n29168 = ~pi787 & ~n29063;
  assign n29169 = pi787 & ~n29072;
  assign n29170 = ~n29168 & ~n29169;
  assign n29171 = ~pi644 & n29170;
  assign n29172 = pi715 & ~n29171;
  assign n29173 = ~n29167 & n29172;
  assign n29174 = ~n17652 & ~n29046;
  assign n29175 = n17652 & n29009;
  assign n29176 = ~n29174 & ~n29175;
  assign n29177 = pi644 & ~n29176;
  assign n29178 = ~pi644 & n29009;
  assign n29179 = ~pi715 & ~n29178;
  assign n29180 = ~n29177 & n29179;
  assign n29181 = pi1160 & ~n29180;
  assign n29182 = ~n29173 & n29181;
  assign n29183 = ~pi644 & n29166;
  assign n29184 = pi644 & n29170;
  assign n29185 = ~pi715 & ~n29184;
  assign n29186 = ~n29183 & n29185;
  assign n29187 = ~pi644 & ~n29176;
  assign n29188 = pi644 & n29009;
  assign n29189 = pi715 & ~n29188;
  assign n29190 = ~n29187 & n29189;
  assign n29191 = ~pi1160 & ~n29190;
  assign n29192 = ~n29186 & n29191;
  assign n29193 = ~n29182 & ~n29192;
  assign n29194 = pi790 & ~n29193;
  assign n29195 = ~pi790 & n29166;
  assign n29196 = pi832 & ~n29195;
  assign n29197 = ~n29194 & n29196;
  assign po343 = ~n29008 & ~n29197;
  assign n29199 = pi187 & ~n3267;
  assign n29200 = ~pi770 & ~n19223;
  assign n29201 = ~n20851 & ~n29200;
  assign n29202 = ~pi187 & ~n29201;
  assign n29203 = ~pi187 & ~n19217;
  assign n29204 = ~pi770 & ~n29203;
  assign n29205 = ~n24271 & n29204;
  assign n29206 = ~n29202 & ~n29205;
  assign n29207 = ~pi726 & ~n29206;
  assign n29208 = ~pi187 & n19236;
  assign n29209 = pi187 & n19241;
  assign n29210 = pi770 & ~n19243;
  assign n29211 = ~n29209 & n29210;
  assign n29212 = ~n29208 & n29211;
  assign n29213 = pi187 & n19253;
  assign n29214 = ~pi187 & ~n19261;
  assign n29215 = ~pi770 & ~n29214;
  assign n29216 = ~n29213 & n29215;
  assign n29217 = pi726 & ~n29216;
  assign n29218 = ~n29212 & n29217;
  assign n29219 = n3267 & ~n29218;
  assign n29220 = ~n29207 & n29219;
  assign n29221 = ~n29199 & ~n29220;
  assign n29222 = ~pi625 & n29221;
  assign n29223 = n3267 & n29206;
  assign n29224 = ~n29199 & ~n29223;
  assign n29225 = pi625 & n29224;
  assign n29226 = ~pi1153 & ~n29225;
  assign n29227 = ~n29222 & n29226;
  assign n29228 = ~pi187 & n17972;
  assign n29229 = pi187 & ~n17976;
  assign n29230 = ~pi38 & ~n29229;
  assign n29231 = ~n29228 & n29230;
  assign n29232 = ~pi187 & ~n17280;
  assign n29233 = n17392 & ~n29232;
  assign n29234 = pi726 & ~n29233;
  assign n29235 = ~n29231 & n29234;
  assign n29236 = ~pi187 & ~pi726;
  assign n29237 = ~n17399 & n29236;
  assign n29238 = n3267 & ~n29237;
  assign n29239 = ~n29235 & n29238;
  assign n29240 = ~n29199 & ~n29239;
  assign n29241 = pi625 & n29240;
  assign n29242 = ~pi187 & ~n17406;
  assign n29243 = ~pi625 & n29242;
  assign n29244 = pi1153 & ~n29243;
  assign n29245 = ~n29241 & n29244;
  assign n29246 = ~pi608 & ~n29245;
  assign n29247 = ~n29227 & n29246;
  assign n29248 = pi625 & n29221;
  assign n29249 = ~pi625 & n29224;
  assign n29250 = pi1153 & ~n29249;
  assign n29251 = ~n29248 & n29250;
  assign n29252 = ~pi625 & n29240;
  assign n29253 = pi625 & n29242;
  assign n29254 = ~pi1153 & ~n29253;
  assign n29255 = ~n29252 & n29254;
  assign n29256 = pi608 & ~n29255;
  assign n29257 = ~n29251 & n29256;
  assign n29258 = ~n29247 & ~n29257;
  assign n29259 = pi778 & ~n29258;
  assign n29260 = ~pi778 & n29221;
  assign n29261 = ~n29259 & ~n29260;
  assign n29262 = ~pi609 & ~n29261;
  assign n29263 = ~pi778 & ~n29240;
  assign n29264 = ~n29245 & ~n29255;
  assign n29265 = pi778 & ~n29264;
  assign n29266 = ~n29263 & ~n29265;
  assign n29267 = pi609 & n29266;
  assign n29268 = ~pi1155 & ~n29267;
  assign n29269 = ~n29262 & n29268;
  assign n29270 = ~n17439 & ~n29242;
  assign n29271 = ~n17438 & ~n29224;
  assign n29272 = pi609 & n29271;
  assign n29273 = ~n29270 & ~n29272;
  assign n29274 = pi1155 & ~n29273;
  assign n29275 = ~pi660 & ~n29274;
  assign n29276 = ~n29269 & n29275;
  assign n29277 = pi609 & ~n29261;
  assign n29278 = ~pi609 & n29266;
  assign n29279 = pi1155 & ~n29278;
  assign n29280 = ~n29277 & n29279;
  assign n29281 = ~n17451 & ~n29242;
  assign n29282 = ~pi609 & n29271;
  assign n29283 = ~n29281 & ~n29282;
  assign n29284 = ~pi1155 & ~n29283;
  assign n29285 = pi660 & ~n29284;
  assign n29286 = ~n29280 & n29285;
  assign n29287 = ~n29276 & ~n29286;
  assign n29288 = pi785 & ~n29287;
  assign n29289 = ~pi785 & ~n29261;
  assign n29290 = ~n29288 & ~n29289;
  assign n29291 = ~pi618 & ~n29290;
  assign n29292 = ~n17466 & ~n29266;
  assign n29293 = n17466 & ~n29242;
  assign n29294 = ~n29292 & ~n29293;
  assign n29295 = pi618 & n29294;
  assign n29296 = ~pi1154 & ~n29295;
  assign n29297 = ~n29291 & n29296;
  assign n29298 = n17438 & ~n29242;
  assign n29299 = ~n29271 & ~n29298;
  assign n29300 = ~pi785 & ~n29299;
  assign n29301 = ~n29274 & ~n29284;
  assign n29302 = pi785 & ~n29301;
  assign n29303 = ~n29300 & ~n29302;
  assign n29304 = pi618 & n29303;
  assign n29305 = ~pi618 & n29242;
  assign n29306 = pi1154 & ~n29305;
  assign n29307 = ~n29304 & n29306;
  assign n29308 = ~pi627 & ~n29307;
  assign n29309 = ~n29297 & n29308;
  assign n29310 = pi618 & ~n29290;
  assign n29311 = ~pi618 & n29294;
  assign n29312 = pi1154 & ~n29311;
  assign n29313 = ~n29310 & n29312;
  assign n29314 = ~pi618 & n29303;
  assign n29315 = pi618 & n29242;
  assign n29316 = ~pi1154 & ~n29315;
  assign n29317 = ~n29314 & n29316;
  assign n29318 = pi627 & ~n29317;
  assign n29319 = ~n29313 & n29318;
  assign n29320 = ~n29309 & ~n29319;
  assign n29321 = pi781 & ~n29320;
  assign n29322 = ~pi781 & ~n29290;
  assign n29323 = ~n29321 & ~n29322;
  assign n29324 = ~pi619 & ~n29323;
  assign n29325 = ~n17503 & n29294;
  assign n29326 = n17503 & n29242;
  assign n29327 = ~n29325 & ~n29326;
  assign n29328 = pi619 & ~n29327;
  assign n29329 = ~pi1159 & ~n29328;
  assign n29330 = ~n29324 & n29329;
  assign n29331 = ~pi781 & ~n29303;
  assign n29332 = ~n29307 & ~n29317;
  assign n29333 = pi781 & ~n29332;
  assign n29334 = ~n29331 & ~n29333;
  assign n29335 = pi619 & n29334;
  assign n29336 = ~pi619 & n29242;
  assign n29337 = pi1159 & ~n29336;
  assign n29338 = ~n29335 & n29337;
  assign n29339 = ~pi648 & ~n29338;
  assign n29340 = ~n29330 & n29339;
  assign n29341 = pi619 & ~n29323;
  assign n29342 = ~pi619 & ~n29327;
  assign n29343 = pi1159 & ~n29342;
  assign n29344 = ~n29341 & n29343;
  assign n29345 = ~pi619 & n29334;
  assign n29346 = pi619 & n29242;
  assign n29347 = ~pi1159 & ~n29346;
  assign n29348 = ~n29345 & n29347;
  assign n29349 = pi648 & ~n29348;
  assign n29350 = ~n29344 & n29349;
  assign n29351 = ~n29340 & ~n29350;
  assign n29352 = pi789 & ~n29351;
  assign n29353 = ~pi789 & ~n29323;
  assign n29354 = ~n29352 & ~n29353;
  assign n29355 = ~pi788 & n29354;
  assign n29356 = ~pi626 & n29354;
  assign n29357 = n17539 & ~n29242;
  assign n29358 = ~n17539 & n29327;
  assign n29359 = ~n29357 & ~n29358;
  assign n29360 = pi626 & ~n29359;
  assign n29361 = ~pi641 & ~n29360;
  assign n29362 = ~n29356 & n29361;
  assign n29363 = ~pi789 & ~n29334;
  assign n29364 = ~n29338 & ~n29348;
  assign n29365 = pi789 & ~n29364;
  assign n29366 = ~n29363 & ~n29365;
  assign n29367 = ~pi626 & ~n29366;
  assign n29368 = pi626 & ~n29242;
  assign n29369 = pi641 & ~n29368;
  assign n29370 = ~n29367 & n29369;
  assign n29371 = ~pi1158 & ~n29370;
  assign n29372 = ~n29362 & n29371;
  assign n29373 = pi626 & n29354;
  assign n29374 = ~pi626 & ~n29359;
  assign n29375 = pi641 & ~n29374;
  assign n29376 = ~n29373 & n29375;
  assign n29377 = pi626 & ~n29366;
  assign n29378 = ~pi626 & ~n29242;
  assign n29379 = ~pi641 & ~n29378;
  assign n29380 = ~n29377 & n29379;
  assign n29381 = pi1158 & ~n29380;
  assign n29382 = ~n29376 & n29381;
  assign n29383 = ~n29372 & ~n29382;
  assign n29384 = pi788 & ~n29383;
  assign n29385 = ~n29355 & ~n29384;
  assign n29386 = ~pi628 & n29385;
  assign n29387 = ~n17816 & n29366;
  assign n29388 = n17816 & n29242;
  assign n29389 = ~n29387 & ~n29388;
  assign n29390 = pi628 & ~n29389;
  assign n29391 = ~pi1156 & ~n29390;
  assign n29392 = ~n29386 & n29391;
  assign n29393 = ~n17582 & n29359;
  assign n29394 = n17582 & n29242;
  assign n29395 = ~n29393 & ~n29394;
  assign n29396 = pi628 & ~n29395;
  assign n29397 = ~pi628 & n29242;
  assign n29398 = pi1156 & ~n29397;
  assign n29399 = ~n29396 & n29398;
  assign n29400 = ~pi629 & ~n29399;
  assign n29401 = ~n29392 & n29400;
  assign n29402 = pi628 & n29385;
  assign n29403 = ~pi628 & ~n29389;
  assign n29404 = pi1156 & ~n29403;
  assign n29405 = ~n29402 & n29404;
  assign n29406 = ~pi628 & ~n29395;
  assign n29407 = pi628 & n29242;
  assign n29408 = ~pi1156 & ~n29407;
  assign n29409 = ~n29406 & n29408;
  assign n29410 = pi629 & ~n29409;
  assign n29411 = ~n29405 & n29410;
  assign n29412 = ~n29401 & ~n29411;
  assign n29413 = pi792 & ~n29412;
  assign n29414 = ~pi792 & n29385;
  assign n29415 = ~n29413 & ~n29414;
  assign n29416 = ~pi647 & ~n29415;
  assign n29417 = ~n17610 & ~n29389;
  assign n29418 = n17610 & n29242;
  assign n29419 = ~n29417 & ~n29418;
  assign n29420 = pi647 & ~n29419;
  assign n29421 = ~pi1157 & ~n29420;
  assign n29422 = ~n29416 & n29421;
  assign n29423 = ~pi792 & n29395;
  assign n29424 = ~n29399 & ~n29409;
  assign n29425 = pi792 & ~n29424;
  assign n29426 = ~n29423 & ~n29425;
  assign n29427 = pi647 & n29426;
  assign n29428 = ~pi647 & n29242;
  assign n29429 = pi1157 & ~n29428;
  assign n29430 = ~n29427 & n29429;
  assign n29431 = ~pi630 & ~n29430;
  assign n29432 = ~n29422 & n29431;
  assign n29433 = pi647 & ~n29415;
  assign n29434 = ~pi647 & ~n29419;
  assign n29435 = pi1157 & ~n29434;
  assign n29436 = ~n29433 & n29435;
  assign n29437 = ~pi647 & n29426;
  assign n29438 = pi647 & n29242;
  assign n29439 = ~pi1157 & ~n29438;
  assign n29440 = ~n29437 & n29439;
  assign n29441 = pi630 & ~n29440;
  assign n29442 = ~n29436 & n29441;
  assign n29443 = ~n29432 & ~n29442;
  assign n29444 = pi787 & ~n29443;
  assign n29445 = ~pi787 & ~n29415;
  assign n29446 = ~n29444 & ~n29445;
  assign n29447 = ~pi644 & ~n29446;
  assign n29448 = ~pi787 & ~n29426;
  assign n29449 = ~n29430 & ~n29440;
  assign n29450 = pi787 & ~n29449;
  assign n29451 = ~n29448 & ~n29450;
  assign n29452 = pi644 & n29451;
  assign n29453 = ~pi715 & ~n29452;
  assign n29454 = ~n29447 & n29453;
  assign n29455 = n17652 & ~n29242;
  assign n29456 = ~n17652 & n29419;
  assign n29457 = ~n29455 & ~n29456;
  assign n29458 = ~pi644 & n29457;
  assign n29459 = pi644 & n29242;
  assign n29460 = pi715 & ~n29459;
  assign n29461 = ~n29458 & n29460;
  assign n29462 = ~pi1160 & ~n29461;
  assign n29463 = ~n29454 & n29462;
  assign n29464 = pi644 & ~n29446;
  assign n29465 = ~pi644 & n29451;
  assign n29466 = pi715 & ~n29465;
  assign n29467 = ~n29464 & n29466;
  assign n29468 = pi644 & n29457;
  assign n29469 = ~pi644 & n29242;
  assign n29470 = ~pi715 & ~n29469;
  assign n29471 = ~n29468 & n29470;
  assign n29472 = pi1160 & ~n29471;
  assign n29473 = ~n29467 & n29472;
  assign n29474 = pi790 & ~n29473;
  assign n29475 = ~n29463 & n29474;
  assign n29476 = ~pi790 & n29446;
  assign n29477 = ~po1038 & ~n29476;
  assign n29478 = ~n29475 & n29477;
  assign n29479 = ~pi187 & po1038;
  assign n29480 = ~pi832 & ~n29479;
  assign n29481 = ~n29478 & n29480;
  assign n29482 = ~pi187 & ~n2754;
  assign n29483 = ~pi770 & n16784;
  assign n29484 = ~n29482 & ~n29483;
  assign n29485 = ~n17706 & ~n29484;
  assign n29486 = ~pi785 & ~n29485;
  assign n29487 = ~n17711 & ~n29484;
  assign n29488 = pi1155 & ~n29487;
  assign n29489 = ~n17714 & n29485;
  assign n29490 = ~pi1155 & ~n29489;
  assign n29491 = ~n29488 & ~n29490;
  assign n29492 = pi785 & ~n29491;
  assign n29493 = ~n29486 & ~n29492;
  assign n29494 = ~pi781 & ~n29493;
  assign n29495 = ~n17721 & n29493;
  assign n29496 = pi1154 & ~n29495;
  assign n29497 = ~n17724 & n29493;
  assign n29498 = ~pi1154 & ~n29497;
  assign n29499 = ~n29496 & ~n29498;
  assign n29500 = pi781 & ~n29499;
  assign n29501 = ~n29494 & ~n29500;
  assign n29502 = ~pi789 & ~n29501;
  assign n29503 = pi619 & n29501;
  assign n29504 = ~pi619 & n29482;
  assign n29505 = pi1159 & ~n29504;
  assign n29506 = ~n29503 & n29505;
  assign n29507 = ~pi619 & n29501;
  assign n29508 = pi619 & n29482;
  assign n29509 = ~pi1159 & ~n29508;
  assign n29510 = ~n29507 & n29509;
  assign n29511 = ~n29506 & ~n29510;
  assign n29512 = pi789 & ~n29511;
  assign n29513 = ~n29502 & ~n29512;
  assign n29514 = ~n17816 & n29513;
  assign n29515 = n17816 & n29482;
  assign n29516 = ~n29514 & ~n29515;
  assign n29517 = ~n17610 & ~n29516;
  assign n29518 = n17610 & n29482;
  assign n29519 = ~n29517 & ~n29518;
  assign n29520 = ~n20398 & n29519;
  assign n29521 = pi726 & n16786;
  assign n29522 = ~n29482 & ~n29521;
  assign n29523 = ~pi778 & n29522;
  assign n29524 = ~pi625 & n29521;
  assign n29525 = ~n29522 & ~n29524;
  assign n29526 = pi1153 & ~n29525;
  assign n29527 = ~pi1153 & ~n29482;
  assign n29528 = ~n29524 & n29527;
  assign n29529 = ~n29526 & ~n29528;
  assign n29530 = pi778 & ~n29529;
  assign n29531 = ~n29523 & ~n29530;
  assign n29532 = ~n17692 & n29531;
  assign n29533 = ~n17694 & n29532;
  assign n29534 = ~n17696 & n29533;
  assign n29535 = ~n17828 & n29534;
  assign n29536 = ~n17859 & n29535;
  assign n29537 = ~pi647 & n29536;
  assign n29538 = pi647 & n29482;
  assign n29539 = ~pi1157 & ~n29538;
  assign n29540 = ~n29537 & n29539;
  assign n29541 = pi647 & ~n29536;
  assign n29542 = ~pi647 & ~n29482;
  assign n29543 = ~n29541 & ~n29542;
  assign n29544 = pi1157 & ~n29543;
  assign n29545 = ~n29540 & ~n29544;
  assign n29546 = ~n17651 & ~n29545;
  assign n29547 = ~n29520 & ~n29546;
  assign n29548 = pi787 & ~n29547;
  assign n29549 = pi626 & ~n29513;
  assign n29550 = ~pi626 & ~n29482;
  assign n29551 = n17579 & ~n29550;
  assign n29552 = ~n29549 & n29551;
  assign n29553 = n17704 & n29534;
  assign n29554 = ~pi626 & ~n29513;
  assign n29555 = pi626 & ~n29482;
  assign n29556 = n17580 & ~n29555;
  assign n29557 = ~n29554 & n29556;
  assign n29558 = ~n29553 & ~n29557;
  assign n29559 = ~n29552 & n29558;
  assign n29560 = pi788 & ~n29559;
  assign n29561 = ~n16521 & ~n29522;
  assign n29562 = pi625 & n29561;
  assign n29563 = n29484 & ~n29561;
  assign n29564 = ~n29562 & ~n29563;
  assign n29565 = n29527 & ~n29564;
  assign n29566 = ~pi608 & ~n29526;
  assign n29567 = ~n29565 & n29566;
  assign n29568 = pi1153 & n29484;
  assign n29569 = ~n29562 & n29568;
  assign n29570 = pi608 & ~n29528;
  assign n29571 = ~n29569 & n29570;
  assign n29572 = ~n29567 & ~n29571;
  assign n29573 = pi778 & ~n29572;
  assign n29574 = ~pi778 & ~n29563;
  assign n29575 = ~n29573 & ~n29574;
  assign n29576 = ~pi609 & ~n29575;
  assign n29577 = pi609 & n29531;
  assign n29578 = ~pi1155 & ~n29577;
  assign n29579 = ~n29576 & n29578;
  assign n29580 = ~pi660 & ~n29488;
  assign n29581 = ~n29579 & n29580;
  assign n29582 = pi609 & ~n29575;
  assign n29583 = ~pi609 & n29531;
  assign n29584 = pi1155 & ~n29583;
  assign n29585 = ~n29582 & n29584;
  assign n29586 = pi660 & ~n29490;
  assign n29587 = ~n29585 & n29586;
  assign n29588 = ~n29581 & ~n29587;
  assign n29589 = pi785 & ~n29588;
  assign n29590 = ~pi785 & ~n29575;
  assign n29591 = ~n29589 & ~n29590;
  assign n29592 = ~pi618 & ~n29591;
  assign n29593 = pi618 & n29532;
  assign n29594 = ~pi1154 & ~n29593;
  assign n29595 = ~n29592 & n29594;
  assign n29596 = ~pi627 & ~n29496;
  assign n29597 = ~n29595 & n29596;
  assign n29598 = pi618 & ~n29591;
  assign n29599 = ~pi618 & n29532;
  assign n29600 = pi1154 & ~n29599;
  assign n29601 = ~n29598 & n29600;
  assign n29602 = pi627 & ~n29498;
  assign n29603 = ~n29601 & n29602;
  assign n29604 = ~n29597 & ~n29603;
  assign n29605 = pi781 & ~n29604;
  assign n29606 = ~pi781 & ~n29591;
  assign n29607 = ~n29605 & ~n29606;
  assign n29608 = pi619 & ~n29607;
  assign n29609 = ~pi619 & n29533;
  assign n29610 = pi1159 & ~n29609;
  assign n29611 = ~n29608 & n29610;
  assign n29612 = pi648 & ~n29510;
  assign n29613 = ~n29611 & n29612;
  assign n29614 = ~pi619 & ~n29607;
  assign n29615 = pi619 & n29533;
  assign n29616 = ~pi1159 & ~n29615;
  assign n29617 = ~n29614 & n29616;
  assign n29618 = ~pi648 & ~n29506;
  assign n29619 = ~n29617 & n29618;
  assign n29620 = pi789 & ~n29619;
  assign n29621 = ~n29613 & n29620;
  assign n29622 = ~pi789 & n29607;
  assign n29623 = n17817 & ~n29622;
  assign n29624 = ~n29621 & n29623;
  assign n29625 = ~n29560 & ~n29624;
  assign n29626 = ~n20205 & ~n29625;
  assign n29627 = n17856 & ~n29516;
  assign n29628 = n20693 & n29535;
  assign n29629 = ~n29627 & ~n29628;
  assign n29630 = ~pi629 & ~n29629;
  assign n29631 = n20697 & n29535;
  assign n29632 = n17855 & ~n29516;
  assign n29633 = ~n29631 & ~n29632;
  assign n29634 = pi629 & ~n29633;
  assign n29635 = ~n29630 & ~n29634;
  assign n29636 = pi792 & ~n29635;
  assign n29637 = n20207 & ~n29636;
  assign n29638 = ~n29626 & n29637;
  assign n29639 = ~n29548 & ~n29638;
  assign n29640 = pi644 & n29639;
  assign n29641 = ~pi787 & ~n29536;
  assign n29642 = pi787 & ~n29545;
  assign n29643 = ~n29641 & ~n29642;
  assign n29644 = ~pi644 & n29643;
  assign n29645 = pi715 & ~n29644;
  assign n29646 = ~n29640 & n29645;
  assign n29647 = ~n17652 & ~n29519;
  assign n29648 = n17652 & n29482;
  assign n29649 = ~n29647 & ~n29648;
  assign n29650 = pi644 & ~n29649;
  assign n29651 = ~pi644 & n29482;
  assign n29652 = ~pi715 & ~n29651;
  assign n29653 = ~n29650 & n29652;
  assign n29654 = pi1160 & ~n29653;
  assign n29655 = ~n29646 & n29654;
  assign n29656 = ~pi644 & n29639;
  assign n29657 = pi644 & n29643;
  assign n29658 = ~pi715 & ~n29657;
  assign n29659 = ~n29656 & n29658;
  assign n29660 = ~pi644 & ~n29649;
  assign n29661 = pi644 & n29482;
  assign n29662 = pi715 & ~n29661;
  assign n29663 = ~n29660 & n29662;
  assign n29664 = ~pi1160 & ~n29663;
  assign n29665 = ~n29659 & n29664;
  assign n29666 = ~n29655 & ~n29665;
  assign n29667 = pi790 & ~n29666;
  assign n29668 = ~pi790 & n29639;
  assign n29669 = pi832 & ~n29668;
  assign n29670 = ~n29667 & n29669;
  assign po344 = ~n29481 & ~n29670;
  assign n29672 = pi188 & ~n3267;
  assign n29673 = ~pi768 & ~n19223;
  assign n29674 = ~n22171 & ~n29673;
  assign n29675 = ~pi188 & ~n29674;
  assign n29676 = ~pi188 & ~n19217;
  assign n29677 = ~pi768 & ~n29676;
  assign n29678 = ~n24271 & n29677;
  assign n29679 = ~n29675 & ~n29678;
  assign n29680 = ~pi705 & ~n29679;
  assign n29681 = ~pi188 & n19236;
  assign n29682 = pi188 & n19241;
  assign n29683 = pi768 & ~n19243;
  assign n29684 = ~n29682 & n29683;
  assign n29685 = ~n29681 & n29684;
  assign n29686 = pi188 & n19253;
  assign n29687 = ~pi188 & ~n19261;
  assign n29688 = ~pi768 & ~n29687;
  assign n29689 = ~n29686 & n29688;
  assign n29690 = pi705 & ~n29689;
  assign n29691 = ~n29685 & n29690;
  assign n29692 = n3267 & ~n29691;
  assign n29693 = ~n29680 & n29692;
  assign n29694 = ~n29672 & ~n29693;
  assign n29695 = ~pi625 & n29694;
  assign n29696 = n3267 & n29679;
  assign n29697 = ~n29672 & ~n29696;
  assign n29698 = pi625 & n29697;
  assign n29699 = ~pi1153 & ~n29698;
  assign n29700 = ~n29695 & n29699;
  assign n29701 = ~pi188 & n17972;
  assign n29702 = pi188 & ~n17976;
  assign n29703 = ~pi38 & ~n29702;
  assign n29704 = ~n29701 & n29703;
  assign n29705 = ~pi188 & ~n17280;
  assign n29706 = n17392 & ~n29705;
  assign n29707 = pi705 & ~n29706;
  assign n29708 = ~n29704 & n29707;
  assign n29709 = ~pi188 & ~pi705;
  assign n29710 = ~n17399 & n29709;
  assign n29711 = n3267 & ~n29710;
  assign n29712 = ~n29708 & n29711;
  assign n29713 = ~n29672 & ~n29712;
  assign n29714 = pi625 & n29713;
  assign n29715 = ~pi188 & ~n17406;
  assign n29716 = ~pi625 & n29715;
  assign n29717 = pi1153 & ~n29716;
  assign n29718 = ~n29714 & n29717;
  assign n29719 = ~pi608 & ~n29718;
  assign n29720 = ~n29700 & n29719;
  assign n29721 = pi625 & n29694;
  assign n29722 = ~pi625 & n29697;
  assign n29723 = pi1153 & ~n29722;
  assign n29724 = ~n29721 & n29723;
  assign n29725 = ~pi625 & n29713;
  assign n29726 = pi625 & n29715;
  assign n29727 = ~pi1153 & ~n29726;
  assign n29728 = ~n29725 & n29727;
  assign n29729 = pi608 & ~n29728;
  assign n29730 = ~n29724 & n29729;
  assign n29731 = ~n29720 & ~n29730;
  assign n29732 = pi778 & ~n29731;
  assign n29733 = ~pi778 & n29694;
  assign n29734 = ~n29732 & ~n29733;
  assign n29735 = ~pi609 & ~n29734;
  assign n29736 = ~pi778 & ~n29713;
  assign n29737 = ~n29718 & ~n29728;
  assign n29738 = pi778 & ~n29737;
  assign n29739 = ~n29736 & ~n29738;
  assign n29740 = pi609 & n29739;
  assign n29741 = ~pi1155 & ~n29740;
  assign n29742 = ~n29735 & n29741;
  assign n29743 = ~n17439 & ~n29715;
  assign n29744 = ~n17438 & ~n29697;
  assign n29745 = pi609 & n29744;
  assign n29746 = ~n29743 & ~n29745;
  assign n29747 = pi1155 & ~n29746;
  assign n29748 = ~pi660 & ~n29747;
  assign n29749 = ~n29742 & n29748;
  assign n29750 = pi609 & ~n29734;
  assign n29751 = ~pi609 & n29739;
  assign n29752 = pi1155 & ~n29751;
  assign n29753 = ~n29750 & n29752;
  assign n29754 = ~n17451 & ~n29715;
  assign n29755 = ~pi609 & n29744;
  assign n29756 = ~n29754 & ~n29755;
  assign n29757 = ~pi1155 & ~n29756;
  assign n29758 = pi660 & ~n29757;
  assign n29759 = ~n29753 & n29758;
  assign n29760 = ~n29749 & ~n29759;
  assign n29761 = pi785 & ~n29760;
  assign n29762 = ~pi785 & ~n29734;
  assign n29763 = ~n29761 & ~n29762;
  assign n29764 = ~pi618 & ~n29763;
  assign n29765 = ~n17466 & ~n29739;
  assign n29766 = n17466 & ~n29715;
  assign n29767 = ~n29765 & ~n29766;
  assign n29768 = pi618 & n29767;
  assign n29769 = ~pi1154 & ~n29768;
  assign n29770 = ~n29764 & n29769;
  assign n29771 = n17438 & ~n29715;
  assign n29772 = ~n29744 & ~n29771;
  assign n29773 = ~pi785 & ~n29772;
  assign n29774 = ~n29747 & ~n29757;
  assign n29775 = pi785 & ~n29774;
  assign n29776 = ~n29773 & ~n29775;
  assign n29777 = pi618 & n29776;
  assign n29778 = ~pi618 & n29715;
  assign n29779 = pi1154 & ~n29778;
  assign n29780 = ~n29777 & n29779;
  assign n29781 = ~pi627 & ~n29780;
  assign n29782 = ~n29770 & n29781;
  assign n29783 = pi618 & ~n29763;
  assign n29784 = ~pi618 & n29767;
  assign n29785 = pi1154 & ~n29784;
  assign n29786 = ~n29783 & n29785;
  assign n29787 = ~pi618 & n29776;
  assign n29788 = pi618 & n29715;
  assign n29789 = ~pi1154 & ~n29788;
  assign n29790 = ~n29787 & n29789;
  assign n29791 = pi627 & ~n29790;
  assign n29792 = ~n29786 & n29791;
  assign n29793 = ~n29782 & ~n29792;
  assign n29794 = pi781 & ~n29793;
  assign n29795 = ~pi781 & ~n29763;
  assign n29796 = ~n29794 & ~n29795;
  assign n29797 = ~pi619 & ~n29796;
  assign n29798 = ~n17503 & n29767;
  assign n29799 = n17503 & n29715;
  assign n29800 = ~n29798 & ~n29799;
  assign n29801 = pi619 & ~n29800;
  assign n29802 = ~pi1159 & ~n29801;
  assign n29803 = ~n29797 & n29802;
  assign n29804 = ~pi781 & ~n29776;
  assign n29805 = ~n29780 & ~n29790;
  assign n29806 = pi781 & ~n29805;
  assign n29807 = ~n29804 & ~n29806;
  assign n29808 = pi619 & n29807;
  assign n29809 = ~pi619 & n29715;
  assign n29810 = pi1159 & ~n29809;
  assign n29811 = ~n29808 & n29810;
  assign n29812 = ~pi648 & ~n29811;
  assign n29813 = ~n29803 & n29812;
  assign n29814 = pi619 & ~n29796;
  assign n29815 = ~pi619 & ~n29800;
  assign n29816 = pi1159 & ~n29815;
  assign n29817 = ~n29814 & n29816;
  assign n29818 = ~pi619 & n29807;
  assign n29819 = pi619 & n29715;
  assign n29820 = ~pi1159 & ~n29819;
  assign n29821 = ~n29818 & n29820;
  assign n29822 = pi648 & ~n29821;
  assign n29823 = ~n29817 & n29822;
  assign n29824 = ~n29813 & ~n29823;
  assign n29825 = pi789 & ~n29824;
  assign n29826 = ~pi789 & ~n29796;
  assign n29827 = ~n29825 & ~n29826;
  assign n29828 = ~pi788 & n29827;
  assign n29829 = ~pi626 & n29827;
  assign n29830 = n17539 & ~n29715;
  assign n29831 = ~n17539 & n29800;
  assign n29832 = ~n29830 & ~n29831;
  assign n29833 = pi626 & ~n29832;
  assign n29834 = ~pi641 & ~n29833;
  assign n29835 = ~n29829 & n29834;
  assign n29836 = ~pi789 & ~n29807;
  assign n29837 = ~n29811 & ~n29821;
  assign n29838 = pi789 & ~n29837;
  assign n29839 = ~n29836 & ~n29838;
  assign n29840 = ~pi626 & ~n29839;
  assign n29841 = pi626 & ~n29715;
  assign n29842 = pi641 & ~n29841;
  assign n29843 = ~n29840 & n29842;
  assign n29844 = ~pi1158 & ~n29843;
  assign n29845 = ~n29835 & n29844;
  assign n29846 = pi626 & n29827;
  assign n29847 = ~pi626 & ~n29832;
  assign n29848 = pi641 & ~n29847;
  assign n29849 = ~n29846 & n29848;
  assign n29850 = pi626 & ~n29839;
  assign n29851 = ~pi626 & ~n29715;
  assign n29852 = ~pi641 & ~n29851;
  assign n29853 = ~n29850 & n29852;
  assign n29854 = pi1158 & ~n29853;
  assign n29855 = ~n29849 & n29854;
  assign n29856 = ~n29845 & ~n29855;
  assign n29857 = pi788 & ~n29856;
  assign n29858 = ~n29828 & ~n29857;
  assign n29859 = ~pi628 & n29858;
  assign n29860 = ~n17816 & n29839;
  assign n29861 = n17816 & n29715;
  assign n29862 = ~n29860 & ~n29861;
  assign n29863 = pi628 & ~n29862;
  assign n29864 = ~pi1156 & ~n29863;
  assign n29865 = ~n29859 & n29864;
  assign n29866 = ~n17582 & n29832;
  assign n29867 = n17582 & n29715;
  assign n29868 = ~n29866 & ~n29867;
  assign n29869 = pi628 & ~n29868;
  assign n29870 = ~pi628 & n29715;
  assign n29871 = pi1156 & ~n29870;
  assign n29872 = ~n29869 & n29871;
  assign n29873 = ~pi629 & ~n29872;
  assign n29874 = ~n29865 & n29873;
  assign n29875 = pi628 & n29858;
  assign n29876 = ~pi628 & ~n29862;
  assign n29877 = pi1156 & ~n29876;
  assign n29878 = ~n29875 & n29877;
  assign n29879 = ~pi628 & ~n29868;
  assign n29880 = pi628 & n29715;
  assign n29881 = ~pi1156 & ~n29880;
  assign n29882 = ~n29879 & n29881;
  assign n29883 = pi629 & ~n29882;
  assign n29884 = ~n29878 & n29883;
  assign n29885 = ~n29874 & ~n29884;
  assign n29886 = pi792 & ~n29885;
  assign n29887 = ~pi792 & n29858;
  assign n29888 = ~n29886 & ~n29887;
  assign n29889 = ~pi647 & ~n29888;
  assign n29890 = ~n17610 & ~n29862;
  assign n29891 = n17610 & n29715;
  assign n29892 = ~n29890 & ~n29891;
  assign n29893 = pi647 & ~n29892;
  assign n29894 = ~pi1157 & ~n29893;
  assign n29895 = ~n29889 & n29894;
  assign n29896 = ~pi792 & n29868;
  assign n29897 = ~n29872 & ~n29882;
  assign n29898 = pi792 & ~n29897;
  assign n29899 = ~n29896 & ~n29898;
  assign n29900 = pi647 & n29899;
  assign n29901 = ~pi647 & n29715;
  assign n29902 = pi1157 & ~n29901;
  assign n29903 = ~n29900 & n29902;
  assign n29904 = ~pi630 & ~n29903;
  assign n29905 = ~n29895 & n29904;
  assign n29906 = pi647 & ~n29888;
  assign n29907 = ~pi647 & ~n29892;
  assign n29908 = pi1157 & ~n29907;
  assign n29909 = ~n29906 & n29908;
  assign n29910 = ~pi647 & n29899;
  assign n29911 = pi647 & n29715;
  assign n29912 = ~pi1157 & ~n29911;
  assign n29913 = ~n29910 & n29912;
  assign n29914 = pi630 & ~n29913;
  assign n29915 = ~n29909 & n29914;
  assign n29916 = ~n29905 & ~n29915;
  assign n29917 = pi787 & ~n29916;
  assign n29918 = ~pi787 & ~n29888;
  assign n29919 = ~n29917 & ~n29918;
  assign n29920 = ~pi644 & ~n29919;
  assign n29921 = ~pi787 & ~n29899;
  assign n29922 = ~n29903 & ~n29913;
  assign n29923 = pi787 & ~n29922;
  assign n29924 = ~n29921 & ~n29923;
  assign n29925 = pi644 & n29924;
  assign n29926 = ~pi715 & ~n29925;
  assign n29927 = ~n29920 & n29926;
  assign n29928 = n17652 & ~n29715;
  assign n29929 = ~n17652 & n29892;
  assign n29930 = ~n29928 & ~n29929;
  assign n29931 = ~pi644 & n29930;
  assign n29932 = pi644 & n29715;
  assign n29933 = pi715 & ~n29932;
  assign n29934 = ~n29931 & n29933;
  assign n29935 = ~pi1160 & ~n29934;
  assign n29936 = ~n29927 & n29935;
  assign n29937 = pi644 & ~n29919;
  assign n29938 = ~pi644 & n29924;
  assign n29939 = pi715 & ~n29938;
  assign n29940 = ~n29937 & n29939;
  assign n29941 = pi644 & n29930;
  assign n29942 = ~pi644 & n29715;
  assign n29943 = ~pi715 & ~n29942;
  assign n29944 = ~n29941 & n29943;
  assign n29945 = pi1160 & ~n29944;
  assign n29946 = ~n29940 & n29945;
  assign n29947 = pi790 & ~n29946;
  assign n29948 = ~n29936 & n29947;
  assign n29949 = ~pi790 & n29919;
  assign n29950 = ~po1038 & ~n29949;
  assign n29951 = ~n29948 & n29950;
  assign n29952 = ~pi188 & po1038;
  assign n29953 = ~pi832 & ~n29952;
  assign n29954 = ~n29951 & n29953;
  assign n29955 = ~pi188 & ~n2754;
  assign n29956 = ~pi768 & n16784;
  assign n29957 = ~n29955 & ~n29956;
  assign n29958 = ~n17706 & ~n29957;
  assign n29959 = ~pi785 & ~n29958;
  assign n29960 = ~n17711 & ~n29957;
  assign n29961 = pi1155 & ~n29960;
  assign n29962 = ~n17714 & n29958;
  assign n29963 = ~pi1155 & ~n29962;
  assign n29964 = ~n29961 & ~n29963;
  assign n29965 = pi785 & ~n29964;
  assign n29966 = ~n29959 & ~n29965;
  assign n29967 = ~pi781 & ~n29966;
  assign n29968 = ~n17721 & n29966;
  assign n29969 = pi1154 & ~n29968;
  assign n29970 = ~n17724 & n29966;
  assign n29971 = ~pi1154 & ~n29970;
  assign n29972 = ~n29969 & ~n29971;
  assign n29973 = pi781 & ~n29972;
  assign n29974 = ~n29967 & ~n29973;
  assign n29975 = ~pi789 & ~n29974;
  assign n29976 = pi619 & n29974;
  assign n29977 = ~pi619 & n29955;
  assign n29978 = pi1159 & ~n29977;
  assign n29979 = ~n29976 & n29978;
  assign n29980 = ~pi619 & n29974;
  assign n29981 = pi619 & n29955;
  assign n29982 = ~pi1159 & ~n29981;
  assign n29983 = ~n29980 & n29982;
  assign n29984 = ~n29979 & ~n29983;
  assign n29985 = pi789 & ~n29984;
  assign n29986 = ~n29975 & ~n29985;
  assign n29987 = ~n17816 & n29986;
  assign n29988 = n17816 & n29955;
  assign n29989 = ~n29987 & ~n29988;
  assign n29990 = ~n17610 & ~n29989;
  assign n29991 = n17610 & n29955;
  assign n29992 = ~n29990 & ~n29991;
  assign n29993 = ~n20398 & n29992;
  assign n29994 = pi705 & n16786;
  assign n29995 = ~n29955 & ~n29994;
  assign n29996 = ~pi778 & n29995;
  assign n29997 = ~pi625 & n29994;
  assign n29998 = ~n29995 & ~n29997;
  assign n29999 = pi1153 & ~n29998;
  assign n30000 = ~pi1153 & ~n29955;
  assign n30001 = ~n29997 & n30000;
  assign n30002 = ~n29999 & ~n30001;
  assign n30003 = pi778 & ~n30002;
  assign n30004 = ~n29996 & ~n30003;
  assign n30005 = ~n17692 & n30004;
  assign n30006 = ~n17694 & n30005;
  assign n30007 = ~n17696 & n30006;
  assign n30008 = ~n17828 & n30007;
  assign n30009 = ~n17859 & n30008;
  assign n30010 = ~pi647 & n30009;
  assign n30011 = pi647 & n29955;
  assign n30012 = ~pi1157 & ~n30011;
  assign n30013 = ~n30010 & n30012;
  assign n30014 = pi647 & ~n30009;
  assign n30015 = ~pi647 & ~n29955;
  assign n30016 = ~n30014 & ~n30015;
  assign n30017 = pi1157 & ~n30016;
  assign n30018 = ~n30013 & ~n30017;
  assign n30019 = ~n17651 & ~n30018;
  assign n30020 = ~n29993 & ~n30019;
  assign n30021 = pi787 & ~n30020;
  assign n30022 = pi626 & ~n29986;
  assign n30023 = ~pi626 & ~n29955;
  assign n30024 = n17579 & ~n30023;
  assign n30025 = ~n30022 & n30024;
  assign n30026 = n17704 & n30007;
  assign n30027 = ~pi626 & ~n29986;
  assign n30028 = pi626 & ~n29955;
  assign n30029 = n17580 & ~n30028;
  assign n30030 = ~n30027 & n30029;
  assign n30031 = ~n30026 & ~n30030;
  assign n30032 = ~n30025 & n30031;
  assign n30033 = pi788 & ~n30032;
  assign n30034 = ~n16521 & ~n29995;
  assign n30035 = pi625 & n30034;
  assign n30036 = n29957 & ~n30034;
  assign n30037 = ~n30035 & ~n30036;
  assign n30038 = n30000 & ~n30037;
  assign n30039 = ~pi608 & ~n29999;
  assign n30040 = ~n30038 & n30039;
  assign n30041 = pi1153 & n29957;
  assign n30042 = ~n30035 & n30041;
  assign n30043 = pi608 & ~n30001;
  assign n30044 = ~n30042 & n30043;
  assign n30045 = ~n30040 & ~n30044;
  assign n30046 = pi778 & ~n30045;
  assign n30047 = ~pi778 & ~n30036;
  assign n30048 = ~n30046 & ~n30047;
  assign n30049 = ~pi609 & ~n30048;
  assign n30050 = pi609 & n30004;
  assign n30051 = ~pi1155 & ~n30050;
  assign n30052 = ~n30049 & n30051;
  assign n30053 = ~pi660 & ~n29961;
  assign n30054 = ~n30052 & n30053;
  assign n30055 = pi609 & ~n30048;
  assign n30056 = ~pi609 & n30004;
  assign n30057 = pi1155 & ~n30056;
  assign n30058 = ~n30055 & n30057;
  assign n30059 = pi660 & ~n29963;
  assign n30060 = ~n30058 & n30059;
  assign n30061 = ~n30054 & ~n30060;
  assign n30062 = pi785 & ~n30061;
  assign n30063 = ~pi785 & ~n30048;
  assign n30064 = ~n30062 & ~n30063;
  assign n30065 = ~pi618 & ~n30064;
  assign n30066 = pi618 & n30005;
  assign n30067 = ~pi1154 & ~n30066;
  assign n30068 = ~n30065 & n30067;
  assign n30069 = ~pi627 & ~n29969;
  assign n30070 = ~n30068 & n30069;
  assign n30071 = pi618 & ~n30064;
  assign n30072 = ~pi618 & n30005;
  assign n30073 = pi1154 & ~n30072;
  assign n30074 = ~n30071 & n30073;
  assign n30075 = pi627 & ~n29971;
  assign n30076 = ~n30074 & n30075;
  assign n30077 = ~n30070 & ~n30076;
  assign n30078 = pi781 & ~n30077;
  assign n30079 = ~pi781 & ~n30064;
  assign n30080 = ~n30078 & ~n30079;
  assign n30081 = pi619 & ~n30080;
  assign n30082 = ~pi619 & n30006;
  assign n30083 = pi1159 & ~n30082;
  assign n30084 = ~n30081 & n30083;
  assign n30085 = pi648 & ~n29983;
  assign n30086 = ~n30084 & n30085;
  assign n30087 = ~pi619 & ~n30080;
  assign n30088 = pi619 & n30006;
  assign n30089 = ~pi1159 & ~n30088;
  assign n30090 = ~n30087 & n30089;
  assign n30091 = ~pi648 & ~n29979;
  assign n30092 = ~n30090 & n30091;
  assign n30093 = pi789 & ~n30092;
  assign n30094 = ~n30086 & n30093;
  assign n30095 = ~pi789 & n30080;
  assign n30096 = n17817 & ~n30095;
  assign n30097 = ~n30094 & n30096;
  assign n30098 = ~n30033 & ~n30097;
  assign n30099 = ~n20205 & ~n30098;
  assign n30100 = n17856 & ~n29989;
  assign n30101 = n20693 & n30008;
  assign n30102 = ~n30100 & ~n30101;
  assign n30103 = ~pi629 & ~n30102;
  assign n30104 = n20697 & n30008;
  assign n30105 = n17855 & ~n29989;
  assign n30106 = ~n30104 & ~n30105;
  assign n30107 = pi629 & ~n30106;
  assign n30108 = ~n30103 & ~n30107;
  assign n30109 = pi792 & ~n30108;
  assign n30110 = n20207 & ~n30109;
  assign n30111 = ~n30099 & n30110;
  assign n30112 = ~n30021 & ~n30111;
  assign n30113 = pi644 & n30112;
  assign n30114 = ~pi787 & ~n30009;
  assign n30115 = pi787 & ~n30018;
  assign n30116 = ~n30114 & ~n30115;
  assign n30117 = ~pi644 & n30116;
  assign n30118 = pi715 & ~n30117;
  assign n30119 = ~n30113 & n30118;
  assign n30120 = ~n17652 & ~n29992;
  assign n30121 = n17652 & n29955;
  assign n30122 = ~n30120 & ~n30121;
  assign n30123 = pi644 & ~n30122;
  assign n30124 = ~pi644 & n29955;
  assign n30125 = ~pi715 & ~n30124;
  assign n30126 = ~n30123 & n30125;
  assign n30127 = pi1160 & ~n30126;
  assign n30128 = ~n30119 & n30127;
  assign n30129 = ~pi644 & n30112;
  assign n30130 = pi644 & n30116;
  assign n30131 = ~pi715 & ~n30130;
  assign n30132 = ~n30129 & n30131;
  assign n30133 = ~pi644 & ~n30122;
  assign n30134 = pi644 & n29955;
  assign n30135 = pi715 & ~n30134;
  assign n30136 = ~n30133 & n30135;
  assign n30137 = ~pi1160 & ~n30136;
  assign n30138 = ~n30132 & n30137;
  assign n30139 = ~n30128 & ~n30138;
  assign n30140 = pi790 & ~n30139;
  assign n30141 = ~pi790 & n30112;
  assign n30142 = pi832 & ~n30141;
  assign n30143 = ~n30140 & n30142;
  assign po345 = ~n29954 & ~n30143;
  assign n30145 = pi189 & ~n3267;
  assign n30146 = pi189 & ~n16687;
  assign n30147 = ~pi189 & ~n16799;
  assign n30148 = ~pi772 & ~n30147;
  assign n30149 = ~n30146 & n30148;
  assign n30150 = ~pi189 & ~n16879;
  assign n30151 = pi189 & n16944;
  assign n30152 = pi772 & ~n30151;
  assign n30153 = ~n30150 & n30152;
  assign n30154 = pi39 & ~n30153;
  assign n30155 = ~n30149 & n30154;
  assign n30156 = pi189 & ~n17088;
  assign n30157 = ~pi189 & ~n17059;
  assign n30158 = ~pi772 & ~n30157;
  assign n30159 = ~n30156 & n30158;
  assign n30160 = pi189 & n17092;
  assign n30161 = ~pi189 & n17094;
  assign n30162 = pi772 & ~n30161;
  assign n30163 = ~n30160 & n30162;
  assign n30164 = ~pi39 & ~n30163;
  assign n30165 = ~n30159 & n30164;
  assign n30166 = ~pi38 & ~n30165;
  assign n30167 = ~n30155 & n30166;
  assign n30168 = pi772 & n16521;
  assign n30169 = n17280 & ~n30168;
  assign n30170 = ~pi189 & ~n17280;
  assign n30171 = pi38 & ~n30170;
  assign n30172 = ~n30169 & n30171;
  assign n30173 = pi727 & ~n19243;
  assign n30174 = ~n30172 & n30173;
  assign n30175 = ~n30167 & n30174;
  assign n30176 = pi772 & n17240;
  assign n30177 = ~n22064 & ~n30176;
  assign n30178 = pi39 & ~n30177;
  assign n30179 = pi772 & n17042;
  assign n30180 = ~pi772 & n17120;
  assign n30181 = ~pi39 & ~n30180;
  assign n30182 = ~n30179 & n30181;
  assign n30183 = ~n30178 & ~n30182;
  assign n30184 = pi189 & ~n30183;
  assign n30185 = ~pi189 & pi772;
  assign n30186 = n17275 & n30185;
  assign n30187 = ~n30184 & ~n30186;
  assign n30188 = ~pi38 & ~n30187;
  assign n30189 = ~n30172 & ~n30188;
  assign n30190 = n3267 & ~n30189;
  assign n30191 = pi727 & n3267;
  assign n30192 = ~n30190 & ~n30191;
  assign n30193 = ~n30175 & ~n30192;
  assign n30194 = ~n30145 & ~n30193;
  assign n30195 = ~pi625 & n30194;
  assign n30196 = ~n30145 & ~n30190;
  assign n30197 = pi625 & n30196;
  assign n30198 = ~pi1153 & ~n30197;
  assign n30199 = ~n30195 & n30198;
  assign n30200 = pi189 & ~n17406;
  assign n30201 = ~n30191 & ~n30200;
  assign n30202 = pi189 & ~n17972;
  assign n30203 = ~pi189 & n17976;
  assign n30204 = ~pi38 & ~n30203;
  assign n30205 = ~n30202 & n30204;
  assign n30206 = n19802 & ~n30170;
  assign n30207 = n30191 & ~n30206;
  assign n30208 = ~n30205 & n30207;
  assign n30209 = ~n30201 & ~n30208;
  assign n30210 = pi625 & ~n30209;
  assign n30211 = ~pi625 & ~n30200;
  assign n30212 = pi1153 & ~n30211;
  assign n30213 = ~n30210 & n30212;
  assign n30214 = ~pi608 & ~n30213;
  assign n30215 = ~n30199 & n30214;
  assign n30216 = pi625 & n30194;
  assign n30217 = ~pi625 & n30196;
  assign n30218 = pi1153 & ~n30217;
  assign n30219 = ~n30216 & n30218;
  assign n30220 = ~pi625 & ~n30209;
  assign n30221 = pi625 & ~n30200;
  assign n30222 = ~pi1153 & ~n30221;
  assign n30223 = ~n30220 & n30222;
  assign n30224 = pi608 & ~n30223;
  assign n30225 = ~n30219 & n30224;
  assign n30226 = ~n30215 & ~n30225;
  assign n30227 = pi778 & ~n30226;
  assign n30228 = ~pi778 & n30194;
  assign n30229 = ~n30227 & ~n30228;
  assign n30230 = ~pi609 & ~n30229;
  assign n30231 = ~pi778 & n30209;
  assign n30232 = ~n30213 & ~n30223;
  assign n30233 = pi778 & ~n30232;
  assign n30234 = ~n30231 & ~n30233;
  assign n30235 = pi609 & n30234;
  assign n30236 = ~pi1155 & ~n30235;
  assign n30237 = ~n30230 & n30236;
  assign n30238 = n17438 & ~n30200;
  assign n30239 = ~n17438 & n30196;
  assign n30240 = ~n30238 & ~n30239;
  assign n30241 = pi609 & ~n30240;
  assign n30242 = ~pi609 & ~n30200;
  assign n30243 = pi1155 & ~n30242;
  assign n30244 = ~n30241 & n30243;
  assign n30245 = ~pi660 & ~n30244;
  assign n30246 = ~n30237 & n30245;
  assign n30247 = pi609 & ~n30229;
  assign n30248 = ~pi609 & n30234;
  assign n30249 = pi1155 & ~n30248;
  assign n30250 = ~n30247 & n30249;
  assign n30251 = ~pi609 & ~n30240;
  assign n30252 = pi609 & ~n30200;
  assign n30253 = ~pi1155 & ~n30252;
  assign n30254 = ~n30251 & n30253;
  assign n30255 = pi660 & ~n30254;
  assign n30256 = ~n30250 & n30255;
  assign n30257 = ~n30246 & ~n30256;
  assign n30258 = pi785 & ~n30257;
  assign n30259 = ~pi785 & ~n30229;
  assign n30260 = ~n30258 & ~n30259;
  assign n30261 = ~pi618 & ~n30260;
  assign n30262 = n17466 & ~n30200;
  assign n30263 = ~n17466 & n30234;
  assign n30264 = ~n30262 & ~n30263;
  assign n30265 = pi618 & ~n30264;
  assign n30266 = ~pi1154 & ~n30265;
  assign n30267 = ~n30261 & n30266;
  assign n30268 = ~pi785 & n30240;
  assign n30269 = ~n30244 & ~n30254;
  assign n30270 = pi785 & ~n30269;
  assign n30271 = ~n30268 & ~n30270;
  assign n30272 = pi618 & n30271;
  assign n30273 = ~pi618 & ~n30200;
  assign n30274 = pi1154 & ~n30273;
  assign n30275 = ~n30272 & n30274;
  assign n30276 = ~pi627 & ~n30275;
  assign n30277 = ~n30267 & n30276;
  assign n30278 = pi618 & ~n30260;
  assign n30279 = ~pi618 & ~n30264;
  assign n30280 = pi1154 & ~n30279;
  assign n30281 = ~n30278 & n30280;
  assign n30282 = ~pi618 & n30271;
  assign n30283 = pi618 & ~n30200;
  assign n30284 = ~pi1154 & ~n30283;
  assign n30285 = ~n30282 & n30284;
  assign n30286 = pi627 & ~n30285;
  assign n30287 = ~n30281 & n30286;
  assign n30288 = ~n30277 & ~n30287;
  assign n30289 = pi781 & ~n30288;
  assign n30290 = ~pi781 & ~n30260;
  assign n30291 = ~n30289 & ~n30290;
  assign n30292 = ~pi619 & ~n30291;
  assign n30293 = ~n17503 & n30264;
  assign n30294 = n17503 & n30200;
  assign n30295 = ~n30293 & ~n30294;
  assign n30296 = pi619 & n30295;
  assign n30297 = ~pi1159 & ~n30296;
  assign n30298 = ~n30292 & n30297;
  assign n30299 = ~pi781 & ~n30271;
  assign n30300 = ~n30275 & ~n30285;
  assign n30301 = pi781 & ~n30300;
  assign n30302 = ~n30299 & ~n30301;
  assign n30303 = pi619 & n30302;
  assign n30304 = ~pi619 & ~n30200;
  assign n30305 = pi1159 & ~n30304;
  assign n30306 = ~n30303 & n30305;
  assign n30307 = ~pi648 & ~n30306;
  assign n30308 = ~n30298 & n30307;
  assign n30309 = pi619 & ~n30291;
  assign n30310 = ~pi619 & n30295;
  assign n30311 = pi1159 & ~n30310;
  assign n30312 = ~n30309 & n30311;
  assign n30313 = ~pi619 & n30302;
  assign n30314 = pi619 & ~n30200;
  assign n30315 = ~pi1159 & ~n30314;
  assign n30316 = ~n30313 & n30315;
  assign n30317 = pi648 & ~n30316;
  assign n30318 = ~n30312 & n30317;
  assign n30319 = ~n30308 & ~n30318;
  assign n30320 = pi789 & ~n30319;
  assign n30321 = ~pi789 & ~n30291;
  assign n30322 = ~n30320 & ~n30321;
  assign n30323 = ~pi788 & n30322;
  assign n30324 = ~pi626 & n30322;
  assign n30325 = n17539 & ~n30200;
  assign n30326 = ~n17539 & n30295;
  assign n30327 = ~n30325 & ~n30326;
  assign n30328 = pi626 & n30327;
  assign n30329 = ~pi641 & ~n30328;
  assign n30330 = ~n30324 & n30329;
  assign n30331 = ~pi789 & ~n30302;
  assign n30332 = ~n30306 & ~n30316;
  assign n30333 = pi789 & ~n30332;
  assign n30334 = ~n30331 & ~n30333;
  assign n30335 = ~pi626 & ~n30334;
  assign n30336 = pi626 & n30200;
  assign n30337 = pi641 & ~n30336;
  assign n30338 = ~n30335 & n30337;
  assign n30339 = ~pi1158 & ~n30338;
  assign n30340 = ~n30330 & n30339;
  assign n30341 = pi626 & n30322;
  assign n30342 = ~pi626 & n30327;
  assign n30343 = pi641 & ~n30342;
  assign n30344 = ~n30341 & n30343;
  assign n30345 = pi626 & ~n30334;
  assign n30346 = ~pi626 & n30200;
  assign n30347 = ~pi641 & ~n30346;
  assign n30348 = ~n30345 & n30347;
  assign n30349 = pi1158 & ~n30348;
  assign n30350 = ~n30344 & n30349;
  assign n30351 = ~n30340 & ~n30350;
  assign n30352 = pi788 & ~n30351;
  assign n30353 = ~n30323 & ~n30352;
  assign n30354 = ~pi628 & n30353;
  assign n30355 = ~n17816 & ~n30334;
  assign n30356 = n17816 & n30200;
  assign n30357 = ~n30355 & ~n30356;
  assign n30358 = pi628 & n30357;
  assign n30359 = ~pi1156 & ~n30358;
  assign n30360 = ~n30354 & n30359;
  assign n30361 = ~n17582 & n30327;
  assign n30362 = n17582 & n30200;
  assign n30363 = ~n30361 & ~n30362;
  assign n30364 = pi628 & n30363;
  assign n30365 = ~pi628 & ~n30200;
  assign n30366 = pi1156 & ~n30365;
  assign n30367 = ~n30364 & n30366;
  assign n30368 = ~pi629 & ~n30367;
  assign n30369 = ~n30360 & n30368;
  assign n30370 = pi628 & n30353;
  assign n30371 = ~pi628 & n30357;
  assign n30372 = pi1156 & ~n30371;
  assign n30373 = ~n30370 & n30372;
  assign n30374 = ~pi628 & n30363;
  assign n30375 = pi628 & ~n30200;
  assign n30376 = ~pi1156 & ~n30375;
  assign n30377 = ~n30374 & n30376;
  assign n30378 = pi629 & ~n30377;
  assign n30379 = ~n30373 & n30378;
  assign n30380 = ~n30369 & ~n30379;
  assign n30381 = pi792 & ~n30380;
  assign n30382 = ~pi792 & n30353;
  assign n30383 = ~n30381 & ~n30382;
  assign n30384 = ~pi647 & ~n30383;
  assign n30385 = ~n17610 & ~n30357;
  assign n30386 = n17610 & n30200;
  assign n30387 = ~n30385 & ~n30386;
  assign n30388 = pi647 & n30387;
  assign n30389 = ~pi1157 & ~n30388;
  assign n30390 = ~n30384 & n30389;
  assign n30391 = ~pi792 & ~n30363;
  assign n30392 = ~n30367 & ~n30377;
  assign n30393 = pi792 & ~n30392;
  assign n30394 = ~n30391 & ~n30393;
  assign n30395 = pi647 & n30394;
  assign n30396 = ~pi647 & ~n30200;
  assign n30397 = pi1157 & ~n30396;
  assign n30398 = ~n30395 & n30397;
  assign n30399 = ~pi630 & ~n30398;
  assign n30400 = ~n30390 & n30399;
  assign n30401 = pi647 & ~n30383;
  assign n30402 = ~pi647 & n30387;
  assign n30403 = pi1157 & ~n30402;
  assign n30404 = ~n30401 & n30403;
  assign n30405 = ~pi647 & n30394;
  assign n30406 = pi647 & ~n30200;
  assign n30407 = ~pi1157 & ~n30406;
  assign n30408 = ~n30405 & n30407;
  assign n30409 = pi630 & ~n30408;
  assign n30410 = ~n30404 & n30409;
  assign n30411 = ~n30400 & ~n30410;
  assign n30412 = pi787 & ~n30411;
  assign n30413 = ~pi787 & ~n30383;
  assign n30414 = ~n30412 & ~n30413;
  assign n30415 = ~pi644 & ~n30414;
  assign n30416 = ~pi787 & ~n30394;
  assign n30417 = ~n30398 & ~n30408;
  assign n30418 = pi787 & ~n30417;
  assign n30419 = ~n30416 & ~n30418;
  assign n30420 = pi644 & n30419;
  assign n30421 = ~pi715 & ~n30420;
  assign n30422 = ~n30415 & n30421;
  assign n30423 = n17652 & ~n30200;
  assign n30424 = ~n17652 & n30387;
  assign n30425 = ~n30423 & ~n30424;
  assign n30426 = ~pi644 & ~n30425;
  assign n30427 = pi644 & ~n30200;
  assign n30428 = pi715 & ~n30427;
  assign n30429 = ~n30426 & n30428;
  assign n30430 = ~pi1160 & ~n30429;
  assign n30431 = ~n30422 & n30430;
  assign n30432 = pi644 & ~n30414;
  assign n30433 = ~pi644 & n30419;
  assign n30434 = pi715 & ~n30433;
  assign n30435 = ~n30432 & n30434;
  assign n30436 = pi644 & ~n30425;
  assign n30437 = ~pi644 & ~n30200;
  assign n30438 = ~pi715 & ~n30437;
  assign n30439 = ~n30436 & n30438;
  assign n30440 = pi1160 & ~n30439;
  assign n30441 = ~n30435 & n30440;
  assign n30442 = pi790 & ~n30441;
  assign n30443 = ~n30431 & n30442;
  assign n30444 = ~pi790 & n30414;
  assign n30445 = n6286 & ~n30444;
  assign n30446 = ~n30443 & n30445;
  assign n30447 = ~pi189 & ~n6286;
  assign n30448 = ~pi57 & ~n30447;
  assign n30449 = ~n30446 & n30448;
  assign n30450 = pi57 & pi189;
  assign n30451 = ~pi832 & ~n30450;
  assign n30452 = ~n30449 & n30451;
  assign n30453 = pi189 & ~n2754;
  assign n30454 = pi772 & n16784;
  assign n30455 = ~n30453 & ~n30454;
  assign n30456 = pi727 & n16787;
  assign n30457 = n30455 & ~n30456;
  assign n30458 = pi625 & n30456;
  assign n30459 = ~n30457 & ~n30458;
  assign n30460 = ~pi1153 & ~n30459;
  assign n30461 = pi727 & n16786;
  assign n30462 = pi625 & n30461;
  assign n30463 = pi1153 & ~n30453;
  assign n30464 = ~n30462 & n30463;
  assign n30465 = ~pi608 & ~n30464;
  assign n30466 = ~n30460 & n30465;
  assign n30467 = pi1153 & n30455;
  assign n30468 = ~n30458 & n30467;
  assign n30469 = ~n30453 & ~n30461;
  assign n30470 = ~n30462 & ~n30469;
  assign n30471 = ~pi1153 & ~n30470;
  assign n30472 = pi608 & ~n30471;
  assign n30473 = ~n30468 & n30472;
  assign n30474 = ~n30466 & ~n30473;
  assign n30475 = pi778 & ~n30474;
  assign n30476 = ~pi778 & ~n30457;
  assign n30477 = ~n30475 & ~n30476;
  assign n30478 = ~pi609 & ~n30477;
  assign n30479 = ~pi778 & n30469;
  assign n30480 = ~n30464 & ~n30471;
  assign n30481 = pi778 & ~n30480;
  assign n30482 = ~n30479 & ~n30481;
  assign n30483 = pi609 & n30482;
  assign n30484 = ~pi1155 & ~n30483;
  assign n30485 = ~n30478 & n30484;
  assign n30486 = n17439 & n30454;
  assign n30487 = pi1155 & ~n30453;
  assign n30488 = ~n30486 & n30487;
  assign n30489 = ~pi660 & ~n30488;
  assign n30490 = ~n30485 & n30489;
  assign n30491 = pi609 & ~n30477;
  assign n30492 = ~pi609 & n30482;
  assign n30493 = pi1155 & ~n30492;
  assign n30494 = ~n30491 & n30493;
  assign n30495 = n17451 & n30454;
  assign n30496 = ~pi1155 & ~n30453;
  assign n30497 = ~n30495 & n30496;
  assign n30498 = pi660 & ~n30497;
  assign n30499 = ~n30494 & n30498;
  assign n30500 = ~n30490 & ~n30499;
  assign n30501 = pi785 & ~n30500;
  assign n30502 = ~pi785 & ~n30477;
  assign n30503 = ~n30501 & ~n30502;
  assign n30504 = pi618 & ~n30503;
  assign n30505 = ~n17692 & n30482;
  assign n30506 = ~pi618 & n30505;
  assign n30507 = pi1154 & ~n30506;
  assign n30508 = ~n30504 & n30507;
  assign n30509 = ~n20069 & n30454;
  assign n30510 = n20164 & n30509;
  assign n30511 = ~pi1154 & ~n30453;
  assign n30512 = ~n30510 & n30511;
  assign n30513 = pi627 & ~n30512;
  assign n30514 = ~n30508 & n30513;
  assign n30515 = ~pi618 & ~n30503;
  assign n30516 = pi618 & n30505;
  assign n30517 = ~pi1154 & ~n30516;
  assign n30518 = ~n30515 & n30517;
  assign n30519 = n20154 & n30509;
  assign n30520 = pi1154 & ~n30453;
  assign n30521 = ~n30519 & n30520;
  assign n30522 = ~pi627 & ~n30521;
  assign n30523 = ~n30518 & n30522;
  assign n30524 = ~n30514 & ~n30523;
  assign n30525 = pi781 & ~n30524;
  assign n30526 = ~pi781 & ~n30503;
  assign n30527 = ~n23444 & ~n30526;
  assign n30528 = ~n30525 & n30527;
  assign n30529 = n19127 & n30482;
  assign n30530 = ~n23442 & ~n30529;
  assign n30531 = ~n20075 & n30509;
  assign n30532 = n20179 & n30531;
  assign n30533 = n17537 & ~n30532;
  assign n30534 = n20189 & n30531;
  assign n30535 = n17536 & ~n30534;
  assign n30536 = ~n30533 & ~n30535;
  assign n30537 = ~n30530 & n30536;
  assign n30538 = pi789 & ~n30453;
  assign n30539 = ~n30537 & n30538;
  assign n30540 = n17817 & ~n30539;
  assign n30541 = ~n30528 & n30540;
  assign n30542 = ~n17539 & n30529;
  assign n30543 = ~n30453 & ~n30542;
  assign n30544 = n17699 & ~n30543;
  assign n30545 = n20081 & n30509;
  assign n30546 = pi626 & n30545;
  assign n30547 = ~n30453 & ~n30546;
  assign n30548 = pi1158 & ~n30547;
  assign n30549 = ~pi641 & ~n30548;
  assign n30550 = ~n30544 & n30549;
  assign n30551 = n17698 & ~n30543;
  assign n30552 = ~pi626 & n30545;
  assign n30553 = ~n30453 & ~n30552;
  assign n30554 = ~pi1158 & ~n30553;
  assign n30555 = pi641 & ~n30554;
  assign n30556 = ~n30551 & n30555;
  assign n30557 = pi788 & ~n30556;
  assign n30558 = ~n30550 & n30557;
  assign n30559 = ~n20205 & ~n30558;
  assign n30560 = ~n30541 & n30559;
  assign n30561 = ~n17816 & n30545;
  assign n30562 = ~pi629 & n30561;
  assign n30563 = pi628 & ~n30562;
  assign n30564 = n19128 & n30482;
  assign n30565 = pi629 & ~n30564;
  assign n30566 = ~n30563 & ~n30565;
  assign n30567 = ~pi1156 & ~n30566;
  assign n30568 = pi628 & n30564;
  assign n30569 = ~pi628 & ~n30561;
  assign n30570 = pi629 & ~n30569;
  assign n30571 = pi1156 & ~n30570;
  assign n30572 = ~n30568 & n30571;
  assign n30573 = ~n30567 & ~n30572;
  assign n30574 = pi792 & ~n30453;
  assign n30575 = ~n30573 & n30574;
  assign n30576 = ~n30560 & ~n30575;
  assign n30577 = n20207 & ~n30576;
  assign n30578 = ~n17610 & n30561;
  assign n30579 = ~pi630 & n30578;
  assign n30580 = pi647 & ~n30579;
  assign n30581 = ~n19158 & n30564;
  assign n30582 = pi630 & ~n30581;
  assign n30583 = ~n30580 & ~n30582;
  assign n30584 = ~pi1157 & ~n30583;
  assign n30585 = ~pi630 & ~n30581;
  assign n30586 = pi647 & ~n30585;
  assign n30587 = pi630 & n30578;
  assign n30588 = pi1157 & ~n30587;
  assign n30589 = ~n30586 & n30588;
  assign n30590 = ~n30584 & ~n30589;
  assign n30591 = pi787 & ~n30453;
  assign n30592 = ~n30590 & n30591;
  assign n30593 = ~n30577 & ~n30592;
  assign n30594 = pi644 & n30593;
  assign n30595 = ~n19182 & n30581;
  assign n30596 = ~n30453 & ~n30595;
  assign n30597 = ~pi644 & ~n30596;
  assign n30598 = pi715 & ~n30597;
  assign n30599 = ~n30594 & n30598;
  assign n30600 = ~n17816 & n23518;
  assign n30601 = n30545 & n30600;
  assign n30602 = pi644 & n30601;
  assign n30603 = ~pi715 & ~n30453;
  assign n30604 = ~n30602 & n30603;
  assign n30605 = pi1160 & ~n30604;
  assign n30606 = ~n30599 & n30605;
  assign n30607 = ~pi644 & n30593;
  assign n30608 = pi644 & ~n30596;
  assign n30609 = ~pi715 & ~n30608;
  assign n30610 = ~n30607 & n30609;
  assign n30611 = ~pi644 & n30601;
  assign n30612 = pi715 & ~n30453;
  assign n30613 = ~n30611 & n30612;
  assign n30614 = ~pi1160 & ~n30613;
  assign n30615 = ~n30610 & n30614;
  assign n30616 = ~n30606 & ~n30615;
  assign n30617 = pi790 & ~n30616;
  assign n30618 = ~pi790 & n30593;
  assign n30619 = pi832 & ~n30618;
  assign n30620 = ~n30617 & n30619;
  assign po346 = ~n30452 & ~n30620;
  assign n30622 = ~pi190 & ~n2754;
  assign n30623 = pi763 & n16784;
  assign n30624 = ~n30622 & ~n30623;
  assign n30625 = ~n17706 & ~n30624;
  assign n30626 = ~pi785 & ~n30625;
  assign n30627 = n17451 & n30623;
  assign n30628 = n30625 & ~n30627;
  assign n30629 = pi1155 & ~n30628;
  assign n30630 = ~pi1155 & ~n30622;
  assign n30631 = ~n30627 & n30630;
  assign n30632 = ~n30629 & ~n30631;
  assign n30633 = pi785 & ~n30632;
  assign n30634 = ~n30626 & ~n30633;
  assign n30635 = ~pi781 & ~n30634;
  assign n30636 = ~n17721 & n30634;
  assign n30637 = pi1154 & ~n30636;
  assign n30638 = ~n17724 & n30634;
  assign n30639 = ~pi1154 & ~n30638;
  assign n30640 = ~n30637 & ~n30639;
  assign n30641 = pi781 & ~n30640;
  assign n30642 = ~n30635 & ~n30641;
  assign n30643 = ~pi789 & ~n30642;
  assign n30644 = ~n22890 & n30642;
  assign n30645 = pi1159 & ~n30644;
  assign n30646 = ~n22893 & n30642;
  assign n30647 = ~pi1159 & ~n30646;
  assign n30648 = ~n30645 & ~n30647;
  assign n30649 = pi789 & ~n30648;
  assign n30650 = ~n30643 & ~n30649;
  assign n30651 = ~n17816 & n30650;
  assign n30652 = n17816 & n30622;
  assign n30653 = ~n30651 & ~n30652;
  assign n30654 = ~n17610 & ~n30653;
  assign n30655 = n17610 & n30622;
  assign n30656 = ~n30654 & ~n30655;
  assign n30657 = ~n20398 & n30656;
  assign n30658 = pi699 & n16786;
  assign n30659 = ~n30622 & ~n30658;
  assign n30660 = ~pi778 & ~n30659;
  assign n30661 = ~pi625 & n30658;
  assign n30662 = ~n30659 & ~n30661;
  assign n30663 = pi1153 & ~n30662;
  assign n30664 = ~pi1153 & ~n30622;
  assign n30665 = ~n30661 & n30664;
  assign n30666 = pi778 & ~n30665;
  assign n30667 = ~n30663 & n30666;
  assign n30668 = ~n30660 & ~n30667;
  assign n30669 = ~n17692 & ~n30668;
  assign n30670 = ~n17694 & n30669;
  assign n30671 = ~n17696 & n30670;
  assign n30672 = ~n17828 & n30671;
  assign n30673 = ~n17859 & n30672;
  assign n30674 = ~pi647 & n30673;
  assign n30675 = pi647 & n30622;
  assign n30676 = ~pi1157 & ~n30675;
  assign n30677 = ~n30674 & n30676;
  assign n30678 = pi647 & ~n30673;
  assign n30679 = ~pi647 & ~n30622;
  assign n30680 = ~n30678 & ~n30679;
  assign n30681 = pi1157 & ~n30680;
  assign n30682 = ~n30677 & ~n30681;
  assign n30683 = ~n17651 & ~n30682;
  assign n30684 = ~n30657 & ~n30683;
  assign n30685 = pi787 & ~n30684;
  assign n30686 = pi626 & ~n30650;
  assign n30687 = ~pi626 & ~n30622;
  assign n30688 = n17579 & ~n30687;
  assign n30689 = ~n30686 & n30688;
  assign n30690 = n17704 & n30671;
  assign n30691 = ~pi626 & ~n30650;
  assign n30692 = pi626 & ~n30622;
  assign n30693 = n17580 & ~n30692;
  assign n30694 = ~n30691 & n30693;
  assign n30695 = ~n30690 & ~n30694;
  assign n30696 = ~n30689 & n30695;
  assign n30697 = pi788 & ~n30696;
  assign n30698 = ~n16521 & ~n30659;
  assign n30699 = pi625 & n30698;
  assign n30700 = n30624 & ~n30698;
  assign n30701 = ~n30699 & ~n30700;
  assign n30702 = n30664 & ~n30701;
  assign n30703 = ~pi608 & ~n30663;
  assign n30704 = ~n30702 & n30703;
  assign n30705 = pi1153 & n30624;
  assign n30706 = ~n30699 & n30705;
  assign n30707 = pi608 & ~n30665;
  assign n30708 = ~n30706 & n30707;
  assign n30709 = ~n30704 & ~n30708;
  assign n30710 = pi778 & ~n30709;
  assign n30711 = ~pi778 & ~n30700;
  assign n30712 = ~n30710 & ~n30711;
  assign n30713 = ~pi609 & ~n30712;
  assign n30714 = pi609 & ~n30668;
  assign n30715 = ~pi1155 & ~n30714;
  assign n30716 = ~n30713 & n30715;
  assign n30717 = ~pi660 & ~n30629;
  assign n30718 = ~n30716 & n30717;
  assign n30719 = pi609 & ~n30712;
  assign n30720 = ~pi609 & ~n30668;
  assign n30721 = pi1155 & ~n30720;
  assign n30722 = ~n30719 & n30721;
  assign n30723 = pi660 & ~n30631;
  assign n30724 = ~n30722 & n30723;
  assign n30725 = ~n30718 & ~n30724;
  assign n30726 = pi785 & ~n30725;
  assign n30727 = ~pi785 & ~n30712;
  assign n30728 = ~n30726 & ~n30727;
  assign n30729 = ~pi618 & ~n30728;
  assign n30730 = pi618 & n30669;
  assign n30731 = ~pi1154 & ~n30730;
  assign n30732 = ~n30729 & n30731;
  assign n30733 = ~pi627 & ~n30637;
  assign n30734 = ~n30732 & n30733;
  assign n30735 = pi618 & ~n30728;
  assign n30736 = ~pi618 & n30669;
  assign n30737 = pi1154 & ~n30736;
  assign n30738 = ~n30735 & n30737;
  assign n30739 = pi627 & ~n30639;
  assign n30740 = ~n30738 & n30739;
  assign n30741 = ~n30734 & ~n30740;
  assign n30742 = pi781 & ~n30741;
  assign n30743 = ~pi781 & ~n30728;
  assign n30744 = ~n30742 & ~n30743;
  assign n30745 = pi619 & ~n30744;
  assign n30746 = ~pi619 & n30670;
  assign n30747 = pi1159 & ~n30746;
  assign n30748 = ~n30745 & n30747;
  assign n30749 = pi648 & ~n30647;
  assign n30750 = ~n30748 & n30749;
  assign n30751 = ~pi619 & ~n30744;
  assign n30752 = pi619 & n30670;
  assign n30753 = ~pi1159 & ~n30752;
  assign n30754 = ~n30751 & n30753;
  assign n30755 = ~pi648 & ~n30645;
  assign n30756 = ~n30754 & n30755;
  assign n30757 = pi789 & ~n30756;
  assign n30758 = ~n30750 & n30757;
  assign n30759 = ~pi789 & n30744;
  assign n30760 = n17817 & ~n30759;
  assign n30761 = ~n30758 & n30760;
  assign n30762 = ~n30697 & ~n30761;
  assign n30763 = ~n20205 & ~n30762;
  assign n30764 = n17856 & ~n30653;
  assign n30765 = n20693 & n30672;
  assign n30766 = ~n30764 & ~n30765;
  assign n30767 = ~pi629 & ~n30766;
  assign n30768 = n20697 & n30672;
  assign n30769 = n17855 & ~n30653;
  assign n30770 = ~n30768 & ~n30769;
  assign n30771 = pi629 & ~n30770;
  assign n30772 = ~n30767 & ~n30771;
  assign n30773 = pi792 & ~n30772;
  assign n30774 = n20207 & ~n30773;
  assign n30775 = ~n30763 & n30774;
  assign n30776 = ~n30685 & ~n30775;
  assign n30777 = pi644 & n30776;
  assign n30778 = ~pi787 & ~n30673;
  assign n30779 = pi787 & ~n30682;
  assign n30780 = ~n30778 & ~n30779;
  assign n30781 = ~pi644 & n30780;
  assign n30782 = pi715 & ~n30781;
  assign n30783 = ~n30777 & n30782;
  assign n30784 = ~n17652 & ~n30656;
  assign n30785 = n17652 & n30622;
  assign n30786 = ~n30784 & ~n30785;
  assign n30787 = pi644 & ~n30786;
  assign n30788 = ~pi644 & n30622;
  assign n30789 = ~pi715 & ~n30788;
  assign n30790 = ~n30787 & n30789;
  assign n30791 = pi1160 & ~n30790;
  assign n30792 = ~n30783 & n30791;
  assign n30793 = ~pi644 & n30776;
  assign n30794 = pi644 & n30780;
  assign n30795 = ~pi715 & ~n30794;
  assign n30796 = ~n30793 & n30795;
  assign n30797 = ~pi644 & ~n30786;
  assign n30798 = pi644 & n30622;
  assign n30799 = pi715 & ~n30798;
  assign n30800 = ~n30797 & n30799;
  assign n30801 = ~pi1160 & ~n30800;
  assign n30802 = ~n30796 & n30801;
  assign n30803 = ~n30792 & ~n30802;
  assign n30804 = pi790 & ~n30803;
  assign n30805 = ~pi790 & n30776;
  assign n30806 = pi832 & ~n30805;
  assign n30807 = ~n30804 & n30806;
  assign n30808 = ~pi190 & ~n17406;
  assign n30809 = n17539 & ~n30808;
  assign n30810 = pi190 & ~n3267;
  assign n30811 = ~pi190 & n17972;
  assign n30812 = pi190 & ~n17976;
  assign n30813 = ~pi38 & ~n30812;
  assign n30814 = ~n30811 & n30813;
  assign n30815 = ~pi190 & ~n17280;
  assign n30816 = n17392 & ~n30815;
  assign n30817 = pi699 & ~n30816;
  assign n30818 = ~n30814 & n30817;
  assign n30819 = ~pi190 & ~pi699;
  assign n30820 = ~n17399 & n30819;
  assign n30821 = n3267 & ~n30820;
  assign n30822 = ~n30818 & n30821;
  assign n30823 = ~n30810 & ~n30822;
  assign n30824 = ~pi778 & ~n30823;
  assign n30825 = pi625 & n30823;
  assign n30826 = ~pi625 & n30808;
  assign n30827 = pi1153 & ~n30826;
  assign n30828 = ~n30825 & n30827;
  assign n30829 = ~pi625 & n30823;
  assign n30830 = pi625 & n30808;
  assign n30831 = ~pi1153 & ~n30830;
  assign n30832 = ~n30829 & n30831;
  assign n30833 = ~n30828 & ~n30832;
  assign n30834 = pi778 & ~n30833;
  assign n30835 = ~n30824 & ~n30834;
  assign n30836 = ~n17466 & ~n30835;
  assign n30837 = n17466 & ~n30808;
  assign n30838 = ~n30836 & ~n30837;
  assign n30839 = ~n17503 & n30838;
  assign n30840 = n17503 & n30808;
  assign n30841 = ~n30839 & ~n30840;
  assign n30842 = ~n17539 & n30841;
  assign n30843 = ~n30809 & ~n30842;
  assign n30844 = ~n17582 & n30843;
  assign n30845 = n17582 & n30808;
  assign n30846 = ~n30844 & ~n30845;
  assign n30847 = ~pi628 & ~n30846;
  assign n30848 = pi628 & n30808;
  assign n30849 = ~n30847 & ~n30848;
  assign n30850 = ~pi1156 & ~n30849;
  assign n30851 = pi628 & ~n30846;
  assign n30852 = ~pi628 & n30808;
  assign n30853 = ~n30851 & ~n30852;
  assign n30854 = pi1156 & ~n30853;
  assign n30855 = ~n30850 & ~n30854;
  assign n30856 = pi792 & ~n30855;
  assign n30857 = ~pi792 & ~n30846;
  assign n30858 = ~n30856 & ~n30857;
  assign n30859 = ~pi647 & ~n30858;
  assign n30860 = pi647 & n30808;
  assign n30861 = ~n30859 & ~n30860;
  assign n30862 = ~pi1157 & ~n30861;
  assign n30863 = pi647 & ~n30858;
  assign n30864 = ~pi647 & n30808;
  assign n30865 = ~n30863 & ~n30864;
  assign n30866 = pi1157 & ~n30865;
  assign n30867 = ~n30862 & ~n30866;
  assign n30868 = pi787 & ~n30867;
  assign n30869 = ~pi787 & ~n30858;
  assign n30870 = ~n30868 & ~n30869;
  assign n30871 = ~pi644 & ~n30870;
  assign n30872 = pi715 & ~n30871;
  assign n30873 = ~pi763 & n17199;
  assign n30874 = pi190 & n17273;
  assign n30875 = ~n30873 & ~n30874;
  assign n30876 = pi39 & ~n30875;
  assign n30877 = ~pi190 & pi763;
  assign n30878 = n17242 & n30877;
  assign n30879 = pi763 & ~n17246;
  assign n30880 = pi190 & ~n30879;
  assign n30881 = ~n22189 & ~n30880;
  assign n30882 = ~n30878 & n30881;
  assign n30883 = ~n30876 & n30882;
  assign n30884 = ~pi38 & ~n30883;
  assign n30885 = pi763 & n17282;
  assign n30886 = pi38 & ~n30815;
  assign n30887 = ~n30885 & n30886;
  assign n30888 = ~n30884 & ~n30887;
  assign n30889 = n3267 & ~n30888;
  assign n30890 = ~n30810 & ~n30889;
  assign n30891 = ~n17438 & ~n30890;
  assign n30892 = n17438 & ~n30808;
  assign n30893 = ~n30891 & ~n30892;
  assign n30894 = ~pi785 & ~n30893;
  assign n30895 = ~n17439 & ~n30808;
  assign n30896 = pi609 & n30891;
  assign n30897 = ~n30895 & ~n30896;
  assign n30898 = pi1155 & ~n30897;
  assign n30899 = ~n17451 & ~n30808;
  assign n30900 = ~pi609 & n30891;
  assign n30901 = ~n30899 & ~n30900;
  assign n30902 = ~pi1155 & ~n30901;
  assign n30903 = ~n30898 & ~n30902;
  assign n30904 = pi785 & ~n30903;
  assign n30905 = ~n30894 & ~n30904;
  assign n30906 = ~pi781 & ~n30905;
  assign n30907 = pi618 & n30905;
  assign n30908 = ~pi618 & n30808;
  assign n30909 = pi1154 & ~n30908;
  assign n30910 = ~n30907 & n30909;
  assign n30911 = ~pi618 & n30905;
  assign n30912 = pi618 & n30808;
  assign n30913 = ~pi1154 & ~n30912;
  assign n30914 = ~n30911 & n30913;
  assign n30915 = ~n30910 & ~n30914;
  assign n30916 = pi781 & ~n30915;
  assign n30917 = ~n30906 & ~n30916;
  assign n30918 = ~pi789 & ~n30917;
  assign n30919 = pi619 & n30917;
  assign n30920 = ~pi619 & n30808;
  assign n30921 = pi1159 & ~n30920;
  assign n30922 = ~n30919 & n30921;
  assign n30923 = ~pi619 & n30917;
  assign n30924 = pi619 & n30808;
  assign n30925 = ~pi1159 & ~n30924;
  assign n30926 = ~n30923 & n30925;
  assign n30927 = ~n30922 & ~n30926;
  assign n30928 = pi789 & ~n30927;
  assign n30929 = ~n30918 & ~n30928;
  assign n30930 = ~n17816 & n30929;
  assign n30931 = n17816 & n30808;
  assign n30932 = ~n30930 & ~n30931;
  assign n30933 = ~n17610 & ~n30932;
  assign n30934 = n17610 & n30808;
  assign n30935 = ~n30933 & ~n30934;
  assign n30936 = ~n17652 & ~n30935;
  assign n30937 = n17652 & n30808;
  assign n30938 = ~n30936 & ~n30937;
  assign n30939 = pi644 & ~n30938;
  assign n30940 = ~pi644 & n30808;
  assign n30941 = ~pi715 & ~n30940;
  assign n30942 = ~n30939 & n30941;
  assign n30943 = pi1160 & ~n30942;
  assign n30944 = ~n30872 & n30943;
  assign n30945 = pi644 & ~n30870;
  assign n30946 = ~pi715 & ~n30945;
  assign n30947 = ~pi644 & ~n30938;
  assign n30948 = pi644 & n30808;
  assign n30949 = pi715 & ~n30948;
  assign n30950 = ~n30947 & n30949;
  assign n30951 = ~pi1160 & ~n30950;
  assign n30952 = ~n30946 & n30951;
  assign n30953 = ~n30944 & ~n30952;
  assign n30954 = pi790 & ~n30953;
  assign n30955 = pi644 & n30943;
  assign n30956 = ~pi644 & n30951;
  assign n30957 = pi790 & ~n30956;
  assign n30958 = ~n30955 & n30957;
  assign n30959 = ~n20409 & n30932;
  assign n30960 = n17608 & n30849;
  assign n30961 = n17607 & n30853;
  assign n30962 = ~n30960 & ~n30961;
  assign n30963 = ~n30959 & n30962;
  assign n30964 = pi792 & ~n30963;
  assign n30965 = ~pi699 & n30888;
  assign n30966 = ~pi190 & n16687;
  assign n30967 = pi190 & n16799;
  assign n30968 = ~pi763 & ~n30967;
  assign n30969 = ~n30966 & n30968;
  assign n30970 = pi190 & n16879;
  assign n30971 = ~pi190 & ~n16944;
  assign n30972 = pi763 & ~n30971;
  assign n30973 = ~n30970 & n30972;
  assign n30974 = pi39 & ~n30973;
  assign n30975 = ~n30969 & n30974;
  assign n30976 = pi190 & n17059;
  assign n30977 = ~pi190 & n17088;
  assign n30978 = ~pi763 & ~n30977;
  assign n30979 = ~n30976 & n30978;
  assign n30980 = ~pi190 & ~n17092;
  assign n30981 = pi190 & ~n17094;
  assign n30982 = pi763 & ~n30981;
  assign n30983 = ~n30980 & n30982;
  assign n30984 = ~pi39 & ~n30983;
  assign n30985 = ~n30979 & n30984;
  assign n30986 = ~pi38 & ~n30985;
  assign n30987 = ~n30975 & n30986;
  assign n30988 = ~pi763 & n23906;
  assign n30989 = ~n16905 & ~n30988;
  assign n30990 = ~pi39 & ~n30989;
  assign n30991 = ~pi190 & ~n30990;
  assign n30992 = ~n16787 & ~n30623;
  assign n30993 = pi190 & ~n30992;
  assign n30994 = n6234 & n30993;
  assign n30995 = pi38 & ~n30994;
  assign n30996 = ~n30991 & n30995;
  assign n30997 = pi699 & ~n30996;
  assign n30998 = ~n30987 & n30997;
  assign n30999 = n3267 & ~n30998;
  assign n31000 = ~n30965 & n30999;
  assign n31001 = ~n30810 & ~n31000;
  assign n31002 = ~pi625 & n31001;
  assign n31003 = pi625 & n30890;
  assign n31004 = ~pi1153 & ~n31003;
  assign n31005 = ~n31002 & n31004;
  assign n31006 = ~pi608 & ~n30828;
  assign n31007 = ~n31005 & n31006;
  assign n31008 = pi625 & n31001;
  assign n31009 = ~pi625 & n30890;
  assign n31010 = pi1153 & ~n31009;
  assign n31011 = ~n31008 & n31010;
  assign n31012 = pi608 & ~n30832;
  assign n31013 = ~n31011 & n31012;
  assign n31014 = ~n31007 & ~n31013;
  assign n31015 = pi778 & ~n31014;
  assign n31016 = ~pi778 & n31001;
  assign n31017 = ~n31015 & ~n31016;
  assign n31018 = ~pi609 & ~n31017;
  assign n31019 = pi609 & n30835;
  assign n31020 = ~pi1155 & ~n31019;
  assign n31021 = ~n31018 & n31020;
  assign n31022 = ~pi660 & ~n30898;
  assign n31023 = ~n31021 & n31022;
  assign n31024 = pi609 & ~n31017;
  assign n31025 = ~pi609 & n30835;
  assign n31026 = pi1155 & ~n31025;
  assign n31027 = ~n31024 & n31026;
  assign n31028 = pi660 & ~n30902;
  assign n31029 = ~n31027 & n31028;
  assign n31030 = ~n31023 & ~n31029;
  assign n31031 = pi785 & ~n31030;
  assign n31032 = ~pi785 & ~n31017;
  assign n31033 = ~n31031 & ~n31032;
  assign n31034 = ~pi618 & ~n31033;
  assign n31035 = pi618 & n30838;
  assign n31036 = ~pi1154 & ~n31035;
  assign n31037 = ~n31034 & n31036;
  assign n31038 = ~pi627 & ~n30910;
  assign n31039 = ~n31037 & n31038;
  assign n31040 = pi618 & ~n31033;
  assign n31041 = ~pi618 & n30838;
  assign n31042 = pi1154 & ~n31041;
  assign n31043 = ~n31040 & n31042;
  assign n31044 = pi627 & ~n30914;
  assign n31045 = ~n31043 & n31044;
  assign n31046 = ~n31039 & ~n31045;
  assign n31047 = pi781 & ~n31046;
  assign n31048 = ~pi781 & ~n31033;
  assign n31049 = ~n31047 & ~n31048;
  assign n31050 = pi619 & ~n31049;
  assign n31051 = ~pi619 & ~n30841;
  assign n31052 = pi1159 & ~n31051;
  assign n31053 = ~n31050 & n31052;
  assign n31054 = pi648 & ~n30926;
  assign n31055 = ~n31053 & n31054;
  assign n31056 = ~pi619 & ~n31049;
  assign n31057 = pi619 & ~n30841;
  assign n31058 = ~pi1159 & ~n31057;
  assign n31059 = ~n31056 & n31058;
  assign n31060 = ~pi648 & ~n30922;
  assign n31061 = ~n31059 & n31060;
  assign n31062 = pi789 & ~n31061;
  assign n31063 = ~n31055 & n31062;
  assign n31064 = ~pi789 & n31049;
  assign n31065 = n17817 & ~n31064;
  assign n31066 = ~n31063 & n31065;
  assign n31067 = pi626 & ~n30929;
  assign n31068 = ~pi626 & ~n30808;
  assign n31069 = n17579 & ~n31068;
  assign n31070 = ~n31067 & n31069;
  assign n31071 = n17704 & n30843;
  assign n31072 = ~pi626 & ~n30929;
  assign n31073 = pi626 & ~n30808;
  assign n31074 = n17580 & ~n31073;
  assign n31075 = ~n31072 & n31074;
  assign n31076 = ~n31071 & ~n31075;
  assign n31077 = ~n31070 & n31076;
  assign n31078 = pi788 & ~n31077;
  assign n31079 = ~n20205 & ~n31078;
  assign n31080 = ~n31066 & n31079;
  assign n31081 = ~n30964 & ~n31080;
  assign n31082 = n20207 & ~n31081;
  assign n31083 = n17649 & n30865;
  assign n31084 = n17650 & n30861;
  assign n31085 = ~n20398 & n30935;
  assign n31086 = ~n31084 & ~n31085;
  assign n31087 = ~n31083 & n31086;
  assign n31088 = pi787 & ~n31087;
  assign n31089 = ~n31082 & ~n31088;
  assign n31090 = ~n30958 & n31089;
  assign n31091 = ~n30954 & ~n31090;
  assign n31092 = ~po1038 & ~n31091;
  assign n31093 = ~pi190 & po1038;
  assign n31094 = ~pi832 & ~n31093;
  assign n31095 = ~n31092 & n31094;
  assign po347 = ~n30807 & ~n31095;
  assign n31097 = ~pi191 & ~n2754;
  assign n31098 = pi746 & n16784;
  assign n31099 = ~n31097 & ~n31098;
  assign n31100 = ~n17706 & ~n31099;
  assign n31101 = ~pi785 & ~n31100;
  assign n31102 = n17451 & n31098;
  assign n31103 = n31100 & ~n31102;
  assign n31104 = pi1155 & ~n31103;
  assign n31105 = ~pi1155 & ~n31097;
  assign n31106 = ~n31102 & n31105;
  assign n31107 = ~n31104 & ~n31106;
  assign n31108 = pi785 & ~n31107;
  assign n31109 = ~n31101 & ~n31108;
  assign n31110 = ~pi781 & ~n31109;
  assign n31111 = ~n17721 & n31109;
  assign n31112 = pi1154 & ~n31111;
  assign n31113 = ~n17724 & n31109;
  assign n31114 = ~pi1154 & ~n31113;
  assign n31115 = ~n31112 & ~n31114;
  assign n31116 = pi781 & ~n31115;
  assign n31117 = ~n31110 & ~n31116;
  assign n31118 = ~pi789 & ~n31117;
  assign n31119 = ~n22890 & n31117;
  assign n31120 = pi1159 & ~n31119;
  assign n31121 = ~n22893 & n31117;
  assign n31122 = ~pi1159 & ~n31121;
  assign n31123 = ~n31120 & ~n31122;
  assign n31124 = pi789 & ~n31123;
  assign n31125 = ~n31118 & ~n31124;
  assign n31126 = ~n17816 & n31125;
  assign n31127 = n17816 & n31097;
  assign n31128 = ~n31126 & ~n31127;
  assign n31129 = ~n17610 & ~n31128;
  assign n31130 = n17610 & n31097;
  assign n31131 = ~n31129 & ~n31130;
  assign n31132 = ~n20398 & n31131;
  assign n31133 = pi729 & n16786;
  assign n31134 = ~n31097 & ~n31133;
  assign n31135 = ~pi778 & ~n31134;
  assign n31136 = ~pi625 & n31133;
  assign n31137 = ~n31134 & ~n31136;
  assign n31138 = pi1153 & ~n31137;
  assign n31139 = ~pi1153 & ~n31097;
  assign n31140 = ~n31136 & n31139;
  assign n31141 = pi778 & ~n31140;
  assign n31142 = ~n31138 & n31141;
  assign n31143 = ~n31135 & ~n31142;
  assign n31144 = ~n17692 & ~n31143;
  assign n31145 = ~n17694 & n31144;
  assign n31146 = ~n17696 & n31145;
  assign n31147 = ~n17828 & n31146;
  assign n31148 = ~n17859 & n31147;
  assign n31149 = ~pi647 & n31148;
  assign n31150 = pi647 & n31097;
  assign n31151 = ~pi1157 & ~n31150;
  assign n31152 = ~n31149 & n31151;
  assign n31153 = pi647 & ~n31148;
  assign n31154 = ~pi647 & ~n31097;
  assign n31155 = ~n31153 & ~n31154;
  assign n31156 = pi1157 & ~n31155;
  assign n31157 = ~n31152 & ~n31156;
  assign n31158 = ~n17651 & ~n31157;
  assign n31159 = ~n31132 & ~n31158;
  assign n31160 = pi787 & ~n31159;
  assign n31161 = pi626 & ~n31125;
  assign n31162 = ~pi626 & ~n31097;
  assign n31163 = n17579 & ~n31162;
  assign n31164 = ~n31161 & n31163;
  assign n31165 = n17704 & n31146;
  assign n31166 = ~pi626 & ~n31125;
  assign n31167 = pi626 & ~n31097;
  assign n31168 = n17580 & ~n31167;
  assign n31169 = ~n31166 & n31168;
  assign n31170 = ~n31165 & ~n31169;
  assign n31171 = ~n31164 & n31170;
  assign n31172 = pi788 & ~n31171;
  assign n31173 = ~n16521 & ~n31134;
  assign n31174 = pi625 & n31173;
  assign n31175 = n31099 & ~n31173;
  assign n31176 = ~n31174 & ~n31175;
  assign n31177 = n31139 & ~n31176;
  assign n31178 = ~pi608 & ~n31138;
  assign n31179 = ~n31177 & n31178;
  assign n31180 = pi1153 & n31099;
  assign n31181 = ~n31174 & n31180;
  assign n31182 = pi608 & ~n31140;
  assign n31183 = ~n31181 & n31182;
  assign n31184 = ~n31179 & ~n31183;
  assign n31185 = pi778 & ~n31184;
  assign n31186 = ~pi778 & ~n31175;
  assign n31187 = ~n31185 & ~n31186;
  assign n31188 = ~pi609 & ~n31187;
  assign n31189 = pi609 & ~n31143;
  assign n31190 = ~pi1155 & ~n31189;
  assign n31191 = ~n31188 & n31190;
  assign n31192 = ~pi660 & ~n31104;
  assign n31193 = ~n31191 & n31192;
  assign n31194 = pi609 & ~n31187;
  assign n31195 = ~pi609 & ~n31143;
  assign n31196 = pi1155 & ~n31195;
  assign n31197 = ~n31194 & n31196;
  assign n31198 = pi660 & ~n31106;
  assign n31199 = ~n31197 & n31198;
  assign n31200 = ~n31193 & ~n31199;
  assign n31201 = pi785 & ~n31200;
  assign n31202 = ~pi785 & ~n31187;
  assign n31203 = ~n31201 & ~n31202;
  assign n31204 = ~pi618 & ~n31203;
  assign n31205 = pi618 & n31144;
  assign n31206 = ~pi1154 & ~n31205;
  assign n31207 = ~n31204 & n31206;
  assign n31208 = ~pi627 & ~n31112;
  assign n31209 = ~n31207 & n31208;
  assign n31210 = pi618 & ~n31203;
  assign n31211 = ~pi618 & n31144;
  assign n31212 = pi1154 & ~n31211;
  assign n31213 = ~n31210 & n31212;
  assign n31214 = pi627 & ~n31114;
  assign n31215 = ~n31213 & n31214;
  assign n31216 = ~n31209 & ~n31215;
  assign n31217 = pi781 & ~n31216;
  assign n31218 = ~pi781 & ~n31203;
  assign n31219 = ~n31217 & ~n31218;
  assign n31220 = pi619 & ~n31219;
  assign n31221 = ~pi619 & n31145;
  assign n31222 = pi1159 & ~n31221;
  assign n31223 = ~n31220 & n31222;
  assign n31224 = pi648 & ~n31122;
  assign n31225 = ~n31223 & n31224;
  assign n31226 = ~pi619 & ~n31219;
  assign n31227 = pi619 & n31145;
  assign n31228 = ~pi1159 & ~n31227;
  assign n31229 = ~n31226 & n31228;
  assign n31230 = ~pi648 & ~n31120;
  assign n31231 = ~n31229 & n31230;
  assign n31232 = pi789 & ~n31231;
  assign n31233 = ~n31225 & n31232;
  assign n31234 = ~pi789 & n31219;
  assign n31235 = n17817 & ~n31234;
  assign n31236 = ~n31233 & n31235;
  assign n31237 = ~n31172 & ~n31236;
  assign n31238 = ~n20205 & ~n31237;
  assign n31239 = n17856 & ~n31128;
  assign n31240 = n20693 & n31147;
  assign n31241 = ~n31239 & ~n31240;
  assign n31242 = ~pi629 & ~n31241;
  assign n31243 = n20697 & n31147;
  assign n31244 = n17855 & ~n31128;
  assign n31245 = ~n31243 & ~n31244;
  assign n31246 = pi629 & ~n31245;
  assign n31247 = ~n31242 & ~n31246;
  assign n31248 = pi792 & ~n31247;
  assign n31249 = n20207 & ~n31248;
  assign n31250 = ~n31238 & n31249;
  assign n31251 = ~n31160 & ~n31250;
  assign n31252 = pi644 & n31251;
  assign n31253 = ~pi787 & ~n31148;
  assign n31254 = pi787 & ~n31157;
  assign n31255 = ~n31253 & ~n31254;
  assign n31256 = ~pi644 & n31255;
  assign n31257 = pi715 & ~n31256;
  assign n31258 = ~n31252 & n31257;
  assign n31259 = ~n17652 & ~n31131;
  assign n31260 = n17652 & n31097;
  assign n31261 = ~n31259 & ~n31260;
  assign n31262 = pi644 & ~n31261;
  assign n31263 = ~pi644 & n31097;
  assign n31264 = ~pi715 & ~n31263;
  assign n31265 = ~n31262 & n31264;
  assign n31266 = pi1160 & ~n31265;
  assign n31267 = ~n31258 & n31266;
  assign n31268 = ~pi644 & n31251;
  assign n31269 = pi644 & n31255;
  assign n31270 = ~pi715 & ~n31269;
  assign n31271 = ~n31268 & n31270;
  assign n31272 = ~pi644 & ~n31261;
  assign n31273 = pi644 & n31097;
  assign n31274 = pi715 & ~n31273;
  assign n31275 = ~n31272 & n31274;
  assign n31276 = ~pi1160 & ~n31275;
  assign n31277 = ~n31271 & n31276;
  assign n31278 = ~n31267 & ~n31277;
  assign n31279 = pi790 & ~n31278;
  assign n31280 = ~pi790 & n31251;
  assign n31281 = pi832 & ~n31280;
  assign n31282 = ~n31279 & n31281;
  assign n31283 = ~pi191 & ~n17406;
  assign n31284 = n17539 & ~n31283;
  assign n31285 = pi191 & ~n3267;
  assign n31286 = ~pi191 & n17972;
  assign n31287 = pi191 & ~n17976;
  assign n31288 = ~pi38 & ~n31287;
  assign n31289 = ~n31286 & n31288;
  assign n31290 = ~pi191 & ~n17280;
  assign n31291 = n17392 & ~n31290;
  assign n31292 = pi729 & ~n31291;
  assign n31293 = ~n31289 & n31292;
  assign n31294 = ~pi191 & ~pi729;
  assign n31295 = ~n17399 & n31294;
  assign n31296 = n3267 & ~n31295;
  assign n31297 = ~n31293 & n31296;
  assign n31298 = ~n31285 & ~n31297;
  assign n31299 = ~pi778 & ~n31298;
  assign n31300 = pi625 & n31298;
  assign n31301 = ~pi625 & n31283;
  assign n31302 = pi1153 & ~n31301;
  assign n31303 = ~n31300 & n31302;
  assign n31304 = ~pi625 & n31298;
  assign n31305 = pi625 & n31283;
  assign n31306 = ~pi1153 & ~n31305;
  assign n31307 = ~n31304 & n31306;
  assign n31308 = ~n31303 & ~n31307;
  assign n31309 = pi778 & ~n31308;
  assign n31310 = ~n31299 & ~n31309;
  assign n31311 = ~n17466 & ~n31310;
  assign n31312 = n17466 & ~n31283;
  assign n31313 = ~n31311 & ~n31312;
  assign n31314 = ~n17503 & n31313;
  assign n31315 = n17503 & n31283;
  assign n31316 = ~n31314 & ~n31315;
  assign n31317 = ~n17539 & n31316;
  assign n31318 = ~n31284 & ~n31317;
  assign n31319 = ~n17582 & n31318;
  assign n31320 = n17582 & n31283;
  assign n31321 = ~n31319 & ~n31320;
  assign n31322 = ~pi628 & ~n31321;
  assign n31323 = pi628 & n31283;
  assign n31324 = ~n31322 & ~n31323;
  assign n31325 = ~pi1156 & ~n31324;
  assign n31326 = pi628 & ~n31321;
  assign n31327 = ~pi628 & n31283;
  assign n31328 = ~n31326 & ~n31327;
  assign n31329 = pi1156 & ~n31328;
  assign n31330 = ~n31325 & ~n31329;
  assign n31331 = pi792 & ~n31330;
  assign n31332 = ~pi792 & ~n31321;
  assign n31333 = ~n31331 & ~n31332;
  assign n31334 = ~pi647 & ~n31333;
  assign n31335 = pi647 & n31283;
  assign n31336 = ~n31334 & ~n31335;
  assign n31337 = ~pi1157 & ~n31336;
  assign n31338 = pi647 & ~n31333;
  assign n31339 = ~pi647 & n31283;
  assign n31340 = ~n31338 & ~n31339;
  assign n31341 = pi1157 & ~n31340;
  assign n31342 = ~n31337 & ~n31341;
  assign n31343 = pi787 & ~n31342;
  assign n31344 = ~pi787 & ~n31333;
  assign n31345 = ~n31343 & ~n31344;
  assign n31346 = ~pi644 & ~n31345;
  assign n31347 = pi715 & ~n31346;
  assign n31348 = ~pi746 & n17199;
  assign n31349 = pi191 & n17273;
  assign n31350 = ~n31348 & ~n31349;
  assign n31351 = pi39 & ~n31350;
  assign n31352 = ~pi191 & pi746;
  assign n31353 = n17242 & n31352;
  assign n31354 = pi746 & ~n17246;
  assign n31355 = pi191 & ~n31354;
  assign n31356 = ~n22270 & ~n31355;
  assign n31357 = ~n31353 & n31356;
  assign n31358 = ~n31351 & n31357;
  assign n31359 = ~pi38 & ~n31358;
  assign n31360 = pi746 & n17282;
  assign n31361 = pi38 & ~n31290;
  assign n31362 = ~n31360 & n31361;
  assign n31363 = ~n31359 & ~n31362;
  assign n31364 = n3267 & ~n31363;
  assign n31365 = ~n31285 & ~n31364;
  assign n31366 = ~n17438 & ~n31365;
  assign n31367 = n17438 & ~n31283;
  assign n31368 = ~n31366 & ~n31367;
  assign n31369 = ~pi785 & ~n31368;
  assign n31370 = ~n17439 & ~n31283;
  assign n31371 = pi609 & n31366;
  assign n31372 = ~n31370 & ~n31371;
  assign n31373 = pi1155 & ~n31372;
  assign n31374 = ~n17451 & ~n31283;
  assign n31375 = ~pi609 & n31366;
  assign n31376 = ~n31374 & ~n31375;
  assign n31377 = ~pi1155 & ~n31376;
  assign n31378 = ~n31373 & ~n31377;
  assign n31379 = pi785 & ~n31378;
  assign n31380 = ~n31369 & ~n31379;
  assign n31381 = ~pi781 & ~n31380;
  assign n31382 = pi618 & n31380;
  assign n31383 = ~pi618 & n31283;
  assign n31384 = pi1154 & ~n31383;
  assign n31385 = ~n31382 & n31384;
  assign n31386 = ~pi618 & n31380;
  assign n31387 = pi618 & n31283;
  assign n31388 = ~pi1154 & ~n31387;
  assign n31389 = ~n31386 & n31388;
  assign n31390 = ~n31385 & ~n31389;
  assign n31391 = pi781 & ~n31390;
  assign n31392 = ~n31381 & ~n31391;
  assign n31393 = ~pi789 & ~n31392;
  assign n31394 = pi619 & n31392;
  assign n31395 = ~pi619 & n31283;
  assign n31396 = pi1159 & ~n31395;
  assign n31397 = ~n31394 & n31396;
  assign n31398 = ~pi619 & n31392;
  assign n31399 = pi619 & n31283;
  assign n31400 = ~pi1159 & ~n31399;
  assign n31401 = ~n31398 & n31400;
  assign n31402 = ~n31397 & ~n31401;
  assign n31403 = pi789 & ~n31402;
  assign n31404 = ~n31393 & ~n31403;
  assign n31405 = ~n17816 & n31404;
  assign n31406 = n17816 & n31283;
  assign n31407 = ~n31405 & ~n31406;
  assign n31408 = ~n17610 & ~n31407;
  assign n31409 = n17610 & n31283;
  assign n31410 = ~n31408 & ~n31409;
  assign n31411 = ~n17652 & ~n31410;
  assign n31412 = n17652 & n31283;
  assign n31413 = ~n31411 & ~n31412;
  assign n31414 = pi644 & ~n31413;
  assign n31415 = ~pi644 & n31283;
  assign n31416 = ~pi715 & ~n31415;
  assign n31417 = ~n31414 & n31416;
  assign n31418 = pi1160 & ~n31417;
  assign n31419 = ~n31347 & n31418;
  assign n31420 = pi644 & ~n31345;
  assign n31421 = ~pi715 & ~n31420;
  assign n31422 = ~pi644 & ~n31413;
  assign n31423 = pi644 & n31283;
  assign n31424 = pi715 & ~n31423;
  assign n31425 = ~n31422 & n31424;
  assign n31426 = ~pi1160 & ~n31425;
  assign n31427 = ~n31421 & n31426;
  assign n31428 = ~n31419 & ~n31427;
  assign n31429 = pi790 & ~n31428;
  assign n31430 = pi644 & n31418;
  assign n31431 = ~pi644 & n31426;
  assign n31432 = pi790 & ~n31431;
  assign n31433 = ~n31430 & n31432;
  assign n31434 = ~n20409 & n31407;
  assign n31435 = n17608 & n31324;
  assign n31436 = n17607 & n31328;
  assign n31437 = ~n31435 & ~n31436;
  assign n31438 = ~n31434 & n31437;
  assign n31439 = pi792 & ~n31438;
  assign n31440 = ~pi729 & n31363;
  assign n31441 = ~pi191 & n16687;
  assign n31442 = pi191 & n16799;
  assign n31443 = ~pi746 & ~n31442;
  assign n31444 = ~n31441 & n31443;
  assign n31445 = pi191 & n16879;
  assign n31446 = ~pi191 & ~n16944;
  assign n31447 = pi746 & ~n31446;
  assign n31448 = ~n31445 & n31447;
  assign n31449 = pi39 & ~n31448;
  assign n31450 = ~n31444 & n31449;
  assign n31451 = pi191 & n17059;
  assign n31452 = ~pi191 & n17088;
  assign n31453 = ~pi746 & ~n31452;
  assign n31454 = ~n31451 & n31453;
  assign n31455 = ~pi191 & ~n17092;
  assign n31456 = pi191 & ~n17094;
  assign n31457 = pi746 & ~n31456;
  assign n31458 = ~n31455 & n31457;
  assign n31459 = ~pi39 & ~n31458;
  assign n31460 = ~n31454 & n31459;
  assign n31461 = ~pi38 & ~n31460;
  assign n31462 = ~n31450 & n31461;
  assign n31463 = ~pi746 & n23906;
  assign n31464 = ~n16905 & ~n31463;
  assign n31465 = ~pi39 & ~n31464;
  assign n31466 = ~pi191 & ~n31465;
  assign n31467 = ~n16787 & ~n31098;
  assign n31468 = pi191 & ~n31467;
  assign n31469 = n6234 & n31468;
  assign n31470 = pi38 & ~n31469;
  assign n31471 = ~n31466 & n31470;
  assign n31472 = pi729 & ~n31471;
  assign n31473 = ~n31462 & n31472;
  assign n31474 = n3267 & ~n31473;
  assign n31475 = ~n31440 & n31474;
  assign n31476 = ~n31285 & ~n31475;
  assign n31477 = ~pi625 & n31476;
  assign n31478 = pi625 & n31365;
  assign n31479 = ~pi1153 & ~n31478;
  assign n31480 = ~n31477 & n31479;
  assign n31481 = ~pi608 & ~n31303;
  assign n31482 = ~n31480 & n31481;
  assign n31483 = pi625 & n31476;
  assign n31484 = ~pi625 & n31365;
  assign n31485 = pi1153 & ~n31484;
  assign n31486 = ~n31483 & n31485;
  assign n31487 = pi608 & ~n31307;
  assign n31488 = ~n31486 & n31487;
  assign n31489 = ~n31482 & ~n31488;
  assign n31490 = pi778 & ~n31489;
  assign n31491 = ~pi778 & n31476;
  assign n31492 = ~n31490 & ~n31491;
  assign n31493 = ~pi609 & ~n31492;
  assign n31494 = pi609 & n31310;
  assign n31495 = ~pi1155 & ~n31494;
  assign n31496 = ~n31493 & n31495;
  assign n31497 = ~pi660 & ~n31373;
  assign n31498 = ~n31496 & n31497;
  assign n31499 = pi609 & ~n31492;
  assign n31500 = ~pi609 & n31310;
  assign n31501 = pi1155 & ~n31500;
  assign n31502 = ~n31499 & n31501;
  assign n31503 = pi660 & ~n31377;
  assign n31504 = ~n31502 & n31503;
  assign n31505 = ~n31498 & ~n31504;
  assign n31506 = pi785 & ~n31505;
  assign n31507 = ~pi785 & ~n31492;
  assign n31508 = ~n31506 & ~n31507;
  assign n31509 = ~pi618 & ~n31508;
  assign n31510 = pi618 & n31313;
  assign n31511 = ~pi1154 & ~n31510;
  assign n31512 = ~n31509 & n31511;
  assign n31513 = ~pi627 & ~n31385;
  assign n31514 = ~n31512 & n31513;
  assign n31515 = pi618 & ~n31508;
  assign n31516 = ~pi618 & n31313;
  assign n31517 = pi1154 & ~n31516;
  assign n31518 = ~n31515 & n31517;
  assign n31519 = pi627 & ~n31389;
  assign n31520 = ~n31518 & n31519;
  assign n31521 = ~n31514 & ~n31520;
  assign n31522 = pi781 & ~n31521;
  assign n31523 = ~pi781 & ~n31508;
  assign n31524 = ~n31522 & ~n31523;
  assign n31525 = pi619 & ~n31524;
  assign n31526 = ~pi619 & ~n31316;
  assign n31527 = pi1159 & ~n31526;
  assign n31528 = ~n31525 & n31527;
  assign n31529 = pi648 & ~n31401;
  assign n31530 = ~n31528 & n31529;
  assign n31531 = ~pi619 & ~n31524;
  assign n31532 = pi619 & ~n31316;
  assign n31533 = ~pi1159 & ~n31532;
  assign n31534 = ~n31531 & n31533;
  assign n31535 = ~pi648 & ~n31397;
  assign n31536 = ~n31534 & n31535;
  assign n31537 = pi789 & ~n31536;
  assign n31538 = ~n31530 & n31537;
  assign n31539 = ~pi789 & n31524;
  assign n31540 = n17817 & ~n31539;
  assign n31541 = ~n31538 & n31540;
  assign n31542 = pi626 & ~n31404;
  assign n31543 = ~pi626 & ~n31283;
  assign n31544 = n17579 & ~n31543;
  assign n31545 = ~n31542 & n31544;
  assign n31546 = n17704 & n31318;
  assign n31547 = ~pi626 & ~n31404;
  assign n31548 = pi626 & ~n31283;
  assign n31549 = n17580 & ~n31548;
  assign n31550 = ~n31547 & n31549;
  assign n31551 = ~n31546 & ~n31550;
  assign n31552 = ~n31545 & n31551;
  assign n31553 = pi788 & ~n31552;
  assign n31554 = ~n20205 & ~n31553;
  assign n31555 = ~n31541 & n31554;
  assign n31556 = ~n31439 & ~n31555;
  assign n31557 = n20207 & ~n31556;
  assign n31558 = n17649 & n31340;
  assign n31559 = n17650 & n31336;
  assign n31560 = ~n20398 & n31410;
  assign n31561 = ~n31559 & ~n31560;
  assign n31562 = ~n31558 & n31561;
  assign n31563 = pi787 & ~n31562;
  assign n31564 = ~n31557 & ~n31563;
  assign n31565 = ~n31433 & n31564;
  assign n31566 = ~n31429 & ~n31565;
  assign n31567 = ~po1038 & ~n31566;
  assign n31568 = ~pi191 & po1038;
  assign n31569 = ~pi832 & ~n31568;
  assign n31570 = ~n31567 & n31569;
  assign po348 = ~n31282 & ~n31570;
  assign n31572 = ~pi192 & ~n2754;
  assign n31573 = pi764 & n16784;
  assign n31574 = ~n31572 & ~n31573;
  assign n31575 = ~n17706 & ~n31574;
  assign n31576 = ~pi785 & ~n31575;
  assign n31577 = n17451 & n31573;
  assign n31578 = n31575 & ~n31577;
  assign n31579 = pi1155 & ~n31578;
  assign n31580 = ~pi1155 & ~n31572;
  assign n31581 = ~n31577 & n31580;
  assign n31582 = ~n31579 & ~n31581;
  assign n31583 = pi785 & ~n31582;
  assign n31584 = ~n31576 & ~n31583;
  assign n31585 = ~pi781 & ~n31584;
  assign n31586 = ~n17721 & n31584;
  assign n31587 = pi1154 & ~n31586;
  assign n31588 = ~n17724 & n31584;
  assign n31589 = ~pi1154 & ~n31588;
  assign n31590 = ~n31587 & ~n31589;
  assign n31591 = pi781 & ~n31590;
  assign n31592 = ~n31585 & ~n31591;
  assign n31593 = ~pi789 & ~n31592;
  assign n31594 = ~n22890 & n31592;
  assign n31595 = pi1159 & ~n31594;
  assign n31596 = ~n22893 & n31592;
  assign n31597 = ~pi1159 & ~n31596;
  assign n31598 = ~n31595 & ~n31597;
  assign n31599 = pi789 & ~n31598;
  assign n31600 = ~n31593 & ~n31599;
  assign n31601 = ~n17816 & n31600;
  assign n31602 = n17816 & n31572;
  assign n31603 = ~n31601 & ~n31602;
  assign n31604 = ~n17610 & ~n31603;
  assign n31605 = n17610 & n31572;
  assign n31606 = ~n31604 & ~n31605;
  assign n31607 = ~n20398 & n31606;
  assign n31608 = pi691 & n16786;
  assign n31609 = ~n31572 & ~n31608;
  assign n31610 = ~pi778 & ~n31609;
  assign n31611 = ~pi625 & n31608;
  assign n31612 = ~n31609 & ~n31611;
  assign n31613 = pi1153 & ~n31612;
  assign n31614 = ~pi1153 & ~n31572;
  assign n31615 = ~n31611 & n31614;
  assign n31616 = pi778 & ~n31615;
  assign n31617 = ~n31613 & n31616;
  assign n31618 = ~n31610 & ~n31617;
  assign n31619 = ~n17692 & ~n31618;
  assign n31620 = ~n17694 & n31619;
  assign n31621 = ~n17696 & n31620;
  assign n31622 = ~n17828 & n31621;
  assign n31623 = ~n17859 & n31622;
  assign n31624 = ~pi647 & n31623;
  assign n31625 = pi647 & n31572;
  assign n31626 = ~pi1157 & ~n31625;
  assign n31627 = ~n31624 & n31626;
  assign n31628 = pi647 & ~n31623;
  assign n31629 = ~pi647 & ~n31572;
  assign n31630 = ~n31628 & ~n31629;
  assign n31631 = pi1157 & ~n31630;
  assign n31632 = ~n31627 & ~n31631;
  assign n31633 = ~n17651 & ~n31632;
  assign n31634 = ~n31607 & ~n31633;
  assign n31635 = pi787 & ~n31634;
  assign n31636 = pi626 & ~n31600;
  assign n31637 = ~pi626 & ~n31572;
  assign n31638 = n17579 & ~n31637;
  assign n31639 = ~n31636 & n31638;
  assign n31640 = n17704 & n31621;
  assign n31641 = ~pi626 & ~n31600;
  assign n31642 = pi626 & ~n31572;
  assign n31643 = n17580 & ~n31642;
  assign n31644 = ~n31641 & n31643;
  assign n31645 = ~n31640 & ~n31644;
  assign n31646 = ~n31639 & n31645;
  assign n31647 = pi788 & ~n31646;
  assign n31648 = ~n16521 & ~n31609;
  assign n31649 = pi625 & n31648;
  assign n31650 = n31574 & ~n31648;
  assign n31651 = ~n31649 & ~n31650;
  assign n31652 = n31614 & ~n31651;
  assign n31653 = ~pi608 & ~n31613;
  assign n31654 = ~n31652 & n31653;
  assign n31655 = pi1153 & n31574;
  assign n31656 = ~n31649 & n31655;
  assign n31657 = pi608 & ~n31615;
  assign n31658 = ~n31656 & n31657;
  assign n31659 = ~n31654 & ~n31658;
  assign n31660 = pi778 & ~n31659;
  assign n31661 = ~pi778 & ~n31650;
  assign n31662 = ~n31660 & ~n31661;
  assign n31663 = ~pi609 & ~n31662;
  assign n31664 = pi609 & ~n31618;
  assign n31665 = ~pi1155 & ~n31664;
  assign n31666 = ~n31663 & n31665;
  assign n31667 = ~pi660 & ~n31579;
  assign n31668 = ~n31666 & n31667;
  assign n31669 = pi609 & ~n31662;
  assign n31670 = ~pi609 & ~n31618;
  assign n31671 = pi1155 & ~n31670;
  assign n31672 = ~n31669 & n31671;
  assign n31673 = pi660 & ~n31581;
  assign n31674 = ~n31672 & n31673;
  assign n31675 = ~n31668 & ~n31674;
  assign n31676 = pi785 & ~n31675;
  assign n31677 = ~pi785 & ~n31662;
  assign n31678 = ~n31676 & ~n31677;
  assign n31679 = ~pi618 & ~n31678;
  assign n31680 = pi618 & n31619;
  assign n31681 = ~pi1154 & ~n31680;
  assign n31682 = ~n31679 & n31681;
  assign n31683 = ~pi627 & ~n31587;
  assign n31684 = ~n31682 & n31683;
  assign n31685 = pi618 & ~n31678;
  assign n31686 = ~pi618 & n31619;
  assign n31687 = pi1154 & ~n31686;
  assign n31688 = ~n31685 & n31687;
  assign n31689 = pi627 & ~n31589;
  assign n31690 = ~n31688 & n31689;
  assign n31691 = ~n31684 & ~n31690;
  assign n31692 = pi781 & ~n31691;
  assign n31693 = ~pi781 & ~n31678;
  assign n31694 = ~n31692 & ~n31693;
  assign n31695 = pi619 & ~n31694;
  assign n31696 = ~pi619 & n31620;
  assign n31697 = pi1159 & ~n31696;
  assign n31698 = ~n31695 & n31697;
  assign n31699 = pi648 & ~n31597;
  assign n31700 = ~n31698 & n31699;
  assign n31701 = ~pi619 & ~n31694;
  assign n31702 = pi619 & n31620;
  assign n31703 = ~pi1159 & ~n31702;
  assign n31704 = ~n31701 & n31703;
  assign n31705 = ~pi648 & ~n31595;
  assign n31706 = ~n31704 & n31705;
  assign n31707 = pi789 & ~n31706;
  assign n31708 = ~n31700 & n31707;
  assign n31709 = ~pi789 & n31694;
  assign n31710 = n17817 & ~n31709;
  assign n31711 = ~n31708 & n31710;
  assign n31712 = ~n31647 & ~n31711;
  assign n31713 = ~n20205 & ~n31712;
  assign n31714 = n17856 & ~n31603;
  assign n31715 = n20693 & n31622;
  assign n31716 = ~n31714 & ~n31715;
  assign n31717 = ~pi629 & ~n31716;
  assign n31718 = n20697 & n31622;
  assign n31719 = n17855 & ~n31603;
  assign n31720 = ~n31718 & ~n31719;
  assign n31721 = pi629 & ~n31720;
  assign n31722 = ~n31717 & ~n31721;
  assign n31723 = pi792 & ~n31722;
  assign n31724 = n20207 & ~n31723;
  assign n31725 = ~n31713 & n31724;
  assign n31726 = ~n31635 & ~n31725;
  assign n31727 = pi644 & n31726;
  assign n31728 = ~pi787 & ~n31623;
  assign n31729 = pi787 & ~n31632;
  assign n31730 = ~n31728 & ~n31729;
  assign n31731 = ~pi644 & n31730;
  assign n31732 = pi715 & ~n31731;
  assign n31733 = ~n31727 & n31732;
  assign n31734 = ~n17652 & ~n31606;
  assign n31735 = n17652 & n31572;
  assign n31736 = ~n31734 & ~n31735;
  assign n31737 = pi644 & ~n31736;
  assign n31738 = ~pi644 & n31572;
  assign n31739 = ~pi715 & ~n31738;
  assign n31740 = ~n31737 & n31739;
  assign n31741 = pi1160 & ~n31740;
  assign n31742 = ~n31733 & n31741;
  assign n31743 = ~pi644 & n31726;
  assign n31744 = pi644 & n31730;
  assign n31745 = ~pi715 & ~n31744;
  assign n31746 = ~n31743 & n31745;
  assign n31747 = ~pi644 & ~n31736;
  assign n31748 = pi644 & n31572;
  assign n31749 = pi715 & ~n31748;
  assign n31750 = ~n31747 & n31749;
  assign n31751 = ~pi1160 & ~n31750;
  assign n31752 = ~n31746 & n31751;
  assign n31753 = ~n31742 & ~n31752;
  assign n31754 = pi790 & ~n31753;
  assign n31755 = ~pi790 & n31726;
  assign n31756 = pi832 & ~n31755;
  assign n31757 = ~n31754 & n31756;
  assign n31758 = ~pi192 & ~n17406;
  assign n31759 = n17539 & ~n31758;
  assign n31760 = pi192 & ~n3267;
  assign n31761 = ~pi192 & n17972;
  assign n31762 = pi192 & ~n17976;
  assign n31763 = ~pi38 & ~n31762;
  assign n31764 = ~n31761 & n31763;
  assign n31765 = ~pi192 & ~n17280;
  assign n31766 = n17392 & ~n31765;
  assign n31767 = pi691 & ~n31766;
  assign n31768 = ~n31764 & n31767;
  assign n31769 = ~pi192 & ~pi691;
  assign n31770 = ~n17399 & n31769;
  assign n31771 = n3267 & ~n31770;
  assign n31772 = ~n31768 & n31771;
  assign n31773 = ~n31760 & ~n31772;
  assign n31774 = ~pi778 & ~n31773;
  assign n31775 = pi625 & n31773;
  assign n31776 = ~pi625 & n31758;
  assign n31777 = pi1153 & ~n31776;
  assign n31778 = ~n31775 & n31777;
  assign n31779 = ~pi625 & n31773;
  assign n31780 = pi625 & n31758;
  assign n31781 = ~pi1153 & ~n31780;
  assign n31782 = ~n31779 & n31781;
  assign n31783 = ~n31778 & ~n31782;
  assign n31784 = pi778 & ~n31783;
  assign n31785 = ~n31774 & ~n31784;
  assign n31786 = ~n17466 & ~n31785;
  assign n31787 = n17466 & ~n31758;
  assign n31788 = ~n31786 & ~n31787;
  assign n31789 = ~n17503 & n31788;
  assign n31790 = n17503 & n31758;
  assign n31791 = ~n31789 & ~n31790;
  assign n31792 = ~n17539 & n31791;
  assign n31793 = ~n31759 & ~n31792;
  assign n31794 = ~n17582 & n31793;
  assign n31795 = n17582 & n31758;
  assign n31796 = ~n31794 & ~n31795;
  assign n31797 = ~pi628 & ~n31796;
  assign n31798 = pi628 & n31758;
  assign n31799 = ~n31797 & ~n31798;
  assign n31800 = ~pi1156 & ~n31799;
  assign n31801 = pi628 & ~n31796;
  assign n31802 = ~pi628 & n31758;
  assign n31803 = ~n31801 & ~n31802;
  assign n31804 = pi1156 & ~n31803;
  assign n31805 = ~n31800 & ~n31804;
  assign n31806 = pi792 & ~n31805;
  assign n31807 = ~pi792 & ~n31796;
  assign n31808 = ~n31806 & ~n31807;
  assign n31809 = ~pi647 & ~n31808;
  assign n31810 = pi647 & n31758;
  assign n31811 = ~n31809 & ~n31810;
  assign n31812 = ~pi1157 & ~n31811;
  assign n31813 = pi647 & ~n31808;
  assign n31814 = ~pi647 & n31758;
  assign n31815 = ~n31813 & ~n31814;
  assign n31816 = pi1157 & ~n31815;
  assign n31817 = ~n31812 & ~n31816;
  assign n31818 = pi787 & ~n31817;
  assign n31819 = ~pi787 & ~n31808;
  assign n31820 = ~n31818 & ~n31819;
  assign n31821 = ~pi644 & ~n31820;
  assign n31822 = pi715 & ~n31821;
  assign n31823 = ~pi764 & n17199;
  assign n31824 = pi192 & n17273;
  assign n31825 = ~n31823 & ~n31824;
  assign n31826 = pi39 & ~n31825;
  assign n31827 = ~pi192 & pi764;
  assign n31828 = n17242 & n31827;
  assign n31829 = pi764 & ~n17246;
  assign n31830 = pi192 & ~n31829;
  assign n31831 = ~n22431 & ~n31830;
  assign n31832 = ~n31828 & n31831;
  assign n31833 = ~n31826 & n31832;
  assign n31834 = ~pi38 & ~n31833;
  assign n31835 = pi764 & n17282;
  assign n31836 = pi38 & ~n31765;
  assign n31837 = ~n31835 & n31836;
  assign n31838 = ~n31834 & ~n31837;
  assign n31839 = n3267 & ~n31838;
  assign n31840 = ~n31760 & ~n31839;
  assign n31841 = ~n17438 & ~n31840;
  assign n31842 = n17438 & ~n31758;
  assign n31843 = ~n31841 & ~n31842;
  assign n31844 = ~pi785 & ~n31843;
  assign n31845 = ~n17439 & ~n31758;
  assign n31846 = pi609 & n31841;
  assign n31847 = ~n31845 & ~n31846;
  assign n31848 = pi1155 & ~n31847;
  assign n31849 = ~n17451 & ~n31758;
  assign n31850 = ~pi609 & n31841;
  assign n31851 = ~n31849 & ~n31850;
  assign n31852 = ~pi1155 & ~n31851;
  assign n31853 = ~n31848 & ~n31852;
  assign n31854 = pi785 & ~n31853;
  assign n31855 = ~n31844 & ~n31854;
  assign n31856 = ~pi781 & ~n31855;
  assign n31857 = pi618 & n31855;
  assign n31858 = ~pi618 & n31758;
  assign n31859 = pi1154 & ~n31858;
  assign n31860 = ~n31857 & n31859;
  assign n31861 = ~pi618 & n31855;
  assign n31862 = pi618 & n31758;
  assign n31863 = ~pi1154 & ~n31862;
  assign n31864 = ~n31861 & n31863;
  assign n31865 = ~n31860 & ~n31864;
  assign n31866 = pi781 & ~n31865;
  assign n31867 = ~n31856 & ~n31866;
  assign n31868 = ~pi789 & ~n31867;
  assign n31869 = pi619 & n31867;
  assign n31870 = ~pi619 & n31758;
  assign n31871 = pi1159 & ~n31870;
  assign n31872 = ~n31869 & n31871;
  assign n31873 = ~pi619 & n31867;
  assign n31874 = pi619 & n31758;
  assign n31875 = ~pi1159 & ~n31874;
  assign n31876 = ~n31873 & n31875;
  assign n31877 = ~n31872 & ~n31876;
  assign n31878 = pi789 & ~n31877;
  assign n31879 = ~n31868 & ~n31878;
  assign n31880 = ~n17816 & n31879;
  assign n31881 = n17816 & n31758;
  assign n31882 = ~n31880 & ~n31881;
  assign n31883 = ~n17610 & ~n31882;
  assign n31884 = n17610 & n31758;
  assign n31885 = ~n31883 & ~n31884;
  assign n31886 = ~n17652 & ~n31885;
  assign n31887 = n17652 & n31758;
  assign n31888 = ~n31886 & ~n31887;
  assign n31889 = pi644 & ~n31888;
  assign n31890 = ~pi644 & n31758;
  assign n31891 = ~pi715 & ~n31890;
  assign n31892 = ~n31889 & n31891;
  assign n31893 = pi1160 & ~n31892;
  assign n31894 = ~n31822 & n31893;
  assign n31895 = pi644 & ~n31820;
  assign n31896 = ~pi715 & ~n31895;
  assign n31897 = ~pi644 & ~n31888;
  assign n31898 = pi644 & n31758;
  assign n31899 = pi715 & ~n31898;
  assign n31900 = ~n31897 & n31899;
  assign n31901 = ~pi1160 & ~n31900;
  assign n31902 = ~n31896 & n31901;
  assign n31903 = ~n31894 & ~n31902;
  assign n31904 = pi790 & ~n31903;
  assign n31905 = pi644 & n31893;
  assign n31906 = ~pi644 & n31901;
  assign n31907 = pi790 & ~n31906;
  assign n31908 = ~n31905 & n31907;
  assign n31909 = ~n20409 & n31882;
  assign n31910 = n17608 & n31799;
  assign n31911 = n17607 & n31803;
  assign n31912 = ~n31910 & ~n31911;
  assign n31913 = ~n31909 & n31912;
  assign n31914 = pi792 & ~n31913;
  assign n31915 = ~pi691 & n31838;
  assign n31916 = ~pi192 & n16687;
  assign n31917 = pi192 & n16799;
  assign n31918 = ~pi764 & ~n31917;
  assign n31919 = ~n31916 & n31918;
  assign n31920 = pi192 & n16879;
  assign n31921 = ~pi192 & ~n16944;
  assign n31922 = pi764 & ~n31921;
  assign n31923 = ~n31920 & n31922;
  assign n31924 = pi39 & ~n31923;
  assign n31925 = ~n31919 & n31924;
  assign n31926 = pi192 & n17059;
  assign n31927 = ~pi192 & n17088;
  assign n31928 = ~pi764 & ~n31927;
  assign n31929 = ~n31926 & n31928;
  assign n31930 = ~pi192 & ~n17092;
  assign n31931 = pi192 & ~n17094;
  assign n31932 = pi764 & ~n31931;
  assign n31933 = ~n31930 & n31932;
  assign n31934 = ~pi39 & ~n31933;
  assign n31935 = ~n31929 & n31934;
  assign n31936 = ~pi38 & ~n31935;
  assign n31937 = ~n31925 & n31936;
  assign n31938 = ~pi764 & n23906;
  assign n31939 = ~n16905 & ~n31938;
  assign n31940 = ~pi39 & ~n31939;
  assign n31941 = ~pi192 & ~n31940;
  assign n31942 = ~n16787 & ~n31573;
  assign n31943 = pi192 & ~n31942;
  assign n31944 = n6234 & n31943;
  assign n31945 = pi38 & ~n31944;
  assign n31946 = ~n31941 & n31945;
  assign n31947 = pi691 & ~n31946;
  assign n31948 = ~n31937 & n31947;
  assign n31949 = n3267 & ~n31948;
  assign n31950 = ~n31915 & n31949;
  assign n31951 = ~n31760 & ~n31950;
  assign n31952 = ~pi625 & n31951;
  assign n31953 = pi625 & n31840;
  assign n31954 = ~pi1153 & ~n31953;
  assign n31955 = ~n31952 & n31954;
  assign n31956 = ~pi608 & ~n31778;
  assign n31957 = ~n31955 & n31956;
  assign n31958 = pi625 & n31951;
  assign n31959 = ~pi625 & n31840;
  assign n31960 = pi1153 & ~n31959;
  assign n31961 = ~n31958 & n31960;
  assign n31962 = pi608 & ~n31782;
  assign n31963 = ~n31961 & n31962;
  assign n31964 = ~n31957 & ~n31963;
  assign n31965 = pi778 & ~n31964;
  assign n31966 = ~pi778 & n31951;
  assign n31967 = ~n31965 & ~n31966;
  assign n31968 = ~pi609 & ~n31967;
  assign n31969 = pi609 & n31785;
  assign n31970 = ~pi1155 & ~n31969;
  assign n31971 = ~n31968 & n31970;
  assign n31972 = ~pi660 & ~n31848;
  assign n31973 = ~n31971 & n31972;
  assign n31974 = pi609 & ~n31967;
  assign n31975 = ~pi609 & n31785;
  assign n31976 = pi1155 & ~n31975;
  assign n31977 = ~n31974 & n31976;
  assign n31978 = pi660 & ~n31852;
  assign n31979 = ~n31977 & n31978;
  assign n31980 = ~n31973 & ~n31979;
  assign n31981 = pi785 & ~n31980;
  assign n31982 = ~pi785 & ~n31967;
  assign n31983 = ~n31981 & ~n31982;
  assign n31984 = ~pi618 & ~n31983;
  assign n31985 = pi618 & n31788;
  assign n31986 = ~pi1154 & ~n31985;
  assign n31987 = ~n31984 & n31986;
  assign n31988 = ~pi627 & ~n31860;
  assign n31989 = ~n31987 & n31988;
  assign n31990 = pi618 & ~n31983;
  assign n31991 = ~pi618 & n31788;
  assign n31992 = pi1154 & ~n31991;
  assign n31993 = ~n31990 & n31992;
  assign n31994 = pi627 & ~n31864;
  assign n31995 = ~n31993 & n31994;
  assign n31996 = ~n31989 & ~n31995;
  assign n31997 = pi781 & ~n31996;
  assign n31998 = ~pi781 & ~n31983;
  assign n31999 = ~n31997 & ~n31998;
  assign n32000 = pi619 & ~n31999;
  assign n32001 = ~pi619 & ~n31791;
  assign n32002 = pi1159 & ~n32001;
  assign n32003 = ~n32000 & n32002;
  assign n32004 = pi648 & ~n31876;
  assign n32005 = ~n32003 & n32004;
  assign n32006 = ~pi619 & ~n31999;
  assign n32007 = pi619 & ~n31791;
  assign n32008 = ~pi1159 & ~n32007;
  assign n32009 = ~n32006 & n32008;
  assign n32010 = ~pi648 & ~n31872;
  assign n32011 = ~n32009 & n32010;
  assign n32012 = pi789 & ~n32011;
  assign n32013 = ~n32005 & n32012;
  assign n32014 = ~pi789 & n31999;
  assign n32015 = n17817 & ~n32014;
  assign n32016 = ~n32013 & n32015;
  assign n32017 = pi626 & ~n31879;
  assign n32018 = ~pi626 & ~n31758;
  assign n32019 = n17579 & ~n32018;
  assign n32020 = ~n32017 & n32019;
  assign n32021 = n17704 & n31793;
  assign n32022 = ~pi626 & ~n31879;
  assign n32023 = pi626 & ~n31758;
  assign n32024 = n17580 & ~n32023;
  assign n32025 = ~n32022 & n32024;
  assign n32026 = ~n32021 & ~n32025;
  assign n32027 = ~n32020 & n32026;
  assign n32028 = pi788 & ~n32027;
  assign n32029 = ~n20205 & ~n32028;
  assign n32030 = ~n32016 & n32029;
  assign n32031 = ~n31914 & ~n32030;
  assign n32032 = n20207 & ~n32031;
  assign n32033 = n17649 & n31815;
  assign n32034 = n17650 & n31811;
  assign n32035 = ~n20398 & n31885;
  assign n32036 = ~n32034 & ~n32035;
  assign n32037 = ~n32033 & n32036;
  assign n32038 = pi787 & ~n32037;
  assign n32039 = ~n32032 & ~n32038;
  assign n32040 = ~n31908 & n32039;
  assign n32041 = ~n31904 & ~n32040;
  assign n32042 = ~po1038 & ~n32041;
  assign n32043 = ~pi192 & po1038;
  assign n32044 = ~pi832 & ~n32043;
  assign n32045 = ~n32042 & n32044;
  assign po349 = ~n31757 & ~n32045;
  assign n32047 = ~pi193 & ~n2754;
  assign n32048 = pi739 & n16784;
  assign n32049 = ~n32047 & ~n32048;
  assign n32050 = ~n17706 & ~n32049;
  assign n32051 = ~pi785 & ~n32050;
  assign n32052 = n17451 & n32048;
  assign n32053 = n32050 & ~n32052;
  assign n32054 = pi1155 & ~n32053;
  assign n32055 = ~pi1155 & ~n32047;
  assign n32056 = ~n32052 & n32055;
  assign n32057 = ~n32054 & ~n32056;
  assign n32058 = pi785 & ~n32057;
  assign n32059 = ~n32051 & ~n32058;
  assign n32060 = ~pi781 & ~n32059;
  assign n32061 = ~n17721 & n32059;
  assign n32062 = pi1154 & ~n32061;
  assign n32063 = ~n17724 & n32059;
  assign n32064 = ~pi1154 & ~n32063;
  assign n32065 = ~n32062 & ~n32064;
  assign n32066 = pi781 & ~n32065;
  assign n32067 = ~n32060 & ~n32066;
  assign n32068 = ~pi789 & ~n32067;
  assign n32069 = ~n22890 & n32067;
  assign n32070 = pi1159 & ~n32069;
  assign n32071 = ~n22893 & n32067;
  assign n32072 = ~pi1159 & ~n32071;
  assign n32073 = ~n32070 & ~n32072;
  assign n32074 = pi789 & ~n32073;
  assign n32075 = ~n32068 & ~n32074;
  assign n32076 = ~n17816 & n32075;
  assign n32077 = n17816 & n32047;
  assign n32078 = ~n32076 & ~n32077;
  assign n32079 = ~n17610 & ~n32078;
  assign n32080 = n17610 & n32047;
  assign n32081 = ~n32079 & ~n32080;
  assign n32082 = ~n20398 & n32081;
  assign n32083 = pi690 & n16786;
  assign n32084 = ~n32047 & ~n32083;
  assign n32085 = ~pi778 & ~n32084;
  assign n32086 = ~pi625 & n32083;
  assign n32087 = ~n32084 & ~n32086;
  assign n32088 = pi1153 & ~n32087;
  assign n32089 = ~pi1153 & ~n32047;
  assign n32090 = ~n32086 & n32089;
  assign n32091 = pi778 & ~n32090;
  assign n32092 = ~n32088 & n32091;
  assign n32093 = ~n32085 & ~n32092;
  assign n32094 = ~n17692 & ~n32093;
  assign n32095 = ~n17694 & n32094;
  assign n32096 = ~n17696 & n32095;
  assign n32097 = ~n17828 & n32096;
  assign n32098 = ~n17859 & n32097;
  assign n32099 = ~pi647 & n32098;
  assign n32100 = pi647 & n32047;
  assign n32101 = ~pi1157 & ~n32100;
  assign n32102 = ~n32099 & n32101;
  assign n32103 = pi647 & ~n32098;
  assign n32104 = ~pi647 & ~n32047;
  assign n32105 = ~n32103 & ~n32104;
  assign n32106 = pi1157 & ~n32105;
  assign n32107 = ~n32102 & ~n32106;
  assign n32108 = ~n17651 & ~n32107;
  assign n32109 = ~n32082 & ~n32108;
  assign n32110 = pi787 & ~n32109;
  assign n32111 = pi626 & ~n32075;
  assign n32112 = ~pi626 & ~n32047;
  assign n32113 = n17579 & ~n32112;
  assign n32114 = ~n32111 & n32113;
  assign n32115 = n17704 & n32096;
  assign n32116 = ~pi626 & ~n32075;
  assign n32117 = pi626 & ~n32047;
  assign n32118 = n17580 & ~n32117;
  assign n32119 = ~n32116 & n32118;
  assign n32120 = ~n32115 & ~n32119;
  assign n32121 = ~n32114 & n32120;
  assign n32122 = pi788 & ~n32121;
  assign n32123 = ~n16521 & ~n32084;
  assign n32124 = pi625 & n32123;
  assign n32125 = n32049 & ~n32123;
  assign n32126 = ~n32124 & ~n32125;
  assign n32127 = n32089 & ~n32126;
  assign n32128 = ~pi608 & ~n32088;
  assign n32129 = ~n32127 & n32128;
  assign n32130 = pi1153 & n32049;
  assign n32131 = ~n32124 & n32130;
  assign n32132 = pi608 & ~n32090;
  assign n32133 = ~n32131 & n32132;
  assign n32134 = ~n32129 & ~n32133;
  assign n32135 = pi778 & ~n32134;
  assign n32136 = ~pi778 & ~n32125;
  assign n32137 = ~n32135 & ~n32136;
  assign n32138 = ~pi609 & ~n32137;
  assign n32139 = pi609 & ~n32093;
  assign n32140 = ~pi1155 & ~n32139;
  assign n32141 = ~n32138 & n32140;
  assign n32142 = ~pi660 & ~n32054;
  assign n32143 = ~n32141 & n32142;
  assign n32144 = pi609 & ~n32137;
  assign n32145 = ~pi609 & ~n32093;
  assign n32146 = pi1155 & ~n32145;
  assign n32147 = ~n32144 & n32146;
  assign n32148 = pi660 & ~n32056;
  assign n32149 = ~n32147 & n32148;
  assign n32150 = ~n32143 & ~n32149;
  assign n32151 = pi785 & ~n32150;
  assign n32152 = ~pi785 & ~n32137;
  assign n32153 = ~n32151 & ~n32152;
  assign n32154 = ~pi618 & ~n32153;
  assign n32155 = pi618 & n32094;
  assign n32156 = ~pi1154 & ~n32155;
  assign n32157 = ~n32154 & n32156;
  assign n32158 = ~pi627 & ~n32062;
  assign n32159 = ~n32157 & n32158;
  assign n32160 = pi618 & ~n32153;
  assign n32161 = ~pi618 & n32094;
  assign n32162 = pi1154 & ~n32161;
  assign n32163 = ~n32160 & n32162;
  assign n32164 = pi627 & ~n32064;
  assign n32165 = ~n32163 & n32164;
  assign n32166 = ~n32159 & ~n32165;
  assign n32167 = pi781 & ~n32166;
  assign n32168 = ~pi781 & ~n32153;
  assign n32169 = ~n32167 & ~n32168;
  assign n32170 = pi619 & ~n32169;
  assign n32171 = ~pi619 & n32095;
  assign n32172 = pi1159 & ~n32171;
  assign n32173 = ~n32170 & n32172;
  assign n32174 = pi648 & ~n32072;
  assign n32175 = ~n32173 & n32174;
  assign n32176 = ~pi619 & ~n32169;
  assign n32177 = pi619 & n32095;
  assign n32178 = ~pi1159 & ~n32177;
  assign n32179 = ~n32176 & n32178;
  assign n32180 = ~pi648 & ~n32070;
  assign n32181 = ~n32179 & n32180;
  assign n32182 = pi789 & ~n32181;
  assign n32183 = ~n32175 & n32182;
  assign n32184 = ~pi789 & n32169;
  assign n32185 = n17817 & ~n32184;
  assign n32186 = ~n32183 & n32185;
  assign n32187 = ~n32122 & ~n32186;
  assign n32188 = ~n20205 & ~n32187;
  assign n32189 = n17856 & ~n32078;
  assign n32190 = n20693 & n32097;
  assign n32191 = ~n32189 & ~n32190;
  assign n32192 = ~pi629 & ~n32191;
  assign n32193 = n20697 & n32097;
  assign n32194 = n17855 & ~n32078;
  assign n32195 = ~n32193 & ~n32194;
  assign n32196 = pi629 & ~n32195;
  assign n32197 = ~n32192 & ~n32196;
  assign n32198 = pi792 & ~n32197;
  assign n32199 = n20207 & ~n32198;
  assign n32200 = ~n32188 & n32199;
  assign n32201 = ~n32110 & ~n32200;
  assign n32202 = pi644 & n32201;
  assign n32203 = ~pi787 & ~n32098;
  assign n32204 = pi787 & ~n32107;
  assign n32205 = ~n32203 & ~n32204;
  assign n32206 = ~pi644 & n32205;
  assign n32207 = pi715 & ~n32206;
  assign n32208 = ~n32202 & n32207;
  assign n32209 = ~n17652 & ~n32081;
  assign n32210 = n17652 & n32047;
  assign n32211 = ~n32209 & ~n32210;
  assign n32212 = pi644 & ~n32211;
  assign n32213 = ~pi644 & n32047;
  assign n32214 = ~pi715 & ~n32213;
  assign n32215 = ~n32212 & n32214;
  assign n32216 = pi1160 & ~n32215;
  assign n32217 = ~n32208 & n32216;
  assign n32218 = ~pi644 & n32201;
  assign n32219 = pi644 & n32205;
  assign n32220 = ~pi715 & ~n32219;
  assign n32221 = ~n32218 & n32220;
  assign n32222 = ~pi644 & ~n32211;
  assign n32223 = pi644 & n32047;
  assign n32224 = pi715 & ~n32223;
  assign n32225 = ~n32222 & n32224;
  assign n32226 = ~pi1160 & ~n32225;
  assign n32227 = ~n32221 & n32226;
  assign n32228 = ~n32217 & ~n32227;
  assign n32229 = pi790 & ~n32228;
  assign n32230 = ~pi790 & n32201;
  assign n32231 = pi832 & ~n32230;
  assign n32232 = ~n32229 & n32231;
  assign n32233 = ~pi193 & ~n17406;
  assign n32234 = n17539 & ~n32233;
  assign n32235 = pi690 & n3267;
  assign n32236 = n32233 & ~n32235;
  assign n32237 = pi193 & ~n17976;
  assign n32238 = ~pi38 & ~n32237;
  assign n32239 = n3267 & ~n32238;
  assign n32240 = ~pi193 & n17972;
  assign n32241 = ~n32239 & ~n32240;
  assign n32242 = ~pi193 & ~n17280;
  assign n32243 = n17392 & ~n32242;
  assign n32244 = pi690 & ~n32243;
  assign n32245 = ~n32241 & n32244;
  assign n32246 = ~n32236 & ~n32245;
  assign n32247 = ~pi778 & n32246;
  assign n32248 = pi625 & ~n32246;
  assign n32249 = ~pi625 & n32233;
  assign n32250 = pi1153 & ~n32249;
  assign n32251 = ~n32248 & n32250;
  assign n32252 = ~pi625 & ~n32246;
  assign n32253 = pi625 & n32233;
  assign n32254 = ~pi1153 & ~n32253;
  assign n32255 = ~n32252 & n32254;
  assign n32256 = ~n32251 & ~n32255;
  assign n32257 = pi778 & ~n32256;
  assign n32258 = ~n32247 & ~n32257;
  assign n32259 = ~n17466 & ~n32258;
  assign n32260 = n17466 & ~n32233;
  assign n32261 = ~n32259 & ~n32260;
  assign n32262 = ~n17503 & n32261;
  assign n32263 = n17503 & n32233;
  assign n32264 = ~n32262 & ~n32263;
  assign n32265 = ~n17539 & n32264;
  assign n32266 = ~n32234 & ~n32265;
  assign n32267 = ~n17582 & n32266;
  assign n32268 = n17582 & n32233;
  assign n32269 = ~n32267 & ~n32268;
  assign n32270 = ~pi792 & n32269;
  assign n32271 = pi628 & ~n32269;
  assign n32272 = ~pi628 & n32233;
  assign n32273 = pi1156 & ~n32272;
  assign n32274 = ~n32271 & n32273;
  assign n32275 = ~pi628 & ~n32269;
  assign n32276 = pi628 & n32233;
  assign n32277 = ~pi1156 & ~n32276;
  assign n32278 = ~n32275 & n32277;
  assign n32279 = ~n32274 & ~n32278;
  assign n32280 = pi792 & ~n32279;
  assign n32281 = ~n32270 & ~n32280;
  assign n32282 = ~pi647 & ~n32281;
  assign n32283 = pi647 & ~n32233;
  assign n32284 = ~n32282 & ~n32283;
  assign n32285 = ~pi1157 & n32284;
  assign n32286 = pi647 & ~n32281;
  assign n32287 = ~pi647 & ~n32233;
  assign n32288 = ~n32286 & ~n32287;
  assign n32289 = pi1157 & n32288;
  assign n32290 = ~n32285 & ~n32289;
  assign n32291 = pi787 & ~n32290;
  assign n32292 = ~pi787 & n32281;
  assign n32293 = ~n32291 & ~n32292;
  assign n32294 = ~pi644 & ~n32293;
  assign n32295 = pi715 & ~n32294;
  assign n32296 = pi193 & ~n3267;
  assign n32297 = pi739 & n17282;
  assign n32298 = ~n32242 & ~n32297;
  assign n32299 = pi38 & ~n32298;
  assign n32300 = ~pi193 & n17242;
  assign n32301 = pi193 & ~n17275;
  assign n32302 = pi739 & ~n32301;
  assign n32303 = ~n32300 & n32302;
  assign n32304 = ~pi193 & ~pi739;
  assign n32305 = ~n17201 & n32304;
  assign n32306 = ~n32303 & ~n32305;
  assign n32307 = ~pi38 & ~n32306;
  assign n32308 = ~n32299 & ~n32307;
  assign n32309 = n3267 & n32308;
  assign n32310 = ~n32296 & ~n32309;
  assign n32311 = ~n17438 & ~n32310;
  assign n32312 = n17438 & ~n32233;
  assign n32313 = ~n32311 & ~n32312;
  assign n32314 = ~pi785 & ~n32313;
  assign n32315 = ~n17439 & ~n32233;
  assign n32316 = pi609 & n32311;
  assign n32317 = ~n32315 & ~n32316;
  assign n32318 = pi1155 & ~n32317;
  assign n32319 = ~n17451 & ~n32233;
  assign n32320 = ~pi609 & n32311;
  assign n32321 = ~n32319 & ~n32320;
  assign n32322 = ~pi1155 & ~n32321;
  assign n32323 = ~n32318 & ~n32322;
  assign n32324 = pi785 & ~n32323;
  assign n32325 = ~n32314 & ~n32324;
  assign n32326 = ~pi781 & ~n32325;
  assign n32327 = pi618 & n32325;
  assign n32328 = ~pi618 & n32233;
  assign n32329 = pi1154 & ~n32328;
  assign n32330 = ~n32327 & n32329;
  assign n32331 = ~pi618 & n32325;
  assign n32332 = pi618 & n32233;
  assign n32333 = ~pi1154 & ~n32332;
  assign n32334 = ~n32331 & n32333;
  assign n32335 = ~n32330 & ~n32334;
  assign n32336 = pi781 & ~n32335;
  assign n32337 = ~n32326 & ~n32336;
  assign n32338 = ~pi789 & ~n32337;
  assign n32339 = pi619 & n32337;
  assign n32340 = ~pi619 & n32233;
  assign n32341 = pi1159 & ~n32340;
  assign n32342 = ~n32339 & n32341;
  assign n32343 = ~pi619 & n32337;
  assign n32344 = pi619 & n32233;
  assign n32345 = ~pi1159 & ~n32344;
  assign n32346 = ~n32343 & n32345;
  assign n32347 = ~n32342 & ~n32346;
  assign n32348 = pi789 & ~n32347;
  assign n32349 = ~n32338 & ~n32348;
  assign n32350 = ~n17816 & n32349;
  assign n32351 = n17816 & n32233;
  assign n32352 = ~n32350 & ~n32351;
  assign n32353 = ~n17610 & ~n32352;
  assign n32354 = n17610 & n32233;
  assign n32355 = ~n32353 & ~n32354;
  assign n32356 = ~n17652 & ~n32355;
  assign n32357 = n17652 & n32233;
  assign n32358 = ~n32356 & ~n32357;
  assign n32359 = pi644 & ~n32358;
  assign n32360 = ~pi644 & n32233;
  assign n32361 = ~pi715 & ~n32360;
  assign n32362 = ~n32359 & n32361;
  assign n32363 = pi1160 & ~n32362;
  assign n32364 = ~n32295 & n32363;
  assign n32365 = pi644 & ~n32293;
  assign n32366 = ~pi715 & ~n32365;
  assign n32367 = ~pi644 & ~n32358;
  assign n32368 = pi644 & n32233;
  assign n32369 = pi715 & ~n32368;
  assign n32370 = ~n32367 & n32369;
  assign n32371 = ~pi1160 & ~n32370;
  assign n32372 = ~n32366 & n32371;
  assign n32373 = ~n32364 & ~n32372;
  assign n32374 = pi790 & ~n32373;
  assign n32375 = pi644 & n32363;
  assign n32376 = ~pi644 & n32371;
  assign n32377 = pi790 & ~n32376;
  assign n32378 = ~n32375 & n32377;
  assign n32379 = ~n20409 & n32352;
  assign n32380 = ~pi629 & n32274;
  assign n32381 = pi629 & n32278;
  assign n32382 = ~n32380 & ~n32381;
  assign n32383 = ~n32379 & n32382;
  assign n32384 = pi792 & ~n32383;
  assign n32385 = ~pi690 & ~n32308;
  assign n32386 = ~pi193 & n16687;
  assign n32387 = pi193 & n16799;
  assign n32388 = ~pi739 & ~n32387;
  assign n32389 = ~n32386 & n32388;
  assign n32390 = pi193 & n16879;
  assign n32391 = ~pi193 & ~n16944;
  assign n32392 = pi739 & ~n32391;
  assign n32393 = ~n32390 & n32392;
  assign n32394 = pi39 & ~n32393;
  assign n32395 = ~n32389 & n32394;
  assign n32396 = ~pi193 & n17092;
  assign n32397 = pi193 & n17094;
  assign n32398 = pi739 & ~n32397;
  assign n32399 = ~n32396 & n32398;
  assign n32400 = ~pi193 & ~n17088;
  assign n32401 = pi193 & ~n17059;
  assign n32402 = ~pi739 & ~n32401;
  assign n32403 = ~n32400 & n32402;
  assign n32404 = ~n32399 & ~n32403;
  assign n32405 = ~pi39 & ~n32404;
  assign n32406 = ~pi38 & ~n32405;
  assign n32407 = ~n32395 & n32406;
  assign n32408 = ~pi739 & n23906;
  assign n32409 = ~n16905 & ~n32408;
  assign n32410 = ~pi39 & ~n32409;
  assign n32411 = ~pi193 & ~n32410;
  assign n32412 = ~n16787 & ~n32048;
  assign n32413 = pi193 & ~n32412;
  assign n32414 = n6234 & n32413;
  assign n32415 = pi38 & ~n32414;
  assign n32416 = ~n32411 & n32415;
  assign n32417 = pi690 & ~n32416;
  assign n32418 = ~n32407 & n32417;
  assign n32419 = n3267 & ~n32418;
  assign n32420 = ~n32385 & n32419;
  assign n32421 = ~n32296 & ~n32420;
  assign n32422 = ~pi625 & n32421;
  assign n32423 = pi625 & n32310;
  assign n32424 = ~pi1153 & ~n32423;
  assign n32425 = ~n32422 & n32424;
  assign n32426 = ~pi608 & ~n32251;
  assign n32427 = ~n32425 & n32426;
  assign n32428 = pi625 & n32421;
  assign n32429 = ~pi625 & n32310;
  assign n32430 = pi1153 & ~n32429;
  assign n32431 = ~n32428 & n32430;
  assign n32432 = pi608 & ~n32255;
  assign n32433 = ~n32431 & n32432;
  assign n32434 = ~n32427 & ~n32433;
  assign n32435 = pi778 & ~n32434;
  assign n32436 = ~pi778 & n32421;
  assign n32437 = ~n32435 & ~n32436;
  assign n32438 = ~pi609 & ~n32437;
  assign n32439 = pi609 & n32258;
  assign n32440 = ~pi1155 & ~n32439;
  assign n32441 = ~n32438 & n32440;
  assign n32442 = ~pi660 & ~n32318;
  assign n32443 = ~n32441 & n32442;
  assign n32444 = pi609 & ~n32437;
  assign n32445 = ~pi609 & n32258;
  assign n32446 = pi1155 & ~n32445;
  assign n32447 = ~n32444 & n32446;
  assign n32448 = pi660 & ~n32322;
  assign n32449 = ~n32447 & n32448;
  assign n32450 = ~n32443 & ~n32449;
  assign n32451 = pi785 & ~n32450;
  assign n32452 = ~pi785 & ~n32437;
  assign n32453 = ~n32451 & ~n32452;
  assign n32454 = ~pi618 & ~n32453;
  assign n32455 = pi618 & n32261;
  assign n32456 = ~pi1154 & ~n32455;
  assign n32457 = ~n32454 & n32456;
  assign n32458 = ~pi627 & ~n32330;
  assign n32459 = ~n32457 & n32458;
  assign n32460 = pi618 & ~n32453;
  assign n32461 = ~pi618 & n32261;
  assign n32462 = pi1154 & ~n32461;
  assign n32463 = ~n32460 & n32462;
  assign n32464 = pi627 & ~n32334;
  assign n32465 = ~n32463 & n32464;
  assign n32466 = ~n32459 & ~n32465;
  assign n32467 = pi781 & ~n32466;
  assign n32468 = ~pi781 & ~n32453;
  assign n32469 = ~n32467 & ~n32468;
  assign n32470 = pi619 & ~n32469;
  assign n32471 = ~pi619 & ~n32264;
  assign n32472 = pi1159 & ~n32471;
  assign n32473 = ~n32470 & n32472;
  assign n32474 = pi648 & ~n32346;
  assign n32475 = ~n32473 & n32474;
  assign n32476 = ~pi619 & ~n32469;
  assign n32477 = pi619 & ~n32264;
  assign n32478 = ~pi1159 & ~n32477;
  assign n32479 = ~n32476 & n32478;
  assign n32480 = ~pi648 & ~n32342;
  assign n32481 = ~n32479 & n32480;
  assign n32482 = pi789 & ~n32481;
  assign n32483 = ~n32475 & n32482;
  assign n32484 = ~pi789 & n32469;
  assign n32485 = n17817 & ~n32484;
  assign n32486 = ~n32483 & n32485;
  assign n32487 = pi626 & ~n32349;
  assign n32488 = ~pi626 & ~n32233;
  assign n32489 = n17579 & ~n32488;
  assign n32490 = ~n32487 & n32489;
  assign n32491 = n17704 & n32266;
  assign n32492 = ~pi626 & ~n32349;
  assign n32493 = pi626 & ~n32233;
  assign n32494 = n17580 & ~n32493;
  assign n32495 = ~n32492 & n32494;
  assign n32496 = ~n32491 & ~n32495;
  assign n32497 = ~n32490 & n32496;
  assign n32498 = pi788 & ~n32497;
  assign n32499 = ~n20205 & ~n32498;
  assign n32500 = ~n32486 & n32499;
  assign n32501 = ~n32384 & ~n32500;
  assign n32502 = n20207 & ~n32501;
  assign n32503 = ~n20398 & n32355;
  assign n32504 = n17650 & ~n32284;
  assign n32505 = n17649 & ~n32288;
  assign n32506 = ~n32504 & ~n32505;
  assign n32507 = ~n32503 & n32506;
  assign n32508 = pi787 & ~n32507;
  assign n32509 = ~n32502 & ~n32508;
  assign n32510 = ~n32378 & n32509;
  assign n32511 = ~n32374 & ~n32510;
  assign n32512 = ~po1038 & ~n32511;
  assign n32513 = ~pi193 & po1038;
  assign n32514 = ~pi832 & ~n32513;
  assign n32515 = ~n32512 & n32514;
  assign po350 = ~n32232 & ~n32515;
  assign n32517 = pi194 & ~n3267;
  assign n32518 = ~pi194 & n19236;
  assign n32519 = pi194 & ~n24373;
  assign n32520 = ~pi748 & ~n32519;
  assign n32521 = ~n32518 & n32520;
  assign n32522 = pi194 & n19253;
  assign n32523 = ~pi194 & ~n19261;
  assign n32524 = pi748 & ~n32523;
  assign n32525 = ~n32522 & n32524;
  assign n32526 = pi730 & ~n32525;
  assign n32527 = ~n32521 & n32526;
  assign n32528 = ~pi194 & n19223;
  assign n32529 = pi194 & n24271;
  assign n32530 = ~n32528 & ~n32529;
  assign n32531 = pi748 & ~n32530;
  assign n32532 = ~pi194 & ~n17399;
  assign n32533 = ~pi748 & ~n32532;
  assign n32534 = ~n32531 & ~n32533;
  assign n32535 = ~pi730 & n32534;
  assign n32536 = n3267 & ~n32535;
  assign n32537 = ~n32527 & n32536;
  assign n32538 = ~n32517 & ~n32537;
  assign n32539 = ~pi625 & n32538;
  assign n32540 = n3267 & ~n32534;
  assign n32541 = ~n32517 & ~n32540;
  assign n32542 = pi625 & n32541;
  assign n32543 = ~pi1153 & ~n32542;
  assign n32544 = ~n32539 & n32543;
  assign n32545 = pi194 & ~n24209;
  assign n32546 = ~pi194 & n24212;
  assign n32547 = pi730 & ~n32546;
  assign n32548 = ~pi730 & n32532;
  assign n32549 = n3267 & ~n32548;
  assign n32550 = ~n32547 & n32549;
  assign n32551 = ~n32545 & ~n32550;
  assign n32552 = pi625 & n32551;
  assign n32553 = ~pi194 & ~n17406;
  assign n32554 = ~pi625 & n32553;
  assign n32555 = pi1153 & ~n32554;
  assign n32556 = ~n32552 & n32555;
  assign n32557 = ~pi608 & ~n32556;
  assign n32558 = ~n32544 & n32557;
  assign n32559 = pi625 & n32538;
  assign n32560 = ~pi625 & n32541;
  assign n32561 = pi1153 & ~n32560;
  assign n32562 = ~n32559 & n32561;
  assign n32563 = ~pi625 & n32551;
  assign n32564 = pi625 & n32553;
  assign n32565 = ~pi1153 & ~n32564;
  assign n32566 = ~n32563 & n32565;
  assign n32567 = pi608 & ~n32566;
  assign n32568 = ~n32562 & n32567;
  assign n32569 = ~n32558 & ~n32568;
  assign n32570 = pi778 & ~n32569;
  assign n32571 = ~pi778 & n32538;
  assign n32572 = ~n32570 & ~n32571;
  assign n32573 = ~pi609 & ~n32572;
  assign n32574 = ~pi778 & ~n32551;
  assign n32575 = ~n32556 & ~n32566;
  assign n32576 = pi778 & ~n32575;
  assign n32577 = ~n32574 & ~n32576;
  assign n32578 = pi609 & n32577;
  assign n32579 = ~pi1155 & ~n32578;
  assign n32580 = ~n32573 & n32579;
  assign n32581 = ~n17439 & ~n32553;
  assign n32582 = ~n17438 & ~n32541;
  assign n32583 = pi609 & n32582;
  assign n32584 = ~n32581 & ~n32583;
  assign n32585 = pi1155 & ~n32584;
  assign n32586 = ~pi660 & ~n32585;
  assign n32587 = ~n32580 & n32586;
  assign n32588 = pi609 & ~n32572;
  assign n32589 = ~pi609 & n32577;
  assign n32590 = pi1155 & ~n32589;
  assign n32591 = ~n32588 & n32590;
  assign n32592 = ~n17451 & ~n32553;
  assign n32593 = ~pi609 & n32582;
  assign n32594 = ~n32592 & ~n32593;
  assign n32595 = ~pi1155 & ~n32594;
  assign n32596 = pi660 & ~n32595;
  assign n32597 = ~n32591 & n32596;
  assign n32598 = ~n32587 & ~n32597;
  assign n32599 = pi785 & ~n32598;
  assign n32600 = ~pi785 & ~n32572;
  assign n32601 = ~n32599 & ~n32600;
  assign n32602 = ~pi618 & ~n32601;
  assign n32603 = ~n17466 & ~n32577;
  assign n32604 = n17466 & ~n32553;
  assign n32605 = ~n32603 & ~n32604;
  assign n32606 = pi618 & n32605;
  assign n32607 = ~pi1154 & ~n32606;
  assign n32608 = ~n32602 & n32607;
  assign n32609 = n17438 & ~n32553;
  assign n32610 = ~n32582 & ~n32609;
  assign n32611 = ~pi785 & ~n32610;
  assign n32612 = ~n32585 & ~n32595;
  assign n32613 = pi785 & ~n32612;
  assign n32614 = ~n32611 & ~n32613;
  assign n32615 = pi618 & n32614;
  assign n32616 = ~pi618 & n32553;
  assign n32617 = pi1154 & ~n32616;
  assign n32618 = ~n32615 & n32617;
  assign n32619 = ~pi627 & ~n32618;
  assign n32620 = ~n32608 & n32619;
  assign n32621 = pi618 & ~n32601;
  assign n32622 = ~pi618 & n32605;
  assign n32623 = pi1154 & ~n32622;
  assign n32624 = ~n32621 & n32623;
  assign n32625 = ~pi618 & n32614;
  assign n32626 = pi618 & n32553;
  assign n32627 = ~pi1154 & ~n32626;
  assign n32628 = ~n32625 & n32627;
  assign n32629 = pi627 & ~n32628;
  assign n32630 = ~n32624 & n32629;
  assign n32631 = ~n32620 & ~n32630;
  assign n32632 = pi781 & ~n32631;
  assign n32633 = ~pi781 & ~n32601;
  assign n32634 = ~n32632 & ~n32633;
  assign n32635 = ~pi619 & ~n32634;
  assign n32636 = ~n17503 & n32605;
  assign n32637 = n17503 & n32553;
  assign n32638 = ~n32636 & ~n32637;
  assign n32639 = pi619 & ~n32638;
  assign n32640 = ~pi1159 & ~n32639;
  assign n32641 = ~n32635 & n32640;
  assign n32642 = ~pi781 & ~n32614;
  assign n32643 = ~n32618 & ~n32628;
  assign n32644 = pi781 & ~n32643;
  assign n32645 = ~n32642 & ~n32644;
  assign n32646 = pi619 & n32645;
  assign n32647 = ~pi619 & n32553;
  assign n32648 = pi1159 & ~n32647;
  assign n32649 = ~n32646 & n32648;
  assign n32650 = ~pi648 & ~n32649;
  assign n32651 = ~n32641 & n32650;
  assign n32652 = pi619 & ~n32634;
  assign n32653 = ~pi619 & ~n32638;
  assign n32654 = pi1159 & ~n32653;
  assign n32655 = ~n32652 & n32654;
  assign n32656 = ~pi619 & n32645;
  assign n32657 = pi619 & n32553;
  assign n32658 = ~pi1159 & ~n32657;
  assign n32659 = ~n32656 & n32658;
  assign n32660 = pi648 & ~n32659;
  assign n32661 = ~n32655 & n32660;
  assign n32662 = ~n32651 & ~n32661;
  assign n32663 = pi789 & ~n32662;
  assign n32664 = ~pi789 & ~n32634;
  assign n32665 = ~n32663 & ~n32664;
  assign n32666 = ~pi788 & n32665;
  assign n32667 = ~pi626 & n32665;
  assign n32668 = n17539 & ~n32553;
  assign n32669 = ~n17539 & n32638;
  assign n32670 = ~n32668 & ~n32669;
  assign n32671 = pi626 & ~n32670;
  assign n32672 = ~pi641 & ~n32671;
  assign n32673 = ~n32667 & n32672;
  assign n32674 = ~pi789 & ~n32645;
  assign n32675 = ~n32649 & ~n32659;
  assign n32676 = pi789 & ~n32675;
  assign n32677 = ~n32674 & ~n32676;
  assign n32678 = ~pi626 & ~n32677;
  assign n32679 = pi626 & ~n32553;
  assign n32680 = pi641 & ~n32679;
  assign n32681 = ~n32678 & n32680;
  assign n32682 = ~pi1158 & ~n32681;
  assign n32683 = ~n32673 & n32682;
  assign n32684 = pi626 & n32665;
  assign n32685 = ~pi626 & ~n32670;
  assign n32686 = pi641 & ~n32685;
  assign n32687 = ~n32684 & n32686;
  assign n32688 = pi626 & ~n32677;
  assign n32689 = ~pi626 & ~n32553;
  assign n32690 = ~pi641 & ~n32689;
  assign n32691 = ~n32688 & n32690;
  assign n32692 = pi1158 & ~n32691;
  assign n32693 = ~n32687 & n32692;
  assign n32694 = ~n32683 & ~n32693;
  assign n32695 = pi788 & ~n32694;
  assign n32696 = ~n32666 & ~n32695;
  assign n32697 = ~pi628 & n32696;
  assign n32698 = ~n17816 & n32677;
  assign n32699 = n17816 & n32553;
  assign n32700 = ~n32698 & ~n32699;
  assign n32701 = pi628 & ~n32700;
  assign n32702 = ~pi1156 & ~n32701;
  assign n32703 = ~n32697 & n32702;
  assign n32704 = ~n17582 & n32670;
  assign n32705 = n17582 & n32553;
  assign n32706 = ~n32704 & ~n32705;
  assign n32707 = pi628 & ~n32706;
  assign n32708 = ~pi628 & n32553;
  assign n32709 = pi1156 & ~n32708;
  assign n32710 = ~n32707 & n32709;
  assign n32711 = ~pi629 & ~n32710;
  assign n32712 = ~n32703 & n32711;
  assign n32713 = pi628 & n32696;
  assign n32714 = ~pi628 & ~n32700;
  assign n32715 = pi1156 & ~n32714;
  assign n32716 = ~n32713 & n32715;
  assign n32717 = ~pi628 & ~n32706;
  assign n32718 = pi628 & n32553;
  assign n32719 = ~pi1156 & ~n32718;
  assign n32720 = ~n32717 & n32719;
  assign n32721 = pi629 & ~n32720;
  assign n32722 = ~n32716 & n32721;
  assign n32723 = ~n32712 & ~n32722;
  assign n32724 = pi792 & ~n32723;
  assign n32725 = ~pi792 & n32696;
  assign n32726 = ~n32724 & ~n32725;
  assign n32727 = ~pi647 & ~n32726;
  assign n32728 = ~n17610 & ~n32700;
  assign n32729 = n17610 & n32553;
  assign n32730 = ~n32728 & ~n32729;
  assign n32731 = pi647 & ~n32730;
  assign n32732 = ~pi1157 & ~n32731;
  assign n32733 = ~n32727 & n32732;
  assign n32734 = ~pi792 & n32706;
  assign n32735 = ~n32710 & ~n32720;
  assign n32736 = pi792 & ~n32735;
  assign n32737 = ~n32734 & ~n32736;
  assign n32738 = pi647 & n32737;
  assign n32739 = ~pi647 & n32553;
  assign n32740 = pi1157 & ~n32739;
  assign n32741 = ~n32738 & n32740;
  assign n32742 = ~pi630 & ~n32741;
  assign n32743 = ~n32733 & n32742;
  assign n32744 = pi647 & ~n32726;
  assign n32745 = ~pi647 & ~n32730;
  assign n32746 = pi1157 & ~n32745;
  assign n32747 = ~n32744 & n32746;
  assign n32748 = ~pi647 & n32737;
  assign n32749 = pi647 & n32553;
  assign n32750 = ~pi1157 & ~n32749;
  assign n32751 = ~n32748 & n32750;
  assign n32752 = pi630 & ~n32751;
  assign n32753 = ~n32747 & n32752;
  assign n32754 = ~n32743 & ~n32753;
  assign n32755 = pi787 & ~n32754;
  assign n32756 = ~pi787 & ~n32726;
  assign n32757 = ~n32755 & ~n32756;
  assign n32758 = ~pi644 & ~n32757;
  assign n32759 = ~pi787 & ~n32737;
  assign n32760 = ~n32741 & ~n32751;
  assign n32761 = pi787 & ~n32760;
  assign n32762 = ~n32759 & ~n32761;
  assign n32763 = pi644 & n32762;
  assign n32764 = ~pi715 & ~n32763;
  assign n32765 = ~n32758 & n32764;
  assign n32766 = n17652 & ~n32553;
  assign n32767 = ~n17652 & n32730;
  assign n32768 = ~n32766 & ~n32767;
  assign n32769 = ~pi644 & n32768;
  assign n32770 = pi644 & n32553;
  assign n32771 = pi715 & ~n32770;
  assign n32772 = ~n32769 & n32771;
  assign n32773 = ~pi1160 & ~n32772;
  assign n32774 = ~n32765 & n32773;
  assign n32775 = pi644 & ~n32757;
  assign n32776 = ~pi644 & n32762;
  assign n32777 = pi715 & ~n32776;
  assign n32778 = ~n32775 & n32777;
  assign n32779 = pi644 & n32768;
  assign n32780 = ~pi644 & n32553;
  assign n32781 = ~pi715 & ~n32780;
  assign n32782 = ~n32779 & n32781;
  assign n32783 = pi1160 & ~n32782;
  assign n32784 = ~n32778 & n32783;
  assign n32785 = pi790 & ~n32784;
  assign n32786 = ~n32774 & n32785;
  assign n32787 = ~pi790 & n32757;
  assign n32788 = ~po1038 & ~n32787;
  assign n32789 = ~n32786 & n32788;
  assign n32790 = ~pi194 & po1038;
  assign n32791 = ~pi832 & ~n32790;
  assign n32792 = ~n32789 & n32791;
  assign n32793 = ~pi194 & ~n2754;
  assign n32794 = pi748 & n16784;
  assign n32795 = ~n32793 & ~n32794;
  assign n32796 = ~n17706 & ~n32795;
  assign n32797 = ~pi785 & ~n32796;
  assign n32798 = ~n17711 & ~n32795;
  assign n32799 = pi1155 & ~n32798;
  assign n32800 = ~n17714 & n32796;
  assign n32801 = ~pi1155 & ~n32800;
  assign n32802 = ~n32799 & ~n32801;
  assign n32803 = pi785 & ~n32802;
  assign n32804 = ~n32797 & ~n32803;
  assign n32805 = ~pi781 & ~n32804;
  assign n32806 = ~n17721 & n32804;
  assign n32807 = pi1154 & ~n32806;
  assign n32808 = ~n17724 & n32804;
  assign n32809 = ~pi1154 & ~n32808;
  assign n32810 = ~n32807 & ~n32809;
  assign n32811 = pi781 & ~n32810;
  assign n32812 = ~n32805 & ~n32811;
  assign n32813 = ~pi789 & ~n32812;
  assign n32814 = pi619 & n32812;
  assign n32815 = ~pi619 & n32793;
  assign n32816 = pi1159 & ~n32815;
  assign n32817 = ~n32814 & n32816;
  assign n32818 = ~pi619 & n32812;
  assign n32819 = pi619 & n32793;
  assign n32820 = ~pi1159 & ~n32819;
  assign n32821 = ~n32818 & n32820;
  assign n32822 = ~n32817 & ~n32821;
  assign n32823 = pi789 & ~n32822;
  assign n32824 = ~n32813 & ~n32823;
  assign n32825 = ~n17816 & n32824;
  assign n32826 = n17816 & n32793;
  assign n32827 = ~n32825 & ~n32826;
  assign n32828 = ~n17610 & ~n32827;
  assign n32829 = n17610 & n32793;
  assign n32830 = ~n32828 & ~n32829;
  assign n32831 = ~n20398 & n32830;
  assign n32832 = pi730 & n16786;
  assign n32833 = ~n32793 & ~n32832;
  assign n32834 = ~pi778 & n32833;
  assign n32835 = ~pi625 & n32832;
  assign n32836 = ~n32833 & ~n32835;
  assign n32837 = pi1153 & ~n32836;
  assign n32838 = ~pi1153 & ~n32793;
  assign n32839 = ~n32835 & n32838;
  assign n32840 = ~n32837 & ~n32839;
  assign n32841 = pi778 & ~n32840;
  assign n32842 = ~n32834 & ~n32841;
  assign n32843 = ~n17692 & n32842;
  assign n32844 = ~n17694 & n32843;
  assign n32845 = ~n17696 & n32844;
  assign n32846 = ~n17828 & n32845;
  assign n32847 = ~n17859 & n32846;
  assign n32848 = ~pi647 & n32847;
  assign n32849 = pi647 & n32793;
  assign n32850 = ~pi1157 & ~n32849;
  assign n32851 = ~n32848 & n32850;
  assign n32852 = pi647 & ~n32847;
  assign n32853 = ~pi647 & ~n32793;
  assign n32854 = ~n32852 & ~n32853;
  assign n32855 = pi1157 & ~n32854;
  assign n32856 = ~n32851 & ~n32855;
  assign n32857 = ~n17651 & ~n32856;
  assign n32858 = ~n32831 & ~n32857;
  assign n32859 = pi787 & ~n32858;
  assign n32860 = pi626 & ~n32824;
  assign n32861 = ~pi626 & ~n32793;
  assign n32862 = n17579 & ~n32861;
  assign n32863 = ~n32860 & n32862;
  assign n32864 = n17704 & n32845;
  assign n32865 = ~pi626 & ~n32824;
  assign n32866 = pi626 & ~n32793;
  assign n32867 = n17580 & ~n32866;
  assign n32868 = ~n32865 & n32867;
  assign n32869 = ~n32864 & ~n32868;
  assign n32870 = ~n32863 & n32869;
  assign n32871 = pi788 & ~n32870;
  assign n32872 = ~n16521 & ~n32833;
  assign n32873 = pi625 & n32872;
  assign n32874 = n32795 & ~n32872;
  assign n32875 = ~n32873 & ~n32874;
  assign n32876 = n32838 & ~n32875;
  assign n32877 = ~pi608 & ~n32837;
  assign n32878 = ~n32876 & n32877;
  assign n32879 = pi1153 & n32795;
  assign n32880 = ~n32873 & n32879;
  assign n32881 = pi608 & ~n32839;
  assign n32882 = ~n32880 & n32881;
  assign n32883 = ~n32878 & ~n32882;
  assign n32884 = pi778 & ~n32883;
  assign n32885 = ~pi778 & ~n32874;
  assign n32886 = ~n32884 & ~n32885;
  assign n32887 = ~pi609 & ~n32886;
  assign n32888 = pi609 & n32842;
  assign n32889 = ~pi1155 & ~n32888;
  assign n32890 = ~n32887 & n32889;
  assign n32891 = ~pi660 & ~n32799;
  assign n32892 = ~n32890 & n32891;
  assign n32893 = pi609 & ~n32886;
  assign n32894 = ~pi609 & n32842;
  assign n32895 = pi1155 & ~n32894;
  assign n32896 = ~n32893 & n32895;
  assign n32897 = pi660 & ~n32801;
  assign n32898 = ~n32896 & n32897;
  assign n32899 = ~n32892 & ~n32898;
  assign n32900 = pi785 & ~n32899;
  assign n32901 = ~pi785 & ~n32886;
  assign n32902 = ~n32900 & ~n32901;
  assign n32903 = ~pi618 & ~n32902;
  assign n32904 = pi618 & n32843;
  assign n32905 = ~pi1154 & ~n32904;
  assign n32906 = ~n32903 & n32905;
  assign n32907 = ~pi627 & ~n32807;
  assign n32908 = ~n32906 & n32907;
  assign n32909 = pi618 & ~n32902;
  assign n32910 = ~pi618 & n32843;
  assign n32911 = pi1154 & ~n32910;
  assign n32912 = ~n32909 & n32911;
  assign n32913 = pi627 & ~n32809;
  assign n32914 = ~n32912 & n32913;
  assign n32915 = ~n32908 & ~n32914;
  assign n32916 = pi781 & ~n32915;
  assign n32917 = ~pi781 & ~n32902;
  assign n32918 = ~n32916 & ~n32917;
  assign n32919 = pi619 & ~n32918;
  assign n32920 = ~pi619 & n32844;
  assign n32921 = pi1159 & ~n32920;
  assign n32922 = ~n32919 & n32921;
  assign n32923 = pi648 & ~n32821;
  assign n32924 = ~n32922 & n32923;
  assign n32925 = ~pi619 & ~n32918;
  assign n32926 = pi619 & n32844;
  assign n32927 = ~pi1159 & ~n32926;
  assign n32928 = ~n32925 & n32927;
  assign n32929 = ~pi648 & ~n32817;
  assign n32930 = ~n32928 & n32929;
  assign n32931 = pi789 & ~n32930;
  assign n32932 = ~n32924 & n32931;
  assign n32933 = ~pi789 & n32918;
  assign n32934 = n17817 & ~n32933;
  assign n32935 = ~n32932 & n32934;
  assign n32936 = ~n32871 & ~n32935;
  assign n32937 = ~n20205 & ~n32936;
  assign n32938 = n17856 & ~n32827;
  assign n32939 = n20693 & n32846;
  assign n32940 = ~n32938 & ~n32939;
  assign n32941 = ~pi629 & ~n32940;
  assign n32942 = n20697 & n32846;
  assign n32943 = n17855 & ~n32827;
  assign n32944 = ~n32942 & ~n32943;
  assign n32945 = pi629 & ~n32944;
  assign n32946 = ~n32941 & ~n32945;
  assign n32947 = pi792 & ~n32946;
  assign n32948 = n20207 & ~n32947;
  assign n32949 = ~n32937 & n32948;
  assign n32950 = ~n32859 & ~n32949;
  assign n32951 = pi644 & n32950;
  assign n32952 = ~pi787 & ~n32847;
  assign n32953 = pi787 & ~n32856;
  assign n32954 = ~n32952 & ~n32953;
  assign n32955 = ~pi644 & n32954;
  assign n32956 = pi715 & ~n32955;
  assign n32957 = ~n32951 & n32956;
  assign n32958 = ~n17652 & ~n32830;
  assign n32959 = n17652 & n32793;
  assign n32960 = ~n32958 & ~n32959;
  assign n32961 = pi644 & ~n32960;
  assign n32962 = ~pi644 & n32793;
  assign n32963 = ~pi715 & ~n32962;
  assign n32964 = ~n32961 & n32963;
  assign n32965 = pi1160 & ~n32964;
  assign n32966 = ~n32957 & n32965;
  assign n32967 = ~pi644 & n32950;
  assign n32968 = pi644 & n32954;
  assign n32969 = ~pi715 & ~n32968;
  assign n32970 = ~n32967 & n32969;
  assign n32971 = ~pi644 & ~n32960;
  assign n32972 = pi644 & n32793;
  assign n32973 = pi715 & ~n32972;
  assign n32974 = ~n32971 & n32973;
  assign n32975 = ~pi1160 & ~n32974;
  assign n32976 = ~n32970 & n32975;
  assign n32977 = ~n32966 & ~n32976;
  assign n32978 = pi790 & ~n32977;
  assign n32979 = ~pi790 & n32950;
  assign n32980 = pi832 & ~n32979;
  assign n32981 = ~n32978 & n32980;
  assign po351 = ~n32792 & ~n32981;
  assign n32983 = ~n6198 & n16078;
  assign n32984 = ~n11413 & ~n32983;
  assign n32985 = ~n11410 & n16055;
  assign n32986 = n16052 & ~n16433;
  assign n32987 = ~n32985 & ~n32986;
  assign n32988 = n32984 & n32987;
  assign n32989 = pi232 & ~n32988;
  assign n32990 = ~n16430 & ~n32989;
  assign n32991 = pi39 & ~n32990;
  assign n32992 = n13809 & ~n16080;
  assign n32993 = ~pi39 & ~n32992;
  assign n32994 = ~pi138 & n16447;
  assign n32995 = ~pi196 & n32994;
  assign n32996 = pi195 & ~n32995;
  assign n32997 = n10146 & ~n32996;
  assign n32998 = ~n32993 & n32997;
  assign n32999 = ~n32991 & n32998;
  assign n33000 = ~n9358 & ~n16046;
  assign n33001 = pi171 & n13630;
  assign n33002 = ~n33000 & ~n33001;
  assign n33003 = pi299 & ~n33002;
  assign n33004 = pi192 & n16387;
  assign n33005 = ~pi192 & n16375;
  assign n33006 = pi232 & ~n33005;
  assign n33007 = ~n33004 & n33006;
  assign n33008 = ~n33003 & n33007;
  assign n33009 = n16379 & ~n33008;
  assign n33010 = pi192 & n16410;
  assign n33011 = ~pi171 & n9033;
  assign n33012 = ~n16403 & ~n33011;
  assign n33013 = n9028 & ~n33012;
  assign n33014 = n9030 & ~n33013;
  assign n33015 = ~pi192 & n16396;
  assign n33016 = ~n33014 & ~n33015;
  assign n33017 = ~n33010 & n33016;
  assign n33018 = pi232 & ~n33017;
  assign n33019 = ~n16402 & ~n33018;
  assign n33020 = pi39 & ~n33019;
  assign n33021 = n3206 & ~n33020;
  assign n33022 = ~n33009 & n33021;
  assign n33023 = ~pi87 & ~n33022;
  assign n33024 = n16374 & ~n33023;
  assign n33025 = ~pi92 & ~n33024;
  assign n33026 = n16373 & ~n33025;
  assign n33027 = ~pi55 & ~n33026;
  assign n33028 = ~n16425 & ~n33027;
  assign n33029 = n3293 & ~n33028;
  assign n33030 = n9666 & n32996;
  assign n33031 = ~n33029 & n33030;
  assign po352 = n32999 | n33031;
  assign n33033 = ~pi170 & n9033;
  assign n33034 = ~n16403 & ~n33033;
  assign n33035 = n9028 & ~n33034;
  assign n33036 = n9030 & ~n33035;
  assign n33037 = ~n16396 & ~n33036;
  assign n33038 = pi232 & ~n33037;
  assign n33039 = ~n16402 & ~n33038;
  assign n33040 = pi232 & n16410;
  assign n33041 = n33039 & ~n33040;
  assign n33042 = pi39 & ~n33041;
  assign n33043 = ~pi38 & pi194;
  assign n33044 = ~n33042 & n33043;
  assign n33045 = pi39 & ~n33039;
  assign n33046 = ~pi38 & ~pi194;
  assign n33047 = ~n33045 & n33046;
  assign n33048 = ~n33044 & ~n33047;
  assign n33049 = ~n16379 & ~n33048;
  assign n33050 = ~n16387 & n33044;
  assign n33051 = ~n16375 & n33047;
  assign n33052 = ~n33050 & ~n33051;
  assign n33053 = ~n9358 & ~n16155;
  assign n33054 = pi170 & n13630;
  assign n33055 = ~n33053 & ~n33054;
  assign n33056 = pi299 & ~n33055;
  assign n33057 = pi232 & ~n33056;
  assign n33058 = ~n33052 & n33057;
  assign n33059 = ~n33049 & ~n33058;
  assign n33060 = ~pi100 & ~n33059;
  assign n33061 = ~pi87 & ~n33060;
  assign n33062 = n16374 & ~n33061;
  assign n33063 = ~pi92 & ~n33062;
  assign n33064 = n16373 & ~n33063;
  assign n33065 = ~pi55 & ~n33064;
  assign n33066 = ~n16425 & ~n33065;
  assign n33067 = n3293 & ~n33066;
  assign n33068 = n9666 & ~n33067;
  assign n33069 = pi196 & ~n33068;
  assign n33070 = ~pi170 & n9489;
  assign n33071 = ~n16432 & ~n33070;
  assign n33072 = n13047 & ~n33071;
  assign n33073 = n13049 & n16432;
  assign n33074 = pi232 & ~n33073;
  assign n33075 = ~n33072 & n33074;
  assign n33076 = ~n16430 & ~n33075;
  assign n33077 = pi299 & ~n33076;
  assign n33078 = ~n11411 & ~n33077;
  assign n33079 = pi39 & ~n33078;
  assign n33080 = n13809 & ~n16156;
  assign n33081 = ~pi39 & ~n33080;
  assign n33082 = ~pi38 & ~n33081;
  assign n33083 = ~n33079 & n33082;
  assign n33084 = ~pi194 & ~n33083;
  assign n33085 = pi39 & ~n33076;
  assign n33086 = n13809 & n16215;
  assign n33087 = ~pi39 & ~n33086;
  assign n33088 = ~pi38 & ~n33087;
  assign n33089 = ~n33085 & n33088;
  assign n33090 = pi194 & ~n33089;
  assign n33091 = n10143 & ~n33090;
  assign n33092 = ~n33084 & n33091;
  assign n33093 = ~pi196 & ~n33092;
  assign n33094 = ~n32994 & ~n33093;
  assign n33095 = ~n33069 & n33094;
  assign n33096 = pi195 & ~pi196;
  assign n33097 = ~n33068 & n33096;
  assign n33098 = ~n33092 & ~n33096;
  assign n33099 = n32994 & ~n33098;
  assign n33100 = ~n33097 & n33099;
  assign po353 = n33095 | n33100;
  assign n33102 = ~pi767 & pi947;
  assign n33103 = ~pi698 & n20755;
  assign n33104 = ~n33102 & ~n33103;
  assign n33105 = n2754 & ~n33104;
  assign n33106 = ~pi197 & ~n2754;
  assign n33107 = pi832 & ~n33106;
  assign n33108 = ~n33105 & n33107;
  assign n33109 = pi197 & ~n17397;
  assign n33110 = n17280 & ~n33102;
  assign n33111 = pi38 & ~n33110;
  assign n33112 = ~n33109 & n33111;
  assign n33113 = ~pi197 & ~n20840;
  assign n33114 = pi197 & ~n20985;
  assign n33115 = pi299 & ~n33114;
  assign n33116 = ~n33113 & n33115;
  assign n33117 = ~pi197 & ~n17179;
  assign n33118 = n20858 & ~n33117;
  assign n33119 = ~pi767 & ~n33118;
  assign n33120 = ~n33116 & n33119;
  assign n33121 = ~pi197 & pi767;
  assign n33122 = ~n17199 & n33121;
  assign n33123 = pi39 & ~n33122;
  assign n33124 = ~n33120 & n33123;
  assign n33125 = n17120 & n33102;
  assign n33126 = ~pi197 & ~n17120;
  assign n33127 = ~pi39 & ~n33126;
  assign n33128 = ~n33125 & n33127;
  assign n33129 = ~pi38 & ~n33128;
  assign n33130 = ~n33124 & n33129;
  assign n33131 = ~n33112 & ~n33130;
  assign n33132 = pi698 & ~n33131;
  assign n33133 = ~n20906 & n33128;
  assign n33134 = ~pi197 & n20924;
  assign n33135 = pi197 & n20938;
  assign n33136 = ~pi767 & ~n33135;
  assign n33137 = ~n33134 & n33136;
  assign n33138 = ~pi197 & n20884;
  assign n33139 = pi197 & n20900;
  assign n33140 = pi299 & ~n33139;
  assign n33141 = ~n33138 & n33140;
  assign n33142 = n20903 & ~n33117;
  assign n33143 = pi767 & ~n33142;
  assign n33144 = ~n33141 & n33143;
  assign n33145 = pi39 & ~n33144;
  assign n33146 = ~n33137 & n33145;
  assign n33147 = ~n33133 & ~n33146;
  assign n33148 = ~pi38 & ~n33147;
  assign n33149 = pi767 & pi947;
  assign n33150 = ~pi39 & ~n33149;
  assign n33151 = n21067 & n33150;
  assign n33152 = ~pi197 & ~n17280;
  assign n33153 = pi38 & ~n33152;
  assign n33154 = ~n33151 & n33153;
  assign n33155 = ~pi698 & ~n33154;
  assign n33156 = ~n33148 & n33155;
  assign n33157 = ~n33132 & ~n33156;
  assign n33158 = n10143 & ~n33157;
  assign n33159 = ~pi197 & ~n10143;
  assign n33160 = ~pi832 & ~n33159;
  assign n33161 = ~n33158 & n33160;
  assign po354 = ~n33108 & ~n33161;
  assign n33163 = n3181 & ~n17120;
  assign n33164 = n18723 & ~n33163;
  assign n33165 = pi198 & ~n33164;
  assign n33166 = pi198 & ~n16812;
  assign n33167 = ~n6215 & n33166;
  assign n33168 = pi198 & ~n16518;
  assign n33169 = ~po1101 & ~n33168;
  assign n33170 = pi198 & ~n16621;
  assign n33171 = po1101 & ~n33170;
  assign n33172 = ~n33169 & ~n33171;
  assign n33173 = n6215 & n33172;
  assign n33174 = ~n3052 & ~n33173;
  assign n33175 = ~n33167 & n33174;
  assign n33176 = n3052 & ~n33168;
  assign n33177 = ~pi223 & ~n33176;
  assign n33178 = ~n33175 & n33177;
  assign n33179 = pi198 & ~n16569;
  assign n33180 = ~n33169 & n33179;
  assign n33181 = pi198 & n16585;
  assign n33182 = ~n6215 & n33181;
  assign n33183 = ~n33180 & ~n33182;
  assign n33184 = pi223 & ~n33183;
  assign n33185 = ~pi299 & ~n33184;
  assign n33186 = ~n33178 & n33185;
  assign n33187 = ~n6189 & n33166;
  assign n33188 = n6189 & n33172;
  assign n33189 = ~n3329 & ~n33188;
  assign n33190 = ~n33187 & n33189;
  assign n33191 = n3329 & ~n33168;
  assign n33192 = ~pi215 & ~n33191;
  assign n33193 = ~n33190 & n33192;
  assign n33194 = ~n6189 & n33181;
  assign n33195 = ~n33180 & ~n33194;
  assign n33196 = pi215 & ~n33195;
  assign n33197 = pi299 & ~n33196;
  assign n33198 = ~n33193 & n33197;
  assign n33199 = n3267 & n10922;
  assign n33200 = ~n33198 & n33199;
  assign n33201 = ~n33186 & n33200;
  assign n33202 = ~n33165 & ~n33201;
  assign n33203 = n17610 & ~n33202;
  assign n33204 = pi198 & ~n3267;
  assign n33205 = pi198 & ~n17026;
  assign n33206 = pi603 & pi633;
  assign n33207 = ~n33205 & ~n33206;
  assign n33208 = pi198 & ~n17018;
  assign n33209 = ~pi198 & n17083;
  assign n33210 = ~n33208 & ~n33209;
  assign n33211 = n33206 & n33210;
  assign n33212 = ~n33207 & ~n33211;
  assign n33213 = pi299 & n33212;
  assign n33214 = ~n17030 & ~n17034;
  assign n33215 = pi633 & ~n33214;
  assign n33216 = ~n17062 & ~n33215;
  assign n33217 = ~n17039 & ~n33216;
  assign n33218 = ~pi299 & n33217;
  assign n33219 = ~pi39 & ~n33218;
  assign n33220 = ~n33213 & n33219;
  assign n33221 = pi633 & n16518;
  assign n33222 = ~n16520 & n33221;
  assign n33223 = ~n33168 & ~n33222;
  assign n33224 = pi603 & ~n33223;
  assign n33225 = ~pi603 & n33168;
  assign n33226 = ~n33224 & ~n33225;
  assign n33227 = ~n16592 & n33226;
  assign n33228 = n6162 & ~n33223;
  assign n33229 = ~n16542 & n33222;
  assign n33230 = ~n33179 & ~n33229;
  assign n33231 = ~n33228 & n33230;
  assign n33232 = pi603 & ~n33231;
  assign n33233 = n16592 & ~n33225;
  assign n33234 = ~n33232 & n33233;
  assign n33235 = ~n33227 & ~n33234;
  assign n33236 = ~n6160 & n33235;
  assign n33237 = ~n33179 & ~n33232;
  assign n33238 = n6160 & ~n33237;
  assign n33239 = ~n33236 & ~n33238;
  assign n33240 = n6189 & n33239;
  assign n33241 = pi633 & n16848;
  assign n33242 = ~n33181 & ~n33241;
  assign n33243 = ~n6160 & ~n33242;
  assign n33244 = pi198 & n16542;
  assign n33245 = ~n33229 & ~n33244;
  assign n33246 = n17220 & ~n33245;
  assign n33247 = ~n33243 & ~n33246;
  assign n33248 = ~n6189 & n33247;
  assign n33249 = pi215 & ~n33248;
  assign n33250 = ~n33240 & n33249;
  assign n33251 = pi198 & n16619;
  assign n33252 = pi633 & n16656;
  assign n33253 = ~n33251 & ~n33252;
  assign n33254 = ~n6162 & ~n33253;
  assign n33255 = ~n33228 & ~n33254;
  assign n33256 = pi603 & ~n33255;
  assign n33257 = ~pi642 & ~n33256;
  assign n33258 = pi642 & ~n33224;
  assign n33259 = n6156 & ~n33258;
  assign n33260 = ~n33257 & n33259;
  assign n33261 = ~n6156 & n33224;
  assign n33262 = ~n33225 & ~n33261;
  assign n33263 = ~n33260 & n33262;
  assign n33264 = ~n6160 & n33263;
  assign n33265 = ~pi603 & n33170;
  assign n33266 = n6160 & ~n33265;
  assign n33267 = ~n33256 & n33266;
  assign n33268 = ~n33264 & ~n33267;
  assign n33269 = n6189 & n33268;
  assign n33270 = n6162 & n33253;
  assign n33271 = ~n6162 & n33223;
  assign n33272 = pi603 & ~n16592;
  assign n33273 = ~n33271 & n33272;
  assign n33274 = ~n33270 & n33273;
  assign n33275 = pi603 & ~n33253;
  assign n33276 = n16592 & n33275;
  assign n33277 = ~pi603 & n16649;
  assign n33278 = pi198 & n33277;
  assign n33279 = ~n33276 & ~n33278;
  assign n33280 = ~n33274 & n33279;
  assign n33281 = ~n6160 & n33280;
  assign n33282 = n6160 & ~n33251;
  assign n33283 = ~n33275 & n33282;
  assign n33284 = ~n33281 & ~n33283;
  assign n33285 = ~n6189 & n33284;
  assign n33286 = ~n3329 & ~n33285;
  assign n33287 = ~n33269 & n33286;
  assign n33288 = n3329 & n33226;
  assign n33289 = ~pi215 & ~n33288;
  assign n33290 = ~n33287 & n33289;
  assign n33291 = ~n33250 & ~n33290;
  assign n33292 = pi299 & ~n33291;
  assign n33293 = n6215 & n33239;
  assign n33294 = ~n6215 & n33247;
  assign n33295 = pi223 & ~n33294;
  assign n33296 = ~n33293 & n33295;
  assign n33297 = n6215 & n33268;
  assign n33298 = ~n6215 & n33284;
  assign n33299 = ~n3052 & ~n33298;
  assign n33300 = ~n33297 & n33299;
  assign n33301 = n3052 & n33226;
  assign n33302 = ~pi223 & ~n33301;
  assign n33303 = ~n33300 & n33302;
  assign n33304 = ~n33296 & ~n33303;
  assign n33305 = ~pi299 & ~n33304;
  assign n33306 = pi39 & ~n33305;
  assign n33307 = ~n33292 & n33306;
  assign n33308 = ~n33220 & ~n33307;
  assign n33309 = ~pi38 & ~n33308;
  assign n33310 = pi39 & pi198;
  assign n33311 = pi38 & ~n33310;
  assign n33312 = pi198 & ~n16529;
  assign n33313 = pi633 & n16521;
  assign n33314 = n16529 & n33313;
  assign n33315 = ~n33312 & ~n33314;
  assign n33316 = ~pi39 & ~n33315;
  assign n33317 = n33311 & ~n33316;
  assign n33318 = n3267 & ~n33317;
  assign n33319 = ~n33309 & n33318;
  assign n33320 = ~n33204 & ~n33319;
  assign n33321 = ~n17438 & ~n33320;
  assign n33322 = n17438 & ~n33202;
  assign n33323 = ~n33321 & ~n33322;
  assign n33324 = ~pi785 & ~n33323;
  assign n33325 = ~n17439 & ~n33202;
  assign n33326 = pi609 & n33321;
  assign n33327 = ~n33325 & ~n33326;
  assign n33328 = pi1155 & ~n33327;
  assign n33329 = ~n17451 & ~n33202;
  assign n33330 = ~pi609 & n33321;
  assign n33331 = ~n33329 & ~n33330;
  assign n33332 = ~pi1155 & ~n33331;
  assign n33333 = ~n33328 & ~n33332;
  assign n33334 = pi785 & ~n33333;
  assign n33335 = ~n33324 & ~n33334;
  assign n33336 = ~pi781 & ~n33335;
  assign n33337 = pi618 & n33335;
  assign n33338 = ~pi618 & n33202;
  assign n33339 = pi1154 & ~n33338;
  assign n33340 = ~n33337 & n33339;
  assign n33341 = ~pi618 & n33335;
  assign n33342 = pi618 & n33202;
  assign n33343 = ~pi1154 & ~n33342;
  assign n33344 = ~n33341 & n33343;
  assign n33345 = ~n33340 & ~n33344;
  assign n33346 = pi781 & ~n33345;
  assign n33347 = ~n33336 & ~n33346;
  assign n33348 = ~pi789 & ~n33347;
  assign n33349 = pi619 & n33347;
  assign n33350 = ~pi619 & n33202;
  assign n33351 = pi1159 & ~n33350;
  assign n33352 = ~n33349 & n33351;
  assign n33353 = ~pi619 & n33347;
  assign n33354 = pi619 & n33202;
  assign n33355 = ~pi1159 & ~n33354;
  assign n33356 = ~n33353 & n33355;
  assign n33357 = ~n33352 & ~n33356;
  assign n33358 = pi789 & ~n33357;
  assign n33359 = ~n33348 & ~n33358;
  assign n33360 = ~n17816 & n33359;
  assign n33361 = n17816 & n33202;
  assign n33362 = ~n33360 & ~n33361;
  assign n33363 = ~n17610 & n33362;
  assign n33364 = ~n33203 & ~n33363;
  assign n33365 = ~n20398 & ~n33364;
  assign n33366 = ~n19126 & n33202;
  assign n33367 = n17503 & ~n33202;
  assign n33368 = ~n16689 & ~n33168;
  assign n33369 = pi634 & ~n33368;
  assign n33370 = ~n33168 & ~n33369;
  assign n33371 = ~n6162 & n33370;
  assign n33372 = pi634 & n16690;
  assign n33373 = ~n33251 & ~n33372;
  assign n33374 = n6162 & n33373;
  assign n33375 = ~n33371 & ~n33374;
  assign n33376 = ~n6157 & ~n33375;
  assign n33377 = n6157 & n33373;
  assign n33378 = n16513 & ~n33377;
  assign n33379 = ~n33376 & n33378;
  assign n33380 = pi198 & n16655;
  assign n33381 = n6160 & ~n33373;
  assign n33382 = ~n33380 & ~n33381;
  assign n33383 = ~n33379 & n33382;
  assign n33384 = ~n6215 & ~n33383;
  assign n33385 = ~n6157 & n33370;
  assign n33386 = n16513 & ~n33385;
  assign n33387 = n6162 & ~n33370;
  assign n33388 = ~n6162 & ~n33373;
  assign n33389 = ~n33387 & ~n33388;
  assign n33390 = n6157 & n33389;
  assign n33391 = n33386 & ~n33390;
  assign n33392 = n6160 & ~n33389;
  assign n33393 = n6157 & ~n33170;
  assign n33394 = ~n6157 & ~n33168;
  assign n33395 = ~pi680 & ~n33394;
  assign n33396 = ~n33393 & n33395;
  assign n33397 = ~n33392 & ~n33396;
  assign n33398 = ~n33391 & n33397;
  assign n33399 = n6215 & ~n33398;
  assign n33400 = ~n3052 & ~n33399;
  assign n33401 = ~n33384 & n33400;
  assign n33402 = pi680 & n33369;
  assign n33403 = ~n33168 & ~n33402;
  assign n33404 = n3052 & n33403;
  assign n33405 = ~pi223 & ~n33404;
  assign n33406 = ~n33401 & n33405;
  assign n33407 = pi634 & ~n16542;
  assign n33408 = n16689 & n33407;
  assign n33409 = ~n33244 & ~n33408;
  assign n33410 = ~n6162 & ~n33409;
  assign n33411 = ~n33387 & ~n33410;
  assign n33412 = n6157 & n33411;
  assign n33413 = n33386 & ~n33412;
  assign n33414 = ~pi680 & n33181;
  assign n33415 = n33179 & n33414;
  assign n33416 = n6160 & ~n33411;
  assign n33417 = ~n33415 & ~n33416;
  assign n33418 = ~n33413 & n33417;
  assign n33419 = n6215 & n33418;
  assign n33420 = n6162 & n33409;
  assign n33421 = ~n33371 & ~n33420;
  assign n33422 = ~n6157 & ~n33421;
  assign n33423 = n6157 & n33409;
  assign n33424 = n16513 & ~n33423;
  assign n33425 = ~n33422 & n33424;
  assign n33426 = n6160 & ~n33409;
  assign n33427 = ~n33414 & ~n33426;
  assign n33428 = ~n33425 & n33427;
  assign n33429 = ~n6215 & n33428;
  assign n33430 = pi223 & ~n33429;
  assign n33431 = ~n33419 & n33430;
  assign n33432 = ~pi299 & ~n33431;
  assign n33433 = ~n33406 & n33432;
  assign n33434 = n6189 & ~n33398;
  assign n33435 = ~n6189 & ~n33383;
  assign n33436 = ~n3329 & ~n33435;
  assign n33437 = ~n33434 & n33436;
  assign n33438 = n3329 & n33403;
  assign n33439 = ~pi215 & ~n33438;
  assign n33440 = ~n33437 & n33439;
  assign n33441 = n6189 & n33418;
  assign n33442 = ~n6189 & n33428;
  assign n33443 = pi215 & ~n33442;
  assign n33444 = ~n33441 & n33443;
  assign n33445 = pi299 & ~n33444;
  assign n33446 = ~n33440 & n33445;
  assign n33447 = ~n33433 & ~n33446;
  assign n33448 = pi39 & ~n33447;
  assign n33449 = pi634 & pi680;
  assign n33450 = ~pi198 & n17054;
  assign n33451 = pi198 & ~n17074;
  assign n33452 = ~n33450 & ~n33451;
  assign n33453 = n33449 & ~n33452;
  assign n33454 = n33205 & ~n33449;
  assign n33455 = ~n33453 & ~n33454;
  assign n33456 = pi299 & ~n33455;
  assign n33457 = pi198 & n17064;
  assign n33458 = ~n17045 & n33449;
  assign n33459 = ~n33457 & n33458;
  assign n33460 = ~n17062 & ~n33459;
  assign n33461 = ~pi299 & ~n33460;
  assign n33462 = ~pi39 & ~n33461;
  assign n33463 = ~n33456 & n33462;
  assign n33464 = ~n33448 & ~n33463;
  assign n33465 = ~pi38 & ~n33464;
  assign n33466 = pi634 & n16785;
  assign n33467 = n16529 & n33466;
  assign n33468 = ~n33312 & ~n33467;
  assign n33469 = ~pi39 & ~n33468;
  assign n33470 = n33311 & ~n33469;
  assign n33471 = n3267 & ~n33470;
  assign n33472 = ~n33465 & n33471;
  assign n33473 = ~n33204 & ~n33472;
  assign n33474 = ~pi778 & ~n33473;
  assign n33475 = pi625 & n33473;
  assign n33476 = ~pi625 & n33202;
  assign n33477 = pi1153 & ~n33476;
  assign n33478 = ~n33475 & n33477;
  assign n33479 = ~pi625 & n33473;
  assign n33480 = pi625 & n33202;
  assign n33481 = ~pi1153 & ~n33480;
  assign n33482 = ~n33479 & n33481;
  assign n33483 = ~n33478 & ~n33482;
  assign n33484 = pi778 & ~n33483;
  assign n33485 = ~n33474 & ~n33484;
  assign n33486 = ~n17466 & n33485;
  assign n33487 = n17466 & n33202;
  assign n33488 = ~n33486 & ~n33487;
  assign n33489 = ~n17503 & n33488;
  assign n33490 = ~n33367 & ~n33489;
  assign n33491 = ~n17539 & n33490;
  assign n33492 = ~n17582 & n33491;
  assign n33493 = ~n33366 & ~n33492;
  assign n33494 = ~pi792 & n33493;
  assign n33495 = pi628 & ~n33493;
  assign n33496 = ~pi628 & n33202;
  assign n33497 = ~n33495 & ~n33496;
  assign n33498 = pi1156 & n33497;
  assign n33499 = ~pi628 & ~n33493;
  assign n33500 = pi628 & n33202;
  assign n33501 = ~pi1156 & ~n33500;
  assign n33502 = ~n33499 & n33501;
  assign n33503 = ~n33498 & ~n33502;
  assign n33504 = pi792 & ~n33503;
  assign n33505 = ~n33494 & ~n33504;
  assign n33506 = ~pi647 & n33505;
  assign n33507 = pi647 & n33202;
  assign n33508 = ~pi1157 & ~n33507;
  assign n33509 = ~n33506 & n33508;
  assign n33510 = pi647 & ~n33505;
  assign n33511 = ~pi647 & ~n33202;
  assign n33512 = ~n33510 & ~n33511;
  assign n33513 = pi1157 & ~n33512;
  assign n33514 = ~n33509 & ~n33513;
  assign n33515 = ~n17651 & ~n33514;
  assign n33516 = ~n33365 & ~n33515;
  assign n33517 = pi787 & ~n33516;
  assign n33518 = ~n20409 & n33362;
  assign n33519 = pi629 & n33502;
  assign n33520 = n17607 & n33497;
  assign n33521 = ~n33519 & ~n33520;
  assign n33522 = ~n33518 & n33521;
  assign n33523 = pi792 & ~n33522;
  assign n33524 = pi626 & ~n33359;
  assign n33525 = ~pi626 & ~n33202;
  assign n33526 = n17579 & ~n33525;
  assign n33527 = ~n33524 & n33526;
  assign n33528 = n17539 & n33202;
  assign n33529 = ~n33491 & ~n33528;
  assign n33530 = n17704 & ~n33529;
  assign n33531 = ~pi626 & ~n33359;
  assign n33532 = pi626 & ~n33202;
  assign n33533 = n17580 & ~n33532;
  assign n33534 = ~n33531 & n33533;
  assign n33535 = ~n33530 & ~n33534;
  assign n33536 = ~n33527 & n33535;
  assign n33537 = pi788 & ~n33536;
  assign n33538 = ~pi603 & ~n33452;
  assign n33539 = pi198 & ~pi665;
  assign n33540 = pi633 & ~n33539;
  assign n33541 = ~n33450 & n33540;
  assign n33542 = n33210 & n33541;
  assign n33543 = ~n17083 & n33451;
  assign n33544 = ~pi198 & ~pi665;
  assign n33545 = n17018 & n33544;
  assign n33546 = ~pi633 & ~n33545;
  assign n33547 = ~n33543 & n33546;
  assign n33548 = pi603 & ~n33547;
  assign n33549 = ~n33542 & n33548;
  assign n33550 = ~n33538 & ~n33549;
  assign n33551 = n33449 & ~n33550;
  assign n33552 = n33212 & ~n33449;
  assign n33553 = pi299 & ~n33552;
  assign n33554 = ~n33551 & n33553;
  assign n33555 = ~pi634 & n17062;
  assign n33556 = pi634 & n17065;
  assign n33557 = ~n17036 & n33556;
  assign n33558 = ~n33555 & ~n33557;
  assign n33559 = ~pi633 & ~n33558;
  assign n33560 = pi198 & ~pi633;
  assign n33561 = pi634 & ~pi665;
  assign n33562 = ~n33560 & n33561;
  assign n33563 = ~n17029 & n33562;
  assign n33564 = pi603 & ~n33563;
  assign n33565 = ~n33215 & n33564;
  assign n33566 = ~n33559 & n33565;
  assign n33567 = ~pi603 & n33460;
  assign n33568 = pi680 & ~n33567;
  assign n33569 = ~n33566 & n33568;
  assign n33570 = ~pi680 & n33217;
  assign n33571 = ~pi299 & ~n33570;
  assign n33572 = ~n33569 & n33571;
  assign n33573 = ~n33554 & ~n33572;
  assign n33574 = ~pi39 & ~n33573;
  assign n33575 = ~pi680 & n33263;
  assign n33576 = n16717 & n33561;
  assign n33577 = n33223 & ~n33576;
  assign n33578 = n6162 & ~n33577;
  assign n33579 = pi634 & n16696;
  assign n33580 = n33253 & ~n33579;
  assign n33581 = ~n6162 & ~n33580;
  assign n33582 = ~n33578 & ~n33581;
  assign n33583 = pi603 & ~n33582;
  assign n33584 = ~pi642 & n33583;
  assign n33585 = ~pi603 & ~n33370;
  assign n33586 = pi603 & ~n33577;
  assign n33587 = pi642 & n33586;
  assign n33588 = ~n33585 & ~n33587;
  assign n33589 = ~n33584 & n33588;
  assign n33590 = n6156 & ~n33589;
  assign n33591 = ~n33585 & ~n33586;
  assign n33592 = ~n6156 & ~n33591;
  assign n33593 = ~n16512 & ~n33592;
  assign n33594 = ~n33590 & n33593;
  assign n33595 = ~pi603 & ~n33389;
  assign n33596 = n16512 & ~n33595;
  assign n33597 = ~n33583 & n33596;
  assign n33598 = ~n33594 & ~n33597;
  assign n33599 = pi680 & ~n33598;
  assign n33600 = ~n33575 & ~n33599;
  assign n33601 = n6189 & n33600;
  assign n33602 = ~pi603 & n33375;
  assign n33603 = ~n16592 & n33586;
  assign n33604 = ~n33273 & ~n33603;
  assign n33605 = ~n6157 & n33604;
  assign n33606 = ~n6162 & ~n33604;
  assign n33607 = n33580 & ~n33606;
  assign n33608 = ~n33605 & ~n33607;
  assign n33609 = ~n33602 & ~n33608;
  assign n33610 = n16513 & ~n33609;
  assign n33611 = ~pi680 & ~n33280;
  assign n33612 = ~n16521 & ~n33373;
  assign n33613 = ~n33275 & ~n33612;
  assign n33614 = n6160 & ~n33613;
  assign n33615 = ~n33611 & ~n33614;
  assign n33616 = ~n33610 & n33615;
  assign n33617 = ~n6189 & ~n33616;
  assign n33618 = ~n3329 & ~n33617;
  assign n33619 = ~n33601 & n33618;
  assign n33620 = n16667 & n33369;
  assign n33621 = n33226 & ~n33620;
  assign n33622 = n3329 & n33621;
  assign n33623 = ~pi215 & ~n33622;
  assign n33624 = ~n33619 & n33623;
  assign n33625 = n16746 & n33544;
  assign n33626 = n16520 & n33539;
  assign n33627 = ~n33244 & ~n33626;
  assign n33628 = ~n33625 & n33627;
  assign n33629 = pi634 & ~n33628;
  assign n33630 = ~pi634 & n33244;
  assign n33631 = ~n33229 & ~n33630;
  assign n33632 = ~n33629 & n33631;
  assign n33633 = ~n6162 & ~n33632;
  assign n33634 = ~n33578 & ~n33633;
  assign n33635 = pi603 & ~n33634;
  assign n33636 = n16592 & ~n33585;
  assign n33637 = ~n33635 & n33636;
  assign n33638 = ~n16592 & n33591;
  assign n33639 = n16513 & ~n33638;
  assign n33640 = ~n33637 & n33639;
  assign n33641 = ~pi680 & n33235;
  assign n33642 = ~pi603 & ~n33411;
  assign n33643 = ~n33635 & ~n33642;
  assign n33644 = n6160 & ~n33643;
  assign n33645 = ~n33641 & ~n33644;
  assign n33646 = ~n33640 & n33645;
  assign n33647 = n6189 & n33646;
  assign n33648 = ~pi603 & n33421;
  assign n33649 = ~n33606 & ~n33648;
  assign n33650 = pi603 & ~n33632;
  assign n33651 = ~n16592 & n33604;
  assign n33652 = n33650 & ~n33651;
  assign n33653 = n33649 & ~n33652;
  assign n33654 = n16513 & ~n33653;
  assign n33655 = ~pi680 & ~n33242;
  assign n33656 = ~pi603 & ~n33409;
  assign n33657 = ~n33650 & ~n33656;
  assign n33658 = n6160 & ~n33657;
  assign n33659 = ~n33655 & ~n33658;
  assign n33660 = ~n33654 & n33659;
  assign n33661 = ~n6189 & n33660;
  assign n33662 = pi215 & ~n33661;
  assign n33663 = ~n33647 & n33662;
  assign n33664 = ~n33624 & ~n33663;
  assign n33665 = pi299 & ~n33664;
  assign n33666 = n6215 & n33600;
  assign n33667 = ~n6215 & ~n33616;
  assign n33668 = ~n3052 & ~n33667;
  assign n33669 = ~n33666 & n33668;
  assign n33670 = n3052 & n33621;
  assign n33671 = ~pi223 & ~n33670;
  assign n33672 = ~n33669 & n33671;
  assign n33673 = n6215 & n33646;
  assign n33674 = ~n6215 & n33660;
  assign n33675 = pi223 & ~n33674;
  assign n33676 = ~n33673 & n33675;
  assign n33677 = ~n33672 & ~n33676;
  assign n33678 = ~pi299 & ~n33677;
  assign n33679 = pi39 & ~n33678;
  assign n33680 = ~n33665 & n33679;
  assign n33681 = ~n33574 & ~n33680;
  assign n33682 = ~pi38 & ~n33681;
  assign n33683 = pi634 & n17940;
  assign n33684 = ~n33316 & ~n33683;
  assign n33685 = n33311 & n33684;
  assign n33686 = n3267 & ~n33685;
  assign n33687 = ~n33682 & n33686;
  assign n33688 = ~n33204 & ~n33687;
  assign n33689 = ~pi625 & n33688;
  assign n33690 = pi625 & n33320;
  assign n33691 = ~pi1153 & ~n33690;
  assign n33692 = ~n33689 & n33691;
  assign n33693 = ~pi608 & ~n33478;
  assign n33694 = ~n33692 & n33693;
  assign n33695 = pi625 & n33688;
  assign n33696 = ~pi625 & n33320;
  assign n33697 = pi1153 & ~n33696;
  assign n33698 = ~n33695 & n33697;
  assign n33699 = pi608 & ~n33482;
  assign n33700 = ~n33698 & n33699;
  assign n33701 = ~n33694 & ~n33700;
  assign n33702 = pi778 & ~n33701;
  assign n33703 = ~pi778 & n33688;
  assign n33704 = ~n33702 & ~n33703;
  assign n33705 = ~pi609 & ~n33704;
  assign n33706 = pi609 & n33485;
  assign n33707 = ~pi1155 & ~n33706;
  assign n33708 = ~n33705 & n33707;
  assign n33709 = ~pi660 & ~n33328;
  assign n33710 = ~n33708 & n33709;
  assign n33711 = pi609 & ~n33704;
  assign n33712 = ~pi609 & n33485;
  assign n33713 = pi1155 & ~n33712;
  assign n33714 = ~n33711 & n33713;
  assign n33715 = pi660 & ~n33332;
  assign n33716 = ~n33714 & n33715;
  assign n33717 = ~n33710 & ~n33716;
  assign n33718 = pi785 & ~n33717;
  assign n33719 = ~pi785 & ~n33704;
  assign n33720 = ~n33718 & ~n33719;
  assign n33721 = ~pi618 & ~n33720;
  assign n33722 = pi618 & ~n33488;
  assign n33723 = ~pi1154 & ~n33722;
  assign n33724 = ~n33721 & n33723;
  assign n33725 = ~pi627 & ~n33340;
  assign n33726 = ~n33724 & n33725;
  assign n33727 = pi618 & ~n33720;
  assign n33728 = ~pi618 & ~n33488;
  assign n33729 = pi1154 & ~n33728;
  assign n33730 = ~n33727 & n33729;
  assign n33731 = pi627 & ~n33344;
  assign n33732 = ~n33730 & n33731;
  assign n33733 = ~n33726 & ~n33732;
  assign n33734 = pi781 & ~n33733;
  assign n33735 = ~pi781 & ~n33720;
  assign n33736 = ~n33734 & ~n33735;
  assign n33737 = pi619 & ~n33736;
  assign n33738 = ~pi619 & n33490;
  assign n33739 = pi1159 & ~n33738;
  assign n33740 = ~n33737 & n33739;
  assign n33741 = pi648 & ~n33356;
  assign n33742 = ~n33740 & n33741;
  assign n33743 = ~pi619 & ~n33736;
  assign n33744 = pi619 & n33490;
  assign n33745 = ~pi1159 & ~n33744;
  assign n33746 = ~n33743 & n33745;
  assign n33747 = ~pi648 & ~n33352;
  assign n33748 = ~n33746 & n33747;
  assign n33749 = pi789 & ~n33748;
  assign n33750 = ~n33742 & n33749;
  assign n33751 = ~pi789 & n33736;
  assign n33752 = n17817 & ~n33751;
  assign n33753 = ~n33750 & n33752;
  assign n33754 = ~n33537 & ~n33753;
  assign n33755 = ~n33523 & ~n33754;
  assign n33756 = n20205 & n33522;
  assign n33757 = n20207 & ~n33756;
  assign n33758 = ~n33755 & n33757;
  assign n33759 = ~n33517 & ~n33758;
  assign n33760 = ~pi790 & ~n33759;
  assign n33761 = ~pi644 & n33759;
  assign n33762 = ~pi787 & ~n33505;
  assign n33763 = pi787 & ~n33514;
  assign n33764 = ~n33762 & ~n33763;
  assign n33765 = pi644 & n33764;
  assign n33766 = ~pi715 & ~n33765;
  assign n33767 = ~n33761 & n33766;
  assign n33768 = ~n17652 & n33364;
  assign n33769 = n17652 & n33202;
  assign n33770 = ~n33768 & ~n33769;
  assign n33771 = ~pi644 & ~n33770;
  assign n33772 = pi644 & n33202;
  assign n33773 = pi715 & ~n33772;
  assign n33774 = ~n33771 & n33773;
  assign n33775 = ~pi1160 & ~n33774;
  assign n33776 = ~n33767 & n33775;
  assign n33777 = pi644 & n33759;
  assign n33778 = ~pi644 & n33764;
  assign n33779 = pi715 & ~n33778;
  assign n33780 = ~n33777 & n33779;
  assign n33781 = pi644 & ~n33770;
  assign n33782 = ~pi644 & n33202;
  assign n33783 = ~pi715 & ~n33782;
  assign n33784 = ~n33781 & n33783;
  assign n33785 = pi1160 & ~n33784;
  assign n33786 = ~n33780 & n33785;
  assign n33787 = pi790 & ~n33786;
  assign n33788 = ~n33776 & n33787;
  assign n33789 = ~n33760 & ~n33788;
  assign n33790 = ~po1038 & ~n33789;
  assign n33791 = pi198 & po1038;
  assign po355 = n33790 | n33791;
  assign n33793 = pi199 & ~n17406;
  assign n33794 = ~pi617 & ~n33793;
  assign n33795 = ~pi199 & ~n19216;
  assign n33796 = n19222 & ~n33795;
  assign n33797 = pi199 & n17242;
  assign n33798 = ~pi199 & ~n17275;
  assign n33799 = ~pi38 & ~n33798;
  assign n33800 = ~n33797 & n33799;
  assign n33801 = ~n33796 & ~n33800;
  assign n33802 = n3267 & ~n33801;
  assign n33803 = pi199 & ~n3267;
  assign n33804 = pi617 & ~n33803;
  assign n33805 = ~n33802 & n33804;
  assign n33806 = ~n33794 & ~n33805;
  assign n33807 = ~pi637 & n33806;
  assign n33808 = pi199 & n19235;
  assign n33809 = n3267 & ~n24373;
  assign n33810 = ~pi199 & ~n33809;
  assign n33811 = ~pi617 & ~n19231;
  assign n33812 = ~n33810 & n33811;
  assign n33813 = ~n33808 & n33812;
  assign n33814 = n3267 & n19253;
  assign n33815 = ~pi199 & ~n33814;
  assign n33816 = pi199 & n19261;
  assign n33817 = pi617 & ~n33816;
  assign n33818 = ~n33815 & n33817;
  assign n33819 = ~n33803 & ~n33818;
  assign n33820 = ~n33813 & n33819;
  assign n33821 = pi637 & ~n33820;
  assign n33822 = ~n33807 & ~n33821;
  assign n33823 = ~pi625 & n33822;
  assign n33824 = pi625 & ~n33806;
  assign n33825 = ~pi1153 & ~n33824;
  assign n33826 = ~n33823 & n33825;
  assign n33827 = ~pi637 & ~n33793;
  assign n33828 = ~pi199 & ~n17280;
  assign n33829 = n19802 & ~n33828;
  assign n33830 = pi199 & ~n17381;
  assign n33831 = ~pi199 & ~n17332;
  assign n33832 = pi39 & ~n33831;
  assign n33833 = ~n33830 & n33832;
  assign n33834 = ~pi199 & n17057;
  assign n33835 = pi199 & ~n17078;
  assign n33836 = ~pi39 & ~n33835;
  assign n33837 = ~n33834 & n33836;
  assign n33838 = ~pi38 & ~n33837;
  assign n33839 = ~n33833 & n33838;
  assign n33840 = ~n33829 & ~n33839;
  assign n33841 = n3267 & ~n33840;
  assign n33842 = pi637 & ~n33803;
  assign n33843 = ~n33841 & n33842;
  assign n33844 = ~n33827 & ~n33843;
  assign n33845 = pi625 & ~n33844;
  assign n33846 = ~pi625 & ~n33793;
  assign n33847 = pi1153 & ~n33846;
  assign n33848 = ~n33845 & n33847;
  assign n33849 = ~pi608 & ~n33848;
  assign n33850 = ~n33826 & n33849;
  assign n33851 = pi625 & n33822;
  assign n33852 = ~pi625 & ~n33806;
  assign n33853 = pi1153 & ~n33852;
  assign n33854 = ~n33851 & n33853;
  assign n33855 = ~pi625 & ~n33844;
  assign n33856 = pi625 & ~n33793;
  assign n33857 = ~pi1153 & ~n33856;
  assign n33858 = ~n33855 & n33857;
  assign n33859 = pi608 & ~n33858;
  assign n33860 = ~n33854 & n33859;
  assign n33861 = ~n33850 & ~n33860;
  assign n33862 = pi778 & ~n33861;
  assign n33863 = ~pi778 & n33822;
  assign n33864 = ~n33862 & ~n33863;
  assign n33865 = ~pi609 & ~n33864;
  assign n33866 = ~pi778 & n33844;
  assign n33867 = ~n33848 & ~n33858;
  assign n33868 = pi778 & ~n33867;
  assign n33869 = ~n33866 & ~n33868;
  assign n33870 = pi609 & n33869;
  assign n33871 = ~pi1155 & ~n33870;
  assign n33872 = ~n33865 & n33871;
  assign n33873 = ~n17438 & ~n33806;
  assign n33874 = n17438 & ~n33793;
  assign n33875 = ~n33873 & ~n33874;
  assign n33876 = pi609 & ~n33875;
  assign n33877 = ~pi609 & ~n33793;
  assign n33878 = pi1155 & ~n33877;
  assign n33879 = ~n33876 & n33878;
  assign n33880 = ~pi660 & ~n33879;
  assign n33881 = ~n33872 & n33880;
  assign n33882 = pi609 & ~n33864;
  assign n33883 = ~pi609 & n33869;
  assign n33884 = pi1155 & ~n33883;
  assign n33885 = ~n33882 & n33884;
  assign n33886 = ~pi609 & ~n33875;
  assign n33887 = pi609 & ~n33793;
  assign n33888 = ~pi1155 & ~n33887;
  assign n33889 = ~n33886 & n33888;
  assign n33890 = pi660 & ~n33889;
  assign n33891 = ~n33885 & n33890;
  assign n33892 = ~n33881 & ~n33891;
  assign n33893 = pi785 & ~n33892;
  assign n33894 = ~pi785 & ~n33864;
  assign n33895 = ~n33893 & ~n33894;
  assign n33896 = ~pi618 & ~n33895;
  assign n33897 = n17466 & ~n33793;
  assign n33898 = ~n17466 & n33869;
  assign n33899 = ~n33897 & ~n33898;
  assign n33900 = pi618 & ~n33899;
  assign n33901 = ~pi1154 & ~n33900;
  assign n33902 = ~n33896 & n33901;
  assign n33903 = ~pi785 & n33875;
  assign n33904 = ~n33879 & ~n33889;
  assign n33905 = pi785 & ~n33904;
  assign n33906 = ~n33903 & ~n33905;
  assign n33907 = pi618 & n33906;
  assign n33908 = ~pi618 & ~n33793;
  assign n33909 = pi1154 & ~n33908;
  assign n33910 = ~n33907 & n33909;
  assign n33911 = ~pi627 & ~n33910;
  assign n33912 = ~n33902 & n33911;
  assign n33913 = pi618 & ~n33895;
  assign n33914 = ~pi618 & ~n33899;
  assign n33915 = pi1154 & ~n33914;
  assign n33916 = ~n33913 & n33915;
  assign n33917 = ~pi618 & n33906;
  assign n33918 = pi618 & ~n33793;
  assign n33919 = ~pi1154 & ~n33918;
  assign n33920 = ~n33917 & n33919;
  assign n33921 = pi627 & ~n33920;
  assign n33922 = ~n33916 & n33921;
  assign n33923 = ~n33912 & ~n33922;
  assign n33924 = pi781 & ~n33923;
  assign n33925 = ~pi781 & ~n33895;
  assign n33926 = ~n33924 & ~n33925;
  assign n33927 = ~pi619 & ~n33926;
  assign n33928 = ~n17503 & n33899;
  assign n33929 = n17503 & n33793;
  assign n33930 = ~n33928 & ~n33929;
  assign n33931 = pi619 & n33930;
  assign n33932 = ~pi1159 & ~n33931;
  assign n33933 = ~n33927 & n33932;
  assign n33934 = ~pi781 & ~n33906;
  assign n33935 = ~n33910 & ~n33920;
  assign n33936 = pi781 & ~n33935;
  assign n33937 = ~n33934 & ~n33936;
  assign n33938 = pi619 & n33937;
  assign n33939 = ~pi619 & ~n33793;
  assign n33940 = pi1159 & ~n33939;
  assign n33941 = ~n33938 & n33940;
  assign n33942 = ~pi648 & ~n33941;
  assign n33943 = ~n33933 & n33942;
  assign n33944 = pi619 & ~n33926;
  assign n33945 = ~pi619 & n33930;
  assign n33946 = pi1159 & ~n33945;
  assign n33947 = ~n33944 & n33946;
  assign n33948 = ~pi619 & n33937;
  assign n33949 = pi619 & ~n33793;
  assign n33950 = ~pi1159 & ~n33949;
  assign n33951 = ~n33948 & n33950;
  assign n33952 = pi648 & ~n33951;
  assign n33953 = ~n33947 & n33952;
  assign n33954 = ~n33943 & ~n33953;
  assign n33955 = pi789 & ~n33954;
  assign n33956 = ~pi789 & ~n33926;
  assign n33957 = ~n33955 & ~n33956;
  assign n33958 = ~pi788 & n33957;
  assign n33959 = ~pi626 & n33957;
  assign n33960 = n17539 & ~n33793;
  assign n33961 = ~n17539 & n33930;
  assign n33962 = ~n33960 & ~n33961;
  assign n33963 = pi626 & n33962;
  assign n33964 = ~pi641 & ~n33963;
  assign n33965 = ~n33959 & n33964;
  assign n33966 = ~pi789 & ~n33937;
  assign n33967 = ~n33941 & ~n33951;
  assign n33968 = pi789 & ~n33967;
  assign n33969 = ~n33966 & ~n33968;
  assign n33970 = ~pi626 & ~n33969;
  assign n33971 = pi626 & n33793;
  assign n33972 = pi641 & ~n33971;
  assign n33973 = ~n33970 & n33972;
  assign n33974 = ~pi1158 & ~n33973;
  assign n33975 = ~n33965 & n33974;
  assign n33976 = pi626 & n33957;
  assign n33977 = ~pi626 & n33962;
  assign n33978 = pi641 & ~n33977;
  assign n33979 = ~n33976 & n33978;
  assign n33980 = pi626 & ~n33969;
  assign n33981 = ~pi626 & n33793;
  assign n33982 = ~pi641 & ~n33981;
  assign n33983 = ~n33980 & n33982;
  assign n33984 = pi1158 & ~n33983;
  assign n33985 = ~n33979 & n33984;
  assign n33986 = ~n33975 & ~n33985;
  assign n33987 = pi788 & ~n33986;
  assign n33988 = ~n33958 & ~n33987;
  assign n33989 = ~pi628 & n33988;
  assign n33990 = ~n17816 & ~n33969;
  assign n33991 = n17816 & n33793;
  assign n33992 = ~n33990 & ~n33991;
  assign n33993 = pi628 & n33992;
  assign n33994 = ~pi1156 & ~n33993;
  assign n33995 = ~n33989 & n33994;
  assign n33996 = ~n17582 & n33962;
  assign n33997 = n17582 & n33793;
  assign n33998 = ~n33996 & ~n33997;
  assign n33999 = pi628 & n33998;
  assign n34000 = ~pi628 & ~n33793;
  assign n34001 = pi1156 & ~n34000;
  assign n34002 = ~n33999 & n34001;
  assign n34003 = ~pi629 & ~n34002;
  assign n34004 = ~n33995 & n34003;
  assign n34005 = pi628 & n33988;
  assign n34006 = ~pi628 & n33992;
  assign n34007 = pi1156 & ~n34006;
  assign n34008 = ~n34005 & n34007;
  assign n34009 = ~pi628 & n33998;
  assign n34010 = pi628 & ~n33793;
  assign n34011 = ~pi1156 & ~n34010;
  assign n34012 = ~n34009 & n34011;
  assign n34013 = pi629 & ~n34012;
  assign n34014 = ~n34008 & n34013;
  assign n34015 = ~n34004 & ~n34014;
  assign n34016 = pi792 & ~n34015;
  assign n34017 = ~pi792 & n33988;
  assign n34018 = ~n34016 & ~n34017;
  assign n34019 = ~pi647 & ~n34018;
  assign n34020 = ~n17610 & ~n33992;
  assign n34021 = n17610 & n33793;
  assign n34022 = ~n34020 & ~n34021;
  assign n34023 = pi647 & n34022;
  assign n34024 = ~pi1157 & ~n34023;
  assign n34025 = ~n34019 & n34024;
  assign n34026 = ~pi792 & ~n33998;
  assign n34027 = ~n34002 & ~n34012;
  assign n34028 = pi792 & ~n34027;
  assign n34029 = ~n34026 & ~n34028;
  assign n34030 = pi647 & n34029;
  assign n34031 = ~pi647 & ~n33793;
  assign n34032 = pi1157 & ~n34031;
  assign n34033 = ~n34030 & n34032;
  assign n34034 = ~pi630 & ~n34033;
  assign n34035 = ~n34025 & n34034;
  assign n34036 = pi647 & ~n34018;
  assign n34037 = ~pi647 & n34022;
  assign n34038 = pi1157 & ~n34037;
  assign n34039 = ~n34036 & n34038;
  assign n34040 = ~pi647 & n34029;
  assign n34041 = pi647 & ~n33793;
  assign n34042 = ~pi1157 & ~n34041;
  assign n34043 = ~n34040 & n34042;
  assign n34044 = pi630 & ~n34043;
  assign n34045 = ~n34039 & n34044;
  assign n34046 = ~n34035 & ~n34045;
  assign n34047 = pi787 & ~n34046;
  assign n34048 = ~pi787 & ~n34018;
  assign n34049 = ~n34047 & ~n34048;
  assign n34050 = ~pi790 & n34049;
  assign n34051 = ~pi644 & ~n34049;
  assign n34052 = ~pi787 & ~n34029;
  assign n34053 = ~n34033 & ~n34043;
  assign n34054 = pi787 & ~n34053;
  assign n34055 = ~n34052 & ~n34054;
  assign n34056 = pi644 & n34055;
  assign n34057 = ~pi715 & ~n34056;
  assign n34058 = ~n34051 & n34057;
  assign n34059 = n17652 & ~n33793;
  assign n34060 = ~n17652 & n34022;
  assign n34061 = ~n34059 & ~n34060;
  assign n34062 = ~pi644 & ~n34061;
  assign n34063 = pi644 & ~n33793;
  assign n34064 = pi715 & ~n34063;
  assign n34065 = ~n34062 & n34064;
  assign n34066 = ~pi1160 & ~n34065;
  assign n34067 = ~n34058 & n34066;
  assign n34068 = pi644 & ~n34049;
  assign n34069 = ~pi644 & n34055;
  assign n34070 = pi715 & ~n34069;
  assign n34071 = ~n34068 & n34070;
  assign n34072 = pi644 & ~n34061;
  assign n34073 = ~pi644 & ~n33793;
  assign n34074 = ~pi715 & ~n34073;
  assign n34075 = ~n34072 & n34074;
  assign n34076 = pi1160 & ~n34075;
  assign n34077 = ~n34071 & n34076;
  assign n34078 = pi790 & ~n34077;
  assign n34079 = ~n34067 & n34078;
  assign n34080 = ~n34050 & ~n34079;
  assign n34081 = ~po1038 & ~n34080;
  assign n34082 = pi199 & po1038;
  assign po356 = n34081 | n34082;
  assign n34084 = pi200 & ~n17406;
  assign n34085 = ~pi606 & ~n34084;
  assign n34086 = ~pi200 & ~n19216;
  assign n34087 = n19222 & ~n34086;
  assign n34088 = pi200 & n17242;
  assign n34089 = ~pi200 & ~n17275;
  assign n34090 = ~pi38 & ~n34089;
  assign n34091 = ~n34088 & n34090;
  assign n34092 = ~n34087 & ~n34091;
  assign n34093 = n3267 & ~n34092;
  assign n34094 = pi200 & ~n3267;
  assign n34095 = pi606 & ~n34094;
  assign n34096 = ~n34093 & n34095;
  assign n34097 = ~n34085 & ~n34096;
  assign n34098 = ~n17438 & ~n34097;
  assign n34099 = n17438 & ~n34084;
  assign n34100 = ~n34098 & ~n34099;
  assign n34101 = ~pi785 & n34100;
  assign n34102 = pi609 & ~n34100;
  assign n34103 = ~pi609 & ~n34084;
  assign n34104 = pi1155 & ~n34103;
  assign n34105 = ~n34102 & n34104;
  assign n34106 = ~pi609 & ~n34100;
  assign n34107 = pi609 & ~n34084;
  assign n34108 = ~pi1155 & ~n34107;
  assign n34109 = ~n34106 & n34108;
  assign n34110 = ~n34105 & ~n34109;
  assign n34111 = pi785 & ~n34110;
  assign n34112 = ~n34101 & ~n34111;
  assign n34113 = ~pi781 & ~n34112;
  assign n34114 = pi618 & n34112;
  assign n34115 = ~pi618 & ~n34084;
  assign n34116 = pi1154 & ~n34115;
  assign n34117 = ~n34114 & n34116;
  assign n34118 = ~pi618 & n34112;
  assign n34119 = pi618 & ~n34084;
  assign n34120 = ~pi1154 & ~n34119;
  assign n34121 = ~n34118 & n34120;
  assign n34122 = ~n34117 & ~n34121;
  assign n34123 = pi781 & ~n34122;
  assign n34124 = ~n34113 & ~n34123;
  assign n34125 = ~pi789 & ~n34124;
  assign n34126 = pi619 & n34124;
  assign n34127 = ~pi619 & ~n34084;
  assign n34128 = pi1159 & ~n34127;
  assign n34129 = ~n34126 & n34128;
  assign n34130 = ~pi619 & n34124;
  assign n34131 = pi619 & ~n34084;
  assign n34132 = ~pi1159 & ~n34131;
  assign n34133 = ~n34130 & n34132;
  assign n34134 = ~n34129 & ~n34133;
  assign n34135 = pi789 & ~n34134;
  assign n34136 = ~n34125 & ~n34135;
  assign n34137 = ~n17816 & ~n34136;
  assign n34138 = n17816 & n34084;
  assign n34139 = ~n34137 & ~n34138;
  assign n34140 = ~n20409 & ~n34139;
  assign n34141 = n17539 & ~n34084;
  assign n34142 = n17466 & ~n34084;
  assign n34143 = ~pi643 & ~n34084;
  assign n34144 = ~pi200 & ~n17280;
  assign n34145 = n19802 & ~n34144;
  assign n34146 = pi200 & n17365;
  assign n34147 = ~pi200 & n17317;
  assign n34148 = ~pi299 & ~n34147;
  assign n34149 = ~n34146 & n34148;
  assign n34150 = pi200 & n17379;
  assign n34151 = ~pi200 & n17330;
  assign n34152 = pi299 & ~n34151;
  assign n34153 = ~n34150 & n34152;
  assign n34154 = ~n34149 & ~n34153;
  assign n34155 = pi39 & ~n34154;
  assign n34156 = pi200 & n17078;
  assign n34157 = ~pi200 & ~n17057;
  assign n34158 = ~pi39 & ~n34157;
  assign n34159 = ~n34156 & n34158;
  assign n34160 = ~n34155 & ~n34159;
  assign n34161 = ~pi38 & ~n34160;
  assign n34162 = ~n34145 & ~n34161;
  assign n34163 = n3267 & ~n34162;
  assign n34164 = pi643 & ~n34094;
  assign n34165 = ~n34163 & n34164;
  assign n34166 = ~n34143 & ~n34165;
  assign n34167 = ~pi778 & n34166;
  assign n34168 = pi625 & ~n34166;
  assign n34169 = ~pi625 & ~n34084;
  assign n34170 = pi1153 & ~n34169;
  assign n34171 = ~n34168 & n34170;
  assign n34172 = ~pi625 & ~n34166;
  assign n34173 = pi625 & ~n34084;
  assign n34174 = ~pi1153 & ~n34173;
  assign n34175 = ~n34172 & n34174;
  assign n34176 = ~n34171 & ~n34175;
  assign n34177 = pi778 & ~n34176;
  assign n34178 = ~n34167 & ~n34177;
  assign n34179 = ~n17466 & n34178;
  assign n34180 = ~n34142 & ~n34179;
  assign n34181 = ~n17503 & n34180;
  assign n34182 = n17503 & n34084;
  assign n34183 = ~n34181 & ~n34182;
  assign n34184 = ~n17539 & n34183;
  assign n34185 = ~n34141 & ~n34184;
  assign n34186 = ~n17582 & n34185;
  assign n34187 = n17582 & n34084;
  assign n34188 = ~n34186 & ~n34187;
  assign n34189 = pi628 & n34188;
  assign n34190 = ~pi628 & ~n34084;
  assign n34191 = pi1156 & ~n34190;
  assign n34192 = ~n34189 & n34191;
  assign n34193 = ~pi629 & n34192;
  assign n34194 = ~pi628 & n34188;
  assign n34195 = pi628 & ~n34084;
  assign n34196 = ~pi1156 & ~n34195;
  assign n34197 = ~n34194 & n34196;
  assign n34198 = pi629 & n34197;
  assign n34199 = ~n34193 & ~n34198;
  assign n34200 = ~n34140 & n34199;
  assign n34201 = pi792 & ~n34200;
  assign n34202 = ~pi643 & n34097;
  assign n34203 = pi200 & ~n19234;
  assign n34204 = ~pi200 & ~n19240;
  assign n34205 = ~pi38 & ~n34204;
  assign n34206 = ~n34203 & n34205;
  assign n34207 = ~n19230 & n34145;
  assign n34208 = ~n34206 & ~n34207;
  assign n34209 = ~pi606 & n3267;
  assign n34210 = ~n34208 & n34209;
  assign n34211 = pi200 & ~n24482;
  assign n34212 = ~pi200 & ~n19250;
  assign n34213 = ~pi38 & ~n34212;
  assign n34214 = ~n34211 & n34213;
  assign n34215 = ~n19248 & ~n19249;
  assign n34216 = ~pi200 & ~n34215;
  assign n34217 = pi38 & pi200;
  assign n34218 = n19258 & n34217;
  assign n34219 = pi606 & n3267;
  assign n34220 = ~n34218 & n34219;
  assign n34221 = ~n34216 & n34220;
  assign n34222 = ~n34214 & n34221;
  assign n34223 = ~n34094 & ~n34222;
  assign n34224 = ~n34210 & n34223;
  assign n34225 = pi643 & ~n34224;
  assign n34226 = ~n34202 & ~n34225;
  assign n34227 = ~pi625 & n34226;
  assign n34228 = pi625 & ~n34097;
  assign n34229 = ~pi1153 & ~n34228;
  assign n34230 = ~n34227 & n34229;
  assign n34231 = ~pi608 & ~n34171;
  assign n34232 = ~n34230 & n34231;
  assign n34233 = pi625 & n34226;
  assign n34234 = ~pi625 & ~n34097;
  assign n34235 = pi1153 & ~n34234;
  assign n34236 = ~n34233 & n34235;
  assign n34237 = pi608 & ~n34175;
  assign n34238 = ~n34236 & n34237;
  assign n34239 = ~n34232 & ~n34238;
  assign n34240 = pi778 & ~n34239;
  assign n34241 = ~pi778 & n34226;
  assign n34242 = ~n34240 & ~n34241;
  assign n34243 = ~pi609 & ~n34242;
  assign n34244 = pi609 & n34178;
  assign n34245 = ~pi1155 & ~n34244;
  assign n34246 = ~n34243 & n34245;
  assign n34247 = ~pi660 & ~n34105;
  assign n34248 = ~n34246 & n34247;
  assign n34249 = pi609 & ~n34242;
  assign n34250 = ~pi609 & n34178;
  assign n34251 = pi1155 & ~n34250;
  assign n34252 = ~n34249 & n34251;
  assign n34253 = pi660 & ~n34109;
  assign n34254 = ~n34252 & n34253;
  assign n34255 = ~n34248 & ~n34254;
  assign n34256 = pi785 & ~n34255;
  assign n34257 = ~pi785 & ~n34242;
  assign n34258 = ~n34256 & ~n34257;
  assign n34259 = ~pi618 & ~n34258;
  assign n34260 = pi618 & ~n34180;
  assign n34261 = ~pi1154 & ~n34260;
  assign n34262 = ~n34259 & n34261;
  assign n34263 = ~pi627 & ~n34117;
  assign n34264 = ~n34262 & n34263;
  assign n34265 = pi618 & ~n34258;
  assign n34266 = ~pi618 & ~n34180;
  assign n34267 = pi1154 & ~n34266;
  assign n34268 = ~n34265 & n34267;
  assign n34269 = pi627 & ~n34121;
  assign n34270 = ~n34268 & n34269;
  assign n34271 = ~n34264 & ~n34270;
  assign n34272 = pi781 & ~n34271;
  assign n34273 = ~pi781 & ~n34258;
  assign n34274 = ~n34272 & ~n34273;
  assign n34275 = pi619 & ~n34274;
  assign n34276 = ~pi619 & n34183;
  assign n34277 = pi1159 & ~n34276;
  assign n34278 = ~n34275 & n34277;
  assign n34279 = pi648 & ~n34133;
  assign n34280 = ~n34278 & n34279;
  assign n34281 = ~pi619 & ~n34274;
  assign n34282 = pi619 & n34183;
  assign n34283 = ~pi1159 & ~n34282;
  assign n34284 = ~n34281 & n34283;
  assign n34285 = ~pi648 & ~n34129;
  assign n34286 = ~n34284 & n34285;
  assign n34287 = pi789 & ~n34286;
  assign n34288 = ~n34280 & n34287;
  assign n34289 = ~pi789 & n34274;
  assign n34290 = n17817 & ~n34289;
  assign n34291 = ~n34288 & n34290;
  assign n34292 = pi626 & ~n34136;
  assign n34293 = ~pi626 & n34084;
  assign n34294 = n17579 & ~n34293;
  assign n34295 = ~n34292 & n34294;
  assign n34296 = n17704 & ~n34185;
  assign n34297 = ~pi626 & ~n34136;
  assign n34298 = pi626 & n34084;
  assign n34299 = n17580 & ~n34298;
  assign n34300 = ~n34297 & n34299;
  assign n34301 = ~n34296 & ~n34300;
  assign n34302 = ~n34295 & n34301;
  assign n34303 = pi788 & ~n34302;
  assign n34304 = ~n20205 & ~n34303;
  assign n34305 = ~n34291 & n34304;
  assign n34306 = ~n34201 & ~n34305;
  assign n34307 = n20207 & ~n34306;
  assign n34308 = ~pi792 & ~n34188;
  assign n34309 = ~n34192 & ~n34197;
  assign n34310 = pi792 & ~n34309;
  assign n34311 = ~n34308 & ~n34310;
  assign n34312 = pi647 & ~n34311;
  assign n34313 = ~pi647 & n34084;
  assign n34314 = ~n34312 & ~n34313;
  assign n34315 = n17649 & ~n34314;
  assign n34316 = ~pi647 & n34311;
  assign n34317 = pi647 & ~n34084;
  assign n34318 = ~pi1157 & ~n34317;
  assign n34319 = ~n34316 & n34318;
  assign n34320 = pi630 & n34319;
  assign n34321 = ~n17610 & ~n34139;
  assign n34322 = n17610 & n34084;
  assign n34323 = ~n34321 & ~n34322;
  assign n34324 = ~n20398 & ~n34323;
  assign n34325 = ~n34320 & ~n34324;
  assign n34326 = ~n34315 & n34325;
  assign n34327 = pi787 & ~n34326;
  assign n34328 = ~n34307 & ~n34327;
  assign n34329 = ~pi644 & n34328;
  assign n34330 = ~pi787 & ~n34311;
  assign n34331 = pi1157 & ~n34314;
  assign n34332 = ~n34319 & ~n34331;
  assign n34333 = pi787 & ~n34332;
  assign n34334 = ~n34330 & ~n34333;
  assign n34335 = pi644 & n34334;
  assign n34336 = ~pi715 & ~n34335;
  assign n34337 = ~n34329 & n34336;
  assign n34338 = ~n17652 & ~n34323;
  assign n34339 = n17652 & n34084;
  assign n34340 = ~n34338 & ~n34339;
  assign n34341 = ~pi644 & n34340;
  assign n34342 = pi644 & ~n34084;
  assign n34343 = pi715 & ~n34342;
  assign n34344 = ~n34341 & n34343;
  assign n34345 = ~pi1160 & ~n34344;
  assign n34346 = ~n34337 & n34345;
  assign n34347 = pi644 & n34328;
  assign n34348 = ~pi644 & n34334;
  assign n34349 = pi715 & ~n34348;
  assign n34350 = ~n34347 & n34349;
  assign n34351 = pi644 & n34340;
  assign n34352 = ~pi644 & ~n34084;
  assign n34353 = ~pi715 & ~n34352;
  assign n34354 = ~n34351 & n34353;
  assign n34355 = pi1160 & ~n34354;
  assign n34356 = ~n34350 & n34355;
  assign n34357 = ~n34346 & ~n34356;
  assign n34358 = pi790 & ~n34357;
  assign n34359 = ~pi790 & n34328;
  assign n34360 = ~n34358 & ~n34359;
  assign n34361 = ~po1038 & ~n34360;
  assign n34362 = ~pi200 & po1038;
  assign po357 = ~n34361 & ~n34362;
  assign n34364 = pi233 & pi237;
  assign n34365 = pi57 & pi332;
  assign n34366 = pi332 & ~n3293;
  assign n34367 = ~pi59 & ~n34366;
  assign n34368 = pi74 & pi332;
  assign n34369 = ~pi55 & ~n34368;
  assign n34370 = n2516 & n11026;
  assign n34371 = pi468 & n6157;
  assign n34372 = ~pi299 & pi587;
  assign n34373 = ~n20918 & ~n34372;
  assign n34374 = ~pi468 & ~n34373;
  assign n34375 = ~n34371 & ~n34374;
  assign n34376 = n34370 & ~n34375;
  assign n34377 = ~pi332 & ~n34376;
  assign n34378 = n7357 & ~n34377;
  assign n34379 = n3095 & n6599;
  assign n34380 = ~pi332 & ~n34379;
  assign n34381 = n15580 & ~n34380;
  assign n34382 = pi332 & ~n3238;
  assign n34383 = ~n34381 & ~n34382;
  assign n34384 = ~n34378 & n34383;
  assign n34385 = ~pi74 & ~n34384;
  assign n34386 = n34369 & ~n34385;
  assign n34387 = n3268 & n6555;
  assign n34388 = n3095 & n34387;
  assign n34389 = ~pi332 & ~n34388;
  assign n34390 = pi55 & n34389;
  assign n34391 = n3293 & ~n34390;
  assign n34392 = ~n34386 & n34391;
  assign n34393 = n34367 & ~n34392;
  assign n34394 = n6285 & ~n34389;
  assign n34395 = pi332 & ~n6285;
  assign n34396 = pi59 & ~n34395;
  assign n34397 = ~n34394 & n34396;
  assign n34398 = ~pi57 & ~n34397;
  assign n34399 = ~n34393 & n34398;
  assign n34400 = ~n34365 & ~n34399;
  assign n34401 = ~n34364 & ~n34400;
  assign n34402 = ~pi332 & ~n6157;
  assign n34403 = ~pi947 & ~n34402;
  assign n34404 = pi96 & pi210;
  assign n34405 = pi332 & n34404;
  assign n34406 = ~pi70 & ~pi841;
  assign n34407 = pi32 & ~n34406;
  assign n34408 = ~pi32 & ~pi70;
  assign n34409 = ~n34407 & ~n34408;
  assign n34410 = ~pi210 & n34409;
  assign n34411 = ~pi32 & ~pi96;
  assign n34412 = pi70 & n34411;
  assign n34413 = ~pi332 & ~n34412;
  assign n34414 = ~n34410 & n34413;
  assign n34415 = ~n34405 & ~n34414;
  assign n34416 = ~n6162 & n34415;
  assign n34417 = n6157 & ~n34416;
  assign n34418 = n34403 & ~n34417;
  assign n34419 = pi332 & pi468;
  assign n34420 = ~pi468 & ~n34414;
  assign n34421 = ~n34419 & ~n34420;
  assign n34422 = ~n6157 & n34421;
  assign n34423 = n6157 & ~n34415;
  assign n34424 = pi947 & ~n34423;
  assign n34425 = ~n34422 & n34424;
  assign n34426 = ~n34418 & ~n34425;
  assign n34427 = pi57 & ~n34426;
  assign n34428 = ~n3268 & n34426;
  assign n34429 = ~pi95 & n2720;
  assign n34430 = ~pi70 & ~n34429;
  assign n34431 = n34411 & ~n34430;
  assign n34432 = pi210 & n34431;
  assign n34433 = ~pi95 & n2783;
  assign n34434 = ~n34407 & n34433;
  assign n34435 = n2495 & n34434;
  assign n34436 = n2523 & n34435;
  assign n34437 = ~n34409 & ~n34436;
  assign n34438 = ~pi210 & ~n34437;
  assign n34439 = ~pi332 & ~n34438;
  assign n34440 = ~n34432 & n34439;
  assign n34441 = ~n34405 & ~n34440;
  assign n34442 = ~n6162 & n34441;
  assign n34443 = n6157 & ~n34442;
  assign n34444 = n34403 & ~n34443;
  assign n34445 = ~pi468 & ~n34440;
  assign n34446 = ~n34419 & ~n34445;
  assign n34447 = ~n6157 & n34446;
  assign n34448 = n6157 & ~n34441;
  assign n34449 = pi947 & ~n34448;
  assign n34450 = ~n34447 & n34449;
  assign n34451 = ~n34444 & ~n34450;
  assign n34452 = n3268 & n34451;
  assign n34453 = ~n34428 & ~n34452;
  assign n34454 = n6285 & ~n34453;
  assign n34455 = ~n6285 & n34426;
  assign n34456 = pi59 & ~n34455;
  assign n34457 = ~n34454 & n34456;
  assign n34458 = n2516 & n2535;
  assign n34459 = ~pi95 & n2450;
  assign n34460 = n34458 & n34459;
  assign n34461 = ~pi70 & ~n34460;
  assign n34462 = n34411 & ~n34461;
  assign n34463 = pi210 & n34462;
  assign n34464 = n34434 & n34458;
  assign n34465 = ~n34409 & ~n34464;
  assign n34466 = ~pi210 & ~n34465;
  assign n34467 = ~pi332 & ~n34466;
  assign n34468 = ~n34463 & n34467;
  assign n34469 = ~pi468 & ~n34468;
  assign n34470 = ~n34419 & ~n34469;
  assign n34471 = ~n6157 & n34470;
  assign n34472 = ~n34405 & ~n34468;
  assign n34473 = n6157 & ~n34472;
  assign n34474 = pi947 & ~n34473;
  assign n34475 = ~n34471 & n34474;
  assign n34476 = ~n6162 & n34472;
  assign n34477 = n6157 & ~n34476;
  assign n34478 = n34403 & ~n34477;
  assign n34479 = pi299 & ~n34478;
  assign n34480 = ~n34475 & n34479;
  assign n34481 = pi198 & n34462;
  assign n34482 = ~pi198 & ~n34465;
  assign n34483 = ~pi332 & ~n34482;
  assign n34484 = ~n34481 & n34483;
  assign n34485 = ~pi468 & ~n34484;
  assign n34486 = ~n6157 & ~n34419;
  assign n34487 = ~n34485 & n34486;
  assign n34488 = pi96 & pi198;
  assign n34489 = pi332 & n34488;
  assign n34490 = ~n34484 & ~n34489;
  assign n34491 = n6157 & ~n34490;
  assign n34492 = pi587 & ~n34491;
  assign n34493 = ~n34487 & n34492;
  assign n34494 = ~pi587 & ~n34402;
  assign n34495 = ~n6162 & n34490;
  assign n34496 = n6157 & ~n34495;
  assign n34497 = n34494 & ~n34496;
  assign n34498 = ~pi299 & ~n34497;
  assign n34499 = ~n34493 & n34498;
  assign n34500 = ~n34480 & ~n34499;
  assign n34501 = n7357 & ~n34500;
  assign n34502 = pi198 & n34431;
  assign n34503 = ~pi198 & ~n34437;
  assign n34504 = ~pi332 & ~n34503;
  assign n34505 = ~n34502 & n34504;
  assign n34506 = ~n34489 & ~n34505;
  assign n34507 = ~n6162 & n34506;
  assign n34508 = n6157 & ~n34507;
  assign n34509 = n34494 & ~n34508;
  assign n34510 = ~pi468 & ~n34505;
  assign n34511 = n34486 & ~n34510;
  assign n34512 = n6157 & ~n34506;
  assign n34513 = pi587 & ~n34512;
  assign n34514 = ~n34511 & n34513;
  assign n34515 = ~n34509 & ~n34514;
  assign n34516 = ~pi299 & ~n34515;
  assign n34517 = pi299 & ~n34451;
  assign n34518 = n15580 & ~n34517;
  assign n34519 = ~n34516 & n34518;
  assign n34520 = ~n34501 & ~n34519;
  assign n34521 = ~pi74 & ~n34520;
  assign n34522 = pi299 & ~n34426;
  assign n34523 = ~pi74 & n3238;
  assign n34524 = ~pi198 & n34409;
  assign n34525 = n34413 & ~n34524;
  assign n34526 = n6559 & ~n34525;
  assign n34527 = n34402 & ~n34526;
  assign n34528 = ~n34489 & ~n34525;
  assign n34529 = n6157 & ~n34528;
  assign n34530 = ~pi299 & ~n6558;
  assign n34531 = ~n34529 & n34530;
  assign n34532 = ~n34527 & n34531;
  assign n34533 = ~n34523 & ~n34532;
  assign n34534 = ~n34522 & n34533;
  assign n34535 = ~pi55 & ~n34534;
  assign n34536 = ~n34521 & n34535;
  assign n34537 = pi55 & n34453;
  assign n34538 = n3293 & ~n34537;
  assign n34539 = ~n34536 & n34538;
  assign n34540 = ~n3293 & n34426;
  assign n34541 = ~pi59 & ~n34540;
  assign n34542 = ~n34539 & n34541;
  assign n34543 = ~n34457 & ~n34542;
  assign n34544 = ~pi57 & ~n34543;
  assign n34545 = ~n34427 & ~n34544;
  assign n34546 = n34364 & ~n34545;
  assign n34547 = ~n34401 & ~n34546;
  assign n34548 = ~pi201 & ~n34547;
  assign n34549 = ~n6555 & ~n16361;
  assign n34550 = n6598 & ~po1038;
  assign n34551 = ~n34549 & ~n34550;
  assign n34552 = ~n16361 & ~n34404;
  assign n34553 = n16361 & ~n34488;
  assign n34554 = ~n34552 & ~n34553;
  assign n34555 = n34551 & n34554;
  assign n34556 = n34364 & n34555;
  assign n34557 = pi201 & ~n34556;
  assign po358 = ~n34548 & ~n34557;
  assign n34559 = ~pi233 & pi237;
  assign n34560 = ~n34400 & ~n34559;
  assign n34561 = ~n34545 & n34559;
  assign n34562 = ~n34560 & ~n34561;
  assign n34563 = ~pi202 & ~n34562;
  assign n34564 = n34555 & n34559;
  assign n34565 = pi202 & ~n34564;
  assign po359 = ~n34563 & ~n34565;
  assign n34567 = ~pi233 & ~pi237;
  assign n34568 = ~n34400 & ~n34567;
  assign n34569 = ~n34545 & n34567;
  assign n34570 = ~n34568 & ~n34569;
  assign n34571 = ~pi203 & ~n34570;
  assign n34572 = n34555 & n34567;
  assign n34573 = pi203 & ~n34572;
  assign po360 = ~n34571 & ~n34573;
  assign n34575 = ~pi468 & pi602;
  assign n34576 = pi468 & n6160;
  assign n34577 = ~n34575 & ~n34576;
  assign n34578 = ~pi299 & ~n34577;
  assign n34579 = ~n6473 & ~n34578;
  assign n34580 = n3095 & ~n34579;
  assign n34581 = ~pi332 & ~n34580;
  assign n34582 = n15580 & ~n34581;
  assign n34583 = pi299 & ~pi907;
  assign n34584 = ~pi299 & ~pi602;
  assign n34585 = ~pi468 & ~n34584;
  assign n34586 = ~n34583 & n34585;
  assign n34587 = ~n34576 & ~n34586;
  assign n34588 = n34370 & ~n34587;
  assign n34589 = ~pi332 & ~n34588;
  assign n34590 = n7357 & ~n34589;
  assign n34591 = ~n34582 & ~n34590;
  assign n34592 = ~pi74 & ~n34591;
  assign n34593 = n34369 & ~n34382;
  assign n34594 = ~n34592 & n34593;
  assign n34595 = n3268 & n6291;
  assign n34596 = n3095 & n34595;
  assign n34597 = ~pi332 & ~n34596;
  assign n34598 = pi55 & n34597;
  assign n34599 = n3293 & ~n34598;
  assign n34600 = ~n34594 & n34599;
  assign n34601 = n34367 & ~n34600;
  assign n34602 = n6285 & ~n34597;
  assign n34603 = n34396 & ~n34602;
  assign n34604 = ~pi57 & ~n34603;
  assign n34605 = ~n34601 & n34604;
  assign n34606 = ~n34365 & ~n34605;
  assign n34607 = ~n34364 & ~n34606;
  assign n34608 = ~pi332 & ~n6160;
  assign n34609 = ~pi907 & ~n34608;
  assign n34610 = n6160 & ~n34416;
  assign n34611 = n34609 & ~n34610;
  assign n34612 = ~n6160 & n34421;
  assign n34613 = n6160 & ~n34415;
  assign n34614 = pi907 & ~n34613;
  assign n34615 = ~n34612 & n34614;
  assign n34616 = ~n34611 & ~n34615;
  assign n34617 = pi57 & ~n34616;
  assign n34618 = ~n3268 & n34616;
  assign n34619 = ~n6160 & n34446;
  assign n34620 = n6160 & ~n34441;
  assign n34621 = pi907 & ~n34620;
  assign n34622 = ~n34619 & n34621;
  assign n34623 = pi332 & ~n16512;
  assign n34624 = pi680 & ~n34623;
  assign n34625 = ~n34442 & n34624;
  assign n34626 = n34609 & ~n34625;
  assign n34627 = ~n34622 & ~n34626;
  assign n34628 = n3268 & n34627;
  assign n34629 = ~n34618 & ~n34628;
  assign n34630 = n6285 & ~n34629;
  assign n34631 = ~n6285 & n34616;
  assign n34632 = pi59 & ~n34631;
  assign n34633 = ~n34630 & n34632;
  assign n34634 = pi299 & n34627;
  assign n34635 = n6160 & n34488;
  assign n34636 = pi332 & ~n34635;
  assign n34637 = ~pi299 & ~n34636;
  assign n34638 = n6299 & n34506;
  assign n34639 = n34637 & ~n34638;
  assign n34640 = ~n34634 & ~n34639;
  assign n34641 = n15580 & ~n34640;
  assign n34642 = n6299 & n34490;
  assign n34643 = n34637 & ~n34642;
  assign n34644 = ~n6160 & n34470;
  assign n34645 = n6160 & ~n34472;
  assign n34646 = pi907 & ~n34645;
  assign n34647 = ~n34644 & n34646;
  assign n34648 = n6160 & ~n34476;
  assign n34649 = n34609 & ~n34648;
  assign n34650 = pi299 & ~n34649;
  assign n34651 = ~n34647 & n34650;
  assign n34652 = ~n34643 & ~n34651;
  assign n34653 = n7357 & ~n34652;
  assign n34654 = ~n34641 & ~n34653;
  assign n34655 = ~pi74 & ~n34654;
  assign n34656 = pi299 & ~n34616;
  assign n34657 = n34528 & ~n34577;
  assign n34658 = ~n34636 & ~n34657;
  assign n34659 = ~pi299 & ~n34658;
  assign n34660 = ~n34523 & ~n34659;
  assign n34661 = ~n34656 & n34660;
  assign n34662 = ~pi55 & ~n34661;
  assign n34663 = ~n34655 & n34662;
  assign n34664 = pi55 & n34629;
  assign n34665 = n3293 & ~n34664;
  assign n34666 = ~n34663 & n34665;
  assign n34667 = ~n3293 & n34616;
  assign n34668 = ~pi59 & ~n34667;
  assign n34669 = ~n34666 & n34668;
  assign n34670 = ~n34633 & ~n34669;
  assign n34671 = ~pi57 & ~n34670;
  assign n34672 = ~n34617 & ~n34671;
  assign n34673 = n34364 & ~n34672;
  assign n34674 = ~n34607 & ~n34673;
  assign n34675 = ~pi204 & ~n34674;
  assign n34676 = ~n6291 & ~n16361;
  assign n34677 = ~n6299 & n16361;
  assign n34678 = ~n34676 & ~n34677;
  assign n34679 = n34554 & n34678;
  assign n34680 = n34364 & n34679;
  assign n34681 = pi204 & ~n34680;
  assign po361 = ~n34675 & ~n34681;
  assign n34683 = ~n34559 & ~n34606;
  assign n34684 = n34559 & ~n34672;
  assign n34685 = ~n34683 & ~n34684;
  assign n34686 = ~pi205 & ~n34685;
  assign n34687 = n34559 & n34679;
  assign n34688 = pi205 & ~n34687;
  assign po362 = ~n34686 & ~n34688;
  assign n34690 = pi233 & ~pi237;
  assign n34691 = ~n34606 & ~n34690;
  assign n34692 = ~n34672 & n34690;
  assign n34693 = ~n34691 & ~n34692;
  assign n34694 = ~pi206 & ~n34693;
  assign n34695 = n34679 & n34690;
  assign n34696 = pi206 & ~n34695;
  assign po363 = ~n34694 & ~n34696;
  assign n34698 = ~n19038 & n24209;
  assign n34699 = n19128 & n34698;
  assign n34700 = ~n19158 & n34699;
  assign n34701 = pi207 & ~n34700;
  assign n34702 = ~n17406 & n17539;
  assign n34703 = n3267 & n24212;
  assign n34704 = ~pi778 & ~n34703;
  assign n34705 = ~pi625 & ~n17406;
  assign n34706 = pi625 & ~n34703;
  assign n34707 = ~n34705 & ~n34706;
  assign n34708 = pi1153 & ~n34707;
  assign n34709 = pi625 & ~n17406;
  assign n34710 = ~pi625 & ~n34703;
  assign n34711 = ~n34709 & ~n34710;
  assign n34712 = ~pi1153 & ~n34711;
  assign n34713 = ~n34708 & ~n34712;
  assign n34714 = pi778 & ~n34713;
  assign n34715 = ~n34704 & ~n34714;
  assign n34716 = ~n17466 & ~n34715;
  assign n34717 = ~n17406 & n17466;
  assign n34718 = ~n34716 & ~n34717;
  assign n34719 = ~n17503 & n34718;
  assign n34720 = n17406 & n17503;
  assign n34721 = ~n34719 & ~n34720;
  assign n34722 = ~n17539 & n34721;
  assign n34723 = ~n34702 & ~n34722;
  assign n34724 = ~n17582 & n34723;
  assign n34725 = n17406 & n17582;
  assign n34726 = ~n34724 & ~n34725;
  assign n34727 = ~n19158 & ~n34726;
  assign n34728 = n17406 & n17858;
  assign n34729 = ~n34727 & ~n34728;
  assign n34730 = ~pi207 & ~n34729;
  assign n34731 = ~n34701 & ~n34730;
  assign n34732 = pi710 & ~n34731;
  assign n34733 = ~pi207 & ~n17406;
  assign n34734 = ~pi710 & ~n34733;
  assign n34735 = ~n34732 & ~n34734;
  assign n34736 = ~pi647 & n34735;
  assign n34737 = pi647 & n34733;
  assign n34738 = ~pi1157 & ~n34737;
  assign n34739 = ~n34736 & n34738;
  assign n34740 = pi630 & n34739;
  assign n34741 = pi647 & n34735;
  assign n34742 = ~pi647 & n34733;
  assign n34743 = pi1157 & ~n34742;
  assign n34744 = ~n34741 & n34743;
  assign n34745 = ~pi630 & n34744;
  assign n34746 = ~n17406 & n17438;
  assign n34747 = n3267 & n19223;
  assign n34748 = ~n17438 & ~n34747;
  assign n34749 = ~n34746 & ~n34748;
  assign n34750 = ~pi785 & ~n34749;
  assign n34751 = ~n17406 & ~n17451;
  assign n34752 = ~pi609 & n34748;
  assign n34753 = ~n34751 & ~n34752;
  assign n34754 = ~pi1155 & ~n34753;
  assign n34755 = ~n17406 & ~n17439;
  assign n34756 = pi609 & n34748;
  assign n34757 = ~n34755 & ~n34756;
  assign n34758 = pi1155 & ~n34757;
  assign n34759 = ~n34754 & ~n34758;
  assign n34760 = pi785 & ~n34759;
  assign n34761 = ~n34750 & ~n34760;
  assign n34762 = ~pi781 & ~n34761;
  assign n34763 = ~pi618 & n34761;
  assign n34764 = pi618 & n17406;
  assign n34765 = ~pi1154 & ~n34764;
  assign n34766 = ~n34763 & n34765;
  assign n34767 = pi618 & n34761;
  assign n34768 = ~pi618 & n17406;
  assign n34769 = pi1154 & ~n34768;
  assign n34770 = ~n34767 & n34769;
  assign n34771 = ~n34766 & ~n34770;
  assign n34772 = pi781 & ~n34771;
  assign n34773 = ~n34762 & ~n34772;
  assign n34774 = ~pi789 & ~n34773;
  assign n34775 = ~pi619 & n34773;
  assign n34776 = pi619 & n17406;
  assign n34777 = ~pi1159 & ~n34776;
  assign n34778 = ~n34775 & n34777;
  assign n34779 = pi619 & n34773;
  assign n34780 = ~pi619 & n17406;
  assign n34781 = pi1159 & ~n34780;
  assign n34782 = ~n34779 & n34781;
  assign n34783 = ~n34778 & ~n34782;
  assign n34784 = pi789 & ~n34783;
  assign n34785 = ~n34774 & ~n34784;
  assign n34786 = ~n17816 & n34785;
  assign n34787 = n17406 & n17816;
  assign n34788 = ~n34786 & ~n34787;
  assign n34789 = ~n17610 & ~n34788;
  assign n34790 = n17406 & n17610;
  assign n34791 = ~n34789 & ~n34790;
  assign n34792 = ~pi207 & ~n34791;
  assign n34793 = n3267 & ~n24271;
  assign n34794 = ~n17438 & n34793;
  assign n34795 = ~n20069 & n34794;
  assign n34796 = ~n20075 & n34795;
  assign n34797 = ~n20079 & n34796;
  assign n34798 = ~n17816 & n34797;
  assign n34799 = ~n17610 & n34798;
  assign n34800 = pi207 & ~n34799;
  assign n34801 = pi623 & ~n34800;
  assign n34802 = ~n34792 & n34801;
  assign n34803 = ~pi623 & n34733;
  assign n34804 = ~n34802 & ~n34803;
  assign n34805 = ~n20398 & n34804;
  assign n34806 = ~n34745 & ~n34805;
  assign n34807 = ~n34740 & n34806;
  assign n34808 = pi787 & ~n34807;
  assign n34809 = ~pi628 & ~n17406;
  assign n34810 = pi628 & n34726;
  assign n34811 = ~n34809 & ~n34810;
  assign n34812 = ~pi629 & ~n34811;
  assign n34813 = ~n34809 & ~n34812;
  assign n34814 = pi1156 & ~n34813;
  assign n34815 = pi628 & ~n17406;
  assign n34816 = ~pi1156 & n34815;
  assign n34817 = ~pi628 & n34726;
  assign n34818 = ~n34815 & ~n34817;
  assign n34819 = n17608 & ~n34818;
  assign n34820 = ~n34816 & ~n34819;
  assign n34821 = ~n34814 & n34820;
  assign n34822 = pi792 & ~n34821;
  assign n34823 = pi619 & n34721;
  assign n34824 = pi618 & ~n34718;
  assign n34825 = pi609 & ~n34715;
  assign n34826 = n3267 & ~n19236;
  assign n34827 = ~pi778 & ~n34826;
  assign n34828 = pi625 & ~n34826;
  assign n34829 = ~n34705 & ~n34828;
  assign n34830 = pi1153 & ~n34829;
  assign n34831 = pi608 & ~n34712;
  assign n34832 = ~n34830 & n34831;
  assign n34833 = ~pi625 & ~n34826;
  assign n34834 = ~n34709 & ~n34833;
  assign n34835 = ~pi1153 & ~n34834;
  assign n34836 = ~pi608 & ~n34708;
  assign n34837 = ~n34835 & n34836;
  assign n34838 = pi778 & ~n34837;
  assign n34839 = ~n34832 & n34838;
  assign n34840 = ~n34827 & ~n34839;
  assign n34841 = ~pi609 & ~n34840;
  assign n34842 = ~n34825 & ~n34841;
  assign n34843 = ~pi1155 & ~n34842;
  assign n34844 = pi1155 & ~n17406;
  assign n34845 = ~pi660 & ~n34844;
  assign n34846 = ~n34843 & n34845;
  assign n34847 = ~pi609 & ~n34715;
  assign n34848 = pi609 & ~n34840;
  assign n34849 = ~n34847 & ~n34848;
  assign n34850 = pi1155 & ~n34849;
  assign n34851 = ~pi1155 & ~n17406;
  assign n34852 = pi660 & ~n34851;
  assign n34853 = ~n34850 & n34852;
  assign n34854 = ~n34846 & ~n34853;
  assign n34855 = pi785 & ~n34854;
  assign n34856 = ~pi785 & n34840;
  assign n34857 = ~n34855 & ~n34856;
  assign n34858 = ~pi618 & n34857;
  assign n34859 = ~n34824 & ~n34858;
  assign n34860 = ~pi1154 & ~n34859;
  assign n34861 = pi1154 & ~n17406;
  assign n34862 = ~pi627 & ~n34861;
  assign n34863 = ~n34860 & n34862;
  assign n34864 = ~pi618 & ~n34718;
  assign n34865 = pi618 & n34857;
  assign n34866 = ~n34864 & ~n34865;
  assign n34867 = pi1154 & ~n34866;
  assign n34868 = ~pi1154 & ~n17406;
  assign n34869 = pi627 & ~n34868;
  assign n34870 = ~n34867 & n34869;
  assign n34871 = ~n34863 & ~n34870;
  assign n34872 = pi781 & ~n34871;
  assign n34873 = ~pi781 & ~n34857;
  assign n34874 = ~n34872 & ~n34873;
  assign n34875 = ~pi619 & n34874;
  assign n34876 = ~n34823 & ~n34875;
  assign n34877 = ~pi1159 & ~n34876;
  assign n34878 = pi1159 & ~n17406;
  assign n34879 = ~pi648 & ~n34878;
  assign n34880 = ~n34877 & n34879;
  assign n34881 = ~pi619 & n34721;
  assign n34882 = pi619 & n34874;
  assign n34883 = ~n34881 & ~n34882;
  assign n34884 = pi1159 & ~n34883;
  assign n34885 = ~pi1159 & ~n17406;
  assign n34886 = pi648 & ~n34885;
  assign n34887 = ~n34884 & n34886;
  assign n34888 = ~n34880 & ~n34887;
  assign n34889 = pi789 & ~n34888;
  assign n34890 = ~pi789 & ~n34874;
  assign n34891 = ~n34889 & ~n34890;
  assign n34892 = ~pi626 & ~n34891;
  assign n34893 = pi626 & n34723;
  assign n34894 = ~pi641 & ~n34893;
  assign n34895 = ~n34892 & n34894;
  assign n34896 = pi641 & ~n17406;
  assign n34897 = ~pi1158 & ~n34896;
  assign n34898 = ~n34895 & n34897;
  assign n34899 = pi626 & ~n34891;
  assign n34900 = ~pi626 & n34723;
  assign n34901 = pi641 & ~n34900;
  assign n34902 = ~n34899 & n34901;
  assign n34903 = ~pi641 & ~n17406;
  assign n34904 = pi1158 & ~n34903;
  assign n34905 = ~n34902 & n34904;
  assign n34906 = ~n34898 & ~n34905;
  assign n34907 = pi788 & ~n34906;
  assign n34908 = ~pi788 & ~n34891;
  assign n34909 = ~n20205 & ~n34908;
  assign n34910 = ~n34907 & n34909;
  assign n34911 = ~n34822 & ~n34910;
  assign n34912 = ~pi207 & ~n34911;
  assign n34913 = ~pi778 & ~n33809;
  assign n34914 = pi625 & n33809;
  assign n34915 = pi1153 & ~n34914;
  assign n34916 = ~pi625 & n24209;
  assign n34917 = ~pi1153 & ~n34916;
  assign n34918 = pi608 & ~n34917;
  assign n34919 = ~n34915 & n34918;
  assign n34920 = ~pi625 & n33809;
  assign n34921 = ~pi1153 & ~n34920;
  assign n34922 = pi625 & n24209;
  assign n34923 = pi1153 & ~n34922;
  assign n34924 = ~pi608 & ~n34923;
  assign n34925 = ~n34921 & n34924;
  assign n34926 = pi778 & ~n34925;
  assign n34927 = ~n34919 & n34926;
  assign n34928 = ~n34913 & ~n34927;
  assign n34929 = ~pi609 & ~n34928;
  assign n34930 = pi609 & ~n34698;
  assign n34931 = n17463 & ~n34930;
  assign n34932 = ~n34929 & n34931;
  assign n34933 = pi609 & ~n34928;
  assign n34934 = ~pi609 & ~n34698;
  assign n34935 = n17464 & ~n34934;
  assign n34936 = ~n34933 & n34935;
  assign n34937 = ~n34932 & ~n34936;
  assign n34938 = pi785 & ~n34937;
  assign n34939 = ~pi785 & n34928;
  assign n34940 = ~n34938 & ~n34939;
  assign n34941 = pi618 & n34940;
  assign n34942 = ~n17466 & n34698;
  assign n34943 = ~pi618 & ~n34942;
  assign n34944 = n17501 & ~n34943;
  assign n34945 = ~n34941 & n34944;
  assign n34946 = ~pi618 & n34940;
  assign n34947 = pi618 & ~n34942;
  assign n34948 = n17500 & ~n34947;
  assign n34949 = ~n34946 & n34948;
  assign n34950 = pi781 & ~n34949;
  assign n34951 = ~n34945 & n34950;
  assign n34952 = ~pi781 & n34940;
  assign n34953 = ~n23444 & ~n34952;
  assign n34954 = ~n34951 & n34953;
  assign n34955 = n19127 & n34698;
  assign n34956 = n17538 & n20079;
  assign n34957 = n34955 & n34956;
  assign n34958 = ~n34954 & ~n34957;
  assign n34959 = pi626 & n34958;
  assign n34960 = ~n17539 & n34955;
  assign n34961 = ~pi626 & ~n34960;
  assign n34962 = pi641 & ~n34961;
  assign n34963 = pi1158 & n34962;
  assign n34964 = ~n34959 & n34963;
  assign n34965 = ~pi626 & n34958;
  assign n34966 = pi626 & ~n34960;
  assign n34967 = ~pi641 & ~n34966;
  assign n34968 = ~pi1158 & n34967;
  assign n34969 = ~n34965 & n34968;
  assign n34970 = pi788 & ~n34969;
  assign n34971 = ~n34964 & n34970;
  assign n34972 = ~pi788 & n34958;
  assign n34973 = ~n20205 & ~n34972;
  assign n34974 = ~n34971 & n34973;
  assign n34975 = n17610 & n17857;
  assign n34976 = n34699 & n34975;
  assign n34977 = ~n34974 & ~n34976;
  assign n34978 = pi207 & ~n34977;
  assign n34979 = ~pi623 & ~n34978;
  assign n34980 = ~n34912 & n34979;
  assign n34981 = n3267 & n19261;
  assign n34982 = ~pi778 & ~n34981;
  assign n34983 = pi625 & n34747;
  assign n34984 = ~pi625 & n34981;
  assign n34985 = ~pi1153 & ~n34984;
  assign n34986 = ~n34983 & n34985;
  assign n34987 = n34836 & ~n34986;
  assign n34988 = ~pi625 & n34747;
  assign n34989 = pi625 & n34981;
  assign n34990 = pi1153 & ~n34989;
  assign n34991 = ~n34988 & n34990;
  assign n34992 = n34831 & ~n34991;
  assign n34993 = pi778 & ~n34992;
  assign n34994 = ~n34987 & n34993;
  assign n34995 = ~n34982 & ~n34994;
  assign n34996 = ~pi609 & ~n34995;
  assign n34997 = ~n34825 & ~n34996;
  assign n34998 = ~pi1155 & ~n34997;
  assign n34999 = ~pi660 & ~n34758;
  assign n35000 = ~n34998 & n34999;
  assign n35001 = pi609 & ~n34995;
  assign n35002 = ~n34847 & ~n35001;
  assign n35003 = pi1155 & ~n35002;
  assign n35004 = pi660 & ~n34754;
  assign n35005 = ~n35003 & n35004;
  assign n35006 = ~n35000 & ~n35005;
  assign n35007 = pi785 & ~n35006;
  assign n35008 = ~pi785 & n34995;
  assign n35009 = ~n35007 & ~n35008;
  assign n35010 = ~pi618 & n35009;
  assign n35011 = ~n34824 & ~n35010;
  assign n35012 = ~pi1154 & ~n35011;
  assign n35013 = ~pi627 & ~n34770;
  assign n35014 = ~n35012 & n35013;
  assign n35015 = pi618 & n35009;
  assign n35016 = ~n34864 & ~n35015;
  assign n35017 = pi1154 & ~n35016;
  assign n35018 = pi627 & ~n34766;
  assign n35019 = ~n35017 & n35018;
  assign n35020 = ~n35014 & ~n35019;
  assign n35021 = pi781 & ~n35020;
  assign n35022 = ~pi781 & ~n35009;
  assign n35023 = ~n35021 & ~n35022;
  assign n35024 = pi619 & n35023;
  assign n35025 = ~n34881 & ~n35024;
  assign n35026 = pi1159 & ~n35025;
  assign n35027 = pi648 & ~n34778;
  assign n35028 = ~n35026 & n35027;
  assign n35029 = ~pi619 & n35023;
  assign n35030 = ~n34823 & ~n35029;
  assign n35031 = ~pi1159 & ~n35030;
  assign n35032 = ~pi648 & ~n34782;
  assign n35033 = ~n35031 & n35032;
  assign n35034 = pi789 & ~n35033;
  assign n35035 = ~n35028 & n35034;
  assign n35036 = ~pi789 & n35023;
  assign n35037 = n17817 & ~n35036;
  assign n35038 = ~n35035 & n35037;
  assign n35039 = ~n17581 & ~n17703;
  assign n35040 = n34785 & n35039;
  assign n35041 = pi641 & ~n34723;
  assign n35042 = n17698 & ~n34903;
  assign n35043 = ~n35041 & n35042;
  assign n35044 = ~pi641 & ~n34723;
  assign n35045 = n17699 & ~n34896;
  assign n35046 = ~n35044 & n35045;
  assign n35047 = ~n35043 & ~n35046;
  assign n35048 = ~n35040 & n35047;
  assign n35049 = pi788 & ~n35048;
  assign n35050 = ~n20205 & ~n35049;
  assign n35051 = ~n35038 & n35050;
  assign n35052 = pi1156 & n34812;
  assign n35053 = ~n20409 & n34788;
  assign n35054 = ~n34819 & ~n35053;
  assign n35055 = ~n35052 & n35054;
  assign n35056 = pi792 & ~n35055;
  assign n35057 = ~n35051 & ~n35056;
  assign n35058 = ~pi207 & ~n35057;
  assign n35059 = pi1156 & ~n34798;
  assign n35060 = ~pi1156 & ~n34699;
  assign n35061 = n20405 & ~n35060;
  assign n35062 = ~n35059 & n35061;
  assign n35063 = ~pi1156 & ~n34798;
  assign n35064 = pi1156 & ~n34699;
  assign n35065 = n20407 & ~n35064;
  assign n35066 = ~n35063 & n35065;
  assign n35067 = ~n35062 & ~n35066;
  assign n35068 = pi792 & ~n35067;
  assign n35069 = ~pi1159 & ~n34955;
  assign n35070 = pi1159 & ~n34796;
  assign n35071 = pi619 & ~pi648;
  assign n35072 = ~n35070 & n35071;
  assign n35073 = ~n35069 & n35072;
  assign n35074 = pi1159 & ~n34955;
  assign n35075 = ~pi1159 & ~n34796;
  assign n35076 = ~pi619 & pi648;
  assign n35077 = ~n35075 & n35076;
  assign n35078 = ~n35074 & n35077;
  assign n35079 = pi789 & ~n35078;
  assign n35080 = ~n35073 & n35079;
  assign n35081 = pi789 & ~n35080;
  assign n35082 = ~pi1154 & ~n34947;
  assign n35083 = n20072 & n34795;
  assign n35084 = ~pi627 & ~n35083;
  assign n35085 = ~n35082 & n35084;
  assign n35086 = ~pi778 & ~n33814;
  assign n35087 = pi625 & n33814;
  assign n35088 = ~pi625 & n34793;
  assign n35089 = pi1153 & ~n35088;
  assign n35090 = ~n35087 & n35089;
  assign n35091 = n34918 & ~n35090;
  assign n35092 = ~pi625 & n33814;
  assign n35093 = pi625 & n34793;
  assign n35094 = ~pi1153 & ~n35093;
  assign n35095 = ~n35092 & n35094;
  assign n35096 = n34924 & ~n35095;
  assign n35097 = pi778 & ~n35096;
  assign n35098 = ~n35091 & n35097;
  assign n35099 = ~n35086 & ~n35098;
  assign n35100 = ~pi785 & ~n35099;
  assign n35101 = ~pi609 & ~n35099;
  assign n35102 = ~pi1155 & ~n34930;
  assign n35103 = ~n35101 & n35102;
  assign n35104 = n20066 & n34794;
  assign n35105 = ~pi660 & ~n35104;
  assign n35106 = ~n35103 & n35105;
  assign n35107 = pi609 & ~n35099;
  assign n35108 = pi1155 & ~n34934;
  assign n35109 = ~n35107 & n35108;
  assign n35110 = n20067 & n34794;
  assign n35111 = pi660 & ~n35110;
  assign n35112 = ~n35109 & n35111;
  assign n35113 = ~n35106 & ~n35112;
  assign n35114 = pi785 & ~n35113;
  assign n35115 = ~n35100 & ~n35114;
  assign n35116 = pi618 & ~n35115;
  assign n35117 = pi1154 & ~n34943;
  assign n35118 = ~n35116 & n35117;
  assign n35119 = n20073 & n34795;
  assign n35120 = pi627 & ~n35119;
  assign n35121 = ~n35118 & n35120;
  assign n35122 = ~n35085 & ~n35121;
  assign n35123 = pi781 & ~n35122;
  assign n35124 = ~pi618 & ~pi627;
  assign n35125 = pi781 & ~n35124;
  assign n35126 = ~n35115 & ~n35125;
  assign n35127 = ~n23443 & n35080;
  assign n35128 = ~n35126 & ~n35127;
  assign n35129 = ~n35123 & n35128;
  assign n35130 = ~n35081 & ~n35129;
  assign n35131 = ~pi626 & n35130;
  assign n35132 = n34967 & ~n35131;
  assign n35133 = n17701 & n34797;
  assign n35134 = ~pi1158 & ~n35133;
  assign n35135 = ~n35132 & n35134;
  assign n35136 = pi626 & n35130;
  assign n35137 = n34962 & ~n35136;
  assign n35138 = n17702 & n34797;
  assign n35139 = pi1158 & ~n35138;
  assign n35140 = ~n35137 & n35139;
  assign n35141 = ~n35135 & ~n35140;
  assign n35142 = pi788 & ~n35141;
  assign n35143 = ~pi788 & n35130;
  assign n35144 = ~n20205 & ~n35143;
  assign n35145 = ~n35142 & n35144;
  assign n35146 = ~n35068 & ~n35145;
  assign n35147 = pi207 & ~n35146;
  assign n35148 = pi623 & ~n35147;
  assign n35149 = ~n35058 & n35148;
  assign n35150 = pi710 & ~n35149;
  assign n35151 = ~n34980 & n35150;
  assign n35152 = ~pi710 & ~n34804;
  assign n35153 = n20207 & ~n35152;
  assign n35154 = ~n35151 & n35153;
  assign n35155 = ~n34808 & ~n35154;
  assign n35156 = pi644 & n35155;
  assign n35157 = ~pi787 & ~n34735;
  assign n35158 = ~n34739 & ~n34744;
  assign n35159 = pi787 & ~n35158;
  assign n35160 = ~n35157 & ~n35159;
  assign n35161 = ~pi644 & n35160;
  assign n35162 = pi715 & ~n35161;
  assign n35163 = ~n35156 & n35162;
  assign n35164 = n17652 & ~n34733;
  assign n35165 = ~n17652 & n34804;
  assign n35166 = ~n35164 & ~n35165;
  assign n35167 = pi644 & n35166;
  assign n35168 = ~pi644 & n34733;
  assign n35169 = ~pi715 & ~n35168;
  assign n35170 = ~n35167 & n35169;
  assign n35171 = pi1160 & ~n35170;
  assign n35172 = ~n35163 & n35171;
  assign n35173 = ~pi644 & n35155;
  assign n35174 = pi644 & n35160;
  assign n35175 = ~pi715 & ~n35174;
  assign n35176 = ~n35173 & n35175;
  assign n35177 = ~pi644 & n35166;
  assign n35178 = pi644 & n34733;
  assign n35179 = pi715 & ~n35178;
  assign n35180 = ~n35177 & n35179;
  assign n35181 = ~pi1160 & ~n35180;
  assign n35182 = ~n35176 & n35181;
  assign n35183 = ~n35172 & ~n35182;
  assign n35184 = pi790 & ~n35183;
  assign n35185 = ~pi790 & n35155;
  assign n35186 = ~n35184 & ~n35185;
  assign n35187 = ~po1038 & ~n35186;
  assign n35188 = ~pi207 & po1038;
  assign po364 = n35187 | n35188;
  assign n35190 = pi208 & ~n34700;
  assign n35191 = ~pi208 & ~n34729;
  assign n35192 = ~n35190 & ~n35191;
  assign n35193 = pi638 & ~n35192;
  assign n35194 = ~pi208 & ~n17406;
  assign n35195 = ~pi638 & ~n35194;
  assign n35196 = ~n35193 & ~n35195;
  assign n35197 = ~pi647 & n35196;
  assign n35198 = pi647 & n35194;
  assign n35199 = ~pi1157 & ~n35198;
  assign n35200 = ~n35197 & n35199;
  assign n35201 = pi630 & n35200;
  assign n35202 = pi647 & n35196;
  assign n35203 = ~pi647 & n35194;
  assign n35204 = pi1157 & ~n35203;
  assign n35205 = ~n35202 & n35204;
  assign n35206 = ~pi630 & n35205;
  assign n35207 = ~pi208 & ~n34791;
  assign n35208 = pi208 & ~n34799;
  assign n35209 = pi607 & ~n35208;
  assign n35210 = ~n35207 & n35209;
  assign n35211 = ~pi607 & n35194;
  assign n35212 = ~n35210 & ~n35211;
  assign n35213 = ~n20398 & n35212;
  assign n35214 = ~n35206 & ~n35213;
  assign n35215 = ~n35201 & n35214;
  assign n35216 = pi787 & ~n35215;
  assign n35217 = ~pi208 & ~n34911;
  assign n35218 = pi208 & ~n34977;
  assign n35219 = ~pi607 & ~n35218;
  assign n35220 = ~n35217 & n35219;
  assign n35221 = ~pi208 & ~n35057;
  assign n35222 = pi208 & ~n35146;
  assign n35223 = pi607 & ~n35222;
  assign n35224 = ~n35221 & n35223;
  assign n35225 = pi638 & ~n35224;
  assign n35226 = ~n35220 & n35225;
  assign n35227 = ~pi638 & ~n35212;
  assign n35228 = n20207 & ~n35227;
  assign n35229 = ~n35226 & n35228;
  assign n35230 = ~n35216 & ~n35229;
  assign n35231 = pi644 & n35230;
  assign n35232 = ~pi787 & ~n35196;
  assign n35233 = ~n35200 & ~n35205;
  assign n35234 = pi787 & ~n35233;
  assign n35235 = ~n35232 & ~n35234;
  assign n35236 = ~pi644 & n35235;
  assign n35237 = pi715 & ~n35236;
  assign n35238 = ~n35231 & n35237;
  assign n35239 = n17652 & ~n35194;
  assign n35240 = ~n17652 & n35212;
  assign n35241 = ~n35239 & ~n35240;
  assign n35242 = pi644 & n35241;
  assign n35243 = ~pi644 & n35194;
  assign n35244 = ~pi715 & ~n35243;
  assign n35245 = ~n35242 & n35244;
  assign n35246 = pi1160 & ~n35245;
  assign n35247 = ~n35238 & n35246;
  assign n35248 = ~pi644 & n35230;
  assign n35249 = pi644 & n35235;
  assign n35250 = ~pi715 & ~n35249;
  assign n35251 = ~n35248 & n35250;
  assign n35252 = ~pi644 & n35241;
  assign n35253 = pi644 & n35194;
  assign n35254 = pi715 & ~n35253;
  assign n35255 = ~n35252 & n35254;
  assign n35256 = ~pi1160 & ~n35255;
  assign n35257 = ~n35251 & n35256;
  assign n35258 = ~n35247 & ~n35257;
  assign n35259 = pi790 & ~n35258;
  assign n35260 = ~pi790 & n35230;
  assign n35261 = ~n35259 & ~n35260;
  assign n35262 = ~po1038 & ~n35261;
  assign n35263 = ~pi208 & po1038;
  assign po365 = n35262 | n35263;
  assign n35265 = n20207 & ~n34911;
  assign n35266 = ~pi647 & ~n17406;
  assign n35267 = pi647 & n34729;
  assign n35268 = ~n35266 & ~n35267;
  assign n35269 = ~pi630 & ~n35268;
  assign n35270 = ~n35266 & ~n35269;
  assign n35271 = pi1157 & ~n35270;
  assign n35272 = pi647 & ~n17406;
  assign n35273 = ~pi1157 & n35272;
  assign n35274 = ~pi647 & n34729;
  assign n35275 = ~n35272 & ~n35274;
  assign n35276 = n17650 & ~n35275;
  assign n35277 = ~n35273 & ~n35276;
  assign n35278 = ~n35271 & n35277;
  assign n35279 = pi787 & ~n35278;
  assign n35280 = ~n35265 & ~n35279;
  assign n35281 = ~pi644 & ~n35280;
  assign n35282 = ~n19182 & n34729;
  assign n35283 = ~n17406 & n19182;
  assign n35284 = ~n35282 & ~n35283;
  assign n35285 = pi644 & ~n35284;
  assign n35286 = ~pi715 & ~n35285;
  assign n35287 = ~n35281 & n35286;
  assign n35288 = pi715 & n17406;
  assign n35289 = ~pi1160 & ~n35288;
  assign n35290 = ~n35287 & n35289;
  assign n35291 = pi644 & ~n35280;
  assign n35292 = ~pi644 & ~n35284;
  assign n35293 = pi715 & ~n35292;
  assign n35294 = ~n35291 & n35293;
  assign n35295 = ~pi715 & n17406;
  assign n35296 = pi1160 & ~n35295;
  assign n35297 = ~n35294 & n35296;
  assign n35298 = ~n35290 & ~n35297;
  assign n35299 = pi790 & ~n35298;
  assign n35300 = ~pi790 & ~n35280;
  assign n35301 = ~po1038 & ~n35300;
  assign n35302 = ~n35299 & n35301;
  assign n35303 = pi639 & n35302;
  assign n35304 = n10143 & n17399;
  assign n35305 = ~pi639 & n35304;
  assign n35306 = ~pi622 & ~n35305;
  assign n35307 = ~n35303 & n35306;
  assign n35308 = n20207 & ~n35057;
  assign n35309 = pi1157 & n35269;
  assign n35310 = ~n20398 & n34791;
  assign n35311 = ~n35276 & ~n35310;
  assign n35312 = ~n35309 & n35311;
  assign n35313 = pi787 & ~n35312;
  assign n35314 = ~n35308 & ~n35313;
  assign n35315 = ~pi644 & ~n35314;
  assign n35316 = n35286 & ~n35315;
  assign n35317 = ~n17406 & n17652;
  assign n35318 = ~n17652 & n34791;
  assign n35319 = ~n35317 & ~n35318;
  assign n35320 = ~pi644 & ~n35319;
  assign n35321 = pi644 & ~n17406;
  assign n35322 = ~n35320 & ~n35321;
  assign n35323 = pi715 & n35322;
  assign n35324 = ~pi1160 & ~n35323;
  assign n35325 = ~n35316 & n35324;
  assign n35326 = pi644 & ~n35314;
  assign n35327 = n35293 & ~n35326;
  assign n35328 = pi644 & ~n35319;
  assign n35329 = ~pi644 & ~n17406;
  assign n35330 = ~n35328 & ~n35329;
  assign n35331 = ~pi715 & n35330;
  assign n35332 = pi1160 & ~n35331;
  assign n35333 = ~n35327 & n35332;
  assign n35334 = ~n35325 & ~n35333;
  assign n35335 = pi790 & ~n35334;
  assign n35336 = ~pi790 & ~n35314;
  assign n35337 = ~po1038 & ~n35336;
  assign n35338 = ~n35335 & n35337;
  assign n35339 = pi639 & n35338;
  assign n35340 = ~pi1160 & n35322;
  assign n35341 = pi1160 & n35330;
  assign n35342 = pi790 & ~n35341;
  assign n35343 = ~n35340 & n35342;
  assign n35344 = ~pi790 & ~n35319;
  assign n35345 = ~po1038 & ~n35344;
  assign n35346 = ~n35343 & n35345;
  assign n35347 = ~pi639 & n35346;
  assign n35348 = pi622 & ~n35347;
  assign n35349 = ~n35339 & n35348;
  assign n35350 = ~n35307 & ~n35349;
  assign n35351 = ~pi209 & ~n35350;
  assign n35352 = ~n19182 & n34700;
  assign n35353 = pi644 & ~n35352;
  assign n35354 = ~pi715 & ~n35353;
  assign n35355 = ~pi647 & ~n35146;
  assign n35356 = pi647 & n34799;
  assign n35357 = ~pi1157 & ~n35356;
  assign n35358 = ~n35355 & n35357;
  assign n35359 = pi647 & n34700;
  assign n35360 = pi1157 & ~n35359;
  assign n35361 = ~pi630 & ~n35360;
  assign n35362 = ~n35358 & n35361;
  assign n35363 = pi647 & ~n35146;
  assign n35364 = ~pi647 & n34799;
  assign n35365 = pi1157 & ~n35364;
  assign n35366 = ~n35363 & n35365;
  assign n35367 = ~pi647 & n34700;
  assign n35368 = ~pi1157 & ~n35367;
  assign n35369 = pi630 & ~n35368;
  assign n35370 = ~n35366 & n35369;
  assign n35371 = ~n35362 & ~n35370;
  assign n35372 = pi787 & ~n35371;
  assign n35373 = ~pi787 & ~n35146;
  assign n35374 = ~n35372 & ~n35373;
  assign n35375 = ~pi644 & n35374;
  assign n35376 = n35354 & ~n35375;
  assign n35377 = n23518 & n34798;
  assign n35378 = ~pi644 & pi715;
  assign n35379 = n35377 & n35378;
  assign n35380 = ~pi1160 & ~n35379;
  assign n35381 = ~n35376 & n35380;
  assign n35382 = ~pi644 & ~n35352;
  assign n35383 = pi715 & ~n35382;
  assign n35384 = pi644 & n35374;
  assign n35385 = n35383 & ~n35384;
  assign n35386 = pi644 & ~pi715;
  assign n35387 = n35377 & n35386;
  assign n35388 = pi1160 & ~n35387;
  assign n35389 = ~n35385 & n35388;
  assign n35390 = ~n35381 & ~n35389;
  assign n35391 = pi790 & ~n35390;
  assign n35392 = ~pi790 & n35374;
  assign n35393 = ~po1038 & ~n35392;
  assign n35394 = ~n35391 & n35393;
  assign n35395 = pi622 & pi639;
  assign n35396 = ~n35394 & n35395;
  assign n35397 = n20207 & ~n34977;
  assign n35398 = n17652 & n19181;
  assign n35399 = n34700 & n35398;
  assign n35400 = ~n35397 & ~n35399;
  assign n35401 = ~pi644 & n35400;
  assign n35402 = ~pi1160 & n35354;
  assign n35403 = ~n35401 & n35402;
  assign n35404 = pi644 & n35400;
  assign n35405 = pi1160 & n35383;
  assign n35406 = ~n35404 & n35405;
  assign n35407 = pi790 & ~n35406;
  assign n35408 = ~n35403 & n35407;
  assign n35409 = ~pi790 & n35400;
  assign n35410 = ~po1038 & ~n35409;
  assign n35411 = ~n35408 & n35410;
  assign n35412 = ~pi622 & ~n35411;
  assign n35413 = ~pi644 & pi1160;
  assign n35414 = pi644 & ~pi1160;
  assign n35415 = ~n35413 & ~n35414;
  assign n35416 = pi790 & ~n35415;
  assign n35417 = ~po1038 & ~n35416;
  assign n35418 = n35377 & n35417;
  assign n35419 = pi622 & n35418;
  assign n35420 = ~pi639 & ~n35419;
  assign n35421 = pi209 & ~n35420;
  assign n35422 = ~n35412 & n35421;
  assign n35423 = ~n35396 & n35422;
  assign po366 = n35351 | n35423;
  assign n35425 = pi634 & n20755;
  assign n35426 = pi633 & pi947;
  assign n35427 = ~n35425 & ~n35426;
  assign n35428 = n17280 & ~n35427;
  assign n35429 = pi210 & ~n17280;
  assign n35430 = pi38 & ~n35429;
  assign n35431 = ~n35428 & n35430;
  assign n35432 = pi210 & ~n16518;
  assign n35433 = ~po1101 & n35432;
  assign n35434 = pi210 & po1101;
  assign n35435 = ~n16621 & n35434;
  assign n35436 = ~n35433 & ~n35435;
  assign n35437 = ~pi907 & n35436;
  assign n35438 = pi634 & n16518;
  assign n35439 = ~n35432 & ~n35438;
  assign n35440 = ~n6198 & ~n35439;
  assign n35441 = pi907 & ~n35440;
  assign n35442 = pi210 & n16619;
  assign n35443 = pi634 & ~n16619;
  assign n35444 = ~n35442 & ~n35443;
  assign n35445 = n6198 & ~n35444;
  assign n35446 = n35441 & ~n35445;
  assign n35447 = ~pi947 & ~n35446;
  assign n35448 = ~n35437 & n35447;
  assign n35449 = ~n33221 & ~n35432;
  assign n35450 = ~po1101 & n35449;
  assign n35451 = pi947 & ~n35450;
  assign n35452 = po1101 & n35449;
  assign n35453 = ~n6198 & ~n35452;
  assign n35454 = pi633 & ~n16619;
  assign n35455 = ~n35442 & ~n35454;
  assign n35456 = ~n6162 & ~n35455;
  assign n35457 = ~n35453 & ~n35456;
  assign n35458 = n35451 & ~n35457;
  assign n35459 = n6215 & ~n35458;
  assign n35460 = ~n35448 & n35459;
  assign n35461 = n6192 & n35439;
  assign n35462 = pi907 & ~n35461;
  assign n35463 = ~n6192 & n35444;
  assign n35464 = n35462 & ~n35463;
  assign n35465 = pi210 & ~n16812;
  assign n35466 = ~pi907 & n35465;
  assign n35467 = ~n35464 & ~n35466;
  assign n35468 = ~pi947 & ~n35467;
  assign n35469 = n6192 & n35449;
  assign n35470 = pi947 & ~n35469;
  assign n35471 = ~n6192 & n35455;
  assign n35472 = n35470 & ~n35471;
  assign n35473 = ~n6215 & ~n35472;
  assign n35474 = ~n35468 & n35473;
  assign n35475 = ~n35460 & ~n35474;
  assign n35476 = ~n3052 & ~n35475;
  assign n35477 = n16518 & ~n35427;
  assign n35478 = ~n35432 & ~n35477;
  assign n35479 = n3052 & n35478;
  assign n35480 = ~pi223 & ~n35479;
  assign n35481 = ~n35476 & n35480;
  assign n35482 = ~n16569 & n35434;
  assign n35483 = ~n35433 & ~n35482;
  assign n35484 = ~pi907 & n35483;
  assign n35485 = pi210 & n16542;
  assign n35486 = ~n33407 & ~n35485;
  assign n35487 = n6198 & ~n35486;
  assign n35488 = n35441 & ~n35487;
  assign n35489 = ~pi947 & ~n35488;
  assign n35490 = ~n35484 & n35489;
  assign n35491 = pi633 & ~n16542;
  assign n35492 = ~n35485 & ~n35491;
  assign n35493 = ~n6162 & ~n35492;
  assign n35494 = ~n35453 & ~n35493;
  assign n35495 = n35451 & ~n35494;
  assign n35496 = n6215 & ~n35495;
  assign n35497 = ~n35490 & n35496;
  assign n35498 = ~n6192 & n35486;
  assign n35499 = n35462 & ~n35498;
  assign n35500 = n6192 & n16517;
  assign n35501 = n2754 & n35500;
  assign n35502 = n35485 & ~n35501;
  assign n35503 = ~n35499 & ~n35502;
  assign n35504 = ~pi947 & ~n35503;
  assign n35505 = ~n6192 & n35492;
  assign n35506 = n35470 & ~n35505;
  assign n35507 = ~n6215 & ~n35506;
  assign n35508 = ~n35504 & n35507;
  assign n35509 = pi223 & ~n35508;
  assign n35510 = ~n35497 & n35509;
  assign n35511 = ~pi299 & ~n35510;
  assign n35512 = ~n35481 & n35511;
  assign n35513 = ~n6188 & ~n35465;
  assign n35514 = n6188 & n35436;
  assign n35515 = ~pi907 & ~n35514;
  assign n35516 = ~n35513 & n35515;
  assign n35517 = ~n35464 & ~n35516;
  assign n35518 = ~pi947 & ~n35517;
  assign n35519 = ~n3329 & ~n35472;
  assign n35520 = ~n35518 & n35519;
  assign n35521 = n3329 & n35478;
  assign n35522 = ~pi215 & ~n35521;
  assign n35523 = ~n35520 & n35522;
  assign n35524 = n6188 & n35483;
  assign n35525 = ~n6188 & ~n35502;
  assign n35526 = ~pi907 & ~n35525;
  assign n35527 = ~n35524 & n35526;
  assign n35528 = ~n35499 & ~n35527;
  assign n35529 = ~pi947 & ~n35528;
  assign n35530 = ~n35506 & ~n35529;
  assign n35531 = pi215 & ~n35530;
  assign n35532 = pi299 & ~n35531;
  assign n35533 = ~n35523 & n35532;
  assign n35534 = pi39 & ~n35533;
  assign n35535 = ~n35512 & n35534;
  assign n35536 = n17063 & ~n35427;
  assign n35537 = pi210 & ~n17063;
  assign n35538 = ~pi299 & ~n35537;
  assign n35539 = ~n35536 & n35538;
  assign n35540 = ~n17022 & ~n35427;
  assign n35541 = pi299 & ~n35540;
  assign n35542 = ~n17025 & n35541;
  assign n35543 = ~pi39 & ~n35542;
  assign n35544 = ~n35539 & n35543;
  assign n35545 = ~pi38 & ~n35544;
  assign n35546 = ~n35535 & n35545;
  assign n35547 = ~n35431 & ~n35546;
  assign n35548 = n10143 & ~n35547;
  assign n35549 = ~pi210 & ~n10143;
  assign po367 = ~n35548 & ~n35549;
  assign n35551 = n3267 & ~n21475;
  assign n35552 = pi606 & n35551;
  assign n35553 = n3267 & ~n21471;
  assign n35554 = ~pi606 & n35553;
  assign n35555 = pi643 & ~n35554;
  assign n35556 = ~n35552 & n35555;
  assign n35557 = n3267 & ~n20849;
  assign n35558 = pi606 & n35557;
  assign n35559 = ~pi606 & n17406;
  assign n35560 = ~pi643 & ~n35559;
  assign n35561 = ~n35558 & n35560;
  assign n35562 = ~po1038 & ~n35561;
  assign n35563 = ~n35556 & n35562;
  assign n35564 = pi211 & ~n35563;
  assign n35565 = n3267 & n21460;
  assign n35566 = pi606 & ~n35565;
  assign n35567 = n3267 & n21457;
  assign n35568 = ~pi606 & ~n35567;
  assign n35569 = pi643 & ~n35568;
  assign n35570 = ~n35566 & n35569;
  assign n35571 = n3267 & n20873;
  assign n35572 = pi606 & ~pi643;
  assign n35573 = n35571 & n35572;
  assign n35574 = ~n35570 & ~n35573;
  assign n35575 = ~pi211 & ~po1038;
  assign n35576 = ~n35574 & n35575;
  assign po368 = n35564 | n35576;
  assign n35578 = pi607 & n35551;
  assign n35579 = ~pi607 & n35553;
  assign n35580 = pi638 & ~n35579;
  assign n35581 = ~n35578 & n35580;
  assign n35582 = pi607 & n35557;
  assign n35583 = ~pi607 & n17406;
  assign n35584 = ~pi638 & ~n35583;
  assign n35585 = ~n35582 & n35584;
  assign n35586 = ~po1038 & ~n35585;
  assign n35587 = ~n35581 & n35586;
  assign n35588 = ~pi212 & ~n35587;
  assign n35589 = ~pi607 & ~n35567;
  assign n35590 = pi607 & ~n35565;
  assign n35591 = pi638 & ~n35590;
  assign n35592 = ~n35589 & n35591;
  assign n35593 = pi607 & ~pi638;
  assign n35594 = n35571 & n35593;
  assign n35595 = ~n35592 & ~n35594;
  assign n35596 = pi212 & ~po1038;
  assign n35597 = ~n35595 & n35596;
  assign po369 = n35588 | n35597;
  assign n35599 = pi213 & ~po1038;
  assign n35600 = ~pi622 & ~n35567;
  assign n35601 = pi622 & ~n35565;
  assign n35602 = pi639 & ~n35601;
  assign n35603 = ~n35600 & n35602;
  assign n35604 = pi622 & ~pi639;
  assign n35605 = n35571 & n35604;
  assign n35606 = ~n35603 & ~n35605;
  assign n35607 = n35599 & ~n35606;
  assign n35608 = pi639 & n35551;
  assign n35609 = ~pi639 & n35557;
  assign n35610 = pi622 & ~n35609;
  assign n35611 = ~n35608 & n35610;
  assign n35612 = pi639 & n35553;
  assign n35613 = ~pi639 & n17406;
  assign n35614 = ~pi622 & ~n35613;
  assign n35615 = ~n35612 & n35614;
  assign n35616 = ~po1038 & ~n35615;
  assign n35617 = ~n35611 & n35616;
  assign n35618 = ~pi213 & ~n35617;
  assign po370 = n35607 | n35618;
  assign n35620 = pi623 & n35551;
  assign n35621 = ~pi623 & n35553;
  assign n35622 = pi710 & ~n35621;
  assign n35623 = ~n35620 & n35622;
  assign n35624 = pi623 & n35557;
  assign n35625 = ~pi623 & n17406;
  assign n35626 = ~pi710 & ~n35625;
  assign n35627 = ~n35624 & n35626;
  assign n35628 = ~po1038 & ~n35627;
  assign n35629 = ~n35623 & n35628;
  assign n35630 = ~pi214 & ~n35629;
  assign n35631 = ~pi623 & ~n35567;
  assign n35632 = pi623 & ~n35565;
  assign n35633 = pi710 & ~n35632;
  assign n35634 = ~n35631 & n35633;
  assign n35635 = pi623 & ~pi710;
  assign n35636 = n35571 & n35635;
  assign n35637 = ~n35634 & ~n35636;
  assign n35638 = pi214 & ~po1038;
  assign n35639 = ~n35637 & n35638;
  assign po371 = n35630 | n35639;
  assign n35641 = pi215 & ~n10143;
  assign n35642 = ~pi947 & n21149;
  assign n35643 = pi681 & pi907;
  assign n35644 = ~pi947 & n35643;
  assign n35645 = ~n6160 & n16585;
  assign n35646 = n16511 & n17124;
  assign n35647 = ~pi642 & ~n35646;
  assign n35648 = ~n35645 & n35647;
  assign n35649 = pi947 & ~n35648;
  assign n35650 = ~n35644 & ~n35649;
  assign n35651 = ~n35642 & n35650;
  assign n35652 = pi299 & ~n35651;
  assign n35653 = n21217 & ~n35643;
  assign n35654 = ~pi642 & n16621;
  assign n35655 = n6160 & ~n35654;
  assign n35656 = ~n6156 & n16518;
  assign n35657 = ~pi642 & n35656;
  assign n35658 = ~n6160 & ~n35657;
  assign n35659 = ~n16824 & n35658;
  assign n35660 = ~n35655 & ~n35659;
  assign n35661 = n6215 & ~n35660;
  assign n35662 = ~pi642 & n16812;
  assign n35663 = ~n6215 & ~n35662;
  assign n35664 = pi947 & ~n35663;
  assign n35665 = ~n35661 & n35664;
  assign n35666 = ~n3052 & ~n35665;
  assign n35667 = ~n35653 & n35666;
  assign n35668 = n3052 & ~n16518;
  assign n35669 = pi642 & pi947;
  assign n35670 = ~n35644 & ~n35669;
  assign n35671 = n3052 & ~n35670;
  assign n35672 = ~pi223 & ~n35671;
  assign n35673 = ~n35668 & n35672;
  assign n35674 = ~n35667 & n35673;
  assign n35675 = ~n6160 & ~n16575;
  assign n35676 = n6160 & ~n16569;
  assign n35677 = ~pi642 & ~n35676;
  assign n35678 = ~n35675 & n35677;
  assign n35679 = n6215 & ~n35678;
  assign n35680 = ~n6215 & ~n35648;
  assign n35681 = pi947 & ~n35680;
  assign n35682 = ~n35679 & n35681;
  assign n35683 = ~n21232 & ~n35682;
  assign n35684 = pi223 & ~n35644;
  assign n35685 = ~n35683 & n35684;
  assign n35686 = ~pi299 & ~n35685;
  assign n35687 = ~n35674 & n35686;
  assign n35688 = ~n35652 & ~n35687;
  assign n35689 = pi215 & ~n35688;
  assign n35690 = n16637 & n35644;
  assign n35691 = pi642 & ~n16512;
  assign n35692 = n16518 & n35691;
  assign n35693 = pi642 & n16512;
  assign n35694 = ~n17142 & n35693;
  assign n35695 = ~n17163 & n35694;
  assign n35696 = ~n35692 & ~n35695;
  assign n35697 = pi947 & ~n35696;
  assign n35698 = n6215 & ~n35697;
  assign n35699 = ~n35690 & n35698;
  assign n35700 = n16652 & n35643;
  assign n35701 = ~pi947 & ~n35700;
  assign n35702 = ~n6160 & n16649;
  assign n35703 = ~n16811 & ~n35702;
  assign n35704 = n35693 & n35703;
  assign n35705 = ~n16649 & n35691;
  assign n35706 = pi947 & ~n35705;
  assign n35707 = ~n35704 & n35706;
  assign n35708 = ~n35701 & ~n35707;
  assign n35709 = ~n6215 & ~n35708;
  assign n35710 = ~n3052 & ~n35709;
  assign n35711 = ~n35699 & n35710;
  assign n35712 = n16518 & n35671;
  assign n35713 = ~pi223 & ~n35712;
  assign n35714 = ~n35711 & n35713;
  assign n35715 = n6215 & ~n16575;
  assign n35716 = n35643 & ~n35715;
  assign n35717 = ~pi947 & ~n35716;
  assign n35718 = pi947 & ~n16583;
  assign n35719 = n16585 & ~n35718;
  assign n35720 = ~n6215 & n35719;
  assign n35721 = ~n17137 & n35694;
  assign n35722 = pi947 & ~n35692;
  assign n35723 = ~n35721 & n35722;
  assign n35724 = ~n35720 & ~n35723;
  assign n35725 = ~n35717 & n35724;
  assign n35726 = pi223 & ~n35725;
  assign n35727 = ~n35714 & ~n35726;
  assign n35728 = ~pi299 & ~n35727;
  assign n35729 = ~n3329 & n35708;
  assign n35730 = n16736 & ~n35670;
  assign n35731 = pi299 & ~n35730;
  assign n35732 = ~n35729 & n35731;
  assign n35733 = ~pi215 & ~n35732;
  assign n35734 = ~n35728 & n35733;
  assign n35735 = ~n35689 & ~n35734;
  assign n35736 = pi39 & ~n35735;
  assign n35737 = pi215 & ~n17063;
  assign n35738 = n17063 & ~n35670;
  assign n35739 = ~pi299 & ~n35738;
  assign n35740 = ~n35737 & n35739;
  assign n35741 = n17026 & ~n35670;
  assign n35742 = pi215 & ~n17026;
  assign n35743 = pi299 & ~n35742;
  assign n35744 = ~n35741 & n35743;
  assign n35745 = ~pi39 & ~n35744;
  assign n35746 = ~n35740 & n35745;
  assign n35747 = ~pi38 & ~n35746;
  assign n35748 = ~n35736 & n35747;
  assign n35749 = pi215 & ~n17280;
  assign n35750 = n17280 & ~n35670;
  assign n35751 = pi38 & ~n35750;
  assign n35752 = ~n35749 & n35751;
  assign n35753 = n10143 & ~n35752;
  assign n35754 = ~n35748 & n35753;
  assign po372 = n35641 | n35754;
  assign n35756 = pi216 & ~n17280;
  assign n35757 = pi662 & pi907;
  assign n35758 = ~pi947 & n35757;
  assign n35759 = pi614 & pi947;
  assign n35760 = ~n35758 & ~n35759;
  assign n35761 = n17280 & ~n35760;
  assign n35762 = pi38 & ~n35761;
  assign n35763 = ~n35756 & n35762;
  assign n35764 = ~pi947 & n20833;
  assign n35765 = ~pi614 & n16812;
  assign n35766 = pi947 & ~n35765;
  assign n35767 = ~n35758 & ~n35766;
  assign n35768 = ~n35764 & n35767;
  assign n35769 = pi216 & ~n35768;
  assign n35770 = n35703 & n35759;
  assign n35771 = n16652 & n35758;
  assign n35772 = ~n35770 & ~n35771;
  assign n35773 = n5745 & ~n35772;
  assign n35774 = n16736 & ~n35760;
  assign n35775 = ~n35773 & ~n35774;
  assign n35776 = ~n35769 & n35775;
  assign n35777 = ~pi215 & ~n35776;
  assign n35778 = ~pi614 & ~n16542;
  assign n35779 = n16584 & n17157;
  assign n35780 = ~n35778 & ~n35779;
  assign n35781 = pi947 & n35780;
  assign n35782 = pi216 & ~n35758;
  assign n35783 = ~n35781 & n35782;
  assign n35784 = ~n35642 & n35783;
  assign n35785 = ~n16585 & n35757;
  assign n35786 = ~pi947 & ~n35785;
  assign n35787 = ~n17137 & n17165;
  assign n35788 = pi947 & ~n17168;
  assign n35789 = ~n35787 & n35788;
  assign n35790 = pi947 & n16583;
  assign n35791 = ~n35789 & ~n35790;
  assign n35792 = ~n35786 & n35791;
  assign n35793 = ~pi216 & ~n35792;
  assign n35794 = pi215 & ~n35793;
  assign n35795 = ~n35784 & n35794;
  assign n35796 = pi299 & ~n35795;
  assign n35797 = ~n35777 & n35796;
  assign n35798 = pi947 & ~n17162;
  assign n35799 = ~pi947 & n17172;
  assign n35800 = ~n35757 & n35799;
  assign n35801 = ~n35798 & ~n35800;
  assign n35802 = n6215 & ~n35801;
  assign n35803 = ~pi947 & ~n16812;
  assign n35804 = ~n6215 & ~n35758;
  assign n35805 = ~n35766 & n35804;
  assign n35806 = ~n35803 & n35805;
  assign n35807 = ~n3052 & ~n35806;
  assign n35808 = ~n35802 & n35807;
  assign n35809 = n3052 & ~n35760;
  assign n35810 = ~pi223 & ~n35809;
  assign n35811 = ~n35668 & n35810;
  assign n35812 = ~n35808 & n35811;
  assign n35813 = ~pi614 & ~n35676;
  assign n35814 = ~n35675 & n35813;
  assign n35815 = n6215 & ~n35814;
  assign n35816 = ~n6215 & n35780;
  assign n35817 = pi947 & ~n35816;
  assign n35818 = ~n35815 & n35817;
  assign n35819 = ~n21232 & ~n35818;
  assign n35820 = pi223 & ~n35758;
  assign n35821 = ~n35819 & n35820;
  assign n35822 = pi216 & ~n35821;
  assign n35823 = ~n35812 & n35822;
  assign n35824 = n16637 & n35758;
  assign n35825 = pi947 & ~n17169;
  assign n35826 = n6215 & ~n35825;
  assign n35827 = ~n35824 & n35826;
  assign n35828 = ~n6215 & n35772;
  assign n35829 = ~n3052 & ~n35828;
  assign n35830 = ~n35827 & n35829;
  assign n35831 = n16518 & n35809;
  assign n35832 = ~pi223 & ~n35831;
  assign n35833 = ~n35830 & n35832;
  assign n35834 = ~n35715 & n35757;
  assign n35835 = ~pi947 & ~n35834;
  assign n35836 = ~n35720 & ~n35789;
  assign n35837 = ~n35835 & n35836;
  assign n35838 = pi223 & ~n35837;
  assign n35839 = ~pi216 & ~n35838;
  assign n35840 = ~n35833 & n35839;
  assign n35841 = ~pi299 & ~n35840;
  assign n35842 = ~n35823 & n35841;
  assign n35843 = pi39 & ~n35842;
  assign n35844 = ~n35797 & n35843;
  assign n35845 = pi216 & ~n17063;
  assign n35846 = n17063 & ~n35760;
  assign n35847 = ~pi299 & ~n35846;
  assign n35848 = ~n35845 & n35847;
  assign n35849 = n17026 & ~n35760;
  assign n35850 = pi216 & ~n17026;
  assign n35851 = pi299 & ~n35850;
  assign n35852 = ~n35849 & n35851;
  assign n35853 = ~pi39 & ~n35852;
  assign n35854 = ~n35848 & n35853;
  assign n35855 = ~pi38 & ~n35854;
  assign n35856 = ~n35844 & n35855;
  assign n35857 = ~n35763 & ~n35856;
  assign n35858 = n10143 & ~n35857;
  assign n35859 = ~pi216 & ~n10143;
  assign po373 = ~n35858 & ~n35859;
  assign n35861 = ~pi695 & ~n35302;
  assign n35862 = pi695 & ~n35304;
  assign n35863 = ~pi217 & ~n35862;
  assign n35864 = ~n35861 & n35863;
  assign n35865 = ~pi695 & n35411;
  assign n35866 = pi217 & ~n35865;
  assign n35867 = ~pi612 & ~n35866;
  assign n35868 = ~n35864 & n35867;
  assign n35869 = ~pi695 & ~n35338;
  assign n35870 = pi695 & ~n35346;
  assign n35871 = ~pi217 & ~n35870;
  assign n35872 = ~n35869 & n35871;
  assign n35873 = ~pi695 & n35394;
  assign n35874 = pi695 & n35418;
  assign n35875 = pi217 & ~n35874;
  assign n35876 = ~n35873 & n35875;
  assign n35877 = pi612 & ~n35876;
  assign n35878 = ~n35872 & n35877;
  assign po374 = n35868 | n35878;
  assign n35880 = ~n34567 & ~n34606;
  assign n35881 = n34567 & ~n34672;
  assign n35882 = ~n35880 & ~n35881;
  assign n35883 = ~pi218 & ~n35882;
  assign n35884 = n34567 & n34679;
  assign n35885 = pi218 & ~n35884;
  assign po375 = ~n35883 & ~n35885;
  assign n35887 = ~pi219 & ~po1038;
  assign n35888 = ~pi617 & ~n35567;
  assign n35889 = pi617 & ~n35565;
  assign n35890 = pi637 & ~n35889;
  assign n35891 = ~n35888 & n35890;
  assign n35892 = pi617 & ~pi637;
  assign n35893 = n35571 & n35892;
  assign n35894 = ~n35891 & ~n35893;
  assign n35895 = n35887 & ~n35894;
  assign n35896 = pi617 & n35551;
  assign n35897 = ~pi617 & n35553;
  assign n35898 = pi637 & ~n35897;
  assign n35899 = ~n35896 & n35898;
  assign n35900 = pi617 & n35557;
  assign n35901 = ~pi617 & n17406;
  assign n35902 = ~pi637 & ~n35901;
  assign n35903 = ~n35900 & n35902;
  assign n35904 = ~po1038 & ~n35903;
  assign n35905 = ~n35899 & n35904;
  assign n35906 = pi219 & ~n35905;
  assign po376 = n35895 | n35906;
  assign n35908 = ~n34400 & ~n34690;
  assign n35909 = ~n34545 & n34690;
  assign n35910 = ~n35908 & ~n35909;
  assign n35911 = ~pi220 & ~n35910;
  assign n35912 = n34555 & n34690;
  assign n35913 = pi220 & ~n35912;
  assign po377 = ~n35911 & ~n35913;
  assign n35915 = pi221 & ~n17280;
  assign n35916 = pi616 & pi947;
  assign n35917 = pi661 & n20755;
  assign n35918 = ~n35916 & ~n35917;
  assign n35919 = n17280 & ~n35918;
  assign n35920 = pi38 & ~n35919;
  assign n35921 = ~n35915 & n35920;
  assign n35922 = n35703 & n35916;
  assign n35923 = n16652 & n35917;
  assign n35924 = ~n35922 & ~n35923;
  assign n35925 = pi216 & ~n35924;
  assign n35926 = n16518 & ~n35918;
  assign n35927 = ~pi216 & n35926;
  assign n35928 = ~pi221 & ~n35927;
  assign n35929 = ~n35925 & n35928;
  assign n35930 = ~pi215 & ~n35929;
  assign n35931 = ~n6162 & n16635;
  assign n35932 = ~n16648 & ~n35931;
  assign n35933 = n17135 & ~n35932;
  assign n35934 = ~n35662 & ~n35704;
  assign n35935 = n17138 & ~n35934;
  assign n35936 = pi947 & ~n35935;
  assign n35937 = ~n35933 & n35936;
  assign n35938 = pi221 & ~n35917;
  assign n35939 = ~n35937 & n35938;
  assign n35940 = ~n35764 & n35939;
  assign n35941 = n35930 & ~n35940;
  assign n35942 = ~pi616 & ~n35646;
  assign n35943 = ~n35645 & n35942;
  assign n35944 = pi947 & ~n35943;
  assign n35945 = n35938 & ~n35944;
  assign n35946 = ~n35642 & n35945;
  assign n35947 = pi947 & ~n17148;
  assign n35948 = ~n35917 & ~n35947;
  assign n35949 = ~n35719 & ~n35948;
  assign n35950 = ~pi221 & ~n35949;
  assign n35951 = pi215 & ~n35950;
  assign n35952 = ~n35946 & n35951;
  assign n35953 = pi299 & ~n35952;
  assign n35954 = ~n35941 & n35953;
  assign n35955 = n16635 & n17135;
  assign n35956 = n17162 & ~n17166;
  assign n35957 = n17138 & ~n35956;
  assign n35958 = ~n35955 & ~n35957;
  assign n35959 = pi947 & ~n35958;
  assign n35960 = n6215 & ~n35799;
  assign n35961 = ~n35959 & n35960;
  assign n35962 = ~n35803 & ~n35937;
  assign n35963 = ~n6215 & ~n35962;
  assign n35964 = ~n35917 & ~n35963;
  assign n35965 = ~n35961 & n35964;
  assign n35966 = ~n3052 & ~n35965;
  assign n35967 = n3052 & n35926;
  assign n35968 = ~pi223 & ~n35967;
  assign n35969 = ~n35668 & n35968;
  assign n35970 = ~n35966 & n35969;
  assign n35971 = ~pi947 & ~n17132;
  assign n35972 = ~n35944 & ~n35971;
  assign n35973 = ~n6215 & ~n35972;
  assign n35974 = ~pi947 & n17151;
  assign n35975 = pi947 & ~n17141;
  assign n35976 = n6215 & ~n35975;
  assign n35977 = ~n35974 & n35976;
  assign n35978 = pi223 & ~n35917;
  assign n35979 = ~n35977 & n35978;
  assign n35980 = ~n35973 & n35979;
  assign n35981 = pi221 & ~n35980;
  assign n35982 = ~n35970 & n35981;
  assign n35983 = n16637 & n35917;
  assign n35984 = n17144 & ~n17163;
  assign n35985 = ~n17147 & ~n35984;
  assign n35986 = pi947 & ~n35985;
  assign n35987 = n6215 & ~n35986;
  assign n35988 = ~n35983 & n35987;
  assign n35989 = ~n6215 & n35924;
  assign n35990 = ~n3052 & ~n35989;
  assign n35991 = ~n35988 & n35990;
  assign n35992 = n35968 & ~n35991;
  assign n35993 = n35715 & ~n35947;
  assign n35994 = ~n35720 & ~n35948;
  assign n35995 = ~n35993 & n35994;
  assign n35996 = pi223 & ~n35995;
  assign n35997 = ~pi221 & ~n35996;
  assign n35998 = ~n35992 & n35997;
  assign n35999 = ~pi299 & ~n35998;
  assign n36000 = ~n35982 & n35999;
  assign n36001 = pi39 & ~n36000;
  assign n36002 = ~n35954 & n36001;
  assign n36003 = pi221 & ~n17063;
  assign n36004 = n17063 & ~n35918;
  assign n36005 = ~pi299 & ~n36004;
  assign n36006 = ~n36003 & n36005;
  assign n36007 = n17026 & ~n35918;
  assign n36008 = pi221 & ~n17026;
  assign n36009 = pi299 & ~n36008;
  assign n36010 = ~n36007 & n36009;
  assign n36011 = ~pi39 & ~n36010;
  assign n36012 = ~n36006 & n36011;
  assign n36013 = ~pi38 & ~n36012;
  assign n36014 = ~n36002 & n36013;
  assign n36015 = ~n35921 & ~n36014;
  assign n36016 = n10143 & ~n36015;
  assign n36017 = ~pi221 & ~n10143;
  assign po378 = ~n36016 & ~n36017;
  assign n36019 = ~pi223 & ~n17175;
  assign n36020 = ~n17154 & ~n36019;
  assign n36021 = ~pi299 & ~n36020;
  assign n36022 = pi39 & ~n36021;
  assign n36023 = ~n17198 & n36022;
  assign n36024 = ~pi38 & ~n17954;
  assign n36025 = ~n36023 & n36024;
  assign n36026 = n18723 & ~n36025;
  assign n36027 = pi222 & ~n36026;
  assign n36028 = n17816 & ~n36027;
  assign n36029 = pi222 & ~n3267;
  assign n36030 = pi616 & n16521;
  assign n36031 = ~n33277 & ~n36030;
  assign n36032 = n16652 & n36031;
  assign n36033 = ~n16511 & ~n36032;
  assign n36034 = ~n6158 & n36032;
  assign n36035 = n16656 & ~n36030;
  assign n36036 = ~n16695 & ~n36035;
  assign n36037 = n6158 & ~n36036;
  assign n36038 = n16511 & ~n36037;
  assign n36039 = ~n36034 & n36038;
  assign n36040 = ~n36033 & ~n36039;
  assign n36041 = ~n6215 & n36040;
  assign n36042 = pi616 & ~n16713;
  assign n36043 = ~n16636 & ~n36042;
  assign n36044 = ~n16511 & ~n36043;
  assign n36045 = ~n6158 & n36043;
  assign n36046 = n6158 & ~n36030;
  assign n36047 = n16621 & n36046;
  assign n36048 = n16511 & ~n36047;
  assign n36049 = ~n36045 & n36048;
  assign n36050 = ~n36044 & ~n36049;
  assign n36051 = n6215 & n36050;
  assign n36052 = pi222 & ~n36051;
  assign n36053 = ~n36041 & n36052;
  assign n36054 = ~n16649 & n36030;
  assign n36055 = ~n16511 & ~n36054;
  assign n36056 = ~n6158 & n36054;
  assign n36057 = pi616 & n6158;
  assign n36058 = n16657 & n36057;
  assign n36059 = n16511 & ~n36058;
  assign n36060 = ~n36056 & n36059;
  assign n36061 = ~n36055 & ~n36060;
  assign n36062 = ~n6215 & n36061;
  assign n36063 = ~n6160 & n16543;
  assign n36064 = ~n17248 & ~n36063;
  assign n36065 = pi616 & ~n36064;
  assign n36066 = n6215 & n36065;
  assign n36067 = pi224 & ~n36066;
  assign n36068 = ~n36062 & n36067;
  assign n36069 = n16521 & n17146;
  assign n36070 = ~pi224 & ~n36069;
  assign n36071 = ~pi222 & ~n36070;
  assign n36072 = ~n36068 & n36071;
  assign n36073 = ~pi223 & ~n36072;
  assign n36074 = ~n36053 & n36073;
  assign n36075 = ~n16574 & ~n36042;
  assign n36076 = ~n16511 & ~n36075;
  assign n36077 = ~n6158 & n36075;
  assign n36078 = n16569 & n36046;
  assign n36079 = n16511 & ~n36078;
  assign n36080 = ~n36077 & n36079;
  assign n36081 = ~n36076 & ~n36080;
  assign n36082 = n6215 & n36081;
  assign n36083 = pi616 & ~n16740;
  assign n36084 = ~n16585 & ~n36083;
  assign n36085 = ~n17124 & ~n36083;
  assign n36086 = ~n16585 & n36085;
  assign n36087 = n16511 & ~n36086;
  assign n36088 = n36084 & ~n36087;
  assign n36089 = ~n6215 & n36088;
  assign n36090 = pi222 & ~n36089;
  assign n36091 = ~n36082 & n36090;
  assign n36092 = ~n16551 & ~n36063;
  assign n36093 = pi616 & ~n36092;
  assign n36094 = ~pi222 & n36093;
  assign n36095 = ~n17268 & n36094;
  assign n36096 = pi223 & ~n36095;
  assign n36097 = ~n36091 & n36096;
  assign n36098 = ~n36074 & ~n36097;
  assign n36099 = ~pi299 & ~n36098;
  assign n36100 = ~n6189 & n36040;
  assign n36101 = n6189 & n36050;
  assign n36102 = pi222 & ~n36101;
  assign n36103 = ~n36100 & n36102;
  assign n36104 = ~n6189 & ~n36061;
  assign n36105 = n6189 & ~n36065;
  assign n36106 = ~pi222 & ~n36105;
  assign n36107 = ~n36104 & n36106;
  assign n36108 = ~n3329 & ~n36107;
  assign n36109 = ~n36103 & n36108;
  assign n36110 = pi222 & ~n16518;
  assign n36111 = n3329 & ~n36110;
  assign n36112 = ~n36069 & n36111;
  assign n36113 = ~pi215 & ~n36112;
  assign n36114 = ~n36109 & n36113;
  assign n36115 = ~n17258 & n36094;
  assign n36116 = n6189 & n36081;
  assign n36117 = ~n6189 & n36088;
  assign n36118 = pi222 & ~n36117;
  assign n36119 = ~n36116 & n36118;
  assign n36120 = ~n36115 & ~n36119;
  assign n36121 = pi215 & ~n36120;
  assign n36122 = pi299 & ~n36121;
  assign n36123 = ~n36114 & n36122;
  assign n36124 = pi39 & ~n36123;
  assign n36125 = ~n36099 & n36124;
  assign n36126 = pi222 & n17042;
  assign n36127 = ~pi222 & ~n17086;
  assign n36128 = ~pi616 & n17086;
  assign n36129 = ~pi39 & ~n36128;
  assign n36130 = ~n36127 & n36129;
  assign n36131 = ~n36126 & n36130;
  assign n36132 = ~pi38 & ~n36131;
  assign n36133 = ~n36125 & n36132;
  assign n36134 = pi222 & ~n17280;
  assign n36135 = pi38 & ~n36134;
  assign n36136 = pi616 & n17282;
  assign n36137 = n36135 & ~n36136;
  assign n36138 = n3267 & ~n36137;
  assign n36139 = ~n36133 & n36138;
  assign n36140 = ~n36029 & ~n36139;
  assign n36141 = ~n17438 & ~n36140;
  assign n36142 = n17438 & n36027;
  assign n36143 = ~n36141 & ~n36142;
  assign n36144 = ~pi785 & ~n36143;
  assign n36145 = pi609 & n36143;
  assign n36146 = ~pi609 & ~n36027;
  assign n36147 = pi1155 & ~n36146;
  assign n36148 = ~n36145 & n36147;
  assign n36149 = ~pi609 & n36143;
  assign n36150 = pi609 & ~n36027;
  assign n36151 = ~pi1155 & ~n36150;
  assign n36152 = ~n36149 & n36151;
  assign n36153 = ~n36148 & ~n36152;
  assign n36154 = pi785 & ~n36153;
  assign n36155 = ~n36144 & ~n36154;
  assign n36156 = ~pi781 & ~n36155;
  assign n36157 = pi618 & n36155;
  assign n36158 = ~pi618 & ~n36027;
  assign n36159 = pi1154 & ~n36158;
  assign n36160 = ~n36157 & n36159;
  assign n36161 = ~pi618 & n36155;
  assign n36162 = pi618 & ~n36027;
  assign n36163 = ~pi1154 & ~n36162;
  assign n36164 = ~n36161 & n36163;
  assign n36165 = ~n36160 & ~n36164;
  assign n36166 = pi781 & ~n36165;
  assign n36167 = ~n36156 & ~n36166;
  assign n36168 = ~pi789 & ~n36167;
  assign n36169 = pi619 & n36167;
  assign n36170 = ~pi619 & ~n36027;
  assign n36171 = pi1159 & ~n36170;
  assign n36172 = ~n36169 & n36171;
  assign n36173 = ~pi619 & n36167;
  assign n36174 = pi619 & ~n36027;
  assign n36175 = ~pi1159 & ~n36174;
  assign n36176 = ~n36173 & n36175;
  assign n36177 = ~n36172 & ~n36176;
  assign n36178 = pi789 & ~n36177;
  assign n36179 = ~n36168 & ~n36178;
  assign n36180 = ~n17816 & n36179;
  assign n36181 = ~n36028 & ~n36180;
  assign n36182 = ~n20409 & n36181;
  assign n36183 = ~n19126 & ~n36027;
  assign n36184 = ~pi222 & ~n17054;
  assign n36185 = pi661 & pi680;
  assign n36186 = n17054 & ~n36185;
  assign n36187 = pi222 & n17074;
  assign n36188 = pi299 & ~n36187;
  assign n36189 = ~n36186 & n36188;
  assign n36190 = ~n36184 & n36189;
  assign n36191 = ~pi222 & ~n17049;
  assign n36192 = n17049 & ~n36185;
  assign n36193 = pi222 & n17068;
  assign n36194 = ~pi299 & ~n36193;
  assign n36195 = ~n36192 & n36194;
  assign n36196 = ~n36191 & n36195;
  assign n36197 = ~pi39 & ~n36196;
  assign n36198 = ~n36190 & n36197;
  assign n36199 = pi661 & ~n17338;
  assign n36200 = ~pi661 & ~n17172;
  assign n36201 = ~n36199 & ~n36200;
  assign n36202 = n6215 & n36201;
  assign n36203 = ~pi661 & ~n16812;
  assign n36204 = n16652 & ~n16785;
  assign n36205 = pi661 & ~n36204;
  assign n36206 = ~n36203 & ~n36205;
  assign n36207 = ~n6215 & n36206;
  assign n36208 = pi222 & ~n36207;
  assign n36209 = ~n36202 & n36208;
  assign n36210 = pi661 & n17298;
  assign n36211 = ~n6215 & n36210;
  assign n36212 = ~n17303 & n36185;
  assign n36213 = n6215 & n36212;
  assign n36214 = pi224 & ~n36213;
  assign n36215 = ~n36211 & n36214;
  assign n36216 = pi661 & n17323;
  assign n36217 = ~pi224 & ~n36216;
  assign n36218 = ~pi222 & ~n36217;
  assign n36219 = ~n36215 & n36218;
  assign n36220 = ~pi223 & ~n36219;
  assign n36221 = ~n36209 & n36220;
  assign n36222 = ~pi661 & ~n17151;
  assign n36223 = ~n16576 & ~n17356;
  assign n36224 = pi661 & ~n36223;
  assign n36225 = ~n36222 & ~n36224;
  assign n36226 = n6215 & n36225;
  assign n36227 = n16511 & n17127;
  assign n36228 = ~pi661 & n17122;
  assign n36229 = pi661 & ~n17358;
  assign n36230 = ~n36228 & ~n36229;
  assign n36231 = ~n36227 & n36230;
  assign n36232 = ~n6215 & n36231;
  assign n36233 = pi222 & ~n36232;
  assign n36234 = ~n36226 & n36233;
  assign n36235 = ~pi222 & pi661;
  assign n36236 = n17314 & n36235;
  assign n36237 = pi223 & ~n36236;
  assign n36238 = ~n36234 & n36237;
  assign n36239 = ~n36221 & ~n36238;
  assign n36240 = ~pi299 & ~n36239;
  assign n36241 = n6189 & n36201;
  assign n36242 = ~n6189 & n36206;
  assign n36243 = pi222 & ~n36242;
  assign n36244 = ~n36241 & n36243;
  assign n36245 = n6189 & ~n36212;
  assign n36246 = ~n6189 & ~n36210;
  assign n36247 = ~pi222 & ~n36246;
  assign n36248 = ~n36245 & n36247;
  assign n36249 = ~n3329 & ~n36248;
  assign n36250 = ~n36244 & n36249;
  assign n36251 = n36111 & ~n36216;
  assign n36252 = ~pi215 & ~n36251;
  assign n36253 = ~n36250 & n36252;
  assign n36254 = n17327 & n36235;
  assign n36255 = n6189 & n36225;
  assign n36256 = ~n6189 & n36231;
  assign n36257 = pi222 & ~n36256;
  assign n36258 = ~n36255 & n36257;
  assign n36259 = ~n36254 & ~n36258;
  assign n36260 = pi215 & ~n36259;
  assign n36261 = pi299 & ~n36260;
  assign n36262 = ~n36253 & n36261;
  assign n36263 = ~n36240 & ~n36262;
  assign n36264 = pi39 & ~n36263;
  assign n36265 = ~n36198 & ~n36264;
  assign n36266 = ~pi38 & ~n36265;
  assign n36267 = pi661 & n17391;
  assign n36268 = n36135 & ~n36267;
  assign n36269 = n3267 & ~n36268;
  assign n36270 = ~n36266 & n36269;
  assign n36271 = ~n36029 & ~n36270;
  assign n36272 = ~pi778 & ~n36271;
  assign n36273 = pi625 & n36271;
  assign n36274 = ~pi625 & ~n36027;
  assign n36275 = pi1153 & ~n36274;
  assign n36276 = ~n36273 & n36275;
  assign n36277 = ~pi625 & n36271;
  assign n36278 = pi625 & ~n36027;
  assign n36279 = ~pi1153 & ~n36278;
  assign n36280 = ~n36277 & n36279;
  assign n36281 = ~n36276 & ~n36280;
  assign n36282 = pi778 & ~n36281;
  assign n36283 = ~n36272 & ~n36282;
  assign n36284 = ~n17466 & ~n36283;
  assign n36285 = n17466 & n36027;
  assign n36286 = ~n36284 & ~n36285;
  assign n36287 = ~n17503 & ~n36286;
  assign n36288 = n17503 & n36027;
  assign n36289 = ~n36287 & ~n36288;
  assign n36290 = ~n17539 & n36289;
  assign n36291 = ~n17582 & n36290;
  assign n36292 = ~n36183 & ~n36291;
  assign n36293 = ~pi628 & ~n36292;
  assign n36294 = pi628 & ~n36027;
  assign n36295 = n17608 & ~n36294;
  assign n36296 = ~n36293 & n36295;
  assign n36297 = pi628 & ~n36292;
  assign n36298 = ~pi628 & ~n36027;
  assign n36299 = n17607 & ~n36298;
  assign n36300 = ~n36297 & n36299;
  assign n36301 = ~n36296 & ~n36300;
  assign n36302 = ~n36182 & n36301;
  assign n36303 = pi792 & ~n36302;
  assign n36304 = ~pi680 & n36032;
  assign n36305 = n6162 & n16639;
  assign n36306 = ~n16547 & ~n36305;
  assign n36307 = ~n16805 & n36306;
  assign n36308 = pi642 & ~n36307;
  assign n36309 = ~pi603 & n36306;
  assign n36310 = pi603 & n16619;
  assign n36311 = pi603 & n16522;
  assign n36312 = ~n36310 & ~n36311;
  assign n36313 = ~n36309 & n36312;
  assign n36314 = ~pi642 & n36313;
  assign n36315 = n6156 & ~n36314;
  assign n36316 = ~n36308 & n36315;
  assign n36317 = n16744 & n36307;
  assign n36318 = n16818 & ~n36306;
  assign n36319 = pi616 & ~n36318;
  assign n36320 = pi680 & ~n36319;
  assign n36321 = ~n36317 & n36320;
  assign n36322 = ~n36316 & n36321;
  assign n36323 = pi661 & ~n36322;
  assign n36324 = ~n36304 & n36323;
  assign n36325 = ~pi661 & pi681;
  assign n36326 = ~n36032 & n36325;
  assign n36327 = ~n36039 & ~n36326;
  assign n36328 = ~n36324 & n36327;
  assign n36329 = ~n6189 & ~n36328;
  assign n36330 = pi616 & ~n16891;
  assign n36331 = pi680 & ~n36330;
  assign n36332 = ~n16629 & n36331;
  assign n36333 = ~pi680 & n36043;
  assign n36334 = pi661 & ~n36333;
  assign n36335 = ~n36332 & n36334;
  assign n36336 = ~n36043 & n36325;
  assign n36337 = ~n36049 & ~n36336;
  assign n36338 = ~n36335 & n36337;
  assign n36339 = n6189 & ~n36338;
  assign n36340 = pi222 & ~n36339;
  assign n36341 = ~n36329 & n36340;
  assign n36342 = ~pi680 & n36054;
  assign n36343 = pi661 & ~n36342;
  assign n36344 = ~n16706 & ~n36054;
  assign n36345 = pi680 & ~n36344;
  assign n36346 = n36343 & ~n36345;
  assign n36347 = ~n36054 & n36325;
  assign n36348 = ~n36060 & ~n36347;
  assign n36349 = ~n36346 & n36348;
  assign n36350 = ~n6189 & n36349;
  assign n36351 = pi616 & ~n16819;
  assign n36352 = pi680 & ~n16729;
  assign n36353 = ~n36351 & n36352;
  assign n36354 = ~pi680 & n36069;
  assign n36355 = pi661 & ~n36354;
  assign n36356 = ~n36353 & n36355;
  assign n36357 = n16642 & n36057;
  assign n36358 = ~n6158 & n36069;
  assign n36359 = n16511 & ~n36358;
  assign n36360 = ~n36357 & n36359;
  assign n36361 = ~n36069 & n36325;
  assign n36362 = ~n36360 & ~n36361;
  assign n36363 = ~n36356 & n36362;
  assign n36364 = n6189 & n36363;
  assign n36365 = ~pi222 & ~n36364;
  assign n36366 = ~n36350 & n36365;
  assign n36367 = ~n36341 & ~n36366;
  assign n36368 = ~n3329 & ~n36367;
  assign n36369 = ~n36030 & ~n36185;
  assign n36370 = ~pi616 & ~n16714;
  assign n36371 = ~n36351 & ~n36370;
  assign n36372 = ~n36369 & n36371;
  assign n36373 = n36111 & ~n36372;
  assign n36374 = ~pi215 & ~n36373;
  assign n36375 = ~n36368 & n36374;
  assign n36376 = ~pi680 & n36084;
  assign n36377 = ~n16589 & n16818;
  assign n36378 = pi616 & ~n36377;
  assign n36379 = pi680 & ~n36378;
  assign n36380 = n16594 & n36379;
  assign n36381 = pi661 & ~n36380;
  assign n36382 = ~n36376 & n36381;
  assign n36383 = ~n36084 & n36325;
  assign n36384 = ~n36087 & ~n36383;
  assign n36385 = ~n36382 & n36384;
  assign n36386 = ~n6189 & ~n36385;
  assign n36387 = ~n16562 & n36331;
  assign n36388 = ~pi680 & n36075;
  assign n36389 = pi661 & ~n36388;
  assign n36390 = ~n36387 & n36389;
  assign n36391 = ~n36075 & n36325;
  assign n36392 = ~n36080 & ~n36391;
  assign n36393 = ~n36390 & n36392;
  assign n36394 = n6189 & ~n36393;
  assign n36395 = pi222 & ~n36394;
  assign n36396 = ~n36386 & n36395;
  assign n36397 = ~n16588 & ~n16857;
  assign n36398 = pi616 & n36397;
  assign n36399 = pi680 & ~n36398;
  assign n36400 = n16754 & n36399;
  assign n36401 = pi616 & n16588;
  assign n36402 = ~pi680 & n36401;
  assign n36403 = pi661 & ~n36402;
  assign n36404 = ~n36400 & n36403;
  assign n36405 = ~pi661 & ~n36401;
  assign n36406 = ~n16542 & n36069;
  assign n36407 = n6160 & ~n36406;
  assign n36408 = ~n36405 & ~n36407;
  assign n36409 = ~n36404 & n36408;
  assign n36410 = ~n6189 & n36409;
  assign n36411 = n16765 & n36185;
  assign n36412 = ~n36093 & ~n36411;
  assign n36413 = n6189 & ~n36412;
  assign n36414 = ~pi222 & ~n36413;
  assign n36415 = ~n36410 & n36414;
  assign n36416 = pi215 & ~n36415;
  assign n36417 = ~n36396 & n36416;
  assign n36418 = pi299 & ~n36417;
  assign n36419 = ~n36375 & n36418;
  assign n36420 = n36185 & ~n36371;
  assign n36421 = ~n36069 & ~n36185;
  assign n36422 = ~pi222 & ~n36421;
  assign n36423 = ~n36420 & n36422;
  assign n36424 = ~n3306 & ~n36423;
  assign n36425 = ~n6215 & n36349;
  assign n36426 = n6215 & n36363;
  assign n36427 = pi224 & ~n36426;
  assign n36428 = ~n36425 & n36427;
  assign n36429 = ~n36424 & ~n36428;
  assign n36430 = ~n6215 & n36328;
  assign n36431 = n6215 & n36338;
  assign n36432 = pi222 & ~n36431;
  assign n36433 = ~n36430 & n36432;
  assign n36434 = ~n36429 & ~n36433;
  assign n36435 = ~pi223 & ~n36434;
  assign n36436 = ~n6215 & ~n36385;
  assign n36437 = n6215 & ~n36393;
  assign n36438 = pi222 & ~n36437;
  assign n36439 = ~n36436 & n36438;
  assign n36440 = ~n6215 & n36409;
  assign n36441 = n6215 & ~n36412;
  assign n36442 = ~pi222 & ~n36441;
  assign n36443 = ~n36440 & n36442;
  assign n36444 = pi223 & ~n36443;
  assign n36445 = ~n36439 & n36444;
  assign n36446 = ~pi299 & ~n36445;
  assign n36447 = ~n36435 & n36446;
  assign n36448 = pi39 & ~n36447;
  assign n36449 = ~n36419 & n36448;
  assign n36450 = n18457 & ~n36185;
  assign n36451 = ~pi616 & n17084;
  assign n36452 = ~n17019 & n17074;
  assign n36453 = ~n36451 & ~n36452;
  assign n36454 = ~n36450 & n36453;
  assign n36455 = pi222 & ~n36454;
  assign n36456 = pi661 & n18458;
  assign n36457 = pi616 & n17084;
  assign n36458 = ~pi222 & ~n36457;
  assign n36459 = ~n36456 & n36458;
  assign n36460 = ~n36455 & ~n36459;
  assign n36461 = pi299 & ~n36460;
  assign n36462 = pi661 & n18448;
  assign n36463 = pi616 & n17079;
  assign n36464 = ~pi222 & ~n36463;
  assign n36465 = ~n36462 & n36464;
  assign n36466 = n18447 & ~n36185;
  assign n36467 = ~pi616 & n17079;
  assign n36468 = ~n16658 & n17068;
  assign n36469 = ~n36467 & ~n36468;
  assign n36470 = ~n36466 & n36469;
  assign n36471 = pi222 & ~n36470;
  assign n36472 = ~n36465 & ~n36471;
  assign n36473 = ~pi299 & ~n36472;
  assign n36474 = ~pi39 & ~n36473;
  assign n36475 = ~n36461 & n36474;
  assign n36476 = ~pi38 & ~n36475;
  assign n36477 = ~n36449 & n36476;
  assign n36478 = n16529 & n16818;
  assign n36479 = ~pi222 & ~pi616;
  assign n36480 = ~pi39 & pi616;
  assign n36481 = n36185 & n36480;
  assign n36482 = ~n36479 & ~n36481;
  assign n36483 = n36478 & ~n36482;
  assign n36484 = ~pi616 & ~n16667;
  assign n36485 = ~n36369 & ~n36484;
  assign n36486 = n17280 & n36485;
  assign n36487 = ~n36134 & ~n36486;
  assign n36488 = ~n36483 & ~n36487;
  assign n36489 = pi38 & ~n36488;
  assign n36490 = n3267 & ~n36489;
  assign n36491 = ~n36477 & n36490;
  assign n36492 = ~n36029 & ~n36491;
  assign n36493 = ~pi625 & n36492;
  assign n36494 = pi625 & n36140;
  assign n36495 = ~pi1153 & ~n36494;
  assign n36496 = ~n36493 & n36495;
  assign n36497 = ~pi608 & ~n36276;
  assign n36498 = ~n36496 & n36497;
  assign n36499 = pi625 & n36492;
  assign n36500 = ~pi625 & n36140;
  assign n36501 = pi1153 & ~n36500;
  assign n36502 = ~n36499 & n36501;
  assign n36503 = pi608 & ~n36280;
  assign n36504 = ~n36502 & n36503;
  assign n36505 = ~n36498 & ~n36504;
  assign n36506 = pi778 & ~n36505;
  assign n36507 = ~pi778 & n36492;
  assign n36508 = ~n36506 & ~n36507;
  assign n36509 = ~pi609 & ~n36508;
  assign n36510 = pi609 & n36283;
  assign n36511 = ~pi1155 & ~n36510;
  assign n36512 = ~n36509 & n36511;
  assign n36513 = ~pi660 & ~n36148;
  assign n36514 = ~n36512 & n36513;
  assign n36515 = pi609 & ~n36508;
  assign n36516 = ~pi609 & n36283;
  assign n36517 = pi1155 & ~n36516;
  assign n36518 = ~n36515 & n36517;
  assign n36519 = pi660 & ~n36152;
  assign n36520 = ~n36518 & n36519;
  assign n36521 = ~n36514 & ~n36520;
  assign n36522 = pi785 & ~n36521;
  assign n36523 = ~pi785 & ~n36508;
  assign n36524 = ~n36522 & ~n36523;
  assign n36525 = ~pi618 & ~n36524;
  assign n36526 = pi618 & n36286;
  assign n36527 = ~pi1154 & ~n36526;
  assign n36528 = ~n36525 & n36527;
  assign n36529 = ~pi627 & ~n36160;
  assign n36530 = ~n36528 & n36529;
  assign n36531 = pi618 & ~n36524;
  assign n36532 = ~pi618 & n36286;
  assign n36533 = pi1154 & ~n36532;
  assign n36534 = ~n36531 & n36533;
  assign n36535 = pi627 & ~n36164;
  assign n36536 = ~n36534 & n36535;
  assign n36537 = ~n36530 & ~n36536;
  assign n36538 = pi781 & ~n36537;
  assign n36539 = ~pi781 & ~n36524;
  assign n36540 = ~n36538 & ~n36539;
  assign n36541 = pi619 & ~n36540;
  assign n36542 = ~pi619 & n36289;
  assign n36543 = pi1159 & ~n36542;
  assign n36544 = ~n36541 & n36543;
  assign n36545 = pi648 & ~n36176;
  assign n36546 = ~n36544 & n36545;
  assign n36547 = ~pi619 & ~n36540;
  assign n36548 = pi619 & n36289;
  assign n36549 = ~pi1159 & ~n36548;
  assign n36550 = ~n36547 & n36549;
  assign n36551 = ~pi648 & ~n36172;
  assign n36552 = ~n36550 & n36551;
  assign n36553 = pi789 & ~n36552;
  assign n36554 = ~n36546 & n36553;
  assign n36555 = ~pi789 & n36540;
  assign n36556 = pi626 & n36179;
  assign n36557 = ~pi626 & ~n36027;
  assign n36558 = n17579 & ~n36557;
  assign n36559 = ~n36556 & n36558;
  assign n36560 = ~pi626 & n36179;
  assign n36561 = pi626 & ~n36027;
  assign n36562 = n17580 & ~n36561;
  assign n36563 = ~n36560 & n36562;
  assign n36564 = n17539 & ~n36027;
  assign n36565 = n17704 & ~n36564;
  assign n36566 = ~n36290 & n36565;
  assign n36567 = ~n36563 & ~n36566;
  assign n36568 = ~n36559 & n36567;
  assign n36569 = pi788 & ~n36568;
  assign n36570 = ~n36555 & ~n36569;
  assign n36571 = ~n36554 & n36570;
  assign n36572 = ~n17817 & n36568;
  assign n36573 = ~n20205 & ~n36572;
  assign n36574 = ~n36571 & n36573;
  assign n36575 = ~n36303 & ~n36574;
  assign n36576 = n20207 & ~n36575;
  assign n36577 = ~n17610 & n36181;
  assign n36578 = n17610 & n36027;
  assign n36579 = ~n36577 & ~n36578;
  assign n36580 = ~n20398 & ~n36579;
  assign n36581 = ~n19158 & ~n36292;
  assign n36582 = n17858 & ~n36027;
  assign n36583 = ~n36581 & ~n36582;
  assign n36584 = pi647 & ~n36583;
  assign n36585 = ~pi647 & ~n36027;
  assign n36586 = pi1157 & ~n36585;
  assign n36587 = ~n36584 & n36586;
  assign n36588 = ~pi630 & n36587;
  assign n36589 = ~pi647 & ~n36583;
  assign n36590 = pi647 & ~n36027;
  assign n36591 = ~pi1157 & ~n36590;
  assign n36592 = ~n36589 & n36591;
  assign n36593 = pi630 & n36592;
  assign n36594 = ~n36588 & ~n36593;
  assign n36595 = ~n36580 & n36594;
  assign n36596 = pi787 & ~n36595;
  assign n36597 = ~n36576 & ~n36596;
  assign n36598 = pi644 & n36597;
  assign n36599 = ~pi787 & n36583;
  assign n36600 = ~n36587 & ~n36592;
  assign n36601 = pi787 & ~n36600;
  assign n36602 = ~n36599 & ~n36601;
  assign n36603 = ~pi644 & n36602;
  assign n36604 = pi715 & ~n36603;
  assign n36605 = ~n36598 & n36604;
  assign n36606 = n17652 & ~n36027;
  assign n36607 = ~n17652 & n36579;
  assign n36608 = ~n36606 & ~n36607;
  assign n36609 = pi644 & ~n36608;
  assign n36610 = ~pi644 & ~n36027;
  assign n36611 = ~pi715 & ~n36610;
  assign n36612 = ~n36609 & n36611;
  assign n36613 = pi1160 & ~n36612;
  assign n36614 = ~n36605 & n36613;
  assign n36615 = ~pi644 & n36597;
  assign n36616 = pi644 & n36602;
  assign n36617 = ~pi715 & ~n36616;
  assign n36618 = ~n36615 & n36617;
  assign n36619 = ~pi644 & ~n36608;
  assign n36620 = pi644 & ~n36027;
  assign n36621 = pi715 & ~n36620;
  assign n36622 = ~n36619 & n36621;
  assign n36623 = ~pi1160 & ~n36622;
  assign n36624 = ~n36618 & n36623;
  assign n36625 = ~n36614 & ~n36624;
  assign n36626 = pi790 & ~n36625;
  assign n36627 = ~pi790 & n36597;
  assign n36628 = ~n36626 & ~n36627;
  assign n36629 = ~po1038 & ~n36628;
  assign n36630 = ~pi222 & po1038;
  assign po379 = ~n36629 & ~n36630;
  assign n36632 = ~pi299 & ~n17153;
  assign n36633 = pi39 & ~n36632;
  assign n36634 = ~n17198 & n36633;
  assign n36635 = n14755 & ~n17954;
  assign n36636 = ~n36634 & n36635;
  assign n36637 = n18723 & ~n36636;
  assign n36638 = pi223 & ~n36637;
  assign n36639 = n17816 & ~n36638;
  assign n36640 = n17438 & ~n36638;
  assign n36641 = pi223 & ~n3267;
  assign n36642 = pi642 & n16521;
  assign n36643 = n35656 & ~n36642;
  assign n36644 = pi642 & ~n16713;
  assign n36645 = n6156 & ~n36644;
  assign n36646 = ~n16632 & n36645;
  assign n36647 = ~n36643 & ~n36646;
  assign n36648 = pi681 & n36647;
  assign n36649 = ~n6159 & ~n36647;
  assign n36650 = ~n17204 & ~n35654;
  assign n36651 = n6159 & ~n36650;
  assign n36652 = ~pi681 & ~n36651;
  assign n36653 = ~n36649 & n36652;
  assign n36654 = n6189 & ~n36653;
  assign n36655 = ~n36648 & n36654;
  assign n36656 = pi642 & ~n16692;
  assign n36657 = ~pi642 & ~n16652;
  assign n36658 = ~n36656 & ~n36657;
  assign n36659 = pi681 & ~n36658;
  assign n36660 = ~n6159 & n36658;
  assign n36661 = n6159 & ~n16619;
  assign n36662 = ~n36642 & n36661;
  assign n36663 = ~pi681 & ~n36662;
  assign n36664 = ~n36660 & n36663;
  assign n36665 = ~n6189 & ~n36664;
  assign n36666 = ~n36659 & n36665;
  assign n36667 = pi223 & ~n36666;
  assign n36668 = ~n36655 & n36667;
  assign n36669 = n35703 & n36642;
  assign n36670 = ~n20739 & n36669;
  assign n36671 = pi642 & ~n36064;
  assign n36672 = n20739 & n36671;
  assign n36673 = ~pi947 & ~n36672;
  assign n36674 = ~n36670 & n36673;
  assign n36675 = pi947 & ~n36669;
  assign n36676 = ~pi223 & ~n36675;
  assign n36677 = ~n36674 & n36676;
  assign n36678 = ~n3329 & ~n36677;
  assign n36679 = ~n36668 & n36678;
  assign n36680 = pi642 & n16543;
  assign n36681 = pi223 & ~n16518;
  assign n36682 = n3329 & ~n36681;
  assign n36683 = ~n36680 & n36682;
  assign n36684 = ~pi215 & ~n36683;
  assign n36685 = ~n36679 & n36684;
  assign n36686 = ~n6159 & n36680;
  assign n36687 = ~pi681 & ~n36686;
  assign n36688 = pi642 & n6159;
  assign n36689 = n16551 & n36688;
  assign n36690 = n36687 & ~n36689;
  assign n36691 = pi642 & ~n16740;
  assign n36692 = n6159 & ~n36691;
  assign n36693 = ~n16542 & n36692;
  assign n36694 = ~pi681 & ~n36693;
  assign n36695 = n16583 & n36694;
  assign n36696 = ~n36690 & ~n36695;
  assign n36697 = pi642 & n16588;
  assign n36698 = pi681 & ~n36697;
  assign n36699 = n36696 & ~n36698;
  assign n36700 = ~n20739 & n36699;
  assign n36701 = n6189 & ~n36690;
  assign n36702 = n36680 & n36701;
  assign n36703 = ~pi947 & ~n36702;
  assign n36704 = ~n36700 & n36703;
  assign n36705 = pi947 & ~n36699;
  assign n36706 = ~pi223 & ~n36705;
  assign n36707 = ~n36704 & n36706;
  assign n36708 = n16575 & ~n36680;
  assign n36709 = pi681 & ~n36708;
  assign n36710 = ~n6159 & n36708;
  assign n36711 = n16768 & ~n36642;
  assign n36712 = ~pi681 & ~n36711;
  assign n36713 = ~n36710 & n36712;
  assign n36714 = ~n36709 & ~n36713;
  assign n36715 = n6189 & n36714;
  assign n36716 = ~pi642 & n16585;
  assign n36717 = pi642 & ~n16741;
  assign n36718 = ~n36716 & ~n36717;
  assign n36719 = ~n6159 & n36718;
  assign n36720 = n36694 & ~n36719;
  assign n36721 = pi681 & ~n36718;
  assign n36722 = ~n36720 & ~n36721;
  assign n36723 = ~n6189 & n36722;
  assign n36724 = pi223 & ~n36723;
  assign n36725 = ~n36715 & n36724;
  assign n36726 = ~n36707 & ~n36725;
  assign n36727 = pi215 & ~n36726;
  assign n36728 = pi299 & ~n36727;
  assign n36729 = ~n36685 & n36728;
  assign n36730 = ~n6215 & n36669;
  assign n36731 = n6215 & n36671;
  assign n36732 = ~n3052 & ~n36731;
  assign n36733 = ~n36730 & n36732;
  assign n36734 = n3052 & ~n36680;
  assign n36735 = ~pi223 & ~n36734;
  assign n36736 = ~n36733 & n36735;
  assign n36737 = n6215 & n36714;
  assign n36738 = ~n6215 & n36722;
  assign n36739 = pi223 & ~n36738;
  assign n36740 = ~n36737 & n36739;
  assign n36741 = ~pi299 & ~n36740;
  assign n36742 = ~n36736 & n36741;
  assign n36743 = pi39 & ~n36742;
  assign n36744 = ~n36729 & n36743;
  assign n36745 = ~pi223 & pi642;
  assign n36746 = n17079 & n36745;
  assign n36747 = ~pi299 & ~n36746;
  assign n36748 = ~pi642 & n17079;
  assign n36749 = pi223 & ~n36748;
  assign n36750 = n17040 & n36749;
  assign n36751 = n36747 & ~n36750;
  assign n36752 = n17084 & n36745;
  assign n36753 = pi299 & ~n36752;
  assign n36754 = n6155 & n17083;
  assign n36755 = pi223 & ~n36754;
  assign n36756 = ~n17027 & n36755;
  assign n36757 = n36753 & ~n36756;
  assign n36758 = ~pi39 & ~n36757;
  assign n36759 = ~n36751 & n36758;
  assign n36760 = ~pi38 & ~n36759;
  assign n36761 = ~n36744 & n36760;
  assign n36762 = pi39 & pi223;
  assign n36763 = pi38 & ~n36762;
  assign n36764 = n16529 & ~n36642;
  assign n36765 = ~pi223 & ~n16529;
  assign n36766 = ~pi39 & ~n36765;
  assign n36767 = ~n36764 & n36766;
  assign n36768 = n36763 & ~n36767;
  assign n36769 = n3267 & ~n36768;
  assign n36770 = ~n36761 & n36769;
  assign n36771 = ~n36641 & ~n36770;
  assign n36772 = ~n17438 & n36771;
  assign n36773 = ~n36640 & ~n36772;
  assign n36774 = ~pi785 & n36773;
  assign n36775 = pi609 & ~n36773;
  assign n36776 = ~pi609 & ~n36638;
  assign n36777 = pi1155 & ~n36776;
  assign n36778 = ~n36775 & n36777;
  assign n36779 = ~pi609 & ~n36773;
  assign n36780 = pi609 & ~n36638;
  assign n36781 = ~pi1155 & ~n36780;
  assign n36782 = ~n36779 & n36781;
  assign n36783 = ~n36778 & ~n36782;
  assign n36784 = pi785 & ~n36783;
  assign n36785 = ~n36774 & ~n36784;
  assign n36786 = ~pi781 & ~n36785;
  assign n36787 = pi618 & n36785;
  assign n36788 = ~pi618 & ~n36638;
  assign n36789 = pi1154 & ~n36788;
  assign n36790 = ~n36787 & n36789;
  assign n36791 = ~pi618 & n36785;
  assign n36792 = pi618 & ~n36638;
  assign n36793 = ~pi1154 & ~n36792;
  assign n36794 = ~n36791 & n36793;
  assign n36795 = ~n36790 & ~n36794;
  assign n36796 = pi781 & ~n36795;
  assign n36797 = ~n36786 & ~n36796;
  assign n36798 = ~pi789 & ~n36797;
  assign n36799 = pi619 & n36797;
  assign n36800 = ~pi619 & ~n36638;
  assign n36801 = pi1159 & ~n36800;
  assign n36802 = ~n36799 & n36801;
  assign n36803 = ~pi619 & n36797;
  assign n36804 = pi619 & ~n36638;
  assign n36805 = ~pi1159 & ~n36804;
  assign n36806 = ~n36803 & n36805;
  assign n36807 = ~n36802 & ~n36806;
  assign n36808 = pi789 & ~n36807;
  assign n36809 = ~n36798 & ~n36808;
  assign n36810 = ~n17816 & n36809;
  assign n36811 = ~n36639 & ~n36810;
  assign n36812 = ~n17610 & n36811;
  assign n36813 = n17610 & n36638;
  assign n36814 = ~n36812 & ~n36813;
  assign n36815 = ~n20398 & ~n36814;
  assign n36816 = ~n19126 & ~n36638;
  assign n36817 = n17466 & ~n36638;
  assign n36818 = ~pi223 & ~n17054;
  assign n36819 = pi680 & pi681;
  assign n36820 = n17054 & ~n36819;
  assign n36821 = pi223 & n17074;
  assign n36822 = pi299 & ~n36821;
  assign n36823 = ~n36820 & n36822;
  assign n36824 = ~n36818 & n36823;
  assign n36825 = ~pi223 & ~n17049;
  assign n36826 = n17049 & ~n36819;
  assign n36827 = pi223 & n17068;
  assign n36828 = ~pi299 & ~n36827;
  assign n36829 = ~n36826 & n36828;
  assign n36830 = ~n36825 & n36829;
  assign n36831 = ~pi39 & ~n36830;
  assign n36832 = ~n36824 & n36831;
  assign n36833 = pi681 & n17323;
  assign n36834 = n36682 & ~n36833;
  assign n36835 = pi681 & ~n17338;
  assign n36836 = n6189 & ~n17171;
  assign n36837 = ~n36835 & n36836;
  assign n36838 = pi681 & n17298;
  assign n36839 = ~n6189 & ~n36838;
  assign n36840 = n16812 & n36839;
  assign n36841 = pi223 & ~n36840;
  assign n36842 = ~n36837 & n36841;
  assign n36843 = ~n17303 & n36819;
  assign n36844 = n6189 & ~n36843;
  assign n36845 = ~pi223 & ~n36839;
  assign n36846 = ~n36844 & n36845;
  assign n36847 = ~n3329 & ~n36846;
  assign n36848 = ~n36842 & n36847;
  assign n36849 = ~n36834 & ~n36848;
  assign n36850 = ~pi215 & ~n36849;
  assign n36851 = pi681 & ~n17358;
  assign n36852 = ~n17131 & ~n36851;
  assign n36853 = ~n6189 & n36852;
  assign n36854 = pi681 & ~n36223;
  assign n36855 = ~n17150 & ~n36854;
  assign n36856 = n6189 & n36855;
  assign n36857 = pi223 & ~n36856;
  assign n36858 = ~n36853 & n36857;
  assign n36859 = ~pi223 & pi681;
  assign n36860 = n17327 & n36859;
  assign n36861 = pi215 & ~n36860;
  assign n36862 = ~n36858 & n36861;
  assign n36863 = pi299 & ~n36862;
  assign n36864 = ~n36850 & n36863;
  assign n36865 = n3052 & ~n36833;
  assign n36866 = ~n6215 & n36838;
  assign n36867 = n6215 & n36843;
  assign n36868 = ~n3052 & ~n36867;
  assign n36869 = ~n36866 & n36868;
  assign n36870 = ~n36865 & ~n36869;
  assign n36871 = ~pi223 & ~n36870;
  assign n36872 = ~n6215 & ~n36852;
  assign n36873 = n6215 & ~n36855;
  assign n36874 = pi223 & ~n36873;
  assign n36875 = ~n36872 & n36874;
  assign n36876 = ~pi299 & ~n36875;
  assign n36877 = ~n36871 & n36876;
  assign n36878 = pi39 & ~n36877;
  assign n36879 = ~n36864 & n36878;
  assign n36880 = ~n36832 & ~n36879;
  assign n36881 = ~pi38 & ~n36880;
  assign n36882 = pi223 & ~n17280;
  assign n36883 = pi681 & n17391;
  assign n36884 = pi38 & ~n36883;
  assign n36885 = ~n36882 & n36884;
  assign n36886 = n3267 & ~n36885;
  assign n36887 = ~n36881 & n36886;
  assign n36888 = ~n36641 & ~n36887;
  assign n36889 = ~pi778 & ~n36888;
  assign n36890 = pi625 & n36888;
  assign n36891 = ~pi625 & ~n36638;
  assign n36892 = pi1153 & ~n36891;
  assign n36893 = ~n36890 & n36892;
  assign n36894 = ~pi625 & n36888;
  assign n36895 = pi625 & ~n36638;
  assign n36896 = ~pi1153 & ~n36895;
  assign n36897 = ~n36894 & n36896;
  assign n36898 = ~n36893 & ~n36897;
  assign n36899 = pi778 & ~n36898;
  assign n36900 = ~n36889 & ~n36899;
  assign n36901 = ~n17466 & n36900;
  assign n36902 = ~n36817 & ~n36901;
  assign n36903 = ~n17503 & n36902;
  assign n36904 = n17503 & n36638;
  assign n36905 = ~n36903 & ~n36904;
  assign n36906 = ~n17539 & n36905;
  assign n36907 = ~n17582 & n36906;
  assign n36908 = ~n36816 & ~n36907;
  assign n36909 = ~n19158 & ~n36908;
  assign n36910 = n17858 & ~n36638;
  assign n36911 = ~n36909 & ~n36910;
  assign n36912 = pi647 & ~n36911;
  assign n36913 = ~pi647 & ~n36638;
  assign n36914 = pi1157 & ~n36913;
  assign n36915 = ~n36912 & n36914;
  assign n36916 = ~pi630 & n36915;
  assign n36917 = ~pi647 & ~n36911;
  assign n36918 = pi647 & ~n36638;
  assign n36919 = ~pi1157 & ~n36918;
  assign n36920 = ~n36917 & n36919;
  assign n36921 = pi630 & n36920;
  assign n36922 = ~n36916 & ~n36921;
  assign n36923 = ~n36815 & n36922;
  assign n36924 = pi787 & ~n36923;
  assign n36925 = ~n20409 & n36811;
  assign n36926 = ~pi628 & ~n36908;
  assign n36927 = pi628 & ~n36638;
  assign n36928 = n17608 & ~n36927;
  assign n36929 = ~n36926 & n36928;
  assign n36930 = pi628 & ~n36908;
  assign n36931 = ~pi628 & ~n36638;
  assign n36932 = n17607 & ~n36931;
  assign n36933 = ~n36930 & n36932;
  assign n36934 = ~n36929 & ~n36933;
  assign n36935 = ~n36925 & n36934;
  assign n36936 = pi792 & ~n36935;
  assign n36937 = ~pi626 & ~n36809;
  assign n36938 = pi626 & n36638;
  assign n36939 = n17580 & ~n36938;
  assign n36940 = ~n36937 & n36939;
  assign n36941 = n17539 & ~n36638;
  assign n36942 = ~n36906 & ~n36941;
  assign n36943 = n17704 & ~n36942;
  assign n36944 = pi626 & ~n36809;
  assign n36945 = ~pi626 & n36638;
  assign n36946 = n17579 & ~n36945;
  assign n36947 = ~n36944 & n36946;
  assign n36948 = ~n36943 & ~n36947;
  assign n36949 = ~n36940 & n36948;
  assign n36950 = pi788 & ~n36949;
  assign n36951 = ~n16649 & n36642;
  assign n36952 = pi681 & ~n36951;
  assign n36953 = ~n36819 & ~n36952;
  assign n36954 = ~pi642 & ~n6156;
  assign n36955 = ~n16693 & n36954;
  assign n36956 = pi642 & n16806;
  assign n36957 = pi680 & ~n36956;
  assign n36958 = ~n16701 & n36957;
  assign n36959 = ~n36955 & n36958;
  assign n36960 = ~n36953 & ~n36959;
  assign n36961 = ~pi681 & ~n36669;
  assign n36962 = ~n36960 & ~n36961;
  assign n36963 = ~n6189 & ~n36962;
  assign n36964 = n16642 & n36688;
  assign n36965 = n36687 & ~n36964;
  assign n36966 = ~pi680 & ~n36680;
  assign n36967 = ~pi642 & ~n16522;
  assign n36968 = ~n16818 & ~n36967;
  assign n36969 = n35656 & n36968;
  assign n36970 = pi680 & ~n36969;
  assign n36971 = pi642 & ~n16819;
  assign n36972 = n6156 & ~n36971;
  assign n36973 = ~pi642 & ~n16725;
  assign n36974 = n36972 & ~n36973;
  assign n36975 = n36970 & ~n36974;
  assign n36976 = ~n36966 & ~n36975;
  assign n36977 = pi681 & ~n36976;
  assign n36978 = ~n36965 & ~n36977;
  assign n36979 = n6189 & ~n36978;
  assign n36980 = ~pi223 & ~n36979;
  assign n36981 = ~n36963 & n36980;
  assign n36982 = ~n36648 & ~n36819;
  assign n36983 = pi642 & ~n16891;
  assign n36984 = ~n16625 & ~n36983;
  assign n36985 = n6156 & ~n36984;
  assign n36986 = ~n6156 & ~n16518;
  assign n36987 = n36970 & ~n36986;
  assign n36988 = ~n36985 & n36987;
  assign n36989 = ~n36982 & ~n36988;
  assign n36990 = n36654 & ~n36989;
  assign n36991 = ~n36659 & ~n36819;
  assign n36992 = n36307 & n36954;
  assign n36993 = n16592 & ~n36313;
  assign n36994 = pi642 & ~n36318;
  assign n36995 = pi680 & ~n36994;
  assign n36996 = ~n36993 & n36995;
  assign n36997 = ~n36992 & n36996;
  assign n36998 = ~n36991 & ~n36997;
  assign n36999 = n36665 & ~n36998;
  assign n37000 = pi223 & ~n36999;
  assign n37001 = ~n36990 & n37000;
  assign n37002 = ~n3329 & ~n37001;
  assign n37003 = ~n36981 & n37002;
  assign n37004 = n36642 & ~n36819;
  assign n37005 = n36819 & ~n36967;
  assign n37006 = ~n36478 & n37005;
  assign n37007 = ~n37004 & ~n37006;
  assign n37008 = n16518 & ~n37007;
  assign n37009 = n36682 & ~n37008;
  assign n37010 = ~pi215 & ~n37009;
  assign n37011 = ~n37003 & n37010;
  assign n37012 = ~n36709 & ~n36819;
  assign n37013 = ~pi614 & n16558;
  assign n37014 = ~n36983 & ~n37013;
  assign n37015 = ~pi616 & ~n37014;
  assign n37016 = n36987 & ~n37015;
  assign n37017 = ~n37012 & ~n37016;
  assign n37018 = ~n36713 & ~n37017;
  assign n37019 = n6189 & ~n37018;
  assign n37020 = ~n6156 & n16590;
  assign n37021 = pi642 & ~n36377;
  assign n37022 = pi680 & ~n16593;
  assign n37023 = ~n37021 & n37022;
  assign n37024 = ~n37020 & n37023;
  assign n37025 = ~n36721 & ~n36819;
  assign n37026 = ~n37024 & ~n37025;
  assign n37027 = ~n36720 & ~n37026;
  assign n37028 = ~n6189 & ~n37027;
  assign n37029 = pi223 & ~n37028;
  assign n37030 = ~n37019 & n37029;
  assign n37031 = ~n36698 & ~n36819;
  assign n37032 = n16750 & n16857;
  assign n37033 = n16592 & ~n37032;
  assign n37034 = pi642 & n36397;
  assign n37035 = ~n16742 & n36954;
  assign n37036 = pi680 & ~n37035;
  assign n37037 = ~n37034 & n37036;
  assign n37038 = ~n37033 & n37037;
  assign n37039 = ~n37031 & ~n37038;
  assign n37040 = ~n6189 & n36696;
  assign n37041 = ~n37039 & n37040;
  assign n37042 = ~n16751 & n36972;
  assign n37043 = n36970 & ~n37042;
  assign n37044 = ~n36966 & ~n37043;
  assign n37045 = pi681 & ~n37044;
  assign n37046 = n36701 & ~n37045;
  assign n37047 = ~pi223 & ~n37046;
  assign n37048 = ~n37041 & n37047;
  assign n37049 = pi215 & ~n37048;
  assign n37050 = ~n37030 & n37049;
  assign n37051 = pi299 & ~n37050;
  assign n37052 = ~n37011 & n37051;
  assign n37053 = n6215 & n36978;
  assign n37054 = ~n6215 & n36962;
  assign n37055 = ~n3052 & ~n37054;
  assign n37056 = ~n37053 & n37055;
  assign n37057 = n3052 & ~n37008;
  assign n37058 = ~pi223 & ~n37057;
  assign n37059 = ~n37056 & n37058;
  assign n37060 = n6215 & n37018;
  assign n37061 = ~n6215 & n37027;
  assign n37062 = pi223 & ~n37061;
  assign n37063 = ~n37060 & n37062;
  assign n37064 = ~pi299 & ~n37063;
  assign n37065 = ~n37059 & n37064;
  assign n37066 = pi39 & ~n37065;
  assign n37067 = ~n37052 & n37066;
  assign n37068 = n18457 & ~n36819;
  assign n37069 = ~n36452 & n36755;
  assign n37070 = ~n37068 & n37069;
  assign n37071 = n18458 & n36859;
  assign n37072 = n36753 & ~n37071;
  assign n37073 = ~n37070 & n37072;
  assign n37074 = n18447 & ~n36819;
  assign n37075 = ~n36468 & n36749;
  assign n37076 = ~n37074 & n37075;
  assign n37077 = n18448 & n36859;
  assign n37078 = n36747 & ~n37077;
  assign n37079 = ~n37076 & n37078;
  assign n37080 = ~pi39 & ~n37079;
  assign n37081 = ~n37073 & n37080;
  assign n37082 = ~pi38 & ~n37081;
  assign n37083 = ~n37067 & n37082;
  assign n37084 = ~n36882 & n37007;
  assign n37085 = n36766 & ~n37084;
  assign n37086 = n36763 & ~n37085;
  assign n37087 = n3267 & ~n37086;
  assign n37088 = ~n37083 & n37087;
  assign n37089 = ~n36641 & ~n37088;
  assign n37090 = ~pi625 & n37089;
  assign n37091 = pi625 & n36771;
  assign n37092 = ~pi1153 & ~n37091;
  assign n37093 = ~n37090 & n37092;
  assign n37094 = ~pi608 & ~n37093;
  assign n37095 = ~n36893 & n37094;
  assign n37096 = pi625 & n37089;
  assign n37097 = ~pi625 & n36771;
  assign n37098 = pi1153 & ~n37097;
  assign n37099 = ~n37096 & n37098;
  assign n37100 = pi608 & ~n37099;
  assign n37101 = ~n36897 & n37100;
  assign n37102 = ~n37095 & ~n37101;
  assign n37103 = pi778 & ~n37102;
  assign n37104 = ~pi778 & n37089;
  assign n37105 = ~n37103 & ~n37104;
  assign n37106 = ~pi609 & ~n37105;
  assign n37107 = pi609 & n36900;
  assign n37108 = ~pi1155 & ~n37107;
  assign n37109 = ~n37106 & n37108;
  assign n37110 = ~pi660 & ~n36778;
  assign n37111 = ~n37109 & n37110;
  assign n37112 = pi609 & ~n37105;
  assign n37113 = ~pi609 & n36900;
  assign n37114 = pi1155 & ~n37113;
  assign n37115 = ~n37112 & n37114;
  assign n37116 = pi660 & ~n36782;
  assign n37117 = ~n37115 & n37116;
  assign n37118 = ~n37111 & ~n37117;
  assign n37119 = pi785 & ~n37118;
  assign n37120 = ~pi785 & ~n37105;
  assign n37121 = ~n37119 & ~n37120;
  assign n37122 = ~pi618 & ~n37121;
  assign n37123 = pi618 & ~n36902;
  assign n37124 = ~pi1154 & ~n37123;
  assign n37125 = ~n37122 & n37124;
  assign n37126 = ~pi627 & ~n36790;
  assign n37127 = ~n37125 & n37126;
  assign n37128 = pi618 & ~n37121;
  assign n37129 = ~pi618 & ~n36902;
  assign n37130 = pi1154 & ~n37129;
  assign n37131 = ~n37128 & n37130;
  assign n37132 = pi627 & ~n36794;
  assign n37133 = ~n37131 & n37132;
  assign n37134 = ~n37127 & ~n37133;
  assign n37135 = pi781 & ~n37134;
  assign n37136 = ~pi781 & ~n37121;
  assign n37137 = ~n37135 & ~n37136;
  assign n37138 = pi619 & ~n37137;
  assign n37139 = ~pi619 & n36905;
  assign n37140 = pi1159 & ~n37139;
  assign n37141 = ~n37138 & n37140;
  assign n37142 = pi648 & ~n36806;
  assign n37143 = ~n37141 & n37142;
  assign n37144 = ~pi619 & ~n37137;
  assign n37145 = pi619 & n36905;
  assign n37146 = ~pi1159 & ~n37145;
  assign n37147 = ~n37144 & n37146;
  assign n37148 = ~pi648 & ~n36802;
  assign n37149 = ~n37147 & n37148;
  assign n37150 = pi789 & ~n37149;
  assign n37151 = ~n37143 & n37150;
  assign n37152 = ~pi789 & n37137;
  assign n37153 = n17817 & ~n37152;
  assign n37154 = ~n37151 & n37153;
  assign n37155 = ~n36950 & ~n37154;
  assign n37156 = ~n36936 & ~n37155;
  assign n37157 = n20205 & n36935;
  assign n37158 = n20207 & ~n37157;
  assign n37159 = ~n37156 & n37158;
  assign n37160 = ~n36924 & ~n37159;
  assign n37161 = pi644 & n37160;
  assign n37162 = ~pi787 & n36911;
  assign n37163 = ~n36915 & ~n36920;
  assign n37164 = pi787 & ~n37163;
  assign n37165 = ~n37162 & ~n37164;
  assign n37166 = ~pi644 & n37165;
  assign n37167 = pi715 & ~n37166;
  assign n37168 = ~n37161 & n37167;
  assign n37169 = n17652 & ~n36638;
  assign n37170 = ~n17652 & n36814;
  assign n37171 = ~n37169 & ~n37170;
  assign n37172 = pi644 & ~n37171;
  assign n37173 = ~pi644 & ~n36638;
  assign n37174 = ~pi715 & ~n37173;
  assign n37175 = ~n37172 & n37174;
  assign n37176 = pi1160 & ~n37175;
  assign n37177 = ~n37168 & n37176;
  assign n37178 = ~pi644 & n37160;
  assign n37179 = pi644 & n37165;
  assign n37180 = ~pi715 & ~n37179;
  assign n37181 = ~n37178 & n37180;
  assign n37182 = ~pi644 & ~n37171;
  assign n37183 = pi644 & ~n36638;
  assign n37184 = pi715 & ~n37183;
  assign n37185 = ~n37182 & n37184;
  assign n37186 = ~pi1160 & ~n37185;
  assign n37187 = ~n37181 & n37186;
  assign n37188 = ~n37177 & ~n37187;
  assign n37189 = pi790 & ~n37188;
  assign n37190 = ~pi790 & n37160;
  assign n37191 = ~n37189 & ~n37190;
  assign n37192 = ~po1038 & ~n37191;
  assign n37193 = ~pi223 & po1038;
  assign po380 = ~n37192 & ~n37193;
  assign n37195 = pi224 & ~n36026;
  assign n37196 = n17816 & ~n37195;
  assign n37197 = pi224 & ~n3267;
  assign n37198 = pi614 & n16521;
  assign n37199 = n16518 & ~n37198;
  assign n37200 = ~n6157 & ~n37199;
  assign n37201 = ~n16574 & ~n37200;
  assign n37202 = ~n16512 & ~n37201;
  assign n37203 = ~pi680 & ~n37201;
  assign n37204 = pi680 & n37198;
  assign n37205 = ~n17137 & ~n37204;
  assign n37206 = ~n37203 & n37205;
  assign n37207 = n16512 & ~n37206;
  assign n37208 = ~n37202 & ~n37207;
  assign n37209 = n6215 & n37208;
  assign n37210 = pi614 & ~n16741;
  assign n37211 = n16585 & ~n16744;
  assign n37212 = ~n37210 & ~n37211;
  assign n37213 = ~pi680 & ~n37212;
  assign n37214 = pi680 & ~n17219;
  assign n37215 = ~n35778 & n37214;
  assign n37216 = ~n37213 & ~n37215;
  assign n37217 = n16512 & ~n37216;
  assign n37218 = ~n16512 & ~n37212;
  assign n37219 = ~n37217 & ~n37218;
  assign n37220 = ~n6215 & n37219;
  assign n37221 = pi224 & ~n37220;
  assign n37222 = ~n37209 & n37221;
  assign n37223 = pi614 & ~n36092;
  assign n37224 = ~pi224 & n37223;
  assign n37225 = ~n17268 & n37224;
  assign n37226 = pi223 & ~n37225;
  assign n37227 = ~n37222 & n37226;
  assign n37228 = ~n16636 & ~n37200;
  assign n37229 = ~n16512 & ~n37228;
  assign n37230 = ~pi680 & ~n37228;
  assign n37231 = ~n17163 & ~n37204;
  assign n37232 = ~n37230 & n37231;
  assign n37233 = n16512 & ~n37232;
  assign n37234 = ~n37229 & ~n37233;
  assign n37235 = n6215 & n37234;
  assign n37236 = n16652 & ~n37198;
  assign n37237 = ~n16512 & ~n37236;
  assign n37238 = ~pi680 & ~n37236;
  assign n37239 = pi614 & n16657;
  assign n37240 = pi680 & ~n37239;
  assign n37241 = n16619 & n37240;
  assign n37242 = ~n37204 & ~n37241;
  assign n37243 = ~n37238 & n37242;
  assign n37244 = n16512 & ~n37243;
  assign n37245 = ~n37237 & ~n37244;
  assign n37246 = ~n6215 & n37245;
  assign n37247 = pi224 & ~n37246;
  assign n37248 = ~n37235 & n37247;
  assign n37249 = ~n16649 & n37198;
  assign n37250 = ~pi680 & ~n37249;
  assign n37251 = ~n37240 & ~n37250;
  assign n37252 = n16512 & ~n37251;
  assign n37253 = ~n16512 & ~n37249;
  assign n37254 = ~n37252 & ~n37253;
  assign n37255 = ~n6215 & ~n37254;
  assign n37256 = pi614 & ~n36064;
  assign n37257 = n6215 & ~n37256;
  assign n37258 = n5770 & ~n37257;
  assign n37259 = ~n37255 & n37258;
  assign n37260 = pi614 & n16782;
  assign n37261 = ~pi223 & ~n37260;
  assign n37262 = ~n37259 & n37261;
  assign n37263 = ~n37248 & n37262;
  assign n37264 = ~n37227 & ~n37263;
  assign n37265 = ~pi299 & ~n37264;
  assign n37266 = n6189 & n37234;
  assign n37267 = ~n6189 & n37245;
  assign n37268 = pi224 & ~n37267;
  assign n37269 = ~n37266 & n37268;
  assign n37270 = ~n6189 & ~n37254;
  assign n37271 = n6189 & ~n37256;
  assign n37272 = ~pi224 & ~n37271;
  assign n37273 = ~n37270 & n37272;
  assign n37274 = ~n3329 & ~n37273;
  assign n37275 = ~n37269 & n37274;
  assign n37276 = pi224 & ~n16518;
  assign n37277 = n3329 & ~n37276;
  assign n37278 = n16521 & n17167;
  assign n37279 = n37277 & ~n37278;
  assign n37280 = ~pi215 & ~n37279;
  assign n37281 = ~n37275 & n37280;
  assign n37282 = ~n17258 & n37224;
  assign n37283 = n6189 & n37208;
  assign n37284 = ~n6189 & n37219;
  assign n37285 = pi224 & ~n37284;
  assign n37286 = ~n37283 & n37285;
  assign n37287 = ~n37282 & ~n37286;
  assign n37288 = pi215 & ~n37287;
  assign n37289 = pi299 & ~n37288;
  assign n37290 = ~n37281 & n37289;
  assign n37291 = pi39 & ~n37290;
  assign n37292 = ~n37265 & n37291;
  assign n37293 = pi614 & n17084;
  assign n37294 = pi224 & n17018;
  assign n37295 = n37293 & ~n37294;
  assign n37296 = pi224 & ~n17026;
  assign n37297 = ~n37295 & ~n37296;
  assign n37298 = pi299 & n37297;
  assign n37299 = ~pi614 & n17079;
  assign n37300 = pi224 & ~n37299;
  assign n37301 = n17040 & n37300;
  assign n37302 = pi614 & n17079;
  assign n37303 = ~pi224 & n37302;
  assign n37304 = ~pi299 & ~n37303;
  assign n37305 = ~n37301 & n37304;
  assign n37306 = ~pi39 & ~n37305;
  assign n37307 = ~n37298 & n37306;
  assign n37308 = ~pi38 & ~n37307;
  assign n37309 = ~n37292 & n37308;
  assign n37310 = pi224 & ~n17280;
  assign n37311 = pi38 & ~n37310;
  assign n37312 = pi614 & n17282;
  assign n37313 = n37311 & ~n37312;
  assign n37314 = n3267 & ~n37313;
  assign n37315 = ~n37309 & n37314;
  assign n37316 = ~n37197 & ~n37315;
  assign n37317 = ~n17438 & ~n37316;
  assign n37318 = n17438 & n37195;
  assign n37319 = ~n37317 & ~n37318;
  assign n37320 = ~pi785 & ~n37319;
  assign n37321 = pi609 & n37319;
  assign n37322 = ~pi609 & ~n37195;
  assign n37323 = pi1155 & ~n37322;
  assign n37324 = ~n37321 & n37323;
  assign n37325 = ~pi609 & n37319;
  assign n37326 = pi609 & ~n37195;
  assign n37327 = ~pi1155 & ~n37326;
  assign n37328 = ~n37325 & n37327;
  assign n37329 = ~n37324 & ~n37328;
  assign n37330 = pi785 & ~n37329;
  assign n37331 = ~n37320 & ~n37330;
  assign n37332 = ~pi781 & ~n37331;
  assign n37333 = pi618 & n37331;
  assign n37334 = ~pi618 & ~n37195;
  assign n37335 = pi1154 & ~n37334;
  assign n37336 = ~n37333 & n37335;
  assign n37337 = ~pi618 & n37331;
  assign n37338 = pi618 & ~n37195;
  assign n37339 = ~pi1154 & ~n37338;
  assign n37340 = ~n37337 & n37339;
  assign n37341 = ~n37336 & ~n37340;
  assign n37342 = pi781 & ~n37341;
  assign n37343 = ~n37332 & ~n37342;
  assign n37344 = ~pi789 & ~n37343;
  assign n37345 = pi619 & n37343;
  assign n37346 = ~pi619 & ~n37195;
  assign n37347 = pi1159 & ~n37346;
  assign n37348 = ~n37345 & n37347;
  assign n37349 = ~pi619 & n37343;
  assign n37350 = pi619 & ~n37195;
  assign n37351 = ~pi1159 & ~n37350;
  assign n37352 = ~n37349 & n37351;
  assign n37353 = ~n37348 & ~n37352;
  assign n37354 = pi789 & ~n37353;
  assign n37355 = ~n37344 & ~n37354;
  assign n37356 = ~n17816 & n37355;
  assign n37357 = ~n37196 & ~n37356;
  assign n37358 = ~n20409 & n37357;
  assign n37359 = ~n19126 & ~n37195;
  assign n37360 = ~pi224 & ~n17054;
  assign n37361 = pi662 & pi680;
  assign n37362 = n17054 & ~n37361;
  assign n37363 = pi224 & n17074;
  assign n37364 = pi299 & ~n37363;
  assign n37365 = ~n37362 & n37364;
  assign n37366 = ~n37360 & n37365;
  assign n37367 = ~pi224 & ~n17049;
  assign n37368 = n17049 & ~n37361;
  assign n37369 = pi224 & n17068;
  assign n37370 = ~pi299 & ~n37369;
  assign n37371 = ~n37368 & n37370;
  assign n37372 = ~n37367 & n37371;
  assign n37373 = ~pi39 & ~n37372;
  assign n37374 = ~n37366 & n37373;
  assign n37375 = n16689 & n37361;
  assign n37376 = n37277 & ~n37375;
  assign n37377 = pi662 & ~n17338;
  assign n37378 = ~pi662 & ~n17172;
  assign n37379 = ~n37377 & ~n37378;
  assign n37380 = n6189 & n37379;
  assign n37381 = ~n6158 & ~n36204;
  assign n37382 = n16812 & ~n37381;
  assign n37383 = ~n6189 & n37382;
  assign n37384 = pi224 & ~n37383;
  assign n37385 = ~n37380 & n37384;
  assign n37386 = ~n17303 & n37361;
  assign n37387 = n6189 & ~n37386;
  assign n37388 = pi662 & n17298;
  assign n37389 = ~n6189 & ~n37388;
  assign n37390 = ~pi224 & ~n37389;
  assign n37391 = ~n37387 & n37390;
  assign n37392 = ~n3329 & ~n37391;
  assign n37393 = ~n37385 & n37392;
  assign n37394 = ~n37376 & ~n37393;
  assign n37395 = ~pi215 & ~n37394;
  assign n37396 = ~pi662 & ~n17132;
  assign n37397 = pi662 & ~n17358;
  assign n37398 = ~n37396 & ~n37397;
  assign n37399 = ~n6189 & n37398;
  assign n37400 = ~pi662 & ~n17151;
  assign n37401 = pi662 & ~n36223;
  assign n37402 = ~n37400 & ~n37401;
  assign n37403 = n6189 & n37402;
  assign n37404 = pi224 & ~n37403;
  assign n37405 = ~n37399 & n37404;
  assign n37406 = ~pi224 & pi662;
  assign n37407 = n17327 & n37406;
  assign n37408 = pi215 & ~n37407;
  assign n37409 = ~n37405 & n37408;
  assign n37410 = pi299 & ~n37409;
  assign n37411 = ~n37395 & n37410;
  assign n37412 = n6215 & n37379;
  assign n37413 = ~n6215 & n37382;
  assign n37414 = pi224 & ~n37413;
  assign n37415 = ~n37412 & n37414;
  assign n37416 = n6215 & ~n37386;
  assign n37417 = ~n6215 & ~n37388;
  assign n37418 = n5770 & ~n37417;
  assign n37419 = ~n37416 & n37418;
  assign n37420 = pi662 & n17297;
  assign n37421 = ~pi223 & ~n37420;
  assign n37422 = ~n37419 & n37421;
  assign n37423 = ~n37415 & n37422;
  assign n37424 = ~n6215 & n37398;
  assign n37425 = n6215 & n37402;
  assign n37426 = pi224 & ~n37425;
  assign n37427 = ~n37424 & n37426;
  assign n37428 = n17314 & n37406;
  assign n37429 = pi223 & ~n37428;
  assign n37430 = ~n37427 & n37429;
  assign n37431 = ~pi299 & ~n37430;
  assign n37432 = ~n37423 & n37431;
  assign n37433 = pi39 & ~n37432;
  assign n37434 = ~n37411 & n37433;
  assign n37435 = ~n37374 & ~n37434;
  assign n37436 = ~pi38 & ~n37435;
  assign n37437 = pi662 & n17391;
  assign n37438 = n37311 & ~n37437;
  assign n37439 = n3267 & ~n37438;
  assign n37440 = ~n37436 & n37439;
  assign n37441 = ~n37197 & ~n37440;
  assign n37442 = ~pi778 & ~n37441;
  assign n37443 = pi625 & n37441;
  assign n37444 = ~pi625 & ~n37195;
  assign n37445 = pi1153 & ~n37444;
  assign n37446 = ~n37443 & n37445;
  assign n37447 = ~pi625 & n37441;
  assign n37448 = pi625 & ~n37195;
  assign n37449 = ~pi1153 & ~n37448;
  assign n37450 = ~n37447 & n37449;
  assign n37451 = ~n37446 & ~n37450;
  assign n37452 = pi778 & ~n37451;
  assign n37453 = ~n37442 & ~n37452;
  assign n37454 = ~n17466 & ~n37453;
  assign n37455 = n17466 & n37195;
  assign n37456 = ~n37454 & ~n37455;
  assign n37457 = ~n17503 & ~n37456;
  assign n37458 = n17503 & n37195;
  assign n37459 = ~n37457 & ~n37458;
  assign n37460 = ~n17539 & n37459;
  assign n37461 = ~n17582 & n37460;
  assign n37462 = ~n37359 & ~n37461;
  assign n37463 = ~pi628 & ~n37462;
  assign n37464 = pi628 & ~n37195;
  assign n37465 = n17608 & ~n37464;
  assign n37466 = ~n37463 & n37465;
  assign n37467 = pi628 & ~n37462;
  assign n37468 = ~pi628 & ~n37195;
  assign n37469 = n17607 & ~n37468;
  assign n37470 = ~n37467 & n37469;
  assign n37471 = ~n37466 & ~n37470;
  assign n37472 = ~n37358 & n37471;
  assign n37473 = pi792 & ~n37472;
  assign n37474 = pi614 & ~n36318;
  assign n37475 = ~pi614 & pi616;
  assign n37476 = n36307 & n37475;
  assign n37477 = ~n37474 & ~n37476;
  assign n37478 = ~n36316 & n37477;
  assign n37479 = pi680 & ~n37478;
  assign n37480 = ~n37238 & ~n37479;
  assign n37481 = pi662 & ~n37480;
  assign n37482 = ~pi662 & ~n16511;
  assign n37483 = ~n37236 & n37482;
  assign n37484 = ~n37244 & ~n37483;
  assign n37485 = ~n37481 & n37484;
  assign n37486 = pi224 & n37485;
  assign n37487 = n16706 & n37361;
  assign n37488 = ~n37254 & ~n37487;
  assign n37489 = ~pi224 & n37488;
  assign n37490 = ~n6189 & ~n37489;
  assign n37491 = ~n37486 & n37490;
  assign n37492 = ~pi614 & ~n23906;
  assign n37493 = pi614 & ~n36478;
  assign n37494 = ~n37492 & ~n37493;
  assign n37495 = ~n16515 & n37494;
  assign n37496 = pi616 & ~n37495;
  assign n37497 = pi614 & ~n16891;
  assign n37498 = ~n16627 & ~n37497;
  assign n37499 = ~pi616 & ~n37498;
  assign n37500 = ~n37496 & ~n37499;
  assign n37501 = pi680 & ~n37500;
  assign n37502 = ~n37230 & ~n37501;
  assign n37503 = pi662 & ~n37502;
  assign n37504 = ~n37228 & n37482;
  assign n37505 = ~n37233 & ~n37504;
  assign n37506 = ~n37503 & n37505;
  assign n37507 = pi224 & n37506;
  assign n37508 = ~n16714 & n37475;
  assign n37509 = ~n36351 & ~n37508;
  assign n37510 = pi680 & ~n37509;
  assign n37511 = ~n36352 & ~n37278;
  assign n37512 = ~n37510 & ~n37511;
  assign n37513 = pi662 & ~n37512;
  assign n37514 = ~pi662 & ~n37256;
  assign n37515 = ~n37513 & ~n37514;
  assign n37516 = ~pi224 & ~n37515;
  assign n37517 = n6189 & ~n37516;
  assign n37518 = ~n37507 & n37517;
  assign n37519 = ~n3329 & ~n37518;
  assign n37520 = ~n37491 & n37519;
  assign n37521 = n16714 & n37361;
  assign n37522 = ~n37278 & ~n37521;
  assign n37523 = ~pi224 & ~n37522;
  assign n37524 = n37361 & n37494;
  assign n37525 = ~n37198 & ~n37361;
  assign n37526 = n16529 & n37525;
  assign n37527 = pi224 & ~n37526;
  assign n37528 = ~n37524 & n37527;
  assign n37529 = n37277 & ~n37528;
  assign n37530 = ~n37523 & n37529;
  assign n37531 = ~pi215 & ~n37530;
  assign n37532 = ~n37520 & n37531;
  assign n37533 = ~n16560 & ~n37497;
  assign n37534 = ~pi616 & ~n37533;
  assign n37535 = ~n37496 & ~n37534;
  assign n37536 = pi680 & ~n37535;
  assign n37537 = ~n37203 & ~n37536;
  assign n37538 = pi662 & ~n37537;
  assign n37539 = ~n37201 & n37482;
  assign n37540 = ~n37207 & ~n37539;
  assign n37541 = ~n37538 & n37540;
  assign n37542 = n6189 & ~n37541;
  assign n37543 = n16594 & ~n37198;
  assign n37544 = pi680 & ~n37543;
  assign n37545 = ~n37213 & ~n37544;
  assign n37546 = pi662 & ~n37545;
  assign n37547 = ~n37212 & n37482;
  assign n37548 = ~n37217 & ~n37547;
  assign n37549 = ~n37546 & n37548;
  assign n37550 = ~n6189 & ~n37549;
  assign n37551 = pi224 & ~n37550;
  assign n37552 = ~n37542 & n37551;
  assign n37553 = pi680 & n16765;
  assign n37554 = ~n37278 & ~n37553;
  assign n37555 = pi662 & n37554;
  assign n37556 = ~pi662 & ~n37223;
  assign n37557 = ~n37555 & ~n37556;
  assign n37558 = n6189 & n37557;
  assign n37559 = ~n16583 & n37223;
  assign n37560 = ~pi662 & ~n37559;
  assign n37561 = ~pi614 & n16743;
  assign n37562 = pi614 & n36397;
  assign n37563 = pi680 & ~n37562;
  assign n37564 = ~n37561 & n37563;
  assign n37565 = ~n16753 & n37564;
  assign n37566 = pi614 & ~pi680;
  assign n37567 = n16588 & n37566;
  assign n37568 = pi662 & ~n37567;
  assign n37569 = ~n37565 & n37568;
  assign n37570 = ~n37560 & ~n37569;
  assign n37571 = ~n6189 & n37570;
  assign n37572 = ~pi224 & ~n37571;
  assign n37573 = ~n37558 & n37572;
  assign n37574 = pi215 & ~n37573;
  assign n37575 = ~n37552 & n37574;
  assign n37576 = pi299 & ~n37575;
  assign n37577 = ~n37532 & n37576;
  assign n37578 = n6215 & n37506;
  assign n37579 = ~n6215 & n37485;
  assign n37580 = pi224 & ~n37579;
  assign n37581 = ~n37578 & n37580;
  assign n37582 = ~n6215 & n37488;
  assign n37583 = n6215 & ~n37515;
  assign n37584 = n5770 & ~n37583;
  assign n37585 = ~n37582 & n37584;
  assign n37586 = ~pi222 & n37523;
  assign n37587 = ~pi223 & ~n37586;
  assign n37588 = ~n37585 & n37587;
  assign n37589 = ~n37581 & n37588;
  assign n37590 = pi224 & n37541;
  assign n37591 = ~pi224 & ~n37557;
  assign n37592 = n6215 & ~n37591;
  assign n37593 = ~n37590 & n37592;
  assign n37594 = pi224 & n37549;
  assign n37595 = ~pi224 & ~n37570;
  assign n37596 = ~n6215 & ~n37595;
  assign n37597 = ~n37594 & n37596;
  assign n37598 = pi223 & ~n37597;
  assign n37599 = ~n37593 & n37598;
  assign n37600 = ~n37589 & ~n37599;
  assign n37601 = ~pi299 & ~n37600;
  assign n37602 = pi39 & ~n37601;
  assign n37603 = ~n37577 & n37602;
  assign n37604 = n18447 & n37361;
  assign n37605 = ~n37302 & ~n37604;
  assign n37606 = ~pi224 & ~n37605;
  assign n37607 = n18447 & ~n37361;
  assign n37608 = ~n36468 & n37300;
  assign n37609 = ~n37607 & n37608;
  assign n37610 = ~n37606 & ~n37609;
  assign n37611 = ~pi299 & ~n37610;
  assign n37612 = ~pi614 & n17084;
  assign n37613 = ~n36452 & ~n37612;
  assign n37614 = pi224 & ~n37613;
  assign n37615 = ~pi224 & ~n18457;
  assign n37616 = ~n37293 & n37615;
  assign n37617 = ~n37614 & ~n37616;
  assign n37618 = n37361 & ~n37617;
  assign n37619 = n37297 & ~n37361;
  assign n37620 = pi299 & ~n37619;
  assign n37621 = ~n37618 & n37620;
  assign n37622 = ~n37611 & ~n37621;
  assign n37623 = ~pi39 & ~n37622;
  assign n37624 = ~pi38 & ~n37623;
  assign n37625 = ~n37603 & n37624;
  assign n37626 = pi662 & n16667;
  assign n37627 = n17280 & n37626;
  assign n37628 = n37313 & ~n37627;
  assign n37629 = n3267 & ~n37628;
  assign n37630 = ~n37625 & n37629;
  assign n37631 = ~n37197 & ~n37630;
  assign n37632 = ~pi625 & n37631;
  assign n37633 = pi625 & n37316;
  assign n37634 = ~pi1153 & ~n37633;
  assign n37635 = ~n37632 & n37634;
  assign n37636 = ~pi608 & ~n37446;
  assign n37637 = ~n37635 & n37636;
  assign n37638 = pi625 & n37631;
  assign n37639 = ~pi625 & n37316;
  assign n37640 = pi1153 & ~n37639;
  assign n37641 = ~n37638 & n37640;
  assign n37642 = pi608 & ~n37450;
  assign n37643 = ~n37641 & n37642;
  assign n37644 = ~n37637 & ~n37643;
  assign n37645 = pi778 & ~n37644;
  assign n37646 = ~pi778 & n37631;
  assign n37647 = ~n37645 & ~n37646;
  assign n37648 = ~pi609 & ~n37647;
  assign n37649 = pi609 & n37453;
  assign n37650 = ~pi1155 & ~n37649;
  assign n37651 = ~n37648 & n37650;
  assign n37652 = ~pi660 & ~n37324;
  assign n37653 = ~n37651 & n37652;
  assign n37654 = pi609 & ~n37647;
  assign n37655 = ~pi609 & n37453;
  assign n37656 = pi1155 & ~n37655;
  assign n37657 = ~n37654 & n37656;
  assign n37658 = pi660 & ~n37328;
  assign n37659 = ~n37657 & n37658;
  assign n37660 = ~n37653 & ~n37659;
  assign n37661 = pi785 & ~n37660;
  assign n37662 = ~pi785 & ~n37647;
  assign n37663 = ~n37661 & ~n37662;
  assign n37664 = ~pi618 & ~n37663;
  assign n37665 = pi618 & n37456;
  assign n37666 = ~pi1154 & ~n37665;
  assign n37667 = ~n37664 & n37666;
  assign n37668 = ~pi627 & ~n37336;
  assign n37669 = ~n37667 & n37668;
  assign n37670 = pi618 & ~n37663;
  assign n37671 = ~pi618 & n37456;
  assign n37672 = pi1154 & ~n37671;
  assign n37673 = ~n37670 & n37672;
  assign n37674 = pi627 & ~n37340;
  assign n37675 = ~n37673 & n37674;
  assign n37676 = ~n37669 & ~n37675;
  assign n37677 = pi781 & ~n37676;
  assign n37678 = ~pi781 & ~n37663;
  assign n37679 = ~n37677 & ~n37678;
  assign n37680 = pi619 & ~n37679;
  assign n37681 = ~pi619 & n37459;
  assign n37682 = pi1159 & ~n37681;
  assign n37683 = ~n37680 & n37682;
  assign n37684 = pi648 & ~n37352;
  assign n37685 = ~n37683 & n37684;
  assign n37686 = ~pi619 & ~n37679;
  assign n37687 = pi619 & n37459;
  assign n37688 = ~pi1159 & ~n37687;
  assign n37689 = ~n37686 & n37688;
  assign n37690 = ~pi648 & ~n37348;
  assign n37691 = ~n37689 & n37690;
  assign n37692 = pi789 & ~n37691;
  assign n37693 = ~n37685 & n37692;
  assign n37694 = ~pi789 & n37679;
  assign n37695 = n17817 & ~n37694;
  assign n37696 = ~n37693 & n37695;
  assign n37697 = ~pi626 & ~n37355;
  assign n37698 = pi626 & n37195;
  assign n37699 = n17580 & ~n37698;
  assign n37700 = ~n37697 & n37699;
  assign n37701 = n17539 & ~n37195;
  assign n37702 = ~n37460 & ~n37701;
  assign n37703 = n17704 & ~n37702;
  assign n37704 = pi626 & ~n37355;
  assign n37705 = ~pi626 & n37195;
  assign n37706 = n17579 & ~n37705;
  assign n37707 = ~n37704 & n37706;
  assign n37708 = ~n37703 & ~n37707;
  assign n37709 = ~n37700 & n37708;
  assign n37710 = pi788 & ~n37709;
  assign n37711 = ~n20205 & ~n37710;
  assign n37712 = ~n37696 & n37711;
  assign n37713 = ~n37473 & ~n37712;
  assign n37714 = n20207 & ~n37713;
  assign n37715 = ~n17610 & n37357;
  assign n37716 = n17610 & n37195;
  assign n37717 = ~n37715 & ~n37716;
  assign n37718 = ~n20398 & ~n37717;
  assign n37719 = ~n19158 & ~n37462;
  assign n37720 = n17858 & ~n37195;
  assign n37721 = ~n37719 & ~n37720;
  assign n37722 = pi647 & ~n37721;
  assign n37723 = ~pi647 & ~n37195;
  assign n37724 = pi1157 & ~n37723;
  assign n37725 = ~n37722 & n37724;
  assign n37726 = ~pi630 & n37725;
  assign n37727 = ~pi647 & ~n37721;
  assign n37728 = pi647 & ~n37195;
  assign n37729 = ~pi1157 & ~n37728;
  assign n37730 = ~n37727 & n37729;
  assign n37731 = pi630 & n37730;
  assign n37732 = ~n37726 & ~n37731;
  assign n37733 = ~n37718 & n37732;
  assign n37734 = pi787 & ~n37733;
  assign n37735 = ~n37714 & ~n37734;
  assign n37736 = pi644 & n37735;
  assign n37737 = ~pi787 & n37721;
  assign n37738 = ~n37725 & ~n37730;
  assign n37739 = pi787 & ~n37738;
  assign n37740 = ~n37737 & ~n37739;
  assign n37741 = ~pi644 & n37740;
  assign n37742 = pi715 & ~n37741;
  assign n37743 = ~n37736 & n37742;
  assign n37744 = n17652 & ~n37195;
  assign n37745 = ~n17652 & n37717;
  assign n37746 = ~n37744 & ~n37745;
  assign n37747 = pi644 & ~n37746;
  assign n37748 = ~pi644 & ~n37195;
  assign n37749 = ~pi715 & ~n37748;
  assign n37750 = ~n37747 & n37749;
  assign n37751 = pi1160 & ~n37750;
  assign n37752 = ~n37743 & n37751;
  assign n37753 = ~pi644 & n37735;
  assign n37754 = pi644 & n37740;
  assign n37755 = ~pi715 & ~n37754;
  assign n37756 = ~n37753 & n37755;
  assign n37757 = ~pi644 & ~n37746;
  assign n37758 = pi644 & ~n37195;
  assign n37759 = pi715 & ~n37758;
  assign n37760 = ~n37757 & n37759;
  assign n37761 = ~pi1160 & ~n37760;
  assign n37762 = ~n37756 & n37761;
  assign n37763 = ~n37752 & ~n37762;
  assign n37764 = pi790 & ~n37763;
  assign n37765 = ~pi790 & n37735;
  assign n37766 = ~n37764 & ~n37765;
  assign n37767 = ~po1038 & ~n37766;
  assign n37768 = ~pi224 & po1038;
  assign po381 = ~n37767 & ~n37768;
  assign n37770 = ~n6143 & ~n6243;
  assign n37771 = ~pi137 & ~n37770;
  assign n37772 = n6236 & ~n37771;
  assign n37773 = n2921 & ~n11354;
  assign n37774 = ~n2713 & n37773;
  assign n37775 = n2556 & ~n37774;
  assign n37776 = n2554 & ~n37775;
  assign n37777 = ~n2742 & ~n37776;
  assign n37778 = ~pi95 & ~n37777;
  assign n37779 = ~n2727 & ~n37778;
  assign n37780 = pi137 & ~n37779;
  assign n37781 = n2450 & n11354;
  assign n37782 = n2785 & ~n37781;
  assign n37783 = n2747 & ~n37782;
  assign n37784 = ~pi137 & ~n37783;
  assign n37785 = ~n37780 & ~n37784;
  assign n37786 = pi332 & ~n37785;
  assign n37787 = ~n2727 & ~n2744;
  assign n37788 = pi137 & ~n37787;
  assign n37789 = ~n2823 & ~n37788;
  assign n37790 = ~pi332 & ~n37789;
  assign n37791 = ~n37786 & ~n37790;
  assign n37792 = n2988 & n37791;
  assign n37793 = pi1093 & ~n37783;
  assign n37794 = n2747 & n7491;
  assign n37795 = n2450 & ~n7446;
  assign n37796 = ~n2531 & n37795;
  assign n37797 = ~pi32 & ~n37796;
  assign n37798 = n37794 & ~n37797;
  assign n37799 = ~pi1093 & ~n37798;
  assign n37800 = ~n7491 & n37783;
  assign n37801 = n11353 & n37795;
  assign n37802 = n37794 & n37801;
  assign n37803 = ~n37800 & ~n37802;
  assign n37804 = n37799 & n37803;
  assign n37805 = ~n37793 & ~n37804;
  assign n37806 = n11485 & ~n37805;
  assign n37807 = n2822 & ~n7491;
  assign n37808 = n37799 & ~n37807;
  assign n37809 = ~n2767 & n37795;
  assign n37810 = ~pi32 & ~n37809;
  assign n37811 = n37794 & ~n37810;
  assign n37812 = pi1093 & ~n37807;
  assign n37813 = ~n37811 & n37812;
  assign n37814 = ~n37808 & ~n37813;
  assign n37815 = n11452 & ~n37814;
  assign n37816 = n37803 & n37815;
  assign n37817 = ~n37806 & ~n37816;
  assign n37818 = ~n37780 & n37817;
  assign n37819 = pi332 & ~n37818;
  assign n37820 = pi1093 & ~n2822;
  assign n37821 = ~n37808 & ~n37820;
  assign n37822 = n11485 & ~n37821;
  assign n37823 = ~n37815 & ~n37822;
  assign n37824 = ~n37788 & n37823;
  assign n37825 = ~pi332 & ~n37824;
  assign n37826 = ~n37819 & ~n37825;
  assign n37827 = ~n2988 & n37826;
  assign n37828 = ~pi210 & ~n37827;
  assign n37829 = ~n37792 & n37828;
  assign n37830 = ~n2724 & ~n2727;
  assign n37831 = pi137 & ~n37830;
  assign n37832 = ~n2787 & ~n37831;
  assign n37833 = ~pi332 & ~n37832;
  assign n37834 = ~n2501 & ~n37776;
  assign n37835 = ~pi95 & ~n37834;
  assign n37836 = n3020 & ~n37835;
  assign n37837 = ~pi137 & n2502;
  assign n37838 = ~n37782 & n37837;
  assign n37839 = pi332 & ~n37838;
  assign n37840 = ~n37836 & n37839;
  assign n37841 = ~n37833 & ~n37840;
  assign n37842 = pi210 & ~n37841;
  assign n37843 = pi299 & ~n37842;
  assign n37844 = ~n37829 & n37843;
  assign n37845 = ~n6483 & n37826;
  assign n37846 = n6483 & n37791;
  assign n37847 = ~pi198 & ~n37846;
  assign n37848 = ~n37845 & n37847;
  assign n37849 = pi198 & ~n37841;
  assign n37850 = ~pi299 & ~n37849;
  assign n37851 = ~n37848 & n37850;
  assign n37852 = ~n37844 & ~n37851;
  assign n37853 = ~pi39 & ~n37852;
  assign n37854 = pi39 & n3110;
  assign n37855 = ~pi38 & ~n37854;
  assign n37856 = ~n37853 & n37855;
  assign n37857 = pi38 & ~pi137;
  assign n37858 = n6111 & ~n37857;
  assign n37859 = ~n37856 & n37858;
  assign n37860 = ~n37772 & ~n37859;
  assign n37861 = ~pi87 & ~n37860;
  assign n37862 = n3110 & n3207;
  assign n37863 = pi87 & n37862;
  assign n37864 = ~pi75 & ~n37863;
  assign n37865 = ~n37861 & n37864;
  assign n37866 = n7268 & ~n37771;
  assign n37867 = pi75 & ~n37866;
  assign n37868 = ~pi92 & ~n37867;
  assign n37869 = ~n37865 & n37868;
  assign n37870 = pi92 & n3230;
  assign n37871 = n37862 & n37870;
  assign n37872 = ~pi54 & ~n37871;
  assign n37873 = ~n37869 & n37872;
  assign n37874 = n3277 & n37862;
  assign n37875 = pi54 & ~n37874;
  assign n37876 = ~pi74 & ~n37875;
  assign n37877 = ~n37873 & n37876;
  assign n37878 = pi74 & n6105;
  assign n37879 = n37862 & n37878;
  assign n37880 = ~pi55 & ~n37879;
  assign n37881 = ~n37877 & n37880;
  assign n37882 = n7315 & ~n37881;
  assign n37883 = pi56 & n3279;
  assign n37884 = n37862 & n37883;
  assign n37885 = ~n37882 & ~n37884;
  assign n37886 = ~pi62 & ~n37885;
  assign n37887 = n3430 & n37862;
  assign n37888 = pi62 & n37887;
  assign n37889 = n3429 & ~n37888;
  assign n37890 = ~n37886 & n37889;
  assign n37891 = ~pi62 & n37887;
  assign n37892 = ~n3429 & ~n37891;
  assign n37893 = ~n6097 & ~n37892;
  assign po382 = ~n37890 & n37893;
  assign n37895 = pi228 & pi231;
  assign n37896 = ~n2525 & ~n2867;
  assign n37897 = ~pi70 & ~n37896;
  assign n37898 = ~pi51 & ~n37897;
  assign n37899 = n2559 & ~n37898;
  assign n37900 = n2921 & ~n37899;
  assign n37901 = n2556 & ~n37900;
  assign n37902 = n2554 & ~n37901;
  assign n37903 = ~n6150 & ~n37902;
  assign n37904 = ~pi95 & ~n37903;
  assign n37905 = n2788 & ~n37904;
  assign n37906 = ~pi39 & ~n37905;
  assign n37907 = ~pi38 & ~n3350;
  assign n37908 = ~n37906 & n37907;
  assign n37909 = ~pi228 & n37908;
  assign n37910 = ~n37895 & ~n37909;
  assign n37911 = ~pi100 & ~n37910;
  assign n37912 = ~n13914 & ~n37895;
  assign n37913 = pi100 & ~n37912;
  assign n37914 = ~pi87 & ~n37913;
  assign n37915 = ~n37911 & n37914;
  assign n37916 = pi87 & ~n37895;
  assign n37917 = ~n7323 & n37916;
  assign n37918 = ~pi75 & ~n37917;
  assign n37919 = ~n37915 & n37918;
  assign n37920 = ~n13922 & ~n37895;
  assign n37921 = pi75 & ~n37920;
  assign n37922 = ~pi92 & ~n37921;
  assign n37923 = ~n37919 & n37922;
  assign n37924 = pi92 & ~n37895;
  assign n37925 = ~n7349 & n37924;
  assign n37926 = ~n37923 & ~n37925;
  assign n37927 = ~pi54 & ~n37926;
  assign n37928 = pi54 & ~n37895;
  assign n37929 = ~pi74 & ~n37928;
  assign n37930 = ~n37927 & n37929;
  assign n37931 = ~n7358 & ~n37895;
  assign n37932 = pi74 & ~n37931;
  assign n37933 = ~pi55 & ~n37932;
  assign n37934 = ~n37930 & n37933;
  assign n37935 = pi55 & ~n37895;
  assign n37936 = ~pi56 & ~n37935;
  assign n37937 = ~n37934 & n37936;
  assign n37938 = ~n7364 & ~n37895;
  assign n37939 = pi56 & ~n37938;
  assign n37940 = ~pi62 & ~n37939;
  assign n37941 = ~n37937 & n37940;
  assign n37942 = pi62 & ~n37895;
  assign n37943 = ~n7324 & n37942;
  assign n37944 = ~n37941 & ~n37943;
  assign n37945 = n3429 & ~n37944;
  assign n37946 = ~n3429 & ~n37895;
  assign po383 = ~n37945 & ~n37946;
  assign n37948 = n2497 & n6337;
  assign n37949 = n2532 & n10972;
  assign n37950 = n10970 & n37949;
  assign n37951 = ~pi91 & ~n2570;
  assign n37952 = ~n6257 & n10962;
  assign n37953 = n37951 & ~n37952;
  assign n37954 = ~n37950 & n37953;
  assign n37955 = n37948 & ~n37954;
  assign n37956 = ~pi72 & ~n37955;
  assign n37957 = n6361 & ~n37956;
  assign n37958 = pi829 & ~n6173;
  assign n37959 = ~n37957 & n37958;
  assign n37960 = n13008 & ~n13033;
  assign n37961 = n6361 & n37960;
  assign n37962 = ~n6450 & ~n37961;
  assign n37963 = pi1093 & ~n37962;
  assign n37964 = n10962 & n37948;
  assign n37965 = ~n7474 & n37964;
  assign n37966 = n37948 & ~n37951;
  assign n37967 = ~pi72 & ~n37966;
  assign n37968 = ~n8863 & n37967;
  assign n37969 = ~n37965 & n37968;
  assign n37970 = n6361 & ~n37969;
  assign n37971 = ~n37963 & ~n37970;
  assign n37972 = ~n37964 & n37967;
  assign n37973 = n6361 & ~n37972;
  assign n37974 = n10019 & ~n37973;
  assign n37975 = ~n37971 & ~n37974;
  assign n37976 = ~n37959 & n37975;
  assign n37977 = ~pi39 & ~n37976;
  assign po384 = ~n11408 | n37977;
  assign n37979 = ~pi39 & pi228;
  assign n37980 = ~n11357 & ~n11362;
  assign n37981 = pi39 & ~n37980;
  assign n37982 = n6446 & n37981;
  assign n37983 = ~n8864 & ~n10018;
  assign n37984 = ~pi32 & n10181;
  assign n37985 = ~n37983 & n37984;
  assign n37986 = n2541 & n37985;
  assign n37987 = ~n11424 & n37986;
  assign n37988 = ~n37982 & ~n37987;
  assign n37989 = n10146 & ~n37988;
  assign po385 = n37979 | n37989;
  assign n37991 = ~n6110 & n10143;
  assign n37992 = pi824 & ~n17005;
  assign n37993 = pi829 & pi1091;
  assign n37994 = n17009 & n37993;
  assign n37995 = ~pi824 & ~n37994;
  assign n37996 = n37993 & n37995;
  assign n37997 = ~n37992 & ~n37996;
  assign n37998 = n6257 & ~n6442;
  assign n37999 = ~n37997 & n37998;
  assign n38000 = ~n6143 & ~n6442;
  assign n38001 = ~n6442 & ~n37995;
  assign n38002 = ~n37992 & n38001;
  assign n38003 = ~n16972 & ~n38002;
  assign n38004 = ~n38000 & ~n38003;
  assign n38005 = ~n37999 & n38004;
  assign n38006 = ~n7474 & n16972;
  assign n38007 = ~n16989 & ~n38006;
  assign n38008 = n38000 & ~n38007;
  assign n38009 = pi1093 & ~n38008;
  assign n38010 = ~n38005 & n38009;
  assign n38011 = ~n6258 & n16972;
  assign n38012 = n6144 & n16960;
  assign n38013 = ~n16962 & n38012;
  assign n38014 = ~pi40 & ~n38013;
  assign n38015 = n10227 & ~n38014;
  assign n38016 = pi252 & ~n38015;
  assign n38017 = n6258 & ~n16959;
  assign n38018 = ~n38016 & n38017;
  assign n38019 = ~pi1093 & ~n38018;
  assign n38020 = ~n38011 & n38019;
  assign n38021 = ~pi39 & ~n38020;
  assign n38022 = ~n38010 & n38021;
  assign n38023 = ~n6198 & n16517;
  assign n38024 = ~n6171 & n7473;
  assign n38025 = n16514 & ~n38024;
  assign n38026 = n16603 & n38024;
  assign n38027 = pi1091 & ~n38026;
  assign n38028 = ~n38025 & n38027;
  assign n38029 = ~n6438 & n16514;
  assign n38030 = n6438 & n16603;
  assign n38031 = ~pi1091 & ~n38030;
  assign n38032 = ~n38029 & n38031;
  assign n38033 = ~n38028 & ~n38032;
  assign n38034 = ~pi120 & ~n38033;
  assign n38035 = ~n16516 & ~n38034;
  assign n38036 = n6198 & n38035;
  assign n38037 = ~n38023 & ~n38036;
  assign n38038 = n6215 & n38037;
  assign n38039 = ~n6192 & n38035;
  assign n38040 = ~n35500 & ~n38039;
  assign n38041 = ~n6215 & n38040;
  assign n38042 = ~n3052 & ~n38041;
  assign n38043 = ~n38038 & n38042;
  assign n38044 = n3052 & n16517;
  assign n38045 = ~pi223 & ~n38044;
  assign n38046 = ~n38043 & n38045;
  assign n38047 = pi120 & n6176;
  assign n38048 = n16517 & ~n38047;
  assign n38049 = ~n38023 & ~n38048;
  assign n38050 = n6215 & ~n38049;
  assign n38051 = ~n35500 & ~n38048;
  assign n38052 = ~n6215 & ~n38051;
  assign n38053 = pi223 & ~n38052;
  assign n38054 = ~n38050 & n38053;
  assign n38055 = ~pi299 & ~n38054;
  assign n38056 = ~n38046 & n38055;
  assign n38057 = n6189 & n38037;
  assign n38058 = ~n6189 & n38040;
  assign n38059 = ~n3329 & ~n38058;
  assign n38060 = ~n38057 & n38059;
  assign n38061 = ~pi215 & ~n17254;
  assign n38062 = ~n38060 & n38061;
  assign n38063 = n6189 & ~n38049;
  assign n38064 = ~n6189 & ~n38051;
  assign n38065 = pi215 & ~n38064;
  assign n38066 = ~n38063 & n38065;
  assign n38067 = pi299 & ~n38066;
  assign n38068 = ~n38062 & n38067;
  assign n38069 = ~n38056 & ~n38068;
  assign n38070 = pi39 & ~n38069;
  assign n38071 = ~pi38 & ~n38070;
  assign n38072 = ~n38022 & n38071;
  assign po387 = n37991 & ~n38072;
  assign n38074 = ~pi81 & ~n2675;
  assign n38075 = n6322 & ~n38074;
  assign n38076 = n2451 & ~n38075;
  assign n38077 = n2683 & ~n38076;
  assign n38078 = n2594 & ~n38077;
  assign n38079 = n2687 & ~n38078;
  assign n38080 = n2504 & ~n38079;
  assign n38081 = ~n2507 & ~n38080;
  assign n38082 = ~pi86 & ~n38081;
  assign n38083 = n2592 & ~n38082;
  assign n38084 = n2590 & ~n38083;
  assign n38085 = ~n2585 & ~n38084;
  assign n38086 = ~pi108 & ~n38085;
  assign n38087 = n2584 & ~n38086;
  assign n38088 = n2699 & ~n38087;
  assign n38089 = ~n2575 & ~n38088;
  assign n38090 = n2574 & ~n38089;
  assign n38091 = n2573 & ~n38090;
  assign n38092 = n2566 & ~n38091;
  assign n38093 = n2852 & ~n38092;
  assign n38094 = n2547 & ~n38093;
  assign n38095 = n15510 & ~n38094;
  assign n38096 = ~pi70 & ~n38095;
  assign n38097 = ~n2843 & ~n38096;
  assign n38098 = ~pi51 & ~n38097;
  assign n38099 = n2559 & ~n38098;
  assign n38100 = n2921 & ~n38099;
  assign n38101 = n2556 & ~n38100;
  assign n38102 = ~pi1082 & n2553;
  assign n38103 = ~pi32 & ~n38102;
  assign n38104 = ~n38101 & n38103;
  assign n38105 = ~n3360 & ~n38104;
  assign n38106 = ~pi95 & ~n38105;
  assign n38107 = ~n2727 & ~n38106;
  assign n38108 = ~pi39 & ~n38107;
  assign n38109 = ~n7274 & ~n7276;
  assign po950 = ~n6175 | ~n6257;
  assign n38111 = n6436 & ~po950;
  assign n38112 = ~n38109 & n38111;
  assign n38113 = n6167 & n11307;
  assign n38114 = ~n38112 & n38113;
  assign n38115 = ~n3350 & ~n38114;
  assign n38116 = ~n38108 & n38115;
  assign n38117 = ~pi38 & ~n38116;
  assign n38118 = n6111 & ~n38117;
  assign n38119 = ~pi87 & ~n6236;
  assign n38120 = ~n38118 & n38119;
  assign n38121 = ~n6269 & ~n38120;
  assign n38122 = n3237 & ~n38121;
  assign n38123 = n7273 & ~n38122;
  assign n38124 = ~pi54 & ~n38123;
  assign n38125 = ~n7308 & ~n38124;
  assign n38126 = n8839 & ~n38125;
  assign n38127 = n15599 & ~n38126;
  assign n38128 = ~pi56 & ~n38127;
  assign n38129 = ~n6104 & ~n38128;
  assign n38130 = ~pi62 & ~n38129;
  assign n38131 = ~n6280 & ~n38130;
  assign n38132 = n3429 & ~n38131;
  assign po389 = n6100 & ~n38132;
  assign n38134 = ~pi230 & ~pi233;
  assign n38135 = ~pi212 & ~pi214;
  assign n38136 = ~pi211 & ~n38135;
  assign n38137 = pi219 & ~n38136;
  assign n38138 = po1038 & ~n38137;
  assign n38139 = pi1142 & ~n10428;
  assign n38140 = pi211 & pi1143;
  assign n38141 = ~pi211 & pi1144;
  assign n38142 = ~n38140 & ~n38141;
  assign n38143 = ~pi212 & pi214;
  assign n38144 = pi212 & ~pi214;
  assign n38145 = ~n38143 & ~n38144;
  assign n38146 = ~n38142 & ~n38145;
  assign n38147 = ~pi211 & pi1143;
  assign n38148 = n10669 & n38147;
  assign n38149 = ~n38146 & ~n38148;
  assign n38150 = ~pi219 & ~n38149;
  assign n38151 = ~n38139 & ~n38150;
  assign n38152 = n38138 & ~n38151;
  assign n38153 = pi299 & ~n38142;
  assign n38154 = pi199 & pi1142;
  assign n38155 = ~pi200 & ~n38154;
  assign n38156 = ~pi199 & pi1144;
  assign n38157 = n38155 & ~n38156;
  assign n38158 = ~pi199 & pi1143;
  assign n38159 = pi200 & ~n38158;
  assign n38160 = ~n38157 & ~n38159;
  assign n38161 = ~pi299 & ~n38160;
  assign n38162 = ~pi207 & ~n38161;
  assign n38163 = n38155 & ~n38158;
  assign n38164 = pi207 & ~pi299;
  assign n38165 = ~pi199 & pi1142;
  assign n38166 = pi200 & ~n38165;
  assign n38167 = n38164 & ~n38166;
  assign n38168 = ~n38163 & n38167;
  assign n38169 = ~n38162 & ~n38168;
  assign n38170 = pi208 & ~n38169;
  assign n38171 = pi207 & ~pi208;
  assign n38172 = n38160 & n38171;
  assign n38173 = ~n38170 & ~n38172;
  assign n38174 = ~pi299 & ~n38173;
  assign n38175 = ~n38153 & ~n38174;
  assign n38176 = ~pi214 & ~n38174;
  assign n38177 = ~pi212 & ~n38176;
  assign n38178 = ~n38175 & n38177;
  assign n38179 = ~n38153 & n38176;
  assign n38180 = pi211 & pi1142;
  assign n38181 = ~n38147 & ~n38180;
  assign n38182 = pi299 & ~n38181;
  assign n38183 = pi214 & ~n38182;
  assign n38184 = ~n38174 & n38183;
  assign n38185 = pi212 & ~n38184;
  assign n38186 = ~n38179 & n38185;
  assign n38187 = ~pi219 & ~n38186;
  assign n38188 = ~n38178 & n38187;
  assign n38189 = ~pi299 & n38173;
  assign n38190 = pi299 & ~pi1142;
  assign n38191 = n38136 & ~n38190;
  assign n38192 = ~n38189 & n38191;
  assign n38193 = ~n38136 & n38174;
  assign n38194 = pi219 & ~n38193;
  assign n38195 = ~n38192 & n38194;
  assign n38196 = ~po1038 & ~n38195;
  assign n38197 = ~n38188 & n38196;
  assign n38198 = ~n38152 & ~n38197;
  assign n38199 = pi213 & n38198;
  assign n38200 = ~pi211 & pi1156;
  assign n38201 = pi211 & pi1155;
  assign n38202 = ~n38200 & ~n38201;
  assign n38203 = ~pi214 & ~n38202;
  assign n38204 = ~pi211 & pi1155;
  assign n38205 = pi211 & pi1154;
  assign n38206 = ~n38204 & ~n38205;
  assign n38207 = pi214 & ~n38206;
  assign n38208 = ~n38203 & ~n38207;
  assign n38209 = pi212 & ~n38208;
  assign n38210 = ~pi211 & pi1157;
  assign n38211 = pi211 & pi1156;
  assign n38212 = ~n38210 & ~n38211;
  assign n38213 = pi214 & ~n38212;
  assign n38214 = ~pi212 & n38213;
  assign n38215 = ~n38209 & ~n38214;
  assign n38216 = ~pi219 & n38215;
  assign n38217 = ~pi211 & pi214;
  assign n38218 = pi1155 & n38217;
  assign n38219 = ~pi212 & ~n38218;
  assign n38220 = ~pi211 & pi1154;
  assign n38221 = ~pi214 & ~n38220;
  assign n38222 = ~pi211 & pi1153;
  assign n38223 = n10669 & ~n38222;
  assign n38224 = ~n38221 & ~n38223;
  assign n38225 = ~n38219 & n38224;
  assign n38226 = pi219 & ~n38225;
  assign n38227 = po1038 & ~n38226;
  assign n38228 = ~n38216 & n38227;
  assign n38229 = ~pi213 & ~n38228;
  assign n38230 = ~pi219 & pi299;
  assign n38231 = ~n38215 & n38230;
  assign n38232 = pi299 & pi1155;
  assign n38233 = n38143 & n38232;
  assign n38234 = pi299 & pi1154;
  assign n38235 = ~pi214 & ~n38234;
  assign n38236 = pi299 & pi1153;
  assign n38237 = pi214 & ~n38236;
  assign n38238 = pi212 & ~n38237;
  assign n38239 = ~n38235 & n38238;
  assign n38240 = ~n38233 & ~n38239;
  assign n38241 = ~pi211 & pi219;
  assign n38242 = ~n38240 & n38241;
  assign n38243 = ~n38231 & ~n38242;
  assign n38244 = ~n38174 & n38243;
  assign n38245 = ~po1038 & ~n38244;
  assign n38246 = n38229 & ~n38245;
  assign n38247 = pi209 & ~n38246;
  assign n38248 = ~n38199 & n38247;
  assign n38249 = ~pi200 & pi1155;
  assign n38250 = pi199 & n38249;
  assign n38251 = ~pi299 & n38250;
  assign n38252 = ~pi1156 & ~n38251;
  assign n38253 = ~pi200 & ~pi1155;
  assign n38254 = pi199 & pi200;
  assign n38255 = ~n10758 & ~n38254;
  assign n38256 = ~pi299 & n38255;
  assign n38257 = ~n38253 & n38256;
  assign n38258 = ~n38252 & n38257;
  assign n38259 = pi207 & n38258;
  assign n38260 = ~pi208 & ~n38259;
  assign n38261 = ~pi299 & ~n38254;
  assign n38262 = pi1153 & ~n38261;
  assign n38263 = pi1154 & ~n38262;
  assign n38264 = n11311 & n38249;
  assign n38265 = ~pi1153 & ~n11311;
  assign n38266 = pi1154 & n38255;
  assign n38267 = ~n38265 & n38266;
  assign n38268 = ~n38264 & ~n38267;
  assign n38269 = n38263 & ~n38268;
  assign n38270 = ~pi200 & ~pi299;
  assign n38271 = pi199 & ~pi1153;
  assign n38272 = n38270 & ~n38271;
  assign n38273 = ~pi199 & ~pi1155;
  assign n38274 = ~pi1154 & ~n38273;
  assign n38275 = n38272 & n38274;
  assign n38276 = ~n38269 & ~n38275;
  assign n38277 = pi207 & n38276;
  assign n38278 = pi200 & ~pi299;
  assign n38279 = ~pi199 & pi1155;
  assign n38280 = n38278 & n38279;
  assign n38281 = ~pi1154 & ~n38280;
  assign n38282 = pi200 & ~n38279;
  assign n38283 = n10761 & ~n38282;
  assign n38284 = ~n38281 & n38283;
  assign n38285 = pi200 & ~pi1155;
  assign n38286 = n11311 & ~n38285;
  assign n38287 = pi1156 & n38286;
  assign n38288 = ~n38284 & ~n38287;
  assign n38289 = ~n10564 & n38288;
  assign n38290 = ~n38277 & ~n38289;
  assign n38291 = pi208 & ~n38290;
  assign n38292 = ~n38260 & ~n38291;
  assign n38293 = ~pi1157 & ~n38292;
  assign n38294 = pi199 & ~pi1155;
  assign n38295 = pi1156 & ~n38294;
  assign n38296 = n38261 & n38295;
  assign n38297 = ~pi1156 & ~n38294;
  assign n38298 = n38270 & n38297;
  assign n38299 = ~n38296 & ~n38298;
  assign n38300 = pi207 & ~n38299;
  assign n38301 = ~pi208 & ~n38300;
  assign n38302 = ~n38291 & ~n38301;
  assign n38303 = pi1157 & ~n38302;
  assign n38304 = ~n38293 & ~n38303;
  assign n38305 = pi211 & ~n38304;
  assign n38306 = ~pi214 & ~n38304;
  assign n38307 = ~pi212 & ~n38306;
  assign n38308 = pi1155 & ~n11321;
  assign n38309 = n38256 & ~n38271;
  assign n38310 = ~n38308 & ~n38309;
  assign n38311 = ~pi1154 & n38278;
  assign n38312 = ~n38310 & ~n38311;
  assign n38313 = pi207 & ~n38312;
  assign n38314 = ~pi207 & ~n38232;
  assign n38315 = n38288 & n38314;
  assign n38316 = pi208 & ~n38315;
  assign n38317 = ~n38313 & n38316;
  assign n38318 = ~pi208 & ~n38314;
  assign n38319 = ~pi299 & n38252;
  assign n38320 = ~pi299 & ~n38255;
  assign n38321 = ~pi1155 & ~n11311;
  assign n38322 = ~n38320 & ~n38321;
  assign n38323 = ~n38319 & n38322;
  assign n38324 = n38318 & n38323;
  assign n38325 = pi1155 & ~n38278;
  assign n38326 = ~n11311 & ~n38325;
  assign n38327 = pi1156 & ~n38326;
  assign n38328 = pi199 & ~pi200;
  assign n38329 = ~pi299 & ~n38328;
  assign n38330 = ~pi1155 & ~n38329;
  assign n38331 = ~pi1156 & ~n38278;
  assign n38332 = ~n38330 & n38331;
  assign n38333 = ~n38327 & ~n38332;
  assign n38334 = pi1157 & n38318;
  assign n38335 = ~n38333 & n38334;
  assign n38336 = ~n38324 & ~n38335;
  assign n38337 = ~n38317 & n38336;
  assign n38338 = n38217 & n38337;
  assign n38339 = n38307 & ~n38338;
  assign n38340 = ~pi1155 & ~n10761;
  assign n38341 = ~n38325 & ~n38340;
  assign n38342 = n11321 & ~n38249;
  assign n38343 = pi1156 & ~n38342;
  assign n38344 = n38341 & ~n38343;
  assign n38345 = pi207 & n38344;
  assign n38346 = ~pi207 & ~pi299;
  assign n38347 = ~pi208 & ~n38346;
  assign n38348 = ~n38345 & n38347;
  assign n38349 = pi1157 & ~n38348;
  assign n38350 = ~pi299 & ~n11381;
  assign n38351 = pi1156 & ~n38250;
  assign n38352 = n38350 & n38351;
  assign n38353 = ~n38252 & ~n38352;
  assign n38354 = ~pi299 & ~n38353;
  assign n38355 = n38347 & ~n38354;
  assign n38356 = ~pi1157 & ~n38355;
  assign n38357 = pi299 & ~pi1153;
  assign n38358 = ~n38356 & ~n38357;
  assign n38359 = ~n38349 & n38358;
  assign n38360 = pi1153 & ~n38329;
  assign n38361 = n38268 & ~n38360;
  assign n38362 = pi207 & ~n38361;
  assign n38363 = ~n38308 & ~n38340;
  assign n38364 = pi1156 & ~n38363;
  assign n38365 = pi1155 & ~n38320;
  assign n38366 = ~n38330 & ~n38365;
  assign n38367 = pi1154 & ~n38366;
  assign n38368 = ~n38364 & ~n38367;
  assign n38369 = pi299 & ~pi1155;
  assign n38370 = pi1155 & ~n38350;
  assign n38371 = ~n38369 & ~n38370;
  assign n38372 = n38368 & n38371;
  assign n38373 = ~pi207 & ~n38357;
  assign n38374 = ~n38372 & n38373;
  assign n38375 = ~n38362 & ~n38374;
  assign n38376 = pi208 & ~n38375;
  assign n38377 = n38217 & ~n38376;
  assign n38378 = ~n38359 & n38377;
  assign n38379 = ~pi211 & ~pi214;
  assign n38380 = n38288 & ~n38367;
  assign n38381 = ~pi207 & ~n38380;
  assign n38382 = ~pi299 & n38310;
  assign n38383 = pi1154 & ~n38382;
  assign n38384 = ~n38275 & ~n38383;
  assign n38385 = pi207 & ~n38384;
  assign n38386 = ~n38381 & ~n38385;
  assign n38387 = pi208 & ~n38386;
  assign n38388 = pi299 & ~pi1154;
  assign n38389 = pi1157 & ~n38388;
  assign n38390 = ~n38234 & ~n38259;
  assign n38391 = ~pi208 & ~n38390;
  assign n38392 = ~n38389 & ~n38391;
  assign n38393 = ~n38349 & ~n38392;
  assign n38394 = ~n38387 & ~n38393;
  assign n38395 = n38379 & n38394;
  assign n38396 = pi212 & ~n38395;
  assign n38397 = ~n38378 & n38396;
  assign n38398 = ~n38339 & ~n38397;
  assign n38399 = ~n38305 & ~n38398;
  assign n38400 = pi219 & ~n38399;
  assign n38401 = ~pi207 & n38372;
  assign n38402 = n38164 & n38361;
  assign n38403 = pi208 & ~n38402;
  assign n38404 = ~n38401 & n38403;
  assign n38405 = n38349 & ~n38404;
  assign n38406 = ~pi211 & ~n38405;
  assign n38407 = ~n38293 & n38406;
  assign n38408 = pi207 & ~n38276;
  assign n38409 = ~n38284 & ~n38364;
  assign n38410 = ~n38164 & ~n38409;
  assign n38411 = ~n38408 & ~n38410;
  assign n38412 = pi208 & ~n38411;
  assign n38413 = ~n38252 & n38355;
  assign n38414 = ~pi208 & pi1157;
  assign n38415 = pi299 & pi1156;
  assign n38416 = ~n38300 & ~n38415;
  assign n38417 = n38414 & ~n38416;
  assign n38418 = ~n38413 & ~n38417;
  assign n38419 = ~n38412 & n38418;
  assign n38420 = pi211 & ~n38419;
  assign n38421 = pi214 & ~n38420;
  assign n38422 = ~n38407 & n38421;
  assign n38423 = n38307 & ~n38422;
  assign n38424 = n10426 & ~n38394;
  assign n38425 = ~n10426 & ~n38379;
  assign n38426 = ~n38337 & n38425;
  assign n38427 = n38379 & ~n38419;
  assign n38428 = ~n38426 & ~n38427;
  assign n38429 = ~n38424 & n38428;
  assign n38430 = pi212 & ~n38429;
  assign n38431 = ~pi219 & ~n38430;
  assign n38432 = ~n38423 & n38431;
  assign n38433 = ~po1038 & ~n38432;
  assign n38434 = ~n38400 & n38433;
  assign n38435 = n38229 & ~n38434;
  assign n38436 = ~pi211 & n10669;
  assign n38437 = pi299 & pi1143;
  assign n38438 = ~pi299 & ~n38409;
  assign n38439 = ~n38437 & ~n38438;
  assign n38440 = ~pi207 & n38439;
  assign n38441 = n38277 & ~n38437;
  assign n38442 = pi208 & ~n38441;
  assign n38443 = ~n38440 & n38442;
  assign n38444 = pi299 & ~pi1143;
  assign n38445 = ~pi1157 & n38355;
  assign n38446 = ~n38444 & n38445;
  assign n38447 = ~n38296 & n38341;
  assign n38448 = ~n38346 & ~n38444;
  assign n38449 = ~n38447 & n38448;
  assign n38450 = n38414 & n38449;
  assign n38451 = ~n38446 & ~n38450;
  assign n38452 = ~n38443 & n38451;
  assign n38453 = n38436 & n38452;
  assign n38454 = pi299 & pi1144;
  assign n38455 = ~n38438 & ~n38454;
  assign n38456 = ~pi207 & n38455;
  assign n38457 = n38277 & ~n38454;
  assign n38458 = pi208 & ~n38457;
  assign n38459 = ~n38456 & n38458;
  assign n38460 = pi299 & ~pi1144;
  assign n38461 = n38445 & ~n38460;
  assign n38462 = ~n38346 & ~n38460;
  assign n38463 = ~n38447 & n38462;
  assign n38464 = n38414 & n38463;
  assign n38465 = ~n38461 & ~n38464;
  assign n38466 = ~n38459 & n38465;
  assign n38467 = ~pi211 & ~n38466;
  assign n38468 = ~n10669 & ~n38135;
  assign n38469 = pi211 & ~n38452;
  assign n38470 = n38468 & ~n38469;
  assign n38471 = ~n38467 & n38470;
  assign n38472 = ~n38453 & ~n38471;
  assign n38473 = ~pi219 & ~n38472;
  assign n38474 = ~pi219 & ~n38135;
  assign n38475 = ~n38136 & ~n38474;
  assign n38476 = ~n38304 & n38475;
  assign n38477 = ~pi299 & n38312;
  assign n38478 = pi299 & pi1142;
  assign n38479 = pi207 & ~n38478;
  assign n38480 = ~n38477 & n38479;
  assign n38481 = ~pi207 & ~n38478;
  assign n38482 = ~n38438 & n38481;
  assign n38483 = pi208 & ~n38482;
  assign n38484 = ~n38480 & n38483;
  assign n38485 = ~n38190 & ~n38356;
  assign n38486 = ~n38349 & n38485;
  assign n38487 = ~n10428 & ~n38475;
  assign n38488 = ~n38486 & n38487;
  assign n38489 = ~n38484 & n38488;
  assign n38490 = ~po1038 & ~n38489;
  assign n38491 = ~n38476 & n38490;
  assign n38492 = ~n38473 & n38491;
  assign n38493 = pi213 & ~n38152;
  assign n38494 = ~n38492 & n38493;
  assign n38495 = ~pi209 & ~n38494;
  assign n38496 = ~n38435 & n38495;
  assign n38497 = ~n38248 & ~n38496;
  assign n38498 = pi230 & ~n38497;
  assign po390 = n38134 | n38498;
  assign n38500 = pi1153 & ~n38379;
  assign n38501 = ~n38217 & ~n38221;
  assign n38502 = ~n38500 & ~n38501;
  assign n38503 = pi212 & ~n38502;
  assign n38504 = pi211 & pi1153;
  assign n38505 = ~n38220 & ~n38504;
  assign n38506 = n38143 & ~n38505;
  assign n38507 = ~pi219 & ~n38506;
  assign n38508 = ~n38503 & n38507;
  assign n38509 = n38138 & ~n38508;
  assign n38510 = pi1152 & ~n38509;
  assign n38511 = ~pi207 & ~pi208;
  assign n38512 = ~n10564 & ~n38511;
  assign n38513 = ~pi1154 & ~n38264;
  assign n38514 = ~pi199 & n38253;
  assign n38515 = n38261 & ~n38514;
  assign n38516 = ~n38513 & n38515;
  assign n38517 = pi207 & n38516;
  assign n38518 = ~n38512 & ~n38517;
  assign n38519 = ~n38289 & ~n38518;
  assign n38520 = ~pi214 & ~n38519;
  assign n38521 = ~pi212 & ~n38520;
  assign n38522 = ~pi207 & n38234;
  assign n38523 = pi207 & ~n38380;
  assign n38524 = ~n38522 & ~n38523;
  assign n38525 = ~pi208 & ~n38524;
  assign n38526 = ~pi1155 & n10758;
  assign n38527 = ~n38254 & ~n38526;
  assign n38528 = ~pi299 & ~n38527;
  assign n38529 = ~n38513 & ~n38528;
  assign n38530 = pi207 & n38529;
  assign n38531 = ~n38381 & ~n38530;
  assign n38532 = pi208 & ~n38531;
  assign n38533 = ~n38525 & ~n38532;
  assign n38534 = ~pi211 & ~n38533;
  assign n38535 = pi207 & n38371;
  assign n38536 = n38368 & n38535;
  assign n38537 = n38347 & ~n38536;
  assign n38538 = n38164 & ~n38529;
  assign n38539 = pi208 & ~n38538;
  assign n38540 = ~n38401 & n38539;
  assign n38541 = ~n38537 & ~n38540;
  assign n38542 = ~n38357 & ~n38541;
  assign n38543 = pi211 & n38542;
  assign n38544 = ~n38534 & ~n38543;
  assign n38545 = pi214 & n38544;
  assign n38546 = n38521 & ~n38545;
  assign n38547 = ~pi219 & ~n38546;
  assign n38548 = ~pi214 & ~n38544;
  assign n38549 = ~pi211 & ~n38542;
  assign n38550 = pi214 & ~n38549;
  assign n38551 = ~n38541 & n38550;
  assign n38552 = ~n38548 & ~n38551;
  assign n38553 = pi212 & ~n38552;
  assign n38554 = n38547 & ~n38553;
  assign n38555 = ~n38136 & n38519;
  assign n38556 = pi219 & ~n38555;
  assign n38557 = n38136 & ~n38541;
  assign n38558 = n38556 & ~n38557;
  assign n38559 = ~po1038 & ~n38558;
  assign n38560 = ~n38554 & n38559;
  assign n38561 = n38510 & ~n38560;
  assign n38562 = ~n10669 & n38505;
  assign n38563 = n38474 & ~n38562;
  assign n38564 = ~n38223 & n38563;
  assign n38565 = po1038 & n38564;
  assign n38566 = ~pi1152 & ~n38565;
  assign n38567 = pi211 & ~n38519;
  assign n38568 = n38550 & ~n38567;
  assign n38569 = ~n38548 & ~n38568;
  assign n38570 = pi212 & ~n38569;
  assign n38571 = n38547 & ~n38570;
  assign n38572 = pi219 & ~n38519;
  assign n38573 = ~po1038 & ~n38572;
  assign n38574 = ~n38571 & n38573;
  assign n38575 = n38566 & ~n38574;
  assign n38576 = ~pi213 & ~n38575;
  assign n38577 = ~n38561 & n38576;
  assign n38578 = ~n38410 & ~n38517;
  assign n38579 = pi208 & ~n38578;
  assign n38580 = n38347 & ~n38409;
  assign n38581 = ~n38579 & ~n38580;
  assign n38582 = ~pi211 & ~n38581;
  assign n38583 = ~n38232 & ~n38519;
  assign n38584 = pi211 & ~n38583;
  assign n38585 = ~n38582 & ~n38584;
  assign n38586 = ~pi214 & n38585;
  assign n38587 = pi211 & ~n38533;
  assign n38588 = ~pi211 & ~n38583;
  assign n38589 = pi214 & ~n38588;
  assign n38590 = ~n38587 & n38589;
  assign n38591 = pi212 & ~n38590;
  assign n38592 = ~n38586 & n38591;
  assign n38593 = pi214 & n38585;
  assign n38594 = n38521 & ~n38593;
  assign n38595 = ~pi219 & ~n38594;
  assign n38596 = ~n38592 & n38595;
  assign n38597 = ~n38135 & n38534;
  assign n38598 = n38556 & ~n38597;
  assign n38599 = n35599 & ~n38598;
  assign n38600 = ~n38596 & n38599;
  assign n38601 = pi209 & ~n38600;
  assign n38602 = ~n38577 & n38601;
  assign n38603 = ~pi199 & pi1153;
  assign n38604 = pi200 & n38603;
  assign n38605 = ~pi299 & n38604;
  assign n38606 = pi1154 & ~n38278;
  assign n38607 = ~n38605 & ~n38606;
  assign n38608 = n38329 & n38607;
  assign n38609 = n38347 & ~n38608;
  assign n38610 = ~pi207 & n38608;
  assign n38611 = ~pi200 & ~pi1153;
  assign n38612 = ~pi199 & ~n38611;
  assign n38613 = ~pi299 & ~n38612;
  assign n38614 = ~n38328 & n38613;
  assign n38615 = pi207 & n38614;
  assign n38616 = pi208 & ~n38615;
  assign n38617 = ~n38610 & n38616;
  assign n38618 = ~n38609 & ~n38617;
  assign n38619 = ~pi211 & n38618;
  assign n38620 = ~pi299 & n10758;
  assign n38621 = ~pi1153 & ~n38620;
  assign n38622 = n38263 & ~n38621;
  assign n38623 = ~pi199 & ~pi1153;
  assign n38624 = n38256 & ~n38623;
  assign n38625 = ~n38622 & ~n38624;
  assign n38626 = ~n10564 & n38625;
  assign n38627 = ~pi1153 & n10758;
  assign n38628 = n38261 & ~n38627;
  assign n38629 = n10564 & ~n38628;
  assign n38630 = ~n38511 & ~n38629;
  assign n38631 = ~n38626 & n38630;
  assign n38632 = pi211 & ~n38631;
  assign n38633 = ~n38619 & ~n38632;
  assign n38634 = ~n38135 & n38633;
  assign n38635 = pi219 & ~n38135;
  assign n38636 = pi219 & ~n38631;
  assign n38637 = ~n38635 & ~n38636;
  assign n38638 = ~n38634 & ~n38637;
  assign n38639 = ~po1038 & ~n38638;
  assign n38640 = ~pi214 & ~n38631;
  assign n38641 = ~pi212 & ~n38640;
  assign n38642 = ~n38234 & ~n38631;
  assign n38643 = ~pi211 & ~n38642;
  assign n38644 = ~pi1153 & ~n38270;
  assign n38645 = ~n38320 & ~n38644;
  assign n38646 = pi1154 & ~n11321;
  assign n38647 = ~n38644 & n38646;
  assign n38648 = ~n38645 & ~n38647;
  assign n38649 = ~pi207 & ~n38648;
  assign n38650 = ~pi1153 & ~n10761;
  assign n38651 = ~pi299 & n38254;
  assign n38652 = pi207 & ~n38651;
  assign n38653 = ~n38650 & n38652;
  assign n38654 = ~n38649 & ~n38653;
  assign n38655 = pi208 & ~n38654;
  assign n38656 = n38347 & ~n38648;
  assign n38657 = ~n38655 & ~n38656;
  assign n38658 = pi211 & ~n38657;
  assign n38659 = ~n38643 & ~n38658;
  assign n38660 = pi214 & n38659;
  assign n38661 = n38641 & ~n38660;
  assign n38662 = ~pi214 & n38659;
  assign n38663 = pi211 & ~n38618;
  assign n38664 = ~pi211 & ~n38657;
  assign n38665 = pi214 & ~n38664;
  assign n38666 = ~n38663 & n38665;
  assign n38667 = pi212 & ~n38666;
  assign n38668 = ~n38662 & n38667;
  assign n38669 = ~pi219 & ~n38668;
  assign n38670 = ~n38661 & n38669;
  assign n38671 = n38639 & ~n38670;
  assign n38672 = n38510 & ~n38671;
  assign n38673 = pi1153 & ~pi1154;
  assign n38674 = ~n38350 & n38673;
  assign n38675 = ~n38647 & ~n38674;
  assign n38676 = n38347 & ~n38675;
  assign n38677 = pi207 & ~n10761;
  assign n38678 = pi1153 & n38677;
  assign n38679 = n38164 & ~n38678;
  assign n38680 = pi208 & ~n38679;
  assign n38681 = n38675 & ~n38678;
  assign n38682 = n38680 & ~n38681;
  assign n38683 = ~n38676 & ~n38682;
  assign n38684 = n38436 & n38683;
  assign n38685 = pi1154 & ~n10761;
  assign n38686 = ~n38605 & ~n38685;
  assign n38687 = ~pi299 & n38686;
  assign n38688 = pi207 & n38687;
  assign n38689 = n38347 & ~n38688;
  assign n38690 = ~pi207 & n38687;
  assign n38691 = n38680 & ~n38690;
  assign n38692 = ~n38689 & ~n38691;
  assign n38693 = ~n38388 & ~n38690;
  assign n38694 = ~n38692 & n38693;
  assign n38695 = ~pi211 & ~n38694;
  assign n38696 = pi211 & n38683;
  assign n38697 = ~n38695 & ~n38696;
  assign n38698 = n38468 & ~n38697;
  assign n38699 = ~n38684 & ~n38698;
  assign n38700 = ~pi219 & ~n38699;
  assign n38701 = ~pi200 & pi207;
  assign n38702 = ~n38512 & ~n38701;
  assign n38703 = n11311 & ~n38702;
  assign n38704 = ~n38692 & n38703;
  assign n38705 = pi219 & ~n38704;
  assign n38706 = ~po1038 & ~n38705;
  assign n38707 = ~n38217 & ~n38468;
  assign n38708 = ~n38704 & n38707;
  assign n38709 = n38706 & ~n38708;
  assign n38710 = ~n38700 & n38709;
  assign n38711 = n38566 & ~n38710;
  assign n38712 = ~n38672 & ~n38711;
  assign n38713 = ~pi213 & n38712;
  assign n38714 = ~pi1152 & ~po1038;
  assign n38715 = pi211 & ~n38694;
  assign n38716 = ~n38232 & ~n38704;
  assign n38717 = ~pi211 & n38716;
  assign n38718 = n10669 & ~n38717;
  assign n38719 = ~n38715 & n38718;
  assign n38720 = pi211 & n38716;
  assign n38721 = ~pi211 & ~n38415;
  assign n38722 = ~n38704 & n38721;
  assign n38723 = ~n38145 & ~n38722;
  assign n38724 = ~n38720 & n38723;
  assign n38725 = ~n38719 & ~n38724;
  assign n38726 = ~pi219 & ~n38725;
  assign n38727 = n38135 & n38704;
  assign n38728 = pi211 & ~n38704;
  assign n38729 = n38635 & ~n38728;
  assign n38730 = ~n38695 & n38729;
  assign n38731 = ~n38727 & ~n38730;
  assign n38732 = ~n38726 & n38731;
  assign n38733 = n38714 & ~n38732;
  assign n38734 = ~pi212 & n38640;
  assign n38735 = ~n38632 & ~n38642;
  assign n38736 = ~n38734 & n38735;
  assign n38737 = pi219 & n38736;
  assign n38738 = pi211 & ~n38642;
  assign n38739 = ~n38369 & ~n38610;
  assign n38740 = ~n38618 & n38739;
  assign n38741 = ~pi211 & n38740;
  assign n38742 = n10669 & ~n38741;
  assign n38743 = ~n38738 & n38742;
  assign n38744 = pi211 & n38740;
  assign n38745 = ~n38415 & n38625;
  assign n38746 = ~pi207 & ~n38745;
  assign n38747 = pi207 & ~n38614;
  assign n38748 = pi299 & ~pi1156;
  assign n38749 = n38747 & ~n38748;
  assign n38750 = pi208 & ~n38749;
  assign n38751 = ~n38746 & n38750;
  assign n38752 = ~pi208 & ~n38415;
  assign n38753 = ~n38631 & n38752;
  assign n38754 = ~pi211 & ~n38753;
  assign n38755 = ~n38751 & n38754;
  assign n38756 = ~n38145 & ~n38755;
  assign n38757 = ~n38744 & n38756;
  assign n38758 = ~pi219 & ~n38734;
  assign n38759 = ~n38757 & n38758;
  assign n38760 = ~n38743 & n38759;
  assign n38761 = ~n38737 & ~n38760;
  assign n38762 = pi1152 & ~po1038;
  assign n38763 = ~n38761 & n38762;
  assign n38764 = ~n38733 & ~n38763;
  assign n38765 = pi213 & ~n38764;
  assign n38766 = ~pi209 & ~n38765;
  assign n38767 = ~n38713 & n38766;
  assign n38768 = ~n38602 & ~n38767;
  assign n38769 = pi214 & ~n38202;
  assign n38770 = ~pi212 & n38769;
  assign n38771 = ~pi219 & ~n38770;
  assign n38772 = ~n38209 & n38771;
  assign n38773 = pi219 & ~n38220;
  assign n38774 = pi213 & ~n38773;
  assign n38775 = n38138 & n38774;
  assign n38776 = ~n38772 & n38775;
  assign n38777 = ~n38768 & ~n38776;
  assign n38778 = pi230 & ~n38777;
  assign n38779 = ~pi230 & pi234;
  assign po391 = n38778 | n38779;
  assign n38781 = ~pi1156 & n38280;
  assign n38782 = ~n38364 & ~n38781;
  assign n38783 = pi207 & ~n38782;
  assign n38784 = ~pi207 & n38353;
  assign n38785 = ~n38783 & ~n38784;
  assign n38786 = pi208 & ~n38785;
  assign n38787 = ~n38413 & ~n38786;
  assign n38788 = ~pi1157 & ~n38787;
  assign n38789 = pi208 & pi1157;
  assign n38790 = ~n38298 & ~n38343;
  assign n38791 = ~pi207 & ~n38790;
  assign n38792 = ~n38783 & ~n38791;
  assign n38793 = n38789 & ~n38792;
  assign n38794 = ~n38417 & ~n38793;
  assign n38795 = ~n38788 & n38794;
  assign n38796 = ~pi211 & ~n38795;
  assign n38797 = ~n38287 & ~n38370;
  assign n38798 = pi207 & ~n38797;
  assign n38799 = ~pi207 & n38323;
  assign n38800 = ~n38798 & ~n38799;
  assign n38801 = pi208 & ~n38800;
  assign n38802 = ~n38324 & ~n38801;
  assign n38803 = ~pi1157 & ~n38802;
  assign n38804 = ~pi207 & ~n38333;
  assign n38805 = ~n38798 & ~n38804;
  assign n38806 = n38789 & ~n38805;
  assign n38807 = ~n38335 & ~n38806;
  assign n38808 = ~n38803 & n38807;
  assign n38809 = pi211 & ~n38808;
  assign n38810 = n10669 & ~n38809;
  assign n38811 = ~n38796 & n38810;
  assign n38812 = n10564 & ~n38287;
  assign n38813 = ~n38781 & n38812;
  assign n38814 = ~pi207 & ~n38258;
  assign n38815 = ~n38813 & ~n38814;
  assign n38816 = ~n38260 & n38815;
  assign n38817 = ~pi1157 & ~n38816;
  assign n38818 = ~pi207 & n38299;
  assign n38819 = ~n38813 & ~n38818;
  assign n38820 = ~n38301 & n38819;
  assign n38821 = pi1157 & ~n38820;
  assign n38822 = ~n38817 & ~n38821;
  assign n38823 = n38135 & ~n38822;
  assign n38824 = pi211 & ~n38795;
  assign n38825 = ~pi207 & n38344;
  assign n38826 = pi208 & ~n38825;
  assign n38827 = ~n38364 & n38535;
  assign n38828 = n38826 & ~n38827;
  assign n38829 = ~n38348 & ~n38828;
  assign n38830 = pi1157 & n38829;
  assign n38831 = ~pi211 & ~n38817;
  assign n38832 = ~n38830 & n38831;
  assign n38833 = n38468 & ~n38832;
  assign n38834 = ~n38824 & n38833;
  assign n38835 = ~n38823 & ~n38834;
  assign n38836 = ~n38811 & n38835;
  assign n38837 = ~pi219 & ~n38836;
  assign n38838 = ~pi211 & n38808;
  assign n38839 = pi211 & ~n38822;
  assign n38840 = ~n38145 & ~n38839;
  assign n38841 = ~n38838 & n38840;
  assign n38842 = n38145 & n38822;
  assign n38843 = pi219 & ~n38842;
  assign n38844 = ~n38841 & n38843;
  assign n38845 = pi209 & ~n38844;
  assign n38846 = ~n38837 & n38845;
  assign n38847 = ~pi1154 & ~n38605;
  assign n38848 = pi200 & ~pi1153;
  assign n38849 = n11311 & ~n38848;
  assign n38850 = ~n38847 & n38849;
  assign n38851 = n10564 & ~n38850;
  assign n38852 = ~n38276 & ~n38511;
  assign n38853 = ~n10564 & ~n38852;
  assign n38854 = ~n38851 & ~n38853;
  assign n38855 = ~pi1157 & n38854;
  assign n38856 = n38347 & ~n38402;
  assign n38857 = n38346 & n38361;
  assign n38858 = pi208 & ~n38857;
  assign n38859 = ~n38688 & n38858;
  assign n38860 = ~n38856 & ~n38859;
  assign n38861 = pi1157 & ~n38860;
  assign n38862 = ~pi211 & ~n38861;
  assign n38863 = ~n38855 & n38862;
  assign n38864 = ~n38415 & ~n38854;
  assign n38865 = pi211 & n38864;
  assign n38866 = ~n38863 & ~n38865;
  assign n38867 = n38468 & ~n38866;
  assign n38868 = ~pi211 & ~n38864;
  assign n38869 = n38312 & n38318;
  assign n38870 = ~pi207 & ~n38312;
  assign n38871 = ~n38321 & ~n38687;
  assign n38872 = pi207 & ~n38871;
  assign n38873 = pi208 & ~n38872;
  assign n38874 = ~n38870 & n38873;
  assign n38875 = ~n38869 & ~n38874;
  assign n38876 = pi211 & ~n38875;
  assign n38877 = n10669 & ~n38876;
  assign n38878 = ~n38868 & n38877;
  assign n38879 = n38135 & ~n38854;
  assign n38880 = ~n38878 & ~n38879;
  assign n38881 = ~n38867 & n38880;
  assign n38882 = ~pi219 & ~n38881;
  assign n38883 = ~pi211 & n38875;
  assign n38884 = pi211 & ~n38854;
  assign n38885 = ~n38145 & ~n38884;
  assign n38886 = ~n38883 & n38885;
  assign n38887 = n38145 & n38854;
  assign n38888 = pi219 & ~n38887;
  assign n38889 = ~n38886 & n38888;
  assign n38890 = ~pi209 & ~n38889;
  assign n38891 = ~n38882 & n38890;
  assign n38892 = ~n38846 & ~n38891;
  assign n38893 = ~po1038 & ~n38892;
  assign n38894 = ~pi214 & ~n38212;
  assign n38895 = ~n38769 & ~n38894;
  assign n38896 = pi212 & ~n38895;
  assign n38897 = ~pi219 & ~n38896;
  assign n38898 = ~n38214 & n38897;
  assign n38899 = pi219 & ~n38204;
  assign n38900 = pi219 & ~n38468;
  assign n38901 = ~n38899 & ~n38900;
  assign n38902 = po1038 & n38901;
  assign n38903 = ~n38898 & n38902;
  assign n38904 = pi213 & ~n38903;
  assign n38905 = ~n38893 & n38904;
  assign n38906 = pi1157 & ~n38829;
  assign n38907 = pi299 & ~pi1157;
  assign n38908 = ~n38788 & ~n38907;
  assign n38909 = ~n38906 & n38908;
  assign n38910 = ~n38357 & ~n38909;
  assign n38911 = ~pi211 & ~n38910;
  assign n38912 = n38840 & ~n38911;
  assign n38913 = n38843 & ~n38912;
  assign n38914 = pi211 & n38910;
  assign n38915 = ~n38281 & ~n38371;
  assign n38916 = ~n38287 & ~n38915;
  assign n38917 = pi207 & ~n38916;
  assign n38918 = pi1154 & ~n38352;
  assign n38919 = ~n38257 & ~n38918;
  assign n38920 = ~pi207 & ~n38319;
  assign n38921 = ~n38919 & n38920;
  assign n38922 = ~n38917 & ~n38921;
  assign n38923 = pi208 & ~n38922;
  assign n38924 = ~n38391 & ~n38923;
  assign n38925 = ~pi1157 & ~n38924;
  assign n38926 = n38389 & ~n38829;
  assign n38927 = ~n38925 & ~n38926;
  assign n38928 = ~pi211 & ~n38927;
  assign n38929 = n10669 & ~n38928;
  assign n38930 = ~n38914 & n38929;
  assign n38931 = pi211 & n38927;
  assign n38932 = ~n38838 & ~n38931;
  assign n38933 = n38468 & ~n38932;
  assign n38934 = ~n38823 & ~n38933;
  assign n38935 = ~n38930 & n38934;
  assign n38936 = ~pi219 & ~n38935;
  assign n38937 = ~n38913 & ~n38936;
  assign n38938 = pi209 & ~n38937;
  assign n38939 = n38347 & ~n38361;
  assign n38940 = ~pi207 & ~n38361;
  assign n38941 = n38675 & ~n38940;
  assign n38942 = n38858 & ~n38941;
  assign n38943 = ~n38939 & ~n38942;
  assign n38944 = ~pi211 & n38943;
  assign n38945 = n38885 & ~n38944;
  assign n38946 = n38888 & ~n38945;
  assign n38947 = pi207 & ~n38686;
  assign n38948 = ~pi207 & ~n38384;
  assign n38949 = ~n38947 & ~n38948;
  assign n38950 = pi208 & ~n38949;
  assign n38951 = n38347 & ~n38384;
  assign n38952 = ~n38950 & ~n38951;
  assign n38953 = pi211 & n38952;
  assign n38954 = ~n38883 & ~n38953;
  assign n38955 = ~n38145 & ~n38954;
  assign n38956 = ~pi211 & ~n38952;
  assign n38957 = pi211 & ~n38943;
  assign n38958 = n10669 & ~n38957;
  assign n38959 = ~n38956 & n38958;
  assign n38960 = ~n38879 & ~n38959;
  assign n38961 = ~n38955 & n38960;
  assign n38962 = ~pi219 & ~n38961;
  assign n38963 = ~n38946 & ~n38962;
  assign n38964 = ~pi209 & ~n38963;
  assign n38965 = ~po1038 & ~n38964;
  assign n38966 = ~n38938 & n38965;
  assign n38967 = n10669 & ~n38505;
  assign n38968 = ~n38206 & n38468;
  assign n38969 = ~pi219 & ~n38968;
  assign n38970 = ~n38967 & n38969;
  assign n38971 = pi219 & ~n38222;
  assign n38972 = po1038 & ~n38971;
  assign n38973 = ~n38900 & n38972;
  assign n38974 = ~n38970 & n38973;
  assign n38975 = ~pi213 & ~n38974;
  assign n38976 = ~n38966 & n38975;
  assign n38977 = ~n38905 & ~n38976;
  assign n38978 = pi230 & ~n38977;
  assign n38979 = ~pi230 & ~pi235;
  assign po392 = ~n38978 & ~n38979;
  assign n38981 = ~pi100 & n37908;
  assign n38982 = n38119 & ~n38981;
  assign n38983 = ~n6269 & ~n38982;
  assign n38984 = ~pi75 & ~n38983;
  assign n38985 = ~n7269 & ~n38984;
  assign n38986 = ~pi92 & ~n38985;
  assign n38987 = n13563 & ~n38986;
  assign n38988 = ~pi74 & ~n38987;
  assign n38989 = n6108 & ~n38988;
  assign n38990 = ~pi56 & ~n38989;
  assign n38991 = ~n6104 & ~n38990;
  assign n38992 = ~pi62 & ~n38991;
  assign po393 = n13571 & ~n38992;
  assign n38994 = ~pi211 & pi1145;
  assign n38995 = pi211 & pi1144;
  assign n38996 = ~n38994 & ~n38995;
  assign n38997 = ~n10669 & n38996;
  assign n38998 = n10669 & n38142;
  assign n38999 = ~n38135 & ~n38998;
  assign n39000 = ~n38997 & n38999;
  assign n39001 = ~pi219 & ~n39000;
  assign n39002 = pi219 & ~n38147;
  assign n39003 = n38138 & ~n39002;
  assign n39004 = ~n39001 & n39003;
  assign n39005 = n38230 & n39000;
  assign n39006 = pi199 & pi1143;
  assign n39007 = ~pi200 & ~n39006;
  assign n39008 = ~n38156 & n39007;
  assign n39009 = pi208 & n38164;
  assign n39010 = ~n38159 & n39009;
  assign n39011 = ~n39008 & n39010;
  assign n39012 = ~pi199 & pi1145;
  assign n39013 = n39007 & ~n39012;
  assign n39014 = pi200 & ~n38156;
  assign n39015 = n38512 & ~n39014;
  assign n39016 = ~n39013 & n39015;
  assign n39017 = ~n39011 & ~n39016;
  assign n39018 = ~pi299 & ~n39017;
  assign n39019 = pi299 & n38635;
  assign n39020 = n38147 & n39019;
  assign n39021 = ~n39018 & ~n39020;
  assign n39022 = ~n39005 & n39021;
  assign n39023 = ~po1038 & ~n39022;
  assign n39024 = ~n39004 & ~n39023;
  assign n39025 = pi213 & n39024;
  assign n39026 = pi211 & pi1157;
  assign n39027 = ~pi211 & pi1158;
  assign n39028 = ~n39026 & ~n39027;
  assign n39029 = n38143 & ~n39028;
  assign n39030 = n38897 & ~n39029;
  assign n39031 = ~pi219 & po1038;
  assign n39032 = n38143 & n38200;
  assign n39033 = po1038 & n39032;
  assign n39034 = ~n39031 & ~n39033;
  assign n39035 = pi214 & n38220;
  assign n39036 = pi1155 & n38379;
  assign n39037 = ~n39035 & ~n39036;
  assign n39038 = pi212 & ~n39037;
  assign n39039 = po1038 & n39038;
  assign n39040 = n39034 & ~n39039;
  assign n39041 = ~n39030 & ~n39040;
  assign n39042 = ~pi213 & ~n39041;
  assign n39043 = n38230 & ~n39030;
  assign n39044 = n38143 & n38415;
  assign n39045 = ~pi214 & ~n38232;
  assign n39046 = pi214 & ~n38234;
  assign n39047 = pi212 & ~n39046;
  assign n39048 = ~n39045 & n39047;
  assign n39049 = ~n39044 & ~n39048;
  assign n39050 = n38241 & ~n39049;
  assign n39051 = ~n39018 & ~n39050;
  assign n39052 = ~n39043 & n39051;
  assign n39053 = ~po1038 & ~n39052;
  assign n39054 = n39042 & ~n39053;
  assign n39055 = pi209 & ~n39054;
  assign n39056 = ~n39025 & n39055;
  assign n39057 = pi207 & n38288;
  assign n39058 = pi208 & ~n38814;
  assign n39059 = ~n39057 & n39058;
  assign n39060 = pi1158 & n38620;
  assign n39061 = ~pi199 & ~pi1158;
  assign n39062 = pi1156 & ~n39061;
  assign n39063 = ~n39060 & ~n39062;
  assign n39064 = n38701 & ~n39063;
  assign n39065 = ~n10564 & n38270;
  assign n39066 = ~n38511 & n39065;
  assign n39067 = n39064 & n39066;
  assign n39068 = ~n39059 & ~n39067;
  assign n39069 = ~pi1157 & ~n39068;
  assign n39070 = pi1156 & n38328;
  assign n39071 = ~pi200 & ~pi1158;
  assign n39072 = ~pi199 & ~n39071;
  assign n39073 = ~n39070 & ~n39072;
  assign n39074 = n38164 & ~n39073;
  assign n39075 = ~pi208 & n39074;
  assign n39076 = pi208 & ~n38818;
  assign n39077 = ~n39057 & n39076;
  assign n39078 = ~n39075 & ~n39077;
  assign n39079 = pi1157 & ~n39078;
  assign n39080 = ~n39069 & ~n39079;
  assign n39081 = ~pi214 & n39080;
  assign n39082 = ~pi212 & ~n39081;
  assign n39083 = ~pi299 & n39073;
  assign n39084 = n38347 & ~n39083;
  assign n39085 = ~n38536 & n38826;
  assign n39086 = ~n39084 & ~n39085;
  assign n39087 = pi1157 & ~n39086;
  assign n39088 = ~n39069 & ~n39087;
  assign n39089 = pi211 & n39088;
  assign n39090 = pi1158 & n38372;
  assign n39091 = ~pi1158 & n38288;
  assign n39092 = pi207 & ~n39091;
  assign n39093 = ~n39090 & n39092;
  assign n39094 = ~pi207 & ~n38344;
  assign n39095 = pi299 & ~pi1158;
  assign n39096 = n39094 & ~n39095;
  assign n39097 = ~n39093 & ~n39096;
  assign n39098 = n38789 & ~n39097;
  assign n39099 = ~pi207 & ~n39095;
  assign n39100 = ~n38354 & n39099;
  assign n39101 = pi208 & ~n39100;
  assign n39102 = ~n39093 & n39101;
  assign n39103 = ~pi299 & ~n38677;
  assign n39104 = pi1158 & ~n39103;
  assign n39105 = n38164 & n39070;
  assign n39106 = ~pi208 & ~n39105;
  assign n39107 = ~n39104 & n39106;
  assign n39108 = ~pi1157 & ~n39107;
  assign n39109 = ~n39102 & n39108;
  assign n39110 = n38256 & ~n38331;
  assign n39111 = pi1157 & ~n39060;
  assign n39112 = ~n39110 & n39111;
  assign n39113 = pi207 & ~n39112;
  assign n39114 = ~n39104 & ~n39113;
  assign n39115 = n38414 & ~n39114;
  assign n39116 = ~pi211 & ~n39115;
  assign n39117 = ~n39109 & n39116;
  assign n39118 = ~n39098 & n39117;
  assign n39119 = ~n39089 & ~n39118;
  assign n39120 = pi214 & ~n39119;
  assign n39121 = n39082 & ~n39120;
  assign n39122 = n38379 & ~n39088;
  assign n39123 = pi207 & ~n38409;
  assign n39124 = pi208 & ~n38784;
  assign n39125 = ~n39123 & n39124;
  assign n39126 = n38752 & ~n39064;
  assign n39127 = ~pi1157 & ~n39126;
  assign n39128 = ~n39125 & n39127;
  assign n39129 = ~n38791 & ~n39123;
  assign n39130 = n38789 & ~n39129;
  assign n39131 = ~n38415 & ~n39074;
  assign n39132 = n38414 & ~n39131;
  assign n39133 = ~n39130 & ~n39132;
  assign n39134 = ~n39128 & n39133;
  assign n39135 = n38425 & ~n39134;
  assign n39136 = ~n38232 & n38288;
  assign n39137 = pi207 & ~n39136;
  assign n39138 = ~n38799 & ~n39137;
  assign n39139 = pi208 & ~n39138;
  assign n39140 = ~pi208 & n38232;
  assign n39141 = ~n39067 & ~n39140;
  assign n39142 = ~n39139 & n39141;
  assign n39143 = ~pi1157 & ~n39142;
  assign n39144 = ~n38804 & ~n39137;
  assign n39145 = n38789 & ~n39144;
  assign n39146 = ~n39064 & ~n39072;
  assign n39147 = n38164 & ~n39146;
  assign n39148 = ~n38232 & ~n39147;
  assign n39149 = n38414 & ~n39148;
  assign n39150 = ~n39145 & ~n39149;
  assign n39151 = ~n39143 & n39150;
  assign n39152 = n10426 & ~n39151;
  assign n39153 = ~n39135 & ~n39152;
  assign n39154 = ~n39122 & n39153;
  assign n39155 = pi212 & ~n39154;
  assign n39156 = ~pi219 & ~n39155;
  assign n39157 = ~n39121 & n39156;
  assign n39158 = ~n38136 & n39080;
  assign n39159 = n38143 & n39134;
  assign n39160 = ~pi214 & ~n39151;
  assign n39161 = ~n38388 & n39094;
  assign n39162 = pi1157 & ~n39161;
  assign n39163 = ~pi1157 & ~n39067;
  assign n39164 = ~n38921 & n39163;
  assign n39165 = ~n39162 & ~n39164;
  assign n39166 = pi208 & ~n38523;
  assign n39167 = ~n39165 & n39166;
  assign n39168 = ~pi299 & ~n38701;
  assign n39169 = ~pi208 & ~n39168;
  assign n39170 = ~n38414 & ~n39169;
  assign n39171 = n39147 & ~n39170;
  assign n39172 = ~pi208 & ~n39171;
  assign n39173 = ~n38234 & n39172;
  assign n39174 = pi214 & ~n39173;
  assign n39175 = ~n39167 & n39174;
  assign n39176 = pi212 & ~n39175;
  assign n39177 = ~n39160 & n39176;
  assign n39178 = ~n39159 & ~n39177;
  assign n39179 = ~pi211 & ~n39178;
  assign n39180 = ~n39158 & ~n39179;
  assign n39181 = pi219 & ~n39180;
  assign n39182 = ~po1038 & ~n39181;
  assign n39183 = ~n39157 & n39182;
  assign n39184 = n39042 & ~n39183;
  assign n39185 = pi299 & pi1145;
  assign n39186 = ~n38438 & ~n39185;
  assign n39187 = pi207 & ~n39186;
  assign n39188 = ~pi200 & pi1157;
  assign n39189 = ~pi199 & n39188;
  assign n39190 = n38354 & ~n39189;
  assign n39191 = pi299 & ~pi1145;
  assign n39192 = ~pi207 & ~n39191;
  assign n39193 = ~n39190 & n39192;
  assign n39194 = pi208 & ~n39193;
  assign n39195 = ~n39187 & n39194;
  assign n39196 = n39172 & ~n39185;
  assign n39197 = ~n39195 & ~n39196;
  assign n39198 = ~pi211 & ~n39197;
  assign n39199 = ~n38454 & n39172;
  assign n39200 = pi207 & ~n38455;
  assign n39201 = ~pi207 & ~n38460;
  assign n39202 = ~n39190 & n39201;
  assign n39203 = pi208 & ~n39202;
  assign n39204 = ~n39200 & n39203;
  assign n39205 = ~n39199 & ~n39204;
  assign n39206 = pi211 & ~n39205;
  assign n39207 = ~n39198 & ~n39206;
  assign n39208 = ~pi214 & ~n39207;
  assign n39209 = ~n38437 & n39172;
  assign n39210 = pi207 & ~n38439;
  assign n39211 = ~pi207 & ~n38444;
  assign n39212 = ~n39190 & n39211;
  assign n39213 = pi208 & ~n39212;
  assign n39214 = ~n39210 & n39213;
  assign n39215 = ~n39209 & ~n39214;
  assign n39216 = pi211 & n39215;
  assign n39217 = ~pi211 & n39205;
  assign n39218 = pi214 & ~n39217;
  assign n39219 = ~n39216 & n39218;
  assign n39220 = pi212 & ~n39219;
  assign n39221 = ~n39208 & n39220;
  assign n39222 = pi214 & ~n39207;
  assign n39223 = n39082 & ~n39222;
  assign n39224 = ~pi219 & ~n39223;
  assign n39225 = ~n39221 & n39224;
  assign n39226 = n38136 & ~n39215;
  assign n39227 = ~n39158 & ~n39226;
  assign n39228 = pi219 & ~n39227;
  assign n39229 = ~po1038 & ~n39228;
  assign n39230 = ~n39225 & n39229;
  assign n39231 = pi213 & ~n39004;
  assign n39232 = ~n39230 & n39231;
  assign n39233 = ~pi209 & ~n39232;
  assign n39234 = ~n39184 & n39233;
  assign n39235 = ~n39056 & ~n39234;
  assign n39236 = pi230 & ~n39235;
  assign n39237 = ~pi230 & ~pi237;
  assign po394 = n39236 | n39237;
  assign n39239 = ~pi211 & ~pi1153;
  assign n39240 = pi219 & n39239;
  assign n39241 = n38138 & ~n39240;
  assign n39242 = ~n38970 & n39241;
  assign n39243 = n38255 & n39009;
  assign n39244 = ~n39066 & ~n39243;
  assign n39245 = ~n38627 & ~n39244;
  assign n39246 = ~n38232 & ~n39245;
  assign n39247 = n38379 & n39246;
  assign n39248 = n38164 & ~n38255;
  assign n39249 = pi208 & ~n39248;
  assign n39250 = pi200 & n38346;
  assign n39251 = n39249 & ~n39250;
  assign n39252 = ~n39169 & ~n39251;
  assign n39253 = ~n38650 & ~n39252;
  assign n39254 = n10426 & ~n39253;
  assign n39255 = ~n38234 & n38425;
  assign n39256 = ~n39245 & n39255;
  assign n39257 = pi212 & ~n39256;
  assign n39258 = ~n39254 & n39257;
  assign n39259 = ~n39247 & n39258;
  assign n39260 = ~pi219 & ~n39259;
  assign n39261 = ~pi299 & ~n39253;
  assign n39262 = pi299 & n38206;
  assign n39263 = n38512 & n38620;
  assign n39264 = pi1153 & n39263;
  assign n39265 = n38261 & ~n38511;
  assign n39266 = ~n39263 & n39265;
  assign n39267 = ~pi214 & ~n39266;
  assign n39268 = ~n39264 & n39267;
  assign n39269 = ~pi212 & ~n39268;
  assign n39270 = ~n39262 & n39269;
  assign n39271 = ~n39261 & n39270;
  assign n39272 = n39260 & ~n39271;
  assign n39273 = pi1151 & ~po1038;
  assign n39274 = ~pi211 & ~n39252;
  assign n39275 = pi211 & ~n39244;
  assign n39276 = ~n39274 & ~n39275;
  assign n39277 = ~n38650 & ~n39276;
  assign n39278 = n38135 & ~n39245;
  assign n39279 = n39277 & ~n39278;
  assign n39280 = pi219 & ~n39279;
  assign n39281 = n39273 & ~n39280;
  assign n39282 = ~n39272 & n39281;
  assign n39283 = ~n38234 & ~n39264;
  assign n39284 = ~pi211 & ~n39283;
  assign n39285 = n10758 & n38512;
  assign n39286 = ~pi299 & ~n39285;
  assign n39287 = n38504 & ~n39286;
  assign n39288 = n10669 & ~n39287;
  assign n39289 = ~n39284 & n39288;
  assign n39290 = pi299 & ~n38206;
  assign n39291 = ~n38145 & ~n39290;
  assign n39292 = ~n39264 & n39291;
  assign n39293 = ~n39289 & ~n39292;
  assign n39294 = ~pi219 & ~n39293;
  assign n39295 = ~pi1151 & ~po1038;
  assign n39296 = ~n12978 & ~n39286;
  assign n39297 = ~pi214 & ~n39263;
  assign n39298 = ~pi212 & n39297;
  assign n39299 = n39296 & ~n39298;
  assign n39300 = pi1153 & n39299;
  assign n39301 = ~n38474 & ~n39300;
  assign n39302 = n39295 & ~n39301;
  assign n39303 = ~n39294 & n39302;
  assign n39304 = ~pi1152 & ~n39303;
  assign n39305 = ~n39282 & n39304;
  assign n39306 = pi1153 & ~n39286;
  assign n39307 = ~n38512 & ~n38677;
  assign n39308 = ~n10564 & n38350;
  assign n39309 = ~n39307 & ~n39308;
  assign n39310 = n39286 & n39309;
  assign n39311 = ~n39306 & ~n39310;
  assign n39312 = pi211 & ~n39311;
  assign n39313 = n38347 & ~n38613;
  assign n39314 = pi200 & pi207;
  assign n39315 = ~pi199 & ~n39314;
  assign n39316 = ~pi299 & ~n39315;
  assign n39317 = pi208 & ~n39316;
  assign n39318 = ~pi207 & n38613;
  assign n39319 = n39317 & ~n39318;
  assign n39320 = ~n39313 & ~n39319;
  assign n39321 = ~pi211 & ~n38388;
  assign n39322 = ~n39320 & n39321;
  assign n39323 = ~n39312 & ~n39322;
  assign n39324 = n10669 & ~n39323;
  assign n39325 = ~n38145 & ~n39320;
  assign n39326 = ~n39262 & n39325;
  assign n39327 = ~n39324 & ~n39326;
  assign n39328 = ~pi219 & ~n39327;
  assign n39329 = ~pi211 & n38236;
  assign n39330 = ~n38135 & n39329;
  assign n39331 = n38703 & ~n39320;
  assign n39332 = ~n39330 & ~n39331;
  assign n39333 = ~n38474 & ~n39332;
  assign n39334 = ~n39328 & ~n39333;
  assign n39335 = n39295 & ~n39334;
  assign n39336 = ~pi299 & ~n39265;
  assign n39337 = ~n10564 & n38614;
  assign n39338 = ~n39336 & ~n39337;
  assign n39339 = ~pi211 & n39338;
  assign n39340 = ~n38369 & n39339;
  assign n39341 = pi211 & n39338;
  assign n39342 = ~n38388 & n39341;
  assign n39343 = ~n39340 & ~n39342;
  assign n39344 = ~n38145 & ~n39343;
  assign n39345 = ~n39266 & ~n39287;
  assign n39346 = ~n39322 & n39345;
  assign n39347 = n10669 & ~n39346;
  assign n39348 = ~pi214 & n39269;
  assign n39349 = ~pi219 & ~n39348;
  assign n39350 = ~n39347 & n39349;
  assign n39351 = ~n39344 & n39350;
  assign n39352 = pi219 & ~n39266;
  assign n39353 = ~n39300 & n39352;
  assign n39354 = n39273 & ~n39353;
  assign n39355 = ~n39351 & n39354;
  assign n39356 = pi1152 & ~n39355;
  assign n39357 = ~n39335 & n39356;
  assign n39358 = ~n39305 & ~n39357;
  assign n39359 = ~pi209 & ~n39358;
  assign n39360 = pi1153 & ~n38320;
  assign n39361 = ~n38622 & ~n39360;
  assign n39362 = n38164 & n39361;
  assign n39363 = pi208 & ~n39362;
  assign n39364 = ~n38164 & n38384;
  assign n39365 = n39363 & ~n39364;
  assign n39366 = ~n38951 & ~n39365;
  assign n39367 = pi211 & ~n39366;
  assign n39368 = ~n38164 & ~n38312;
  assign n39369 = n39363 & ~n39368;
  assign n39370 = ~n38869 & ~n39369;
  assign n39371 = ~pi211 & ~n39370;
  assign n39372 = n38143 & ~n39371;
  assign n39373 = ~n39367 & n39372;
  assign n39374 = n38425 & ~n39366;
  assign n39375 = n38379 & ~n39370;
  assign n39376 = ~n38857 & n39363;
  assign n39377 = ~n38856 & ~n39376;
  assign n39378 = ~n38265 & ~n38857;
  assign n39379 = ~n39377 & n39378;
  assign n39380 = n10426 & n39379;
  assign n39381 = pi212 & ~n39380;
  assign n39382 = ~n39375 & n39381;
  assign n39383 = ~n39374 & n39382;
  assign n39384 = ~n39373 & ~n39383;
  assign n39385 = ~pi219 & ~n39384;
  assign n39386 = ~pi299 & ~n39362;
  assign n39387 = n10564 & ~n39386;
  assign n39388 = ~n38853 & ~n39387;
  assign n39389 = pi211 & n39388;
  assign n39390 = ~pi211 & n39379;
  assign n39391 = ~n39389 & ~n39390;
  assign n39392 = n38635 & n39391;
  assign n39393 = ~pi214 & ~n39388;
  assign n39394 = ~pi212 & n39393;
  assign n39395 = ~po1038 & ~n39394;
  assign n39396 = ~n39392 & n39395;
  assign n39397 = ~n39385 & n39396;
  assign n39398 = pi209 & ~n39397;
  assign n39399 = ~n39359 & ~n39398;
  assign n39400 = ~n39242 & ~n39399;
  assign n39401 = pi213 & ~n39400;
  assign n39402 = ~n10427 & n38474;
  assign n39403 = po1038 & n39402;
  assign n39404 = ~n10669 & ~n39239;
  assign n39405 = ~n38436 & ~n39404;
  assign n39406 = n39403 & ~n39405;
  assign n39407 = ~n10428 & n38138;
  assign n39408 = pi1151 & ~n39407;
  assign n39409 = ~n39406 & n39408;
  assign n39410 = ~pi211 & ~n39377;
  assign n39411 = ~n39389 & ~n39410;
  assign n39412 = ~n38135 & n39411;
  assign n39413 = ~n39394 & ~n39412;
  assign n39414 = pi219 & ~n39413;
  assign n39415 = ~po1038 & ~n39414;
  assign n39416 = pi211 & ~n39377;
  assign n39417 = ~n39390 & ~n39416;
  assign n39418 = pi214 & n39417;
  assign n39419 = ~pi212 & ~n39393;
  assign n39420 = ~n39418 & n39419;
  assign n39421 = ~pi219 & ~n39420;
  assign n39422 = ~pi214 & ~n39417;
  assign n39423 = pi214 & ~n39377;
  assign n39424 = ~n39422 & ~n39423;
  assign n39425 = pi212 & ~n39424;
  assign n39426 = n39421 & ~n39425;
  assign n39427 = n39415 & ~n39426;
  assign n39428 = n39409 & ~n39427;
  assign n39429 = ~pi1151 & ~n39406;
  assign n39430 = pi214 & ~n39411;
  assign n39431 = ~n39422 & ~n39430;
  assign n39432 = pi212 & ~n39431;
  assign n39433 = n39421 & ~n39432;
  assign n39434 = pi219 & ~n39388;
  assign n39435 = ~po1038 & ~n39434;
  assign n39436 = ~n39433 & n39435;
  assign n39437 = n39429 & ~n39436;
  assign n39438 = pi1152 & ~n39437;
  assign n39439 = ~n39428 & n39438;
  assign n39440 = pi214 & n39391;
  assign n39441 = ~n39393 & ~n39440;
  assign n39442 = ~pi212 & ~n39441;
  assign n39443 = ~pi211 & n39388;
  assign n39444 = ~n39416 & ~n39443;
  assign n39445 = pi214 & ~n39444;
  assign n39446 = ~pi214 & ~n39391;
  assign n39447 = pi212 & ~n39446;
  assign n39448 = ~n39445 & n39447;
  assign n39449 = ~n39442 & ~n39448;
  assign n39450 = ~pi219 & ~n39449;
  assign n39451 = n39415 & ~n39450;
  assign n39452 = n10672 & n38474;
  assign n39453 = po1038 & n39452;
  assign n39454 = ~n39407 & ~n39453;
  assign n39455 = pi1151 & n39454;
  assign n39456 = po1038 & ~n39452;
  assign n39457 = pi1151 & ~n39456;
  assign n39458 = ~pi1153 & n39457;
  assign n39459 = ~n39455 & ~n39458;
  assign n39460 = ~n39451 & ~n39459;
  assign n39461 = pi1153 & n39453;
  assign n39462 = ~pi1151 & ~n39461;
  assign n39463 = ~pi219 & n38468;
  assign n39464 = n39391 & n39463;
  assign n39465 = ~n39388 & ~n39463;
  assign n39466 = ~po1038 & ~n39465;
  assign n39467 = ~n39464 & n39466;
  assign n39468 = n39462 & ~n39467;
  assign n39469 = ~pi1152 & ~n39468;
  assign n39470 = ~n39460 & n39469;
  assign n39471 = pi209 & ~n39470;
  assign n39472 = ~n39439 & n39471;
  assign n39473 = ~pi214 & n39277;
  assign n39474 = ~n12978 & ~n39264;
  assign n39475 = ~n39245 & n39474;
  assign n39476 = pi214 & ~n39475;
  assign n39477 = pi212 & ~n39476;
  assign n39478 = ~n39473 & n39477;
  assign n39479 = ~pi212 & ~n39279;
  assign n39480 = ~n39478 & ~n39479;
  assign n39481 = ~pi219 & ~n39480;
  assign n39482 = ~pi211 & pi299;
  assign n39483 = ~n39245 & ~n39482;
  assign n39484 = ~n39278 & ~n39483;
  assign n39485 = pi219 & ~n39484;
  assign n39486 = ~po1038 & ~n39485;
  assign n39487 = ~n39481 & n39486;
  assign n39488 = ~n39459 & ~n39487;
  assign n39489 = n39297 & n39300;
  assign n39490 = ~pi214 & n12978;
  assign n39491 = pi212 & ~n39490;
  assign n39492 = ~n39474 & n39491;
  assign n39493 = ~pi219 & ~n39492;
  assign n39494 = n38143 & n39329;
  assign n39495 = ~n39263 & ~n39494;
  assign n39496 = n39493 & n39495;
  assign n39497 = ~n39489 & n39496;
  assign n39498 = pi219 & ~n39263;
  assign n39499 = ~po1038 & ~n39498;
  assign n39500 = n39300 & n39499;
  assign n39501 = ~n39497 & n39500;
  assign n39502 = n39462 & ~n39501;
  assign n39503 = ~pi1152 & ~n39502;
  assign n39504 = ~n39488 & n39503;
  assign n39505 = ~n39264 & ~n39266;
  assign n39506 = ~n39339 & n39505;
  assign n39507 = pi214 & n39506;
  assign n39508 = ~n39268 & ~n39507;
  assign n39509 = ~pi212 & ~n39508;
  assign n39510 = ~n39506 & ~n39509;
  assign n39511 = pi219 & ~n39510;
  assign n39512 = ~po1038 & ~n39511;
  assign n39513 = ~n39306 & ~n39341;
  assign n39514 = n39267 & n39513;
  assign n39515 = pi214 & ~n39338;
  assign n39516 = pi212 & ~n39515;
  assign n39517 = ~n39514 & n39516;
  assign n39518 = pi214 & ~n39266;
  assign n39519 = n39513 & n39518;
  assign n39520 = n39269 & ~n39519;
  assign n39521 = ~pi219 & ~n39520;
  assign n39522 = ~n39517 & n39521;
  assign n39523 = n39512 & ~n39522;
  assign n39524 = n39409 & ~n39523;
  assign n39525 = pi219 & ~n39331;
  assign n39526 = ~po1038 & ~n39525;
  assign n39527 = ~pi211 & n39311;
  assign n39528 = n39325 & ~n39527;
  assign n39529 = ~n38468 & n39331;
  assign n39530 = pi299 & n38436;
  assign n39531 = ~pi219 & ~n39530;
  assign n39532 = ~n39529 & n39531;
  assign n39533 = ~n39528 & n39532;
  assign n39534 = n39526 & ~n39533;
  assign n39535 = n39429 & ~n39534;
  assign n39536 = pi1152 & ~n39535;
  assign n39537 = ~n39524 & n39536;
  assign n39538 = ~n39504 & ~n39537;
  assign n39539 = ~pi209 & n39538;
  assign n39540 = ~pi213 & ~n39539;
  assign n39541 = ~n39472 & n39540;
  assign n39542 = ~n39401 & ~n39541;
  assign n39543 = pi230 & ~n39542;
  assign n39544 = ~pi230 & pi238;
  assign po395 = n39543 | n39544;
  assign n39546 = n38171 & ~n38288;
  assign n39547 = ~pi214 & n39546;
  assign n39548 = ~pi212 & ~n39547;
  assign n39549 = ~pi219 & n39548;
  assign n39550 = pi299 & pi1158;
  assign n39551 = ~n38171 & n39550;
  assign n39552 = ~pi208 & n39093;
  assign n39553 = ~n39551 & ~n39552;
  assign n39554 = ~pi211 & ~n39553;
  assign n39555 = pi208 & pi299;
  assign n39556 = pi1157 & ~n39555;
  assign n39557 = ~n38537 & n39556;
  assign n39558 = ~pi1157 & ~n39546;
  assign n39559 = pi211 & ~n39558;
  assign n39560 = ~n39557 & n39559;
  assign n39561 = ~n39554 & ~n39560;
  assign n39562 = pi214 & ~n39561;
  assign n39563 = n39549 & ~n39562;
  assign n39564 = pi219 & n39548;
  assign n39565 = pi211 & ~n39546;
  assign n39566 = pi214 & ~n39565;
  assign n39567 = ~n38580 & n38721;
  assign n39568 = n39566 & ~n39567;
  assign n39569 = n39564 & ~n39568;
  assign n39570 = pi212 & ~n39546;
  assign n39571 = ~po1038 & ~n39570;
  assign n39572 = ~pi209 & n39571;
  assign n39573 = ~n39569 & n39572;
  assign n39574 = ~n39563 & n39573;
  assign n39575 = ~pi214 & n39171;
  assign n39576 = ~pi212 & ~n39575;
  assign n39577 = ~pi219 & n39576;
  assign n39578 = ~n39084 & n39556;
  assign n39579 = ~n39163 & ~n39578;
  assign n39580 = pi211 & ~n39579;
  assign n39581 = pi214 & ~n39580;
  assign n39582 = ~pi211 & ~n39550;
  assign n39583 = ~n39171 & n39582;
  assign n39584 = n39581 & ~n39583;
  assign n39585 = n39577 & ~n39584;
  assign n39586 = pi219 & n39576;
  assign n39587 = pi211 & ~n39171;
  assign n39588 = n38721 & ~n39171;
  assign n39589 = pi214 & ~n39588;
  assign n39590 = ~n39587 & n39589;
  assign n39591 = n39586 & ~n39590;
  assign n39592 = pi212 & ~n39171;
  assign n39593 = ~po1038 & ~n39592;
  assign n39594 = pi209 & n39593;
  assign n39595 = ~n39591 & n39594;
  assign n39596 = ~n39585 & n39595;
  assign n39597 = ~pi219 & ~n39029;
  assign n39598 = ~n39034 & ~n39597;
  assign n39599 = pi213 & ~n39598;
  assign n39600 = ~n39596 & n39599;
  assign n39601 = ~n39574 & n39600;
  assign n39602 = ~pi211 & ~n38234;
  assign n39603 = ~n39171 & n39602;
  assign n39604 = pi214 & ~n39587;
  assign n39605 = ~n39603 & n39604;
  assign n39606 = n39586 & ~n39605;
  assign n39607 = pi211 & ~n38232;
  assign n39608 = ~n39171 & n39607;
  assign n39609 = n39589 & ~n39608;
  assign n39610 = n39577 & ~n39609;
  assign n39611 = n39593 & ~n39610;
  assign n39612 = ~n39606 & n39611;
  assign n39613 = pi209 & ~n39612;
  assign n39614 = ~n38234 & ~n38525;
  assign n39615 = n39566 & ~n39614;
  assign n39616 = n39564 & ~n39615;
  assign n39617 = ~n39546 & n39607;
  assign n39618 = pi214 & ~n39617;
  assign n39619 = ~n39567 & n39618;
  assign n39620 = n39549 & ~n39619;
  assign n39621 = n39571 & ~n39620;
  assign n39622 = ~n39616 & n39621;
  assign n39623 = ~pi209 & ~n39622;
  assign n39624 = ~n39613 & ~n39623;
  assign n39625 = po1038 & ~n38773;
  assign n39626 = n38143 & ~n38771;
  assign n39627 = n39625 & n39626;
  assign n39628 = ~pi213 & ~n39627;
  assign n39629 = ~n39624 & n39628;
  assign n39630 = ~n39601 & ~n39629;
  assign n39631 = pi230 & ~n39630;
  assign n39632 = ~pi230 & ~pi239;
  assign po396 = ~n39631 & ~n39632;
  assign n39634 = ~po1038 & n38703;
  assign n39635 = ~n39499 & ~n39634;
  assign n39636 = ~pi214 & ~n38703;
  assign n39637 = ~pi212 & ~n39636;
  assign n39638 = ~pi299 & ~n38703;
  assign n39639 = n39637 & ~n39638;
  assign n39640 = ~pi219 & ~n39639;
  assign n39641 = ~pi211 & ~n39638;
  assign n39642 = pi211 & n38703;
  assign n39643 = pi214 & ~n39642;
  assign n39644 = ~n39641 & n39643;
  assign n39645 = pi212 & ~n39644;
  assign n39646 = ~n39638 & n39645;
  assign n39647 = n39640 & ~n39646;
  assign n39648 = ~n39635 & ~n39647;
  assign n39649 = ~n39403 & ~n39648;
  assign n39650 = ~pi1147 & n39649;
  assign n39651 = pi299 & ~n38135;
  assign n39652 = ~po1038 & ~n38137;
  assign n39653 = n39651 & n39652;
  assign n39654 = ~po1038 & n39265;
  assign n39655 = ~n39653 & ~n39654;
  assign n39656 = ~n38135 & n38138;
  assign n39657 = n39655 & ~n39656;
  assign n39658 = pi1147 & n39657;
  assign n39659 = pi1149 & ~n39658;
  assign n39660 = ~n39650 & n39659;
  assign n39661 = pi211 & n38143;
  assign n39662 = pi212 & n38425;
  assign n39663 = ~n39661 & ~n39662;
  assign n39664 = n39031 & ~n39663;
  assign n39665 = pi299 & n10426;
  assign n39666 = ~n39310 & ~n39665;
  assign n39667 = ~pi212 & ~n39666;
  assign n39668 = ~pi219 & ~n39667;
  assign n39669 = ~pi299 & ~n39309;
  assign n39670 = pi214 & ~n39669;
  assign n39671 = ~pi214 & n39310;
  assign n39672 = ~pi212 & ~n39671;
  assign n39673 = ~n39670 & n39672;
  assign n39674 = ~pi211 & ~n39669;
  assign n39675 = ~n39310 & ~n39674;
  assign n39676 = pi214 & ~n39675;
  assign n39677 = pi212 & ~n39676;
  assign n39678 = ~pi214 & ~n39669;
  assign n39679 = n39677 & ~n39678;
  assign n39680 = ~n39673 & ~n39679;
  assign n39681 = ~n12978 & ~n39310;
  assign n39682 = ~n39670 & n39681;
  assign n39683 = pi212 & ~n39682;
  assign n39684 = n39680 & n39683;
  assign n39685 = n39668 & ~n39684;
  assign n39686 = pi219 & ~n39310;
  assign n39687 = ~po1038 & ~n39686;
  assign n39688 = ~n39685 & n39687;
  assign n39689 = ~n39664 & ~n39688;
  assign n39690 = ~pi1147 & n39689;
  assign n39691 = pi212 & ~n38379;
  assign n39692 = ~pi219 & ~n39661;
  assign n39693 = ~n39691 & n39692;
  assign n39694 = n39653 & ~n39693;
  assign n39695 = ~po1038 & n39266;
  assign n39696 = n38138 & ~n39693;
  assign n39697 = ~n39695 & ~n39696;
  assign n39698 = ~n39694 & n39697;
  assign n39699 = pi1147 & n39698;
  assign n39700 = ~pi1149 & ~n39699;
  assign n39701 = ~n39690 & n39700;
  assign n39702 = ~n39660 & ~n39701;
  assign n39703 = pi1148 & ~n39702;
  assign n39704 = ~pi211 & ~n39244;
  assign n39705 = pi211 & ~n39252;
  assign n39706 = pi214 & ~n39705;
  assign n39707 = ~n39704 & n39706;
  assign n39708 = n10669 & ~n39707;
  assign n39709 = ~pi214 & n39244;
  assign n39710 = ~pi212 & ~n39709;
  assign n39711 = pi214 & n39276;
  assign n39712 = n39710 & ~n39711;
  assign n39713 = ~pi219 & ~n39712;
  assign n39714 = pi212 & ~n39707;
  assign n39715 = ~n39276 & n39714;
  assign n39716 = n39713 & ~n39715;
  assign n39717 = ~n39708 & n39716;
  assign n39718 = pi212 & ~n39276;
  assign n39719 = pi219 & ~n39718;
  assign n39720 = ~n39712 & n39719;
  assign n39721 = ~po1038 & ~n39720;
  assign n39722 = ~n39717 & n39721;
  assign n39723 = n39454 & ~n39722;
  assign n39724 = pi1147 & n39723;
  assign n39725 = n16361 & n39285;
  assign n39726 = ~pi211 & n38468;
  assign n39727 = ~pi219 & ~n16361;
  assign n39728 = n39726 & n39727;
  assign n39729 = ~n39725 & ~n39728;
  assign n39730 = ~pi1147 & n39729;
  assign n39731 = pi1149 & ~n39730;
  assign n39732 = ~n39724 & n39731;
  assign n39733 = ~pi212 & ~n39665;
  assign n39734 = ~n39266 & n39733;
  assign n39735 = ~n39266 & ~n39482;
  assign n39736 = ~n39267 & ~n39735;
  assign n39737 = n39491 & ~n39736;
  assign n39738 = ~n39734 & ~n39737;
  assign n39739 = ~pi219 & ~n39738;
  assign n39740 = n38329 & ~n39314;
  assign n39741 = pi208 & ~n39740;
  assign n39742 = ~pi199 & ~n39741;
  assign n39743 = n39266 & ~n39742;
  assign n39744 = ~pi299 & ~n39743;
  assign n39745 = ~pi219 & n39744;
  assign n39746 = ~n39739 & ~n39745;
  assign n39747 = ~pi211 & ~n39746;
  assign n39748 = pi214 & ~n39296;
  assign n39749 = ~pi211 & n39297;
  assign n39750 = pi212 & ~n39286;
  assign n39751 = ~n39749 & n39750;
  assign n39752 = ~n39748 & n39751;
  assign n39753 = ~pi212 & ~n39286;
  assign n39754 = ~n39297 & n39753;
  assign n39755 = ~n39482 & n39754;
  assign n39756 = ~pi219 & ~n39755;
  assign n39757 = ~n39752 & n39756;
  assign n39758 = n39499 & ~n39757;
  assign n39759 = ~n39655 & ~n39758;
  assign n39760 = ~n39744 & n39759;
  assign n39761 = ~n39747 & n39760;
  assign n39762 = ~n39407 & ~n39761;
  assign n39763 = pi1147 & ~pi1149;
  assign n39764 = ~n39762 & n39763;
  assign n39765 = ~n39732 & ~n39764;
  assign n39766 = ~pi1148 & ~n39765;
  assign n39767 = ~n39703 & ~n39766;
  assign n39768 = pi213 & ~n39767;
  assign n39769 = ~po1038 & n39310;
  assign n39770 = ~pi211 & pi1146;
  assign n39771 = pi211 & pi1145;
  assign n39772 = ~n39770 & ~n39771;
  assign n39773 = pi214 & ~n39772;
  assign n39774 = pi211 & pi1146;
  assign n39775 = ~pi214 & n39774;
  assign n39776 = ~n39773 & ~n39775;
  assign n39777 = pi212 & ~n39776;
  assign n39778 = n38143 & n39774;
  assign n39779 = ~n39777 & ~n39778;
  assign n39780 = ~n38635 & n39779;
  assign n39781 = po1038 & n38994;
  assign n39782 = ~n39031 & ~n39781;
  assign n39783 = ~n39780 & ~n39782;
  assign n39784 = ~pi1147 & ~n39783;
  assign n39785 = ~pi211 & n39185;
  assign n39786 = pi219 & ~n39785;
  assign n39787 = n39652 & ~n39786;
  assign n39788 = pi219 & n39787;
  assign n39789 = pi299 & ~n39779;
  assign n39790 = n35887 & n39789;
  assign n39791 = ~n39788 & ~n39790;
  assign n39792 = n39784 & n39791;
  assign n39793 = ~n39769 & n39792;
  assign n39794 = pi1147 & ~n39453;
  assign n39795 = ~n39783 & n39794;
  assign n39796 = ~n39695 & ~n39787;
  assign n39797 = pi299 & pi1146;
  assign n39798 = pi211 & n39797;
  assign n39799 = ~n39482 & ~n39798;
  assign n39800 = ~n39266 & n39799;
  assign n39801 = n38468 & ~n39800;
  assign n39802 = n38135 & n39266;
  assign n39803 = ~pi219 & ~n39802;
  assign n39804 = pi299 & ~n39772;
  assign n39805 = ~n39266 & ~n39804;
  assign n39806 = n10669 & ~n39805;
  assign n39807 = n39803 & ~n39806;
  assign n39808 = ~n39801 & n39807;
  assign n39809 = ~n39796 & ~n39808;
  assign n39810 = n39795 & ~n39809;
  assign n39811 = pi1148 & ~n39810;
  assign n39812 = ~n39793 & n39811;
  assign n39813 = ~pi1146 & n12978;
  assign n39814 = n38468 & ~n39813;
  assign n39815 = ~n39806 & ~n39814;
  assign n39816 = ~pi219 & ~n39744;
  assign n39817 = ~n39815 & n39816;
  assign n39818 = n38994 & n39019;
  assign n39819 = ~n38474 & n39743;
  assign n39820 = ~n39818 & ~n39819;
  assign n39821 = ~n39817 & n39820;
  assign n39822 = ~po1038 & ~n39821;
  assign n39823 = n39795 & ~n39822;
  assign n39824 = ~pi1148 & ~n39792;
  assign n39825 = ~n39823 & n39824;
  assign n39826 = ~n39812 & ~n39825;
  assign n39827 = ~pi1149 & ~n39826;
  assign n39828 = pi219 & n39244;
  assign n39829 = ~po1038 & ~n39828;
  assign n39830 = ~n39787 & ~n39829;
  assign n39831 = ~n39275 & ~n39798;
  assign n39832 = ~n39274 & n39831;
  assign n39833 = ~pi214 & n39832;
  assign n39834 = pi214 & ~n39804;
  assign n39835 = n39244 & n39834;
  assign n39836 = pi212 & ~n39835;
  assign n39837 = ~n39833 & n39836;
  assign n39838 = pi214 & n39832;
  assign n39839 = n39710 & ~n39838;
  assign n39840 = ~pi219 & ~n39839;
  assign n39841 = ~n39837 & n39840;
  assign n39842 = ~n39830 & ~n39841;
  assign n39843 = n39795 & ~n39842;
  assign n39844 = ~n39725 & n39792;
  assign n39845 = ~pi1148 & ~n39844;
  assign n39846 = ~n39843 & n39845;
  assign n39847 = ~n38135 & n39641;
  assign n39848 = ~n38136 & n38703;
  assign n39849 = pi219 & ~n39848;
  assign n39850 = ~n39847 & n39849;
  assign n39851 = ~po1038 & ~n39850;
  assign n39852 = n11311 & n39851;
  assign n39853 = ~n39787 & ~n39852;
  assign n39854 = pi212 & ~n39638;
  assign n39855 = ~n38703 & n39776;
  assign n39856 = n39854 & ~n39855;
  assign n39857 = ~pi212 & n38703;
  assign n39858 = ~pi219 & ~n39857;
  assign n39859 = n39637 & n39798;
  assign n39860 = n39858 & ~n39859;
  assign n39861 = ~n39856 & n39860;
  assign n39862 = ~n39853 & ~n39861;
  assign n39863 = n39784 & ~n39862;
  assign n39864 = n39791 & n39795;
  assign n39865 = pi219 & ~n39265;
  assign n39866 = ~po1038 & ~n39865;
  assign n39867 = pi212 & ~n39336;
  assign n39868 = pi211 & ~n39265;
  assign n39869 = pi214 & n39868;
  assign n39870 = n39867 & ~n39869;
  assign n39871 = pi214 & pi299;
  assign n39872 = ~n39265 & ~n39871;
  assign n39873 = ~pi212 & ~n39872;
  assign n39874 = ~pi219 & ~n39873;
  assign n39875 = ~n39870 & n39874;
  assign n39876 = n39866 & ~n39875;
  assign n39877 = pi299 & n39691;
  assign n39878 = ~n39868 & ~n39877;
  assign n39879 = n39876 & n39878;
  assign n39880 = n39864 & ~n39879;
  assign n39881 = pi1148 & ~n39880;
  assign n39882 = ~n39863 & n39881;
  assign n39883 = ~n39846 & ~n39882;
  assign n39884 = pi1149 & ~n39883;
  assign n39885 = ~n39827 & ~n39884;
  assign n39886 = ~pi213 & ~n39885;
  assign n39887 = pi209 & ~n39886;
  assign n39888 = ~n39768 & n39887;
  assign n39889 = pi199 & pi1145;
  assign n39890 = ~pi200 & ~n39889;
  assign n39891 = ~pi199 & pi1146;
  assign n39892 = n39890 & ~n39891;
  assign n39893 = pi200 & ~n39012;
  assign n39894 = n38164 & ~n39893;
  assign n39895 = ~n39892 & n39894;
  assign n39896 = ~n38512 & ~n39895;
  assign n39897 = pi200 & ~n39891;
  assign n39898 = ~pi299 & ~n39897;
  assign n39899 = ~n39890 & n39898;
  assign n39900 = ~n10564 & ~n39899;
  assign n39901 = ~n39896 & ~n39900;
  assign n39902 = ~pi1147 & ~po1038;
  assign n39903 = n39901 & n39902;
  assign n39904 = ~pi200 & n38329;
  assign n39905 = n39900 & ~n39904;
  assign n39906 = ~n39896 & ~n39905;
  assign n39907 = ~n38136 & n39906;
  assign n39908 = pi219 & ~n39907;
  assign n39909 = pi208 & n39797;
  assign n39910 = ~n39906 & ~n39909;
  assign n39911 = ~pi299 & n39910;
  assign n39912 = ~pi211 & ~n39911;
  assign n39913 = ~n38135 & n39912;
  assign n39914 = n39908 & ~n39913;
  assign n39915 = ~po1038 & ~n39914;
  assign n39916 = pi211 & ~n39911;
  assign n39917 = ~n39901 & ~n39909;
  assign n39918 = ~pi299 & n39917;
  assign n39919 = pi214 & ~n39918;
  assign n39920 = ~n39916 & ~n39919;
  assign n39921 = pi212 & ~n39920;
  assign n39922 = n10426 & ~n39911;
  assign n39923 = ~pi219 & ~n39906;
  assign n39924 = ~n39922 & n39923;
  assign n39925 = ~n39921 & n39924;
  assign n39926 = n39915 & ~n39925;
  assign n39927 = ~pi214 & ~n39906;
  assign n39928 = ~n39912 & n39927;
  assign n39929 = pi214 & ~n39906;
  assign n39930 = ~n39916 & n39929;
  assign n39931 = pi212 & ~n39930;
  assign n39932 = ~n39928 & n39931;
  assign n39933 = ~n39906 & ~n39912;
  assign n39934 = ~pi212 & ~n39927;
  assign n39935 = ~n39933 & n39934;
  assign n39936 = ~pi219 & ~n39935;
  assign n39937 = ~n39932 & n39936;
  assign n39938 = n39926 & ~n39937;
  assign n39939 = ~n39407 & ~n39938;
  assign n39940 = pi1147 & ~n39939;
  assign n39941 = ~n39903 & ~n39940;
  assign n39942 = ~pi1149 & ~n39941;
  assign n39943 = n39915 & ~n39937;
  assign n39944 = n39454 & ~n39943;
  assign n39945 = pi1147 & ~n39944;
  assign n39946 = ~pi1147 & n39452;
  assign n39947 = ~n39903 & ~n39946;
  assign n39948 = n16361 & n39452;
  assign n39949 = n39917 & n39948;
  assign n39950 = ~n39947 & ~n39949;
  assign n39951 = ~n39945 & ~n39950;
  assign n39952 = pi1149 & ~n39951;
  assign n39953 = ~pi1148 & ~n39952;
  assign n39954 = ~n39942 & n39953;
  assign n39955 = pi214 & n39933;
  assign n39956 = ~n39918 & ~n39955;
  assign n39957 = pi212 & ~n39956;
  assign n39958 = ~pi212 & ~n39901;
  assign n39959 = ~n39919 & n39958;
  assign n39960 = ~n39957 & ~n39959;
  assign n39961 = ~pi219 & ~n39960;
  assign n39962 = pi219 & ~n39901;
  assign n39963 = ~po1038 & ~n39962;
  assign n39964 = ~n39961 & n39963;
  assign n39965 = ~n39925 & n39964;
  assign n39966 = ~pi1147 & ~n39664;
  assign n39967 = ~n39965 & n39966;
  assign n39968 = pi1147 & ~n39696;
  assign n39969 = ~n39926 & n39968;
  assign n39970 = ~pi1149 & ~n39969;
  assign n39971 = ~n39967 & n39970;
  assign n39972 = ~pi1147 & ~n39403;
  assign n39973 = ~n39964 & n39972;
  assign n39974 = ~n39651 & n39923;
  assign n39975 = n39915 & ~n39974;
  assign n39976 = pi1147 & ~n39656;
  assign n39977 = ~n39975 & n39976;
  assign n39978 = pi1149 & ~n39977;
  assign n39979 = ~n39973 & n39978;
  assign n39980 = pi1148 & ~n39979;
  assign n39981 = ~n39971 & n39980;
  assign n39982 = pi213 & ~n39981;
  assign n39983 = ~n39954 & n39982;
  assign n39984 = ~n39798 & ~n39901;
  assign n39985 = ~pi214 & ~n39901;
  assign n39986 = ~pi212 & ~n39985;
  assign n39987 = ~n39984 & n39986;
  assign n39988 = ~pi219 & ~n39987;
  assign n39989 = n39834 & ~n39901;
  assign n39990 = ~pi214 & n39984;
  assign n39991 = pi212 & ~n39990;
  assign n39992 = ~n39989 & n39991;
  assign n39993 = n39988 & ~n39992;
  assign n39994 = ~n39818 & n39962;
  assign n39995 = ~po1038 & ~n39994;
  assign n39996 = ~n39993 & n39995;
  assign n39997 = n39784 & ~n39996;
  assign n39998 = ~n39191 & n39916;
  assign n39999 = n39834 & n39910;
  assign n40000 = ~n39922 & ~n39999;
  assign n40001 = ~n39998 & ~n40000;
  assign n40002 = ~pi214 & n39799;
  assign n40003 = n39910 & n40002;
  assign n40004 = pi212 & ~n40003;
  assign n40005 = ~n40001 & n40004;
  assign n40006 = ~n39935 & n39988;
  assign n40007 = ~n40005 & n40006;
  assign n40008 = ~n39653 & n39975;
  assign n40009 = ~n39787 & ~n40008;
  assign n40010 = ~n40007 & ~n40009;
  assign n40011 = n39795 & ~n40010;
  assign n40012 = ~n39997 & ~n40011;
  assign n40013 = ~pi213 & n40012;
  assign n40014 = ~pi209 & ~n40013;
  assign n40015 = ~n39983 & n40014;
  assign n40016 = ~n39888 & ~n40015;
  assign n40017 = pi230 & ~n40016;
  assign n40018 = ~pi230 & ~pi240;
  assign po397 = ~n40017 & ~n40018;
  assign n40020 = n39338 & n39452;
  assign n40021 = n39505 & ~n40020;
  assign n40022 = pi1152 & ~n40021;
  assign n40023 = ~po1038 & ~n40022;
  assign n40024 = n39457 & ~n40023;
  assign n40025 = n39264 & n39295;
  assign n40026 = n38230 & n39726;
  assign n40027 = ~n39245 & ~n40026;
  assign n40028 = n39457 & ~n40027;
  assign n40029 = ~n40025 & ~n40028;
  assign n40030 = ~pi1152 & ~n40029;
  assign n40031 = pi1152 & n39295;
  assign n40032 = n39331 & n40031;
  assign n40033 = ~n40030 & ~n40032;
  assign n40034 = ~n40024 & n40033;
  assign n40035 = ~pi1150 & ~n40034;
  assign n40036 = pi1151 & ~n39403;
  assign n40037 = pi219 & ~n39264;
  assign n40038 = ~po1038 & ~n40037;
  assign n40039 = ~n39695 & ~n40038;
  assign n40040 = ~pi214 & n39252;
  assign n40041 = pi212 & ~n40040;
  assign n40042 = ~n39711 & n40041;
  assign n40043 = n39269 & ~n39709;
  assign n40044 = ~n40042 & ~n40043;
  assign n40045 = ~n39261 & ~n40044;
  assign n40046 = ~pi219 & ~n40045;
  assign n40047 = ~pi1152 & ~n39828;
  assign n40048 = ~n40046 & n40047;
  assign n40049 = n39269 & ~n39515;
  assign n40050 = ~pi219 & ~n40049;
  assign n40051 = pi212 & n39338;
  assign n40052 = n40050 & ~n40051;
  assign n40053 = pi1152 & ~n40052;
  assign n40054 = ~n39870 & n40050;
  assign n40055 = n40053 & ~n40054;
  assign n40056 = ~n40048 & ~n40055;
  assign n40057 = ~n40039 & ~n40056;
  assign n40058 = n40036 & ~n40057;
  assign n40059 = ~pi1151 & ~n39664;
  assign n40060 = ~n39264 & n39493;
  assign n40061 = ~pi299 & n40060;
  assign n40062 = ~n39757 & ~n40061;
  assign n40063 = n40038 & n40062;
  assign n40064 = ~pi1152 & ~n40063;
  assign n40065 = ~n39331 & ~n40062;
  assign n40066 = n39526 & ~n40065;
  assign n40067 = pi1152 & ~n40066;
  assign n40068 = ~n40064 & ~n40067;
  assign n40069 = n40059 & ~n40068;
  assign n40070 = pi1150 & ~n40069;
  assign n40071 = ~n40058 & n40070;
  assign n40072 = ~n40035 & ~n40071;
  assign n40073 = ~pi1149 & ~n40072;
  assign n40074 = ~n38425 & n39338;
  assign n40075 = pi212 & n39505;
  assign n40076 = ~n40074 & n40075;
  assign n40077 = ~n39509 & ~n40076;
  assign n40078 = ~pi219 & ~n40077;
  assign n40079 = pi1152 & ~n40078;
  assign n40080 = n39512 & n40079;
  assign n40081 = ~pi214 & ~n39483;
  assign n40082 = n39477 & ~n40081;
  assign n40083 = ~pi212 & ~n39484;
  assign n40084 = ~n40082 & ~n40083;
  assign n40085 = ~pi219 & ~n40084;
  assign n40086 = ~pi1152 & n39486;
  assign n40087 = ~n40085 & n40086;
  assign n40088 = n39455 & ~n40087;
  assign n40089 = ~n40080 & n40088;
  assign n40090 = ~n39331 & n39493;
  assign n40091 = pi219 & ~n39482;
  assign n40092 = n39652 & ~n40091;
  assign n40093 = ~n40038 & ~n40092;
  assign n40094 = ~n39526 & n40093;
  assign n40095 = pi1152 & ~n40094;
  assign n40096 = ~n40090 & n40095;
  assign n40097 = ~pi1151 & ~n39407;
  assign n40098 = ~n40060 & ~n40093;
  assign n40099 = ~pi1152 & n40098;
  assign n40100 = n40097 & ~n40099;
  assign n40101 = ~n40096 & n40100;
  assign n40102 = ~pi1150 & ~n40101;
  assign n40103 = ~n40089 & n40102;
  assign n40104 = n39512 & n40053;
  assign n40105 = pi1151 & ~n39656;
  assign n40106 = ~n39261 & ~n39278;
  assign n40107 = ~pi219 & ~n40106;
  assign n40108 = n40086 & ~n40107;
  assign n40109 = n40105 & ~n40108;
  assign n40110 = ~n40104 & n40109;
  assign n40111 = ~pi1151 & ~n39696;
  assign n40112 = pi211 & ~n39638;
  assign n40113 = ~n38703 & ~n40112;
  assign n40114 = ~n39636 & ~n40113;
  assign n40115 = ~n39751 & ~n40114;
  assign n40116 = ~n39320 & ~n40115;
  assign n40117 = ~pi219 & ~n40116;
  assign n40118 = ~n40094 & ~n40117;
  assign n40119 = pi1152 & ~n40118;
  assign n40120 = n40064 & ~n40098;
  assign n40121 = ~n40119 & ~n40120;
  assign n40122 = n40111 & ~n40121;
  assign n40123 = pi1150 & ~n40122;
  assign n40124 = ~n40110 & n40123;
  assign n40125 = ~n40103 & ~n40124;
  assign n40126 = pi1149 & ~n40125;
  assign n40127 = ~n40073 & ~n40126;
  assign n40128 = ~pi213 & ~n40127;
  assign n40129 = pi213 & ~n39538;
  assign n40130 = pi209 & ~n40129;
  assign n40131 = ~n40128 & n40130;
  assign n40132 = ~n38357 & n39274;
  assign n40133 = n11050 & ~n40132;
  assign n40134 = n39722 & ~n40133;
  assign n40135 = ~n39459 & ~n40134;
  assign n40136 = pi299 & n39239;
  assign n40137 = ~n39743 & ~n40026;
  assign n40138 = ~po1038 & ~n40137;
  assign n40139 = ~n40136 & n40138;
  assign n40140 = n39462 & ~n40139;
  assign n40141 = ~pi1152 & ~n40140;
  assign n40142 = ~n40135 & n40141;
  assign n40143 = ~n39707 & ~n39709;
  assign n40144 = ~pi219 & ~n39877;
  assign n40145 = ~n39279 & n40144;
  assign n40146 = ~n40143 & n40145;
  assign n40147 = n39721 & ~n40146;
  assign n40148 = n39409 & ~n40147;
  assign n40149 = ~n39651 & ~n39743;
  assign n40150 = ~n38256 & n39405;
  assign n40151 = ~n40149 & ~n40150;
  assign n40152 = ~pi219 & ~n40151;
  assign n40153 = pi219 & ~n39743;
  assign n40154 = ~po1038 & ~n40153;
  assign n40155 = ~n40152 & n40154;
  assign n40156 = n39429 & ~n40155;
  assign n40157 = pi1152 & ~n40156;
  assign n40158 = ~n40148 & n40157;
  assign n40159 = ~pi1150 & ~n40158;
  assign n40160 = ~n40142 & n40159;
  assign n40161 = ~pi219 & ~n39265;
  assign n40162 = ~n39877 & n40161;
  assign n40163 = ~pi1153 & n40162;
  assign n40164 = pi299 & n10427;
  assign n40165 = ~pi219 & ~n40164;
  assign n40166 = n40092 & ~n40165;
  assign n40167 = ~n39879 & ~n40166;
  assign n40168 = ~n40163 & ~n40167;
  assign n40169 = ~pi211 & n40162;
  assign n40170 = ~n39655 & ~n40169;
  assign n40171 = n39409 & ~n40170;
  assign n40172 = ~n40168 & n40171;
  assign n40173 = ~po1038 & ~n39352;
  assign n40174 = ~pi299 & ~n39266;
  assign n40175 = ~n38145 & ~n40136;
  assign n40176 = ~n40174 & n40175;
  assign n40177 = n10669 & ~n39735;
  assign n40178 = n39803 & ~n40177;
  assign n40179 = ~n40176 & n40178;
  assign n40180 = n40173 & ~n40179;
  assign n40181 = n39429 & ~n40180;
  assign n40182 = pi1152 & ~n40181;
  assign n40183 = ~n40172 & n40182;
  assign n40184 = ~n39459 & ~n40168;
  assign n40185 = pi1153 & n40026;
  assign n40186 = n39462 & ~n40185;
  assign n40187 = ~pi1152 & ~n40186;
  assign n40188 = ~pi1151 & ~n39695;
  assign n40189 = ~pi1152 & ~n40188;
  assign n40190 = ~n40187 & ~n40189;
  assign n40191 = ~n40184 & ~n40190;
  assign n40192 = pi1150 & ~n40191;
  assign n40193 = ~n40183 & n40192;
  assign n40194 = pi1149 & ~n40193;
  assign n40195 = ~n40160 & n40194;
  assign n40196 = n39527 & ~n39751;
  assign n40197 = n39680 & ~n40196;
  assign n40198 = ~pi219 & ~n40197;
  assign n40199 = n39687 & ~n40198;
  assign n40200 = n39429 & ~n40199;
  assign n40201 = ~pi214 & n40113;
  assign n40202 = n39645 & ~n40201;
  assign n40203 = ~pi219 & ~n40202;
  assign n40204 = ~n40114 & n40203;
  assign n40205 = n39851 & ~n40204;
  assign n40206 = pi214 & n40113;
  assign n40207 = n39636 & ~n39641;
  assign n40208 = pi212 & ~n40207;
  assign n40209 = ~n40206 & n40208;
  assign n40210 = n39637 & ~n39644;
  assign n40211 = ~pi219 & ~n40210;
  assign n40212 = ~n40209 & n40211;
  assign n40213 = n39851 & ~n40212;
  assign n40214 = ~pi1153 & n40204;
  assign n40215 = n40213 & ~n40214;
  assign n40216 = ~n40205 & ~n40215;
  assign n40217 = n39409 & n40216;
  assign n40218 = pi1152 & ~n40217;
  assign n40219 = ~n40200 & n40218;
  assign n40220 = ~n39459 & ~n40215;
  assign n40221 = n39463 & ~n39675;
  assign n40222 = n39310 & ~n39463;
  assign n40223 = ~po1038 & ~n40222;
  assign n40224 = ~n40221 & n40223;
  assign n40225 = ~po1038 & ~n38357;
  assign n40226 = ~n40224 & n40225;
  assign n40227 = n39462 & ~n40226;
  assign n40228 = ~pi1152 & ~n40227;
  assign n40229 = ~n40220 & n40228;
  assign n40230 = pi1150 & ~n40229;
  assign n40231 = ~n40219 & n40230;
  assign n40232 = pi219 & ~n39299;
  assign n40233 = ~po1038 & ~n40232;
  assign n40234 = ~n39751 & n39756;
  assign n40235 = n40233 & ~n40234;
  assign n40236 = ~n39497 & n40233;
  assign n40237 = n39409 & ~n40236;
  assign n40238 = ~n40235 & n40237;
  assign n40239 = pi299 & n39402;
  assign n40240 = ~n39405 & n40239;
  assign n40241 = n39429 & ~n40240;
  assign n40242 = pi1152 & ~n40241;
  assign n40243 = ~n40238 & n40242;
  assign n40244 = ~n39459 & ~n40236;
  assign n40245 = n40187 & ~n40244;
  assign n40246 = ~pi1150 & ~n40245;
  assign n40247 = ~n40243 & n40246;
  assign n40248 = ~pi1149 & ~n40247;
  assign n40249 = ~n40231 & n40248;
  assign n40250 = ~n40195 & ~n40249;
  assign n40251 = pi213 & ~n40250;
  assign n40252 = ~n39688 & n40059;
  assign n40253 = ~n39648 & n40036;
  assign n40254 = pi1150 & ~n40253;
  assign n40255 = ~n40252 & n40254;
  assign n40256 = ~pi1150 & pi1151;
  assign n40257 = ~n39729 & n40256;
  assign n40258 = ~pi1149 & ~n40257;
  assign n40259 = ~n40255 & n40258;
  assign n40260 = n39455 & ~n39722;
  assign n40261 = ~n39761 & n40097;
  assign n40262 = ~pi1150 & ~n40261;
  assign n40263 = ~n40260 & n40262;
  assign n40264 = ~pi1151 & n39698;
  assign n40265 = n39655 & n40105;
  assign n40266 = pi1150 & ~n40265;
  assign n40267 = ~n40264 & n40266;
  assign n40268 = pi1149 & ~n40267;
  assign n40269 = ~n40263 & n40268;
  assign n40270 = ~n40259 & ~n40269;
  assign n40271 = ~pi213 & n40270;
  assign n40272 = ~pi209 & ~n40271;
  assign n40273 = ~n40251 & n40272;
  assign n40274 = ~n40131 & ~n40273;
  assign n40275 = pi230 & ~n40274;
  assign n40276 = ~pi230 & ~pi241;
  assign po398 = ~n40275 & ~n40276;
  assign n40278 = ~pi230 & ~pi242;
  assign n40279 = ~pi299 & ~n39014;
  assign n40280 = pi199 & pi1144;
  assign n40281 = ~pi200 & ~n40280;
  assign n40282 = ~n39012 & n40281;
  assign n40283 = n40279 & ~n40282;
  assign n40284 = pi207 & ~n40283;
  assign n40285 = ~n39891 & n40281;
  assign n40286 = ~pi299 & ~n39893;
  assign n40287 = ~n40285 & n40286;
  assign n40288 = ~pi207 & ~n40287;
  assign n40289 = pi208 & ~n40288;
  assign n40290 = ~n40284 & n40289;
  assign n40291 = n38512 & n40287;
  assign n40292 = ~n40290 & ~n40291;
  assign n40293 = ~n39804 & n40292;
  assign n40294 = ~pi214 & n40293;
  assign n40295 = ~n38454 & n40292;
  assign n40296 = pi211 & ~n40295;
  assign n40297 = ~n39185 & n40292;
  assign n40298 = ~pi211 & ~n40297;
  assign n40299 = pi214 & ~n40298;
  assign n40300 = ~n40296 & n40299;
  assign n40301 = pi212 & ~n40300;
  assign n40302 = ~n40294 & n40301;
  assign n40303 = ~pi214 & n40292;
  assign n40304 = ~pi212 & ~n40303;
  assign n40305 = ~n40293 & n40304;
  assign n40306 = ~pi219 & ~n40305;
  assign n40307 = ~n40302 & n40306;
  assign n40308 = ~n38136 & ~n40292;
  assign n40309 = pi219 & ~n40308;
  assign n40310 = n38136 & ~n40295;
  assign n40311 = n40309 & ~n40310;
  assign n40312 = ~po1038 & ~n40311;
  assign n40313 = ~n40307 & n40312;
  assign n40314 = pi214 & ~n38996;
  assign n40315 = ~pi214 & ~n39772;
  assign n40316 = ~n40314 & ~n40315;
  assign n40317 = pi212 & ~n40316;
  assign n40318 = ~pi212 & n39773;
  assign n40319 = ~pi219 & ~n40318;
  assign n40320 = ~n40317 & n40319;
  assign n40321 = pi219 & ~n38141;
  assign n40322 = ~n38137 & ~n40321;
  assign n40323 = ~n40320 & n40322;
  assign n40324 = po1038 & n40323;
  assign n40325 = ~n40313 & ~n40324;
  assign n40326 = pi213 & n40325;
  assign n40327 = pi211 & ~n40291;
  assign n40328 = n38171 & n40287;
  assign n40329 = n38136 & ~n38478;
  assign n40330 = ~n40328 & n40329;
  assign n40331 = ~n40327 & ~n40330;
  assign n40332 = pi219 & ~n40331;
  assign n40333 = n38135 & ~n40291;
  assign n40334 = n10669 & ~n38182;
  assign n40335 = ~n38153 & n38468;
  assign n40336 = ~n40334 & ~n40335;
  assign n40337 = ~pi219 & ~n40328;
  assign n40338 = ~n40336 & n40337;
  assign n40339 = ~n40333 & ~n40338;
  assign n40340 = ~n40332 & n40339;
  assign n40341 = ~n40290 & ~n40340;
  assign n40342 = ~po1038 & ~n40341;
  assign n40343 = ~pi213 & ~n38152;
  assign n40344 = ~n40342 & n40343;
  assign n40345 = ~n40326 & ~n40344;
  assign n40346 = pi209 & ~n40345;
  assign n40347 = ~pi213 & ~n38198;
  assign n40348 = pi299 & ~n40323;
  assign n40349 = ~po1038 & ~n40348;
  assign n40350 = ~n38189 & n40349;
  assign n40351 = ~n40324 & ~n40350;
  assign n40352 = pi213 & ~n40351;
  assign n40353 = ~pi209 & ~n40352;
  assign n40354 = ~n40347 & n40353;
  assign n40355 = ~n40346 & ~n40354;
  assign n40356 = pi230 & ~n40355;
  assign po399 = ~n40278 & ~n40356;
  assign n40358 = pi243 & ~pi1091;
  assign n40359 = ~pi83 & ~pi85;
  assign n40360 = pi314 & ~n40359;
  assign n40361 = pi802 & n40360;
  assign n40362 = pi276 & n40361;
  assign n40363 = ~pi1091 & ~n40362;
  assign n40364 = pi271 & ~n40363;
  assign n40365 = ~pi1091 & ~n40364;
  assign n40366 = pi273 & ~n40365;
  assign n40367 = ~pi1091 & ~n40366;
  assign n40368 = ~pi200 & ~n40367;
  assign n40369 = pi199 & ~n40367;
  assign n40370 = ~pi81 & n40359;
  assign n40371 = pi314 & ~n40370;
  assign n40372 = pi802 & n40371;
  assign n40373 = pi276 & n40372;
  assign n40374 = ~pi1091 & n40373;
  assign n40375 = pi271 & n40374;
  assign n40376 = pi273 & n40375;
  assign n40377 = ~n40366 & ~n40376;
  assign n40378 = ~pi1091 & n40377;
  assign n40379 = ~pi199 & ~n40378;
  assign n40380 = ~n40369 & ~n40379;
  assign n40381 = n40374 & ~n40380;
  assign n40382 = ~pi299 & ~n40381;
  assign n40383 = ~n40369 & n40382;
  assign n40384 = ~n40368 & n40383;
  assign n40385 = pi299 & ~n40376;
  assign n40386 = ~n40384 & ~n40385;
  assign n40387 = ~n40358 & ~n40386;
  assign n40388 = ~pi200 & ~n40374;
  assign n40389 = ~n40380 & ~n40388;
  assign n40390 = ~pi299 & ~n40389;
  assign n40391 = ~n40369 & n40390;
  assign n40392 = ~pi1091 & n40362;
  assign n40393 = pi271 & n40392;
  assign n40394 = pi273 & n40393;
  assign n40395 = pi299 & ~n40394;
  assign n40396 = ~n40368 & n40382;
  assign n40397 = ~n40379 & n40396;
  assign n40398 = ~n40395 & ~n40397;
  assign n40399 = ~n40391 & n40398;
  assign n40400 = pi299 & n40367;
  assign n40401 = ~n40396 & ~n40400;
  assign n40402 = pi243 & ~n40401;
  assign n40403 = ~n40399 & n40402;
  assign n40404 = pi1155 & ~n40403;
  assign n40405 = ~n40376 & n40400;
  assign n40406 = ~n40397 & ~n40405;
  assign n40407 = pi1155 & n40406;
  assign n40408 = ~n40404 & ~n40407;
  assign n40409 = ~n40385 & ~n40390;
  assign n40410 = ~pi243 & n40409;
  assign n40411 = ~n40384 & n40410;
  assign n40412 = ~n40408 & ~n40411;
  assign n40413 = ~n40379 & n40390;
  assign n40414 = ~n40384 & ~n40413;
  assign n40415 = ~n40405 & n40414;
  assign n40416 = ~pi243 & ~n40415;
  assign n40417 = ~n40385 & ~n40391;
  assign n40418 = pi243 & ~n40397;
  assign n40419 = n40417 & n40418;
  assign n40420 = ~n40416 & ~n40419;
  assign n40421 = ~pi1155 & ~n40420;
  assign n40422 = ~n40412 & ~n40421;
  assign n40423 = ~n40387 & n40422;
  assign n40424 = pi1156 & ~n40423;
  assign n40425 = ~n40400 & ~n40413;
  assign n40426 = ~pi243 & ~n40425;
  assign n40427 = ~pi1155 & ~n40426;
  assign n40428 = ~n40382 & ~n40385;
  assign n40429 = ~pi1155 & n40428;
  assign n40430 = ~n40427 & ~n40429;
  assign n40431 = ~n40385 & ~n40396;
  assign n40432 = pi243 & n40431;
  assign n40433 = ~n40383 & n40432;
  assign n40434 = ~n40430 & ~n40433;
  assign n40435 = ~pi1156 & ~n40434;
  assign n40436 = ~n40390 & ~n40405;
  assign n40437 = ~pi243 & ~n40436;
  assign n40438 = pi1155 & ~n40437;
  assign n40439 = ~n40432 & n40438;
  assign n40440 = n40435 & ~n40439;
  assign n40441 = pi1157 & ~n40440;
  assign n40442 = ~n40424 & n40441;
  assign n40443 = ~n40379 & n40382;
  assign n40444 = ~n40405 & ~n40443;
  assign n40445 = pi243 & ~n40444;
  assign n40446 = ~n40383 & ~n40385;
  assign n40447 = ~pi243 & n40446;
  assign n40448 = ~n40445 & ~n40447;
  assign n40449 = ~pi1091 & n40448;
  assign n40450 = ~pi1155 & ~n40449;
  assign n40451 = ~pi1156 & ~n40450;
  assign n40452 = pi1155 & ~n40358;
  assign n40453 = n40369 & n40452;
  assign n40454 = ~n40439 & ~n40453;
  assign n40455 = n40451 & n40454;
  assign n40456 = ~pi1155 & n40431;
  assign n40457 = ~n40374 & n40456;
  assign n40458 = pi1156 & ~n40457;
  assign n40459 = n40448 & n40458;
  assign n40460 = ~pi1157 & ~n40459;
  assign n40461 = ~n40455 & n40460;
  assign n40462 = pi211 & ~n40461;
  assign n40463 = ~n40442 & n40462;
  assign n40464 = pi1156 & ~n40422;
  assign n40465 = ~n40396 & ~n40405;
  assign n40466 = pi243 & ~n40465;
  assign n40467 = ~n40410 & ~n40466;
  assign n40468 = n40435 & n40467;
  assign n40469 = pi1157 & ~n40468;
  assign n40470 = ~n40464 & n40469;
  assign n40471 = n40448 & n40467;
  assign n40472 = pi1155 & ~n40471;
  assign n40473 = n40451 & ~n40472;
  assign n40474 = ~pi1155 & n40465;
  assign n40475 = ~n40409 & n40474;
  assign n40476 = n40459 & ~n40475;
  assign n40477 = ~pi1157 & ~n40476;
  assign n40478 = ~n40473 & n40477;
  assign n40479 = ~pi211 & ~n40478;
  assign n40480 = ~n40470 & n40479;
  assign n40481 = ~pi219 & ~n40480;
  assign n40482 = ~n40463 & n40481;
  assign n40483 = pi253 & pi254;
  assign n40484 = pi267 & n40483;
  assign n40485 = ~pi263 & n40484;
  assign n40486 = ~n40384 & ~n40400;
  assign n40487 = ~pi243 & n40486;
  assign n40488 = ~n40390 & ~n40395;
  assign n40489 = n40487 & n40488;
  assign n40490 = n40404 & ~n40489;
  assign n40491 = pi243 & ~n40399;
  assign n40492 = ~n40487 & ~n40491;
  assign n40493 = ~n40387 & ~n40426;
  assign n40494 = ~n40492 & n40493;
  assign n40495 = ~pi1155 & ~n40494;
  assign n40496 = ~n40490 & ~n40495;
  assign n40497 = pi1156 & ~n40496;
  assign n40498 = ~n40395 & ~n40413;
  assign n40499 = ~pi243 & ~n40498;
  assign n40500 = pi243 & ~n40383;
  assign n40501 = ~pi1155 & ~n40500;
  assign n40502 = ~n40499 & n40501;
  assign n40503 = ~pi243 & pi1155;
  assign n40504 = n40488 & n40503;
  assign n40505 = ~pi1156 & ~n40504;
  assign n40506 = ~n40402 & n40505;
  assign n40507 = ~n40502 & n40506;
  assign n40508 = n38210 & ~n40507;
  assign n40509 = ~n40497 & n40508;
  assign n40510 = pi243 & n40398;
  assign n40511 = n40438 & ~n40510;
  assign n40512 = ~n40427 & ~n40511;
  assign n40513 = ~n40492 & ~n40512;
  assign n40514 = pi1156 & ~n40513;
  assign n40515 = ~n40395 & ~n40396;
  assign n40516 = pi243 & n40515;
  assign n40517 = ~n40437 & ~n40516;
  assign n40518 = pi1155 & ~n40517;
  assign n40519 = ~n40383 & n40515;
  assign n40520 = pi243 & n40519;
  assign n40521 = ~n40426 & ~n40520;
  assign n40522 = ~n40518 & n40521;
  assign n40523 = ~pi1156 & ~n40522;
  assign n40524 = n39026 & ~n40523;
  assign n40525 = ~n40514 & n40524;
  assign n40526 = ~n40395 & ~n40443;
  assign n40527 = pi1155 & n40526;
  assign n40528 = ~n40390 & n40526;
  assign n40529 = ~n40527 & ~n40528;
  assign n40530 = pi243 & ~n40529;
  assign n40531 = ~n40383 & ~n40400;
  assign n40532 = ~pi243 & ~n40531;
  assign n40533 = ~n40457 & n40532;
  assign n40534 = ~n40530 & ~n40533;
  assign n40535 = pi1156 & ~n40534;
  assign n40536 = ~n40443 & n40516;
  assign n40537 = ~n40391 & ~n40400;
  assign n40538 = ~pi243 & ~n40537;
  assign n40539 = pi1155 & ~n40538;
  assign n40540 = ~n40536 & n40539;
  assign n40541 = ~pi243 & ~pi1091;
  assign n40542 = ~n40382 & ~n40395;
  assign n40543 = n40541 & ~n40542;
  assign n40544 = ~pi1155 & ~n40543;
  assign n40545 = pi243 & n40542;
  assign n40546 = n40544 & ~n40545;
  assign n40547 = ~pi1156 & ~n40546;
  assign n40548 = ~n40540 & n40547;
  assign n40549 = ~pi1157 & ~n40548;
  assign n40550 = ~n40535 & n40549;
  assign n40551 = ~n40525 & ~n40550;
  assign n40552 = ~n40509 & n40551;
  assign n40553 = pi219 & ~n40552;
  assign n40554 = n40485 & ~n40553;
  assign n40555 = ~n40482 & n40554;
  assign n40556 = ~pi299 & pi1091;
  assign n40557 = n38527 & n40556;
  assign n40558 = ~n40541 & ~n40557;
  assign n40559 = pi1156 & ~n40558;
  assign n40560 = pi1156 & ~n38651;
  assign n40561 = pi1091 & ~n38620;
  assign n40562 = n40560 & n40561;
  assign n40563 = ~n40559 & ~n40562;
  assign n40564 = ~pi299 & n38328;
  assign n40565 = pi1091 & ~n40564;
  assign n40566 = ~n40358 & ~n40565;
  assign n40567 = ~n40452 & ~n40541;
  assign n40568 = n38270 & ~n40567;
  assign n40569 = ~n40566 & ~n40568;
  assign n40570 = ~pi1156 & ~n40569;
  assign n40571 = n40563 & ~n40570;
  assign n40572 = pi1157 & ~n40571;
  assign n40573 = pi199 & pi1091;
  assign n40574 = ~pi299 & n40573;
  assign n40575 = n40452 & ~n40574;
  assign n40576 = pi1156 & ~n40575;
  assign n40577 = ~pi1155 & ~n40358;
  assign n40578 = ~n11381 & n40556;
  assign n40579 = n40577 & ~n40578;
  assign n40580 = n40576 & ~n40579;
  assign n40581 = ~n40561 & ~n40567;
  assign n40582 = ~pi1156 & ~n40581;
  assign n40583 = ~pi1157 & ~n40582;
  assign n40584 = ~n40580 & n40583;
  assign n40585 = ~n40572 & ~n40584;
  assign n40586 = pi211 & ~n40585;
  assign n40587 = pi200 & pi1091;
  assign n40588 = ~pi299 & n40587;
  assign n40589 = n40452 & ~n40588;
  assign n40590 = ~n40566 & ~n40589;
  assign n40591 = ~n40559 & n40590;
  assign n40592 = pi1157 & n40591;
  assign n40593 = pi1091 & ~n11382;
  assign n40594 = n40577 & ~n40593;
  assign n40595 = ~n40575 & ~n40594;
  assign n40596 = pi200 & ~pi1156;
  assign n40597 = n40556 & n40596;
  assign n40598 = ~n40595 & ~n40597;
  assign n40599 = ~pi1157 & ~n40598;
  assign n40600 = ~pi211 & ~n40599;
  assign n40601 = ~n40592 & n40600;
  assign n40602 = ~n40586 & ~n40601;
  assign n40603 = ~pi219 & ~n40602;
  assign n40604 = n39026 & ~n40559;
  assign n40605 = ~n40570 & n40604;
  assign n40606 = pi219 & ~n40605;
  assign n40607 = pi299 & pi1091;
  assign n40608 = n40598 & ~n40607;
  assign n40609 = ~pi1157 & ~n40608;
  assign n40610 = pi1091 & n38329;
  assign n40611 = n40577 & ~n40610;
  assign n40612 = ~n40589 & ~n40611;
  assign n40613 = ~pi1156 & ~n40612;
  assign n40614 = n38210 & ~n40613;
  assign n40615 = n40563 & n40614;
  assign n40616 = ~n40609 & ~n40615;
  assign n40617 = n40606 & n40616;
  assign n40618 = ~n40603 & ~n40617;
  assign n40619 = ~n40485 & ~n40618;
  assign n40620 = ~po1038 & ~n40619;
  assign n40621 = ~n40555 & n40620;
  assign n40622 = ~pi243 & n40367;
  assign n40623 = pi243 & n40394;
  assign n40624 = n38210 & ~n40358;
  assign n40625 = ~n40392 & n40624;
  assign n40626 = ~n40623 & ~n40625;
  assign n40627 = ~n40622 & n40626;
  assign n40628 = pi219 & ~n40627;
  assign n40629 = n40358 & n40377;
  assign n40630 = ~pi243 & n40376;
  assign n40631 = ~n38204 & ~n38211;
  assign n40632 = pi1091 & n40631;
  assign n40633 = ~pi219 & ~n40632;
  assign n40634 = ~n40630 & n40633;
  assign n40635 = ~n40629 & n40634;
  assign n40636 = ~n40628 & ~n40635;
  assign n40637 = n40485 & ~n40636;
  assign n40638 = ~pi219 & ~n40631;
  assign n40639 = pi1157 & n38241;
  assign n40640 = ~n40638 & ~n40639;
  assign n40641 = pi1091 & ~n40640;
  assign n40642 = ~n40541 & ~n40641;
  assign n40643 = ~n40485 & ~n40642;
  assign n40644 = po1038 & ~n40643;
  assign n40645 = ~n40637 & n40644;
  assign n40646 = pi272 & pi283;
  assign n40647 = pi275 & n40646;
  assign n40648 = pi268 & n40647;
  assign n40649 = ~n40645 & n40648;
  assign n40650 = ~n40621 & n40649;
  assign n40651 = ~po1038 & n40618;
  assign n40652 = po1038 & n40642;
  assign n40653 = ~n40648 & ~n40652;
  assign n40654 = ~n40651 & n40653;
  assign n40655 = ~pi230 & ~n40654;
  assign n40656 = ~n40650 & n40655;
  assign n40657 = pi199 & ~n39188;
  assign n40658 = ~n38526 & ~n40596;
  assign n40659 = ~n40657 & n40658;
  assign n40660 = n16361 & n40659;
  assign n40661 = ~n16361 & ~n40640;
  assign n40662 = pi230 & ~n40661;
  assign n40663 = ~n40660 & n40662;
  assign po400 = ~n40656 & ~n40663;
  assign n40665 = ~pi230 & ~pi244;
  assign n40666 = pi213 & ~n40012;
  assign n40667 = pi299 & ~n38996;
  assign n40668 = ~n39906 & ~n40667;
  assign n40669 = ~pi214 & n40668;
  assign n40670 = n38142 & n39871;
  assign n40671 = pi212 & ~n40670;
  assign n40672 = ~n40669 & n40671;
  assign n40673 = ~n39918 & n40672;
  assign n40674 = n39934 & ~n40668;
  assign n40675 = ~n39959 & n40674;
  assign n40676 = ~pi219 & ~n40675;
  assign n40677 = ~n40673 & n40676;
  assign n40678 = n38136 & n38437;
  assign n40679 = ~n39963 & ~n40678;
  assign n40680 = n39902 & ~n40679;
  assign n40681 = ~n40677 & n40680;
  assign n40682 = ~n39911 & n40672;
  assign n40683 = ~pi219 & ~n40674;
  assign n40684 = ~n40682 & n40683;
  assign n40685 = pi299 & n39002;
  assign n40686 = pi1147 & ~n40685;
  assign n40687 = n39915 & n40686;
  assign n40688 = ~n40684 & n40687;
  assign n40689 = ~pi213 & ~n39004;
  assign n40690 = ~n40688 & n40689;
  assign n40691 = ~n40681 & n40690;
  assign n40692 = ~n40666 & ~n40691;
  assign n40693 = pi209 & ~n40692;
  assign n40694 = n39784 & ~n39790;
  assign n40695 = ~n39795 & ~n40694;
  assign n40696 = n39784 & ~n39789;
  assign n40697 = n10669 & ~n39804;
  assign n40698 = ~n10669 & n39799;
  assign n40699 = n38474 & ~n40698;
  assign n40700 = ~n40697 & n40699;
  assign n40701 = ~n40696 & n40700;
  assign n40702 = ~n39018 & ~n39818;
  assign n40703 = ~n40701 & n40702;
  assign n40704 = ~po1038 & ~n40703;
  assign n40705 = ~n40695 & ~n40704;
  assign n40706 = pi213 & ~n40705;
  assign n40707 = ~pi213 & ~n39024;
  assign n40708 = ~pi209 & ~n40707;
  assign n40709 = ~n40706 & n40708;
  assign n40710 = ~n40693 & ~n40709;
  assign n40711 = pi230 & ~n40710;
  assign po401 = ~n40665 & ~n40711;
  assign n40713 = pi1146 & n39407;
  assign n40714 = pi1147 & ~n39403;
  assign n40715 = ~n40713 & n40714;
  assign n40716 = ~n39797 & n40292;
  assign n40717 = n38136 & ~n40716;
  assign n40718 = n40309 & ~n40717;
  assign n40719 = ~po1038 & ~n40718;
  assign n40720 = ~pi299 & n40297;
  assign n40721 = ~pi211 & ~n40720;
  assign n40722 = n40292 & ~n40721;
  assign n40723 = pi214 & ~n39798;
  assign n40724 = pi299 & ~n40723;
  assign n40725 = n40722 & ~n40724;
  assign n40726 = pi212 & ~n40725;
  assign n40727 = n40304 & ~n40720;
  assign n40728 = ~pi219 & ~n40727;
  assign n40729 = ~n40726 & n40728;
  assign n40730 = n40719 & ~n40729;
  assign n40731 = n40715 & ~n40730;
  assign n40732 = ~pi1147 & ~n40713;
  assign n40733 = ~n39453 & n40732;
  assign n40734 = n40292 & n40723;
  assign n40735 = pi212 & ~n40734;
  assign n40736 = ~pi214 & n40722;
  assign n40737 = n40735 & ~n40736;
  assign n40738 = n40304 & ~n40722;
  assign n40739 = ~pi219 & ~n40738;
  assign n40740 = ~n40737 & n40739;
  assign n40741 = n40719 & ~n40740;
  assign n40742 = n40733 & ~n40741;
  assign n40743 = pi1148 & ~n40742;
  assign n40744 = ~n40731 & n40743;
  assign n40745 = ~pi219 & ~n39774;
  assign n40746 = n40292 & n40745;
  assign n40747 = n40741 & ~n40746;
  assign n40748 = n40732 & ~n40747;
  assign n40749 = ~n39968 & ~n40715;
  assign n40750 = ~n12978 & n40292;
  assign n40751 = n40304 & ~n40750;
  assign n40752 = ~pi219 & ~n40751;
  assign n40753 = ~pi214 & n40750;
  assign n40754 = n40726 & ~n40753;
  assign n40755 = n40752 & ~n40754;
  assign n40756 = n40719 & ~n40755;
  assign n40757 = ~n40749 & ~n40756;
  assign n40758 = ~pi1148 & ~n40757;
  assign n40759 = ~n40748 & n40758;
  assign n40760 = ~n40744 & ~n40759;
  assign n40761 = pi213 & ~n40760;
  assign n40762 = ~pi213 & ~n40325;
  assign n40763 = ~pi209 & ~n40762;
  assign n40764 = ~n40761 & n40763;
  assign n40765 = pi199 & pi1146;
  assign n40766 = n38328 & ~n40765;
  assign n40767 = ~pi299 & ~n40766;
  assign n40768 = n39066 & n40767;
  assign n40769 = ~pi200 & ~n40765;
  assign n40770 = n39898 & ~n40769;
  assign n40771 = n39741 & n40770;
  assign n40772 = ~n39797 & ~n40771;
  assign n40773 = ~n40768 & n40772;
  assign n40774 = ~pi299 & ~n40773;
  assign n40775 = ~pi214 & ~n40774;
  assign n40776 = ~pi212 & ~n40775;
  assign n40777 = ~n10564 & ~n39066;
  assign n40778 = n40770 & ~n40777;
  assign n40779 = pi211 & ~n40778;
  assign n40780 = ~pi299 & ~n40770;
  assign n40781 = ~n40773 & ~n40780;
  assign n40782 = ~pi299 & ~n40781;
  assign n40783 = ~pi211 & n40782;
  assign n40784 = ~n40779 & ~n40783;
  assign n40785 = ~n40774 & ~n40784;
  assign n40786 = n40776 & ~n40785;
  assign n40787 = ~pi219 & ~n40786;
  assign n40788 = n40723 & ~n40774;
  assign n40789 = ~pi214 & n40785;
  assign n40790 = pi212 & ~n40789;
  assign n40791 = ~n40788 & n40790;
  assign n40792 = n40787 & ~n40791;
  assign n40793 = ~n38136 & n40774;
  assign n40794 = pi219 & ~n40793;
  assign n40795 = n38136 & ~n40773;
  assign n40796 = n40794 & ~n40795;
  assign n40797 = ~po1038 & ~n40796;
  assign n40798 = ~n40792 & n40797;
  assign n40799 = n40733 & ~n40798;
  assign n40800 = n39898 & ~n40766;
  assign n40801 = pi208 & n40800;
  assign n40802 = ~n38512 & ~n40801;
  assign n40803 = ~n38254 & n40767;
  assign n40804 = ~n40802 & n40803;
  assign n40805 = ~n10564 & n40769;
  assign n40806 = n40804 & ~n40805;
  assign n40807 = ~n39797 & ~n40806;
  assign n40808 = ~n38135 & n40806;
  assign n40809 = ~n38136 & ~n40808;
  assign n40810 = ~n40807 & ~n40809;
  assign n40811 = pi219 & ~n40804;
  assign n40812 = ~n40810 & n40811;
  assign n40813 = ~po1038 & ~n40812;
  assign n40814 = ~n40165 & ~n40745;
  assign n40815 = ~n40804 & ~n40814;
  assign n40816 = ~pi299 & n40807;
  assign n40817 = ~pi214 & ~n40804;
  assign n40818 = ~pi212 & ~n40817;
  assign n40819 = ~n39870 & ~n40818;
  assign n40820 = ~n40816 & ~n40819;
  assign n40821 = n40815 & ~n40820;
  assign n40822 = n40813 & ~n40821;
  assign n40823 = n40715 & ~n40822;
  assign n40824 = pi1148 & ~n40823;
  assign n40825 = ~n40799 & n40824;
  assign n40826 = ~n12978 & ~n40806;
  assign n40827 = pi214 & ~n40826;
  assign n40828 = ~pi214 & n40806;
  assign n40829 = ~pi212 & ~n40828;
  assign n40830 = ~n40827 & n40829;
  assign n40831 = ~pi214 & ~n40826;
  assign n40832 = pi214 & ~n40816;
  assign n40833 = ~pi299 & ~n40804;
  assign n40834 = ~pi211 & ~n40833;
  assign n40835 = ~n40804 & ~n40834;
  assign n40836 = n40832 & ~n40835;
  assign n40837 = pi212 & ~n40836;
  assign n40838 = ~n40831 & n40837;
  assign n40839 = ~n40830 & ~n40838;
  assign n40840 = ~pi219 & ~n40839;
  assign n40841 = ~pi1146 & ~n38425;
  assign n40842 = n39877 & ~n40841;
  assign n40843 = n40840 & ~n40842;
  assign n40844 = ~pi212 & n40828;
  assign n40845 = pi219 & ~n40844;
  assign n40846 = ~n40810 & n40845;
  assign n40847 = ~po1038 & ~n40846;
  assign n40848 = ~n40843 & n40847;
  assign n40849 = ~n40749 & ~n40848;
  assign n40850 = pi219 & ~n40778;
  assign n40851 = ~n38635 & ~n40850;
  assign n40852 = ~n38135 & ~n40779;
  assign n40853 = n40781 & n40852;
  assign n40854 = ~n40851 & ~n40853;
  assign n40855 = ~po1038 & ~n40854;
  assign n40856 = ~n40778 & ~n40814;
  assign n40857 = n40855 & ~n40856;
  assign n40858 = n40732 & ~n40857;
  assign n40859 = ~pi1148 & ~n40858;
  assign n40860 = ~n40849 & n40859;
  assign n40861 = ~n40825 & ~n40860;
  assign n40862 = pi213 & ~n40861;
  assign n40863 = ~pi214 & n40778;
  assign n40864 = ~n39804 & ~n40774;
  assign n40865 = pi214 & ~n40782;
  assign n40866 = ~n40864 & n40865;
  assign n40867 = ~n40863 & ~n40866;
  assign n40868 = ~pi212 & ~n40867;
  assign n40869 = pi299 & ~n40316;
  assign n40870 = ~n40774 & ~n40869;
  assign n40871 = pi212 & ~n40870;
  assign n40872 = ~n40780 & n40871;
  assign n40873 = ~pi219 & ~n40872;
  assign n40874 = ~n40868 & n40873;
  assign n40875 = ~n38135 & ~n38460;
  assign n40876 = n40784 & n40875;
  assign n40877 = ~n40851 & ~n40876;
  assign n40878 = n39902 & ~n40877;
  assign n40879 = ~n40874 & n40878;
  assign n40880 = ~n38454 & ~n40804;
  assign n40881 = ~n40809 & ~n40880;
  assign n40882 = n40820 & n40881;
  assign n40883 = n40845 & ~n40882;
  assign n40884 = pi1147 & ~po1038;
  assign n40885 = ~n40804 & ~n40869;
  assign n40886 = pi212 & ~n40885;
  assign n40887 = ~n40816 & n40886;
  assign n40888 = ~pi219 & ~n40887;
  assign n40889 = ~pi212 & n40804;
  assign n40890 = pi299 & n40318;
  assign n40891 = ~n40889 & ~n40890;
  assign n40892 = ~n40816 & ~n40891;
  assign n40893 = n40888 & ~n40892;
  assign n40894 = n40884 & ~n40893;
  assign n40895 = ~n40883 & n40894;
  assign n40896 = ~pi1148 & ~n40324;
  assign n40897 = ~n40895 & n40896;
  assign n40898 = ~n40879 & n40897;
  assign n40899 = ~pi299 & n40773;
  assign n40900 = n38136 & ~n40899;
  assign n40901 = ~n38460 & n40900;
  assign n40902 = n40794 & ~n40901;
  assign n40903 = n39902 & ~n40902;
  assign n40904 = ~n40774 & ~n40890;
  assign n40905 = n40873 & n40904;
  assign n40906 = n40903 & ~n40905;
  assign n40907 = ~pi219 & ~n40886;
  assign n40908 = n40891 & n40907;
  assign n40909 = ~n38136 & n40804;
  assign n40910 = pi219 & ~n40909;
  assign n40911 = ~n40881 & n40910;
  assign n40912 = n40884 & ~n40911;
  assign n40913 = ~n40908 & n40912;
  assign n40914 = pi1148 & ~n40324;
  assign n40915 = ~n40913 & n40914;
  assign n40916 = ~n40906 & n40915;
  assign n40917 = ~pi213 & ~n40916;
  assign n40918 = ~n40898 & n40917;
  assign n40919 = pi209 & ~n40918;
  assign n40920 = ~n40862 & n40919;
  assign n40921 = ~n40764 & ~n40920;
  assign n40922 = pi230 & ~n40921;
  assign n40923 = ~pi230 & ~pi245;
  assign po402 = ~n40922 & ~n40923;
  assign n40925 = ~n40715 & ~n40733;
  assign n40926 = pi219 & ~n39797;
  assign n40927 = n39652 & ~n40926;
  assign n40928 = n39695 & ~n39742;
  assign n40929 = ~n40927 & ~n40928;
  assign n40930 = ~n39744 & ~n39813;
  assign n40931 = n38145 & ~n40930;
  assign n40932 = ~n40149 & ~n40931;
  assign n40933 = ~pi219 & ~n40932;
  assign n40934 = ~n40929 & ~n40933;
  assign n40935 = ~n40925 & ~n40934;
  assign n40936 = ~pi212 & n39736;
  assign n40937 = ~pi219 & ~n40936;
  assign n40938 = ~n39752 & n39867;
  assign n40939 = n40937 & ~n40938;
  assign n40940 = ~n39745 & ~n40939;
  assign n40941 = n40733 & ~n40940;
  assign n40942 = ~pi1150 & ~n40941;
  assign n40943 = ~n40935 & n40942;
  assign n40944 = ~n39829 & ~n40927;
  assign n40945 = ~n39838 & n40041;
  assign n40946 = ~pi212 & ~n39244;
  assign n40947 = ~pi219 & ~n40946;
  assign n40948 = ~n39754 & n40947;
  assign n40949 = ~n40945 & n40948;
  assign n40950 = ~n40944 & ~n40949;
  assign n40951 = n40715 & ~n40950;
  assign n40952 = n40143 & n40945;
  assign n40953 = n39716 & ~n40952;
  assign n40954 = ~n40944 & ~n40953;
  assign n40955 = n40733 & ~n40954;
  assign n40956 = pi1150 & ~n40955;
  assign n40957 = ~n40951 & n40956;
  assign n40958 = ~n40943 & ~n40957;
  assign n40959 = pi1148 & ~n40958;
  assign n40960 = n40814 & n40927;
  assign n40961 = n40732 & ~n40960;
  assign n40962 = ~n40749 & ~n40927;
  assign n40963 = ~n40961 & ~n40962;
  assign n40964 = pi1150 & n39725;
  assign n40965 = ~n40963 & ~n40964;
  assign n40966 = pi1150 & n39263;
  assign n40967 = pi299 & ~n39663;
  assign n40968 = ~n40814 & ~n40967;
  assign n40969 = ~n40966 & n40968;
  assign n40970 = ~n40749 & n40969;
  assign n40971 = ~pi1148 & ~n40970;
  assign n40972 = ~n40965 & n40971;
  assign n40973 = ~n40959 & ~n40972;
  assign n40974 = ~pi1149 & ~n40973;
  assign n40975 = ~pi1146 & n39686;
  assign n40976 = n39652 & ~n39669;
  assign n40977 = ~n39687 & ~n40976;
  assign n40978 = ~n40975 & ~n40977;
  assign n40979 = n39685 & ~n40814;
  assign n40980 = n40978 & ~n40979;
  assign n40981 = ~n40749 & ~n40980;
  assign n40982 = ~n39310 & n40165;
  assign n40983 = ~n40977 & ~n40982;
  assign n40984 = ~pi1146 & ~n39310;
  assign n40985 = n40983 & ~n40984;
  assign n40986 = n40732 & ~n40985;
  assign n40987 = ~pi1150 & ~n40986;
  assign n40988 = ~n40981 & n40987;
  assign n40989 = ~n39852 & ~n40927;
  assign n40990 = ~n40204 & ~n40989;
  assign n40991 = ~n39647 & ~n40204;
  assign n40992 = ~n39797 & ~n40991;
  assign n40993 = n40990 & ~n40992;
  assign n40994 = ~n39634 & ~n40993;
  assign n40995 = n40213 & ~n40994;
  assign n40996 = n40732 & ~n40995;
  assign n40997 = ~n40749 & ~n40993;
  assign n40998 = pi1150 & ~n40997;
  assign n40999 = ~n40996 & n40998;
  assign n41000 = ~pi1148 & ~n40999;
  assign n41001 = ~n40988 & n41000;
  assign n41002 = ~n39695 & ~n40927;
  assign n41003 = ~n39735 & n40938;
  assign n41004 = ~n39738 & ~n41003;
  assign n41005 = ~n40733 & ~n41004;
  assign n41006 = ~pi214 & n39735;
  assign n41007 = pi212 & ~n41006;
  assign n41008 = ~n39266 & n40723;
  assign n41009 = n41007 & ~n41008;
  assign n41010 = n40937 & ~n41009;
  assign n41011 = ~n41005 & n41010;
  assign n41012 = ~n41002 & ~n41011;
  assign n41013 = ~n40925 & ~n41012;
  assign n41014 = ~pi1150 & ~n41013;
  assign n41015 = ~n39879 & ~n40960;
  assign n41016 = n40733 & n41015;
  assign n41017 = pi1146 & n39653;
  assign n41018 = n40715 & ~n41017;
  assign n41019 = ~n39876 & n41018;
  assign n41020 = pi1150 & ~n41019;
  assign n41021 = ~n41016 & n41020;
  assign n41022 = pi1148 & ~n41021;
  assign n41023 = ~n41014 & n41022;
  assign n41024 = pi1149 & ~n41023;
  assign n41025 = ~n41001 & n41024;
  assign n41026 = ~n40974 & ~n41025;
  assign n41027 = ~pi213 & ~n41026;
  assign n41028 = pi1150 & n39657;
  assign n41029 = ~pi1150 & n39698;
  assign n41030 = pi1149 & ~n41029;
  assign n41031 = ~n41028 & n41030;
  assign n41032 = pi1150 & n39723;
  assign n41033 = ~pi1150 & n39762;
  assign n41034 = ~pi1149 & ~n41033;
  assign n41035 = ~n41032 & n41034;
  assign n41036 = ~n41031 & ~n41035;
  assign n41037 = pi1148 & ~n41036;
  assign n41038 = ~pi1150 & n39689;
  assign n41039 = pi1150 & n39649;
  assign n41040 = pi1149 & ~n41039;
  assign n41041 = ~n41038 & n41040;
  assign n41042 = ~pi1149 & pi1150;
  assign n41043 = ~n39729 & n41042;
  assign n41044 = ~n41041 & ~n41043;
  assign n41045 = ~pi1148 & ~n41044;
  assign n41046 = ~n41037 & ~n41045;
  assign n41047 = pi213 & ~n41046;
  assign n41048 = pi209 & ~n41047;
  assign n41049 = ~n41027 & n41048;
  assign n41050 = ~pi212 & ~n40863;
  assign n41051 = ~n12978 & ~n40778;
  assign n41052 = pi214 & ~n41051;
  assign n41053 = n41050 & ~n41052;
  assign n41054 = ~pi214 & ~n41051;
  assign n41055 = pi214 & n40784;
  assign n41056 = pi212 & ~n41055;
  assign n41057 = ~n41054 & n41056;
  assign n41058 = ~n41053 & ~n41057;
  assign n41059 = ~pi219 & ~n41058;
  assign n41060 = n39902 & ~n40850;
  assign n41061 = ~n41059 & n41060;
  assign n41062 = pi219 & ~n40806;
  assign n41063 = n40884 & ~n41062;
  assign n41064 = ~n40840 & n41063;
  assign n41065 = ~pi1150 & ~n39664;
  assign n41066 = ~n41064 & n41065;
  assign n41067 = ~n41061 & n41066;
  assign n41068 = ~n40865 & n41050;
  assign n41069 = ~pi214 & ~n40782;
  assign n41070 = n41056 & ~n41069;
  assign n41071 = ~n41068 & ~n41070;
  assign n41072 = ~pi219 & ~n41071;
  assign n41073 = ~n40850 & ~n41072;
  assign n41074 = ~pi1147 & ~n41073;
  assign n41075 = ~pi219 & ~n40820;
  assign n41076 = ~n41062 & ~n41075;
  assign n41077 = pi1147 & ~n41076;
  assign n41078 = ~po1038 & ~n41077;
  assign n41079 = ~n41074 & n41078;
  assign n41080 = pi1150 & ~n39403;
  assign n41081 = ~n41079 & n41080;
  assign n41082 = ~n41067 & ~n41081;
  assign n41083 = pi1149 & ~n41082;
  assign n41084 = pi1150 & n39452;
  assign n41085 = ~pi1147 & n40781;
  assign n41086 = n16361 & ~n41085;
  assign n41087 = n41084 & ~n41086;
  assign n41088 = pi1147 & ~n40806;
  assign n41089 = n40778 & ~n41084;
  assign n41090 = ~pi1147 & ~n41089;
  assign n41091 = ~po1038 & ~n41090;
  assign n41092 = ~n41088 & n41091;
  assign n41093 = ~pi1149 & ~n41092;
  assign n41094 = ~n41087 & n41093;
  assign n41095 = ~n41083 & ~n41094;
  assign n41096 = ~pi1148 & ~n41095;
  assign n41097 = n40794 & ~n40900;
  assign n41098 = n39902 & ~n41097;
  assign n41099 = ~n40774 & n41051;
  assign n41100 = pi214 & n41099;
  assign n41101 = n40790 & ~n41100;
  assign n41102 = n40787 & ~n41101;
  assign n41103 = n41098 & ~n41102;
  assign n41104 = ~n38135 & n40834;
  assign n41105 = n40910 & ~n41104;
  assign n41106 = n40884 & ~n41105;
  assign n41107 = pi214 & ~n12978;
  assign n41108 = ~n40804 & n41107;
  assign n41109 = pi212 & ~n41108;
  assign n41110 = ~pi214 & n40835;
  assign n41111 = n41109 & ~n41110;
  assign n41112 = n40818 & ~n40835;
  assign n41113 = ~pi219 & ~n41112;
  assign n41114 = ~n41111 & n41113;
  assign n41115 = n41106 & ~n41114;
  assign n41116 = pi1150 & n39454;
  assign n41117 = ~n41115 & n41116;
  assign n41118 = ~n41103 & n41117;
  assign n41119 = n40165 & ~n40774;
  assign n41120 = n41098 & ~n41119;
  assign n41121 = ~pi1150 & ~n39407;
  assign n41122 = ~pi211 & n40161;
  assign n41123 = n41115 & ~n41122;
  assign n41124 = n41121 & ~n41123;
  assign n41125 = ~n41120 & n41124;
  assign n41126 = ~pi1149 & ~n41125;
  assign n41127 = ~n41118 & n41126;
  assign n41128 = pi299 & ~n38475;
  assign n41129 = ~n40804 & ~n41128;
  assign n41130 = n6286 & ~n41129;
  assign n41131 = ~n6286 & ~n38475;
  assign n41132 = ~pi57 & pi1147;
  assign n41133 = ~n41131 & n41132;
  assign n41134 = ~n41130 & n41133;
  assign n41135 = pi57 & n38475;
  assign n41136 = n6286 & ~n38474;
  assign n41137 = n40793 & n41136;
  assign n41138 = ~n38475 & ~n40899;
  assign n41139 = ~pi57 & ~pi1147;
  assign n41140 = ~n41131 & n41139;
  assign n41141 = ~n41138 & n41140;
  assign n41142 = ~n41137 & n41141;
  assign n41143 = ~n41135 & ~n41142;
  assign n41144 = ~n41134 & n41143;
  assign n41145 = pi1150 & ~n41144;
  assign n41146 = ~n40865 & n41099;
  assign n41147 = pi212 & ~n41146;
  assign n41148 = n40776 & ~n41100;
  assign n41149 = ~pi219 & ~n41148;
  assign n41150 = ~n41147 & n41149;
  assign n41151 = n41098 & ~n41150;
  assign n41152 = ~n40169 & n40884;
  assign n41153 = ~n41129 & n41152;
  assign n41154 = ~pi1150 & ~n39696;
  assign n41155 = ~n41153 & n41154;
  assign n41156 = ~n41151 & n41155;
  assign n41157 = pi1149 & ~n41156;
  assign n41158 = ~n41145 & n41157;
  assign n41159 = pi1148 & ~n41158;
  assign n41160 = ~n41127 & n41159;
  assign n41161 = pi213 & ~n41160;
  assign n41162 = ~n41096 & n41161;
  assign n41163 = ~pi213 & ~n40861;
  assign n41164 = ~pi209 & ~n41163;
  assign n41165 = ~n41162 & n41164;
  assign n41166 = ~n41049 & ~n41165;
  assign n41167 = pi230 & ~n41166;
  assign n41168 = ~pi230 & ~pi246;
  assign po403 = ~n41167 & ~n41168;
  assign n41170 = ~pi1147 & ~n40252;
  assign n41171 = pi1151 & ~n39664;
  assign n41172 = ~n39635 & n40991;
  assign n41173 = n41171 & ~n41172;
  assign n41174 = n41170 & ~n41173;
  assign n41175 = n39668 & ~n39683;
  assign n41176 = ~n40977 & ~n41175;
  assign n41177 = ~n39696 & ~n41176;
  assign n41178 = ~pi1151 & n41177;
  assign n41179 = pi1151 & ~n39696;
  assign n41180 = ~n40205 & n41179;
  assign n41181 = pi1147 & ~n41180;
  assign n41182 = ~n41178 & n41181;
  assign n41183 = ~pi1149 & ~n41182;
  assign n41184 = ~n41174 & n41183;
  assign n41185 = ~pi1151 & ~n39403;
  assign n41186 = n40937 & ~n41003;
  assign n41187 = n40173 & ~n41186;
  assign n41188 = ~n39739 & n40173;
  assign n41189 = ~n41187 & ~n41188;
  assign n41190 = n41185 & n41189;
  assign n41191 = ~n39876 & n40036;
  assign n41192 = ~pi1147 & ~n41191;
  assign n41193 = ~n41190 & n41192;
  assign n41194 = pi1147 & ~n40265;
  assign n41195 = ~n39653 & ~n39656;
  assign n41196 = n40188 & n41195;
  assign n41197 = n41194 & ~n41196;
  assign n41198 = pi1149 & ~n41197;
  assign n41199 = ~n41193 & n41198;
  assign n41200 = pi1150 & ~n41199;
  assign n41201 = ~n41184 & n41200;
  assign n41202 = pi212 & ~n39252;
  assign n41203 = n40948 & ~n41202;
  assign n41204 = n39721 & ~n41203;
  assign n41205 = n40105 & ~n41204;
  assign n41206 = pi1147 & ~n41205;
  assign n41207 = n38145 & ~n39736;
  assign n41208 = ~n39744 & n40154;
  assign n41209 = ~n41207 & n41208;
  assign n41210 = ~pi1151 & ~n39656;
  assign n41211 = ~n41209 & n41210;
  assign n41212 = ~n39760 & n41211;
  assign n41213 = n41206 & ~n41212;
  assign n41214 = ~n40042 & n40948;
  assign n41215 = n39829 & ~n41214;
  assign n41216 = ~n39403 & ~n41215;
  assign n41217 = pi1151 & n41216;
  assign n41218 = n41185 & ~n41209;
  assign n41219 = ~pi1147 & ~n41218;
  assign n41220 = ~n41217 & n41219;
  assign n41221 = pi1149 & ~n41220;
  assign n41222 = ~n41213 & n41221;
  assign n41223 = ~n40235 & n41179;
  assign n41224 = ~n39694 & n40111;
  assign n41225 = pi1147 & ~n41224;
  assign n41226 = ~n41223 & n41225;
  assign n41227 = ~n39663 & n39727;
  assign n41228 = ~pi1151 & ~n41227;
  assign n41229 = ~pi1147 & ~n41228;
  assign n41230 = ~n39758 & n41171;
  assign n41231 = n41229 & ~n41230;
  assign n41232 = ~pi1149 & ~n41231;
  assign n41233 = ~n41226 & n41232;
  assign n41234 = ~pi1150 & ~n41233;
  assign n41235 = ~n41222 & n41234;
  assign n41236 = ~n41201 & ~n41235;
  assign n41237 = pi1148 & ~n41236;
  assign n41238 = pi1147 & ~n40260;
  assign n41239 = ~pi1151 & n39454;
  assign n41240 = ~n39760 & n41239;
  assign n41241 = n41238 & ~n41240;
  assign n41242 = ~n39716 & n39829;
  assign n41243 = ~n39453 & ~n41242;
  assign n41244 = pi1151 & n41243;
  assign n41245 = ~pi1151 & ~n39453;
  assign n41246 = ~n40138 & n41245;
  assign n41247 = ~pi1147 & ~n41246;
  assign n41248 = ~n41244 & n41247;
  assign n41249 = ~pi1150 & ~n41248;
  assign n41250 = ~n41241 & n41249;
  assign n41251 = ~n41187 & n41245;
  assign n41252 = pi1151 & ~n39453;
  assign n41253 = ~n39879 & n41252;
  assign n41254 = ~pi1147 & ~n41253;
  assign n41255 = ~n41251 & n41254;
  assign n41256 = n39455 & n40167;
  assign n41257 = pi1147 & ~n41256;
  assign n41258 = n39454 & ~n39759;
  assign n41259 = ~pi1151 & n41258;
  assign n41260 = n41257 & ~n41259;
  assign n41261 = pi1150 & ~n41260;
  assign n41262 = ~n41255 & n41261;
  assign n41263 = ~n41250 & ~n41262;
  assign n41264 = pi1149 & ~n41263;
  assign n41265 = n40205 & ~n40212;
  assign n41266 = n39408 & ~n41265;
  assign n41267 = ~n39407 & ~n40983;
  assign n41268 = ~pi1151 & n41267;
  assign n41269 = pi1147 & ~n41268;
  assign n41270 = ~n41266 & n41269;
  assign n41271 = ~pi1151 & ~n39769;
  assign n41272 = ~pi1147 & ~n41271;
  assign n41273 = pi1151 & ~n39634;
  assign n41274 = n41272 & ~n41273;
  assign n41275 = pi1150 & ~n41274;
  assign n41276 = ~n41270 & n41275;
  assign n41277 = ~n39263 & n40165;
  assign n41278 = n40233 & ~n41277;
  assign n41279 = n39408 & ~n41278;
  assign n41280 = n40097 & ~n40166;
  assign n41281 = pi1147 & ~n41280;
  assign n41282 = ~n41279 & n41281;
  assign n41283 = ~pi1147 & pi1151;
  assign n41284 = n39725 & n41283;
  assign n41285 = ~pi1150 & ~n41284;
  assign n41286 = ~n41282 & n41285;
  assign n41287 = ~n41276 & ~n41286;
  assign n41288 = ~pi1149 & ~n41287;
  assign n41289 = ~pi1148 & ~n41288;
  assign n41290 = ~n41264 & n41289;
  assign n41291 = ~n41237 & ~n41290;
  assign n41292 = ~pi213 & ~n41291;
  assign n41293 = pi213 & n40270;
  assign n41294 = pi209 & ~n41293;
  assign n41295 = ~n41292 & n41294;
  assign n41296 = ~n41187 & n41252;
  assign n41297 = pi1147 & ~n40188;
  assign n41298 = ~n41296 & n41297;
  assign n41299 = ~n39456 & ~n40224;
  assign n41300 = n41272 & n41299;
  assign n41301 = ~pi1150 & ~n41300;
  assign n41302 = ~n41298 & n41301;
  assign n41303 = n39680 & n39687;
  assign n41304 = n40036 & ~n41303;
  assign n41305 = n41170 & ~n41304;
  assign n41306 = n40036 & n41189;
  assign n41307 = n40059 & ~n41188;
  assign n41308 = pi1147 & ~n41307;
  assign n41309 = ~n41306 & n41308;
  assign n41310 = pi1150 & ~n41309;
  assign n41311 = ~n41305 & n41310;
  assign n41312 = ~n41302 & ~n41311;
  assign n41313 = ~pi1149 & ~n41312;
  assign n41314 = ~n39654 & n41280;
  assign n41315 = n41257 & ~n41314;
  assign n41316 = ~pi1150 & ~n41315;
  assign n41317 = n40097 & ~n41265;
  assign n41318 = n39454 & ~n40213;
  assign n41319 = ~pi1147 & ~n41318;
  assign n41320 = ~n41317 & n41319;
  assign n41321 = n41316 & ~n41320;
  assign n41322 = n40111 & ~n40205;
  assign n41323 = n41195 & n41273;
  assign n41324 = ~pi1147 & ~n41323;
  assign n41325 = ~n41322 & n41324;
  assign n41326 = ~n39696 & ~n40170;
  assign n41327 = ~pi1151 & n41326;
  assign n41328 = n41194 & ~n41327;
  assign n41329 = pi1150 & ~n41328;
  assign n41330 = ~n41325 & n41329;
  assign n41331 = ~n41321 & ~n41330;
  assign n41332 = pi1149 & ~n41331;
  assign n41333 = pi1148 & ~n41332;
  assign n41334 = ~n41313 & n41333;
  assign n41335 = ~pi219 & ~n39751;
  assign n41336 = ~n40143 & n41335;
  assign n41337 = n39721 & ~n41336;
  assign n41338 = ~n39717 & n41337;
  assign n41339 = n40097 & ~n41338;
  assign n41340 = n41238 & ~n41339;
  assign n41341 = n39299 & n39499;
  assign n41342 = ~n10669 & n41341;
  assign n41343 = ~n41278 & ~n41342;
  assign n41344 = n39455 & n41343;
  assign n41345 = n40097 & ~n41278;
  assign n41346 = ~pi1147 & ~n41345;
  assign n41347 = ~n41344 & n41346;
  assign n41348 = ~pi1150 & ~n41347;
  assign n41349 = ~n41340 & n41348;
  assign n41350 = ~n39696 & ~n41337;
  assign n41351 = ~pi1151 & n41350;
  assign n41352 = n41206 & ~n41351;
  assign n41353 = n40111 & ~n40235;
  assign n41354 = n40105 & ~n41341;
  assign n41355 = ~n40235 & n41354;
  assign n41356 = ~pi1147 & ~n41355;
  assign n41357 = ~n41353 & n41356;
  assign n41358 = pi1150 & ~n41357;
  assign n41359 = ~n41352 & n41358;
  assign n41360 = ~n41349 & ~n41359;
  assign n41361 = pi1149 & ~n41360;
  assign n41362 = n39746 & n40154;
  assign n41363 = ~n39664 & ~n41362;
  assign n41364 = ~pi1151 & n41363;
  assign n41365 = n40036 & ~n41209;
  assign n41366 = pi1147 & ~n41365;
  assign n41367 = ~n41364 & n41366;
  assign n41368 = ~n16361 & n39402;
  assign n41369 = pi1151 & ~n41368;
  assign n41370 = n41229 & ~n41369;
  assign n41371 = pi1150 & ~n41370;
  assign n41372 = ~n41367 & n41371;
  assign n41373 = ~n39453 & ~n40138;
  assign n41374 = ~pi1151 & ~n40928;
  assign n41375 = pi1147 & ~n41374;
  assign n41376 = ~n41373 & n41375;
  assign n41377 = n39728 & n41283;
  assign n41378 = ~pi1150 & ~n41377;
  assign n41379 = ~n41376 & n41378;
  assign n41380 = ~n41372 & ~n41379;
  assign n41381 = ~pi1149 & ~n41380;
  assign n41382 = ~pi1148 & ~n41381;
  assign n41383 = ~n41361 & n41382;
  assign n41384 = ~n41334 & ~n41383;
  assign n41385 = pi213 & ~n41384;
  assign n41386 = ~pi213 & ~n39767;
  assign n41387 = ~pi209 & ~n41386;
  assign n41388 = ~n41385 & n41387;
  assign n41389 = ~n41295 & ~n41388;
  assign n41390 = pi230 & ~n41389;
  assign n41391 = ~pi230 & ~pi247;
  assign po404 = ~n41390 & ~n41391;
  assign n41393 = pi1152 & ~n40265;
  assign n41394 = ~n41204 & n41210;
  assign n41395 = n41393 & ~n41394;
  assign n41396 = pi1151 & ~n39695;
  assign n41397 = n41195 & n41396;
  assign n41398 = ~pi1152 & ~n41397;
  assign n41399 = ~n41212 & n41398;
  assign n41400 = pi1150 & ~n41399;
  assign n41401 = ~n41395 & n41400;
  assign n41402 = pi1151 & n41177;
  assign n41403 = ~pi1152 & ~n41224;
  assign n41404 = ~n41402 & n41403;
  assign n41405 = pi1152 & ~n41353;
  assign n41406 = ~n41180 & n41405;
  assign n41407 = ~pi1150 & ~n41406;
  assign n41408 = ~n41404 & n41407;
  assign n41409 = pi1148 & ~n41408;
  assign n41410 = ~n41401 & n41409;
  assign n41411 = ~n39688 & n41171;
  assign n41412 = ~pi1152 & ~n41411;
  assign n41413 = ~n41228 & n41412;
  assign n41414 = ~n39758 & n40059;
  assign n41415 = pi1152 & ~n41414;
  assign n41416 = ~n41173 & n41415;
  assign n41417 = ~pi1150 & ~n41416;
  assign n41418 = ~n41413 & n41417;
  assign n41419 = ~pi1152 & ~n41218;
  assign n41420 = ~n41306 & n41419;
  assign n41421 = ~pi1151 & n41216;
  assign n41422 = pi1152 & ~n41191;
  assign n41423 = ~n41421 & n41422;
  assign n41424 = pi1150 & ~n41423;
  assign n41425 = ~n41420 & n41424;
  assign n41426 = ~pi1148 & ~n41425;
  assign n41427 = ~n41418 & n41426;
  assign n41428 = ~n41410 & ~n41427;
  assign n41429 = pi1149 & ~n41428;
  assign n41430 = ~n39722 & n41239;
  assign n41431 = pi1152 & ~n41430;
  assign n41432 = ~n41256 & n41431;
  assign n41433 = ~pi1152 & ~n41258;
  assign n41434 = ~n41240 & n41433;
  assign n41435 = ~n41432 & ~n41434;
  assign n41436 = pi1150 & ~n41435;
  assign n41437 = ~n41266 & ~n41345;
  assign n41438 = pi1152 & ~n41437;
  assign n41439 = ~n41267 & ~n41280;
  assign n41440 = ~pi1152 & ~n41439;
  assign n41441 = ~pi1150 & ~n41440;
  assign n41442 = ~n41438 & n41441;
  assign n41443 = pi1148 & ~n41442;
  assign n41444 = ~n41436 & n41443;
  assign n41445 = ~pi1151 & n41243;
  assign n41446 = pi1152 & ~n41253;
  assign n41447 = ~n41445 & n41446;
  assign n41448 = ~pi1152 & ~n41246;
  assign n41449 = ~n41296 & n41448;
  assign n41450 = pi1150 & ~n41449;
  assign n41451 = ~n41447 & n41450;
  assign n41452 = ~pi1151 & ~n39725;
  assign n41453 = pi1152 & ~n41273;
  assign n41454 = ~n41452 & n41453;
  assign n41455 = pi1151 & ~pi1152;
  assign n41456 = n39769 & n41455;
  assign n41457 = ~pi1150 & ~n41456;
  assign n41458 = ~n41454 & n41457;
  assign n41459 = ~n41451 & ~n41458;
  assign n41460 = ~pi1148 & ~n41459;
  assign n41461 = ~pi1149 & ~n41460;
  assign n41462 = ~n41444 & n41461;
  assign n41463 = ~n41429 & ~n41462;
  assign n41464 = ~pi213 & ~n41463;
  assign n41465 = ~n39689 & n41455;
  assign n41466 = ~pi1151 & ~n39728;
  assign n41467 = ~n39725 & n41466;
  assign n41468 = pi1152 & ~n41467;
  assign n41469 = ~n40253 & n41468;
  assign n41470 = ~pi1150 & ~n41469;
  assign n41471 = ~n41465 & n41470;
  assign n41472 = n41393 & ~n41430;
  assign n41473 = pi1151 & n39698;
  assign n41474 = ~pi1152 & ~n41473;
  assign n41475 = ~n40261 & n41474;
  assign n41476 = pi1150 & ~n41475;
  assign n41477 = ~n41472 & n41476;
  assign n41478 = ~n41471 & ~n41477;
  assign n41479 = pi213 & n41478;
  assign n41480 = pi209 & ~n41479;
  assign n41481 = ~n41464 & n41480;
  assign n41482 = pi1151 & n41350;
  assign n41483 = ~pi1152 & ~n41339;
  assign n41484 = ~n41482 & n41483;
  assign n41485 = ~n41205 & n41431;
  assign n41486 = pi1150 & ~n41485;
  assign n41487 = ~n41484 & n41486;
  assign n41488 = pi1152 & ~n41246;
  assign n41489 = ~n41365 & n41488;
  assign n41490 = ~pi1150 & ~n41489;
  assign n41491 = ~pi1152 & ~n41374;
  assign n41492 = ~n41363 & n41491;
  assign n41493 = n41490 & ~n41492;
  assign n41494 = ~pi1149 & ~n41493;
  assign n41495 = ~n41487 & n41494;
  assign n41496 = pi1152 & ~n41251;
  assign n41497 = ~n41306 & n41496;
  assign n41498 = n41171 & ~n41188;
  assign n41499 = n40189 & ~n41498;
  assign n41500 = ~pi1150 & ~n41499;
  assign n41501 = ~n41497 & n41500;
  assign n41502 = n40167 & n41239;
  assign n41503 = n41393 & ~n41502;
  assign n41504 = pi1151 & n41326;
  assign n41505 = ~pi1152 & ~n41314;
  assign n41506 = ~n41504 & n41505;
  assign n41507 = pi1150 & ~n41506;
  assign n41508 = ~n41503 & n41507;
  assign n41509 = pi1149 & ~n41508;
  assign n41510 = ~n41501 & n41509;
  assign n41511 = pi1148 & ~n41510;
  assign n41512 = ~n41495 & n41511;
  assign n41513 = ~n41271 & n41412;
  assign n41514 = ~pi1151 & ~n41299;
  assign n41515 = pi1152 & ~n41514;
  assign n41516 = ~n41304 & n41515;
  assign n41517 = ~pi1150 & ~n41516;
  assign n41518 = ~n41513 & n41517;
  assign n41519 = ~pi1152 & ~n41180;
  assign n41520 = ~n41317 & n41519;
  assign n41521 = ~pi1151 & n41318;
  assign n41522 = pi1152 & ~n41323;
  assign n41523 = ~n41521 & n41522;
  assign n41524 = pi1150 & ~n41523;
  assign n41525 = ~n41520 & n41524;
  assign n41526 = pi1149 & ~n41525;
  assign n41527 = ~n41518 & n41526;
  assign n41528 = n41239 & n41343;
  assign n41529 = pi1152 & ~n41355;
  assign n41530 = ~n41528 & n41529;
  assign n41531 = ~pi1152 & ~n41345;
  assign n41532 = ~n41223 & n41531;
  assign n41533 = pi1150 & ~n41532;
  assign n41534 = ~n41530 & n41533;
  assign n41535 = pi1152 & ~n41369;
  assign n41536 = ~n41466 & n41535;
  assign n41537 = n41227 & n41455;
  assign n41538 = ~pi1150 & ~n41537;
  assign n41539 = ~n41536 & n41538;
  assign n41540 = ~pi1149 & ~n41539;
  assign n41541 = ~n41534 & n41540;
  assign n41542 = ~pi1148 & ~n41541;
  assign n41543 = ~n41527 & n41542;
  assign n41544 = pi213 & ~n41543;
  assign n41545 = ~n41512 & n41544;
  assign n41546 = ~pi213 & ~n41046;
  assign n41547 = ~pi209 & ~n41546;
  assign n41548 = ~n41545 & n41547;
  assign n41549 = ~n41481 & ~n41548;
  assign n41550 = pi230 & ~n41549;
  assign n41551 = ~pi230 & ~pi248;
  assign po405 = ~n41550 & ~n41551;
  assign n41553 = ~pi213 & n41478;
  assign n41554 = pi299 & n38505;
  assign n41555 = ~n39744 & ~n41554;
  assign n41556 = ~n39267 & n41555;
  assign n41557 = ~pi212 & ~n41556;
  assign n41558 = ~pi214 & n41555;
  assign n41559 = pi214 & ~n39735;
  assign n41560 = n39253 & n41559;
  assign n41561 = pi212 & ~n41560;
  assign n41562 = ~n41558 & n41561;
  assign n41563 = ~n41557 & ~n41562;
  assign n41564 = ~pi219 & ~n41563;
  assign n41565 = n6286 & ~n40153;
  assign n41566 = ~n41564 & n41565;
  assign n41567 = ~n6286 & n38564;
  assign n41568 = ~pi57 & ~pi1151;
  assign n41569 = ~n41567 & n41568;
  assign n41570 = ~n41566 & n41569;
  assign n41571 = pi57 & ~n38564;
  assign n41572 = ~n40174 & ~n41554;
  assign n41573 = ~pi214 & ~n41572;
  assign n41574 = ~n39329 & n39518;
  assign n41575 = pi212 & ~n41574;
  assign n41576 = ~n41573 & n41575;
  assign n41577 = ~pi219 & ~n41576;
  assign n41578 = n39269 & n41572;
  assign n41579 = n41577 & ~n41578;
  assign n41580 = n6286 & ~n39352;
  assign n41581 = ~n41579 & n41580;
  assign n41582 = ~pi57 & pi1151;
  assign n41583 = ~n41567 & n41582;
  assign n41584 = ~n41581 & n41583;
  assign n41585 = ~n41571 & ~n41584;
  assign n41586 = ~n41570 & n41585;
  assign n41587 = ~pi1152 & ~n41586;
  assign n41588 = n39706 & ~n40132;
  assign n41589 = ~n39265 & n41573;
  assign n41590 = n40041 & ~n41589;
  assign n41591 = ~n41588 & n41590;
  assign n41592 = n39754 & ~n41554;
  assign n41593 = n40947 & ~n41592;
  assign n41594 = ~n41591 & n41593;
  assign n41595 = ~pi1151 & ~n41594;
  assign n41596 = n39721 & n41595;
  assign n41597 = pi299 & ~n38505;
  assign n41598 = ~n10669 & n41597;
  assign n41599 = ~n38503 & ~n41598;
  assign n41600 = n39651 & ~n41599;
  assign n41601 = n40161 & ~n41600;
  assign n41602 = ~n39866 & ~n40092;
  assign n41603 = pi1151 & ~n41602;
  assign n41604 = ~n41601 & n41603;
  assign n41605 = n38510 & ~n41604;
  assign n41606 = ~n41596 & n41605;
  assign n41607 = pi1150 & ~n41606;
  assign n41608 = ~n41587 & n41607;
  assign n41609 = ~n38357 & ~n39669;
  assign n41610 = pi211 & n41609;
  assign n41611 = ~n38388 & n39674;
  assign n41612 = n38468 & ~n41611;
  assign n41613 = ~n41610 & n41612;
  assign n41614 = ~n38357 & n39680;
  assign n41615 = ~n38468 & ~n41614;
  assign n41616 = ~n41613 & ~n41615;
  assign n41617 = ~pi219 & ~n41616;
  assign n41618 = pi1151 & n39687;
  assign n41619 = ~n41617 & n41618;
  assign n41620 = ~n39329 & ~n41598;
  assign n41621 = n38563 & n39295;
  assign n41622 = ~n41620 & n41621;
  assign n41623 = n38566 & ~n41622;
  assign n41624 = ~n41619 & n41623;
  assign n41625 = ~n11321 & n38347;
  assign n41626 = ~n39317 & ~n41625;
  assign n41627 = ~pi211 & ~n38357;
  assign n41628 = ~n41626 & n41627;
  assign n41629 = ~n40112 & ~n41628;
  assign n41630 = pi214 & n41629;
  assign n41631 = n39636 & ~n41597;
  assign n41632 = pi212 & ~n41631;
  assign n41633 = ~n41630 & n41632;
  assign n41634 = n39858 & ~n41592;
  assign n41635 = ~n41633 & n41634;
  assign n41636 = n39273 & ~n39850;
  assign n41637 = ~n41635 & n41636;
  assign n41638 = ~pi1151 & n41278;
  assign n41639 = n38510 & ~n41622;
  assign n41640 = ~n41638 & n41639;
  assign n41641 = ~n41637 & n41640;
  assign n41642 = ~pi1150 & ~n41641;
  assign n41643 = ~n41624 & n41642;
  assign n41644 = ~n41608 & ~n41643;
  assign n41645 = pi213 & ~n41644;
  assign n41646 = ~pi209 & ~n41645;
  assign n41647 = ~n41553 & n41646;
  assign n41648 = ~n38704 & ~n39665;
  assign n41649 = ~pi212 & ~n41648;
  assign n41650 = ~pi219 & ~n41649;
  assign n41651 = pi212 & ~n40201;
  assign n41652 = ~n38692 & n41651;
  assign n41653 = n41650 & ~n41652;
  assign n41654 = n40991 & ~n41653;
  assign n41655 = n38706 & n41654;
  assign n41656 = n41171 & ~n41655;
  assign n41657 = n38704 & n38714;
  assign n41658 = ~n41455 & ~n41657;
  assign n41659 = ~n41656 & ~n41658;
  assign n41660 = pi214 & n38618;
  assign n41661 = n38641 & ~n41660;
  assign n41662 = ~pi219 & ~n41661;
  assign n41663 = pi214 & ~n38633;
  assign n41664 = ~pi214 & n38618;
  assign n41665 = pi212 & ~n41664;
  assign n41666 = ~n41663 & n41665;
  assign n41667 = n41662 & ~n41666;
  assign n41668 = ~po1038 & ~n38636;
  assign n41669 = ~n41667 & n41668;
  assign n41670 = n40036 & ~n41669;
  assign n41671 = ~n38633 & n39463;
  assign n41672 = ~n38631 & ~n39463;
  assign n41673 = ~po1038 & ~n41672;
  assign n41674 = ~n41671 & n41673;
  assign n41675 = n41245 & ~n41674;
  assign n41676 = pi1152 & ~n41675;
  assign n41677 = ~n41670 & n41676;
  assign n41678 = ~n41659 & ~n41677;
  assign n41679 = ~pi1150 & ~n41678;
  assign n41680 = n38705 & ~n41128;
  assign n41681 = ~po1038 & ~n41680;
  assign n41682 = ~n41653 & n41681;
  assign n41683 = n41179 & ~n41682;
  assign n41684 = ~n38704 & n40165;
  assign n41685 = n41681 & ~n41684;
  assign n41686 = n40097 & ~n41685;
  assign n41687 = ~pi1152 & ~n41686;
  assign n41688 = ~n41683 & n41687;
  assign n41689 = ~n38640 & ~n41663;
  assign n41690 = ~pi212 & ~n41689;
  assign n41691 = ~pi214 & n38633;
  assign n41692 = ~pi211 & n38631;
  assign n41693 = ~n38663 & ~n41692;
  assign n41694 = pi214 & ~n41693;
  assign n41695 = pi212 & ~n41694;
  assign n41696 = ~n41691 & n41695;
  assign n41697 = ~n41690 & ~n41696;
  assign n41698 = ~pi219 & ~n41697;
  assign n41699 = n38639 & ~n41698;
  assign n41700 = n41239 & ~n41699;
  assign n41701 = pi212 & ~n38618;
  assign n41702 = n41662 & ~n41701;
  assign n41703 = n38639 & ~n41702;
  assign n41704 = n40105 & ~n41703;
  assign n41705 = pi1152 & ~n41704;
  assign n41706 = ~n41700 & n41705;
  assign n41707 = ~n41688 & ~n41706;
  assign n41708 = pi1150 & ~n41707;
  assign n41709 = ~n41679 & ~n41708;
  assign n41710 = ~pi213 & ~n41709;
  assign n41711 = pi213 & n38712;
  assign n41712 = pi209 & ~n41711;
  assign n41713 = ~n41710 & n41712;
  assign n41714 = ~n41647 & ~n41713;
  assign n41715 = pi230 & ~n41714;
  assign n41716 = ~pi230 & ~pi249;
  assign po406 = ~n41715 & ~n41716;
  assign n41718 = n3276 & n11448;
  assign n41719 = ~n6236 & ~n41718;
  assign n41720 = ~pi75 & ~n41719;
  assign n41721 = n7300 & n8925;
  assign n41722 = ~n41720 & ~n41721;
  assign n41723 = ~pi87 & ~pi250;
  assign n41724 = n8841 & n41723;
  assign po407 = ~n41722 & n41724;
  assign n41726 = pi897 & n10758;
  assign n41727 = ~pi476 & n11381;
  assign n41728 = ~n41726 & ~n41727;
  assign n41729 = pi200 & pi1039;
  assign n41730 = ~pi200 & pi1053;
  assign n41731 = ~pi199 & ~n41730;
  assign n41732 = ~n41729 & n41731;
  assign n41733 = ~n41728 & ~n41732;
  assign n41734 = pi251 & n41728;
  assign po408 = n41733 | n41734;
  assign n41736 = ~pi979 & ~pi984;
  assign n41737 = pi1001 & n41736;
  assign n41738 = n6168 & n41737;
  assign n41739 = ~n6171 & n41738;
  assign n41740 = n6435 & n41739;
  assign n41741 = ~pi252 & ~n41740;
  assign n41742 = pi1092 & ~pi1093;
  assign n41743 = ~n41741 & n41742;
  assign n41744 = n6447 & ~n41743;
  assign n41745 = n6446 & n41743;
  assign n41746 = ~n41744 & ~n41745;
  assign n41747 = ~n6192 & n41746;
  assign n41748 = n6192 & n11488;
  assign n41749 = ~n41747 & ~n41748;
  assign n41750 = ~n6215 & ~n41749;
  assign n41751 = ~n6198 & n11488;
  assign n41752 = n6198 & n41746;
  assign n41753 = ~n41751 & ~n41752;
  assign n41754 = n6215 & ~n41753;
  assign n41755 = ~pi299 & ~n41754;
  assign n41756 = ~n41750 & n41755;
  assign n41757 = ~n6189 & ~n41749;
  assign n41758 = n6189 & ~n41753;
  assign n41759 = pi299 & ~n41758;
  assign n41760 = ~n41757 & n41759;
  assign n41761 = n10923 & ~n41760;
  assign n41762 = ~n41756 & n41761;
  assign n41763 = ~n10923 & n11488;
  assign n41764 = ~n8830 & ~n41763;
  assign n41765 = ~n41762 & n41764;
  assign n41766 = n10922 & n41738;
  assign n41767 = n20983 & n41766;
  assign n41768 = n6175 & n41767;
  assign n41769 = ~n38109 & n41768;
  assign n41770 = n6435 & n41769;
  assign n41771 = ~pi252 & ~n41770;
  assign n41772 = ~pi57 & pi1092;
  assign n41773 = ~n41771 & n41772;
  assign n41774 = pi57 & n11487;
  assign n41775 = n8830 & ~n41774;
  assign n41776 = ~n41773 & n41775;
  assign po409 = ~n41765 & ~n41776;
  assign n41778 = ~n12978 & ~n38230;
  assign n41779 = ~n38329 & n41778;
  assign n41780 = ~po1038 & n41779;
  assign n41781 = ~pi211 & po1038;
  assign n41782 = pi219 & n41781;
  assign n41783 = ~n41780 & ~n41782;
  assign n41784 = pi1153 & ~n41783;
  assign n41785 = ~pi1151 & ~n41784;
  assign n41786 = pi1153 & ~n38278;
  assign n41787 = ~n38650 & ~n41786;
  assign n41788 = n10670 & n41787;
  assign n41789 = pi211 & ~n38272;
  assign n41790 = ~n41788 & ~n41789;
  assign n41791 = ~n38265 & ~n38278;
  assign n41792 = n38241 & ~n41791;
  assign n41793 = ~po1038 & ~n41792;
  assign n41794 = n41790 & n41793;
  assign n41795 = ~n11383 & n38972;
  assign n41796 = pi1151 & ~n41795;
  assign n41797 = ~n41794 & n41796;
  assign n41798 = ~n41785 & ~n41797;
  assign n41799 = ~pi1152 & ~n41798;
  assign n41800 = n38241 & n39360;
  assign n41801 = ~pi1151 & ~n11384;
  assign n41802 = ~n38309 & n41801;
  assign n41803 = ~n41800 & n41802;
  assign n41804 = ~n38270 & ~n39482;
  assign n41805 = pi1153 & ~n41804;
  assign n41806 = ~n11311 & ~n38230;
  assign n41807 = pi1151 & n41806;
  assign n41808 = ~n41805 & n41807;
  assign n41809 = ~po1038 & ~n41808;
  assign n41810 = ~n41803 & n41809;
  assign n41811 = ~pi1151 & n10670;
  assign n41812 = n38972 & ~n41811;
  assign n41813 = pi1152 & ~n41812;
  assign n41814 = ~n41810 & n41813;
  assign n41815 = ~n41799 & ~n41814;
  assign n41816 = pi230 & ~n41815;
  assign n41817 = ~n40391 & ~n40405;
  assign n41818 = ~pi211 & n40385;
  assign n41819 = n41817 & ~n41818;
  assign n41820 = ~n40384 & n40425;
  assign n41821 = n41819 & n41820;
  assign n41822 = pi1153 & ~n41821;
  assign n41823 = ~pi1153 & ~n40531;
  assign n41824 = pi219 & ~n41823;
  assign n41825 = ~n41822 & n41824;
  assign n41826 = ~n40385 & n40414;
  assign n41827 = ~n40425 & ~n41826;
  assign n41828 = ~pi1153 & n41827;
  assign n41829 = ~n40414 & ~n41828;
  assign n41830 = ~pi219 & n40446;
  assign n41831 = ~n41829 & n41830;
  assign n41832 = pi253 & ~n41831;
  assign n41833 = ~n41825 & n41832;
  assign n41834 = ~n40396 & n40531;
  assign n41835 = ~pi211 & n41834;
  assign n41836 = ~n40398 & ~n41835;
  assign n41837 = pi1153 & ~n41836;
  assign n41838 = ~n40526 & ~n41837;
  assign n41839 = pi219 & n41838;
  assign n41840 = pi1153 & n40401;
  assign n41841 = ~pi219 & ~n40444;
  assign n41842 = ~n41840 & n41841;
  assign n41843 = ~pi253 & ~n41842;
  assign n41844 = ~n41839 & n41843;
  assign n41845 = ~n41833 & ~n41844;
  assign n41846 = ~po1038 & ~n41845;
  assign n41847 = pi219 & pi1091;
  assign n41848 = ~n38222 & n41847;
  assign n41849 = ~pi219 & ~n40376;
  assign n41850 = ~n41848 & ~n41849;
  assign n41851 = ~pi211 & ~n40367;
  assign n41852 = pi219 & ~n40394;
  assign n41853 = ~n41851 & n41852;
  assign n41854 = n41850 & ~n41853;
  assign n41855 = ~pi253 & ~n41854;
  assign n41856 = ~pi219 & ~n40378;
  assign n41857 = ~n40394 & ~n41848;
  assign n41858 = ~n41856 & n41857;
  assign n41859 = pi253 & ~n41858;
  assign n41860 = po1038 & ~n41859;
  assign n41861 = ~n41855 & n41860;
  assign n41862 = ~pi211 & ~n40376;
  assign n41863 = n41856 & ~n41862;
  assign n41864 = ~pi219 & ~n41863;
  assign n41865 = po1038 & n41864;
  assign n41866 = ~n40367 & n41865;
  assign n41867 = pi1151 & ~n41866;
  assign n41868 = ~n41861 & n41867;
  assign n41869 = ~n41846 & n41868;
  assign n41870 = ~n40397 & n41819;
  assign n41871 = ~n41828 & n41870;
  assign n41872 = pi219 & ~n40383;
  assign n41873 = ~n41871 & ~n41872;
  assign n41874 = ~n41839 & ~n41873;
  assign n41875 = ~pi253 & ~n41874;
  assign n41876 = ~n40386 & ~n41835;
  assign n41877 = n41856 & ~n41876;
  assign n41878 = ~n41829 & n41877;
  assign n41879 = pi219 & n40486;
  assign n41880 = ~n40498 & n41822;
  assign n41881 = n41879 & ~n41880;
  assign n41882 = ~n41878 & ~n41881;
  assign n41883 = pi253 & ~n41882;
  assign n41884 = ~po1038 & ~n41883;
  assign n41885 = ~n41875 & n41884;
  assign n41886 = ~pi1151 & ~n41885;
  assign n41887 = ~n41869 & ~n41886;
  assign n41888 = n41849 & ~n41851;
  assign n41889 = n41856 & ~n41888;
  assign n41890 = pi219 & ~n40367;
  assign n41891 = po1038 & ~n41890;
  assign n41892 = ~n41889 & n41891;
  assign n41893 = ~n40367 & n41892;
  assign n41894 = ~n41861 & ~n41893;
  assign n41895 = ~n41887 & n41894;
  assign n41896 = pi1152 & ~n41895;
  assign n41897 = pi219 & ~n41838;
  assign n41898 = ~n41842 & n41877;
  assign n41899 = ~n41897 & ~n41898;
  assign n41900 = ~n40396 & ~n41899;
  assign n41901 = ~pi253 & ~n41900;
  assign n41902 = pi1153 & ~n40436;
  assign n41903 = n41819 & n41856;
  assign n41904 = ~n41902 & n41903;
  assign n41905 = ~n40488 & ~n41821;
  assign n41906 = pi1153 & n41905;
  assign n41907 = ~pi1153 & ~n40537;
  assign n41908 = pi219 & ~n41907;
  assign n41909 = ~n41906 & n41908;
  assign n41910 = ~n41904 & ~n41909;
  assign n41911 = pi253 & ~n41910;
  assign n41912 = ~po1038 & ~n41911;
  assign n41913 = ~n41901 & n41912;
  assign n41914 = n41868 & ~n41913;
  assign n41915 = ~n40383 & n41897;
  assign n41916 = ~pi1153 & ~n40428;
  assign n41917 = ~n40396 & ~n41916;
  assign n41918 = n41830 & n41917;
  assign n41919 = ~pi253 & ~n41918;
  assign n41920 = ~n41915 & n41919;
  assign n41921 = ~n40498 & ~n41821;
  assign n41922 = ~pi1091 & ~n40526;
  assign n41923 = ~pi1153 & ~n41922;
  assign n41924 = ~pi219 & ~n41827;
  assign n41925 = ~n41923 & ~n41924;
  assign n41926 = n41921 & n41925;
  assign n41927 = pi253 & ~n41926;
  assign n41928 = ~po1038 & ~n41927;
  assign n41929 = ~n41920 & n41928;
  assign n41930 = ~pi1151 & ~n41861;
  assign n41931 = ~n41929 & n41930;
  assign n41932 = ~pi1152 & ~n41931;
  assign n41933 = ~n41914 & n41932;
  assign n41934 = ~n41896 & ~n41933;
  assign n41935 = n40648 & ~n41934;
  assign n41936 = pi1091 & ~n41790;
  assign n41937 = pi1091 & n38241;
  assign n41938 = ~n38621 & ~n40588;
  assign n41939 = n41937 & ~n41938;
  assign n41940 = ~n41936 & ~n41939;
  assign n41941 = pi253 & ~n41940;
  assign n41942 = ~n12981 & ~n41805;
  assign n41943 = pi1091 & ~n41942;
  assign n41944 = ~pi253 & ~n41943;
  assign n41945 = ~po1038 & ~n41944;
  assign n41946 = ~n41941 & n41945;
  assign n41947 = ~pi253 & ~pi1091;
  assign n41948 = po1038 & ~n41947;
  assign n41949 = pi211 & pi1091;
  assign n41950 = pi1091 & ~pi1153;
  assign n41951 = pi219 & n41950;
  assign n41952 = ~n41949 & ~n41951;
  assign n41953 = n41948 & n41952;
  assign n41954 = pi1151 & ~n41953;
  assign n41955 = ~n41946 & n41954;
  assign n41956 = ~n41848 & n41948;
  assign n41957 = pi219 & n41956;
  assign n41958 = pi1091 & pi1153;
  assign n41959 = n41780 & n41958;
  assign n41960 = pi253 & ~pi1091;
  assign n41961 = ~pi1151 & ~n41960;
  assign n41962 = ~n41959 & n41961;
  assign n41963 = ~n41957 & n41962;
  assign n41964 = ~n41955 & ~n41963;
  assign n41965 = ~pi1152 & ~n41964;
  assign n41966 = n11383 & n40556;
  assign n41967 = ~n38309 & n41966;
  assign n41968 = pi253 & ~n41967;
  assign n41969 = ~n38255 & n40556;
  assign n41970 = pi1153 & ~n41969;
  assign n41971 = n38241 & ~n41970;
  assign n41972 = n40593 & n41971;
  assign n41973 = n41968 & ~n41972;
  assign n41974 = pi1091 & n38309;
  assign n41975 = pi211 & ~n40607;
  assign n41976 = ~n41974 & n41975;
  assign n41977 = pi1091 & n39360;
  assign n41978 = pi1091 & n38278;
  assign n41979 = n38623 & n41978;
  assign n41980 = n38241 & ~n41979;
  assign n41981 = ~n41977 & n41980;
  assign n41982 = ~pi253 & ~n41981;
  assign n41983 = ~n41976 & n41982;
  assign n41984 = ~n41973 & ~n41983;
  assign n41985 = ~n11383 & ~n38241;
  assign n41986 = ~n41960 & n41985;
  assign n41987 = ~n41974 & n41986;
  assign n41988 = n39295 & ~n41987;
  assign n41989 = ~n41984 & n41988;
  assign n41990 = n41804 & ~n41960;
  assign n41991 = ~n41950 & ~n41990;
  assign n41992 = n41806 & ~n41991;
  assign n41993 = ~po1038 & ~n41947;
  assign n41994 = ~n41992 & n41993;
  assign n41995 = ~n41956 & ~n41994;
  assign n41996 = pi1151 & ~n41995;
  assign n41997 = ~pi211 & pi1091;
  assign n41998 = ~pi219 & n41997;
  assign n41999 = n41956 & ~n41998;
  assign n42000 = pi1152 & ~n41999;
  assign n42001 = ~n41996 & n42000;
  assign n42002 = ~n41989 & n42001;
  assign n42003 = ~n40648 & ~n42002;
  assign n42004 = ~n41965 & n42003;
  assign n42005 = ~pi230 & ~n42004;
  assign n42006 = ~n41935 & n42005;
  assign po410 = ~n41816 & ~n42006;
  assign n42008 = pi1154 & n38645;
  assign n42009 = ~n38674 & ~n42008;
  assign n42010 = n11383 & ~n42009;
  assign n42011 = pi299 & n38241;
  assign n42012 = ~n11383 & n38624;
  assign n42013 = ~n42011 & ~n42012;
  assign n42014 = ~n38847 & ~n42013;
  assign n42015 = ~n42010 & ~n42014;
  assign n42016 = ~po1038 & ~n42015;
  assign n42017 = ~pi219 & ~n38504;
  assign n42018 = ~n38773 & ~n42017;
  assign n42019 = po1038 & n42018;
  assign n42020 = ~pi1152 & ~n42019;
  assign n42021 = ~n42016 & n42020;
  assign n42022 = ~n38262 & ~n38644;
  assign n42023 = n38205 & ~n42022;
  assign n42024 = n38607 & ~n38849;
  assign n42025 = ~n42023 & ~n42024;
  assign n42026 = pi219 & ~n42025;
  assign n42027 = ~pi200 & pi1154;
  assign n42028 = n11321 & ~n42027;
  assign n42029 = n38644 & ~n39482;
  assign n42030 = ~n42028 & ~n42029;
  assign n42031 = ~pi219 & ~n42030;
  assign n42032 = ~po1038 & ~n42031;
  assign n42033 = ~n42026 & n42032;
  assign n42034 = n11383 & ~n38504;
  assign n42035 = n39625 & ~n42034;
  assign n42036 = pi1152 & ~n42035;
  assign n42037 = ~n42033 & n42036;
  assign n42038 = ~n42021 & ~n42037;
  assign n42039 = pi230 & ~n42038;
  assign n42040 = ~pi1153 & n40425;
  assign n42041 = n41876 & ~n42040;
  assign n42042 = n41819 & ~n42041;
  assign n42043 = ~pi1154 & n42042;
  assign n42044 = n40386 & n40436;
  assign n42045 = pi1153 & ~n42044;
  assign n42046 = pi1154 & ~n40390;
  assign n42047 = n41819 & n42046;
  assign n42048 = ~n42045 & n42047;
  assign n42049 = pi254 & ~n42048;
  assign n42050 = ~n42043 & n42049;
  assign n42051 = ~n40397 & n40537;
  assign n42052 = pi1154 & n42051;
  assign n42053 = ~n40444 & ~n42052;
  assign n42054 = ~n40431 & ~n41818;
  assign n42055 = ~pi1153 & n42054;
  assign n42056 = ~pi254 & ~n42055;
  assign n42057 = ~n42053 & n42056;
  assign n42058 = ~n42050 & ~n42057;
  assign n42059 = ~pi219 & ~n42058;
  assign n42060 = pi1154 & ~n41822;
  assign n42061 = ~n41905 & n42060;
  assign n42062 = pi1153 & ~n40531;
  assign n42063 = ~pi1154 & ~n41907;
  assign n42064 = ~n42062 & n42063;
  assign n42065 = pi254 & ~n42064;
  assign n42066 = ~n42061 & n42065;
  assign n42067 = ~pi1153 & ~n40542;
  assign n42068 = n40528 & ~n42067;
  assign n42069 = ~pi1154 & ~n42068;
  assign n42070 = ~n40396 & n40526;
  assign n42071 = n42069 & ~n42070;
  assign n42072 = ~n41823 & n42051;
  assign n42073 = n38220 & ~n42072;
  assign n42074 = ~n40368 & n42073;
  assign n42075 = pi1153 & n40398;
  assign n42076 = n38205 & ~n40515;
  assign n42077 = ~n42075 & n42076;
  assign n42078 = ~pi254 & ~n42077;
  assign n42079 = ~n42074 & n42078;
  assign n42080 = ~n42071 & n42079;
  assign n42081 = ~n42066 & ~n42080;
  assign n42082 = pi219 & ~n42081;
  assign n42083 = pi253 & ~n42082;
  assign n42084 = ~n42059 & n42083;
  assign n42085 = ~pi211 & n38650;
  assign n42086 = ~pi1153 & ~n40561;
  assign n42087 = pi1153 & ~n40574;
  assign n42088 = ~pi1154 & ~n42087;
  assign n42089 = ~n42086 & n42088;
  assign n42090 = ~n42085 & n42089;
  assign n42091 = pi1153 & ~n11321;
  assign n42092 = pi1091 & n38205;
  assign n42093 = ~n38270 & n42092;
  assign n42094 = ~n42091 & n42093;
  assign n42095 = ~n42090 & ~n42094;
  assign n42096 = ~pi219 & ~n42095;
  assign n42097 = pi1154 & n41997;
  assign n42098 = ~n41847 & ~n42097;
  assign n42099 = ~n42025 & ~n42098;
  assign n42100 = ~n42096 & ~n42099;
  assign n42101 = pi254 & ~n42100;
  assign n42102 = ~pi254 & ~pi1091;
  assign n42103 = pi1154 & ~n41804;
  assign n42104 = pi219 & ~n38849;
  assign n42105 = ~n42103 & n42104;
  assign n42106 = ~n42031 & ~n42105;
  assign n42107 = ~pi254 & ~n42106;
  assign n42108 = ~n42102 & ~n42107;
  assign n42109 = ~n42101 & n42108;
  assign n42110 = ~pi253 & ~n42109;
  assign n42111 = ~po1038 & ~n42110;
  assign n42112 = ~n42084 & n42111;
  assign n42113 = n41888 & ~n41958;
  assign n42114 = pi1091 & n38773;
  assign n42115 = ~pi254 & ~n42114;
  assign n42116 = ~n41853 & n42115;
  assign n42117 = ~n42113 & n42116;
  assign n42118 = ~pi211 & ~n40392;
  assign n42119 = n41890 & ~n42118;
  assign n42120 = ~pi219 & n40376;
  assign n42121 = ~n42119 & ~n42120;
  assign n42122 = n11383 & n41950;
  assign n42123 = pi254 & ~n42122;
  assign n42124 = ~n42114 & n42123;
  assign n42125 = n42121 & n42124;
  assign n42126 = pi253 & ~n42125;
  assign n42127 = ~n42117 & n42126;
  assign n42128 = pi1091 & ~n42018;
  assign n42129 = po1038 & ~n42102;
  assign n42130 = ~n42128 & n42129;
  assign n42131 = po1038 & n41998;
  assign n42132 = ~n42130 & ~n42131;
  assign n42133 = pi253 & po1038;
  assign n42134 = n42132 & ~n42133;
  assign n42135 = ~n42127 & ~n42134;
  assign n42136 = pi1152 & ~n42135;
  assign n42137 = ~n42112 & n42136;
  assign n42138 = ~pi1154 & ~n40519;
  assign n42139 = ~pi1154 & ~n42138;
  assign n42140 = ~n41820 & ~n42040;
  assign n42141 = ~n42139 & n42140;
  assign n42142 = n38220 & ~n40498;
  assign n42143 = pi219 & ~n42142;
  assign n42144 = ~n42141 & n42143;
  assign n42145 = pi1154 & n40413;
  assign n42146 = ~pi219 & ~n42145;
  assign n42147 = ~n42041 & n42146;
  assign n42148 = ~n42144 & ~n42147;
  assign n42149 = pi254 & ~n42148;
  assign n42150 = n40399 & ~n41823;
  assign n42151 = n38205 & ~n42150;
  assign n42152 = pi219 & ~n42073;
  assign n42153 = ~n42069 & n42152;
  assign n42154 = ~n42151 & n42153;
  assign n42155 = ~n40390 & n40444;
  assign n42156 = ~n41916 & n42155;
  assign n42157 = ~n40396 & n40446;
  assign n42158 = pi1154 & ~n42157;
  assign n42159 = ~n42156 & n42158;
  assign n42160 = ~pi1154 & ~n42156;
  assign n42161 = pi1154 & n40391;
  assign n42162 = ~n40385 & ~n42161;
  assign n42163 = ~pi211 & ~n42162;
  assign n42164 = ~pi219 & ~n42163;
  assign n42165 = ~n42160 & n42164;
  assign n42166 = ~n42159 & n42165;
  assign n42167 = ~pi254 & ~n42166;
  assign n42168 = ~n42154 & n42167;
  assign n42169 = ~n42149 & ~n42168;
  assign n42170 = pi253 & ~n42169;
  assign n42171 = n40564 & n41950;
  assign n42172 = ~n41977 & ~n42171;
  assign n42173 = pi211 & ~n42088;
  assign n42174 = ~n42172 & n42173;
  assign n42175 = pi1091 & n38624;
  assign n42176 = pi1154 & ~n42175;
  assign n42177 = n11382 & n41958;
  assign n42178 = ~pi1154 & ~n42177;
  assign n42179 = ~pi211 & ~n42178;
  assign n42180 = ~n42176 & n42179;
  assign n42181 = ~n42174 & ~n42180;
  assign n42182 = ~pi219 & ~n42181;
  assign n42183 = pi211 & n42176;
  assign n42184 = ~pi1153 & ~n38329;
  assign n42185 = pi1091 & n42184;
  assign n42186 = n38220 & ~n42185;
  assign n42187 = ~n41977 & n42186;
  assign n42188 = pi219 & ~n42178;
  assign n42189 = ~n42187 & n42188;
  assign n42190 = ~n42183 & n42189;
  assign n42191 = ~n42182 & ~n42190;
  assign n42192 = ~pi254 & ~n42191;
  assign n42193 = pi1091 & ~n11383;
  assign n42194 = ~n38605 & n42193;
  assign n42195 = ~pi1154 & ~n42194;
  assign n42196 = pi1091 & ~n38256;
  assign n42197 = ~n39360 & n40565;
  assign n42198 = ~n42196 & ~n42197;
  assign n42199 = n41985 & ~n42198;
  assign n42200 = n40610 & n41971;
  assign n42201 = pi1154 & ~n42200;
  assign n42202 = ~n42199 & n42201;
  assign n42203 = ~n42195 & ~n42202;
  assign n42204 = pi1091 & ~pi1154;
  assign n42205 = n38350 & n42204;
  assign n42206 = ~n42197 & ~n42205;
  assign n42207 = n11383 & ~n42206;
  assign n42208 = pi254 & ~n42207;
  assign n42209 = ~n42203 & n42208;
  assign n42210 = ~n42192 & ~n42209;
  assign n42211 = ~pi253 & n42210;
  assign n42212 = ~po1038 & ~n42211;
  assign n42213 = ~n42170 & n42212;
  assign n42214 = ~n42130 & ~n42133;
  assign n42215 = ~n41864 & n42117;
  assign n42216 = ~n41889 & n42125;
  assign n42217 = pi253 & ~n42216;
  assign n42218 = ~n42215 & n42217;
  assign n42219 = ~n42214 & ~n42218;
  assign n42220 = ~pi1152 & ~n42219;
  assign n42221 = ~n42213 & n42220;
  assign n42222 = n40648 & ~n42221;
  assign n42223 = ~n42137 & n42222;
  assign n42224 = ~po1038 & ~n42210;
  assign n42225 = ~pi1152 & ~n42130;
  assign n42226 = ~n42224 & n42225;
  assign n42227 = ~po1038 & n42109;
  assign n42228 = pi1152 & n42132;
  assign n42229 = ~n42227 & n42228;
  assign n42230 = ~n40648 & ~n42229;
  assign n42231 = ~n42226 & n42230;
  assign n42232 = ~pi230 & ~n42231;
  assign n42233 = ~n42223 & n42232;
  assign po411 = ~n42039 & ~n42233;
  assign n42235 = ~pi200 & pi1049;
  assign n42236 = pi200 & pi1036;
  assign n42237 = ~n42235 & ~n42236;
  assign n42238 = ~n41728 & n42237;
  assign n42239 = ~pi255 & n41728;
  assign po412 = ~n42238 & ~n42239;
  assign n42241 = ~pi200 & pi1048;
  assign n42242 = pi200 & pi1070;
  assign n42243 = ~n42241 & ~n42242;
  assign n42244 = ~n41728 & n42243;
  assign n42245 = ~pi256 & n41728;
  assign po413 = ~n42244 & ~n42245;
  assign n42247 = ~pi200 & pi1084;
  assign n42248 = pi200 & pi1065;
  assign n42249 = ~n42247 & ~n42248;
  assign n42250 = ~n41728 & n42249;
  assign n42251 = ~pi257 & n41728;
  assign po414 = ~n42250 & ~n42251;
  assign n42253 = ~pi200 & pi1072;
  assign n42254 = pi200 & pi1062;
  assign n42255 = ~n42253 & ~n42254;
  assign n42256 = ~n41728 & n42255;
  assign n42257 = ~pi258 & n41728;
  assign po415 = ~n42256 & ~n42257;
  assign n42259 = ~pi200 & pi1059;
  assign n42260 = pi200 & pi1069;
  assign n42261 = ~n42259 & ~n42260;
  assign n42262 = ~n41728 & n42261;
  assign n42263 = ~pi259 & n41728;
  assign po416 = ~n42262 & ~n42263;
  assign n42265 = pi200 & pi1067;
  assign n42266 = ~pi200 & pi1044;
  assign n42267 = ~pi199 & ~n42266;
  assign n42268 = ~n42265 & n42267;
  assign n42269 = ~n41728 & ~n42268;
  assign n42270 = pi260 & n41728;
  assign po417 = n42269 | n42270;
  assign n42272 = pi200 & pi1040;
  assign n42273 = ~pi200 & pi1037;
  assign n42274 = ~pi199 & ~n42273;
  assign n42275 = ~n42272 & n42274;
  assign n42276 = ~n41728 & ~n42275;
  assign n42277 = pi261 & n41728;
  assign po418 = n42276 | n42277;
  assign n42279 = pi1093 & pi1142;
  assign n42280 = ~pi262 & ~pi1093;
  assign n42281 = ~n42279 & ~n42280;
  assign n42282 = ~pi228 & ~n42281;
  assign n42283 = pi123 & pi262;
  assign n42284 = ~pi123 & ~pi1142;
  assign n42285 = pi228 & ~n42284;
  assign n42286 = ~n42283 & n42285;
  assign n42287 = ~n42282 & ~n42286;
  assign n42288 = ~pi228 & ~pi1093;
  assign n42289 = pi123 & pi228;
  assign n42290 = ~n42288 & ~n42289;
  assign n42291 = ~pi262 & ~n42290;
  assign n42292 = ~n40239 & ~n42291;
  assign n42293 = pi199 & n42290;
  assign n42294 = n38164 & ~n42293;
  assign n42295 = n42292 & ~n42294;
  assign n42296 = ~n42287 & ~n42295;
  assign n42297 = ~pi207 & n42291;
  assign n42298 = ~pi208 & ~n42297;
  assign n42299 = ~n40239 & ~n42298;
  assign n42300 = ~n42296 & ~n42299;
  assign n42301 = pi299 & ~n42292;
  assign n42302 = ~n39315 & n42290;
  assign n42303 = ~pi299 & ~n42302;
  assign n42304 = ~n42287 & n42303;
  assign n42305 = pi208 & ~n42304;
  assign n42306 = ~n42301 & n42305;
  assign n42307 = ~po1038 & ~n42306;
  assign n42308 = ~n42300 & n42307;
  assign n42309 = ~n39402 & n42290;
  assign n42310 = po1038 & ~n42287;
  assign n42311 = ~n42309 & n42310;
  assign po419 = n42308 | n42311;
  assign n42313 = pi1154 & ~n40407;
  assign n42314 = ~n40456 & n42313;
  assign n42315 = ~pi1154 & ~n40429;
  assign n42316 = pi1155 & n42155;
  assign n42317 = n42315 & ~n42316;
  assign n42318 = ~n40474 & n42313;
  assign n42319 = ~pi1156 & ~n42145;
  assign n42320 = ~n42318 & n42319;
  assign n42321 = ~pi1156 & ~n42320;
  assign n42322 = ~n42317 & ~n42321;
  assign n42323 = pi1156 & n42157;
  assign n42324 = ~n42322 & ~n42323;
  assign n42325 = ~n42314 & ~n42324;
  assign n42326 = pi211 & ~n42325;
  assign n42327 = n40409 & ~n40443;
  assign n42328 = pi1155 & n42327;
  assign n42329 = n42315 & ~n42328;
  assign n42330 = n42320 & ~n42329;
  assign n42331 = ~n42157 & n42329;
  assign n42332 = pi1156 & ~n42331;
  assign n42333 = ~n42318 & n42332;
  assign n42334 = ~pi211 & ~n42333;
  assign n42335 = ~n42330 & n42334;
  assign n42336 = ~pi219 & ~n42335;
  assign n42337 = ~n42326 & n42336;
  assign n42338 = ~n40401 & ~n40527;
  assign n42339 = ~n40399 & ~n42161;
  assign n42340 = ~n42338 & ~n42339;
  assign n42341 = ~n40443 & n42340;
  assign n42342 = ~pi1156 & ~n42341;
  assign n42343 = n38211 & ~n42340;
  assign n42344 = ~pi1155 & ~n41834;
  assign n42345 = pi1155 & ~n42051;
  assign n42346 = ~pi1154 & ~n42345;
  assign n42347 = ~n42344 & n42346;
  assign n42348 = pi1154 & ~n42338;
  assign n42349 = n38200 & ~n42348;
  assign n42350 = ~n42347 & n42349;
  assign n42351 = pi219 & ~n42350;
  assign n42352 = ~n42343 & n42351;
  assign n42353 = ~n42342 & n42352;
  assign n42354 = pi263 & ~n42353;
  assign n42355 = ~n42337 & n42354;
  assign n42356 = ~pi1155 & n41922;
  assign n42357 = ~n40444 & n42356;
  assign n42358 = pi1155 & ~n40386;
  assign n42359 = ~pi1154 & ~n42358;
  assign n42360 = ~n42357 & n42359;
  assign n42361 = ~pi1156 & ~n42360;
  assign n42362 = pi1155 & ~n40446;
  assign n42363 = pi1154 & ~n42362;
  assign n42364 = n41817 & n42363;
  assign n42365 = n42361 & ~n42364;
  assign n42366 = ~n41827 & n42359;
  assign n42367 = pi1156 & ~n42366;
  assign n42368 = n40436 & n42363;
  assign n42369 = n42367 & ~n42368;
  assign n42370 = pi211 & ~n42369;
  assign n42371 = ~n42365 & n42370;
  assign n42372 = pi1155 & ~n40486;
  assign n42373 = ~pi1154 & ~n42372;
  assign n42374 = n40425 & n42373;
  assign n42375 = n40417 & n42363;
  assign n42376 = ~n40388 & n42375;
  assign n42377 = ~n42374 & ~n42376;
  assign n42378 = n42367 & n42377;
  assign n42379 = ~n42356 & n42373;
  assign n42380 = ~n42375 & ~n42379;
  assign n42381 = n42361 & n42380;
  assign n42382 = ~pi211 & ~n42381;
  assign n42383 = ~n42378 & n42382;
  assign n42384 = ~pi219 & ~n42383;
  assign n42385 = ~n42371 & n42384;
  assign n42386 = pi1155 & n40384;
  assign n42387 = pi1154 & n40537;
  assign n42388 = ~n42386 & n42387;
  assign n42389 = ~n42379 & ~n42388;
  assign n42390 = ~pi1156 & ~n42389;
  assign n42391 = ~n40390 & n42388;
  assign n42392 = ~n42374 & ~n42391;
  assign n42393 = n38211 & ~n42392;
  assign n42394 = ~pi1154 & n40526;
  assign n42395 = ~n40488 & ~n42394;
  assign n42396 = n38200 & ~n42386;
  assign n42397 = ~n42395 & n42396;
  assign n42398 = pi219 & ~n42397;
  assign n42399 = ~n42393 & n42398;
  assign n42400 = ~n42390 & n42399;
  assign n42401 = ~pi263 & ~n42400;
  assign n42402 = ~n42385 & n42401;
  assign n42403 = n40484 & ~n42402;
  assign n42404 = ~n42355 & n42403;
  assign n42405 = pi1155 & ~n38651;
  assign n42406 = n40588 & ~n42405;
  assign n42407 = ~pi1154 & n42196;
  assign n42408 = ~n42406 & ~n42407;
  assign n42409 = ~n40607 & n42408;
  assign n42410 = n38211 & ~n42409;
  assign n42411 = ~n40561 & ~n42204;
  assign n42412 = ~pi1156 & ~n38280;
  assign n42413 = ~n42411 & n42412;
  assign n42414 = pi219 & ~n42413;
  assign n42415 = ~n38280 & ~n38685;
  assign n42416 = n38200 & n40610;
  assign n42417 = n42415 & n42416;
  assign n42418 = n42414 & ~n42417;
  assign n42419 = ~n42410 & n42418;
  assign n42420 = ~pi211 & ~n42408;
  assign n42421 = ~pi199 & ~pi1154;
  assign n42422 = n38270 & ~n42421;
  assign n42423 = n41949 & ~n42422;
  assign n42424 = ~n38370 & n42423;
  assign n42425 = ~n42420 & ~n42424;
  assign n42426 = pi1156 & ~n42425;
  assign n42427 = ~n38370 & ~n42411;
  assign n42428 = pi211 & n42427;
  assign n42429 = n41997 & n42415;
  assign n42430 = ~n42428 & ~n42429;
  assign n42431 = ~pi1156 & ~n42430;
  assign n42432 = ~pi219 & ~n42431;
  assign n42433 = ~n42426 & n42432;
  assign n42434 = ~n42419 & ~n42433;
  assign n42435 = ~pi263 & ~n42434;
  assign n42436 = ~pi1154 & ~n38366;
  assign n42437 = ~n38340 & n42436;
  assign n42438 = ~n38270 & ~n38308;
  assign n42439 = pi1154 & ~n42438;
  assign n42440 = pi1156 & ~n42439;
  assign n42441 = ~n42437 & n42440;
  assign n42442 = ~pi1156 & n42427;
  assign n42443 = pi211 & ~n42442;
  assign n42444 = ~n42441 & n42443;
  assign n42445 = ~n38285 & n39110;
  assign n42446 = ~n38685 & ~n42445;
  assign n42447 = ~pi211 & ~n42446;
  assign n42448 = ~pi219 & ~n42447;
  assign n42449 = ~n42444 & n42448;
  assign n42450 = pi1154 & ~n38282;
  assign n42451 = pi1156 & ~n42450;
  assign n42452 = ~pi299 & ~n42451;
  assign n42453 = ~n38283 & ~n39482;
  assign n42454 = ~n42452 & n42453;
  assign n42455 = pi1156 & ~n42454;
  assign n42456 = ~n42415 & n42452;
  assign n42457 = pi219 & ~n42456;
  assign n42458 = ~n42455 & n42457;
  assign n42459 = pi263 & pi1091;
  assign n42460 = ~n42458 & n42459;
  assign n42461 = ~n42449 & n42460;
  assign n42462 = ~n42435 & ~n42461;
  assign n42463 = ~n40484 & ~n42462;
  assign n42464 = ~po1038 & ~n42463;
  assign n42465 = ~n42404 & n42464;
  assign n42466 = pi211 & n40367;
  assign n42467 = ~pi211 & ~n42204;
  assign n42468 = ~n38201 & ~n42467;
  assign n42469 = ~n42466 & n42468;
  assign n42470 = ~n40376 & ~n42469;
  assign n42471 = ~pi219 & ~n42470;
  assign n42472 = ~pi263 & ~n42119;
  assign n42473 = ~n42471 & n42472;
  assign n42474 = ~n38201 & ~n42097;
  assign n42475 = ~n42466 & ~n42474;
  assign n42476 = n41849 & ~n42475;
  assign n42477 = pi263 & ~n41853;
  assign n42478 = ~n42476 & n42477;
  assign n42479 = ~n42473 & ~n42478;
  assign n42480 = pi219 & ~n38200;
  assign n42481 = pi1091 & n42480;
  assign n42482 = n40484 & ~n42481;
  assign n42483 = ~n42479 & n42482;
  assign n42484 = ~pi219 & ~n38201;
  assign n42485 = ~n38220 & n42484;
  assign n42486 = ~n42480 & ~n42485;
  assign n42487 = pi1091 & ~n42486;
  assign n42488 = pi263 & ~pi1091;
  assign n42489 = ~n42487 & ~n42488;
  assign n42490 = ~n40484 & n42489;
  assign n42491 = po1038 & ~n42490;
  assign n42492 = ~n42483 & n42491;
  assign n42493 = n40648 & ~n42492;
  assign n42494 = ~n42465 & n42493;
  assign n42495 = ~po1038 & n42462;
  assign n42496 = po1038 & ~n42489;
  assign n42497 = ~n40648 & ~n42496;
  assign n42498 = ~n42495 & n42497;
  assign n42499 = ~pi230 & ~n42498;
  assign n42500 = ~n42494 & n42499;
  assign n42501 = ~n38281 & n38286;
  assign n42502 = ~pi1156 & ~n42501;
  assign n42503 = ~pi299 & ~n38282;
  assign n42504 = ~pi200 & n42421;
  assign n42505 = n42503 & ~n42504;
  assign n42506 = ~n42502 & n42505;
  assign n42507 = ~n38232 & ~n42506;
  assign n42508 = pi211 & ~n42507;
  assign n42509 = n42448 & ~n42508;
  assign n42510 = pi1156 & n39482;
  assign n42511 = pi219 & ~n42510;
  assign n42512 = ~n42506 & n42511;
  assign n42513 = ~po1038 & ~n42512;
  assign n42514 = ~n42509 & n42513;
  assign n42515 = po1038 & n42486;
  assign n42516 = pi230 & ~n42515;
  assign n42517 = ~n42514 & n42516;
  assign po420 = ~n42500 & ~n42517;
  assign n42519 = pi264 & ~n40371;
  assign n42520 = ~pi796 & n40371;
  assign n42521 = ~pi1091 & ~n42520;
  assign n42522 = ~n42519 & n42521;
  assign n42523 = pi1091 & pi1142;
  assign n42524 = ~n42522 & ~n42523;
  assign n42525 = pi200 & ~n42524;
  assign n42526 = pi1091 & pi1141;
  assign n42527 = ~n42522 & ~n42526;
  assign n42528 = ~pi200 & ~n42527;
  assign n42529 = ~pi199 & ~n42528;
  assign n42530 = ~n42525 & n42529;
  assign n42531 = pi264 & ~n40360;
  assign n42532 = ~pi796 & n40360;
  assign n42533 = ~pi1091 & ~n42532;
  assign n42534 = ~n42531 & n42533;
  assign n42535 = pi1091 & pi1143;
  assign n42536 = ~pi200 & n42535;
  assign n42537 = pi199 & ~n42536;
  assign n42538 = ~n42534 & n42537;
  assign n42539 = n16361 & ~n42538;
  assign n42540 = ~n42530 & n42539;
  assign n42541 = pi211 & ~n42524;
  assign n42542 = ~pi211 & ~n42527;
  assign n42543 = ~pi219 & ~n42542;
  assign n42544 = ~n42541 & n42543;
  assign n42545 = pi219 & ~n41997;
  assign n42546 = ~n39002 & ~n42545;
  assign n42547 = ~n42534 & ~n42546;
  assign n42548 = ~n16361 & ~n42547;
  assign n42549 = ~n42544 & n42548;
  assign n42550 = ~n42540 & ~n42549;
  assign n42551 = ~pi230 & ~n42550;
  assign n42552 = ~pi199 & pi1141;
  assign n42553 = n39007 & ~n42552;
  assign n42554 = ~n38166 & ~n42553;
  assign n42555 = n16361 & ~n42554;
  assign n42556 = ~pi211 & pi1141;
  assign n42557 = ~pi219 & ~n38180;
  assign n42558 = ~n42556 & n42557;
  assign n42559 = ~n39002 & ~n42558;
  assign n42560 = ~n16361 & ~n42559;
  assign n42561 = pi230 & ~n42560;
  assign n42562 = ~n42555 & n42561;
  assign po421 = n42551 | n42562;
  assign n42564 = pi265 & ~n40371;
  assign n42565 = ~pi819 & n40371;
  assign n42566 = ~pi1091 & ~n42565;
  assign n42567 = ~n42564 & n42566;
  assign n42568 = ~n42535 & ~n42567;
  assign n42569 = pi200 & ~n42568;
  assign n42570 = ~n42523 & ~n42567;
  assign n42571 = ~pi200 & ~n42570;
  assign n42572 = ~pi199 & ~n42571;
  assign n42573 = ~n42569 & n42572;
  assign n42574 = pi265 & ~n40360;
  assign n42575 = ~pi819 & n40360;
  assign n42576 = ~pi1091 & ~n42575;
  assign n42577 = ~n42574 & n42576;
  assign n42578 = pi1091 & pi1144;
  assign n42579 = ~pi200 & n42578;
  assign n42580 = pi199 & ~n42579;
  assign n42581 = ~n42577 & n42580;
  assign n42582 = n16361 & ~n42581;
  assign n42583 = ~n42573 & n42582;
  assign n42584 = pi211 & ~n42568;
  assign n42585 = ~pi211 & ~n42570;
  assign n42586 = ~pi219 & ~n42585;
  assign n42587 = ~n42584 & n42586;
  assign n42588 = ~n40321 & ~n42545;
  assign n42589 = ~n42577 & ~n42588;
  assign n42590 = ~n16361 & ~n42589;
  assign n42591 = ~n42587 & n42590;
  assign n42592 = ~n42583 & ~n42591;
  assign n42593 = ~pi230 & ~n42592;
  assign n42594 = ~n38165 & n40281;
  assign n42595 = ~n38159 & ~n42594;
  assign n42596 = n16361 & ~n42595;
  assign n42597 = ~pi211 & pi1142;
  assign n42598 = ~pi219 & ~n38140;
  assign n42599 = ~n42597 & n42598;
  assign n42600 = ~n40321 & ~n42599;
  assign n42601 = ~n16361 & ~n42600;
  assign n42602 = pi230 & ~n42601;
  assign n42603 = ~n42596 & n42602;
  assign po422 = n42593 | n42603;
  assign n42605 = ~pi211 & pi1136;
  assign n42606 = pi219 & ~n42605;
  assign n42607 = pi211 & ~pi1135;
  assign n42608 = ~n42606 & ~n42607;
  assign n42609 = ~n10670 & n42608;
  assign n42610 = pi299 & n42609;
  assign n42611 = pi199 & pi1136;
  assign n42612 = ~pi200 & ~n42611;
  assign n42613 = ~pi199 & pi1135;
  assign n42614 = pi200 & ~n42613;
  assign n42615 = ~pi299 & ~n42614;
  assign n42616 = ~n42612 & n42615;
  assign n42617 = ~n42610 & ~n42616;
  assign n42618 = ~po1038 & ~n42617;
  assign n42619 = po1038 & n42609;
  assign n42620 = pi230 & ~n42619;
  assign n42621 = ~n42618 & n42620;
  assign n42622 = ~pi948 & n40371;
  assign n42623 = ~pi266 & ~n40371;
  assign n42624 = ~pi1091 & ~n42623;
  assign n42625 = ~n42622 & n42624;
  assign n42626 = ~pi199 & ~n42625;
  assign n42627 = pi1091 & pi1136;
  assign n42628 = ~pi948 & n40360;
  assign n42629 = ~pi266 & ~n40360;
  assign n42630 = ~pi1091 & ~n42629;
  assign n42631 = ~n42628 & n42630;
  assign n42632 = pi199 & ~n42631;
  assign n42633 = ~n42627 & n42632;
  assign n42634 = ~n42626 & ~n42633;
  assign n42635 = ~pi200 & n42634;
  assign n42636 = pi1091 & pi1135;
  assign n42637 = n42626 & ~n42636;
  assign n42638 = pi200 & ~n42632;
  assign n42639 = ~n42637 & n42638;
  assign n42640 = ~n42635 & ~n42639;
  assign n42641 = n16361 & ~n42640;
  assign n42642 = ~n42545 & ~n42606;
  assign n42643 = ~n42631 & ~n42642;
  assign n42644 = ~n16361 & ~n42643;
  assign n42645 = ~pi219 & ~n42625;
  assign n42646 = pi1135 & n41949;
  assign n42647 = n42645 & ~n42646;
  assign n42648 = n42644 & ~n42647;
  assign n42649 = ~pi230 & ~n42648;
  assign n42650 = ~n42641 & n42649;
  assign n42651 = ~n42621 & ~n42650;
  assign n42652 = ~pi1134 & ~n42651;
  assign n42653 = ~n16361 & n42608;
  assign n42654 = ~n39904 & ~n42616;
  assign n42655 = ~po1038 & ~n42654;
  assign n42656 = pi230 & ~n42655;
  assign n42657 = ~n42653 & n42656;
  assign n42658 = ~pi199 & pi1091;
  assign n42659 = ~n42634 & ~n42658;
  assign n42660 = ~pi200 & ~n42659;
  assign n42661 = ~n42639 & ~n42660;
  assign n42662 = n16361 & ~n42661;
  assign n42663 = pi1091 & ~n42607;
  assign n42664 = n42645 & ~n42663;
  assign n42665 = n42644 & ~n42664;
  assign n42666 = ~pi230 & ~n42665;
  assign n42667 = ~n42662 & n42666;
  assign n42668 = ~n42657 & ~n42667;
  assign n42669 = pi1134 & ~n42668;
  assign po423 = ~n42652 & ~n42669;
  assign n42671 = ~n42067 & n42070;
  assign n42672 = n42138 & ~n42671;
  assign n42673 = pi1154 & pi1155;
  assign n42674 = ~n40399 & n42673;
  assign n42675 = ~n42075 & n42674;
  assign n42676 = ~n42672 & ~n42675;
  assign n42677 = pi211 & ~n42676;
  assign n42678 = n38204 & ~n41834;
  assign n42679 = ~n41840 & n42678;
  assign n42680 = ~n42052 & n42679;
  assign n42681 = n40526 & n42046;
  assign n42682 = ~pi1155 & ~n42681;
  assign n42683 = ~n42671 & n42682;
  assign n42684 = ~pi267 & ~n42683;
  assign n42685 = ~n42680 & n42684;
  assign n42686 = ~n42677 & n42685;
  assign n42687 = n40486 & ~n42062;
  assign n42688 = pi1154 & ~n42687;
  assign n42689 = ~pi1154 & ~n40537;
  assign n42690 = ~n41923 & n42689;
  assign n42691 = ~pi1155 & ~n42690;
  assign n42692 = ~n42688 & n42691;
  assign n42693 = pi1155 & ~n41902;
  assign n42694 = n40384 & ~n42394;
  assign n42695 = n42693 & ~n42694;
  assign n42696 = ~n41921 & n42695;
  assign n42697 = pi267 & ~n42696;
  assign n42698 = ~n42692 & n42697;
  assign n42699 = ~n42686 & ~n42698;
  assign n42700 = pi219 & ~n42699;
  assign n42701 = ~n41840 & ~n42157;
  assign n42702 = n42345 & n42701;
  assign n42703 = pi1154 & ~n42702;
  assign n42704 = ~pi1153 & ~n40446;
  assign n42705 = ~pi1154 & ~n42704;
  assign n42706 = pi1155 & ~n42705;
  assign n42707 = n40431 & ~n42706;
  assign n42708 = ~n42703 & ~n42707;
  assign n42709 = ~pi1155 & ~n42155;
  assign n42710 = ~n42671 & n42709;
  assign n42711 = pi211 & ~n42710;
  assign n42712 = ~n42708 & n42711;
  assign n42713 = pi1153 & ~n40444;
  assign n42714 = ~pi1155 & ~n42713;
  assign n42715 = ~pi1153 & ~n42327;
  assign n42716 = n42714 & ~n42715;
  assign n42717 = pi1155 & ~n42701;
  assign n42718 = pi1154 & ~n42328;
  assign n42719 = ~n42717 & n42718;
  assign n42720 = ~n42716 & n42719;
  assign n42721 = n41917 & n42714;
  assign n42722 = ~pi1154 & ~n42717;
  assign n42723 = ~n42721 & n42722;
  assign n42724 = ~pi211 & ~n42723;
  assign n42725 = ~n42720 & n42724;
  assign n42726 = ~pi267 & ~n42725;
  assign n42727 = ~n42712 & n42726;
  assign n42728 = n41826 & n42693;
  assign n42729 = ~pi1153 & n40465;
  assign n42730 = ~n40446 & ~n42729;
  assign n42731 = ~pi1155 & n40386;
  assign n42732 = ~n42730 & n42731;
  assign n42733 = pi1154 & ~n42732;
  assign n42734 = ~n42728 & n42733;
  assign n42735 = ~pi1153 & n40444;
  assign n42736 = ~pi1154 & ~n42735;
  assign n42737 = ~n40417 & n42736;
  assign n42738 = ~pi1155 & ~n42737;
  assign n42739 = ~n40436 & n42736;
  assign n42740 = ~n42738 & n42739;
  assign n42741 = ~n42734 & ~n42740;
  assign n42742 = pi211 & ~n42741;
  assign n42743 = pi1154 & n42730;
  assign n42744 = n42738 & ~n42743;
  assign n42745 = ~n40409 & ~n42040;
  assign n42746 = pi1154 & n40384;
  assign n42747 = pi1155 & ~n42746;
  assign n42748 = ~n42745 & n42747;
  assign n42749 = ~pi211 & ~n42748;
  assign n42750 = ~n42744 & n42749;
  assign n42751 = pi267 & ~n42750;
  assign n42752 = ~n42742 & n42751;
  assign n42753 = ~pi219 & ~n42752;
  assign n42754 = ~n42727 & n42753;
  assign n42755 = ~n42700 & ~n42754;
  assign n42756 = n40483 & ~n42755;
  assign n42757 = ~n38330 & ~n40565;
  assign n42758 = pi1153 & ~n10761;
  assign n42759 = pi1091 & ~n42758;
  assign n42760 = ~n42757 & n42759;
  assign n42761 = ~pi1154 & n42760;
  assign n42762 = ~pi219 & ~n42761;
  assign n42763 = pi1155 & n38628;
  assign n42764 = pi1154 & ~n42763;
  assign n42765 = pi1091 & n42764;
  assign n42766 = ~n11382 & ~n42087;
  assign n42767 = n42765 & n42766;
  assign n42768 = n42762 & ~n42767;
  assign n42769 = pi1091 & n42405;
  assign n42770 = ~n42086 & n42769;
  assign n42771 = pi1154 & ~n42770;
  assign n42772 = ~pi299 & n38612;
  assign n42773 = pi1091 & ~n42772;
  assign n42774 = n42771 & n42773;
  assign n42775 = ~n41786 & ~n42184;
  assign n42776 = ~n38330 & n42204;
  assign n42777 = ~n42775 & n42776;
  assign n42778 = n42204 & ~n42777;
  assign n42779 = pi219 & ~n42778;
  assign n42780 = ~n42774 & n42779;
  assign n42781 = ~n42768 & ~n42780;
  assign n42782 = ~pi211 & ~n42781;
  assign n42783 = ~pi1155 & ~n38613;
  assign n42784 = ~n38365 & ~n42783;
  assign n42785 = ~n12979 & ~n42784;
  assign n42786 = n42765 & ~n42785;
  assign n42787 = pi1153 & n38620;
  assign n42788 = n42204 & ~n42787;
  assign n42789 = ~n42757 & n42788;
  assign n42790 = pi211 & ~n42789;
  assign n42791 = ~n42786 & n42790;
  assign n42792 = ~n42782 & ~n42791;
  assign n42793 = pi267 & ~n42792;
  assign n42794 = ~n38311 & ~n38342;
  assign n42795 = ~n38650 & n42794;
  assign n42796 = pi1091 & n42795;
  assign n42797 = ~pi211 & ~n42796;
  assign n42798 = pi1091 & ~pi1155;
  assign n42799 = ~n38613 & n42798;
  assign n42800 = n38205 & ~n42799;
  assign n42801 = ~n42770 & n42800;
  assign n42802 = ~pi219 & ~n42801;
  assign n42803 = ~n42797 & n42802;
  assign n42804 = n42772 & n42798;
  assign n42805 = n42771 & ~n42804;
  assign n42806 = pi1154 & ~n42805;
  assign n42807 = ~pi211 & ~n42777;
  assign n42808 = ~n42806 & n42807;
  assign n42809 = n42405 & n42764;
  assign n42810 = ~n42805 & ~n42809;
  assign n42811 = pi211 & ~n42810;
  assign n42812 = pi219 & ~n42811;
  assign n42813 = ~n42808 & n42812;
  assign n42814 = ~n42803 & ~n42813;
  assign n42815 = pi211 & ~pi1154;
  assign n42816 = n40556 & ~n42760;
  assign n42817 = n42815 & ~n42816;
  assign n42818 = ~pi267 & ~n42817;
  assign n42819 = ~n42814 & n42818;
  assign n42820 = ~n42793 & ~n42819;
  assign n42821 = ~n40483 & ~n42820;
  assign n42822 = ~po1038 & ~n42821;
  assign n42823 = ~n42756 & n42822;
  assign n42824 = pi267 & n42121;
  assign n42825 = ~pi267 & ~n40378;
  assign n42826 = ~n41853 & n42825;
  assign n42827 = n40483 & ~n42826;
  assign n42828 = ~n42824 & n42827;
  assign n42829 = ~pi219 & ~n38205;
  assign n42830 = ~n38222 & n42829;
  assign n42831 = ~n38899 & ~n42830;
  assign n42832 = pi1091 & ~n42831;
  assign n42833 = ~pi267 & ~pi1091;
  assign n42834 = ~n40483 & n42833;
  assign n42835 = ~n42832 & ~n42834;
  assign n42836 = ~n42828 & n42835;
  assign n42837 = po1038 & ~n42836;
  assign n42838 = n40648 & ~n42837;
  assign n42839 = ~n42823 & n42838;
  assign n42840 = ~po1038 & n42820;
  assign n42841 = ~n42832 & ~n42833;
  assign n42842 = po1038 & ~n42841;
  assign n42843 = ~n40648 & ~n42842;
  assign n42844 = ~n42840 & n42843;
  assign n42845 = ~pi230 & ~n42844;
  assign n42846 = ~n42839 & n42845;
  assign n42847 = pi219 & ~n38628;
  assign n42848 = ~pi1155 & n42787;
  assign n42849 = ~pi1154 & ~n42848;
  assign n42850 = ~n38613 & ~n42849;
  assign n42851 = n38270 & ~n38623;
  assign n42852 = pi1155 & n42851;
  assign n42853 = ~n42850 & ~n42852;
  assign n42854 = ~n42847 & ~n42853;
  assign n42855 = pi211 & ~n42854;
  assign n42856 = ~pi199 & pi1154;
  assign n42857 = pi200 & ~n42856;
  assign n42858 = ~n38321 & ~n38627;
  assign n42859 = ~n42857 & n42858;
  assign n42860 = ~n38232 & ~n42859;
  assign n42861 = pi219 & ~n42860;
  assign n42862 = ~pi219 & n42795;
  assign n42863 = ~pi211 & ~n42862;
  assign n42864 = ~n42861 & n42863;
  assign n42865 = ~po1038 & ~n42864;
  assign n42866 = ~n42855 & n42865;
  assign n42867 = po1038 & n42831;
  assign n42868 = pi230 & ~n42867;
  assign n42869 = ~n42866 & n42868;
  assign po424 = ~n42846 & ~n42869;
  assign n42871 = ~n41863 & n41891;
  assign n42872 = ~po1038 & ~n41821;
  assign n42873 = ~n41819 & ~n41872;
  assign n42874 = ~pi219 & n40465;
  assign n42875 = n41836 & ~n42874;
  assign n42876 = ~n42873 & ~n42875;
  assign n42877 = n42872 & ~n42876;
  assign n42878 = ~n42871 & ~n42877;
  assign n42879 = ~pi1151 & ~n42878;
  assign n42880 = ~po1038 & ~n41830;
  assign n42881 = pi219 & n40531;
  assign n42882 = n42880 & ~n42881;
  assign n42883 = n41891 & ~n42120;
  assign n42884 = ~n42882 & ~n42883;
  assign n42885 = pi1151 & ~n42884;
  assign n42886 = ~n42879 & ~n42885;
  assign n42887 = pi268 & ~n42886;
  assign n42888 = po1038 & ~n41853;
  assign n42889 = ~n41888 & n42888;
  assign n42890 = po1038 & ~n42119;
  assign n42891 = ~n41856 & n42890;
  assign n42892 = n42889 & ~n42891;
  assign n42893 = pi219 & ~n40395;
  assign n42894 = ~n41877 & ~n42893;
  assign n42895 = ~n40396 & ~n42894;
  assign n42896 = ~po1038 & ~n40443;
  assign n42897 = n42895 & n42896;
  assign n42898 = ~n42892 & ~n42897;
  assign n42899 = ~pi1151 & n42898;
  assign n42900 = ~n40367 & ~n42884;
  assign n42901 = ~n40542 & n42880;
  assign n42902 = pi219 & po1038;
  assign n42903 = ~n40394 & n42902;
  assign n42904 = ~n41849 & ~n42903;
  assign n42905 = ~n42901 & n42904;
  assign n42906 = ~n42900 & ~n42905;
  assign n42907 = pi1151 & n42906;
  assign n42908 = ~pi268 & ~n42907;
  assign n42909 = ~n42899 & n42908;
  assign n42910 = ~n42887 & ~n42909;
  assign n42911 = ~pi1152 & ~n42910;
  assign n42912 = ~n41863 & n42890;
  assign n42913 = ~n40488 & ~n41924;
  assign n42914 = n42876 & ~n42913;
  assign n42915 = ~po1038 & ~n42914;
  assign n42916 = ~n40394 & ~n41905;
  assign n42917 = n42915 & ~n42916;
  assign n42918 = ~n42912 & ~n42917;
  assign n42919 = ~pi1151 & ~n42918;
  assign n42920 = ~n40363 & n42872;
  assign n42921 = n42884 & ~n42891;
  assign n42922 = ~n42920 & n42921;
  assign n42923 = pi1151 & ~n42922;
  assign n42924 = pi268 & ~n42923;
  assign n42925 = ~n42919 & n42924;
  assign n42926 = ~n41835 & ~n42895;
  assign n42927 = ~po1038 & ~n42926;
  assign n42928 = ~n42889 & ~n42927;
  assign n42929 = ~pi1151 & ~n42928;
  assign n42930 = ~po1038 & ~n42875;
  assign n42931 = ~n41864 & n42888;
  assign n42932 = ~n42892 & ~n42931;
  assign n42933 = ~n42930 & n42932;
  assign n42934 = pi1151 & ~n42933;
  assign n42935 = ~pi268 & ~n42934;
  assign n42936 = ~n42929 & n42935;
  assign n42937 = pi1152 & ~n42936;
  assign n42938 = ~n42925 & n42937;
  assign n42939 = ~n42911 & ~n42938;
  assign n42940 = pi1150 & ~n42939;
  assign n42941 = ~po1038 & n42876;
  assign n42942 = ~n42931 & ~n42941;
  assign n42943 = pi1151 & ~n42942;
  assign n42944 = ~n41849 & n42888;
  assign n42945 = ~n42882 & n42930;
  assign n42946 = ~n42944 & ~n42945;
  assign n42947 = ~pi1151 & ~n42946;
  assign n42948 = pi1152 & ~n42947;
  assign n42949 = ~n42943 & n42948;
  assign n42950 = ~n41865 & ~n42903;
  assign n42951 = ~n42915 & n42950;
  assign n42952 = pi1151 & n42951;
  assign n42953 = ~pi1151 & n42905;
  assign n42954 = ~pi1152 & ~n42953;
  assign n42955 = ~n42952 & n42954;
  assign n42956 = ~n42949 & ~n42955;
  assign n42957 = ~pi268 & ~n42956;
  assign n42958 = ~n41889 & n42890;
  assign n42959 = pi219 & ~n41921;
  assign n42960 = ~n41877 & ~n42959;
  assign n42961 = n40414 & ~n42960;
  assign n42962 = ~po1038 & ~n42961;
  assign n42963 = ~n42958 & ~n42962;
  assign n42964 = pi1151 & n42963;
  assign n42965 = ~po1038 & ~n41924;
  assign n42966 = ~n42959 & n42965;
  assign n42967 = ~n42891 & ~n42966;
  assign n42968 = ~pi1151 & n42967;
  assign n42969 = pi1152 & ~n42968;
  assign n42970 = ~n42964 & n42969;
  assign n42971 = ~po1038 & ~n41879;
  assign n42972 = ~n41877 & n42971;
  assign n42973 = ~n41892 & ~n42972;
  assign n42974 = pi1151 & n42973;
  assign n42975 = n40367 & ~n42884;
  assign n42976 = ~pi1151 & ~n42975;
  assign n42977 = ~pi1152 & ~n42976;
  assign n42978 = ~n42974 & n42977;
  assign n42979 = pi268 & ~n42978;
  assign n42980 = ~n42970 & n42979;
  assign n42981 = ~pi1150 & ~n42980;
  assign n42982 = ~n42957 & n42981;
  assign n42983 = ~n42940 & ~n42982;
  assign n42984 = n40647 & ~n42983;
  assign n42985 = pi268 & pi1152;
  assign n42986 = ~pi199 & n16361;
  assign n42987 = ~n39727 & ~n42986;
  assign n42988 = ~pi211 & ~n16361;
  assign n42989 = ~po1038 & n38270;
  assign n42990 = ~n42988 & ~n42989;
  assign n42991 = pi1152 & ~n42990;
  assign n42992 = n42987 & ~n42991;
  assign n42993 = ~pi1151 & n42990;
  assign n42994 = pi1150 & ~n42993;
  assign n42995 = ~n42992 & n42994;
  assign n42996 = ~n42985 & n42995;
  assign n42997 = ~n16361 & n41985;
  assign n42998 = ~po1038 & n38320;
  assign n42999 = ~n42997 & ~n42998;
  assign n43000 = pi1151 & ~n42999;
  assign n43001 = pi1152 & n43000;
  assign n43002 = ~po1038 & ~n11385;
  assign n43003 = po1038 & n11383;
  assign n43004 = ~n43002 & ~n43003;
  assign n43005 = pi1151 & ~n43004;
  assign n43006 = ~pi1152 & ~n43005;
  assign n43007 = ~pi1151 & n41783;
  assign n43008 = ~pi1150 & ~n43007;
  assign n43009 = ~n43006 & n43008;
  assign n43010 = ~n43001 & n43009;
  assign n43011 = ~n42996 & ~n43010;
  assign n43012 = pi1091 & ~n43011;
  assign n43013 = pi1152 & n42995;
  assign n43014 = pi1091 & ~n43013;
  assign n43015 = pi268 & ~n43014;
  assign n43016 = ~n43012 & ~n43015;
  assign n43017 = ~n40647 & ~n43016;
  assign n43018 = ~pi230 & ~n43017;
  assign n43019 = ~n42984 & n43018;
  assign n43020 = pi230 & ~n42995;
  assign n43021 = ~n43010 & n43020;
  assign po425 = ~n43019 & ~n43021;
  assign n43023 = ~pi199 & pi1137;
  assign n43024 = pi200 & ~n43023;
  assign n43025 = ~pi199 & pi1136;
  assign n43026 = pi199 & pi1138;
  assign n43027 = ~pi200 & ~n43026;
  assign n43028 = ~n43025 & n43027;
  assign n43029 = ~n43024 & ~n43028;
  assign n43030 = n16361 & ~n43029;
  assign n43031 = ~pi211 & pi1138;
  assign n43032 = pi219 & n43031;
  assign n43033 = pi211 & pi1137;
  assign n43034 = ~n42605 & ~n43033;
  assign n43035 = ~pi219 & ~n43034;
  assign n43036 = ~n43032 & ~n43035;
  assign n43037 = ~n16361 & n43036;
  assign n43038 = ~n43030 & ~n43037;
  assign n43039 = pi230 & ~n43038;
  assign n43040 = ~pi200 & n42627;
  assign n43041 = pi1137 & n40587;
  assign n43042 = ~n43040 & ~n43041;
  assign n43043 = n42986 & n43042;
  assign n43044 = pi1091 & ~n43034;
  assign n43045 = n39727 & ~n43044;
  assign n43046 = ~n43043 & ~n43045;
  assign n43047 = pi269 & ~n40371;
  assign n43048 = ~pi817 & n40371;
  assign n43049 = ~pi1091 & ~n43048;
  assign n43050 = ~n43047 & n43049;
  assign n43051 = ~n43046 & ~n43050;
  assign n43052 = pi269 & ~n40360;
  assign n43053 = ~pi817 & n40360;
  assign n43054 = ~pi1091 & ~n43053;
  assign n43055 = ~n43052 & n43054;
  assign n43056 = pi1138 & n41997;
  assign n43057 = pi219 & ~n16361;
  assign n43058 = ~n43056 & n43057;
  assign n43059 = ~pi200 & pi1091;
  assign n43060 = pi1138 & n43059;
  assign n43061 = pi199 & ~n43060;
  assign n43062 = n16361 & n43061;
  assign n43063 = ~n43058 & ~n43062;
  assign n43064 = ~n43055 & ~n43063;
  assign n43065 = ~n43051 & ~n43064;
  assign n43066 = ~pi230 & ~n43065;
  assign po426 = ~n43039 & ~n43066;
  assign n43068 = pi270 & ~n40371;
  assign n43069 = ~pi805 & n40371;
  assign n43070 = ~pi1091 & ~n43069;
  assign n43071 = ~n43068 & n43070;
  assign n43072 = ~pi211 & pi1139;
  assign n43073 = pi211 & pi1140;
  assign n43074 = ~n43072 & ~n43073;
  assign n43075 = pi1091 & ~n43074;
  assign n43076 = n39727 & ~n43075;
  assign n43077 = pi1091 & pi1140;
  assign n43078 = pi200 & n43077;
  assign n43079 = pi1139 & n43059;
  assign n43080 = ~n43078 & ~n43079;
  assign n43081 = n42986 & n43080;
  assign n43082 = ~n43076 & ~n43081;
  assign n43083 = ~n43071 & ~n43082;
  assign n43084 = pi270 & ~n40360;
  assign n43085 = ~pi805 & n40360;
  assign n43086 = ~pi1091 & ~n43085;
  assign n43087 = ~n43084 & n43086;
  assign n43088 = n41997 & n42556;
  assign n43089 = n43057 & ~n43088;
  assign n43090 = ~pi200 & n42526;
  assign n43091 = pi199 & ~n43090;
  assign n43092 = n16361 & n43091;
  assign n43093 = ~n43089 & ~n43092;
  assign n43094 = ~n43087 & ~n43093;
  assign n43095 = ~pi230 & ~n43094;
  assign n43096 = ~n43083 & n43095;
  assign n43097 = ~pi199 & pi1140;
  assign n43098 = pi200 & ~n43097;
  assign n43099 = ~pi199 & pi1139;
  assign n43100 = pi199 & pi1141;
  assign n43101 = ~pi200 & ~n43100;
  assign n43102 = ~n43099 & n43101;
  assign n43103 = ~n43098 & ~n43102;
  assign n43104 = n16361 & ~n43103;
  assign n43105 = pi219 & ~n42556;
  assign n43106 = ~pi219 & n43074;
  assign n43107 = ~n43105 & ~n43106;
  assign n43108 = ~n16361 & ~n43107;
  assign n43109 = pi230 & ~n43108;
  assign n43110 = ~n43104 & n43109;
  assign po427 = n43096 | n43110;
  assign n43112 = ~pi271 & ~n40392;
  assign n43113 = ~n40364 & ~n43112;
  assign n43114 = pi219 & ~n43113;
  assign n43115 = pi1091 & pi1146;
  assign n43116 = ~n40374 & ~n43113;
  assign n43117 = ~n40375 & ~n43116;
  assign n43118 = ~n43115 & ~n43117;
  assign n43119 = ~pi211 & n43115;
  assign n43120 = ~n43118 & ~n43119;
  assign n43121 = pi1091 & n38994;
  assign n43122 = ~pi219 & ~n43121;
  assign n43123 = ~n43120 & n43122;
  assign n43124 = ~n43114 & ~n43123;
  assign n43125 = ~pi211 & pi1147;
  assign n43126 = n41847 & n43125;
  assign n43127 = ~n16361 & ~n43126;
  assign n43128 = ~n43124 & n43127;
  assign n43129 = pi199 & ~n43113;
  assign n43130 = ~pi199 & n43118;
  assign n43131 = ~n43129 & ~n43130;
  assign n43132 = pi200 & ~n43131;
  assign n43133 = pi1091 & pi1145;
  assign n43134 = ~pi199 & ~n43133;
  assign n43135 = ~n43117 & n43134;
  assign n43136 = ~n43129 & ~n43135;
  assign n43137 = pi1147 & n40573;
  assign n43138 = ~pi200 & ~n43137;
  assign n43139 = ~n43136 & n43138;
  assign n43140 = ~n43132 & ~n43139;
  assign n43141 = n16361 & ~n43140;
  assign n43142 = ~n43128 & ~n43141;
  assign n43143 = ~pi230 & ~n43142;
  assign n43144 = ~pi200 & ~n39012;
  assign n43145 = n39898 & ~n43144;
  assign n43146 = pi1147 & n41779;
  assign n43147 = ~n39785 & ~n39798;
  assign n43148 = ~pi219 & ~n43147;
  assign n43149 = ~n43146 & ~n43148;
  assign n43150 = ~n43145 & n43149;
  assign n43151 = ~po1038 & ~n43150;
  assign n43152 = pi219 & ~n43125;
  assign n43153 = ~n38994 & n40745;
  assign n43154 = ~n43152 & ~n43153;
  assign n43155 = po1038 & n43154;
  assign n43156 = pi230 & ~n43155;
  assign n43157 = ~n43151 & n43156;
  assign po428 = ~n43143 & ~n43157;
  assign n43159 = pi1150 & ~n42933;
  assign n43160 = ~pi1150 & ~n42906;
  assign n43161 = pi1149 & ~n43160;
  assign n43162 = ~n43159 & n43161;
  assign n43163 = pi1150 & ~n42928;
  assign n43164 = ~pi1150 & ~n42898;
  assign n43165 = ~pi1149 & ~n43164;
  assign n43166 = ~n43163 & n43165;
  assign n43167 = ~n43162 & ~n43166;
  assign n43168 = pi1148 & ~n43167;
  assign n43169 = ~pi1150 & ~n42951;
  assign n43170 = pi1150 & n42942;
  assign n43171 = pi1149 & ~n43170;
  assign n43172 = ~n43169 & n43171;
  assign n43173 = pi1150 & n42946;
  assign n43174 = ~pi1150 & ~n42905;
  assign n43175 = ~pi1149 & ~n43174;
  assign n43176 = ~n43173 & n43175;
  assign n43177 = ~pi1148 & ~n43176;
  assign n43178 = ~n43172 & n43177;
  assign n43179 = ~n43168 & ~n43178;
  assign n43180 = pi283 & ~n43179;
  assign n43181 = po1038 & n10670;
  assign n43182 = ~n12982 & ~n43181;
  assign n43183 = ~pi1150 & n43182;
  assign n43184 = ~n42990 & ~n43183;
  assign n43185 = ~pi1149 & ~n43184;
  assign n43186 = pi1149 & ~pi1150;
  assign n43187 = ~n42990 & ~n43186;
  assign n43188 = n42987 & ~n43187;
  assign n43189 = ~n43185 & ~n43188;
  assign n43190 = pi1148 & n43189;
  assign n43191 = pi1091 & n43190;
  assign n43192 = pi1150 & ~n41783;
  assign n43193 = ~pi1149 & ~n43192;
  assign n43194 = ~pi1148 & ~n43193;
  assign n43195 = ~pi1150 & ~n43004;
  assign n43196 = pi1149 & ~n42999;
  assign n43197 = ~n43186 & ~n43196;
  assign n43198 = ~n43195 & ~n43197;
  assign n43199 = n43194 & ~n43198;
  assign n43200 = pi1091 & n43199;
  assign n43201 = ~pi283 & ~n43200;
  assign n43202 = ~n43191 & n43201;
  assign n43203 = ~pi272 & ~n43202;
  assign n43204 = ~n43180 & n43203;
  assign n43205 = pi1150 & n42922;
  assign n43206 = ~pi1150 & n42884;
  assign n43207 = pi1149 & ~n43206;
  assign n43208 = ~n43205 & n43207;
  assign n43209 = pi1150 & n42918;
  assign n43210 = ~pi1150 & n42878;
  assign n43211 = ~pi1149 & ~n43210;
  assign n43212 = ~n43209 & n43211;
  assign n43213 = ~n43208 & ~n43212;
  assign n43214 = pi1148 & ~n43213;
  assign n43215 = pi1150 & n42967;
  assign n43216 = ~pi1150 & ~n42975;
  assign n43217 = ~pi1149 & ~n43216;
  assign n43218 = ~n43215 & n43217;
  assign n43219 = pi1150 & n42963;
  assign n43220 = ~pi1150 & n42973;
  assign n43221 = pi1149 & ~n43220;
  assign n43222 = ~n43219 & n43221;
  assign n43223 = ~n43218 & ~n43222;
  assign n43224 = ~pi1148 & ~n43223;
  assign n43225 = pi283 & ~n43224;
  assign n43226 = ~n43214 & n43225;
  assign n43227 = pi1091 & n43202;
  assign n43228 = pi272 & ~n43227;
  assign n43229 = ~n43226 & n43228;
  assign n43230 = ~pi230 & ~n43229;
  assign n43231 = ~n43204 & n43230;
  assign n43232 = pi230 & ~n43190;
  assign n43233 = ~n43199 & n43232;
  assign po429 = ~n43231 & ~n43233;
  assign n43235 = ~pi273 & ~n40393;
  assign n43236 = ~n40366 & ~n43235;
  assign n43237 = pi219 & ~n43236;
  assign n43238 = ~pi273 & ~n40375;
  assign n43239 = n40377 & ~n43238;
  assign n43240 = ~pi219 & ~n43119;
  assign n43241 = ~n43239 & n43240;
  assign n43242 = ~n43237 & ~n43241;
  assign n43243 = pi299 & n43242;
  assign n43244 = ~pi200 & n43115;
  assign n43245 = ~pi199 & ~n43244;
  assign n43246 = ~n43239 & n43245;
  assign n43247 = pi199 & ~n43236;
  assign n43248 = ~pi299 & ~n43247;
  assign n43249 = ~n43246 & n43248;
  assign n43250 = ~n43243 & ~n43249;
  assign n43251 = ~n11384 & ~n40528;
  assign n43252 = pi1091 & ~n43251;
  assign n43253 = n43250 & ~n43252;
  assign n43254 = ~po1038 & ~n43253;
  assign n43255 = pi1091 & n41892;
  assign n43256 = ~n43254 & ~n43255;
  assign n43257 = pi1147 & ~n43256;
  assign n43258 = po1038 & n43242;
  assign n43259 = n39902 & ~n43250;
  assign n43260 = ~pi1148 & ~n43259;
  assign n43261 = ~n41937 & ~n43242;
  assign n43262 = pi299 & ~n43261;
  assign n43263 = n40574 & ~n43132;
  assign n43264 = ~n43249 & ~n43263;
  assign n43265 = ~n43262 & n43264;
  assign n43266 = ~po1038 & ~n43265;
  assign n43267 = n41781 & n41847;
  assign n43268 = pi1148 & ~n43267;
  assign n43269 = ~n43266 & n43268;
  assign n43270 = ~n43260 & ~n43269;
  assign n43271 = ~n43258 & ~n43270;
  assign n43272 = ~n43257 & n43271;
  assign n43273 = ~pi230 & ~n43272;
  assign n43274 = ~pi1146 & n10670;
  assign n43275 = pi1147 & n39727;
  assign n43276 = ~n42988 & ~n43275;
  assign n43277 = ~n43274 & ~n43276;
  assign n43278 = ~pi1146 & n10758;
  assign n43279 = ~pi199 & pi1147;
  assign n43280 = pi200 & ~n43279;
  assign n43281 = ~n43278 & ~n43280;
  assign n43282 = n16361 & n43281;
  assign n43283 = pi1148 & ~n43282;
  assign n43284 = ~n43277 & n43283;
  assign n43285 = ~pi211 & ~n39797;
  assign n43286 = n39727 & ~n43285;
  assign n43287 = n42986 & ~n43278;
  assign n43288 = ~n43286 & ~n43287;
  assign n43289 = pi1147 & ~n43288;
  assign n43290 = pi1146 & ~n40884;
  assign n43291 = ~n43182 & n43290;
  assign n43292 = ~pi1148 & ~n43291;
  assign n43293 = ~n43289 & n43292;
  assign n43294 = pi230 & ~n43293;
  assign n43295 = ~n43284 & n43294;
  assign po430 = n43273 | n43295;
  assign n43297 = pi274 & ~n40371;
  assign n43298 = ~pi659 & n40371;
  assign n43299 = ~pi1091 & ~n43298;
  assign n43300 = ~n43297 & n43299;
  assign n43301 = ~n42535 & ~n43300;
  assign n43302 = ~pi211 & ~n43301;
  assign n43303 = ~n42578 & ~n43300;
  assign n43304 = pi211 & ~n43303;
  assign n43305 = ~pi219 & ~n43304;
  assign n43306 = ~n43302 & n43305;
  assign n43307 = pi274 & ~n40360;
  assign n43308 = ~pi659 & n40360;
  assign n43309 = ~pi1091 & ~n43308;
  assign n43310 = ~n43307 & n43309;
  assign n43311 = pi219 & ~n43121;
  assign n43312 = ~n43310 & n43311;
  assign n43313 = ~n16361 & ~n43312;
  assign n43314 = ~n43306 & n43313;
  assign n43315 = ~pi200 & ~n43301;
  assign n43316 = pi200 & ~n43303;
  assign n43317 = ~pi199 & ~n43316;
  assign n43318 = ~n43315 & n43317;
  assign n43319 = ~pi200 & n43133;
  assign n43320 = pi199 & ~n43319;
  assign n43321 = ~n43310 & n43320;
  assign n43322 = n16361 & ~n43321;
  assign n43323 = ~n43318 & n43322;
  assign n43324 = ~pi230 & ~n43323;
  assign n43325 = ~n43314 & n43324;
  assign n43326 = ~pi219 & ~n38147;
  assign n43327 = ~n38995 & n43326;
  assign n43328 = ~n39782 & ~n43327;
  assign n43329 = ~n38230 & ~n39785;
  assign n43330 = ~n43327 & ~n43329;
  assign n43331 = ~n38158 & n39890;
  assign n43332 = n40279 & ~n43331;
  assign n43333 = ~n43330 & ~n43332;
  assign n43334 = ~po1038 & ~n43333;
  assign n43335 = pi230 & ~n43334;
  assign n43336 = ~n43328 & n43335;
  assign po431 = ~n43325 & ~n43336;
  assign n43338 = ~pi1151 & n43004;
  assign n43339 = pi1150 & ~n43338;
  assign n43340 = ~n43000 & n43339;
  assign n43341 = n40256 & ~n41783;
  assign n43342 = ~pi1149 & ~n43341;
  assign n43343 = ~n43340 & n43342;
  assign n43344 = pi1151 & ~n42990;
  assign n43345 = pi1149 & n42987;
  assign n43346 = ~n43344 & n43345;
  assign n43347 = n42990 & n43186;
  assign n43348 = ~n43346 & ~n43347;
  assign n43349 = ~n43343 & n43348;
  assign n43350 = pi1091 & ~n43349;
  assign n43351 = pi275 & n43350;
  assign n43352 = pi1091 & n43349;
  assign n43353 = ~pi275 & ~n43352;
  assign n43354 = ~n40646 & ~n43353;
  assign n43355 = ~n43351 & n43354;
  assign n43356 = pi1151 & ~n42918;
  assign n43357 = ~pi1150 & ~n42879;
  assign n43358 = ~n43356 & n43357;
  assign n43359 = pi1150 & n42884;
  assign n43360 = ~n42923 & n43359;
  assign n43361 = pi275 & ~n43360;
  assign n43362 = ~n43358 & n43361;
  assign n43363 = ~pi1150 & ~n42928;
  assign n43364 = pi1151 & ~n43159;
  assign n43365 = ~n43363 & n43364;
  assign n43366 = pi1150 & ~n42906;
  assign n43367 = ~pi1151 & ~n43366;
  assign n43368 = ~n43164 & n43367;
  assign n43369 = ~pi275 & ~n43368;
  assign n43370 = ~n43365 & n43369;
  assign n43371 = pi1149 & ~n43370;
  assign n43372 = ~n43362 & n43371;
  assign n43373 = ~pi1150 & n42946;
  assign n43374 = pi1151 & ~n43170;
  assign n43375 = ~n43373 & n43374;
  assign n43376 = pi1150 & ~n42951;
  assign n43377 = ~pi1151 & ~n43174;
  assign n43378 = ~n43376 & n43377;
  assign n43379 = ~n43375 & ~n43378;
  assign n43380 = ~pi275 & ~n43379;
  assign n43381 = ~pi1150 & n42967;
  assign n43382 = ~n43219 & ~n43381;
  assign n43383 = pi1151 & ~n43382;
  assign n43384 = pi1150 & n42973;
  assign n43385 = ~n43216 & ~n43384;
  assign n43386 = ~pi1151 & ~n43385;
  assign n43387 = pi275 & ~n43386;
  assign n43388 = ~n43383 & n43387;
  assign n43389 = ~pi1149 & ~n43388;
  assign n43390 = ~n43380 & n43389;
  assign n43391 = n40646 & ~n43390;
  assign n43392 = ~n43372 & n43391;
  assign n43393 = ~n43355 & ~n43392;
  assign n43394 = ~pi230 & ~n43393;
  assign n43395 = pi230 & n43349;
  assign po432 = n43394 | n43395;
  assign n43397 = ~pi276 & ~n40361;
  assign n43398 = n40363 & ~n43397;
  assign n43399 = n43057 & ~n43119;
  assign n43400 = pi199 & ~n43244;
  assign n43401 = n16361 & n43400;
  assign n43402 = ~n43399 & ~n43401;
  assign n43403 = ~n43398 & ~n43402;
  assign n43404 = ~pi1091 & ~n40373;
  assign n43405 = ~pi276 & ~n40372;
  assign n43406 = n43404 & ~n43405;
  assign n43407 = ~n38141 & ~n39771;
  assign n43408 = pi1091 & ~n43407;
  assign n43409 = n39727 & ~n43408;
  assign n43410 = pi1145 & n40587;
  assign n43411 = ~n42579 & ~n43410;
  assign n43412 = n42986 & n43411;
  assign n43413 = ~n43409 & ~n43412;
  assign n43414 = ~n43406 & ~n43413;
  assign n43415 = ~pi230 & ~n43414;
  assign n43416 = ~n43403 & n43415;
  assign n43417 = ~pi219 & ~n43407;
  assign n43418 = pi1146 & n38241;
  assign n43419 = ~n43417 & ~n43418;
  assign n43420 = ~n16361 & n43419;
  assign n43421 = ~n38156 & n40769;
  assign n43422 = ~n39893 & ~n43421;
  assign n43423 = n16361 & ~n43422;
  assign n43424 = pi230 & ~n43423;
  assign n43425 = ~n43420 & n43424;
  assign po433 = n43416 | n43425;
  assign n43427 = pi277 & ~n40371;
  assign n43428 = ~pi820 & n40371;
  assign n43429 = ~pi1091 & ~n43428;
  assign n43430 = ~n43427 & n43429;
  assign n43431 = ~n42526 & ~n43430;
  assign n43432 = pi200 & ~n43431;
  assign n43433 = ~n43077 & ~n43430;
  assign n43434 = ~pi200 & ~n43433;
  assign n43435 = ~pi199 & ~n43434;
  assign n43436 = ~n43432 & n43435;
  assign n43437 = pi277 & ~n40360;
  assign n43438 = ~pi820 & n40360;
  assign n43439 = ~pi1091 & ~n43438;
  assign n43440 = ~n43437 & n43439;
  assign n43441 = ~pi200 & n42523;
  assign n43442 = pi199 & ~n43441;
  assign n43443 = ~n43440 & n43442;
  assign n43444 = n16361 & ~n43443;
  assign n43445 = ~n43436 & n43444;
  assign n43446 = pi211 & ~n43431;
  assign n43447 = ~pi211 & ~n43433;
  assign n43448 = ~pi219 & ~n43447;
  assign n43449 = ~n43446 & n43448;
  assign n43450 = pi219 & ~n42597;
  assign n43451 = ~n42545 & ~n43450;
  assign n43452 = ~n43440 & ~n43451;
  assign n43453 = ~n16361 & ~n43452;
  assign n43454 = ~n43449 & n43453;
  assign n43455 = ~n43445 & ~n43454;
  assign n43456 = ~pi230 & ~n43455;
  assign n43457 = n38155 & ~n43097;
  assign n43458 = pi200 & ~n42552;
  assign n43459 = ~n43457 & ~n43458;
  assign n43460 = n16361 & ~n43459;
  assign n43461 = ~pi211 & pi1140;
  assign n43462 = pi211 & pi1141;
  assign n43463 = ~pi219 & ~n43462;
  assign n43464 = ~n43461 & n43463;
  assign n43465 = ~n43450 & ~n43464;
  assign n43466 = ~n16361 & ~n43465;
  assign n43467 = pi230 & ~n43466;
  assign n43468 = ~n43460 & n43467;
  assign po434 = n43456 | n43468;
  assign n43470 = ~pi976 & n40360;
  assign n43471 = ~pi278 & ~n40360;
  assign n43472 = ~pi1091 & ~n43471;
  assign n43473 = ~n43470 & n43472;
  assign n43474 = pi199 & ~n43473;
  assign n43475 = pi1091 & ~pi1132;
  assign n43476 = pi278 & ~n40371;
  assign n43477 = pi976 & n40371;
  assign n43478 = ~pi1091 & ~n43477;
  assign n43479 = ~n43476 & n43478;
  assign n43480 = ~n43475 & ~n43479;
  assign n43481 = ~pi199 & ~n43480;
  assign n43482 = ~n43474 & ~n43481;
  assign n43483 = ~pi200 & ~n43482;
  assign n43484 = pi1091 & ~pi1133;
  assign n43485 = ~n43479 & ~n43484;
  assign n43486 = ~pi199 & ~n43485;
  assign n43487 = ~n43474 & ~n43486;
  assign n43488 = pi200 & ~n43487;
  assign n43489 = ~pi299 & ~n43488;
  assign n43490 = ~n43483 & n43489;
  assign n43491 = pi219 & ~n43473;
  assign n43492 = pi211 & ~pi1133;
  assign n43493 = ~pi211 & ~pi1132;
  assign n43494 = ~n43492 & ~n43493;
  assign n43495 = pi1091 & ~n43494;
  assign n43496 = ~n43479 & ~n43495;
  assign n43497 = ~pi219 & ~n43496;
  assign n43498 = ~n43491 & ~n43497;
  assign n43499 = pi299 & n43498;
  assign n43500 = ~n43490 & ~n43499;
  assign n43501 = ~po1038 & ~n43500;
  assign n43502 = po1038 & n43498;
  assign n43503 = ~pi230 & ~n43502;
  assign n43504 = ~n43501 & n43503;
  assign n43505 = ~pi199 & pi1132;
  assign n43506 = ~pi200 & ~n43505;
  assign n43507 = ~pi199 & pi1133;
  assign n43508 = pi200 & ~n43507;
  assign n43509 = ~pi299 & ~n43508;
  assign n43510 = ~n43506 & n43509;
  assign n43511 = n38230 & n43494;
  assign n43512 = ~n43510 & ~n43511;
  assign n43513 = ~po1038 & ~n43512;
  assign n43514 = n39031 & n43494;
  assign n43515 = pi230 & ~n43514;
  assign n43516 = ~n43513 & n43515;
  assign n43517 = ~n43504 & ~n43516;
  assign n43518 = ~pi1134 & ~n43517;
  assign n43519 = n10758 & ~n43505;
  assign n43520 = n43509 & ~n43519;
  assign n43521 = ~n42011 & ~n43511;
  assign n43522 = ~n43520 & n43521;
  assign n43523 = ~po1038 & ~n43522;
  assign n43524 = pi230 & ~n43523;
  assign n43525 = ~n41782 & ~n43514;
  assign n43526 = n43524 & n43525;
  assign n43527 = ~n40573 & n43483;
  assign n43528 = n43489 & ~n43527;
  assign n43529 = n12979 & n41997;
  assign n43530 = ~n43499 & ~n43529;
  assign n43531 = ~n43528 & n43530;
  assign n43532 = ~po1038 & ~n43531;
  assign n43533 = ~n43267 & n43503;
  assign n43534 = ~n43532 & n43533;
  assign n43535 = ~n43526 & ~n43534;
  assign n43536 = pi1134 & ~n43535;
  assign po435 = ~n43518 & ~n43536;
  assign n43538 = ~pi958 & n40360;
  assign n43539 = ~pi279 & ~n40360;
  assign n43540 = ~pi1091 & ~n43539;
  assign n43541 = ~n43538 & n43540;
  assign n43542 = pi1135 & n43059;
  assign n43543 = ~n43541 & ~n43542;
  assign n43544 = pi199 & ~n43543;
  assign n43545 = pi279 & ~n40371;
  assign n43546 = pi958 & n40371;
  assign n43547 = ~pi1091 & ~n43546;
  assign n43548 = ~n43545 & n43547;
  assign n43549 = ~pi1133 & n43059;
  assign n43550 = ~pi199 & ~n43549;
  assign n43551 = ~n43548 & n43550;
  assign n43552 = ~n43544 & ~n43551;
  assign n43553 = n16361 & ~n43552;
  assign n43554 = ~n40587 & n43553;
  assign n43555 = ~n41949 & ~n43484;
  assign n43556 = ~n43548 & n43555;
  assign n43557 = ~pi219 & ~n43556;
  assign n43558 = pi1135 & n41997;
  assign n43559 = pi219 & ~n43558;
  assign n43560 = ~n43541 & n43559;
  assign n43561 = ~n16361 & ~n43560;
  assign n43562 = ~n43557 & n43561;
  assign n43563 = ~pi230 & ~n43562;
  assign n43564 = ~n43554 & n43563;
  assign n43565 = pi199 & pi1135;
  assign n43566 = ~n43507 & ~n43565;
  assign n43567 = n38270 & ~n43566;
  assign n43568 = pi1135 & n38241;
  assign n43569 = ~pi211 & ~pi1133;
  assign n43570 = ~pi219 & ~n43569;
  assign n43571 = ~pi211 & n43570;
  assign n43572 = ~n43568 & ~n43571;
  assign n43573 = pi299 & ~n43572;
  assign n43574 = ~n43567 & ~n43573;
  assign n43575 = ~po1038 & ~n43574;
  assign n43576 = po1038 & ~n43572;
  assign n43577 = pi230 & ~n43576;
  assign n43578 = ~n43575 & n43577;
  assign n43579 = ~n43564 & ~n43578;
  assign n43580 = ~pi1134 & ~n43579;
  assign n43581 = ~pi1133 & n10758;
  assign n43582 = ~pi200 & pi1135;
  assign n43583 = pi199 & ~n43582;
  assign n43584 = ~n43581 & ~n43583;
  assign n43585 = n16361 & ~n43584;
  assign n43586 = ~n43568 & ~n43570;
  assign n43587 = ~n16361 & n43586;
  assign n43588 = ~n43585 & ~n43587;
  assign n43589 = pi230 & ~n43588;
  assign n43590 = pi1091 & ~n43569;
  assign n43591 = n39727 & n43590;
  assign n43592 = ~n43553 & ~n43591;
  assign n43593 = n43563 & n43592;
  assign n43594 = ~n43589 & ~n43593;
  assign n43595 = pi1134 & ~n43594;
  assign po436 = ~n43580 & ~n43595;
  assign n43597 = ~pi211 & pi1135;
  assign n43598 = pi211 & pi1136;
  assign n43599 = ~n43597 & ~n43598;
  assign n43600 = pi1091 & n43599;
  assign n43601 = pi914 & n40371;
  assign n43602 = ~pi280 & ~n40371;
  assign n43603 = ~pi1091 & ~n43602;
  assign n43604 = ~n43601 & n43603;
  assign n43605 = ~n43600 & ~n43604;
  assign n43606 = ~pi219 & ~n43605;
  assign n43607 = ~pi211 & pi1137;
  assign n43608 = pi219 & ~n43607;
  assign n43609 = ~n42545 & ~n43608;
  assign n43610 = pi280 & ~n40360;
  assign n43611 = ~pi914 & n40360;
  assign n43612 = ~pi1091 & ~n43611;
  assign n43613 = ~n43610 & n43612;
  assign n43614 = ~n43609 & ~n43613;
  assign n43615 = ~n43606 & ~n43614;
  assign n43616 = ~n16361 & ~n43615;
  assign n43617 = pi200 & pi1136;
  assign n43618 = pi1091 & ~n43582;
  assign n43619 = ~n43617 & n43618;
  assign n43620 = ~pi199 & ~n43619;
  assign n43621 = ~n43604 & n43620;
  assign n43622 = pi1137 & n43059;
  assign n43623 = ~n43613 & ~n43622;
  assign n43624 = pi199 & ~n43623;
  assign n43625 = n16361 & ~n43624;
  assign n43626 = ~n43621 & n43625;
  assign n43627 = ~n43616 & ~n43626;
  assign n43628 = ~pi230 & ~n43627;
  assign n43629 = ~pi219 & n43599;
  assign n43630 = ~n43608 & ~n43629;
  assign n43631 = ~n16361 & n43630;
  assign n43632 = pi200 & ~n43025;
  assign n43633 = pi199 & pi1137;
  assign n43634 = ~pi200 & ~n42613;
  assign n43635 = ~n43633 & n43634;
  assign n43636 = ~n43632 & ~n43635;
  assign n43637 = n16361 & n43636;
  assign n43638 = pi230 & ~n43637;
  assign n43639 = ~n43631 & n43638;
  assign po437 = ~n43628 & ~n43639;
  assign n43641 = ~pi199 & pi1138;
  assign n43642 = pi200 & ~n43641;
  assign n43643 = pi199 & pi1139;
  assign n43644 = ~pi200 & ~n43023;
  assign n43645 = ~n43643 & n43644;
  assign n43646 = ~n43642 & ~n43645;
  assign n43647 = n16361 & ~n43646;
  assign n43648 = pi219 & n43072;
  assign n43649 = pi211 & pi1138;
  assign n43650 = ~n43607 & ~n43649;
  assign n43651 = ~pi219 & ~n43650;
  assign n43652 = ~n43648 & ~n43651;
  assign n43653 = ~n16361 & n43652;
  assign n43654 = ~n43647 & ~n43653;
  assign n43655 = pi230 & ~n43654;
  assign n43656 = pi281 & ~n40371;
  assign n43657 = ~pi830 & n40371;
  assign n43658 = ~pi1091 & ~n43657;
  assign n43659 = ~n43656 & n43658;
  assign n43660 = pi1091 & ~n43650;
  assign n43661 = n39727 & ~n43660;
  assign n43662 = pi1138 & n40587;
  assign n43663 = ~n43622 & ~n43662;
  assign n43664 = n42986 & n43663;
  assign n43665 = ~n43661 & ~n43664;
  assign n43666 = ~n43659 & ~n43665;
  assign n43667 = pi281 & ~n40360;
  assign n43668 = ~pi830 & n40360;
  assign n43669 = ~pi1091 & ~n43668;
  assign n43670 = ~n43667 & n43669;
  assign n43671 = pi1139 & n41997;
  assign n43672 = n43057 & ~n43671;
  assign n43673 = pi199 & ~n43079;
  assign n43674 = n16361 & n43673;
  assign n43675 = ~n43672 & ~n43674;
  assign n43676 = ~n43670 & ~n43675;
  assign n43677 = ~n43666 & ~n43676;
  assign n43678 = ~pi230 & ~n43677;
  assign po438 = ~n43655 & ~n43678;
  assign n43680 = pi200 & ~n43099;
  assign n43681 = pi199 & pi1140;
  assign n43682 = ~pi200 & ~n43641;
  assign n43683 = ~n43681 & n43682;
  assign n43684 = ~n43680 & ~n43683;
  assign n43685 = n16361 & ~n43684;
  assign n43686 = pi219 & n43461;
  assign n43687 = pi211 & pi1139;
  assign n43688 = ~n43031 & ~n43687;
  assign n43689 = ~pi219 & ~n43688;
  assign n43690 = ~n43686 & ~n43689;
  assign n43691 = ~n16361 & n43690;
  assign n43692 = ~n43685 & ~n43691;
  assign n43693 = pi230 & ~n43692;
  assign n43694 = pi282 & ~n40371;
  assign n43695 = ~pi836 & n40371;
  assign n43696 = ~pi1091 & ~n43695;
  assign n43697 = ~n43694 & n43696;
  assign n43698 = pi1091 & ~n43688;
  assign n43699 = n39727 & ~n43698;
  assign n43700 = pi1139 & n40587;
  assign n43701 = ~n43060 & ~n43700;
  assign n43702 = n42986 & n43701;
  assign n43703 = ~n43699 & ~n43702;
  assign n43704 = ~n43697 & ~n43703;
  assign n43705 = pi282 & ~n40360;
  assign n43706 = ~pi836 & n40360;
  assign n43707 = ~pi1091 & ~n43706;
  assign n43708 = ~n43705 & n43707;
  assign n43709 = pi1140 & n41997;
  assign n43710 = n43057 & ~n43709;
  assign n43711 = ~pi200 & n43077;
  assign n43712 = pi199 & ~n43711;
  assign n43713 = n16361 & n43712;
  assign n43714 = ~n43710 & ~n43713;
  assign n43715 = ~n43708 & ~n43714;
  assign n43716 = ~n43704 & ~n43715;
  assign n43717 = ~pi230 & ~n43716;
  assign po439 = ~n43693 & ~n43717;
  assign n43719 = pi1147 & ~n42987;
  assign n43720 = ~pi1149 & n43004;
  assign n43721 = ~n43719 & n43720;
  assign n43722 = pi1147 & ~n43182;
  assign n43723 = n43196 & ~n43722;
  assign n43724 = pi1148 & ~n43723;
  assign n43725 = ~n43721 & n43724;
  assign n43726 = pi1149 & ~n41783;
  assign n43727 = ~n43722 & ~n43726;
  assign n43728 = ~pi1148 & ~n43727;
  assign n43729 = pi230 & ~n43728;
  assign n43730 = ~n43725 & n43729;
  assign n43731 = ~pi1147 & ~n42951;
  assign n43732 = pi1147 & n42906;
  assign n43733 = ~pi1149 & ~n43732;
  assign n43734 = ~n43731 & n43733;
  assign n43735 = ~pi1147 & n42942;
  assign n43736 = pi1147 & n42933;
  assign n43737 = pi1149 & ~n43736;
  assign n43738 = ~n43735 & n43737;
  assign n43739 = pi1148 & ~n43738;
  assign n43740 = ~n43734 & n43739;
  assign n43741 = pi1147 & n42928;
  assign n43742 = ~pi1147 & n42946;
  assign n43743 = pi1149 & ~n43742;
  assign n43744 = ~n43741 & n43743;
  assign n43745 = pi1147 & n42898;
  assign n43746 = ~pi1147 & ~n42905;
  assign n43747 = ~pi1149 & ~n43746;
  assign n43748 = ~n43745 & n43747;
  assign n43749 = ~pi1148 & ~n43748;
  assign n43750 = ~n43744 & n43749;
  assign n43751 = ~pi283 & ~n43750;
  assign n43752 = ~n43740 & n43751;
  assign n43753 = pi1147 & n42918;
  assign n43754 = ~pi1147 & n42967;
  assign n43755 = ~pi1148 & ~n43754;
  assign n43756 = ~n43753 & n43755;
  assign n43757 = ~pi1147 & n42963;
  assign n43758 = pi1147 & n42922;
  assign n43759 = pi1148 & ~n43758;
  assign n43760 = ~n43757 & n43759;
  assign n43761 = pi1149 & ~n43760;
  assign n43762 = ~n43756 & n43761;
  assign n43763 = pi1147 & n42878;
  assign n43764 = ~pi1147 & ~n42975;
  assign n43765 = ~pi1148 & ~n43764;
  assign n43766 = ~n43763 & n43765;
  assign n43767 = ~pi1147 & n42973;
  assign n43768 = pi1147 & n42884;
  assign n43769 = pi1148 & ~n43768;
  assign n43770 = ~n43767 & n43769;
  assign n43771 = ~pi1149 & ~n43770;
  assign n43772 = ~n43766 & n43771;
  assign n43773 = pi283 & ~n43772;
  assign n43774 = ~n43762 & n43773;
  assign n43775 = ~pi230 & ~n43774;
  assign n43776 = ~n43752 & n43775;
  assign po440 = ~n43730 & ~n43776;
  assign n43778 = ~pi284 & ~n42290;
  assign n43779 = pi1143 & n42290;
  assign n43780 = ~n39729 & n43779;
  assign po441 = n43778 | n43780;
  assign n43782 = n3268 & ~n10361;
  assign n43783 = ~n8021 & n43782;
  assign n43784 = pi286 & n43783;
  assign n43785 = pi288 & pi289;
  assign n43786 = n43784 & n43785;
  assign n43787 = pi285 & n43782;
  assign n43788 = ~n43786 & ~n43787;
  assign n43789 = pi285 & n43786;
  assign n43790 = ~po1038 & ~n43789;
  assign n43791 = ~n43788 & n43790;
  assign n43792 = ~po1038 & n43786;
  assign n43793 = ~pi286 & n8021;
  assign n43794 = ~pi288 & n43793;
  assign n43795 = pi285 & ~pi289;
  assign n43796 = n43794 & n43795;
  assign n43797 = pi285 & ~n43796;
  assign n43798 = ~n43792 & n43797;
  assign n43799 = ~n43791 & ~n43798;
  assign po442 = ~pi793 & ~n43799;
  assign n43801 = ~pi286 & ~n43783;
  assign n43802 = pi288 & ~n43784;
  assign n43803 = ~n43801 & n43802;
  assign n43804 = ~pi288 & ~n7696;
  assign n43805 = n8021 & ~n43782;
  assign n43806 = pi286 & ~n43805;
  assign n43807 = ~n43782 & n43793;
  assign n43808 = ~n43806 & ~n43807;
  assign n43809 = n43804 & ~n43808;
  assign n43810 = ~po1038 & ~n43809;
  assign n43811 = ~n43803 & n43810;
  assign n43812 = n8021 & n43804;
  assign n43813 = ~pi286 & n43812;
  assign n43814 = pi286 & ~n43812;
  assign n43815 = po1038 & ~n43814;
  assign n43816 = ~n43813 & n43815;
  assign n43817 = ~pi793 & ~n43816;
  assign po443 = ~n43811 & n43817;
  assign n43819 = ~pi287 & pi457;
  assign po444 = ~pi332 & ~n43819;
  assign n43821 = pi288 & ~n8021;
  assign n43822 = ~n43812 & ~n43821;
  assign po637 = ~po1038 & n43782;
  assign n43824 = n43822 & ~po637;
  assign n43825 = ~n43822 & po637;
  assign n43826 = ~pi793 & ~n43825;
  assign po445 = ~n43824 & n43826;
  assign n43828 = pi289 & ~n43807;
  assign n43829 = n43795 & n43807;
  assign n43830 = ~pi288 & ~n43829;
  assign n43831 = ~n43828 & n43830;
  assign n43832 = ~pi289 & n43802;
  assign n43833 = ~n43786 & ~n43832;
  assign n43834 = ~n43831 & n43833;
  assign n43835 = ~po1038 & ~n43834;
  assign n43836 = pi289 & ~n43794;
  assign n43837 = po1038 & ~n43836;
  assign n43838 = ~n43796 & n43837;
  assign n43839 = ~pi793 & ~n43838;
  assign po446 = ~n43835 & n43839;
  assign n43841 = ~pi290 & pi476;
  assign n43842 = ~pi476 & ~pi1048;
  assign po447 = ~n43841 & ~n43842;
  assign n43844 = ~pi291 & pi476;
  assign n43845 = ~pi476 & ~pi1049;
  assign po448 = ~n43844 & ~n43845;
  assign n43847 = ~pi292 & pi476;
  assign n43848 = ~pi476 & ~pi1084;
  assign po449 = ~n43847 & ~n43848;
  assign n43850 = ~pi293 & pi476;
  assign n43851 = ~pi476 & ~pi1059;
  assign po450 = ~n43850 & ~n43851;
  assign n43853 = ~pi294 & pi476;
  assign n43854 = ~pi476 & ~pi1072;
  assign po451 = ~n43853 & ~n43854;
  assign n43856 = ~pi295 & pi476;
  assign n43857 = ~pi476 & ~pi1053;
  assign po452 = ~n43856 & ~n43857;
  assign n43859 = ~pi296 & pi476;
  assign n43860 = ~pi476 & ~pi1037;
  assign po453 = ~n43859 & ~n43860;
  assign n43862 = ~pi297 & pi476;
  assign n43863 = ~pi476 & ~pi1044;
  assign po454 = ~n43862 & ~n43863;
  assign n43865 = ~pi478 & pi1044;
  assign n43866 = pi298 & pi478;
  assign po455 = n43865 | n43866;
  assign n43868 = pi54 & n3095;
  assign n43869 = ~pi54 & n13069;
  assign n43870 = n13327 & n43869;
  assign n43871 = ~n43868 & ~n43870;
  assign n43872 = n3242 & n8840;
  assign n43873 = ~n43871 & n43872;
  assign n43874 = ~pi39 & ~n43873;
  assign po456 = ~n11209 & ~n43874;
  assign n43876 = pi57 & ~pi59;
  assign n43877 = n10088 & n43876;
  assign n43878 = ~pi312 & n43877;
  assign n43879 = pi300 & ~n43878;
  assign n43880 = ~pi300 & n43878;
  assign n43881 = ~pi55 & ~n43880;
  assign po457 = n43879 | ~n43881;
  assign n43883 = ~pi301 & n43881;
  assign n43884 = ~pi55 & pi301;
  assign n43885 = n43880 & n43884;
  assign po458 = n43883 | n43885;
  assign n43887 = n5777 & ~po1038;
  assign n43888 = n5788 & ~n16361;
  assign n43889 = ~n43887 & ~n43888;
  assign n43890 = ~pi1148 & n43889;
  assign n43891 = ~pi222 & ~pi223;
  assign n43892 = pi937 & ~n43891;
  assign n43893 = pi273 & n3306;
  assign n43894 = ~n43892 & ~n43893;
  assign n43895 = n43887 & n43894;
  assign n43896 = n3330 & ~n16361;
  assign n43897 = ~n43895 & ~n43896;
  assign n43898 = pi237 & ~n43897;
  assign n43899 = ~n3052 & n43895;
  assign n43900 = ~pi215 & n3324;
  assign n43901 = ~pi273 & n43900;
  assign n43902 = pi833 & n8039;
  assign n43903 = ~pi937 & n43902;
  assign n43904 = ~n43901 & ~n43903;
  assign n43905 = ~n16361 & ~n43904;
  assign n43906 = ~n43899 & ~n43905;
  assign n43907 = ~n43898 & n43906;
  assign po459 = ~n43890 & n43907;
  assign n43909 = ~pi478 & pi1049;
  assign n43910 = pi303 & pi478;
  assign po460 = n43909 | n43910;
  assign n43912 = ~pi478 & pi1048;
  assign n43913 = pi304 & pi478;
  assign po461 = n43912 | n43913;
  assign n43915 = ~pi478 & pi1084;
  assign n43916 = pi305 & pi478;
  assign po462 = n43915 | n43916;
  assign n43918 = ~pi478 & pi1059;
  assign n43919 = pi306 & pi478;
  assign po463 = n43918 | n43919;
  assign n43921 = ~pi478 & pi1053;
  assign n43922 = pi307 & pi478;
  assign po464 = n43921 | n43922;
  assign n43924 = ~pi478 & pi1037;
  assign n43925 = pi308 & pi478;
  assign po465 = n43924 | n43925;
  assign n43927 = ~pi478 & pi1072;
  assign n43928 = pi309 & pi478;
  assign po466 = n43927 | n43928;
  assign n43930 = pi1147 & n43889;
  assign n43931 = pi222 & ~pi934;
  assign n43932 = ~pi271 & n3306;
  assign n43933 = ~n43931 & ~n43932;
  assign n43934 = n43887 & n43933;
  assign n43935 = ~n43896 & ~n43934;
  assign n43936 = pi934 & ~n3136;
  assign n43937 = pi271 & n3324;
  assign n43938 = ~n43936 & ~n43937;
  assign n43939 = n43888 & ~n43938;
  assign n43940 = n43935 & ~n43939;
  assign n43941 = ~n43930 & n43940;
  assign n43942 = ~pi233 & ~n43941;
  assign n43943 = n43888 & n43938;
  assign n43944 = n43887 & ~n43933;
  assign n43945 = n3100 & n16361;
  assign n43946 = pi1147 & ~n43945;
  assign n43947 = ~n43944 & n43946;
  assign n43948 = ~n43943 & n43947;
  assign n43949 = ~n43896 & ~n43945;
  assign n43950 = ~n43889 & n43949;
  assign n43951 = ~pi1147 & n43950;
  assign n43952 = ~n43940 & n43951;
  assign n43953 = ~n43948 & ~n43952;
  assign n43954 = pi233 & ~n43953;
  assign po467 = n43942 | n43954;
  assign n43956 = ~pi55 & ~pi311;
  assign n43957 = ~n43885 & ~n43956;
  assign n43958 = ~pi311 & n43885;
  assign po468 = ~n43957 & ~n43958;
  assign n43960 = pi312 & ~n43877;
  assign n43961 = ~n43878 & ~n43960;
  assign po469 = ~pi55 & ~n43961;
  assign n43963 = ~n10350 & ~n13360;
  assign n43964 = po740 & ~n13367;
  assign n43965 = n10112 & ~n43964;
  assign po634 = n43963 | ~n43965;
  assign n43967 = ~pi954 & po634;
  assign n43968 = pi313 & pi954;
  assign po470 = ~n43967 & ~n43968;
  assign n43970 = n6536 & n8840;
  assign n43971 = n14354 & ~n43970;
  assign n43972 = ~pi39 & ~n14423;
  assign n43973 = pi39 & ~n15186;
  assign n43974 = n3206 & ~n43973;
  assign n43975 = ~n43972 & n43974;
  assign n43976 = ~n15480 & ~n43975;
  assign n43977 = n3277 & n10109;
  assign n43978 = ~n43976 & n43977;
  assign n43979 = ~n43971 & ~n43978;
  assign n43980 = n14348 & n14349;
  assign po471 = ~n43979 & n43980;
  assign n43982 = ~pi340 & n43782;
  assign n43983 = ~po1038 & n43982;
  assign n43984 = pi315 & ~n43983;
  assign n43985 = pi1080 & n43983;
  assign po472 = n43984 | n43985;
  assign n43987 = pi316 & ~n43983;
  assign n43988 = pi1047 & n43983;
  assign po473 = n43987 | n43988;
  assign n43990 = ~pi330 & po637;
  assign n43991 = pi317 & ~n43990;
  assign n43992 = pi1078 & n43990;
  assign po474 = n43991 | n43992;
  assign n43994 = ~pi341 & n43782;
  assign n43995 = ~po1038 & n43994;
  assign n43996 = pi318 & ~n43995;
  assign n43997 = pi1074 & n43995;
  assign po475 = n43996 | n43997;
  assign n43999 = pi319 & ~n43995;
  assign n44000 = pi1072 & n43995;
  assign po476 = n43999 | n44000;
  assign n44002 = pi320 & ~n43983;
  assign n44003 = pi1048 & n43983;
  assign po477 = n44002 | n44003;
  assign n44005 = pi321 & ~n43983;
  assign n44006 = pi1058 & n43983;
  assign po478 = n44005 | n44006;
  assign n44008 = pi322 & ~n43983;
  assign n44009 = pi1051 & n43983;
  assign po479 = n44008 | n44009;
  assign n44011 = pi323 & ~n43983;
  assign n44012 = pi1065 & n43983;
  assign po480 = n44011 | n44012;
  assign n44014 = pi324 & ~n43995;
  assign n44015 = pi1086 & n43995;
  assign po481 = n44014 | n44015;
  assign n44017 = pi325 & ~n43995;
  assign n44018 = pi1063 & n43995;
  assign po482 = n44017 | n44018;
  assign n44020 = pi326 & ~n43995;
  assign n44021 = pi1057 & n43995;
  assign po483 = n44020 | n44021;
  assign n44023 = pi327 & ~n43983;
  assign n44024 = pi1040 & n43983;
  assign po484 = n44023 | n44024;
  assign n44026 = pi328 & ~n43995;
  assign n44027 = pi1058 & n43995;
  assign po485 = n44026 | n44027;
  assign n44029 = pi329 & ~n43995;
  assign n44030 = pi1043 & n43995;
  assign po486 = n44029 | n44030;
  assign n44032 = pi1092 & ~n10018;
  assign n44033 = po1038 & n44032;
  assign n44034 = ~pi330 & n44033;
  assign n44035 = ~po1038 & n44032;
  assign n44036 = ~pi330 & ~n43782;
  assign n44037 = ~n43982 & ~n44036;
  assign n44038 = n44035 & ~n44037;
  assign po487 = n44034 | n44038;
  assign n44040 = ~pi331 & n44033;
  assign n44041 = ~pi331 & ~n43782;
  assign n44042 = ~n43994 & ~n44041;
  assign n44043 = n44035 & ~n44042;
  assign po488 = n44040 | n44043;
  assign n44045 = n10942 & n13090;
  assign n44046 = ~n10942 & ~n13020;
  assign n44047 = n7437 & ~n44046;
  assign n44048 = ~pi70 & ~n44047;
  assign n44049 = pi332 & n9512;
  assign n44050 = ~n44048 & n44049;
  assign n44051 = ~n44045 & ~n44050;
  assign n44052 = ~pi39 & ~n44051;
  assign n44053 = pi39 & n10376;
  assign n44054 = ~pi38 & ~n44053;
  assign n44055 = ~n44052 & n44054;
  assign po489 = n37991 & ~n44055;
  assign n44057 = pi333 & ~n43995;
  assign n44058 = pi1040 & n43995;
  assign po490 = n44057 | n44058;
  assign n44060 = pi334 & ~n43995;
  assign n44061 = pi1065 & n43995;
  assign po491 = n44060 | n44061;
  assign n44063 = pi335 & ~n43995;
  assign n44064 = pi1069 & n43995;
  assign po492 = n44063 | n44064;
  assign n44066 = pi336 & ~n43990;
  assign n44067 = pi1070 & n43990;
  assign po493 = n44066 | n44067;
  assign n44069 = pi337 & ~n43990;
  assign n44070 = pi1044 & n43990;
  assign po494 = n44069 | n44070;
  assign n44072 = pi338 & ~n43990;
  assign n44073 = pi1072 & n43990;
  assign po495 = n44072 | n44073;
  assign n44075 = pi339 & ~n43990;
  assign n44076 = pi1086 & n43990;
  assign po496 = n44075 | n44076;
  assign n44078 = pi340 & n44033;
  assign n44079 = ~pi331 & n43782;
  assign n44080 = ~pi340 & ~n43782;
  assign n44081 = n44035 & ~n44080;
  assign n44082 = ~n44079 & n44081;
  assign po497 = ~n44078 & ~n44082;
  assign n44084 = ~pi341 & ~po637;
  assign n44085 = ~n43990 & ~n44084;
  assign po498 = n44032 & ~n44085;
  assign n44087 = pi342 & ~n43983;
  assign n44088 = pi1049 & n43983;
  assign po499 = n44087 | n44088;
  assign n44090 = pi343 & ~n43983;
  assign n44091 = pi1062 & n43983;
  assign po500 = n44090 | n44091;
  assign n44093 = pi344 & ~n43983;
  assign n44094 = pi1069 & n43983;
  assign po501 = n44093 | n44094;
  assign n44096 = pi345 & ~n43983;
  assign n44097 = pi1039 & n43983;
  assign po502 = n44096 | n44097;
  assign n44099 = pi346 & ~n43983;
  assign n44100 = pi1067 & n43983;
  assign po503 = n44099 | n44100;
  assign n44102 = pi347 & ~n43983;
  assign n44103 = pi1055 & n43983;
  assign po504 = n44102 | n44103;
  assign n44105 = pi348 & ~n43983;
  assign n44106 = pi1087 & n43983;
  assign po505 = n44105 | n44106;
  assign n44108 = pi349 & ~n43983;
  assign n44109 = pi1043 & n43983;
  assign po506 = n44108 | n44109;
  assign n44111 = pi350 & ~n43983;
  assign n44112 = pi1035 & n43983;
  assign po507 = n44111 | n44112;
  assign n44114 = pi351 & ~n43983;
  assign n44115 = pi1079 & n43983;
  assign po508 = n44114 | n44115;
  assign n44117 = pi352 & ~n43983;
  assign n44118 = pi1078 & n43983;
  assign po509 = n44117 | n44118;
  assign n44120 = pi353 & ~n43983;
  assign n44121 = pi1063 & n43983;
  assign po510 = n44120 | n44121;
  assign n44123 = pi354 & ~n43983;
  assign n44124 = pi1045 & n43983;
  assign po511 = n44123 | n44124;
  assign n44126 = pi355 & ~n43983;
  assign n44127 = pi1084 & n43983;
  assign po512 = n44126 | n44127;
  assign n44129 = pi356 & ~n43983;
  assign n44130 = pi1081 & n43983;
  assign po513 = n44129 | n44130;
  assign n44132 = pi357 & ~n43983;
  assign n44133 = pi1076 & n43983;
  assign po514 = n44132 | n44133;
  assign n44135 = pi358 & ~n43983;
  assign n44136 = pi1071 & n43983;
  assign po515 = n44135 | n44136;
  assign n44138 = pi359 & ~n43983;
  assign n44139 = pi1068 & n43983;
  assign po516 = n44138 | n44139;
  assign n44141 = pi360 & ~n43983;
  assign n44142 = pi1042 & n43983;
  assign po517 = n44141 | n44142;
  assign n44144 = pi361 & ~n43983;
  assign n44145 = pi1059 & n43983;
  assign po518 = n44144 | n44145;
  assign n44147 = pi362 & ~n43983;
  assign n44148 = pi1070 & n43983;
  assign po519 = n44147 | n44148;
  assign n44150 = pi363 & ~n43990;
  assign n44151 = pi1049 & n43990;
  assign po520 = n44150 | n44151;
  assign n44153 = pi364 & ~n43990;
  assign n44154 = pi1062 & n43990;
  assign po521 = n44153 | n44154;
  assign n44156 = pi365 & ~n43990;
  assign n44157 = pi1065 & n43990;
  assign po522 = n44156 | n44157;
  assign n44159 = pi366 & ~n43990;
  assign n44160 = pi1069 & n43990;
  assign po523 = n44159 | n44160;
  assign n44162 = pi367 & ~n43990;
  assign n44163 = pi1039 & n43990;
  assign po524 = n44162 | n44163;
  assign n44165 = pi368 & ~n43990;
  assign n44166 = pi1067 & n43990;
  assign po525 = n44165 | n44166;
  assign n44168 = pi369 & ~n43990;
  assign n44169 = pi1080 & n43990;
  assign po526 = n44168 | n44169;
  assign n44171 = pi370 & ~n43990;
  assign n44172 = pi1055 & n43990;
  assign po527 = n44171 | n44172;
  assign n44174 = pi371 & ~n43990;
  assign n44175 = pi1051 & n43990;
  assign po528 = n44174 | n44175;
  assign n44177 = pi372 & ~n43990;
  assign n44178 = pi1048 & n43990;
  assign po529 = n44177 | n44178;
  assign n44180 = pi373 & ~n43990;
  assign n44181 = pi1087 & n43990;
  assign po530 = n44180 | n44181;
  assign n44183 = pi374 & ~n43990;
  assign n44184 = pi1035 & n43990;
  assign po531 = n44183 | n44184;
  assign n44186 = pi375 & ~n43990;
  assign n44187 = pi1047 & n43990;
  assign po532 = n44186 | n44187;
  assign n44189 = pi376 & ~n43990;
  assign n44190 = pi1079 & n43990;
  assign po533 = n44189 | n44190;
  assign n44192 = pi377 & ~n43990;
  assign n44193 = pi1074 & n43990;
  assign po534 = n44192 | n44193;
  assign n44195 = pi378 & ~n43990;
  assign n44196 = pi1063 & n43990;
  assign po535 = n44195 | n44196;
  assign n44198 = pi379 & ~n43990;
  assign n44199 = pi1045 & n43990;
  assign po536 = n44198 | n44199;
  assign n44201 = pi380 & ~n43990;
  assign n44202 = pi1084 & n43990;
  assign po537 = n44201 | n44202;
  assign n44204 = pi381 & ~n43990;
  assign n44205 = pi1081 & n43990;
  assign po538 = n44204 | n44205;
  assign n44207 = pi382 & ~n43990;
  assign n44208 = pi1076 & n43990;
  assign po539 = n44207 | n44208;
  assign n44210 = pi383 & ~n43990;
  assign n44211 = pi1071 & n43990;
  assign po540 = n44210 | n44211;
  assign n44213 = pi384 & ~n43990;
  assign n44214 = pi1068 & n43990;
  assign po541 = n44213 | n44214;
  assign n44216 = pi385 & ~n43990;
  assign n44217 = pi1042 & n43990;
  assign po542 = n44216 | n44217;
  assign n44219 = pi386 & ~n43990;
  assign n44220 = pi1059 & n43990;
  assign po543 = n44219 | n44220;
  assign n44222 = pi387 & ~n43990;
  assign n44223 = pi1053 & n43990;
  assign po544 = n44222 | n44223;
  assign n44225 = pi388 & ~n43990;
  assign n44226 = pi1037 & n43990;
  assign po545 = n44225 | n44226;
  assign n44228 = pi389 & ~n43990;
  assign n44229 = pi1036 & n43990;
  assign po546 = n44228 | n44229;
  assign n44231 = pi390 & ~n43995;
  assign n44232 = pi1049 & n43995;
  assign po547 = n44231 | n44232;
  assign n44234 = pi391 & ~n43995;
  assign n44235 = pi1062 & n43995;
  assign po548 = n44234 | n44235;
  assign n44237 = pi392 & ~n43995;
  assign n44238 = pi1039 & n43995;
  assign po549 = n44237 | n44238;
  assign n44240 = pi393 & ~n43995;
  assign n44241 = pi1067 & n43995;
  assign po550 = n44240 | n44241;
  assign n44243 = pi394 & ~n43995;
  assign n44244 = pi1080 & n43995;
  assign po551 = n44243 | n44244;
  assign n44246 = pi395 & ~n43995;
  assign n44247 = pi1055 & n43995;
  assign po552 = n44246 | n44247;
  assign n44249 = pi396 & ~n43995;
  assign n44250 = pi1051 & n43995;
  assign po553 = n44249 | n44250;
  assign n44252 = pi397 & ~n43995;
  assign n44253 = pi1048 & n43995;
  assign po554 = n44252 | n44253;
  assign n44255 = pi398 & ~n43995;
  assign n44256 = pi1087 & n43995;
  assign po555 = n44255 | n44256;
  assign n44258 = pi399 & ~n43995;
  assign n44259 = pi1047 & n43995;
  assign po556 = n44258 | n44259;
  assign n44261 = pi400 & ~n43995;
  assign n44262 = pi1035 & n43995;
  assign po557 = n44261 | n44262;
  assign n44264 = pi401 & ~n43995;
  assign n44265 = pi1079 & n43995;
  assign po558 = n44264 | n44265;
  assign n44267 = pi402 & ~n43995;
  assign n44268 = pi1078 & n43995;
  assign po559 = n44267 | n44268;
  assign n44270 = pi403 & ~n43995;
  assign n44271 = pi1045 & n43995;
  assign po560 = n44270 | n44271;
  assign n44273 = pi404 & ~n43995;
  assign n44274 = pi1084 & n43995;
  assign po561 = n44273 | n44274;
  assign n44276 = pi405 & ~n43995;
  assign n44277 = pi1081 & n43995;
  assign po562 = n44276 | n44277;
  assign n44279 = pi406 & ~n43995;
  assign n44280 = pi1076 & n43995;
  assign po563 = n44279 | n44280;
  assign n44282 = pi407 & ~n43995;
  assign n44283 = pi1071 & n43995;
  assign po564 = n44282 | n44283;
  assign n44285 = pi408 & ~n43995;
  assign n44286 = pi1068 & n43995;
  assign po565 = n44285 | n44286;
  assign n44288 = pi409 & ~n43995;
  assign n44289 = pi1042 & n43995;
  assign po566 = n44288 | n44289;
  assign n44291 = pi410 & ~n43995;
  assign n44292 = pi1059 & n43995;
  assign po567 = n44291 | n44292;
  assign n44294 = pi411 & ~n43995;
  assign n44295 = pi1053 & n43995;
  assign po568 = n44294 | n44295;
  assign n44297 = pi412 & ~n43995;
  assign n44298 = pi1037 & n43995;
  assign po569 = n44297 | n44298;
  assign n44300 = pi413 & ~n43995;
  assign n44301 = pi1036 & n43995;
  assign po570 = n44300 | n44301;
  assign n44303 = ~po1038 & n44079;
  assign n44304 = pi414 & ~n44303;
  assign n44305 = pi1049 & n44303;
  assign po571 = n44304 | n44305;
  assign n44307 = pi415 & ~n44303;
  assign n44308 = pi1062 & n44303;
  assign po572 = n44307 | n44308;
  assign n44310 = pi416 & ~n44303;
  assign n44311 = pi1069 & n44303;
  assign po573 = n44310 | n44311;
  assign n44313 = pi417 & ~n44303;
  assign n44314 = pi1039 & n44303;
  assign po574 = n44313 | n44314;
  assign n44316 = pi418 & ~n44303;
  assign n44317 = pi1067 & n44303;
  assign po575 = n44316 | n44317;
  assign n44319 = pi419 & ~n44303;
  assign n44320 = pi1080 & n44303;
  assign po576 = n44319 | n44320;
  assign n44322 = pi420 & ~n44303;
  assign n44323 = pi1055 & n44303;
  assign po577 = n44322 | n44323;
  assign n44325 = pi421 & ~n44303;
  assign n44326 = pi1051 & n44303;
  assign po578 = n44325 | n44326;
  assign n44328 = pi422 & ~n44303;
  assign n44329 = pi1048 & n44303;
  assign po579 = n44328 | n44329;
  assign n44331 = pi423 & ~n44303;
  assign n44332 = pi1087 & n44303;
  assign po580 = n44331 | n44332;
  assign n44334 = pi424 & ~n44303;
  assign n44335 = pi1047 & n44303;
  assign po581 = n44334 | n44335;
  assign n44337 = pi425 & ~n44303;
  assign n44338 = pi1035 & n44303;
  assign po582 = n44337 | n44338;
  assign n44340 = pi426 & ~n44303;
  assign n44341 = pi1079 & n44303;
  assign po583 = n44340 | n44341;
  assign n44343 = pi427 & ~n44303;
  assign n44344 = pi1078 & n44303;
  assign po584 = n44343 | n44344;
  assign n44346 = pi428 & ~n44303;
  assign n44347 = pi1045 & n44303;
  assign po585 = n44346 | n44347;
  assign n44349 = pi429 & ~n44303;
  assign n44350 = pi1084 & n44303;
  assign po586 = n44349 | n44350;
  assign n44352 = pi430 & ~n44303;
  assign n44353 = pi1076 & n44303;
  assign po587 = n44352 | n44353;
  assign n44355 = pi431 & ~n44303;
  assign n44356 = pi1071 & n44303;
  assign po588 = n44355 | n44356;
  assign n44358 = pi432 & ~n44303;
  assign n44359 = pi1068 & n44303;
  assign po589 = n44358 | n44359;
  assign n44361 = pi433 & ~n44303;
  assign n44362 = pi1042 & n44303;
  assign po590 = n44361 | n44362;
  assign n44364 = pi434 & ~n44303;
  assign n44365 = pi1059 & n44303;
  assign po591 = n44364 | n44365;
  assign n44367 = pi435 & ~n44303;
  assign n44368 = pi1053 & n44303;
  assign po592 = n44367 | n44368;
  assign n44370 = pi436 & ~n44303;
  assign n44371 = pi1037 & n44303;
  assign po593 = n44370 | n44371;
  assign n44373 = pi437 & ~n44303;
  assign n44374 = pi1070 & n44303;
  assign po594 = n44373 | n44374;
  assign n44376 = pi438 & ~n44303;
  assign n44377 = pi1036 & n44303;
  assign po595 = n44376 | n44377;
  assign n44379 = pi439 & ~n43990;
  assign n44380 = pi1057 & n43990;
  assign po596 = n44379 | n44380;
  assign n44382 = pi440 & ~n43990;
  assign n44383 = pi1043 & n43990;
  assign po597 = n44382 | n44383;
  assign n44385 = pi441 & ~n43983;
  assign n44386 = pi1044 & n43983;
  assign po598 = n44385 | n44386;
  assign n44388 = pi442 & ~n43990;
  assign n44389 = pi1058 & n43990;
  assign po599 = n44388 | n44389;
  assign n44391 = pi443 & ~n44303;
  assign n44392 = pi1044 & n44303;
  assign po600 = n44391 | n44392;
  assign n44394 = pi444 & ~n44303;
  assign n44395 = pi1072 & n44303;
  assign po601 = n44394 | n44395;
  assign n44397 = pi445 & ~n44303;
  assign n44398 = pi1081 & n44303;
  assign po602 = n44397 | n44398;
  assign n44400 = pi446 & ~n44303;
  assign n44401 = pi1086 & n44303;
  assign po603 = n44400 | n44401;
  assign n44403 = pi447 & ~n43990;
  assign n44404 = pi1040 & n43990;
  assign po604 = n44403 | n44404;
  assign n44406 = pi448 & ~n44303;
  assign n44407 = pi1074 & n44303;
  assign po605 = n44406 | n44407;
  assign n44409 = pi449 & ~n44303;
  assign n44410 = pi1057 & n44303;
  assign po606 = n44409 | n44410;
  assign n44412 = pi450 & ~n43983;
  assign n44413 = pi1036 & n43983;
  assign po607 = n44412 | n44413;
  assign n44415 = pi451 & ~n44303;
  assign n44416 = pi1063 & n44303;
  assign po608 = n44415 | n44416;
  assign n44418 = pi452 & ~n43983;
  assign n44419 = pi1053 & n43983;
  assign po609 = n44418 | n44419;
  assign n44421 = pi453 & ~n44303;
  assign n44422 = pi1040 & n44303;
  assign po610 = n44421 | n44422;
  assign n44424 = pi454 & ~n44303;
  assign n44425 = pi1043 & n44303;
  assign po611 = n44424 | n44425;
  assign n44427 = pi455 & ~n43983;
  assign n44428 = pi1037 & n43983;
  assign po612 = n44427 | n44428;
  assign n44430 = pi456 & ~n43995;
  assign n44431 = pi1044 & n43995;
  assign po613 = n44430 | n44431;
  assign n44433 = pi594 & pi600;
  assign n44434 = pi597 & n44433;
  assign n44435 = pi601 & n44434;
  assign n44436 = ~pi804 & ~pi810;
  assign n44437 = ~pi595 & n44436;
  assign n44438 = ~pi599 & pi810;
  assign n44439 = pi596 & ~n44438;
  assign n44440 = pi804 & ~n44439;
  assign n44441 = pi595 & pi815;
  assign n44442 = ~n44440 & n44441;
  assign n44443 = ~n44437 & ~n44442;
  assign n44444 = n44435 & ~n44443;
  assign n44445 = ~pi601 & ~n44436;
  assign n44446 = pi600 & ~pi810;
  assign n44447 = pi804 & ~n44446;
  assign n44448 = ~pi815 & ~n44447;
  assign n44449 = ~n44445 & n44448;
  assign n44450 = ~n44444 & ~n44449;
  assign n44451 = pi605 & ~n44450;
  assign n44452 = pi990 & n44433;
  assign n44453 = ~pi815 & n44447;
  assign n44454 = n44452 & n44453;
  assign n44455 = ~n44451 & ~n44454;
  assign po614 = pi821 & ~n44455;
  assign n44457 = pi458 & ~n43983;
  assign n44458 = pi1072 & n43983;
  assign po615 = n44457 | n44458;
  assign n44460 = pi459 & ~n44303;
  assign n44461 = pi1058 & n44303;
  assign po616 = n44460 | n44461;
  assign n44463 = pi460 & ~n43983;
  assign n44464 = pi1086 & n43983;
  assign po617 = n44463 | n44464;
  assign n44466 = pi461 & ~n43983;
  assign n44467 = pi1057 & n43983;
  assign po618 = n44466 | n44467;
  assign n44469 = pi462 & ~n43983;
  assign n44470 = pi1074 & n43983;
  assign po619 = n44469 | n44470;
  assign n44472 = pi463 & ~n43995;
  assign n44473 = pi1070 & n43995;
  assign po620 = n44472 | n44473;
  assign n44475 = pi464 & ~n44303;
  assign n44476 = pi1065 & n44303;
  assign po621 = n44475 | n44476;
  assign n44478 = ~n5768 & ~n5777;
  assign n44479 = pi1157 & n44478;
  assign n44480 = ~n11334 & ~n11337;
  assign n44481 = ~pi243 & ~n44480;
  assign n44482 = pi926 & ~n44478;
  assign n44483 = ~n44481 & ~n44482;
  assign n44484 = ~n44479 & n44483;
  assign n44485 = ~pi299 & n43891;
  assign n44486 = ~n11360 & ~n44485;
  assign n44487 = ~pi243 & pi1157;
  assign n44488 = ~n44486 & ~n44487;
  assign n44489 = ~n44481 & n44488;
  assign n44490 = ~n3475 & ~n11361;
  assign n44491 = pi926 & n44487;
  assign n44492 = ~n44490 & n44491;
  assign n44493 = ~n44489 & ~n44492;
  assign n44494 = ~n44484 & n44493;
  assign n44495 = ~po1038 & ~n44494;
  assign n44496 = ~pi243 & n43900;
  assign n44497 = po1038 & ~n44496;
  assign n44498 = pi926 & n43902;
  assign n44499 = pi1157 & ~n5788;
  assign n44500 = ~n44498 & ~n44499;
  assign n44501 = n44497 & n44500;
  assign po622 = ~n44495 & ~n44501;
  assign n44503 = po1038 & ~n43900;
  assign n44504 = ~po1038 & n44480;
  assign n44505 = ~n44503 & ~n44504;
  assign n44506 = ~pi943 & ~n44505;
  assign n44507 = pi943 & ~n43950;
  assign n44508 = ~n44506 & ~n44507;
  assign n44509 = ~pi1151 & ~n44508;
  assign n44510 = pi943 & pi1151;
  assign n44511 = ~n43949 & n44510;
  assign n44512 = ~n43889 & n44506;
  assign n44513 = ~po1038 & ~n44486;
  assign n44514 = n3136 & po1038;
  assign n44515 = ~n44513 & ~n44514;
  assign n44516 = ~pi275 & ~n44515;
  assign n44517 = ~n44512 & ~n44516;
  assign n44518 = ~n44511 & n44517;
  assign po623 = ~n44509 & n44518;
  assign n44520 = pi40 & ~pi287;
  assign n44521 = n41737 & n44520;
  assign n44522 = po950 & n44521;
  assign n44523 = ~n10111 & ~n44522;
  assign n44524 = ~pi102 & ~n13297;
  assign n44525 = n8859 & n10108;
  assign n44526 = n16953 & n44525;
  assign n44527 = ~n44524 & n44526;
  assign n44528 = n16951 & n44527;
  assign n44529 = n44521 & ~n44528;
  assign n44530 = ~n44521 & n44528;
  assign n44531 = ~n44529 & ~n44530;
  assign n44532 = ~n6258 & ~n44531;
  assign n44533 = n6258 & n44528;
  assign n44534 = ~n44532 & ~n44533;
  assign n44535 = ~n7538 & ~n44534;
  assign n44536 = n7538 & ~n44531;
  assign n44537 = pi1091 & ~n44536;
  assign n44538 = ~n44535 & n44537;
  assign n44539 = ~n7474 & ~n44531;
  assign n44540 = n7474 & n44528;
  assign n44541 = ~n44539 & ~n44540;
  assign n44542 = pi1093 & ~n44541;
  assign n44543 = ~pi1093 & ~n44534;
  assign n44544 = ~pi1091 & ~n44543;
  assign n44545 = ~n44542 & n44544;
  assign n44546 = ~n44538 & ~n44545;
  assign n44547 = n3222 & n43970;
  assign n44548 = ~n44546 & n44547;
  assign po624 = ~n44523 & ~n44548;
  assign n44550 = n10146 & n11277;
  assign n44551 = pi38 & ~pi39;
  assign n44552 = n10143 & n44551;
  assign n44553 = n8921 & n44552;
  assign n44554 = pi468 & ~n44553;
  assign po625 = n44550 | n44554;
  assign n44556 = pi1156 & n44478;
  assign n44557 = ~pi263 & ~n44480;
  assign n44558 = pi942 & ~n44478;
  assign n44559 = ~n44557 & ~n44558;
  assign n44560 = ~n44556 & n44559;
  assign n44561 = ~pi263 & pi1156;
  assign n44562 = ~n44486 & ~n44561;
  assign n44563 = ~n44557 & n44562;
  assign n44564 = pi942 & n44561;
  assign n44565 = ~n44490 & n44564;
  assign n44566 = ~n44563 & ~n44565;
  assign n44567 = ~n44560 & n44566;
  assign n44568 = ~po1038 & ~n44567;
  assign n44569 = ~pi263 & n43900;
  assign n44570 = po1038 & ~n44569;
  assign n44571 = pi1156 & ~n5788;
  assign n44572 = pi942 & n43902;
  assign n44573 = ~n44571 & ~n44572;
  assign n44574 = n44570 & n44573;
  assign po626 = ~n44568 & ~n44574;
  assign n44576 = pi1155 & n44478;
  assign n44577 = pi267 & ~n44480;
  assign n44578 = pi925 & ~n44478;
  assign n44579 = ~n44577 & ~n44578;
  assign n44580 = ~n44576 & n44579;
  assign n44581 = pi267 & pi1155;
  assign n44582 = ~n44486 & ~n44581;
  assign n44583 = ~n44577 & n44582;
  assign n44584 = pi925 & n44581;
  assign n44585 = ~n44490 & n44584;
  assign n44586 = ~n44583 & ~n44585;
  assign n44587 = ~n44580 & n44586;
  assign n44588 = ~po1038 & ~n44587;
  assign n44589 = pi267 & n43900;
  assign n44590 = po1038 & ~n44589;
  assign n44591 = pi1155 & ~n5788;
  assign n44592 = pi925 & n43902;
  assign n44593 = ~n44591 & ~n44592;
  assign n44594 = n44590 & n44593;
  assign po627 = ~n44588 & ~n44594;
  assign n44596 = pi1153 & n44478;
  assign n44597 = pi253 & ~n44480;
  assign n44598 = pi941 & ~n44478;
  assign n44599 = ~n44597 & ~n44598;
  assign n44600 = ~n44596 & n44599;
  assign n44601 = pi253 & pi1153;
  assign n44602 = ~n44486 & ~n44601;
  assign n44603 = ~n44597 & n44602;
  assign n44604 = pi941 & n44601;
  assign n44605 = ~n44490 & n44604;
  assign n44606 = ~n44603 & ~n44605;
  assign n44607 = ~n44600 & n44606;
  assign n44608 = ~po1038 & ~n44607;
  assign n44609 = pi253 & n43900;
  assign n44610 = po1038 & ~n44609;
  assign n44611 = pi1153 & ~n5788;
  assign n44612 = pi941 & n43902;
  assign n44613 = ~n44611 & ~n44612;
  assign n44614 = n44610 & n44613;
  assign po628 = ~n44608 & ~n44614;
  assign n44616 = pi1154 & n44478;
  assign n44617 = pi254 & ~n44480;
  assign n44618 = pi923 & ~n44478;
  assign n44619 = ~n44617 & ~n44618;
  assign n44620 = ~n44616 & n44619;
  assign n44621 = pi254 & pi1154;
  assign n44622 = ~n44486 & ~n44621;
  assign n44623 = ~n44617 & n44622;
  assign n44624 = pi923 & n44621;
  assign n44625 = ~n44490 & n44624;
  assign n44626 = ~n44623 & ~n44625;
  assign n44627 = ~n44620 & n44626;
  assign n44628 = ~po1038 & ~n44627;
  assign n44629 = pi254 & n43900;
  assign n44630 = po1038 & ~n44629;
  assign n44631 = pi1154 & ~n5788;
  assign n44632 = pi923 & n43902;
  assign n44633 = ~n44631 & ~n44632;
  assign n44634 = n44630 & n44633;
  assign po629 = ~n44628 & ~n44634;
  assign n44636 = ~pi922 & ~n44505;
  assign n44637 = pi922 & ~n43950;
  assign n44638 = ~n44636 & ~n44637;
  assign n44639 = ~pi1152 & ~n44638;
  assign n44640 = pi922 & pi1152;
  assign n44641 = ~n43949 & n44640;
  assign n44642 = ~n43889 & n44636;
  assign n44643 = ~pi268 & ~n44515;
  assign n44644 = ~n44642 & ~n44643;
  assign n44645 = ~n44641 & n44644;
  assign po630 = ~n44639 & n44645;
  assign n44647 = ~pi931 & ~n44505;
  assign n44648 = pi931 & ~n43950;
  assign n44649 = ~n44647 & ~n44648;
  assign n44650 = ~pi1150 & ~n44649;
  assign n44651 = pi931 & pi1150;
  assign n44652 = ~n43949 & n44651;
  assign n44653 = ~n43889 & n44647;
  assign n44654 = ~pi272 & ~n44515;
  assign n44655 = ~n44653 & ~n44654;
  assign n44656 = ~n44652 & n44655;
  assign po631 = ~n44650 & n44656;
  assign n44658 = ~pi936 & ~n44505;
  assign n44659 = pi936 & ~n43950;
  assign n44660 = ~n44658 & ~n44659;
  assign n44661 = ~pi1149 & ~n44660;
  assign n44662 = pi936 & pi1149;
  assign n44663 = ~n43949 & n44662;
  assign n44664 = ~n43889 & n44658;
  assign n44665 = ~pi283 & ~n44515;
  assign n44666 = ~n44664 & ~n44665;
  assign n44667 = ~n44663 & n44666;
  assign po632 = ~n44661 & n44667;
  assign n44669 = pi71 & n43003;
  assign n44670 = pi71 & ~n11385;
  assign n44671 = n11385 & n12965;
  assign n44672 = n10097 & ~n11385;
  assign n44673 = n10093 & n44672;
  assign n44674 = ~n44671 & ~n44673;
  assign n44675 = n3268 & n10108;
  assign n44676 = ~n44674 & n44675;
  assign n44677 = n12973 & n44676;
  assign n44678 = ~n44670 & ~n44677;
  assign n44679 = ~po1038 & ~n44678;
  assign po633 = n44669 | n44679;
  assign po635 = pi71 & ~n43182;
  assign n44682 = pi481 & ~n34556;
  assign n44683 = pi248 & n34556;
  assign po638 = n44682 | n44683;
  assign n44685 = pi482 & ~n34572;
  assign n44686 = pi249 & n34572;
  assign po639 = n44685 | n44686;
  assign n44688 = pi483 & ~n34695;
  assign n44689 = pi242 & n34695;
  assign po640 = n44688 | n44689;
  assign n44691 = pi484 & ~n34695;
  assign n44692 = pi249 & n34695;
  assign po641 = n44691 | n44692;
  assign n44694 = pi485 & ~n35884;
  assign n44695 = pi234 & n35884;
  assign po642 = n44694 | n44695;
  assign n44697 = pi486 & ~n35884;
  assign n44698 = pi244 & n35884;
  assign po643 = n44697 | n44698;
  assign n44700 = pi487 & ~n34556;
  assign n44701 = pi246 & n34556;
  assign po644 = n44700 | n44701;
  assign n44703 = pi488 & ~n34556;
  assign n44704 = ~pi239 & n34556;
  assign po645 = ~n44703 & ~n44704;
  assign n44706 = pi489 & ~n35884;
  assign n44707 = pi242 & n35884;
  assign po646 = n44706 | n44707;
  assign n44709 = pi490 & ~n34695;
  assign n44710 = pi241 & n34695;
  assign po647 = n44709 | n44710;
  assign n44712 = pi491 & ~n34695;
  assign n44713 = pi238 & n34695;
  assign po648 = n44712 | n44713;
  assign n44715 = pi492 & ~n34695;
  assign n44716 = pi240 & n34695;
  assign po649 = n44715 | n44716;
  assign n44718 = pi493 & ~n34695;
  assign n44719 = pi244 & n34695;
  assign po650 = n44718 | n44719;
  assign n44721 = pi494 & ~n34695;
  assign n44722 = ~pi239 & n34695;
  assign po651 = ~n44721 & ~n44722;
  assign n44724 = pi495 & ~n34695;
  assign n44725 = pi235 & n34695;
  assign po652 = n44724 | n44725;
  assign n44727 = pi496 & ~n34687;
  assign n44728 = pi249 & n34687;
  assign po653 = n44727 | n44728;
  assign n44730 = pi497 & ~n34687;
  assign n44731 = ~pi239 & n34687;
  assign po654 = ~n44730 & ~n44731;
  assign n44733 = pi498 & ~n34572;
  assign n44734 = pi238 & n34572;
  assign po655 = n44733 | n44734;
  assign n44736 = pi499 & ~n34687;
  assign n44737 = pi246 & n34687;
  assign po656 = n44736 | n44737;
  assign n44739 = pi500 & ~n34687;
  assign n44740 = pi241 & n34687;
  assign po657 = n44739 | n44740;
  assign n44742 = pi501 & ~n34687;
  assign n44743 = pi248 & n34687;
  assign po658 = n44742 | n44743;
  assign n44745 = pi502 & ~n34687;
  assign n44746 = pi247 & n34687;
  assign po659 = n44745 | n44746;
  assign n44748 = pi503 & ~n34687;
  assign n44749 = pi245 & n34687;
  assign po660 = n44748 | n44749;
  assign n44751 = pi504 & ~n34680;
  assign n44752 = pi242 & n34680;
  assign po661 = n44751 | n44752;
  assign n44754 = ~pi234 & n34678;
  assign n44755 = n34687 & n44754;
  assign n44756 = pi505 & ~n44755;
  assign n44757 = pi234 & n34679;
  assign n44758 = ~pi505 & n34559;
  assign n44759 = n44757 & n44758;
  assign po662 = n44756 | n44759;
  assign n44761 = pi506 & ~n34680;
  assign n44762 = pi241 & n34680;
  assign po663 = n44761 | n44762;
  assign n44764 = pi507 & ~n34680;
  assign n44765 = pi238 & n34680;
  assign po664 = n44764 | n44765;
  assign n44767 = pi508 & ~n34680;
  assign n44768 = pi247 & n34680;
  assign po665 = n44767 | n44768;
  assign n44770 = pi509 & ~n34680;
  assign n44771 = pi245 & n34680;
  assign po666 = n44770 | n44771;
  assign n44773 = pi510 & ~n34556;
  assign n44774 = pi242 & n34556;
  assign po667 = n44773 | n44774;
  assign n44776 = ~pi234 & n34551;
  assign n44777 = n34556 & ~n44776;
  assign n44778 = pi511 & ~n34556;
  assign po668 = n44777 | n44778;
  assign n44780 = pi512 & ~n34556;
  assign n44781 = pi235 & n34556;
  assign po669 = n44780 | n44781;
  assign n44783 = pi513 & ~n34556;
  assign n44784 = pi244 & n34556;
  assign po670 = n44783 | n44784;
  assign n44786 = pi514 & ~n34556;
  assign n44787 = pi245 & n34556;
  assign po671 = n44786 | n44787;
  assign n44789 = pi515 & ~n34556;
  assign n44790 = pi240 & n34556;
  assign po672 = n44789 | n44790;
  assign n44792 = pi516 & ~n34556;
  assign n44793 = pi247 & n34556;
  assign po673 = n44792 | n44793;
  assign n44795 = pi517 & ~n34556;
  assign n44796 = pi238 & n34556;
  assign po674 = n44795 | n44796;
  assign n44798 = n34564 & n44776;
  assign n44799 = pi518 & ~n44798;
  assign n44800 = pi234 & n34555;
  assign n44801 = ~pi518 & n34559;
  assign n44802 = n44800 & n44801;
  assign po675 = n44799 | n44802;
  assign n44804 = pi519 & ~n34564;
  assign n44805 = ~pi239 & n34564;
  assign po676 = ~n44804 & ~n44805;
  assign n44807 = pi520 & ~n34564;
  assign n44808 = pi246 & n34564;
  assign po677 = n44807 | n44808;
  assign n44810 = pi521 & ~n34564;
  assign n44811 = pi248 & n34564;
  assign po678 = n44810 | n44811;
  assign n44813 = pi522 & ~n34564;
  assign n44814 = pi238 & n34564;
  assign po679 = n44813 | n44814;
  assign n44816 = n35912 & n44776;
  assign n44817 = pi523 & ~n44816;
  assign n44818 = ~pi523 & n34690;
  assign n44819 = n44800 & n44818;
  assign po680 = n44817 | n44819;
  assign n44821 = pi524 & ~n35912;
  assign n44822 = ~pi239 & n35912;
  assign po681 = ~n44821 & ~n44822;
  assign n44824 = pi525 & ~n35912;
  assign n44825 = pi245 & n35912;
  assign po682 = n44824 | n44825;
  assign n44827 = pi526 & ~n35912;
  assign n44828 = pi246 & n35912;
  assign po683 = n44827 | n44828;
  assign n44830 = pi527 & ~n35912;
  assign n44831 = pi247 & n35912;
  assign po684 = n44830 | n44831;
  assign n44833 = pi528 & ~n35912;
  assign n44834 = pi249 & n35912;
  assign po685 = n44833 | n44834;
  assign n44836 = pi529 & ~n35912;
  assign n44837 = pi238 & n35912;
  assign po686 = n44836 | n44837;
  assign n44839 = pi530 & ~n35912;
  assign n44840 = pi240 & n35912;
  assign po687 = n44839 | n44840;
  assign n44842 = pi531 & ~n34572;
  assign n44843 = pi235 & n34572;
  assign po688 = n44842 | n44843;
  assign n44845 = pi532 & ~n34572;
  assign n44846 = pi247 & n34572;
  assign po689 = n44845 | n44846;
  assign n44848 = pi533 & ~n34680;
  assign n44849 = pi235 & n34680;
  assign po690 = n44848 | n44849;
  assign n44851 = pi534 & ~n34680;
  assign n44852 = ~pi239 & n34680;
  assign po691 = ~n44851 & ~n44852;
  assign n44854 = pi535 & ~n34680;
  assign n44855 = pi240 & n34680;
  assign po692 = n44854 | n44855;
  assign n44857 = pi536 & ~n34680;
  assign n44858 = pi246 & n34680;
  assign po693 = n44857 | n44858;
  assign n44860 = pi537 & ~n34680;
  assign n44861 = pi248 & n34680;
  assign po694 = n44860 | n44861;
  assign n44863 = pi538 & ~n34680;
  assign n44864 = pi249 & n34680;
  assign po695 = n44863 | n44864;
  assign n44866 = pi539 & ~n34687;
  assign n44867 = pi242 & n34687;
  assign po696 = n44866 | n44867;
  assign n44869 = pi540 & ~n34687;
  assign n44870 = pi235 & n34687;
  assign po697 = n44869 | n44870;
  assign n44872 = pi541 & ~n34687;
  assign n44873 = pi244 & n34687;
  assign po698 = n44872 | n44873;
  assign n44875 = pi542 & ~n34687;
  assign n44876 = pi240 & n34687;
  assign po699 = n44875 | n44876;
  assign n44878 = pi543 & ~n34687;
  assign n44879 = pi238 & n34687;
  assign po700 = n44878 | n44879;
  assign n44881 = n34695 & n44754;
  assign n44882 = pi544 & ~n44881;
  assign n44883 = ~pi544 & n34690;
  assign n44884 = n44757 & n44883;
  assign po701 = n44882 | n44884;
  assign n44886 = pi545 & ~n34695;
  assign n44887 = pi245 & n34695;
  assign po702 = n44886 | n44887;
  assign n44889 = pi546 & ~n34695;
  assign n44890 = pi246 & n34695;
  assign po703 = n44889 | n44890;
  assign n44892 = pi547 & ~n34695;
  assign n44893 = pi247 & n34695;
  assign po704 = n44892 | n44893;
  assign n44895 = pi548 & ~n34695;
  assign n44896 = pi248 & n34695;
  assign po705 = n44895 | n44896;
  assign n44898 = pi549 & ~n35884;
  assign n44899 = pi235 & n35884;
  assign po706 = n44898 | n44899;
  assign n44901 = pi550 & ~n35884;
  assign n44902 = ~pi239 & n35884;
  assign po707 = ~n44901 & ~n44902;
  assign n44904 = pi551 & ~n35884;
  assign n44905 = pi240 & n35884;
  assign po708 = n44904 | n44905;
  assign n44907 = pi552 & ~n35884;
  assign n44908 = pi247 & n35884;
  assign po709 = n44907 | n44908;
  assign n44910 = pi553 & ~n35884;
  assign n44911 = pi241 & n35884;
  assign po710 = n44910 | n44911;
  assign n44913 = pi554 & ~n35884;
  assign n44914 = pi248 & n35884;
  assign po711 = n44913 | n44914;
  assign n44916 = pi555 & ~n35884;
  assign n44917 = pi249 & n35884;
  assign po712 = n44916 | n44917;
  assign n44919 = pi556 & ~n34572;
  assign n44920 = pi242 & n34572;
  assign po713 = n44919 | n44920;
  assign n44922 = n34680 & n44754;
  assign n44923 = pi557 & ~n44922;
  assign n44924 = ~pi557 & n34364;
  assign n44925 = n44757 & n44924;
  assign po714 = n44923 | n44925;
  assign n44927 = pi558 & ~n34680;
  assign n44928 = pi244 & n34680;
  assign po715 = n44927 | n44928;
  assign n44930 = pi559 & ~n34556;
  assign n44931 = pi241 & n34556;
  assign po716 = n44930 | n44931;
  assign n44933 = pi560 & ~n34572;
  assign n44934 = pi240 & n34572;
  assign po717 = n44933 | n44934;
  assign n44936 = pi561 & ~n34564;
  assign n44937 = pi247 & n34564;
  assign po718 = n44936 | n44937;
  assign n44939 = pi562 & ~n34572;
  assign n44940 = pi241 & n34572;
  assign po719 = n44939 | n44940;
  assign n44942 = pi563 & ~n35884;
  assign n44943 = pi246 & n35884;
  assign po720 = n44942 | n44943;
  assign n44945 = pi564 & ~n34572;
  assign n44946 = pi246 & n34572;
  assign po721 = n44945 | n44946;
  assign n44948 = pi565 & ~n34572;
  assign n44949 = pi248 & n34572;
  assign po722 = n44948 | n44949;
  assign n44951 = pi566 & ~n34572;
  assign n44952 = pi244 & n34572;
  assign po723 = n44951 | n44952;
  assign n44954 = ~pi567 & pi1092;
  assign n44955 = ~pi1093 & n44954;
  assign n44956 = pi680 & n17371;
  assign n44957 = ~n19038 & n44956;
  assign n44958 = ~n44955 & ~n44957;
  assign n44959 = n19127 & ~n44958;
  assign n44960 = ~n17539 & n44959;
  assign n44961 = pi603 & ~n17438;
  assign n44962 = n16740 & ~n20069;
  assign n44963 = ~n20075 & n44962;
  assign n44964 = n44961 & n44963;
  assign n44965 = pi619 & n44964;
  assign n44966 = ~n44955 & ~n44965;
  assign n44967 = pi1159 & ~n44966;
  assign n44968 = ~pi619 & n44964;
  assign n44969 = ~n44955 & ~n44968;
  assign n44970 = ~pi1159 & ~n44969;
  assign n44971 = pi789 & ~n44970;
  assign n44972 = ~n44967 & n44971;
  assign n44973 = ~n44964 & n44966;
  assign n44974 = ~n44972 & ~n44973;
  assign n44975 = ~n44960 & ~n44974;
  assign n44976 = n17817 & ~n44975;
  assign n44977 = n35039 & n44974;
  assign n44978 = pi641 & n44960;
  assign n44979 = ~n44955 & ~n44978;
  assign n44980 = n17698 & ~n44979;
  assign n44981 = ~pi641 & n44960;
  assign n44982 = ~n44955 & ~n44981;
  assign n44983 = n17699 & ~n44982;
  assign n44984 = ~n44980 & ~n44983;
  assign n44985 = ~n44977 & n44984;
  assign n44986 = pi788 & ~n44985;
  assign n44987 = ~n44976 & ~n44986;
  assign n44988 = ~n20205 & ~n44987;
  assign n44989 = ~n17816 & n44974;
  assign n44990 = n17816 & n44955;
  assign n44991 = ~n44989 & ~n44990;
  assign n44992 = n17855 & ~n44991;
  assign n44993 = n19128 & ~n44958;
  assign n44994 = ~pi628 & n44993;
  assign n44995 = ~n44955 & ~n44994;
  assign n44996 = ~pi1156 & ~n44995;
  assign n44997 = pi629 & ~n44996;
  assign n44998 = ~n44992 & n44997;
  assign n44999 = n17856 & ~n44991;
  assign n45000 = pi628 & n44993;
  assign n45001 = ~n44955 & ~n45000;
  assign n45002 = pi1156 & ~n45001;
  assign n45003 = ~pi629 & ~n45002;
  assign n45004 = ~n44999 & n45003;
  assign n45005 = pi792 & ~n45004;
  assign n45006 = ~n44998 & n45005;
  assign n45007 = ~n44988 & ~n45006;
  assign n45008 = ~pi647 & ~n45007;
  assign n45009 = ~n17610 & ~n44991;
  assign n45010 = ~n44955 & ~n45009;
  assign n45011 = pi647 & ~n45010;
  assign n45012 = ~pi1157 & ~n45011;
  assign n45013 = ~n45008 & n45012;
  assign n45014 = ~n19158 & n44993;
  assign n45015 = pi647 & n45014;
  assign n45016 = pi1157 & ~n44955;
  assign n45017 = ~n45015 & n45016;
  assign n45018 = ~pi630 & ~n45017;
  assign n45019 = ~n45013 & n45018;
  assign n45020 = pi647 & ~n45007;
  assign n45021 = ~pi647 & ~n45010;
  assign n45022 = pi1157 & ~n45021;
  assign n45023 = ~n45020 & n45022;
  assign n45024 = ~pi647 & n45014;
  assign n45025 = ~pi1157 & ~n44955;
  assign n45026 = ~n45024 & n45025;
  assign n45027 = pi630 & ~n45026;
  assign n45028 = ~n45023 & n45027;
  assign n45029 = ~n45019 & ~n45028;
  assign n45030 = pi787 & ~n45029;
  assign n45031 = ~pi787 & ~n45007;
  assign n45032 = ~n45030 & ~n45031;
  assign n45033 = ~pi790 & ~n45032;
  assign n45034 = ~pi644 & ~n45032;
  assign n45035 = ~n19182 & n45014;
  assign n45036 = ~n44955 & ~n45035;
  assign n45037 = pi644 & ~n45036;
  assign n45038 = ~pi715 & ~n45037;
  assign n45039 = ~n45034 & n45038;
  assign n45040 = ~n17652 & n45009;
  assign n45041 = ~pi644 & n45040;
  assign n45042 = pi715 & ~n44955;
  assign n45043 = ~n45041 & n45042;
  assign n45044 = ~n45039 & ~n45043;
  assign n45045 = ~pi1160 & ~n45044;
  assign n45046 = pi644 & n45032;
  assign n45047 = ~pi644 & n45036;
  assign n45048 = pi715 & ~n45047;
  assign n45049 = ~n45046 & n45048;
  assign n45050 = pi644 & n45040;
  assign n45051 = ~n44955 & ~n45050;
  assign n45052 = ~pi715 & ~n45051;
  assign n45053 = pi1160 & ~n45052;
  assign n45054 = ~n45049 & n45053;
  assign n45055 = pi790 & ~n45054;
  assign n45056 = ~n45045 & n45055;
  assign n45057 = ~n45033 & ~n45056;
  assign n45058 = pi230 & ~n45057;
  assign n45059 = ~pi230 & n44954;
  assign po724 = n45058 | n45059;
  assign n45061 = pi568 & ~n34572;
  assign n45062 = pi245 & n34572;
  assign po725 = n45061 | n45062;
  assign n45064 = pi569 & ~n34572;
  assign n45065 = ~pi239 & n34572;
  assign po726 = ~n45064 & ~n45065;
  assign n45067 = n34572 & n44776;
  assign n45068 = pi570 & ~n45067;
  assign n45069 = ~pi570 & n34567;
  assign n45070 = n44800 & n45069;
  assign po727 = n45068 | n45070;
  assign n45072 = pi571 & ~n35912;
  assign n45073 = pi241 & n35912;
  assign po728 = n45072 | n45073;
  assign n45075 = pi572 & ~n35912;
  assign n45076 = pi244 & n35912;
  assign po729 = n45075 | n45076;
  assign n45078 = pi573 & ~n35912;
  assign n45079 = pi242 & n35912;
  assign po730 = n45078 | n45079;
  assign n45081 = pi574 & ~n34564;
  assign n45082 = pi241 & n34564;
  assign po731 = n45081 | n45082;
  assign n45084 = pi575 & ~n35912;
  assign n45085 = pi235 & n35912;
  assign po732 = n45084 | n45085;
  assign n45087 = pi576 & ~n35912;
  assign n45088 = pi248 & n35912;
  assign po733 = n45087 | n45088;
  assign n45090 = pi577 & ~n35884;
  assign n45091 = pi238 & n35884;
  assign po734 = n45090 | n45091;
  assign n45093 = pi578 & ~n34564;
  assign n45094 = pi249 & n34564;
  assign po735 = n45093 | n45094;
  assign n45096 = pi579 & ~n34556;
  assign n45097 = pi249 & n34556;
  assign po736 = n45096 | n45097;
  assign n45099 = pi580 & ~n35884;
  assign n45100 = pi245 & n35884;
  assign po737 = n45099 | n45100;
  assign n45102 = pi581 & ~n34564;
  assign n45103 = pi235 & n34564;
  assign po738 = n45102 | n45103;
  assign n45105 = pi582 & ~n34564;
  assign n45106 = pi240 & n34564;
  assign po739 = n45105 | n45106;
  assign n45108 = pi584 & ~n34564;
  assign n45109 = pi245 & n34564;
  assign po741 = n45108 | n45109;
  assign n45111 = pi585 & ~n34564;
  assign n45112 = pi244 & n34564;
  assign po742 = n45111 | n45112;
  assign n45114 = pi586 & ~n34564;
  assign n45115 = pi242 & n34564;
  assign po743 = n45114 | n45115;
  assign n45117 = ~pi230 & pi587;
  assign n45118 = pi230 & n16521;
  assign n45119 = ~n20069 & n45118;
  assign n45120 = ~n35416 & n45119;
  assign n45121 = n20081 & n45120;
  assign n45122 = n30600 & n45121;
  assign po744 = n45117 | n45122;
  assign n45124 = ~pi123 & n12135;
  assign n45125 = ~pi591 & n45124;
  assign n45126 = ~pi588 & ~n45124;
  assign n45127 = n44032 & ~n45126;
  assign po745 = ~n45125 & n45127;
  assign n45129 = ~pi201 & n34551;
  assign n45130 = ~pi204 & n34678;
  assign n45131 = pi233 & ~n45130;
  assign n45132 = ~n45129 & n45131;
  assign n45133 = ~pi202 & n34551;
  assign n45134 = ~pi205 & n34678;
  assign n45135 = ~pi233 & ~n45134;
  assign n45136 = ~n45133 & n45135;
  assign n45137 = ~n45132 & ~n45136;
  assign n45138 = pi237 & ~n45137;
  assign n45139 = ~pi220 & n34551;
  assign n45140 = ~pi206 & n34678;
  assign n45141 = pi233 & ~n45140;
  assign n45142 = ~n45139 & n45141;
  assign n45143 = ~pi203 & n34551;
  assign n45144 = ~pi218 & n34678;
  assign n45145 = ~pi233 & ~n45144;
  assign n45146 = ~n45143 & n45145;
  assign n45147 = ~n45142 & ~n45146;
  assign n45148 = ~pi237 & ~n45147;
  assign po746 = ~n45138 & ~n45148;
  assign n45150 = pi590 & ~n45124;
  assign n45151 = pi588 & n45124;
  assign n45152 = n44032 & ~n45151;
  assign po747 = n45150 | ~n45152;
  assign n45154 = ~pi592 & n45124;
  assign n45155 = ~pi591 & ~n45124;
  assign n45156 = n44032 & ~n45155;
  assign po748 = ~n45154 & n45156;
  assign n45158 = ~pi590 & n45124;
  assign n45159 = ~pi592 & ~n45124;
  assign n45160 = n44032 & ~n45159;
  assign po749 = ~n45158 & n45160;
  assign n45162 = pi234 & n34678;
  assign n45163 = pi557 & ~n45162;
  assign n45164 = pi246 & pi536;
  assign n45165 = ~pi246 & ~pi536;
  assign n45166 = ~n45164 & ~n45165;
  assign n45167 = ~pi557 & ~n44754;
  assign n45168 = ~n45166 & ~n45167;
  assign n45169 = ~n45163 & n45168;
  assign n45170 = ~pi538 & n45169;
  assign n45171 = ~pi249 & ~n45170;
  assign n45172 = pi538 & n45169;
  assign n45173 = pi249 & ~n45172;
  assign n45174 = ~n45171 & ~n45173;
  assign n45175 = ~pi537 & n45174;
  assign n45176 = ~pi248 & ~n45175;
  assign n45177 = pi537 & n45174;
  assign n45178 = pi248 & ~n45177;
  assign n45179 = ~n45176 & ~n45178;
  assign n45180 = pi241 & pi506;
  assign n45181 = ~pi241 & ~pi506;
  assign n45182 = ~n45180 & ~n45181;
  assign n45183 = n45179 & ~n45182;
  assign n45184 = pi240 & pi535;
  assign n45185 = ~pi240 & ~pi535;
  assign n45186 = ~n45184 & ~n45185;
  assign n45187 = n45183 & ~n45186;
  assign n45188 = pi534 & n45187;
  assign n45189 = ~pi239 & ~n45188;
  assign n45190 = ~pi534 & n45187;
  assign n45191 = pi239 & ~n45190;
  assign n45192 = ~n45189 & ~n45191;
  assign n45193 = pi504 & n45192;
  assign n45194 = pi242 & ~n45193;
  assign n45195 = ~pi504 & n45192;
  assign n45196 = ~pi242 & ~n45195;
  assign n45197 = ~n45194 & ~n45196;
  assign n45198 = pi533 & n45197;
  assign n45199 = pi235 & ~n45198;
  assign n45200 = ~pi533 & n45197;
  assign n45201 = ~pi235 & ~n45200;
  assign n45202 = ~n45199 & ~n45201;
  assign n45203 = pi558 & n45202;
  assign n45204 = pi244 & ~n45203;
  assign n45205 = ~pi558 & n45202;
  assign n45206 = ~pi244 & ~n45205;
  assign n45207 = ~n45204 & ~n45206;
  assign n45208 = pi509 & n45207;
  assign n45209 = pi245 & ~n45208;
  assign n45210 = ~pi509 & n45207;
  assign n45211 = ~pi245 & ~n45210;
  assign n45212 = ~n45209 & ~n45211;
  assign n45213 = pi508 & n45212;
  assign n45214 = pi247 & ~n45213;
  assign n45215 = pi248 & pi481;
  assign n45216 = ~pi248 & ~pi481;
  assign n45217 = ~n45215 & ~n45216;
  assign n45218 = pi234 & n34551;
  assign n45219 = pi511 & ~n45218;
  assign n45220 = pi246 & pi487;
  assign n45221 = ~pi246 & ~pi487;
  assign n45222 = ~n45220 & ~n45221;
  assign n45223 = ~pi511 & ~n44776;
  assign n45224 = ~n45222 & ~n45223;
  assign n45225 = ~n45219 & n45224;
  assign n45226 = ~pi249 & ~pi579;
  assign n45227 = pi249 & pi579;
  assign n45228 = ~n45226 & ~n45227;
  assign n45229 = n45225 & ~n45228;
  assign n45230 = ~n45217 & n45229;
  assign n45231 = pi559 & n45230;
  assign n45232 = pi241 & ~n45231;
  assign n45233 = ~pi559 & n45230;
  assign n45234 = ~pi241 & ~n45233;
  assign n45235 = ~n45232 & ~n45234;
  assign n45236 = pi515 & n45235;
  assign n45237 = pi240 & ~n45236;
  assign n45238 = ~pi579 & ~n45229;
  assign n45239 = ~n45171 & n45225;
  assign n45240 = pi579 & ~n45239;
  assign n45241 = ~n45238 & ~n45240;
  assign n45242 = ~n45174 & ~n45241;
  assign n45243 = ~pi537 & ~n45242;
  assign n45244 = pi537 & n45229;
  assign n45245 = ~pi248 & ~n45244;
  assign n45246 = ~n45243 & n45245;
  assign n45247 = ~n45178 & ~n45246;
  assign n45248 = ~pi481 & ~n45247;
  assign n45249 = pi537 & ~n45242;
  assign n45250 = ~pi537 & n45229;
  assign n45251 = pi248 & ~n45250;
  assign n45252 = ~n45249 & n45251;
  assign n45253 = ~n45176 & ~n45252;
  assign n45254 = pi481 & ~n45253;
  assign n45255 = ~n45248 & ~n45254;
  assign n45256 = ~pi559 & n45255;
  assign n45257 = pi559 & n45179;
  assign n45258 = ~pi241 & ~n45257;
  assign n45259 = ~n45256 & n45258;
  assign n45260 = ~n45232 & ~n45259;
  assign n45261 = ~pi506 & ~n45260;
  assign n45262 = pi559 & n45255;
  assign n45263 = ~pi559 & n45179;
  assign n45264 = pi241 & ~n45263;
  assign n45265 = ~n45262 & n45264;
  assign n45266 = ~n45234 & ~n45265;
  assign n45267 = pi506 & ~n45266;
  assign n45268 = ~n45261 & ~n45267;
  assign n45269 = ~pi515 & n45268;
  assign n45270 = pi515 & n45183;
  assign n45271 = ~pi240 & ~n45270;
  assign n45272 = ~n45269 & n45271;
  assign n45273 = ~n45237 & ~n45272;
  assign n45274 = ~pi535 & ~n45273;
  assign n45275 = ~pi515 & n45235;
  assign n45276 = ~pi240 & ~n45275;
  assign n45277 = pi515 & n45268;
  assign n45278 = ~pi515 & n45183;
  assign n45279 = pi240 & ~n45278;
  assign n45280 = ~n45277 & n45279;
  assign n45281 = ~n45276 & ~n45280;
  assign n45282 = pi535 & ~n45281;
  assign n45283 = ~n45274 & ~n45282;
  assign n45284 = ~pi534 & n45283;
  assign n45285 = ~n45237 & ~n45276;
  assign n45286 = pi534 & n45285;
  assign n45287 = pi239 & ~n45286;
  assign n45288 = ~n45284 & n45287;
  assign n45289 = ~n45189 & ~n45288;
  assign n45290 = ~pi488 & ~n45289;
  assign n45291 = pi534 & n45283;
  assign n45292 = ~pi534 & n45285;
  assign n45293 = ~pi239 & ~n45292;
  assign n45294 = ~n45291 & n45293;
  assign n45295 = ~n45191 & ~n45294;
  assign n45296 = pi488 & ~n45295;
  assign n45297 = ~n45290 & ~n45296;
  assign n45298 = ~pi504 & n45297;
  assign n45299 = ~pi239 & pi488;
  assign n45300 = pi239 & ~pi488;
  assign n45301 = ~n45299 & ~n45300;
  assign n45302 = n45285 & ~n45301;
  assign n45303 = pi504 & n45302;
  assign n45304 = ~pi242 & ~n45303;
  assign n45305 = ~n45298 & n45304;
  assign n45306 = ~n45194 & ~n45305;
  assign n45307 = ~pi510 & ~n45306;
  assign n45308 = pi504 & n45297;
  assign n45309 = ~pi504 & n45302;
  assign n45310 = pi242 & ~n45309;
  assign n45311 = ~n45308 & n45310;
  assign n45312 = ~n45196 & ~n45311;
  assign n45313 = pi510 & ~n45312;
  assign n45314 = ~n45307 & ~n45313;
  assign n45315 = ~pi533 & n45314;
  assign n45316 = pi242 & pi510;
  assign n45317 = ~pi242 & ~pi510;
  assign n45318 = ~n45316 & ~n45317;
  assign n45319 = n45302 & ~n45318;
  assign n45320 = pi533 & n45319;
  assign n45321 = ~pi235 & ~n45320;
  assign n45322 = ~n45315 & n45321;
  assign n45323 = ~n45199 & ~n45322;
  assign n45324 = ~pi512 & ~n45323;
  assign n45325 = pi533 & n45314;
  assign n45326 = ~pi533 & n45319;
  assign n45327 = pi235 & ~n45326;
  assign n45328 = ~n45325 & n45327;
  assign n45329 = ~n45201 & ~n45328;
  assign n45330 = pi512 & ~n45329;
  assign n45331 = ~n45324 & ~n45330;
  assign n45332 = ~pi558 & n45331;
  assign n45333 = pi235 & pi512;
  assign n45334 = ~pi235 & ~pi512;
  assign n45335 = ~n45333 & ~n45334;
  assign n45336 = n45319 & ~n45335;
  assign n45337 = pi558 & n45336;
  assign n45338 = ~pi244 & ~n45337;
  assign n45339 = ~n45332 & n45338;
  assign n45340 = ~n45204 & ~n45339;
  assign n45341 = ~pi513 & ~n45340;
  assign n45342 = pi558 & n45331;
  assign n45343 = ~pi558 & n45336;
  assign n45344 = pi244 & ~n45343;
  assign n45345 = ~n45342 & n45344;
  assign n45346 = ~n45206 & ~n45345;
  assign n45347 = pi513 & ~n45346;
  assign n45348 = ~n45341 & ~n45347;
  assign n45349 = ~pi509 & n45348;
  assign n45350 = pi244 & pi513;
  assign n45351 = ~pi244 & ~pi513;
  assign n45352 = ~n45350 & ~n45351;
  assign n45353 = n45336 & ~n45352;
  assign n45354 = pi509 & n45353;
  assign n45355 = ~pi245 & ~n45354;
  assign n45356 = ~n45349 & n45355;
  assign n45357 = ~n45209 & ~n45356;
  assign n45358 = ~pi514 & ~n45357;
  assign n45359 = pi509 & n45348;
  assign n45360 = ~pi509 & n45353;
  assign n45361 = pi245 & ~n45360;
  assign n45362 = ~n45359 & n45361;
  assign n45363 = ~n45211 & ~n45362;
  assign n45364 = pi514 & ~n45363;
  assign n45365 = ~n45358 & ~n45364;
  assign n45366 = ~pi508 & n45365;
  assign n45367 = pi245 & pi514;
  assign n45368 = ~pi245 & ~pi514;
  assign n45369 = ~n45367 & ~n45368;
  assign n45370 = n45353 & ~n45369;
  assign n45371 = pi508 & n45370;
  assign n45372 = ~pi247 & ~n45371;
  assign n45373 = ~n45366 & n45372;
  assign n45374 = ~n45214 & ~n45373;
  assign n45375 = ~pi516 & ~n45374;
  assign n45376 = ~pi508 & n45212;
  assign n45377 = ~pi247 & ~n45376;
  assign n45378 = pi508 & n45365;
  assign n45379 = ~pi508 & n45370;
  assign n45380 = pi247 & ~n45379;
  assign n45381 = ~n45378 & n45380;
  assign n45382 = ~n45377 & ~n45381;
  assign n45383 = pi516 & ~n45382;
  assign n45384 = ~n45375 & ~n45383;
  assign n45385 = ~pi238 & n45384;
  assign n45386 = ~pi517 & ~n45385;
  assign n45387 = ~n45214 & ~n45377;
  assign n45388 = ~pi238 & n45387;
  assign n45389 = pi247 & pi516;
  assign n45390 = ~pi247 & ~pi516;
  assign n45391 = ~n45389 & ~n45390;
  assign n45392 = n45370 & ~n45391;
  assign n45393 = pi238 & n45392;
  assign n45394 = pi517 & ~n45393;
  assign n45395 = ~n45388 & n45394;
  assign n45396 = ~pi507 & ~n45395;
  assign n45397 = ~n45386 & n45396;
  assign n45398 = pi238 & n45384;
  assign n45399 = pi517 & ~n45398;
  assign n45400 = pi238 & n45387;
  assign n45401 = ~pi238 & n45392;
  assign n45402 = ~pi517 & ~n45401;
  assign n45403 = ~n45400 & n45402;
  assign n45404 = pi507 & ~n45403;
  assign n45405 = ~n45399 & n45404;
  assign n45406 = ~n45397 & ~n45405;
  assign n45407 = pi233 & ~n45406;
  assign n45408 = pi240 & pi542;
  assign n45409 = ~pi240 & ~pi542;
  assign n45410 = ~n45408 & ~n45409;
  assign n45411 = ~pi505 & ~n44754;
  assign n45412 = pi505 & ~n45162;
  assign n45413 = ~pi246 & ~pi499;
  assign n45414 = pi246 & pi499;
  assign n45415 = ~n45413 & ~n45414;
  assign n45416 = ~pi248 & ~pi501;
  assign n45417 = pi248 & pi501;
  assign n45418 = ~n45416 & ~n45417;
  assign n45419 = pi249 & ~pi496;
  assign n45420 = ~pi249 & pi496;
  assign n45421 = ~n45419 & ~n45420;
  assign n45422 = ~n45418 & n45421;
  assign n45423 = ~n45415 & n45422;
  assign n45424 = ~n45412 & n45423;
  assign n45425 = ~n45411 & n45424;
  assign n45426 = ~pi241 & ~pi500;
  assign n45427 = pi241 & pi500;
  assign n45428 = ~n45426 & ~n45427;
  assign n45429 = n45425 & ~n45428;
  assign n45430 = ~n45410 & n45429;
  assign n45431 = pi497 & n45430;
  assign n45432 = ~pi239 & ~n45431;
  assign n45433 = ~pi497 & n45430;
  assign n45434 = pi239 & ~n45433;
  assign n45435 = ~n45432 & ~n45434;
  assign n45436 = pi539 & n45435;
  assign n45437 = pi242 & ~n45436;
  assign n45438 = ~pi539 & n45435;
  assign n45439 = ~pi242 & ~n45438;
  assign n45440 = ~n45437 & ~n45439;
  assign n45441 = pi540 & n45440;
  assign n45442 = pi235 & ~n45441;
  assign n45443 = ~pi540 & n45440;
  assign n45444 = ~pi235 & ~n45443;
  assign n45445 = ~n45442 & ~n45444;
  assign n45446 = pi244 & pi541;
  assign n45447 = ~pi244 & ~pi541;
  assign n45448 = ~n45446 & ~n45447;
  assign n45449 = n45445 & ~n45448;
  assign n45450 = pi245 & pi503;
  assign n45451 = ~pi245 & ~pi503;
  assign n45452 = ~n45450 & ~n45451;
  assign n45453 = n45449 & ~n45452;
  assign n45454 = ~pi502 & n45453;
  assign n45455 = ~pi247 & ~n45454;
  assign n45456 = pi502 & n45453;
  assign n45457 = pi247 & ~n45456;
  assign n45458 = ~n45455 & ~n45457;
  assign n45459 = ~pi238 & n45458;
  assign n45460 = ~pi518 & ~n44776;
  assign n45461 = pi518 & ~n45218;
  assign n45462 = pi249 & ~pi578;
  assign n45463 = ~pi249 & pi578;
  assign n45464 = ~n45462 & ~n45463;
  assign n45465 = pi248 & ~pi521;
  assign n45466 = ~pi248 & pi521;
  assign n45467 = ~n45465 & ~n45466;
  assign n45468 = n45464 & n45467;
  assign n45469 = pi241 & pi574;
  assign n45470 = ~pi241 & ~pi574;
  assign n45471 = ~n45469 & ~n45470;
  assign n45472 = pi246 & ~pi520;
  assign n45473 = ~pi246 & pi520;
  assign n45474 = ~n45472 & ~n45473;
  assign n45475 = ~n45471 & n45474;
  assign n45476 = n45468 & n45475;
  assign n45477 = ~n45461 & n45476;
  assign n45478 = ~n45460 & n45477;
  assign n45479 = pi582 & n45478;
  assign n45480 = pi240 & ~n45479;
  assign n45481 = ~pi582 & n45478;
  assign n45482 = ~pi240 & ~n45481;
  assign n45483 = ~n45480 & ~n45482;
  assign n45484 = ~pi239 & pi519;
  assign n45485 = pi239 & ~pi519;
  assign n45486 = ~n45484 & ~n45485;
  assign n45487 = n45483 & ~n45486;
  assign n45488 = pi242 & pi586;
  assign n45489 = ~pi242 & ~pi586;
  assign n45490 = ~n45488 & ~n45489;
  assign n45491 = n45487 & ~n45490;
  assign n45492 = pi235 & pi581;
  assign n45493 = ~pi235 & ~pi581;
  assign n45494 = ~n45492 & ~n45493;
  assign n45495 = n45491 & ~n45494;
  assign n45496 = pi585 & n45495;
  assign n45497 = pi244 & ~n45496;
  assign n45498 = ~pi585 & n45495;
  assign n45499 = ~pi244 & ~n45498;
  assign n45500 = ~n45497 & ~n45499;
  assign n45501 = pi584 & n45500;
  assign n45502 = pi245 & ~n45501;
  assign n45503 = ~pi584 & n45500;
  assign n45504 = ~pi245 & ~n45503;
  assign n45505 = ~n45502 & ~n45504;
  assign n45506 = ~pi247 & ~pi561;
  assign n45507 = pi247 & pi561;
  assign n45508 = ~n45506 & ~n45507;
  assign n45509 = n45505 & ~n45508;
  assign n45510 = pi238 & n45509;
  assign n45511 = pi522 & ~n45510;
  assign n45512 = ~n45459 & n45511;
  assign n45513 = ~pi543 & ~n45512;
  assign n45514 = ~pi238 & n45509;
  assign n45515 = ~pi522 & ~n45514;
  assign n45516 = ~n45459 & n45515;
  assign n45517 = n45513 & ~n45516;
  assign n45518 = pi238 & n45458;
  assign n45519 = ~n45510 & ~n45518;
  assign n45520 = pi522 & n45519;
  assign n45521 = n45515 & ~n45518;
  assign n45522 = pi543 & ~n45521;
  assign n45523 = ~n45520 & n45522;
  assign n45524 = ~n45517 & ~n45523;
  assign n45525 = ~pi233 & ~n45524;
  assign n45526 = pi237 & ~n45525;
  assign n45527 = ~n45407 & n45526;
  assign n45528 = ~pi240 & ~pi492;
  assign n45529 = pi240 & pi492;
  assign n45530 = ~n45528 & ~n45529;
  assign n45531 = pi241 & pi490;
  assign n45532 = ~pi241 & ~pi490;
  assign n45533 = ~n45531 & ~n45532;
  assign n45534 = pi544 & ~n45162;
  assign n45535 = ~pi544 & ~n44754;
  assign n45536 = pi246 & pi546;
  assign n45537 = ~pi246 & ~pi546;
  assign n45538 = ~n45536 & ~n45537;
  assign n45539 = pi248 & pi548;
  assign n45540 = ~pi248 & ~pi548;
  assign n45541 = ~n45539 & ~n45540;
  assign n45542 = pi249 & pi484;
  assign n45543 = ~pi249 & ~pi484;
  assign n45544 = ~n45542 & ~n45543;
  assign n45545 = ~n45541 & ~n45544;
  assign n45546 = ~n45538 & n45545;
  assign n45547 = ~n45535 & n45546;
  assign n45548 = ~n45534 & n45547;
  assign n45549 = ~n45533 & n45548;
  assign n45550 = ~n45530 & n45549;
  assign n45551 = pi494 & n45550;
  assign n45552 = ~pi239 & ~n45551;
  assign n45553 = ~pi494 & n45550;
  assign n45554 = pi239 & ~n45553;
  assign n45555 = ~n45552 & ~n45554;
  assign n45556 = pi483 & n45555;
  assign n45557 = pi242 & ~n45556;
  assign n45558 = ~pi483 & n45555;
  assign n45559 = ~pi242 & ~n45558;
  assign n45560 = ~n45557 & ~n45559;
  assign n45561 = pi495 & n45560;
  assign n45562 = pi235 & ~n45561;
  assign n45563 = ~pi495 & n45560;
  assign n45564 = ~pi235 & ~n45563;
  assign n45565 = ~n45562 & ~n45564;
  assign n45566 = pi244 & pi493;
  assign n45567 = ~pi244 & ~pi493;
  assign n45568 = ~n45566 & ~n45567;
  assign n45569 = n45565 & ~n45568;
  assign n45570 = pi545 & n45569;
  assign n45571 = pi245 & ~n45570;
  assign n45572 = ~pi545 & n45569;
  assign n45573 = ~pi245 & ~n45572;
  assign n45574 = ~n45571 & ~n45573;
  assign n45575 = pi547 & n45574;
  assign n45576 = pi247 & ~n45575;
  assign n45577 = ~pi547 & n45574;
  assign n45578 = ~pi247 & ~n45577;
  assign n45579 = ~n45576 & ~n45578;
  assign n45580 = ~pi238 & n45579;
  assign n45581 = ~pi523 & ~n44776;
  assign n45582 = pi523 & ~n45218;
  assign n45583 = pi246 & pi526;
  assign n45584 = ~pi246 & ~pi526;
  assign n45585 = ~n45583 & ~n45584;
  assign n45586 = pi248 & pi576;
  assign n45587 = ~pi248 & ~pi576;
  assign n45588 = ~n45586 & ~n45587;
  assign n45589 = pi249 & pi528;
  assign n45590 = ~pi249 & ~pi528;
  assign n45591 = ~n45589 & ~n45590;
  assign n45592 = ~n45588 & ~n45591;
  assign n45593 = ~n45585 & n45592;
  assign n45594 = ~n45582 & n45593;
  assign n45595 = ~n45581 & n45594;
  assign n45596 = pi571 & n45595;
  assign n45597 = pi241 & ~n45596;
  assign n45598 = ~pi571 & n45595;
  assign n45599 = ~pi241 & ~n45598;
  assign n45600 = ~n45597 & ~n45599;
  assign n45601 = ~pi530 & n45600;
  assign n45602 = ~pi240 & ~n45601;
  assign n45603 = pi530 & n45600;
  assign n45604 = pi240 & ~n45603;
  assign n45605 = ~n45602 & ~n45604;
  assign n45606 = ~pi239 & pi524;
  assign n45607 = pi239 & ~pi524;
  assign n45608 = ~n45606 & ~n45607;
  assign n45609 = n45605 & ~n45608;
  assign n45610 = pi242 & pi573;
  assign n45611 = ~pi242 & ~pi573;
  assign n45612 = ~n45610 & ~n45611;
  assign n45613 = n45609 & ~n45612;
  assign n45614 = pi235 & pi575;
  assign n45615 = ~pi235 & ~pi575;
  assign n45616 = ~n45614 & ~n45615;
  assign n45617 = n45613 & ~n45616;
  assign n45618 = pi572 & n45617;
  assign n45619 = pi244 & ~n45618;
  assign n45620 = ~pi572 & n45617;
  assign n45621 = ~pi244 & ~n45620;
  assign n45622 = ~n45619 & ~n45621;
  assign n45623 = pi245 & pi525;
  assign n45624 = ~pi245 & ~pi525;
  assign n45625 = ~n45623 & ~n45624;
  assign n45626 = n45622 & ~n45625;
  assign n45627 = pi247 & pi527;
  assign n45628 = ~pi247 & ~pi527;
  assign n45629 = ~n45627 & ~n45628;
  assign n45630 = n45626 & ~n45629;
  assign n45631 = pi238 & n45630;
  assign n45632 = pi529 & ~n45631;
  assign n45633 = ~n45580 & n45632;
  assign n45634 = ~pi491 & ~n45633;
  assign n45635 = ~pi238 & n45630;
  assign n45636 = ~pi529 & ~n45635;
  assign n45637 = ~n45580 & n45636;
  assign n45638 = n45634 & ~n45637;
  assign n45639 = pi238 & n45579;
  assign n45640 = ~n45631 & ~n45639;
  assign n45641 = pi529 & n45640;
  assign n45642 = n45636 & ~n45639;
  assign n45643 = pi491 & ~n45642;
  assign n45644 = ~n45641 & n45643;
  assign n45645 = ~n45638 & ~n45644;
  assign n45646 = pi233 & ~n45645;
  assign n45647 = ~pi485 & ~n44754;
  assign n45648 = pi485 & ~n45162;
  assign n45649 = pi248 & ~pi554;
  assign n45650 = ~pi248 & pi554;
  assign n45651 = ~n45649 & ~n45650;
  assign n45652 = ~pi246 & pi563;
  assign n45653 = pi246 & ~pi563;
  assign n45654 = ~n45652 & ~n45653;
  assign n45655 = n45651 & n45654;
  assign n45656 = pi240 & pi551;
  assign n45657 = ~pi240 & ~pi551;
  assign n45658 = ~n45656 & ~n45657;
  assign n45659 = pi249 & ~pi555;
  assign n45660 = ~pi249 & pi555;
  assign n45661 = ~n45659 & ~n45660;
  assign n45662 = pi241 & ~pi553;
  assign n45663 = ~pi241 & pi553;
  assign n45664 = ~n45662 & ~n45663;
  assign n45665 = n45661 & n45664;
  assign n45666 = ~n45658 & n45665;
  assign n45667 = n45655 & n45666;
  assign n45668 = ~n45648 & n45667;
  assign n45669 = ~n45647 & n45668;
  assign n45670 = pi550 & n45669;
  assign n45671 = ~pi239 & ~n45670;
  assign n45672 = ~pi550 & n45669;
  assign n45673 = pi239 & ~n45672;
  assign n45674 = ~n45671 & ~n45673;
  assign n45675 = ~pi489 & n45674;
  assign n45676 = ~pi242 & ~n45675;
  assign n45677 = pi489 & n45674;
  assign n45678 = pi242 & ~n45677;
  assign n45679 = ~n45676 & ~n45678;
  assign n45680 = pi549 & n45679;
  assign n45681 = pi235 & ~n45680;
  assign n45682 = ~pi549 & n45679;
  assign n45683 = ~pi235 & ~n45682;
  assign n45684 = ~n45681 & ~n45683;
  assign n45685 = pi486 & n45684;
  assign n45686 = pi244 & ~n45685;
  assign n45687 = ~pi486 & n45684;
  assign n45688 = ~pi244 & ~n45687;
  assign n45689 = ~n45686 & ~n45688;
  assign n45690 = pi245 & pi580;
  assign n45691 = ~pi245 & ~pi580;
  assign n45692 = ~n45690 & ~n45691;
  assign n45693 = n45689 & ~n45692;
  assign n45694 = pi552 & n45693;
  assign n45695 = pi247 & ~n45694;
  assign n45696 = ~pi552 & n45693;
  assign n45697 = ~pi247 & ~n45696;
  assign n45698 = ~n45695 & ~n45697;
  assign n45699 = ~pi242 & ~pi556;
  assign n45700 = pi242 & pi556;
  assign n45701 = ~n45699 & ~n45700;
  assign n45702 = ~pi570 & ~n44776;
  assign n45703 = pi570 & ~n45218;
  assign n45704 = pi241 & pi562;
  assign n45705 = ~pi241 & ~pi562;
  assign n45706 = ~n45704 & ~n45705;
  assign n45707 = ~pi249 & pi482;
  assign n45708 = ~pi246 & pi564;
  assign n45709 = pi249 & ~pi482;
  assign n45710 = ~n45708 & ~n45709;
  assign n45711 = ~n45707 & n45710;
  assign n45712 = ~n45706 & n45711;
  assign n45713 = ~n45703 & n45712;
  assign n45714 = ~n45702 & n45713;
  assign n45715 = pi240 & pi560;
  assign n45716 = ~pi240 & ~pi560;
  assign n45717 = ~n45715 & ~n45716;
  assign n45718 = pi246 & ~pi564;
  assign n45719 = pi248 & ~pi565;
  assign n45720 = ~pi248 & pi565;
  assign n45721 = ~n45719 & ~n45720;
  assign n45722 = ~n45718 & n45721;
  assign n45723 = ~n45717 & n45722;
  assign n45724 = n45714 & n45723;
  assign n45725 = ~pi239 & pi569;
  assign n45726 = pi239 & ~pi569;
  assign n45727 = ~n45725 & ~n45726;
  assign n45728 = n45724 & ~n45727;
  assign n45729 = ~n45701 & n45728;
  assign n45730 = pi235 & pi531;
  assign n45731 = ~pi235 & ~pi531;
  assign n45732 = ~n45730 & ~n45731;
  assign n45733 = n45729 & ~n45732;
  assign n45734 = pi244 & pi566;
  assign n45735 = ~pi244 & ~pi566;
  assign n45736 = ~n45734 & ~n45735;
  assign n45737 = n45733 & ~n45736;
  assign n45738 = pi568 & n45737;
  assign n45739 = pi245 & ~n45738;
  assign n45740 = ~pi568 & n45737;
  assign n45741 = ~pi245 & ~n45740;
  assign n45742 = ~n45739 & ~n45741;
  assign n45743 = pi247 & pi532;
  assign n45744 = ~pi247 & ~pi532;
  assign n45745 = ~n45743 & ~n45744;
  assign n45746 = n45742 & ~n45745;
  assign n45747 = ~n45698 & ~n45746;
  assign n45748 = ~pi238 & ~n45747;
  assign n45749 = ~pi577 & ~n45748;
  assign n45750 = pi238 & n45698;
  assign n45751 = ~pi238 & n45746;
  assign n45752 = pi577 & ~n45751;
  assign n45753 = ~n45750 & n45752;
  assign n45754 = ~pi498 & ~n45753;
  assign n45755 = ~n45749 & n45754;
  assign n45756 = pi238 & ~n45747;
  assign n45757 = pi577 & ~n45756;
  assign n45758 = ~pi238 & n45698;
  assign n45759 = pi238 & n45746;
  assign n45760 = ~pi577 & ~n45759;
  assign n45761 = ~n45758 & n45760;
  assign n45762 = pi498 & ~n45761;
  assign n45763 = ~n45757 & n45762;
  assign n45764 = ~n45755 & ~n45763;
  assign n45765 = ~pi233 & ~n45764;
  assign n45766 = ~pi237 & ~n45765;
  assign n45767 = ~n45646 & n45766;
  assign po750 = ~n45527 & ~n45767;
  assign n45769 = ~pi806 & n44452;
  assign n45770 = ~pi332 & ~pi806;
  assign n45771 = pi990 & n45770;
  assign n45772 = pi600 & n45771;
  assign n45773 = ~pi332 & pi594;
  assign n45774 = ~n45772 & ~n45773;
  assign po751 = ~n45769 & ~n45774;
  assign n45776 = pi605 & ~pi806;
  assign n45777 = n44435 & n45776;
  assign n45778 = pi595 & n45777;
  assign n45779 = ~pi595 & ~n45777;
  assign n45780 = ~pi332 & ~n45779;
  assign po752 = ~n45778 & n45780;
  assign n45782 = ~pi332 & pi596;
  assign n45783 = pi595 & n44434;
  assign n45784 = n45771 & n45783;
  assign n45785 = ~n45782 & ~n45784;
  assign n45786 = pi596 & n45784;
  assign po753 = ~n45785 & ~n45786;
  assign n45788 = pi597 & n45769;
  assign n45789 = ~pi597 & ~n45769;
  assign n45790 = ~pi332 & ~n45789;
  assign po754 = ~n45788 & n45790;
  assign n45792 = ~pi882 & ~po1038;
  assign n45793 = pi947 & n45792;
  assign n45794 = pi598 & ~n45793;
  assign n45795 = pi740 & pi780;
  assign n45796 = n6157 & n45795;
  assign po755 = n45794 | n45796;
  assign n45798 = ~pi332 & pi599;
  assign n45799 = ~n45786 & ~n45798;
  assign n45800 = pi599 & n45786;
  assign po756 = ~n45799 & ~n45800;
  assign n45802 = ~pi332 & pi600;
  assign n45803 = ~n45771 & ~n45802;
  assign po757 = ~n45772 & ~n45803;
  assign n45805 = ~pi601 & pi806;
  assign n45806 = ~pi806 & ~pi989;
  assign n45807 = ~pi332 & ~n45806;
  assign po758 = ~n45805 & n45807;
  assign n45809 = ~pi230 & pi602;
  assign n45810 = pi230 & n16785;
  assign n45811 = ~n17858 & n45810;
  assign n45812 = pi715 & pi1160;
  assign n45813 = ~pi715 & ~pi1160;
  assign n45814 = pi790 & ~n45813;
  assign n45815 = ~n45812 & n45814;
  assign n45816 = ~n19038 & ~n19182;
  assign n45817 = ~n45815 & n45816;
  assign n45818 = n45811 & n45817;
  assign n45819 = n19128 & n45818;
  assign po759 = n45809 | n45819;
  assign n45821 = ~pi980 & pi1038;
  assign n45822 = pi1060 & n45821;
  assign n45823 = pi952 & ~pi1061;
  assign n45824 = n45822 & n45823;
  assign po897 = pi832 & n45824;
  assign n45826 = ~pi603 & ~po897;
  assign n45827 = pi832 & ~pi1100;
  assign n45828 = n45824 & n45827;
  assign n45829 = ~pi966 & ~n45828;
  assign n45830 = ~n45826 & n45829;
  assign n45831 = pi871 & pi966;
  assign n45832 = pi872 & pi966;
  assign n45833 = ~n45831 & ~n45832;
  assign po760 = n45830 | ~n45833;
  assign n45835 = pi823 & n16512;
  assign n45836 = ~pi779 & n45835;
  assign n45837 = ~pi299 & pi983;
  assign n45838 = pi907 & n45837;
  assign n45839 = pi604 & ~n45838;
  assign n45840 = ~n45835 & n45839;
  assign po761 = n45836 | n45840;
  assign n45842 = ~pi605 & ~n45770;
  assign n45843 = ~pi332 & ~n45776;
  assign po762 = ~n45842 & n45843;
  assign n45845 = ~pi606 & ~po897;
  assign n45846 = ~pi1104 & po897;
  assign n45847 = ~n45845 & ~n45846;
  assign n45848 = ~pi966 & ~n45847;
  assign n45849 = ~pi837 & pi966;
  assign po763 = ~n45848 & ~n45849;
  assign n45851 = ~pi1107 & po897;
  assign n45852 = ~pi607 & ~po897;
  assign n45853 = ~pi966 & ~n45852;
  assign po764 = ~n45851 & n45853;
  assign n45855 = ~pi1116 & po897;
  assign n45856 = ~pi608 & ~po897;
  assign n45857 = ~pi966 & ~n45856;
  assign po765 = ~n45855 & n45857;
  assign n45859 = ~pi1118 & po897;
  assign n45860 = ~pi609 & ~po897;
  assign n45861 = ~pi966 & ~n45860;
  assign po766 = ~n45859 & n45861;
  assign n45863 = ~pi1113 & po897;
  assign n45864 = ~pi610 & ~po897;
  assign n45865 = ~pi966 & ~n45864;
  assign po767 = ~n45863 & n45865;
  assign n45867 = ~pi1114 & po897;
  assign n45868 = ~pi611 & ~po897;
  assign n45869 = ~pi966 & ~n45868;
  assign po768 = ~n45867 & n45869;
  assign n45871 = ~pi1111 & po897;
  assign n45872 = ~pi612 & ~po897;
  assign n45873 = ~pi966 & ~n45872;
  assign po769 = ~n45871 & n45873;
  assign n45875 = ~pi1115 & po897;
  assign n45876 = ~pi613 & ~po897;
  assign n45877 = ~pi966 & ~n45876;
  assign po770 = ~n45875 & n45877;
  assign n45879 = ~pi1102 & po897;
  assign n45880 = ~pi614 & ~po897;
  assign n45881 = ~pi966 & ~n45880;
  assign n45882 = ~n45879 & n45881;
  assign po771 = n45831 | n45882;
  assign n45884 = pi907 & n45792;
  assign n45885 = ~pi615 & ~n45884;
  assign n45886 = pi779 & pi797;
  assign n45887 = n6160 & n45886;
  assign po772 = n45885 | n45887;
  assign n45889 = ~pi1101 & po897;
  assign n45890 = ~pi616 & ~po897;
  assign n45891 = ~pi966 & ~n45890;
  assign n45892 = ~n45889 & n45891;
  assign po773 = n45832 | n45892;
  assign n45894 = ~pi617 & ~po897;
  assign n45895 = ~pi1105 & po897;
  assign n45896 = ~n45894 & ~n45895;
  assign n45897 = ~pi966 & ~n45896;
  assign n45898 = ~pi850 & pi966;
  assign po774 = ~n45897 & ~n45898;
  assign n45900 = ~pi1117 & po897;
  assign n45901 = ~pi618 & ~po897;
  assign n45902 = ~pi966 & ~n45901;
  assign po775 = ~n45900 & n45902;
  assign n45904 = ~pi1122 & po897;
  assign n45905 = ~pi619 & ~po897;
  assign n45906 = ~pi966 & ~n45905;
  assign po776 = ~n45904 & n45906;
  assign n45908 = ~pi1112 & po897;
  assign n45909 = ~pi620 & ~po897;
  assign n45910 = ~pi966 & ~n45909;
  assign po777 = ~n45908 & n45910;
  assign n45912 = ~pi1108 & po897;
  assign n45913 = ~pi621 & ~po897;
  assign n45914 = ~pi966 & ~n45913;
  assign po778 = ~n45912 & n45914;
  assign n45916 = ~pi1109 & po897;
  assign n45917 = ~pi622 & ~po897;
  assign n45918 = ~pi966 & ~n45917;
  assign po779 = ~n45916 & n45918;
  assign n45920 = ~pi1106 & po897;
  assign n45921 = ~pi623 & ~po897;
  assign n45922 = ~pi966 & ~n45921;
  assign po780 = ~n45920 & n45922;
  assign n45924 = pi831 & n16592;
  assign n45925 = ~pi780 & n45924;
  assign n45926 = pi947 & n45837;
  assign n45927 = pi624 & ~n45926;
  assign n45928 = ~n45924 & n45927;
  assign po781 = n45925 | n45928;
  assign n45930 = pi832 & ~pi973;
  assign n45931 = ~pi1054 & pi1066;
  assign n45932 = pi1088 & n45931;
  assign n45933 = n45930 & n45932;
  assign po954 = ~pi953 & n45933;
  assign n45935 = ~pi1116 & po954;
  assign n45936 = ~pi625 & ~po954;
  assign n45937 = ~pi962 & ~n45936;
  assign po782 = ~n45935 & n45937;
  assign n45939 = ~pi1121 & po897;
  assign n45940 = ~pi626 & ~po897;
  assign n45941 = ~pi966 & ~n45940;
  assign po783 = ~n45939 & n45941;
  assign n45943 = ~pi1117 & po954;
  assign n45944 = ~pi627 & ~po954;
  assign n45945 = ~pi962 & ~n45944;
  assign po784 = ~n45943 & n45945;
  assign n45947 = ~pi1119 & po954;
  assign n45948 = ~pi628 & ~po954;
  assign n45949 = ~pi962 & ~n45948;
  assign po785 = ~n45947 & n45949;
  assign n45951 = ~pi1119 & po897;
  assign n45952 = ~pi629 & ~po897;
  assign n45953 = ~pi966 & ~n45952;
  assign po786 = ~n45951 & n45953;
  assign n45955 = ~pi1120 & po897;
  assign n45956 = ~pi630 & ~po897;
  assign n45957 = ~pi966 & ~n45956;
  assign po787 = ~n45955 & n45957;
  assign n45959 = pi631 & ~po954;
  assign n45960 = ~pi1113 & po954;
  assign n45961 = ~pi962 & ~n45960;
  assign po788 = ~n45959 & n45961;
  assign n45963 = pi632 & ~po954;
  assign n45964 = ~pi1115 & po954;
  assign n45965 = ~pi962 & ~n45964;
  assign po789 = ~n45963 & n45965;
  assign n45967 = ~pi1110 & po897;
  assign n45968 = ~pi633 & ~po897;
  assign n45969 = ~pi966 & ~n45968;
  assign po790 = ~n45967 & n45969;
  assign n45971 = ~pi1110 & po954;
  assign n45972 = ~pi634 & ~po954;
  assign n45973 = ~pi962 & ~n45972;
  assign po791 = ~n45971 & n45973;
  assign n45975 = pi635 & ~po954;
  assign n45976 = ~pi1112 & po954;
  assign n45977 = ~pi962 & ~n45976;
  assign po792 = ~n45975 & n45977;
  assign n45979 = ~pi1127 & po897;
  assign n45980 = ~pi636 & ~po897;
  assign n45981 = ~pi966 & ~n45980;
  assign po793 = ~n45979 & n45981;
  assign n45983 = ~pi1105 & po954;
  assign n45984 = ~pi637 & ~po954;
  assign n45985 = ~pi962 & ~n45984;
  assign po794 = ~n45983 & n45985;
  assign n45987 = ~pi1107 & po954;
  assign n45988 = ~pi638 & ~po954;
  assign n45989 = ~pi962 & ~n45988;
  assign po795 = ~n45987 & n45989;
  assign n45991 = ~pi1109 & po954;
  assign n45992 = ~pi639 & ~po954;
  assign n45993 = ~pi962 & ~n45992;
  assign po796 = ~n45991 & n45993;
  assign n45995 = ~pi1128 & po897;
  assign n45996 = ~pi640 & ~po897;
  assign n45997 = ~pi966 & ~n45996;
  assign po797 = ~n45995 & n45997;
  assign n45999 = ~pi1121 & po954;
  assign n46000 = ~pi641 & ~po954;
  assign n46001 = ~pi962 & ~n46000;
  assign po798 = ~n45999 & n46001;
  assign n46003 = ~pi1103 & po897;
  assign n46004 = ~pi642 & ~po897;
  assign n46005 = ~pi966 & ~n46004;
  assign po799 = ~n46003 & n46005;
  assign n46007 = ~pi1104 & po954;
  assign n46008 = ~pi643 & ~po954;
  assign n46009 = ~pi962 & ~n46008;
  assign po800 = ~n46007 & n46009;
  assign n46011 = ~pi1123 & po897;
  assign n46012 = ~pi644 & ~po897;
  assign n46013 = ~pi966 & ~n46012;
  assign po801 = ~n46011 & n46013;
  assign n46015 = ~pi1125 & po897;
  assign n46016 = ~pi645 & ~po897;
  assign n46017 = ~pi966 & ~n46016;
  assign po802 = ~n46015 & n46017;
  assign n46019 = pi646 & ~po954;
  assign n46020 = ~pi1114 & po954;
  assign n46021 = ~pi962 & ~n46020;
  assign po803 = ~n46019 & n46021;
  assign n46023 = ~pi1120 & po954;
  assign n46024 = ~pi647 & ~po954;
  assign n46025 = ~pi962 & ~n46024;
  assign po804 = ~n46023 & n46025;
  assign n46027 = ~pi1122 & po954;
  assign n46028 = ~pi648 & ~po954;
  assign n46029 = ~pi962 & ~n46028;
  assign po805 = ~n46027 & n46029;
  assign n46031 = pi649 & ~po954;
  assign n46032 = ~pi1126 & po954;
  assign n46033 = ~pi962 & ~n46032;
  assign po806 = ~n46031 & n46033;
  assign n46035 = pi650 & ~po954;
  assign n46036 = ~pi1127 & po954;
  assign n46037 = ~pi962 & ~n46036;
  assign po807 = ~n46035 & n46037;
  assign n46039 = ~pi1130 & po897;
  assign n46040 = ~pi651 & ~po897;
  assign n46041 = ~pi966 & ~n46040;
  assign po808 = ~n46039 & n46041;
  assign n46043 = ~pi1131 & po897;
  assign n46044 = ~pi652 & ~po897;
  assign n46045 = ~pi966 & ~n46044;
  assign po809 = ~n46043 & n46045;
  assign n46047 = ~pi1129 & po897;
  assign n46048 = ~pi653 & ~po897;
  assign n46049 = ~pi966 & ~n46048;
  assign po810 = ~n46047 & n46049;
  assign n46051 = pi654 & ~po954;
  assign n46052 = ~pi1130 & po954;
  assign n46053 = ~pi962 & ~n46052;
  assign po811 = ~n46051 & n46053;
  assign n46055 = pi655 & ~po954;
  assign n46056 = ~pi1124 & po954;
  assign n46057 = ~pi962 & ~n46056;
  assign po812 = ~n46055 & n46057;
  assign n46059 = ~pi1126 & po897;
  assign n46060 = ~pi656 & ~po897;
  assign n46061 = ~pi966 & ~n46060;
  assign po813 = ~n46059 & n46061;
  assign n46063 = pi657 & ~po954;
  assign n46064 = ~pi1131 & po954;
  assign n46065 = ~pi962 & ~n46064;
  assign po814 = ~n46063 & n46065;
  assign n46067 = ~pi1124 & po897;
  assign n46068 = ~pi658 & ~po897;
  assign n46069 = ~pi966 & ~n46068;
  assign po815 = ~n46067 & n46069;
  assign n46071 = pi266 & pi992;
  assign n46072 = ~pi280 & n46071;
  assign n46073 = ~pi269 & n46072;
  assign n46074 = ~pi281 & n46073;
  assign n46075 = ~pi270 & ~pi277;
  assign n46076 = ~pi282 & n46075;
  assign n46077 = n46074 & n46076;
  assign n46078 = ~pi264 & n46077;
  assign n46079 = ~pi265 & n46078;
  assign po959 = ~pi274 & n46079;
  assign n46081 = pi274 & ~n46079;
  assign po816 = ~po959 & ~n46081;
  assign n46083 = ~pi1118 & po954;
  assign n46084 = ~pi660 & ~po954;
  assign n46085 = ~pi962 & ~n46084;
  assign po817 = ~n46083 & n46085;
  assign n46087 = ~pi1101 & po954;
  assign n46088 = ~pi661 & ~po954;
  assign n46089 = ~pi962 & ~n46088;
  assign po818 = ~n46087 & n46089;
  assign n46091 = ~pi1102 & po954;
  assign n46092 = ~pi662 & ~po954;
  assign n46093 = ~pi962 & ~n46092;
  assign po819 = ~n46091 & n46093;
  assign n46095 = pi199 & ~pi1065;
  assign n46096 = ~pi223 & ~pi224;
  assign n46097 = ~pi199 & ~pi257;
  assign n46098 = ~n46096 & ~n46097;
  assign n46099 = ~n46095 & n46098;
  assign n46100 = ~pi591 & pi592;
  assign n46101 = pi365 & n46100;
  assign n46102 = pi334 & pi591;
  assign n46103 = ~pi592 & n46102;
  assign n46104 = ~n46101 & ~n46103;
  assign n46105 = ~pi590 & ~n46104;
  assign n46106 = ~pi591 & ~pi592;
  assign n46107 = pi590 & n46106;
  assign n46108 = pi323 & n46107;
  assign n46109 = ~pi588 & ~n46108;
  assign n46110 = ~n46105 & n46109;
  assign n46111 = ~pi592 & n8558;
  assign n46112 = pi464 & n46111;
  assign n46113 = pi588 & ~n46112;
  assign n46114 = n46096 & ~n46113;
  assign n46115 = ~n46110 & n46114;
  assign n46116 = ~n46099 & ~n46115;
  assign n46117 = n8830 & ~n46116;
  assign n46118 = ~pi1137 & ~pi1138;
  assign n46119 = ~pi1134 & n46118;
  assign n46120 = ~pi634 & pi1136;
  assign n46121 = ~pi784 & ~pi1136;
  assign n46122 = pi1135 & ~n46121;
  assign n46123 = ~n46120 & n46122;
  assign n46124 = ~pi633 & pi1136;
  assign n46125 = ~pi815 & ~pi1136;
  assign n46126 = ~pi1135 & ~n46125;
  assign n46127 = ~n46124 & n46126;
  assign n46128 = ~n46123 & ~n46127;
  assign n46129 = n46119 & ~n46128;
  assign n46130 = pi1135 & n46118;
  assign n46131 = pi1136 & ~n46130;
  assign n46132 = ~pi766 & n46131;
  assign n46133 = pi1135 & ~pi1136;
  assign n46134 = pi1134 & n46118;
  assign n46135 = ~n46133 & n46134;
  assign n46136 = ~pi855 & ~pi1136;
  assign n46137 = ~pi700 & pi1135;
  assign n46138 = ~n46136 & ~n46137;
  assign n46139 = n46135 & n46138;
  assign n46140 = ~n46132 & n46139;
  assign n46141 = ~n46129 & ~n46140;
  assign n46142 = ~n8830 & ~n46141;
  assign po820 = n46117 | n46142;
  assign n46144 = ~pi590 & pi591;
  assign n46145 = pi404 & n46144;
  assign n46146 = ~pi590 & pi592;
  assign n46147 = ~pi588 & ~n46146;
  assign n46148 = ~n46145 & n46147;
  assign n46149 = pi380 & ~pi591;
  assign n46150 = pi592 & ~n46149;
  assign n46151 = ~n46148 & ~n46150;
  assign n46152 = pi355 & n46107;
  assign n46153 = ~n46151 & ~n46152;
  assign n46154 = pi429 & n46111;
  assign n46155 = pi588 & ~n46154;
  assign n46156 = n46096 & ~n46155;
  assign n46157 = ~n46153 & n46156;
  assign n46158 = pi199 & ~pi1084;
  assign n46159 = ~pi199 & ~pi292;
  assign n46160 = ~n46096 & ~n46159;
  assign n46161 = ~n46158 & n46160;
  assign n46162 = ~n46157 & ~n46161;
  assign n46163 = n8830 & ~n46162;
  assign n46164 = pi662 & pi1135;
  assign n46165 = pi614 & ~pi1135;
  assign n46166 = pi1136 & ~n46165;
  assign n46167 = ~n46164 & n46166;
  assign n46168 = pi785 & pi1135;
  assign n46169 = pi811 & ~pi1135;
  assign n46170 = ~pi1136 & ~n46169;
  assign n46171 = ~n46168 & n46170;
  assign n46172 = ~n46167 & ~n46171;
  assign n46173 = ~pi1134 & ~n46172;
  assign n46174 = ~pi727 & pi1135;
  assign n46175 = ~pi772 & ~pi1135;
  assign n46176 = pi1136 & ~n46175;
  assign n46177 = ~n46174 & n46176;
  assign n46178 = ~pi1135 & ~pi1136;
  assign n46179 = pi872 & n46178;
  assign n46180 = pi1134 & ~n46179;
  assign n46181 = ~n46177 & n46180;
  assign n46182 = ~n8830 & n46118;
  assign n46183 = ~n46181 & n46182;
  assign n46184 = ~n46173 & n46183;
  assign po821 = n46163 | n46184;
  assign n46186 = ~pi1108 & po954;
  assign n46187 = ~pi665 & ~po954;
  assign n46188 = ~pi962 & ~n46187;
  assign po822 = ~n46186 & n46188;
  assign n46190 = ~pi638 & pi1135;
  assign n46191 = ~pi607 & ~pi1135;
  assign n46192 = pi1136 & ~n46191;
  assign n46193 = ~n46190 & n46192;
  assign n46194 = pi799 & ~pi1135;
  assign n46195 = ~pi790 & pi1135;
  assign n46196 = ~pi1136 & ~n46195;
  assign n46197 = ~n46194 & n46196;
  assign n46198 = ~n46193 & ~n46197;
  assign n46199 = n46119 & ~n46198;
  assign n46200 = ~pi764 & n46131;
  assign n46201 = ~pi691 & pi1135;
  assign n46202 = ~pi873 & ~pi1136;
  assign n46203 = ~n46201 & ~n46202;
  assign n46204 = n46135 & n46203;
  assign n46205 = ~n46200 & n46204;
  assign n46206 = ~n46199 & ~n46205;
  assign n46207 = ~n8830 & ~n46206;
  assign n46208 = pi199 & ~pi1044;
  assign n46209 = ~pi199 & ~pi297;
  assign n46210 = ~n46096 & ~n46209;
  assign n46211 = ~n46208 & n46210;
  assign n46212 = pi456 & n46144;
  assign n46213 = n46147 & ~n46212;
  assign n46214 = pi337 & ~pi591;
  assign n46215 = pi592 & ~n46214;
  assign n46216 = ~n46213 & ~n46215;
  assign n46217 = pi441 & n46107;
  assign n46218 = ~n46216 & ~n46217;
  assign n46219 = pi443 & n46111;
  assign n46220 = pi588 & ~n46219;
  assign n46221 = n46096 & ~n46220;
  assign n46222 = ~n46218 & n46221;
  assign n46223 = ~n46211 & ~n46222;
  assign n46224 = n8830 & ~n46223;
  assign po823 = n46207 | n46224;
  assign n46226 = pi319 & n46144;
  assign n46227 = n46147 & ~n46226;
  assign n46228 = pi338 & ~pi591;
  assign n46229 = pi592 & ~n46228;
  assign n46230 = ~n46227 & ~n46229;
  assign n46231 = pi458 & n46107;
  assign n46232 = ~n46230 & ~n46231;
  assign n46233 = pi444 & n46111;
  assign n46234 = pi588 & ~n46233;
  assign n46235 = n46096 & ~n46234;
  assign n46236 = ~n46232 & n46235;
  assign n46237 = pi199 & ~pi1072;
  assign n46238 = ~pi199 & ~pi294;
  assign n46239 = ~n46096 & ~n46238;
  assign n46240 = ~n46237 & n46239;
  assign n46241 = ~n46236 & ~n46240;
  assign n46242 = n8830 & ~n46241;
  assign n46243 = pi681 & pi1136;
  assign n46244 = pi792 & ~pi1136;
  assign n46245 = pi1135 & ~n46244;
  assign n46246 = ~n46243 & n46245;
  assign n46247 = pi642 & pi1136;
  assign n46248 = ~pi809 & ~pi1136;
  assign n46249 = ~pi1135 & ~n46248;
  assign n46250 = ~n46247 & n46249;
  assign n46251 = ~n46246 & ~n46250;
  assign n46252 = ~pi1134 & ~n46251;
  assign n46253 = ~pi699 & pi1135;
  assign n46254 = ~pi763 & ~pi1135;
  assign n46255 = pi1136 & ~n46254;
  assign n46256 = ~n46253 & n46255;
  assign n46257 = pi871 & n46178;
  assign n46258 = pi1134 & ~n46257;
  assign n46259 = ~n46256 & n46258;
  assign n46260 = n46182 & ~n46259;
  assign n46261 = ~n46252 & n46260;
  assign po824 = n46242 | n46261;
  assign n46263 = ~pi680 & pi1135;
  assign n46264 = ~pi603 & ~pi1135;
  assign n46265 = pi1136 & ~n46264;
  assign n46266 = ~n46263 & n46265;
  assign n46267 = ~pi778 & pi1135;
  assign n46268 = ~pi981 & ~pi1135;
  assign n46269 = ~pi1136 & ~n46268;
  assign n46270 = ~n46267 & n46269;
  assign n46271 = ~n46266 & ~n46270;
  assign n46272 = n46119 & ~n46271;
  assign n46273 = ~pi759 & n46131;
  assign n46274 = ~pi696 & pi1135;
  assign n46275 = ~pi837 & ~pi1136;
  assign n46276 = ~n46274 & ~n46275;
  assign n46277 = n46135 & n46276;
  assign n46278 = ~n46273 & n46277;
  assign n46279 = ~n46272 & ~n46278;
  assign n46280 = ~n8830 & ~n46279;
  assign n46281 = pi199 & ~pi1049;
  assign n46282 = ~pi199 & ~pi291;
  assign n46283 = ~n46096 & ~n46282;
  assign n46284 = ~n46281 & n46283;
  assign n46285 = pi390 & n46144;
  assign n46286 = n46147 & ~n46285;
  assign n46287 = pi363 & ~pi591;
  assign n46288 = pi592 & ~n46287;
  assign n46289 = ~n46286 & ~n46288;
  assign n46290 = pi342 & n46107;
  assign n46291 = ~n46289 & ~n46290;
  assign n46292 = pi414 & n46111;
  assign n46293 = pi588 & ~n46292;
  assign n46294 = n46096 & ~n46293;
  assign n46295 = ~n46291 & n46294;
  assign n46296 = ~n46284 & ~n46295;
  assign n46297 = n8830 & ~n46296;
  assign po825 = n46280 | n46297;
  assign n46299 = pi669 & ~po954;
  assign n46300 = ~pi1125 & po954;
  assign n46301 = ~pi962 & ~n46300;
  assign po826 = ~n46299 & n46301;
  assign n46303 = pi199 & ~pi1062;
  assign n46304 = ~pi199 & ~pi258;
  assign n46305 = ~n46096 & ~n46304;
  assign n46306 = ~n46303 & n46305;
  assign n46307 = pi364 & n46100;
  assign n46308 = pi391 & pi591;
  assign n46309 = ~pi592 & n46308;
  assign n46310 = ~n46307 & ~n46309;
  assign n46311 = ~pi590 & ~n46310;
  assign n46312 = pi343 & n46107;
  assign n46313 = ~pi588 & ~n46312;
  assign n46314 = ~n46311 & n46313;
  assign n46315 = pi415 & n46111;
  assign n46316 = pi588 & ~n46315;
  assign n46317 = n46096 & ~n46316;
  assign n46318 = ~n46314 & n46317;
  assign n46319 = ~n46306 & ~n46318;
  assign n46320 = n8830 & ~n46319;
  assign n46321 = pi745 & n46131;
  assign n46322 = pi723 & pi1135;
  assign n46323 = ~pi852 & ~pi1136;
  assign n46324 = ~n46322 & ~n46323;
  assign n46325 = n46135 & n46324;
  assign n46326 = ~n46321 & n46325;
  assign n46327 = pi1136 & n46118;
  assign n46328 = ~pi612 & ~pi1135;
  assign n46329 = pi695 & pi1135;
  assign n46330 = ~pi1134 & ~n46329;
  assign n46331 = ~n46328 & n46330;
  assign n46332 = n46327 & n46331;
  assign n46333 = ~n46326 & ~n46332;
  assign n46334 = ~n8830 & ~n46333;
  assign po827 = n46320 | n46334;
  assign n46336 = pi199 & ~pi1040;
  assign n46337 = ~pi199 & ~pi261;
  assign n46338 = ~n46096 & ~n46337;
  assign n46339 = ~n46336 & n46338;
  assign n46340 = pi447 & n46100;
  assign n46341 = pi333 & pi591;
  assign n46342 = ~pi592 & n46341;
  assign n46343 = ~n46340 & ~n46342;
  assign n46344 = ~pi590 & ~n46343;
  assign n46345 = pi327 & n46107;
  assign n46346 = ~pi588 & ~n46345;
  assign n46347 = ~n46344 & n46346;
  assign n46348 = pi453 & n46111;
  assign n46349 = pi588 & ~n46348;
  assign n46350 = n46096 & ~n46349;
  assign n46351 = ~n46347 & n46350;
  assign n46352 = ~n46339 & ~n46351;
  assign n46353 = n8830 & ~n46352;
  assign n46354 = pi741 & n46131;
  assign n46355 = pi724 & pi1135;
  assign n46356 = ~pi865 & ~pi1136;
  assign n46357 = ~n46355 & ~n46356;
  assign n46358 = n46135 & n46357;
  assign n46359 = ~n46354 & n46358;
  assign n46360 = ~pi611 & ~pi1135;
  assign n46361 = pi646 & pi1135;
  assign n46362 = ~pi1134 & ~n46361;
  assign n46363 = ~n46360 & n46362;
  assign n46364 = n46327 & n46363;
  assign n46365 = ~n46359 & ~n46364;
  assign n46366 = ~n8830 & ~n46365;
  assign po828 = n46353 | n46366;
  assign n46368 = ~pi661 & pi1135;
  assign n46369 = ~pi616 & ~pi1135;
  assign n46370 = pi1136 & ~n46369;
  assign n46371 = ~n46368 & n46370;
  assign n46372 = ~pi781 & pi1135;
  assign n46373 = ~pi808 & ~pi1135;
  assign n46374 = ~pi1136 & ~n46373;
  assign n46375 = ~n46372 & n46374;
  assign n46376 = ~n46371 & ~n46375;
  assign n46377 = n46119 & ~n46376;
  assign n46378 = ~pi758 & n46131;
  assign n46379 = ~pi736 & pi1135;
  assign n46380 = ~pi850 & ~pi1136;
  assign n46381 = ~n46379 & ~n46380;
  assign n46382 = n46135 & n46381;
  assign n46383 = ~n46378 & n46382;
  assign n46384 = ~n46377 & ~n46383;
  assign n46385 = ~n8830 & ~n46384;
  assign n46386 = pi199 & ~pi1048;
  assign n46387 = ~pi199 & ~pi290;
  assign n46388 = ~n46096 & ~n46387;
  assign n46389 = ~n46386 & n46388;
  assign n46390 = pi397 & n46144;
  assign n46391 = n46147 & ~n46390;
  assign n46392 = pi372 & ~pi591;
  assign n46393 = pi592 & ~n46392;
  assign n46394 = ~n46391 & ~n46393;
  assign n46395 = pi320 & n46107;
  assign n46396 = ~n46394 & ~n46395;
  assign n46397 = pi422 & n46111;
  assign n46398 = pi588 & ~n46397;
  assign n46399 = n46096 & ~n46398;
  assign n46400 = ~n46396 & n46399;
  assign n46401 = ~n46389 & ~n46400;
  assign n46402 = n8830 & ~n46401;
  assign po829 = n46385 | n46402;
  assign n46404 = ~pi637 & pi1135;
  assign n46405 = ~pi617 & ~pi1135;
  assign n46406 = pi1136 & ~n46405;
  assign n46407 = ~n46404 & n46406;
  assign n46408 = pi814 & ~pi1135;
  assign n46409 = ~pi788 & pi1135;
  assign n46410 = ~pi1136 & ~n46409;
  assign n46411 = ~n46408 & n46410;
  assign n46412 = ~n46407 & ~n46411;
  assign n46413 = n46119 & ~n46412;
  assign n46414 = ~pi749 & n46131;
  assign n46415 = ~pi706 & pi1135;
  assign n46416 = ~pi866 & ~pi1136;
  assign n46417 = ~n46415 & ~n46416;
  assign n46418 = n46135 & n46417;
  assign n46419 = ~n46414 & n46418;
  assign n46420 = ~n46413 & ~n46419;
  assign n46421 = ~n8830 & ~n46420;
  assign n46422 = pi199 & ~pi1053;
  assign n46423 = ~pi199 & ~pi295;
  assign n46424 = ~n46096 & ~n46423;
  assign n46425 = ~n46422 & n46424;
  assign n46426 = pi411 & n46144;
  assign n46427 = n46147 & ~n46426;
  assign n46428 = pi387 & ~pi591;
  assign n46429 = pi592 & ~n46428;
  assign n46430 = ~n46427 & ~n46429;
  assign n46431 = pi452 & n46107;
  assign n46432 = ~n46430 & ~n46431;
  assign n46433 = pi435 & n46111;
  assign n46434 = pi588 & ~n46433;
  assign n46435 = n46096 & ~n46434;
  assign n46436 = ~n46432 & n46435;
  assign n46437 = ~n46425 & ~n46436;
  assign n46438 = n8830 & ~n46437;
  assign po830 = n46421 | n46438;
  assign n46440 = pi199 & ~pi1070;
  assign n46441 = ~pi199 & ~pi256;
  assign n46442 = ~n46096 & ~n46441;
  assign n46443 = ~n46440 & n46442;
  assign n46444 = pi336 & n46100;
  assign n46445 = pi463 & pi591;
  assign n46446 = ~pi592 & n46445;
  assign n46447 = ~n46444 & ~n46446;
  assign n46448 = ~pi590 & ~n46447;
  assign n46449 = pi362 & n46107;
  assign n46450 = ~pi588 & ~n46449;
  assign n46451 = ~n46448 & n46450;
  assign n46452 = pi437 & n46111;
  assign n46453 = pi588 & ~n46452;
  assign n46454 = n46096 & ~n46453;
  assign n46455 = ~n46451 & n46454;
  assign n46456 = ~n46443 & ~n46455;
  assign n46457 = n8830 & ~n46456;
  assign n46458 = pi639 & pi1135;
  assign n46459 = pi622 & ~pi1135;
  assign n46460 = pi1136 & ~n46459;
  assign n46461 = ~n46458 & n46460;
  assign n46462 = pi783 & pi1135;
  assign n46463 = pi804 & ~pi1135;
  assign n46464 = ~pi1136 & ~n46463;
  assign n46465 = ~n46462 & n46464;
  assign n46466 = ~n46461 & ~n46465;
  assign n46467 = ~pi1134 & ~n46466;
  assign n46468 = ~pi735 & pi1135;
  assign n46469 = ~pi743 & ~pi1135;
  assign n46470 = pi1136 & ~n46469;
  assign n46471 = ~n46468 & n46470;
  assign n46472 = pi859 & n46178;
  assign n46473 = pi1134 & ~n46472;
  assign n46474 = ~n46471 & n46473;
  assign n46475 = n46182 & ~n46474;
  assign n46476 = ~n46467 & n46475;
  assign po831 = n46457 | n46476;
  assign n46478 = pi876 & n46178;
  assign n46479 = ~pi730 & pi1135;
  assign n46480 = ~pi748 & ~pi1135;
  assign n46481 = pi1136 & ~n46480;
  assign n46482 = ~n46479 & n46481;
  assign n46483 = ~n46478 & ~n46482;
  assign n46484 = n46134 & ~n46483;
  assign n46485 = ~pi710 & pi1135;
  assign n46486 = pi1136 & ~n46485;
  assign n46487 = pi789 & n46133;
  assign n46488 = ~pi803 & ~pi1135;
  assign n46489 = ~n46487 & ~n46488;
  assign n46490 = ~n46486 & n46489;
  assign n46491 = ~pi623 & n46131;
  assign n46492 = n46119 & ~n46491;
  assign n46493 = ~n46490 & n46492;
  assign n46494 = ~n46484 & ~n46493;
  assign n46495 = ~n8830 & ~n46494;
  assign n46496 = pi199 & ~pi1037;
  assign n46497 = ~pi199 & ~pi296;
  assign n46498 = ~n46096 & ~n46497;
  assign n46499 = ~n46496 & n46498;
  assign n46500 = pi412 & n46144;
  assign n46501 = n46147 & ~n46500;
  assign n46502 = pi388 & ~pi591;
  assign n46503 = pi592 & ~n46502;
  assign n46504 = ~n46501 & ~n46503;
  assign n46505 = pi455 & n46107;
  assign n46506 = ~n46504 & ~n46505;
  assign n46507 = pi436 & n46111;
  assign n46508 = pi588 & ~n46507;
  assign n46509 = n46096 & ~n46508;
  assign n46510 = ~n46506 & n46509;
  assign n46511 = ~n46499 & ~n46510;
  assign n46512 = n8830 & ~n46511;
  assign po832 = n46495 | n46512;
  assign n46514 = ~pi643 & pi1135;
  assign n46515 = ~pi606 & ~pi1135;
  assign n46516 = pi1136 & ~n46515;
  assign n46517 = ~n46514 & n46516;
  assign n46518 = pi812 & ~pi1135;
  assign n46519 = ~pi787 & pi1135;
  assign n46520 = ~pi1136 & ~n46519;
  assign n46521 = ~n46518 & n46520;
  assign n46522 = ~n46517 & ~n46521;
  assign n46523 = n46119 & ~n46522;
  assign n46524 = ~pi746 & n46131;
  assign n46525 = ~pi729 & pi1135;
  assign n46526 = ~pi881 & ~pi1136;
  assign n46527 = ~n46525 & ~n46526;
  assign n46528 = n46135 & n46527;
  assign n46529 = ~n46524 & n46528;
  assign n46530 = ~n46523 & ~n46529;
  assign n46531 = ~n8830 & ~n46530;
  assign n46532 = pi199 & ~pi1059;
  assign n46533 = ~pi199 & ~pi293;
  assign n46534 = ~n46096 & ~n46533;
  assign n46535 = ~n46532 & n46534;
  assign n46536 = pi410 & n46144;
  assign n46537 = n46147 & ~n46536;
  assign n46538 = pi386 & ~pi591;
  assign n46539 = pi592 & ~n46538;
  assign n46540 = ~n46537 & ~n46539;
  assign n46541 = pi361 & n46107;
  assign n46542 = ~n46540 & ~n46541;
  assign n46543 = pi434 & n46111;
  assign n46544 = pi588 & ~n46543;
  assign n46545 = n46096 & ~n46544;
  assign n46546 = ~n46542 & n46545;
  assign n46547 = ~n46535 & ~n46546;
  assign n46548 = n8830 & ~n46547;
  assign po833 = n46531 | n46548;
  assign n46550 = pi199 & ~pi1069;
  assign n46551 = ~pi199 & ~pi259;
  assign n46552 = ~n46096 & ~n46551;
  assign n46553 = ~n46550 & n46552;
  assign n46554 = pi366 & n46100;
  assign n46555 = pi335 & pi591;
  assign n46556 = ~pi592 & n46555;
  assign n46557 = ~n46554 & ~n46556;
  assign n46558 = ~pi590 & ~n46557;
  assign n46559 = pi344 & n46107;
  assign n46560 = ~pi588 & ~n46559;
  assign n46561 = ~n46558 & n46560;
  assign n46562 = pi416 & n46111;
  assign n46563 = pi588 & ~n46562;
  assign n46564 = n46096 & ~n46563;
  assign n46565 = ~n46561 & n46564;
  assign n46566 = ~n46553 & ~n46565;
  assign n46567 = n8830 & ~n46566;
  assign n46568 = pi742 & n46131;
  assign n46569 = pi704 & pi1135;
  assign n46570 = ~pi870 & ~pi1136;
  assign n46571 = ~n46569 & ~n46570;
  assign n46572 = n46135 & n46571;
  assign n46573 = ~n46568 & n46572;
  assign n46574 = ~pi620 & ~pi1135;
  assign n46575 = pi635 & pi1135;
  assign n46576 = ~pi1134 & ~n46575;
  assign n46577 = ~n46574 & n46576;
  assign n46578 = n46327 & n46577;
  assign n46579 = ~n46573 & ~n46578;
  assign n46580 = ~n8830 & ~n46579;
  assign po834 = n46567 | n46580;
  assign n46582 = pi199 & ~pi1067;
  assign n46583 = ~pi199 & ~pi260;
  assign n46584 = ~n46096 & ~n46583;
  assign n46585 = ~n46582 & n46584;
  assign n46586 = pi368 & n46100;
  assign n46587 = pi393 & pi591;
  assign n46588 = ~pi592 & n46587;
  assign n46589 = ~n46586 & ~n46588;
  assign n46590 = ~pi590 & ~n46589;
  assign n46591 = pi346 & n46107;
  assign n46592 = ~pi588 & ~n46591;
  assign n46593 = ~n46590 & n46592;
  assign n46594 = pi418 & n46111;
  assign n46595 = pi588 & ~n46594;
  assign n46596 = n46096 & ~n46595;
  assign n46597 = ~n46593 & n46596;
  assign n46598 = ~n46585 & ~n46597;
  assign n46599 = n8830 & ~n46598;
  assign n46600 = pi760 & n46131;
  assign n46601 = pi688 & pi1135;
  assign n46602 = ~pi856 & ~pi1136;
  assign n46603 = ~n46601 & ~n46602;
  assign n46604 = n46135 & n46603;
  assign n46605 = ~n46600 & n46604;
  assign n46606 = ~pi613 & ~pi1135;
  assign n46607 = pi632 & pi1135;
  assign n46608 = ~pi1134 & ~n46607;
  assign n46609 = ~n46606 & n46608;
  assign n46610 = n46327 & n46609;
  assign n46611 = ~n46605 & ~n46610;
  assign n46612 = ~n8830 & ~n46611;
  assign po835 = n46599 | n46612;
  assign n46614 = pi199 & ~pi1036;
  assign n46615 = ~pi199 & ~pi255;
  assign n46616 = ~n46096 & ~n46615;
  assign n46617 = ~n46614 & n46616;
  assign n46618 = pi389 & n46100;
  assign n46619 = pi413 & pi591;
  assign n46620 = ~pi592 & n46619;
  assign n46621 = ~n46618 & ~n46620;
  assign n46622 = ~pi590 & ~n46621;
  assign n46623 = pi450 & n46107;
  assign n46624 = ~pi588 & ~n46623;
  assign n46625 = ~n46622 & n46624;
  assign n46626 = pi438 & n46111;
  assign n46627 = pi588 & ~n46626;
  assign n46628 = n46096 & ~n46627;
  assign n46629 = ~n46625 & n46628;
  assign n46630 = ~n46617 & ~n46629;
  assign n46631 = n8830 & ~n46630;
  assign n46632 = ~pi665 & pi1136;
  assign n46633 = ~pi791 & ~pi1136;
  assign n46634 = pi1135 & ~n46633;
  assign n46635 = ~n46632 & n46634;
  assign n46636 = ~pi621 & pi1136;
  assign n46637 = ~pi810 & ~pi1136;
  assign n46638 = ~pi1135 & ~n46637;
  assign n46639 = ~n46636 & n46638;
  assign n46640 = ~n46635 & ~n46639;
  assign n46641 = n46119 & ~n46640;
  assign n46642 = ~pi739 & n46131;
  assign n46643 = ~pi874 & ~pi1136;
  assign n46644 = ~pi690 & pi1135;
  assign n46645 = ~n46643 & ~n46644;
  assign n46646 = n46135 & n46645;
  assign n46647 = ~n46642 & n46646;
  assign n46648 = ~n46641 & ~n46647;
  assign n46649 = ~n8830 & ~n46648;
  assign po836 = n46631 | n46649;
  assign n46651 = ~pi1100 & po954;
  assign n46652 = ~pi680 & ~po954;
  assign n46653 = ~pi962 & ~n46652;
  assign po837 = ~n46651 & n46653;
  assign n46655 = ~pi1103 & po954;
  assign n46656 = ~pi681 & ~po954;
  assign n46657 = ~pi962 & ~n46656;
  assign po838 = ~n46655 & n46657;
  assign n46659 = pi199 & ~pi1039;
  assign n46660 = ~pi199 & ~pi251;
  assign n46661 = ~n46096 & ~n46660;
  assign n46662 = ~n46659 & n46661;
  assign n46663 = pi367 & n46100;
  assign n46664 = pi392 & pi591;
  assign n46665 = ~pi592 & n46664;
  assign n46666 = ~n46663 & ~n46665;
  assign n46667 = ~pi590 & ~n46666;
  assign n46668 = pi345 & n46107;
  assign n46669 = ~pi588 & ~n46668;
  assign n46670 = ~n46667 & n46669;
  assign n46671 = pi417 & n46111;
  assign n46672 = pi588 & ~n46671;
  assign n46673 = n46096 & ~n46672;
  assign n46674 = ~n46670 & n46673;
  assign n46675 = ~n46662 & ~n46674;
  assign n46676 = n8830 & ~n46675;
  assign n46677 = pi757 & n46131;
  assign n46678 = pi686 & pi1135;
  assign n46679 = ~pi848 & ~pi1136;
  assign n46680 = ~n46678 & ~n46679;
  assign n46681 = n46135 & n46680;
  assign n46682 = ~n46677 & n46681;
  assign n46683 = ~pi610 & ~pi1135;
  assign n46684 = pi631 & pi1135;
  assign n46685 = ~pi1134 & ~n46684;
  assign n46686 = ~n46683 & n46685;
  assign n46687 = n46327 & n46686;
  assign n46688 = ~n46682 & ~n46687;
  assign n46689 = ~n8830 & ~n46688;
  assign po839 = n46676 | n46689;
  assign po980 = pi953 & n45933;
  assign n46692 = pi684 & ~po980;
  assign n46693 = ~pi1130 & po980;
  assign n46694 = ~pi962 & ~n46693;
  assign po841 = ~n46692 & n46694;
  assign n46696 = pi590 & ~pi592;
  assign n46697 = pi357 & n46696;
  assign n46698 = pi382 & n46146;
  assign n46699 = ~n46697 & ~n46698;
  assign n46700 = ~pi591 & ~n46699;
  assign n46701 = pi406 & ~pi592;
  assign n46702 = n46144 & n46701;
  assign n46703 = ~n46700 & ~n46702;
  assign n46704 = ~pi588 & ~n46703;
  assign n46705 = pi588 & ~pi590;
  assign n46706 = pi430 & n46106;
  assign n46707 = n46705 & n46706;
  assign n46708 = ~n46704 & ~n46707;
  assign n46709 = n46096 & ~n46708;
  assign n46710 = pi199 & ~pi1076;
  assign n46711 = ~n46096 & ~n46710;
  assign n46712 = ~n42268 & n46711;
  assign n46713 = ~n46709 & ~n46712;
  assign n46714 = n8830 & ~n46713;
  assign n46715 = pi860 & n46178;
  assign n46716 = pi728 & pi1135;
  assign n46717 = pi744 & ~pi1135;
  assign n46718 = pi1136 & ~n46717;
  assign n46719 = ~n46716 & n46718;
  assign n46720 = ~n46715 & ~n46719;
  assign n46721 = n46134 & ~n46720;
  assign n46722 = pi1136 & ~n46118;
  assign n46723 = ~pi1134 & ~n46722;
  assign n46724 = pi657 & pi1135;
  assign n46725 = ~pi652 & ~pi1135;
  assign n46726 = pi1136 & ~n46725;
  assign n46727 = ~n46724 & n46726;
  assign n46728 = pi813 & n46118;
  assign n46729 = n46178 & n46728;
  assign n46730 = ~n46727 & ~n46729;
  assign n46731 = n46723 & ~n46730;
  assign n46732 = ~n46721 & ~n46731;
  assign n46733 = ~n8830 & ~n46732;
  assign po842 = n46714 | n46733;
  assign n46735 = pi686 & ~po980;
  assign n46736 = ~pi1113 & po980;
  assign n46737 = ~pi962 & ~n46736;
  assign po843 = ~n46735 & n46737;
  assign n46739 = ~pi1127 & po980;
  assign n46740 = ~pi687 & ~po980;
  assign n46741 = ~pi962 & ~n46740;
  assign po844 = ~n46739 & n46741;
  assign n46743 = pi688 & ~po980;
  assign n46744 = ~pi1115 & po980;
  assign n46745 = ~pi962 & ~n46744;
  assign po845 = ~n46743 & n46745;
  assign n46747 = pi351 & n46696;
  assign n46748 = pi376 & n46146;
  assign n46749 = ~n46747 & ~n46748;
  assign n46750 = ~pi591 & ~n46749;
  assign n46751 = pi401 & ~pi592;
  assign n46752 = n46144 & n46751;
  assign n46753 = ~n46750 & ~n46752;
  assign n46754 = ~pi588 & ~n46753;
  assign n46755 = pi426 & n46106;
  assign n46756 = n46705 & n46755;
  assign n46757 = ~n46754 & ~n46756;
  assign n46758 = n46096 & ~n46757;
  assign n46759 = ~pi199 & n42237;
  assign n46760 = pi199 & ~pi1079;
  assign n46761 = ~n46096 & ~n46760;
  assign n46762 = ~n46759 & n46761;
  assign n46763 = ~n46758 & ~n46762;
  assign n46764 = n8830 & ~n46763;
  assign n46765 = pi798 & n46178;
  assign n46766 = pi655 & pi1135;
  assign n46767 = ~pi658 & ~pi1135;
  assign n46768 = pi1136 & ~n46767;
  assign n46769 = ~n46766 & n46768;
  assign n46770 = ~n46765 & ~n46769;
  assign n46771 = n46119 & ~n46770;
  assign n46772 = pi752 & n46131;
  assign n46773 = ~pi703 & pi1135;
  assign n46774 = ~pi843 & ~pi1136;
  assign n46775 = ~n46773 & ~n46774;
  assign n46776 = n46135 & n46775;
  assign n46777 = ~n46772 & n46776;
  assign n46778 = ~n46771 & ~n46777;
  assign n46779 = ~n8830 & ~n46778;
  assign po846 = n46764 | n46779;
  assign n46781 = ~pi1108 & po980;
  assign n46782 = ~pi690 & ~po980;
  assign n46783 = ~pi962 & ~n46782;
  assign po847 = ~n46781 & n46783;
  assign n46785 = ~pi1107 & po980;
  assign n46786 = ~pi691 & ~po980;
  assign n46787 = ~pi962 & ~n46786;
  assign po848 = ~n46785 & n46787;
  assign n46789 = pi352 & n46696;
  assign n46790 = pi317 & n46146;
  assign n46791 = ~n46789 & ~n46790;
  assign n46792 = ~pi591 & ~n46791;
  assign n46793 = pi402 & ~pi592;
  assign n46794 = n46144 & n46793;
  assign n46795 = ~n46792 & ~n46794;
  assign n46796 = ~pi588 & ~n46795;
  assign n46797 = pi427 & n46106;
  assign n46798 = n46705 & n46797;
  assign n46799 = ~n46796 & ~n46798;
  assign n46800 = n46096 & ~n46799;
  assign n46801 = ~pi199 & n42249;
  assign n46802 = pi199 & ~pi1078;
  assign n46803 = ~n46096 & ~n46802;
  assign n46804 = ~n46801 & n46803;
  assign n46805 = ~n46800 & ~n46804;
  assign n46806 = n8830 & ~n46805;
  assign n46807 = pi649 & pi1135;
  assign n46808 = ~pi656 & ~pi1135;
  assign n46809 = pi1136 & ~n46808;
  assign n46810 = ~n46807 & n46809;
  assign n46811 = pi801 & n46178;
  assign n46812 = ~pi1134 & ~n46811;
  assign n46813 = ~n46810 & n46812;
  assign n46814 = pi770 & ~pi1135;
  assign n46815 = ~pi726 & pi1135;
  assign n46816 = pi1136 & ~n46815;
  assign n46817 = ~n46814 & n46816;
  assign n46818 = pi844 & n46178;
  assign n46819 = pi1134 & ~n46818;
  assign n46820 = ~n46817 & n46819;
  assign n46821 = n46182 & ~n46820;
  assign n46822 = ~n46813 & n46821;
  assign po849 = n46806 | n46822;
  assign n46824 = pi693 & ~po954;
  assign n46825 = ~pi1129 & po954;
  assign n46826 = ~pi962 & ~n46825;
  assign po850 = ~n46824 & n46826;
  assign n46828 = pi694 & ~po980;
  assign n46829 = ~pi1128 & po980;
  assign n46830 = ~pi962 & ~n46829;
  assign po851 = ~n46828 & n46830;
  assign n46832 = pi695 & ~po954;
  assign n46833 = ~pi1111 & po954;
  assign n46834 = ~pi962 & ~n46833;
  assign po852 = ~n46832 & n46834;
  assign n46836 = ~pi1100 & po980;
  assign n46837 = ~pi696 & ~po980;
  assign n46838 = ~pi962 & ~n46837;
  assign po853 = ~n46836 & n46838;
  assign n46840 = pi697 & ~po980;
  assign n46841 = ~pi1129 & po980;
  assign n46842 = ~pi962 & ~n46841;
  assign po854 = ~n46840 & n46842;
  assign n46844 = pi698 & ~po980;
  assign n46845 = ~pi1116 & po980;
  assign n46846 = ~pi962 & ~n46845;
  assign po855 = ~n46844 & n46846;
  assign n46848 = ~pi1103 & po980;
  assign n46849 = ~pi699 & ~po980;
  assign n46850 = ~pi962 & ~n46849;
  assign po856 = ~n46848 & n46850;
  assign n46852 = ~pi1110 & po980;
  assign n46853 = ~pi700 & ~po980;
  assign n46854 = ~pi962 & ~n46853;
  assign po857 = ~n46852 & n46854;
  assign n46856 = pi701 & ~po980;
  assign n46857 = ~pi1123 & po980;
  assign n46858 = ~pi962 & ~n46857;
  assign po858 = ~n46856 & n46858;
  assign n46860 = pi702 & ~po980;
  assign n46861 = ~pi1117 & po980;
  assign n46862 = ~pi962 & ~n46861;
  assign po859 = ~n46860 & n46862;
  assign n46864 = ~pi1124 & po980;
  assign n46865 = ~pi703 & ~po980;
  assign n46866 = ~pi962 & ~n46865;
  assign po860 = ~n46864 & n46866;
  assign n46868 = pi704 & ~po980;
  assign n46869 = ~pi1112 & po980;
  assign n46870 = ~pi962 & ~n46869;
  assign po861 = ~n46868 & n46870;
  assign n46872 = ~pi1125 & po980;
  assign n46873 = ~pi705 & ~po980;
  assign n46874 = ~pi962 & ~n46873;
  assign po862 = ~n46872 & n46874;
  assign n46876 = ~pi1105 & po980;
  assign n46877 = ~pi706 & ~po980;
  assign n46878 = ~pi962 & ~n46877;
  assign po863 = ~n46876 & n46878;
  assign n46880 = pi370 & n46100;
  assign n46881 = pi395 & pi591;
  assign n46882 = ~pi592 & n46881;
  assign n46883 = ~n46880 & ~n46882;
  assign n46884 = ~pi590 & ~n46883;
  assign n46885 = pi347 & n46107;
  assign n46886 = ~n46884 & ~n46885;
  assign n46887 = ~pi588 & n46096;
  assign n46888 = ~n46886 & n46887;
  assign n46889 = ~pi200 & ~pi304;
  assign n46890 = pi200 & ~pi1048;
  assign n46891 = ~n46889 & ~n46890;
  assign n46892 = ~pi199 & ~n46891;
  assign n46893 = pi199 & ~pi1055;
  assign n46894 = ~n46096 & ~n46893;
  assign n46895 = ~n46892 & n46894;
  assign n46896 = n46096 & n46111;
  assign n46897 = pi420 & pi588;
  assign n46898 = n46896 & n46897;
  assign n46899 = ~n46895 & ~n46898;
  assign n46900 = ~n46888 & n46899;
  assign n46901 = n8830 & ~n46900;
  assign n46902 = ~pi618 & ~pi1135;
  assign n46903 = ~pi627 & pi1135;
  assign n46904 = ~pi1134 & ~n46903;
  assign n46905 = ~n46902 & n46904;
  assign n46906 = n46327 & n46905;
  assign n46907 = pi753 & n46131;
  assign n46908 = pi702 & pi1135;
  assign n46909 = ~pi847 & ~pi1136;
  assign n46910 = ~n46908 & ~n46909;
  assign n46911 = n46135 & n46910;
  assign n46912 = ~n46907 & n46911;
  assign n46913 = ~n46906 & ~n46912;
  assign n46914 = ~n8830 & ~n46913;
  assign po864 = n46901 | n46914;
  assign n46916 = n46096 & n46100;
  assign n46917 = pi442 & n46916;
  assign n46918 = ~pi592 & n46096;
  assign n46919 = pi328 & pi591;
  assign n46920 = n46918 & n46919;
  assign n46921 = ~n46917 & ~n46920;
  assign n46922 = ~pi590 & ~n46921;
  assign n46923 = pi321 & n46096;
  assign n46924 = n46107 & n46923;
  assign n46925 = ~n46922 & ~n46924;
  assign n46926 = ~pi588 & ~n46925;
  assign n46927 = ~pi200 & ~pi305;
  assign n46928 = pi200 & ~pi1084;
  assign n46929 = ~n46927 & ~n46928;
  assign n46930 = ~pi199 & ~n46929;
  assign n46931 = pi199 & ~pi1058;
  assign n46932 = ~n46096 & ~n46931;
  assign n46933 = ~n46930 & n46932;
  assign n46934 = n46096 & n46106;
  assign n46935 = pi459 & n46705;
  assign n46936 = n46934 & n46935;
  assign n46937 = n8830 & ~n46936;
  assign n46938 = ~n46933 & n46937;
  assign n46939 = ~n46926 & n46938;
  assign n46940 = pi754 & n46131;
  assign n46941 = n46118 & ~n46133;
  assign n46942 = ~pi857 & ~pi1136;
  assign n46943 = pi709 & pi1135;
  assign n46944 = pi1134 & ~n46943;
  assign n46945 = ~n46942 & n46944;
  assign n46946 = n46941 & n46945;
  assign n46947 = ~n46940 & n46946;
  assign n46948 = ~pi660 & pi1135;
  assign n46949 = ~pi609 & ~pi1135;
  assign n46950 = ~pi1134 & ~n46949;
  assign n46951 = ~n46948 & n46950;
  assign n46952 = n46327 & n46951;
  assign n46953 = ~n8830 & ~n46952;
  assign n46954 = ~n46947 & n46953;
  assign po865 = ~n46939 & ~n46954;
  assign n46956 = pi709 & ~po980;
  assign n46957 = ~pi1118 & po980;
  assign n46958 = ~pi962 & ~n46957;
  assign po866 = ~n46956 & n46958;
  assign n46960 = ~pi1106 & po954;
  assign n46961 = ~pi710 & ~po954;
  assign n46962 = ~pi962 & ~n46961;
  assign po867 = ~n46960 & n46962;
  assign n46964 = pi373 & n46100;
  assign n46965 = pi398 & pi591;
  assign n46966 = ~pi592 & n46965;
  assign n46967 = ~n46964 & ~n46966;
  assign n46968 = ~pi590 & ~n46967;
  assign n46969 = pi348 & n46107;
  assign n46970 = ~n46968 & ~n46969;
  assign n46971 = n46887 & ~n46970;
  assign n46972 = ~pi200 & ~pi306;
  assign n46973 = pi200 & ~pi1059;
  assign n46974 = ~n46972 & ~n46973;
  assign n46975 = ~pi199 & ~n46974;
  assign n46976 = pi199 & ~pi1087;
  assign n46977 = ~n46096 & ~n46976;
  assign n46978 = ~n46975 & n46977;
  assign n46979 = pi423 & pi588;
  assign n46980 = n46896 & n46979;
  assign n46981 = ~n46978 & ~n46980;
  assign n46982 = ~n46971 & n46981;
  assign n46983 = n8830 & ~n46982;
  assign n46984 = ~pi630 & ~pi1135;
  assign n46985 = ~pi647 & pi1135;
  assign n46986 = ~pi1134 & ~n46985;
  assign n46987 = ~n46984 & n46986;
  assign n46988 = n46327 & n46987;
  assign n46989 = pi755 & n46131;
  assign n46990 = pi725 & pi1135;
  assign n46991 = ~pi858 & ~pi1136;
  assign n46992 = ~n46990 & ~n46991;
  assign n46993 = n46135 & n46992;
  assign n46994 = ~n46989 & n46993;
  assign n46995 = ~n46988 & ~n46994;
  assign n46996 = ~n8830 & ~n46995;
  assign po868 = n46983 | n46996;
  assign n46998 = pi751 & n46131;
  assign n46999 = ~pi842 & ~pi1136;
  assign n47000 = pi701 & pi1135;
  assign n47001 = pi1134 & ~n47000;
  assign n47002 = ~n46999 & n47001;
  assign n47003 = n46941 & n47002;
  assign n47004 = ~n46998 & n47003;
  assign n47005 = ~pi644 & ~pi1135;
  assign n47006 = ~pi715 & pi1135;
  assign n47007 = ~pi1134 & ~n47006;
  assign n47008 = ~n47005 & n47007;
  assign n47009 = n46327 & n47008;
  assign n47010 = ~n47004 & ~n47009;
  assign n47011 = ~n8830 & ~n47010;
  assign n47012 = pi374 & n46100;
  assign n47013 = pi400 & pi591;
  assign n47014 = ~pi592 & n47013;
  assign n47015 = ~n47012 & ~n47014;
  assign n47016 = ~pi590 & ~n47015;
  assign n47017 = pi350 & n46107;
  assign n47018 = ~n47016 & ~n47017;
  assign n47019 = ~pi588 & ~n47018;
  assign n47020 = pi425 & n46106;
  assign n47021 = n46705 & n47020;
  assign n47022 = n46096 & ~n47021;
  assign n47023 = ~n47019 & n47022;
  assign n47024 = pi1044 & n11381;
  assign n47025 = pi298 & n10758;
  assign n47026 = pi199 & pi1035;
  assign n47027 = ~n46096 & ~n47026;
  assign n47028 = ~n47025 & n47027;
  assign n47029 = ~n47024 & n47028;
  assign n47030 = n8830 & ~n47029;
  assign n47031 = ~n47023 & n47030;
  assign po869 = n47011 | n47031;
  assign n47033 = pi371 & n46100;
  assign n47034 = pi396 & pi591;
  assign n47035 = ~pi592 & n47034;
  assign n47036 = ~n47033 & ~n47035;
  assign n47037 = ~pi590 & ~n47036;
  assign n47038 = pi322 & n46107;
  assign n47039 = ~n47037 & ~n47038;
  assign n47040 = n46887 & ~n47039;
  assign n47041 = ~pi200 & ~pi309;
  assign n47042 = pi200 & ~pi1072;
  assign n47043 = ~n47041 & ~n47042;
  assign n47044 = ~pi199 & ~n47043;
  assign n47045 = pi199 & ~pi1051;
  assign n47046 = ~n46096 & ~n47045;
  assign n47047 = ~n47044 & n47046;
  assign n47048 = pi421 & pi588;
  assign n47049 = n46896 & n47048;
  assign n47050 = ~n47047 & ~n47049;
  assign n47051 = ~n47040 & n47050;
  assign n47052 = n8830 & ~n47051;
  assign n47053 = ~pi629 & ~pi1135;
  assign n47054 = ~pi628 & pi1135;
  assign n47055 = ~pi1134 & ~n47054;
  assign n47056 = ~n47053 & n47055;
  assign n47057 = n46327 & n47056;
  assign n47058 = pi756 & n46131;
  assign n47059 = pi734 & pi1135;
  assign n47060 = ~pi854 & ~pi1136;
  assign n47061 = ~n47059 & ~n47060;
  assign n47062 = n46135 & n47061;
  assign n47063 = ~n47058 & n47062;
  assign n47064 = ~n47057 & ~n47063;
  assign n47065 = ~n8830 & ~n47064;
  assign po870 = n47052 | n47065;
  assign n47067 = pi461 & n46696;
  assign n47068 = pi439 & n46146;
  assign n47069 = ~n47067 & ~n47068;
  assign n47070 = ~pi591 & ~n47069;
  assign n47071 = pi326 & ~pi592;
  assign n47072 = n46144 & n47071;
  assign n47073 = ~n47070 & ~n47072;
  assign n47074 = ~pi588 & ~n47073;
  assign n47075 = pi449 & n46106;
  assign n47076 = n46705 & n47075;
  assign n47077 = ~n47074 & ~n47076;
  assign n47078 = n46096 & ~n47077;
  assign n47079 = pi199 & ~pi1057;
  assign n47080 = ~n46096 & ~n47079;
  assign n47081 = ~n41732 & n47080;
  assign n47082 = ~n47078 & ~n47081;
  assign n47083 = n8830 & ~n47082;
  assign n47084 = pi867 & n46178;
  assign n47085 = pi697 & pi1135;
  assign n47086 = pi762 & ~pi1135;
  assign n47087 = pi1136 & ~n47086;
  assign n47088 = ~n47085 & n47087;
  assign n47089 = ~n47084 & ~n47088;
  assign n47090 = n46134 & ~n47089;
  assign n47091 = pi693 & pi1135;
  assign n47092 = ~pi653 & ~pi1135;
  assign n47093 = pi1136 & ~n47092;
  assign n47094 = ~n47091 & n47093;
  assign n47095 = pi816 & n46118;
  assign n47096 = n46178 & n47095;
  assign n47097 = ~n47094 & ~n47096;
  assign n47098 = n46723 & ~n47097;
  assign n47099 = ~n47090 & ~n47098;
  assign n47100 = ~n8830 & ~n47099;
  assign po871 = n47083 | n47100;
  assign n47102 = ~pi1123 & po954;
  assign n47103 = ~pi715 & ~po954;
  assign n47104 = ~pi962 & ~n47103;
  assign po872 = ~n47102 & n47104;
  assign n47106 = pi440 & n46916;
  assign n47107 = pi329 & pi591;
  assign n47108 = n46918 & n47107;
  assign n47109 = ~n47106 & ~n47108;
  assign n47110 = ~pi590 & ~n47109;
  assign n47111 = pi349 & n46096;
  assign n47112 = n46107 & n47111;
  assign n47113 = ~n47110 & ~n47112;
  assign n47114 = ~pi588 & ~n47113;
  assign n47115 = ~pi200 & ~pi307;
  assign n47116 = pi200 & ~pi1053;
  assign n47117 = ~n47115 & ~n47116;
  assign n47118 = ~pi199 & ~n47117;
  assign n47119 = pi199 & ~pi1043;
  assign n47120 = ~n46096 & ~n47119;
  assign n47121 = ~n47118 & n47120;
  assign n47122 = pi454 & n46705;
  assign n47123 = n46934 & n47122;
  assign n47124 = n8830 & ~n47123;
  assign n47125 = ~n47121 & n47124;
  assign n47126 = ~n47114 & n47125;
  assign n47127 = pi761 & n46131;
  assign n47128 = ~pi845 & ~pi1136;
  assign n47129 = pi738 & pi1135;
  assign n47130 = pi1134 & ~n47129;
  assign n47131 = ~n47128 & n47130;
  assign n47132 = n46941 & n47131;
  assign n47133 = ~n47127 & n47132;
  assign n47134 = ~pi641 & pi1135;
  assign n47135 = ~pi626 & ~pi1135;
  assign n47136 = ~pi1134 & ~n47135;
  assign n47137 = ~n47134 & n47136;
  assign n47138 = n46327 & n47137;
  assign n47139 = ~n8830 & ~n47138;
  assign n47140 = ~n47133 & n47139;
  assign po873 = ~n47126 & ~n47140;
  assign n47142 = pi318 & pi591;
  assign n47143 = ~pi592 & n47142;
  assign n47144 = ~pi591 & n7749;
  assign n47145 = ~n47143 & ~n47144;
  assign n47146 = ~pi590 & ~n47145;
  assign n47147 = pi462 & n46107;
  assign n47148 = ~n47146 & ~n47147;
  assign n47149 = n46887 & ~n47148;
  assign n47150 = ~pi199 & n42243;
  assign n47151 = pi199 & ~pi1074;
  assign n47152 = ~n46096 & ~n47151;
  assign n47153 = ~n47150 & n47152;
  assign n47154 = pi448 & pi588;
  assign n47155 = n46896 & n47154;
  assign n47156 = ~n47153 & ~n47155;
  assign n47157 = ~n47149 & n47156;
  assign n47158 = n8830 & ~n47157;
  assign n47159 = pi768 & n46131;
  assign n47160 = ~pi839 & ~pi1136;
  assign n47161 = ~pi705 & pi1135;
  assign n47162 = pi1134 & ~n47161;
  assign n47163 = ~n47160 & n47162;
  assign n47164 = n46941 & n47163;
  assign n47165 = ~n47159 & n47164;
  assign n47166 = pi800 & n46178;
  assign n47167 = pi669 & pi1135;
  assign n47168 = ~pi645 & ~pi1135;
  assign n47169 = pi1136 & ~n47168;
  assign n47170 = ~n47167 & n47169;
  assign n47171 = ~n47166 & ~n47170;
  assign n47172 = n46119 & ~n47171;
  assign n47173 = ~n47165 & ~n47172;
  assign n47174 = ~n8830 & ~n47173;
  assign po874 = n47158 | n47174;
  assign n47176 = pi369 & n46916;
  assign n47177 = pi394 & pi591;
  assign n47178 = n46918 & n47177;
  assign n47179 = ~n47176 & ~n47178;
  assign n47180 = ~pi590 & ~n47179;
  assign n47181 = pi315 & n46096;
  assign n47182 = n46107 & n47181;
  assign n47183 = ~n47180 & ~n47182;
  assign n47184 = ~pi588 & ~n47183;
  assign n47185 = ~pi200 & ~pi303;
  assign n47186 = pi200 & ~pi1049;
  assign n47187 = ~n47185 & ~n47186;
  assign n47188 = ~pi199 & ~n47187;
  assign n47189 = pi199 & ~pi1080;
  assign n47190 = ~n46096 & ~n47189;
  assign n47191 = ~n47188 & n47190;
  assign n47192 = pi419 & n46705;
  assign n47193 = n46934 & n47192;
  assign n47194 = n8830 & ~n47193;
  assign n47195 = ~n47191 & n47194;
  assign n47196 = ~n47184 & n47195;
  assign n47197 = pi767 & n46131;
  assign n47198 = ~pi853 & ~pi1136;
  assign n47199 = pi698 & pi1135;
  assign n47200 = pi1134 & ~n47199;
  assign n47201 = ~n47198 & n47200;
  assign n47202 = n46941 & n47201;
  assign n47203 = ~n47197 & n47202;
  assign n47204 = ~pi625 & pi1135;
  assign n47205 = ~pi608 & ~pi1135;
  assign n47206 = ~pi1134 & ~n47205;
  assign n47207 = ~n47204 & n47206;
  assign n47208 = n46327 & n47207;
  assign n47209 = ~n8830 & ~n47208;
  assign n47210 = ~n47203 & n47209;
  assign po875 = ~n47196 & ~n47210;
  assign n47212 = pi378 & n46100;
  assign n47213 = pi325 & pi591;
  assign n47214 = ~pi592 & n47213;
  assign n47215 = ~n47212 & ~n47214;
  assign n47216 = ~pi590 & ~n47215;
  assign n47217 = pi353 & n46107;
  assign n47218 = ~n47216 & ~n47217;
  assign n47219 = n46887 & ~n47218;
  assign n47220 = ~pi199 & n42255;
  assign n47221 = pi199 & ~pi1063;
  assign n47222 = ~n46096 & ~n47221;
  assign n47223 = ~n47220 & n47222;
  assign n47224 = pi451 & pi588;
  assign n47225 = n46896 & n47224;
  assign n47226 = ~n47223 & ~n47225;
  assign n47227 = ~n47219 & n47226;
  assign n47228 = n8830 & ~n47227;
  assign n47229 = pi774 & n46131;
  assign n47230 = ~pi868 & ~pi1136;
  assign n47231 = ~pi687 & pi1135;
  assign n47232 = pi1134 & ~n47231;
  assign n47233 = ~n47230 & n47232;
  assign n47234 = n46941 & n47233;
  assign n47235 = ~n47229 & n47234;
  assign n47236 = pi807 & n46178;
  assign n47237 = pi650 & pi1135;
  assign n47238 = ~pi636 & ~pi1135;
  assign n47239 = pi1136 & ~n47238;
  assign n47240 = ~n47237 & n47239;
  assign n47241 = ~n47236 & ~n47240;
  assign n47242 = n46119 & ~n47241;
  assign n47243 = ~n47235 & ~n47242;
  assign n47244 = ~n8830 & ~n47243;
  assign po876 = n47228 | n47244;
  assign n47246 = pi356 & n46696;
  assign n47247 = pi381 & n46146;
  assign n47248 = ~n47246 & ~n47247;
  assign n47249 = ~pi591 & ~n47248;
  assign n47250 = pi405 & ~pi592;
  assign n47251 = n46144 & n47250;
  assign n47252 = ~n47249 & ~n47251;
  assign n47253 = ~pi588 & ~n47252;
  assign n47254 = pi445 & n46106;
  assign n47255 = n46705 & n47254;
  assign n47256 = ~n47253 & ~n47255;
  assign n47257 = n46096 & ~n47256;
  assign n47258 = pi199 & ~pi1081;
  assign n47259 = ~n46096 & ~n47258;
  assign n47260 = ~n42275 & n47259;
  assign n47261 = ~n47257 & ~n47260;
  assign n47262 = n8830 & ~n47261;
  assign n47263 = pi880 & n46178;
  assign n47264 = pi684 & pi1135;
  assign n47265 = pi750 & ~pi1135;
  assign n47266 = pi1136 & ~n47265;
  assign n47267 = ~n47264 & n47266;
  assign n47268 = ~n47263 & ~n47267;
  assign n47269 = n46134 & ~n47268;
  assign n47270 = pi654 & pi1135;
  assign n47271 = ~pi651 & ~pi1135;
  assign n47272 = pi1136 & ~n47271;
  assign n47273 = ~n47270 & n47272;
  assign n47274 = pi794 & n46118;
  assign n47275 = n46178 & n47274;
  assign n47276 = ~n47273 & ~n47275;
  assign n47277 = n46723 & ~n47276;
  assign n47278 = ~n47269 & ~n47277;
  assign n47279 = ~n8830 & ~n47278;
  assign po877 = n47262 | n47279;
  assign n47281 = pi747 & pi773;
  assign n47282 = pi769 & n47281;
  assign n47283 = ~pi721 & ~n47282;
  assign n47284 = pi721 & n47282;
  assign n47285 = pi775 & ~n47284;
  assign n47286 = ~n47283 & n47285;
  assign n47287 = pi721 & pi813;
  assign n47288 = ~pi773 & ~pi801;
  assign n47289 = pi773 & pi801;
  assign n47290 = ~n47288 & ~n47289;
  assign n47291 = ~pi771 & ~pi800;
  assign n47292 = pi771 & pi800;
  assign n47293 = ~n47291 & ~n47292;
  assign n47294 = ~pi769 & ~pi794;
  assign n47295 = pi769 & pi794;
  assign n47296 = ~n47294 & ~n47295;
  assign n47297 = ~pi765 & ~pi798;
  assign n47298 = pi765 & pi798;
  assign n47299 = ~n47297 & ~n47298;
  assign n47300 = pi807 & ~n47299;
  assign n47301 = pi747 & n47300;
  assign n47302 = ~pi747 & ~pi807;
  assign n47303 = ~n47299 & n47302;
  assign n47304 = ~n47301 & ~n47303;
  assign n47305 = ~n47296 & ~n47304;
  assign n47306 = ~n47293 & n47305;
  assign n47307 = ~n47290 & n47306;
  assign n47308 = n47287 & n47307;
  assign n47309 = ~n47293 & n47300;
  assign n47310 = ~pi721 & ~pi813;
  assign n47311 = pi794 & pi801;
  assign n47312 = n47310 & n47311;
  assign n47313 = n47309 & n47312;
  assign n47314 = ~n47308 & ~n47313;
  assign n47315 = pi816 & ~n47314;
  assign n47316 = n47286 & ~n47315;
  assign n47317 = pi795 & ~n47316;
  assign n47318 = ~pi945 & pi988;
  assign n47319 = pi731 & n47318;
  assign n47320 = pi721 & ~pi775;
  assign n47321 = ~n47286 & ~n47320;
  assign n47322 = n47319 & ~n47321;
  assign n47323 = ~n47317 & n47322;
  assign n47324 = ~pi775 & ~pi816;
  assign n47325 = pi775 & pi816;
  assign n47326 = ~n47324 & ~n47325;
  assign n47327 = n47308 & ~n47326;
  assign n47328 = n47320 & ~n47327;
  assign n47329 = pi721 & ~n47319;
  assign n47330 = ~pi731 & ~pi795;
  assign n47331 = pi731 & pi795;
  assign n47332 = ~n47330 & ~n47331;
  assign n47333 = ~n47287 & ~n47310;
  assign n47334 = ~n47326 & ~n47333;
  assign n47335 = ~n47332 & n47334;
  assign po978 = n47307 & n47335;
  assign n47337 = n47329 & ~po978;
  assign n47338 = ~n47328 & ~n47337;
  assign po878 = n47323 | ~n47338;
  assign n47340 = pi379 & n46100;
  assign n47341 = pi403 & pi591;
  assign n47342 = ~pi592 & n47341;
  assign n47343 = ~n47340 & ~n47342;
  assign n47344 = ~pi590 & ~n47343;
  assign n47345 = pi354 & n46107;
  assign n47346 = ~n47344 & ~n47345;
  assign n47347 = n46887 & ~n47346;
  assign n47348 = ~pi199 & n42261;
  assign n47349 = pi199 & ~pi1045;
  assign n47350 = ~n46096 & ~n47349;
  assign n47351 = ~n47348 & n47350;
  assign n47352 = pi428 & pi588;
  assign n47353 = n46896 & n47352;
  assign n47354 = ~n47351 & ~n47353;
  assign n47355 = ~n47347 & n47354;
  assign n47356 = n8830 & ~n47355;
  assign n47357 = ~pi851 & pi1134;
  assign n47358 = ~pi795 & ~pi1134;
  assign n47359 = ~pi1136 & ~n47358;
  assign n47360 = ~n47357 & n47359;
  assign n47361 = pi776 & pi1134;
  assign n47362 = ~pi640 & ~pi1134;
  assign n47363 = pi1136 & ~n47362;
  assign n47364 = ~n47361 & n47363;
  assign n47365 = ~n47360 & ~n47364;
  assign n47366 = ~pi1135 & ~n47365;
  assign n47367 = pi732 & ~pi1134;
  assign n47368 = pi694 & pi1134;
  assign n47369 = pi1135 & pi1136;
  assign n47370 = ~n47368 & n47369;
  assign n47371 = ~n47367 & n47370;
  assign n47372 = ~n47366 & ~n47371;
  assign n47373 = n46182 & ~n47372;
  assign po879 = n47356 | n47373;
  assign n47375 = pi723 & ~po980;
  assign n47376 = ~pi1111 & po980;
  assign n47377 = ~pi962 & ~n47376;
  assign po880 = ~n47375 & n47377;
  assign n47379 = pi724 & ~po980;
  assign n47380 = ~pi1114 & po980;
  assign n47381 = ~pi962 & ~n47380;
  assign po881 = ~n47379 & n47381;
  assign n47383 = pi725 & ~po980;
  assign n47384 = ~pi1120 & po980;
  assign n47385 = ~pi962 & ~n47384;
  assign po882 = ~n47383 & n47385;
  assign n47387 = ~pi1126 & po980;
  assign n47388 = ~pi726 & ~po980;
  assign n47389 = ~pi962 & ~n47388;
  assign po883 = ~n47387 & n47389;
  assign n47391 = ~pi1102 & po980;
  assign n47392 = ~pi727 & ~po980;
  assign n47393 = ~pi962 & ~n47392;
  assign po884 = ~n47391 & n47393;
  assign n47395 = pi728 & ~po980;
  assign n47396 = ~pi1131 & po980;
  assign n47397 = ~pi962 & ~n47396;
  assign po885 = ~n47395 & n47397;
  assign n47399 = ~pi1104 & po980;
  assign n47400 = ~pi729 & ~po980;
  assign n47401 = ~pi962 & ~n47400;
  assign po886 = ~n47399 & n47401;
  assign n47403 = ~pi1106 & po980;
  assign n47404 = ~pi730 & ~po980;
  assign n47405 = ~pi962 & ~n47404;
  assign po887 = ~n47403 & n47405;
  assign n47407 = n47307 & ~n47333;
  assign n47408 = pi795 & ~n47326;
  assign n47409 = n47407 & n47408;
  assign n47410 = ~n47281 & ~n47409;
  assign n47411 = n47319 & ~n47410;
  assign n47412 = pi731 & ~n47409;
  assign n47413 = ~pi795 & pi801;
  assign n47414 = ~n47296 & n47413;
  assign n47415 = n47334 & n47414;
  assign n47416 = n47309 & n47415;
  assign n47417 = n47281 & ~n47416;
  assign n47418 = ~pi731 & ~n47417;
  assign n47419 = n47318 & ~n47418;
  assign n47420 = ~n47412 & ~n47419;
  assign po888 = ~n47411 & ~n47420;
  assign n47422 = pi732 & ~po954;
  assign n47423 = ~pi1128 & po954;
  assign n47424 = ~pi962 & ~n47423;
  assign po889 = ~n47422 & n47424;
  assign n47426 = pi375 & n46916;
  assign n47427 = pi399 & pi591;
  assign n47428 = n46918 & n47427;
  assign n47429 = ~n47426 & ~n47428;
  assign n47430 = ~pi590 & ~n47429;
  assign n47431 = pi316 & n46096;
  assign n47432 = n46107 & n47431;
  assign n47433 = ~n47430 & ~n47432;
  assign n47434 = ~pi588 & ~n47433;
  assign n47435 = ~pi200 & ~pi308;
  assign n47436 = pi200 & ~pi1037;
  assign n47437 = ~n47435 & ~n47436;
  assign n47438 = ~pi199 & ~n47437;
  assign n47439 = pi199 & ~pi1047;
  assign n47440 = ~n46096 & ~n47439;
  assign n47441 = ~n47438 & n47440;
  assign n47442 = pi424 & n46705;
  assign n47443 = n46934 & n47442;
  assign n47444 = n8830 & ~n47443;
  assign n47445 = ~n47441 & n47444;
  assign n47446 = ~n47434 & n47445;
  assign n47447 = pi777 & n46131;
  assign n47448 = ~pi838 & ~pi1136;
  assign n47449 = pi737 & pi1135;
  assign n47450 = pi1134 & ~n47449;
  assign n47451 = ~n47448 & n47450;
  assign n47452 = n46941 & n47451;
  assign n47453 = ~n47447 & n47452;
  assign n47454 = ~pi648 & pi1135;
  assign n47455 = ~pi619 & ~pi1135;
  assign n47456 = ~pi1134 & ~n47455;
  assign n47457 = ~n47454 & n47456;
  assign n47458 = n46327 & n47457;
  assign n47459 = ~n8830 & ~n47458;
  assign n47460 = ~n47453 & n47459;
  assign po890 = ~n47446 & ~n47460;
  assign n47462 = pi734 & ~po980;
  assign n47463 = ~pi1119 & po980;
  assign n47464 = ~pi962 & ~n47463;
  assign po891 = ~n47462 & n47464;
  assign n47466 = ~pi1109 & po980;
  assign n47467 = ~pi735 & ~po980;
  assign n47468 = ~pi962 & ~n47467;
  assign po892 = ~n47466 & n47468;
  assign n47470 = ~pi1101 & po980;
  assign n47471 = ~pi736 & ~po980;
  assign n47472 = ~pi962 & ~n47471;
  assign po893 = ~n47470 & n47472;
  assign n47474 = pi737 & ~po980;
  assign n47475 = ~pi1122 & po980;
  assign n47476 = ~pi962 & ~n47475;
  assign po894 = ~n47474 & n47476;
  assign n47478 = pi738 & ~po980;
  assign n47479 = ~pi1121 & po980;
  assign n47480 = ~pi962 & ~n47479;
  assign po895 = ~n47478 & n47480;
  assign n47482 = ~pi952 & ~pi1061;
  assign n47483 = n45822 & n47482;
  assign po988 = pi832 & n47483;
  assign n47485 = pi739 & ~po988;
  assign n47486 = pi1108 & po988;
  assign n47487 = ~pi966 & ~n47486;
  assign po896 = n47485 | ~n47487;
  assign n47489 = pi1114 & po988;
  assign n47490 = ~pi741 & ~po988;
  assign n47491 = ~pi966 & ~n47490;
  assign po898 = n47489 | ~n47491;
  assign n47493 = pi1112 & po988;
  assign n47494 = ~pi742 & ~po988;
  assign n47495 = ~pi966 & ~n47494;
  assign po899 = n47493 | ~n47495;
  assign n47497 = pi743 & ~po988;
  assign n47498 = pi1109 & po988;
  assign n47499 = ~pi966 & ~n47498;
  assign po900 = n47497 | ~n47499;
  assign n47501 = pi1131 & po988;
  assign n47502 = ~pi744 & ~po988;
  assign n47503 = ~pi966 & ~n47502;
  assign po901 = n47501 | ~n47503;
  assign n47505 = pi1111 & po988;
  assign n47506 = ~pi745 & ~po988;
  assign n47507 = ~pi966 & ~n47506;
  assign po902 = n47505 | ~n47507;
  assign n47509 = pi746 & ~po988;
  assign n47510 = pi1104 & po988;
  assign n47511 = ~pi966 & ~n47510;
  assign po903 = n47509 | ~n47511;
  assign n47513 = pi801 & n47303;
  assign n47514 = pi773 & n47318;
  assign n47515 = ~n47290 & ~n47514;
  assign n47516 = n47300 & n47515;
  assign n47517 = ~n47513 & ~n47516;
  assign n47518 = ~n47293 & ~n47296;
  assign n47519 = n47335 & n47518;
  assign n47520 = ~n47517 & n47519;
  assign n47521 = ~pi747 & ~n47514;
  assign n47522 = n47281 & n47318;
  assign n47523 = ~n47521 & ~n47522;
  assign po904 = ~n47520 & n47523;
  assign n47525 = pi748 & ~po988;
  assign n47526 = pi1106 & po988;
  assign n47527 = ~pi966 & ~n47526;
  assign po905 = n47525 | ~n47527;
  assign n47529 = pi749 & ~po988;
  assign n47530 = pi1105 & po988;
  assign n47531 = ~pi966 & ~n47530;
  assign po906 = n47529 | ~n47531;
  assign n47533 = pi1130 & po988;
  assign n47534 = ~pi750 & ~po988;
  assign n47535 = ~pi966 & ~n47534;
  assign po907 = n47533 | ~n47535;
  assign n47537 = pi1123 & po988;
  assign n47538 = ~pi751 & ~po988;
  assign n47539 = ~pi966 & ~n47538;
  assign po908 = n47537 | ~n47539;
  assign n47541 = pi1124 & po988;
  assign n47542 = ~pi752 & ~po988;
  assign n47543 = ~pi966 & ~n47542;
  assign po909 = n47541 | ~n47543;
  assign n47545 = pi1117 & po988;
  assign n47546 = ~pi753 & ~po988;
  assign n47547 = ~pi966 & ~n47546;
  assign po910 = n47545 | ~n47547;
  assign n47549 = pi1118 & po988;
  assign n47550 = ~pi754 & ~po988;
  assign n47551 = ~pi966 & ~n47550;
  assign po911 = n47549 | ~n47551;
  assign n47553 = pi1120 & po988;
  assign n47554 = ~pi755 & ~po988;
  assign n47555 = ~pi966 & ~n47554;
  assign po912 = n47553 | ~n47555;
  assign n47557 = pi1119 & po988;
  assign n47558 = ~pi756 & ~po988;
  assign n47559 = ~pi966 & ~n47558;
  assign po913 = n47557 | ~n47559;
  assign n47561 = pi1113 & po988;
  assign n47562 = ~pi757 & ~po988;
  assign n47563 = ~pi966 & ~n47562;
  assign po914 = n47561 | ~n47563;
  assign n47565 = pi758 & ~po988;
  assign n47566 = pi1101 & po988;
  assign n47567 = ~pi966 & ~n47566;
  assign po915 = n47565 | ~n47567;
  assign n47569 = ~pi759 & ~po988;
  assign n47570 = n45827 & n47483;
  assign n47571 = ~n47569 & ~n47570;
  assign po916 = pi966 | n47571;
  assign n47573 = pi1115 & po988;
  assign n47574 = ~pi760 & ~po988;
  assign n47575 = ~pi966 & ~n47574;
  assign po917 = n47573 | ~n47575;
  assign n47577 = pi1121 & po988;
  assign n47578 = ~pi761 & ~po988;
  assign n47579 = ~pi966 & ~n47578;
  assign po918 = n47577 | ~n47579;
  assign n47581 = pi1129 & po988;
  assign n47582 = ~pi762 & ~po988;
  assign n47583 = ~pi966 & ~n47582;
  assign po919 = n47581 | ~n47583;
  assign n47585 = pi763 & ~po988;
  assign n47586 = pi1103 & po988;
  assign n47587 = ~pi966 & ~n47586;
  assign po920 = n47585 | ~n47587;
  assign n47589 = pi764 & ~po988;
  assign n47590 = pi1107 & po988;
  assign n47591 = ~pi966 & ~n47590;
  assign po921 = n47589 | ~n47591;
  assign n47593 = pi765 & ~po978;
  assign n47594 = pi945 & ~n47593;
  assign n47595 = ~pi765 & ~n47292;
  assign n47596 = ~n47295 & n47595;
  assign n47597 = ~n47301 & n47596;
  assign n47598 = n47288 & ~n47597;
  assign n47599 = ~n47289 & ~n47598;
  assign n47600 = n47306 & ~n47599;
  assign n47601 = ~pi721 & ~n47600;
  assign n47602 = n47324 & ~n47601;
  assign n47603 = ~n47325 & ~n47602;
  assign n47604 = n47330 & ~n47603;
  assign n47605 = ~n47326 & n47331;
  assign n47606 = ~n47604 & ~n47605;
  assign po963 = n47407 & ~n47606;
  assign n47608 = ~pi765 & ~po963;
  assign n47609 = ~pi945 & ~n47608;
  assign po922 = ~n47594 & ~n47609;
  assign n47611 = pi766 & ~po988;
  assign n47612 = pi1110 & po988;
  assign n47613 = ~pi966 & ~n47612;
  assign po923 = n47611 | ~n47613;
  assign n47615 = pi1116 & po988;
  assign n47616 = ~pi767 & ~po988;
  assign n47617 = ~pi966 & ~n47616;
  assign po924 = n47615 | ~n47617;
  assign n47619 = pi1125 & po988;
  assign n47620 = ~pi768 & ~po988;
  assign n47621 = ~pi966 & ~n47620;
  assign po925 = n47619 | ~n47621;
  assign n47623 = n47325 & n47407;
  assign n47624 = pi794 & ~n47290;
  assign n47625 = ~n47293 & n47624;
  assign n47626 = n47334 & n47625;
  assign n47627 = ~n47304 & n47626;
  assign n47628 = ~pi775 & n47627;
  assign n47629 = ~n47623 & ~n47628;
  assign n47630 = pi795 & ~n47629;
  assign n47631 = pi775 & n47281;
  assign n47632 = pi769 & ~n47631;
  assign n47633 = ~pi769 & n47631;
  assign n47634 = ~n47632 & ~n47633;
  assign n47635 = n47319 & ~n47634;
  assign n47636 = ~n47630 & n47635;
  assign n47637 = pi769 & ~n47319;
  assign n47638 = ~po978 & n47637;
  assign po926 = n47636 | n47638;
  assign n47640 = pi1126 & po988;
  assign n47641 = ~pi770 & ~po988;
  assign n47642 = ~pi966 & ~n47641;
  assign po927 = n47640 | ~n47642;
  assign n47644 = ~pi945 & pi987;
  assign n47645 = ~po963 & n47644;
  assign n47646 = pi771 & pi945;
  assign n47647 = ~po978 & n47646;
  assign po928 = n47645 | n47647;
  assign n47649 = pi772 & ~po988;
  assign n47650 = pi1102 & po988;
  assign n47651 = ~pi966 & ~n47650;
  assign po929 = n47649 | ~n47651;
  assign n47653 = ~pi801 & n47306;
  assign n47654 = po963 & n47653;
  assign n47655 = n47318 & ~n47654;
  assign n47656 = pi773 & ~po978;
  assign n47657 = ~n47655 & ~n47656;
  assign po930 = ~n47514 & ~n47657;
  assign n47659 = pi1127 & po988;
  assign n47660 = ~pi774 & ~po988;
  assign n47661 = ~pi966 & ~n47660;
  assign po931 = n47659 | ~n47661;
  assign n47663 = pi775 & ~po978;
  assign n47664 = pi731 & ~pi945;
  assign n47665 = pi765 & pi771;
  assign n47666 = n47281 & n47665;
  assign n47667 = pi795 & pi800;
  assign n47668 = pi801 & ~pi816;
  assign n47669 = n47667 & n47668;
  assign n47670 = ~n47333 & n47669;
  assign n47671 = n47305 & n47670;
  assign n47672 = n47666 & ~n47671;
  assign n47673 = ~pi775 & ~n47672;
  assign n47674 = n47664 & ~n47673;
  assign n47675 = ~n47663 & ~n47674;
  assign n47676 = ~n47409 & ~n47666;
  assign n47677 = pi775 & n47664;
  assign n47678 = ~n47676 & n47677;
  assign po932 = ~n47675 & ~n47678;
  assign n47680 = pi1128 & po988;
  assign n47681 = ~pi776 & ~po988;
  assign n47682 = ~pi966 & ~n47681;
  assign po933 = n47680 | ~n47682;
  assign n47684 = pi1122 & po988;
  assign n47685 = ~pi777 & ~po988;
  assign n47686 = ~pi966 & ~n47685;
  assign po934 = n47684 | ~n47686;
  assign n47688 = pi832 & pi956;
  assign n47689 = ~pi1046 & ~pi1083;
  assign n47690 = pi1085 & n47689;
  assign n47691 = n47688 & n47690;
  assign n47692 = ~pi968 & n47691;
  assign n47693 = pi778 & ~n47692;
  assign n47694 = pi1100 & n47692;
  assign po935 = n47693 | n47694;
  assign po936 = ~pi779 | n45884;
  assign po937 = ~pi780 | n45793;
  assign n47698 = pi781 & ~n47692;
  assign n47699 = pi1101 & n47692;
  assign po938 = n47698 | n47699;
  assign n47701 = ~n41736 & ~n45837;
  assign po939 = n45792 | ~n47701;
  assign n47703 = pi783 & ~n47692;
  assign n47704 = pi1109 & n47692;
  assign po940 = n47703 | n47704;
  assign n47706 = pi784 & ~n47692;
  assign n47707 = pi1110 & n47692;
  assign po941 = n47706 | n47707;
  assign n47709 = pi785 & ~n47692;
  assign n47710 = pi1102 & n47692;
  assign po942 = n47709 | n47710;
  assign n47712 = pi24 & ~pi954;
  assign n47713 = pi786 & pi954;
  assign po943 = ~n47712 & ~n47713;
  assign n47715 = pi787 & ~n47692;
  assign n47716 = pi1104 & n47692;
  assign po944 = n47715 | n47716;
  assign n47718 = pi788 & ~n47692;
  assign n47719 = pi1105 & n47692;
  assign po945 = n47718 | n47719;
  assign n47721 = pi789 & ~n47692;
  assign n47722 = pi1106 & n47692;
  assign po946 = n47721 | n47722;
  assign n47724 = pi790 & ~n47692;
  assign n47725 = pi1107 & n47692;
  assign po947 = n47724 | n47725;
  assign n47727 = pi791 & ~n47692;
  assign n47728 = pi1108 & n47692;
  assign po948 = n47727 | n47728;
  assign n47730 = pi792 & ~n47692;
  assign n47731 = pi1103 & n47692;
  assign po949 = n47730 | n47731;
  assign n47733 = pi968 & n47691;
  assign n47734 = pi794 & ~n47733;
  assign n47735 = pi1130 & n47733;
  assign po951 = n47734 | n47735;
  assign n47737 = pi795 & ~n47733;
  assign n47738 = pi1128 & n47733;
  assign po952 = n47737 | n47738;
  assign n47740 = pi266 & ~pi269;
  assign n47741 = pi278 & pi279;
  assign n47742 = ~pi280 & n47741;
  assign n47743 = n47740 & n47742;
  assign n47744 = ~pi281 & n47743;
  assign n47745 = n46076 & n47744;
  assign n47746 = pi264 & ~n47745;
  assign n47747 = ~pi264 & n47745;
  assign po953 = ~n47746 & ~n47747;
  assign n47749 = pi798 & ~n47733;
  assign n47750 = pi1124 & n47733;
  assign po955 = n47749 | n47750;
  assign n47752 = pi799 & ~n47733;
  assign n47753 = ~pi1107 & n47733;
  assign po956 = ~n47752 & ~n47753;
  assign n47755 = pi800 & ~n47733;
  assign n47756 = pi1125 & n47733;
  assign po957 = n47755 | n47756;
  assign n47758 = pi801 & ~n47733;
  assign n47759 = pi1126 & n47733;
  assign po958 = n47758 | n47759;
  assign n47761 = pi803 & ~n47733;
  assign n47762 = ~pi1106 & n47733;
  assign po960 = ~n47761 & ~n47762;
  assign n47764 = pi804 & ~n47733;
  assign n47765 = pi1109 & n47733;
  assign po961 = n47764 | n47765;
  assign n47767 = ~pi282 & n46074;
  assign n47768 = ~pi270 & n47767;
  assign n47769 = pi270 & ~n47767;
  assign po962 = ~n47768 & ~n47769;
  assign n47771 = pi807 & ~n47733;
  assign n47772 = pi1127 & n47733;
  assign po964 = n47771 | n47772;
  assign n47774 = pi808 & ~n47733;
  assign n47775 = pi1101 & n47733;
  assign po965 = n47774 | n47775;
  assign n47777 = pi809 & ~n47733;
  assign n47778 = ~pi1103 & n47733;
  assign po966 = ~n47777 & ~n47778;
  assign n47780 = pi810 & ~n47733;
  assign n47781 = pi1108 & n47733;
  assign po967 = n47780 | n47781;
  assign n47783 = pi811 & ~n47733;
  assign n47784 = pi1102 & n47733;
  assign po968 = n47783 | n47784;
  assign n47786 = pi812 & ~n47733;
  assign n47787 = ~pi1104 & n47733;
  assign po969 = ~n47786 & ~n47787;
  assign n47789 = pi813 & ~n47733;
  assign n47790 = pi1131 & n47733;
  assign po970 = n47789 | n47790;
  assign n47792 = pi814 & ~n47733;
  assign n47793 = ~pi1105 & n47733;
  assign po971 = ~n47792 & ~n47793;
  assign n47795 = pi815 & ~n47733;
  assign n47796 = pi1110 & n47733;
  assign po972 = n47795 | n47796;
  assign n47798 = pi816 & ~n47733;
  assign n47799 = pi1129 & n47733;
  assign po973 = n47798 | n47799;
  assign n47801 = pi269 & ~n46072;
  assign po974 = ~n46073 & ~n47801;
  assign n47803 = n8830 & n14080;
  assign po975 = n13933 | n47803;
  assign n47805 = pi265 & ~n46078;
  assign po976 = ~n46079 & ~n47805;
  assign n47807 = pi277 & ~n47768;
  assign po977 = ~n46077 & ~n47807;
  assign po979 = ~pi811 & ~pi893;
  assign n47810 = ~pi982 & ~n10019;
  assign n47811 = n7536 & n8830;
  assign n47812 = ~n47810 & ~n47811;
  assign po981 = n6257 & ~n47812;
  assign n47814 = pi123 & n3100;
  assign n47815 = pi1131 & ~n47814;
  assign n47816 = pi1127 & ~n47814;
  assign n47817 = ~n47815 & ~n47816;
  assign n47818 = ~pi825 & n47814;
  assign n47819 = n47817 & ~n47818;
  assign n47820 = pi1131 & n47816;
  assign n47821 = ~n47819 & ~n47820;
  assign n47822 = pi1124 & ~pi1130;
  assign n47823 = ~pi1124 & pi1130;
  assign n47824 = ~n47822 & ~n47823;
  assign n47825 = ~pi1128 & ~pi1129;
  assign n47826 = pi1128 & pi1129;
  assign n47827 = ~n47825 & ~n47826;
  assign n47828 = ~pi1125 & ~pi1126;
  assign n47829 = pi1125 & pi1126;
  assign n47830 = ~n47828 & ~n47829;
  assign n47831 = n47827 & ~n47830;
  assign n47832 = ~n47827 & n47830;
  assign n47833 = ~n47831 & ~n47832;
  assign n47834 = n47824 & n47833;
  assign n47835 = ~n47824 & ~n47833;
  assign n47836 = ~n47834 & ~n47835;
  assign n47837 = ~n47821 & ~n47836;
  assign n47838 = pi825 & n47814;
  assign n47839 = n47817 & ~n47838;
  assign n47840 = ~n47820 & n47836;
  assign n47841 = ~n47839 & n47840;
  assign po982 = ~n47837 & ~n47841;
  assign n47843 = pi1123 & ~n47814;
  assign n47844 = pi1122 & ~n47814;
  assign n47845 = ~n47843 & ~n47844;
  assign n47846 = ~pi826 & n47814;
  assign n47847 = n47845 & ~n47846;
  assign n47848 = pi1123 & n47844;
  assign n47849 = ~n47847 & ~n47848;
  assign n47850 = pi1118 & ~pi1119;
  assign n47851 = ~pi1118 & pi1119;
  assign n47852 = ~n47850 & ~n47851;
  assign n47853 = ~pi1120 & ~pi1121;
  assign n47854 = pi1120 & pi1121;
  assign n47855 = ~n47853 & ~n47854;
  assign n47856 = ~pi1116 & ~pi1117;
  assign n47857 = pi1116 & pi1117;
  assign n47858 = ~n47856 & ~n47857;
  assign n47859 = n47855 & ~n47858;
  assign n47860 = ~n47855 & n47858;
  assign n47861 = ~n47859 & ~n47860;
  assign n47862 = n47852 & n47861;
  assign n47863 = ~n47852 & ~n47861;
  assign n47864 = ~n47862 & ~n47863;
  assign n47865 = ~n47849 & ~n47864;
  assign n47866 = pi826 & n47814;
  assign n47867 = n47845 & ~n47866;
  assign n47868 = ~n47848 & n47864;
  assign n47869 = ~n47867 & n47868;
  assign po983 = ~n47865 & ~n47869;
  assign n47871 = pi1100 & ~n47814;
  assign n47872 = pi1107 & ~n47814;
  assign n47873 = ~n47871 & ~n47872;
  assign n47874 = ~pi827 & n47814;
  assign n47875 = n47873 & ~n47874;
  assign n47876 = pi1100 & n47872;
  assign n47877 = ~n47875 & ~n47876;
  assign n47878 = pi1103 & ~pi1105;
  assign n47879 = ~pi1103 & pi1105;
  assign n47880 = ~n47878 & ~n47879;
  assign n47881 = ~pi1101 & ~pi1102;
  assign n47882 = pi1101 & pi1102;
  assign n47883 = ~n47881 & ~n47882;
  assign n47884 = ~pi1104 & ~pi1106;
  assign n47885 = pi1104 & pi1106;
  assign n47886 = ~n47884 & ~n47885;
  assign n47887 = n47883 & ~n47886;
  assign n47888 = ~n47883 & n47886;
  assign n47889 = ~n47887 & ~n47888;
  assign n47890 = n47880 & n47889;
  assign n47891 = ~n47880 & ~n47889;
  assign n47892 = ~n47890 & ~n47891;
  assign n47893 = ~n47877 & ~n47892;
  assign n47894 = pi827 & n47814;
  assign n47895 = n47873 & ~n47894;
  assign n47896 = ~n47876 & n47892;
  assign n47897 = ~n47895 & n47896;
  assign po984 = ~n47893 & ~n47897;
  assign n47899 = pi1115 & ~n47814;
  assign n47900 = pi1114 & ~n47814;
  assign n47901 = ~n47899 & ~n47900;
  assign n47902 = ~pi828 & n47814;
  assign n47903 = n47901 & ~n47902;
  assign n47904 = pi1115 & n47900;
  assign n47905 = ~n47903 & ~n47904;
  assign n47906 = pi1110 & ~pi1111;
  assign n47907 = ~pi1110 & pi1111;
  assign n47908 = ~n47906 & ~n47907;
  assign n47909 = ~pi1112 & ~pi1113;
  assign n47910 = pi1112 & pi1113;
  assign n47911 = ~n47909 & ~n47910;
  assign n47912 = ~pi1108 & ~pi1109;
  assign n47913 = pi1108 & pi1109;
  assign n47914 = ~n47912 & ~n47913;
  assign n47915 = n47911 & ~n47914;
  assign n47916 = ~n47911 & n47914;
  assign n47917 = ~n47915 & ~n47916;
  assign n47918 = n47908 & n47917;
  assign n47919 = ~n47908 & ~n47917;
  assign n47920 = ~n47918 & ~n47919;
  assign n47921 = ~n47905 & ~n47920;
  assign n47922 = pi828 & n47814;
  assign n47923 = n47901 & ~n47922;
  assign n47924 = ~n47904 & n47920;
  assign n47925 = ~n47923 & n47924;
  assign po985 = ~n47921 & ~n47925;
  assign n47927 = n8830 & n10018;
  assign n47928 = pi951 & ~n47927;
  assign po986 = pi1092 & ~n47928;
  assign n47930 = pi281 & ~n47743;
  assign po987 = ~n47744 & ~n47930;
  assign n47932 = ~pi832 & pi1091;
  assign n47933 = pi1162 & n47932;
  assign po989 = n8834 & n47933;
  assign n47935 = pi833 & ~n2754;
  assign po990 = n16993 | n47935;
  assign po991 = pi946 & n2754;
  assign n47938 = pi282 & ~n46074;
  assign po992 = ~n47767 & ~n47938;
  assign n47940 = ~pi955 & pi1049;
  assign n47941 = pi837 & pi955;
  assign po993 = n47940 | n47941;
  assign n47943 = ~pi955 & pi1047;
  assign n47944 = pi838 & pi955;
  assign po994 = n47943 | n47944;
  assign n47946 = ~pi955 & pi1074;
  assign n47947 = pi839 & pi955;
  assign po995 = n47946 | n47947;
  assign n47949 = pi840 & ~n2754;
  assign n47950 = pi1196 & n2754;
  assign po996 = n47949 | n47950;
  assign po997 = ~pi33 & n8938;
  assign n47953 = ~pi955 & pi1035;
  assign n47954 = pi842 & pi955;
  assign po998 = n47953 | n47954;
  assign n47956 = ~pi955 & pi1079;
  assign n47957 = pi843 & pi955;
  assign po999 = n47956 | n47957;
  assign n47959 = ~pi955 & pi1078;
  assign n47960 = pi844 & pi955;
  assign po1000 = n47959 | n47960;
  assign n47962 = ~pi955 & pi1043;
  assign n47963 = pi845 & pi955;
  assign po1001 = n47962 | n47963;
  assign n47965 = pi846 & ~n42290;
  assign n47966 = pi1134 & n42290;
  assign po1002 = n47965 | n47966;
  assign n47968 = ~pi955 & pi1055;
  assign n47969 = pi847 & pi955;
  assign po1003 = n47968 | n47969;
  assign n47971 = ~pi955 & pi1039;
  assign n47972 = pi848 & pi955;
  assign po1004 = n47971 | n47972;
  assign n47974 = pi849 & ~n2754;
  assign n47975 = pi1198 & n2754;
  assign po1005 = n47974 | n47975;
  assign n47977 = ~pi955 & pi1048;
  assign n47978 = pi850 & pi955;
  assign po1006 = n47977 | n47978;
  assign n47980 = ~pi955 & pi1045;
  assign n47981 = pi851 & pi955;
  assign po1007 = n47980 | n47981;
  assign n47983 = ~pi955 & pi1062;
  assign n47984 = pi852 & pi955;
  assign po1008 = n47983 | n47984;
  assign n47986 = ~pi955 & pi1080;
  assign n47987 = pi853 & pi955;
  assign po1009 = n47986 | n47987;
  assign n47989 = ~pi955 & pi1051;
  assign n47990 = pi854 & pi955;
  assign po1010 = n47989 | n47990;
  assign n47992 = ~pi955 & pi1065;
  assign n47993 = pi855 & pi955;
  assign po1011 = n47992 | n47993;
  assign n47995 = ~pi955 & pi1067;
  assign n47996 = pi856 & pi955;
  assign po1012 = n47995 | n47996;
  assign n47998 = ~pi955 & pi1058;
  assign n47999 = pi857 & pi955;
  assign po1013 = n47998 | n47999;
  assign n48001 = ~pi955 & pi1087;
  assign n48002 = pi858 & pi955;
  assign po1014 = n48001 | n48002;
  assign n48004 = ~pi955 & pi1070;
  assign n48005 = pi859 & pi955;
  assign po1015 = n48004 | n48005;
  assign n48007 = ~pi955 & pi1076;
  assign n48008 = pi860 & pi955;
  assign po1016 = n48007 | n48008;
  assign n48010 = pi1093 & pi1141;
  assign n48011 = pi861 & ~pi1093;
  assign n48012 = ~n48010 & ~n48011;
  assign n48013 = ~pi228 & ~n48012;
  assign n48014 = pi123 & ~pi861;
  assign n48015 = ~pi123 & ~pi1141;
  assign n48016 = pi228 & ~n48015;
  assign n48017 = ~n48014 & n48016;
  assign po1017 = n48013 | n48017;
  assign n48019 = pi862 & ~n42290;
  assign n48020 = pi1139 & n42290;
  assign po1018 = n48019 | n48020;
  assign n48022 = pi863 & ~n2754;
  assign n48023 = pi1199 & n2754;
  assign po1019 = n48022 | n48023;
  assign n48025 = pi864 & ~n2754;
  assign n48026 = pi1197 & n2754;
  assign po1020 = n48025 | n48026;
  assign n48028 = ~pi955 & pi1040;
  assign n48029 = pi865 & pi955;
  assign po1021 = n48028 | n48029;
  assign n48031 = ~pi955 & pi1053;
  assign n48032 = pi866 & pi955;
  assign po1022 = n48031 | n48032;
  assign n48034 = ~pi955 & pi1057;
  assign n48035 = pi867 & pi955;
  assign po1023 = n48034 | n48035;
  assign n48037 = ~pi955 & pi1063;
  assign n48038 = pi868 & pi955;
  assign po1024 = n48037 | n48038;
  assign n48040 = pi1093 & pi1140;
  assign n48041 = pi869 & ~pi1093;
  assign n48042 = ~n48040 & ~n48041;
  assign n48043 = ~pi228 & ~n48042;
  assign n48044 = pi123 & ~pi869;
  assign n48045 = ~pi123 & ~pi1140;
  assign n48046 = pi228 & ~n48045;
  assign n48047 = ~n48044 & n48046;
  assign po1025 = n48043 | n48047;
  assign n48049 = ~pi955 & pi1069;
  assign n48050 = pi870 & pi955;
  assign po1026 = n48049 | n48050;
  assign n48052 = ~pi955 & pi1072;
  assign n48053 = pi871 & pi955;
  assign po1027 = n48052 | n48053;
  assign n48055 = ~pi955 & pi1084;
  assign n48056 = pi872 & pi955;
  assign po1028 = n48055 | n48056;
  assign n48058 = ~pi955 & pi1044;
  assign n48059 = pi873 & pi955;
  assign po1029 = n48058 | n48059;
  assign n48061 = ~pi955 & pi1036;
  assign n48062 = pi874 & pi955;
  assign po1030 = n48061 | n48062;
  assign n48064 = pi1093 & ~pi1136;
  assign n48065 = ~pi875 & ~pi1093;
  assign n48066 = ~n48064 & ~n48065;
  assign n48067 = ~pi228 & ~n48066;
  assign n48068 = pi123 & pi875;
  assign n48069 = ~pi123 & pi1136;
  assign n48070 = pi228 & ~n48069;
  assign n48071 = ~n48068 & n48070;
  assign po1031 = ~n48067 & ~n48071;
  assign n48073 = ~pi955 & pi1037;
  assign n48074 = pi876 & pi955;
  assign po1032 = n48073 | n48074;
  assign n48076 = pi1093 & pi1138;
  assign n48077 = pi877 & ~pi1093;
  assign n48078 = ~n48076 & ~n48077;
  assign n48079 = ~pi228 & ~n48078;
  assign n48080 = pi123 & ~pi877;
  assign n48081 = ~pi123 & ~pi1138;
  assign n48082 = pi228 & ~n48081;
  assign n48083 = ~n48080 & n48082;
  assign po1033 = n48079 | n48083;
  assign n48085 = pi1093 & pi1137;
  assign n48086 = pi878 & ~pi1093;
  assign n48087 = ~n48085 & ~n48086;
  assign n48088 = ~pi228 & ~n48087;
  assign n48089 = pi123 & ~pi878;
  assign n48090 = ~pi123 & ~pi1137;
  assign n48091 = pi228 & ~n48090;
  assign n48092 = ~n48089 & n48091;
  assign po1034 = n48088 | n48092;
  assign n48094 = pi1093 & pi1135;
  assign n48095 = pi879 & ~pi1093;
  assign n48096 = ~n48094 & ~n48095;
  assign n48097 = ~pi228 & ~n48096;
  assign n48098 = pi123 & ~pi879;
  assign n48099 = ~pi123 & ~pi1135;
  assign n48100 = pi228 & ~n48099;
  assign n48101 = ~n48098 & n48100;
  assign po1035 = n48097 | n48101;
  assign n48103 = ~pi955 & pi1081;
  assign n48104 = pi880 & pi955;
  assign po1036 = n48103 | n48104;
  assign n48106 = ~pi955 & pi1059;
  assign n48107 = pi881 & pi955;
  assign po1037 = n48106 | n48107;
  assign n48109 = ~pi883 & n47814;
  assign po1039 = n47872 | n48109;
  assign n48111 = pi1124 & ~n47814;
  assign n48112 = ~pi884 & n47814;
  assign po1040 = n48111 | n48112;
  assign n48114 = pi1125 & ~n47814;
  assign n48115 = ~pi885 & n47814;
  assign po1041 = n48114 | n48115;
  assign n48117 = pi1109 & ~n47814;
  assign n48118 = ~pi886 & n47814;
  assign po1042 = n48117 | n48118;
  assign n48120 = ~pi887 & n47814;
  assign po1043 = n47871 | n48120;
  assign n48122 = pi1120 & ~n47814;
  assign n48123 = ~pi888 & n47814;
  assign po1044 = n48122 | n48123;
  assign n48125 = pi1103 & ~n47814;
  assign n48126 = ~pi889 & n47814;
  assign po1045 = n48125 | n48126;
  assign n48128 = pi1126 & ~n47814;
  assign n48129 = ~pi890 & n47814;
  assign po1046 = n48128 | n48129;
  assign n48131 = pi1116 & ~n47814;
  assign n48132 = ~pi891 & n47814;
  assign po1047 = n48131 | n48132;
  assign n48134 = pi1101 & ~n47814;
  assign n48135 = ~pi892 & n47814;
  assign po1048 = n48134 | n48135;
  assign n48137 = pi1119 & ~n47814;
  assign n48138 = ~pi894 & n47814;
  assign po1050 = n48137 | n48138;
  assign n48140 = pi1113 & ~n47814;
  assign n48141 = ~pi895 & n47814;
  assign po1051 = n48140 | n48141;
  assign n48143 = pi1118 & ~n47814;
  assign n48144 = ~pi896 & n47814;
  assign po1052 = n48143 | n48144;
  assign n48146 = pi1129 & ~n47814;
  assign n48147 = ~pi898 & n47814;
  assign po1054 = n48146 | n48147;
  assign n48149 = ~pi899 & n47814;
  assign po1055 = n47899 | n48149;
  assign n48151 = pi1110 & ~n47814;
  assign n48152 = ~pi900 & n47814;
  assign po1056 = n48151 | n48152;
  assign n48154 = pi1111 & ~n47814;
  assign n48155 = ~pi902 & n47814;
  assign po1058 = n48154 | n48155;
  assign n48157 = pi1121 & ~n47814;
  assign n48158 = ~pi903 & n47814;
  assign po1059 = n48157 | n48158;
  assign n48160 = ~pi904 & n47814;
  assign po1060 = n47816 | n48160;
  assign n48162 = ~pi905 & n47814;
  assign po1061 = n47815 | n48162;
  assign n48164 = pi1128 & ~n47814;
  assign n48165 = ~pi906 & n47814;
  assign po1062 = n48164 | n48165;
  assign n48167 = ~pi604 & ~pi979;
  assign n48168 = pi615 & pi979;
  assign n48169 = ~n48167 & ~n48168;
  assign n48170 = pi782 & ~n48169;
  assign n48171 = ~pi782 & ~pi907;
  assign n48172 = ~pi598 & pi979;
  assign n48173 = ~pi624 & ~pi979;
  assign n48174 = pi782 & ~n48173;
  assign n48175 = ~n48172 & n48174;
  assign n48176 = ~n48171 & ~n48175;
  assign po1063 = ~n48170 & n48176;
  assign n48178 = ~pi908 & n47814;
  assign po1064 = n47844 | n48178;
  assign n48180 = pi1105 & ~n47814;
  assign n48181 = ~pi909 & n47814;
  assign po1065 = n48180 | n48181;
  assign n48183 = pi1117 & ~n47814;
  assign n48184 = ~pi910 & n47814;
  assign po1066 = n48183 | n48184;
  assign n48186 = pi1130 & ~n47814;
  assign n48187 = ~pi911 & n47814;
  assign po1067 = n48186 | n48187;
  assign n48189 = ~pi912 & n47814;
  assign po1068 = n47900 | n48189;
  assign n48191 = pi1106 & ~n47814;
  assign n48192 = ~pi913 & n47814;
  assign po1069 = n48191 | n48192;
  assign n48194 = pi280 & ~n46071;
  assign po1070 = ~n46072 & ~n48194;
  assign n48196 = pi1108 & ~n47814;
  assign n48197 = ~pi915 & n47814;
  assign po1071 = n48196 | n48197;
  assign n48199 = ~pi916 & n47814;
  assign po1072 = n47843 | n48199;
  assign n48201 = pi1112 & ~n47814;
  assign n48202 = ~pi917 & n47814;
  assign po1073 = n48201 | n48202;
  assign n48204 = pi1104 & ~n47814;
  assign n48205 = ~pi918 & n47814;
  assign po1074 = n48204 | n48205;
  assign n48207 = pi1102 & ~n47814;
  assign n48208 = ~pi919 & n47814;
  assign po1075 = n48207 | n48208;
  assign n48210 = pi1093 & pi1139;
  assign n48211 = pi920 & ~pi1093;
  assign po1076 = n48210 | n48211;
  assign n48213 = pi921 & ~pi1093;
  assign po1077 = n48040 | n48213;
  assign n48215 = ~pi922 & ~pi1093;
  assign n48216 = pi1093 & ~pi1152;
  assign po1078 = ~n48215 & ~n48216;
  assign n48218 = ~pi923 & ~pi1093;
  assign n48219 = pi1093 & ~pi1154;
  assign po1079 = ~n48218 & ~n48219;
  assign n48221 = ~pi300 & pi301;
  assign n48222 = pi311 & ~pi312;
  assign po1080 = n48221 & n48222;
  assign n48224 = ~pi925 & ~pi1093;
  assign n48225 = pi1093 & ~pi1155;
  assign po1081 = ~n48224 & ~n48225;
  assign n48227 = ~pi926 & ~pi1093;
  assign n48228 = pi1093 & ~pi1157;
  assign po1082 = ~n48227 & ~n48228;
  assign n48230 = ~pi927 & ~pi1093;
  assign n48231 = pi1093 & ~pi1145;
  assign po1083 = ~n48230 & ~n48231;
  assign n48233 = ~pi928 & ~pi1093;
  assign po1084 = ~n48064 & ~n48233;
  assign n48235 = ~pi929 & ~pi1093;
  assign n48236 = pi1093 & ~pi1144;
  assign po1085 = ~n48235 & ~n48236;
  assign n48238 = ~pi930 & ~pi1093;
  assign n48239 = pi1093 & ~pi1134;
  assign po1086 = ~n48238 & ~n48239;
  assign n48241 = ~pi931 & ~pi1093;
  assign n48242 = pi1093 & ~pi1150;
  assign po1087 = ~n48241 & ~n48242;
  assign n48244 = pi932 & ~pi1093;
  assign po1088 = n42279 | n48244;
  assign n48246 = pi933 & ~pi1093;
  assign po1089 = n48085 | n48246;
  assign n48248 = ~pi934 & ~pi1093;
  assign n48249 = pi1093 & ~pi1147;
  assign po1090 = ~n48248 & ~n48249;
  assign n48251 = pi935 & ~pi1093;
  assign po1091 = n48010 | n48251;
  assign n48253 = ~pi936 & ~pi1093;
  assign n48254 = pi1093 & ~pi1149;
  assign po1092 = ~n48253 & ~n48254;
  assign n48256 = ~pi937 & ~pi1093;
  assign n48257 = pi1093 & ~pi1148;
  assign po1093 = ~n48256 & ~n48257;
  assign n48259 = pi938 & ~pi1093;
  assign po1094 = n48094 | n48259;
  assign n48261 = ~pi939 & ~pi1093;
  assign n48262 = pi1093 & ~pi1146;
  assign po1095 = ~n48261 & ~n48262;
  assign n48264 = pi940 & ~pi1093;
  assign po1096 = n48076 | n48264;
  assign n48266 = ~pi941 & ~pi1093;
  assign n48267 = pi1093 & ~pi1153;
  assign po1097 = ~n48266 & ~n48267;
  assign n48269 = ~pi942 & ~pi1093;
  assign n48270 = pi1093 & ~pi1156;
  assign po1098 = ~n48269 & ~n48270;
  assign n48272 = ~pi943 & ~pi1093;
  assign n48273 = pi1093 & ~pi1151;
  assign po1099 = ~n48272 & ~n48273;
  assign n48275 = pi1093 & pi1143;
  assign n48276 = pi944 & ~pi1093;
  assign po1100 = n48275 | n48276;
  assign po1102 = pi230 & n2754;
  assign n48279 = ~pi782 & pi947;
  assign po1103 = n48175 | n48279;
  assign n48281 = ~pi266 & ~pi992;
  assign po1104 = ~n46071 & ~n48281;
  assign n48283 = ~pi313 & ~pi954;
  assign n48284 = pi949 & pi954;
  assign po1105 = n48283 | n48284;
  assign po1107 = ~n7536 & n14166;
  assign n48287 = pi957 & pi1092;
  assign po1112 = pi31 | n48287;
  assign po1115 = ~pi782 & pi960;
  assign po1116 = ~pi230 & pi961;
  assign po1118 = ~pi782 & pi963;
  assign po1122 = ~pi230 & pi967;
  assign po1124 = ~pi230 & pi969;
  assign po1125 = ~pi782 & pi970;
  assign po1126 = ~pi230 & pi971;
  assign po1127 = ~pi782 & pi972;
  assign po1128 = ~pi230 & pi974;
  assign po1129 = ~pi782 & pi975;
  assign po1131 = ~pi230 & pi977;
  assign po1132 = ~pi782 & pi978;
  assign po1133 = pi598 | ~pi615;
  assign po1135 = pi824 & pi1092;
  assign po1137 = pi604 | pi624;
  assign po166 = 1'b1;
  assign po170 = ~pi1090;
  assign po1110 = ~pi954;
  assign po1130 = ~pi278;
  assign po1146 = ~pi915;
  assign po1147 = ~pi825;
  assign po1148 = ~pi826;
  assign po1149 = ~pi913;
  assign po1150 = ~pi894;
  assign po1151 = ~pi905;
  assign po1153 = ~pi890;
  assign po1155 = ~pi906;
  assign po1156 = ~pi896;
  assign po1157 = ~pi909;
  assign po1158 = ~pi911;
  assign po1159 = ~pi908;
  assign po1160 = ~pi891;
  assign po1161 = ~pi902;
  assign po1162 = ~pi903;
  assign po1163 = ~pi883;
  assign po1164 = ~pi888;
  assign po1165 = ~pi919;
  assign po1166 = ~pi886;
  assign po1167 = ~pi912;
  assign po1168 = ~pi895;
  assign po1169 = ~pi916;
  assign po1170 = ~pi889;
  assign po1171 = ~pi900;
  assign po1172 = ~pi885;
  assign po1173 = ~pi904;
  assign po1174 = ~pi899;
  assign po1175 = ~pi918;
  assign po1176 = ~pi898;
  assign po1177 = ~pi917;
  assign po1178 = ~pi827;
  assign po1179 = ~pi887;
  assign po1180 = ~pi884;
  assign po1181 = ~pi910;
  assign po1182 = ~pi828;
  assign po1183 = ~pi892;
  assign po0 = pi668;
  assign po1 = pi672;
  assign po2 = pi664;
  assign po3 = pi667;
  assign po4 = pi676;
  assign po5 = pi673;
  assign po6 = pi675;
  assign po7 = pi666;
  assign po8 = pi679;
  assign po9 = pi674;
  assign po10 = pi663;
  assign po11 = pi670;
  assign po12 = pi677;
  assign po13 = pi682;
  assign po14 = pi671;
  assign po15 = pi678;
  assign po16 = pi718;
  assign po17 = pi707;
  assign po18 = pi708;
  assign po19 = pi713;
  assign po20 = pi711;
  assign po21 = pi716;
  assign po22 = pi733;
  assign po23 = pi712;
  assign po24 = pi689;
  assign po25 = pi717;
  assign po26 = pi692;
  assign po27 = pi719;
  assign po28 = pi722;
  assign po29 = pi714;
  assign po30 = pi720;
  assign po31 = pi685;
  assign po32 = pi837;
  assign po33 = pi850;
  assign po34 = pi872;
  assign po35 = pi871;
  assign po36 = pi881;
  assign po37 = pi866;
  assign po38 = pi876;
  assign po39 = pi873;
  assign po40 = pi874;
  assign po41 = pi859;
  assign po42 = pi855;
  assign po43 = pi852;
  assign po44 = pi870;
  assign po45 = pi848;
  assign po46 = pi865;
  assign po47 = pi856;
  assign po48 = pi853;
  assign po49 = pi847;
  assign po50 = pi857;
  assign po51 = pi854;
  assign po52 = pi858;
  assign po53 = pi845;
  assign po54 = pi838;
  assign po55 = pi842;
  assign po56 = pi843;
  assign po57 = pi839;
  assign po58 = pi844;
  assign po59 = pi868;
  assign po60 = pi851;
  assign po61 = pi867;
  assign po62 = pi880;
  assign po63 = pi860;
  assign po64 = pi1030;
  assign po65 = pi1034;
  assign po66 = pi1015;
  assign po67 = pi1020;
  assign po68 = pi1025;
  assign po69 = pi1005;
  assign po70 = pi996;
  assign po71 = pi1012;
  assign po72 = pi993;
  assign po73 = pi1016;
  assign po74 = pi1021;
  assign po75 = pi1010;
  assign po76 = pi1027;
  assign po77 = pi1018;
  assign po78 = pi1017;
  assign po79 = pi1024;
  assign po80 = pi1009;
  assign po81 = pi1032;
  assign po82 = pi1003;
  assign po83 = pi997;
  assign po84 = pi1013;
  assign po85 = pi1011;
  assign po86 = pi1008;
  assign po87 = pi1019;
  assign po88 = pi1031;
  assign po89 = pi1022;
  assign po90 = pi1000;
  assign po91 = pi1023;
  assign po92 = pi1002;
  assign po93 = pi1026;
  assign po94 = pi1006;
  assign po95 = pi998;
  assign po96 = pi31;
  assign po97 = pi80;
  assign po98 = pi893;
  assign po99 = pi467;
  assign po100 = pi78;
  assign po101 = pi112;
  assign po102 = pi13;
  assign po103 = pi25;
  assign po104 = pi226;
  assign po105 = pi127;
  assign po106 = pi822;
  assign po107 = pi808;
  assign po108 = pi227;
  assign po109 = pi477;
  assign po110 = pi834;
  assign po111 = pi229;
  assign po112 = pi12;
  assign po113 = pi11;
  assign po114 = pi10;
  assign po115 = pi9;
  assign po116 = pi8;
  assign po117 = pi7;
  assign po118 = pi6;
  assign po119 = pi5;
  assign po120 = pi4;
  assign po121 = pi3;
  assign po122 = pi0;
  assign po123 = pi2;
  assign po124 = pi1;
  assign po125 = pi310;
  assign po126 = pi302;
  assign po127 = pi475;
  assign po128 = pi474;
  assign po129 = pi466;
  assign po130 = pi473;
  assign po131 = pi471;
  assign po132 = pi472;
  assign po133 = pi470;
  assign po134 = pi469;
  assign po135 = pi465;
  assign po136 = pi1028;
  assign po137 = pi1033;
  assign po138 = pi995;
  assign po139 = pi994;
  assign po140 = pi28;
  assign po141 = pi27;
  assign po142 = pi26;
  assign po143 = pi29;
  assign po144 = pi15;
  assign po145 = pi14;
  assign po146 = pi21;
  assign po147 = pi20;
  assign po148 = pi19;
  assign po149 = pi18;
  assign po150 = pi17;
  assign po151 = pi16;
  assign po152 = pi1096;
  assign po168 = pi228;
  assign po169 = pi22;
  assign po179 = pi1089;
  assign po180 = pi23;
  assign po181 = po167;
  assign po188 = pi37;
  assign po263 = pi117;
  assign po285 = pi131;
  assign po386 = pi232;
  assign po388 = pi236;
  assign po636 = pi583;
  assign po1053 = pi67;
  assign po1108 = pi1134;
  assign po1109 = pi964;
  assign po1111 = pi965;
  assign po1113 = pi991;
  assign po1114 = pi985;
  assign po1117 = pi1014;
  assign po1119 = pi1029;
  assign po1120 = pi1004;
  assign po1121 = pi1007;
  assign po1123 = pi1135;
  assign po1134 = pi1064;
  assign po1136 = pi299;
  assign po1138 = pi1075;
  assign po1139 = pi1052;
  assign po1140 = pi771;
  assign po1141 = pi765;
  assign po1142 = pi605;
  assign po1143 = pi601;
  assign po1144 = pi278;
  assign po1145 = pi279;
  assign po1152 = pi1095;
  assign po1154 = pi1094;
  assign po1184 = pi1187;
  assign po1185 = pi1172;
  assign po1186 = pi1170;
  assign po1187 = pi1138;
  assign po1188 = pi1177;
  assign po1189 = pi1178;
  assign po1190 = pi863;
  assign po1191 = pi1203;
  assign po1192 = pi1185;
  assign po1193 = pi1171;
  assign po1194 = pi1192;
  assign po1195 = pi1137;
  assign po1196 = pi1186;
  assign po1197 = pi1165;
  assign po1198 = pi1164;
  assign po1199 = pi1098;
  assign po1200 = pi1183;
  assign po1201 = pi230;
  assign po1202 = pi1169;
  assign po1203 = pi1136;
  assign po1204 = pi1181;
  assign po1205 = pi849;
  assign po1206 = pi1193;
  assign po1207 = pi1182;
  assign po1208 = pi1168;
  assign po1209 = pi1175;
  assign po1210 = pi1191;
  assign po1211 = pi1099;
  assign po1212 = pi1174;
  assign po1213 = pi1179;
  assign po1214 = pi1202;
  assign po1215 = pi1176;
  assign po1216 = pi1173;
  assign po1217 = pi1201;
  assign po1218 = pi1167;
  assign po1219 = pi840;
  assign po1220 = pi1189;
  assign po1221 = pi1195;
  assign po1222 = pi864;
  assign po1223 = pi1190;
  assign po1224 = pi1188;
  assign po1225 = pi1180;
  assign po1226 = pi1194;
  assign po1227 = pi1097;
  assign po1228 = pi1166;
  assign po1229 = pi1200;
  assign po1230 = pi1184;
endmodule
