module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 ,
    pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 ,
    pi139 , pi140 , pi141 , pi142 , pi143 , pi144 , pi145 ,
    pi146 , pi147 , pi148 , pi149 , pi150 , pi151 , pi152 ,
    pi153 , pi154 , pi155 , pi156 , pi157 , pi158 , pi159 ,
    pi160 , pi161 , pi162 , pi163 , pi164 , pi165 , pi166 ,
    pi167 , pi168 , pi169 , pi170 , pi171 , pi172 , pi173 ,
    pi174 , pi175 , pi176 , pi177 , pi178 , pi179 , pi180 ,
    pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 ,
    pi188 , pi189 , pi190 , pi191 , pi192 , pi193 , pi194 ,
    pi195 , pi196 , pi197 , pi198 , pi199 , pi200 , pi201 ,
    pi202 , pi203 , pi204 , pi205 , pi206 , pi207 , pi208 ,
    pi209 , pi210 , pi211 , pi212 , pi213 , pi214 , pi215 ,
    pi216 , pi217 , pi218 , pi219 , pi220 , pi221 , pi222 ,
    pi223 , pi224 , pi225 , pi226 , pi227 , pi228 , pi229 ,
    pi230 , pi231 , pi232 , pi233 , pi234 , pi235 , pi236 ,
    pi237 , pi238 , pi239 , pi240 , pi241 , pi242 , pi243 ,
    pi244 , pi245 , pi246 , pi247 , pi248 , pi249 , pi250 ,
    pi251 , pi252 , pi253 , pi254 , pi255 , pi256 , pi257 ,
    pi258 , pi259 , pi260 , pi261 , pi262 , pi263 , pi264 ,
    pi265 , pi266 , pi267 , pi268 , pi269 , pi270 , pi271 ,
    pi272 , pi273 , pi274 , pi275 , pi276 , pi277 , pi278 ,
    pi279 , pi280 , pi281 , pi282 , pi283 , pi284 , pi285 ,
    pi286 , pi287 , pi288 , pi289 , pi290 , pi291 , pi292 ,
    pi293 , pi294 , pi295 , pi296 , pi297 , pi298 , pi299 ,
    pi300 , pi301 , pi302 , pi303 , pi304 , pi305 , pi306 ,
    pi307 , pi308 , pi309 , pi310 , pi311 , pi312 , pi313 ,
    pi314 , pi315 , pi316 , pi317 , pi318 , pi319 , pi320 ,
    pi321 , pi322 , pi323 , pi324 , pi325 , pi326 , pi327 ,
    pi328 , pi329 , pi330 , pi331 , pi332 , pi333 , pi334 ,
    pi335 , pi336 , pi337 , pi338 , pi339 , pi340 , pi341 ,
    pi342 , pi343 , pi344 , pi345 , pi346 , pi347 , pi348 ,
    pi349 , pi350 , pi351 , pi352 , pi353 , pi354 , pi355 ,
    pi356 , pi357 , pi358 , pi359 , pi360 , pi361 , pi362 ,
    pi363 , pi364 , pi365 , pi366 , pi367 , pi368 , pi369 ,
    pi370 , pi371 , pi372 , pi373 , pi374 , pi375 , pi376 ,
    pi377 , pi378 , pi379 , pi380 , pi381 , pi382 , pi383 ,
    pi384 , pi385 , pi386 , pi387 , pi388 , pi389 , pi390 ,
    pi391 , pi392 , pi393 , pi394 , pi395 , pi396 , pi397 ,
    pi398 , pi399 , pi400 , pi401 , pi402 , pi403 , pi404 ,
    pi405 , pi406 , pi407 , pi408 , pi409 , pi410 , pi411 ,
    pi412 , pi413 , pi414 , pi415 , pi416 , pi417 , pi418 ,
    pi419 , pi420 , pi421 , pi422 , pi423 , pi424 , pi425 ,
    pi426 , pi427 , pi428 , pi429 , pi430 , pi431 , pi432 ,
    pi433 , pi434 , pi435 , pi436 , pi437 , pi438 , pi439 ,
    pi440 , pi441 , pi442 , pi443 , pi444 , pi445 , pi446 ,
    pi447 , pi448 , pi449 , pi450 , pi451 , pi452 , pi453 ,
    pi454 , pi455 , pi456 , pi457 , pi458 , pi459 , pi460 ,
    pi461 , pi462 , pi463 , pi464 , pi465 , pi466 , pi467 ,
    pi468 , pi469 , pi470 , pi471 , pi472 , pi473 , pi474 ,
    pi475 , pi476 , pi477 , pi478 , pi479 , pi480 , pi481 ,
    pi482 , pi483 , pi484 , pi485 , pi486 , pi487 , pi488 ,
    pi489 , pi490 , pi491 , pi492 , pi493 , pi494 , pi495 ,
    pi496 , pi497 , pi498 , pi499 , pi500 , pi501 , pi502 ,
    pi503 , pi504 , pi505 , pi506 , pi507 , pi508 , pi509 ,
    pi510 , pi511 , pi512 , pi513 , pi514 , pi515 , pi516 ,
    pi517 , pi518 , pi519 , pi520 , pi521 , pi522 , pi523 ,
    pi524 , pi525 , pi526 , pi527 , pi528 , pi529 , pi530 ,
    pi531 , pi532 , pi533 , pi534 , pi535 , pi536 , pi537 ,
    pi538 , pi539 , pi540 , pi541 , pi542 , pi543 , pi544 ,
    pi545 , pi546 , pi547 , pi548 , pi549 , pi550 , pi551 ,
    pi552 , pi553 , pi554 , pi555 , pi556 , pi557 , pi558 ,
    pi559 , pi560 , pi561 , pi562 , pi563 , pi564 , pi565 ,
    pi566 , pi567 , pi568 , pi569 , pi570 , pi571 , pi572 ,
    pi573 , pi574 , pi575 , pi576 , pi577 , pi578 , pi579 ,
    pi580 , pi581 , pi582 , pi583 , pi584 , pi585 , pi586 ,
    pi587 , pi588 , pi589 , pi590 , pi591 , pi592 , pi593 ,
    pi594 , pi595 , pi596 , pi597 , pi598 , pi599 , pi600 ,
    pi601 , pi602 , pi603 , pi604 , pi605 , pi606 , pi607 ,
    pi608 , pi609 , pi610 , pi611 , pi612 , pi613 , pi614 ,
    pi615 , pi616 , pi617 , pi618 , pi619 , pi620 , pi621 ,
    pi622 , pi623 , pi624 , pi625 , pi626 , pi627 , pi628 ,
    pi629 , pi630 , pi631 , pi632 , pi633 , pi634 , pi635 ,
    pi636 , pi637 , pi638 , pi639 , pi640 , pi641 , pi642 ,
    pi643 , pi644 , pi645 , pi646 , pi647 , pi648 , pi649 ,
    pi650 , pi651 , pi652 , pi653 , pi654 , pi655 , pi656 ,
    pi657 , pi658 , pi659 , pi660 , pi661 , pi662 , pi663 ,
    pi664 , pi665 , pi666 , pi667 , pi668 , pi669 , pi670 ,
    pi671 , pi672 , pi673 , pi674 , pi675 , pi676 , pi677 ,
    pi678 , pi679 , pi680 , pi681 , pi682 , pi683 , pi684 ,
    pi685 , pi686 , pi687 , pi688 , pi689 , pi690 , pi691 ,
    pi692 , pi693 , pi694 , pi695 , pi696 , pi697 , pi698 ,
    pi699 , pi700 , pi701 , pi702 , pi703 , pi704 , pi705 ,
    pi706 , pi707 , pi708 , pi709 , pi710 , pi711 , pi712 ,
    pi713 , pi714 , pi715 , pi716 , pi717 , pi718 , pi719 ,
    pi720 , pi721 , pi722 , pi723 , pi724 , pi725 , pi726 ,
    pi727 , pi728 , pi729 , pi730 , pi731 , pi732 , pi733 ,
    pi734 , pi735 , pi736 , pi737 , pi738 , pi739 , pi740 ,
    pi741 , pi742 , pi743 , pi744 , pi745 , pi746 , pi747 ,
    pi748 , pi749 , pi750 , pi751 , pi752 , pi753 , pi754 ,
    pi755 , pi756 , pi757 , pi758 , pi759 , pi760 , pi761 ,
    pi762 , pi763 , pi764 , pi765 , pi766 , pi767 , pi768 ,
    pi769 , pi770 , pi771 , pi772 , pi773 , pi774 , pi775 ,
    pi776 , pi777 , pi778 , pi779 , pi780 , pi781 , pi782 ,
    pi783 , pi784 , pi785 , pi786 , pi787 , pi788 , pi789 ,
    pi790 , pi791 , pi792 , pi793 , pi794 , pi795 , pi796 ,
    pi797 , pi798 , pi799 , pi800 , pi801 , pi802 , pi803 ,
    pi804 , pi805 , pi806 , pi807 , pi808 , pi809 , pi810 ,
    pi811 , pi812 , pi813 , pi814 , pi815 , pi816 , pi817 ,
    pi818 , pi819 , pi820 , pi821 , pi822 , pi823 , pi824 ,
    pi825 , pi826 , pi827 , pi828 , pi829 , pi830 , pi831 ,
    pi832 , pi833 , pi834 , pi835 , pi836 , pi837 , pi838 ,
    pi839 , pi840 , pi841 , pi842 , pi843 , pi844 , pi845 ,
    pi846 , pi847 , pi848 , pi849 , pi850 , pi851 , pi852 ,
    pi853 , pi854 , pi855 , pi856 , pi857 , pi858 , pi859 ,
    pi860 , pi861 , pi862 , pi863 , pi864 , pi865 , pi866 ,
    pi867 , pi868 , pi869 , pi870 , pi871 , pi872 , pi873 ,
    pi874 , pi875 , pi876 , pi877 , pi878 , pi879 , pi880 ,
    pi881 , pi882 , pi883 , pi884 , pi885 , pi886 , pi887 ,
    pi888 , pi889 , pi890 , pi891 , pi892 , pi893 , pi894 ,
    pi895 , pi896 , pi897 , pi898 , pi899 , pi900 , pi901 ,
    pi902 , pi903 , pi904 , pi905 , pi906 , pi907 , pi908 ,
    pi909 , pi910 , pi911 , pi912 , pi913 , pi914 , pi915 ,
    pi916 , pi917 , pi918 , pi919 , pi920 , pi921 , pi922 ,
    pi923 , pi924 , pi925 , pi926 , pi927 , pi928 , pi929 ,
    pi930 , pi931 , pi932 , pi933 , pi934 , pi935 , pi936 ,
    pi937 , pi938 , pi939 , pi940 , pi941 , pi942 , pi943 ,
    pi944 , pi945 , pi946 , pi947 , pi948 , pi949 , pi950 ,
    pi951 , pi952 , pi953 , pi954 , pi955 , pi956 , pi957 ,
    pi958 , pi959 , pi960 , pi961 , pi962 , pi963 , pi964 ,
    pi965 , pi966 , pi967 , pi968 , pi969 , pi970 , pi971 ,
    pi972 , pi973 , pi974 , pi975 , pi976 , pi977 , pi978 ,
    pi979 , pi980 , pi981 , pi982 , pi983 , pi984 , pi985 ,
    pi986 , pi987 , pi988 , pi989 , pi990 , pi991 , pi992 ,
    pi993 , pi994 , pi995 , pi996 , pi997 , pi998 , pi999 ,
    pi1000 ,
    po0  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 , pi130 ,
    pi131 , pi132 , pi133 , pi134 , pi135 , pi136 , pi137 ,
    pi138 , pi139 , pi140 , pi141 , pi142 , pi143 , pi144 ,
    pi145 , pi146 , pi147 , pi148 , pi149 , pi150 , pi151 ,
    pi152 , pi153 , pi154 , pi155 , pi156 , pi157 , pi158 ,
    pi159 , pi160 , pi161 , pi162 , pi163 , pi164 , pi165 ,
    pi166 , pi167 , pi168 , pi169 , pi170 , pi171 , pi172 ,
    pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 ,
    pi180 , pi181 , pi182 , pi183 , pi184 , pi185 , pi186 ,
    pi187 , pi188 , pi189 , pi190 , pi191 , pi192 , pi193 ,
    pi194 , pi195 , pi196 , pi197 , pi198 , pi199 , pi200 ,
    pi201 , pi202 , pi203 , pi204 , pi205 , pi206 , pi207 ,
    pi208 , pi209 , pi210 , pi211 , pi212 , pi213 , pi214 ,
    pi215 , pi216 , pi217 , pi218 , pi219 , pi220 , pi221 ,
    pi222 , pi223 , pi224 , pi225 , pi226 , pi227 , pi228 ,
    pi229 , pi230 , pi231 , pi232 , pi233 , pi234 , pi235 ,
    pi236 , pi237 , pi238 , pi239 , pi240 , pi241 , pi242 ,
    pi243 , pi244 , pi245 , pi246 , pi247 , pi248 , pi249 ,
    pi250 , pi251 , pi252 , pi253 , pi254 , pi255 , pi256 ,
    pi257 , pi258 , pi259 , pi260 , pi261 , pi262 , pi263 ,
    pi264 , pi265 , pi266 , pi267 , pi268 , pi269 , pi270 ,
    pi271 , pi272 , pi273 , pi274 , pi275 , pi276 , pi277 ,
    pi278 , pi279 , pi280 , pi281 , pi282 , pi283 , pi284 ,
    pi285 , pi286 , pi287 , pi288 , pi289 , pi290 , pi291 ,
    pi292 , pi293 , pi294 , pi295 , pi296 , pi297 , pi298 ,
    pi299 , pi300 , pi301 , pi302 , pi303 , pi304 , pi305 ,
    pi306 , pi307 , pi308 , pi309 , pi310 , pi311 , pi312 ,
    pi313 , pi314 , pi315 , pi316 , pi317 , pi318 , pi319 ,
    pi320 , pi321 , pi322 , pi323 , pi324 , pi325 , pi326 ,
    pi327 , pi328 , pi329 , pi330 , pi331 , pi332 , pi333 ,
    pi334 , pi335 , pi336 , pi337 , pi338 , pi339 , pi340 ,
    pi341 , pi342 , pi343 , pi344 , pi345 , pi346 , pi347 ,
    pi348 , pi349 , pi350 , pi351 , pi352 , pi353 , pi354 ,
    pi355 , pi356 , pi357 , pi358 , pi359 , pi360 , pi361 ,
    pi362 , pi363 , pi364 , pi365 , pi366 , pi367 , pi368 ,
    pi369 , pi370 , pi371 , pi372 , pi373 , pi374 , pi375 ,
    pi376 , pi377 , pi378 , pi379 , pi380 , pi381 , pi382 ,
    pi383 , pi384 , pi385 , pi386 , pi387 , pi388 , pi389 ,
    pi390 , pi391 , pi392 , pi393 , pi394 , pi395 , pi396 ,
    pi397 , pi398 , pi399 , pi400 , pi401 , pi402 , pi403 ,
    pi404 , pi405 , pi406 , pi407 , pi408 , pi409 , pi410 ,
    pi411 , pi412 , pi413 , pi414 , pi415 , pi416 , pi417 ,
    pi418 , pi419 , pi420 , pi421 , pi422 , pi423 , pi424 ,
    pi425 , pi426 , pi427 , pi428 , pi429 , pi430 , pi431 ,
    pi432 , pi433 , pi434 , pi435 , pi436 , pi437 , pi438 ,
    pi439 , pi440 , pi441 , pi442 , pi443 , pi444 , pi445 ,
    pi446 , pi447 , pi448 , pi449 , pi450 , pi451 , pi452 ,
    pi453 , pi454 , pi455 , pi456 , pi457 , pi458 , pi459 ,
    pi460 , pi461 , pi462 , pi463 , pi464 , pi465 , pi466 ,
    pi467 , pi468 , pi469 , pi470 , pi471 , pi472 , pi473 ,
    pi474 , pi475 , pi476 , pi477 , pi478 , pi479 , pi480 ,
    pi481 , pi482 , pi483 , pi484 , pi485 , pi486 , pi487 ,
    pi488 , pi489 , pi490 , pi491 , pi492 , pi493 , pi494 ,
    pi495 , pi496 , pi497 , pi498 , pi499 , pi500 , pi501 ,
    pi502 , pi503 , pi504 , pi505 , pi506 , pi507 , pi508 ,
    pi509 , pi510 , pi511 , pi512 , pi513 , pi514 , pi515 ,
    pi516 , pi517 , pi518 , pi519 , pi520 , pi521 , pi522 ,
    pi523 , pi524 , pi525 , pi526 , pi527 , pi528 , pi529 ,
    pi530 , pi531 , pi532 , pi533 , pi534 , pi535 , pi536 ,
    pi537 , pi538 , pi539 , pi540 , pi541 , pi542 , pi543 ,
    pi544 , pi545 , pi546 , pi547 , pi548 , pi549 , pi550 ,
    pi551 , pi552 , pi553 , pi554 , pi555 , pi556 , pi557 ,
    pi558 , pi559 , pi560 , pi561 , pi562 , pi563 , pi564 ,
    pi565 , pi566 , pi567 , pi568 , pi569 , pi570 , pi571 ,
    pi572 , pi573 , pi574 , pi575 , pi576 , pi577 , pi578 ,
    pi579 , pi580 , pi581 , pi582 , pi583 , pi584 , pi585 ,
    pi586 , pi587 , pi588 , pi589 , pi590 , pi591 , pi592 ,
    pi593 , pi594 , pi595 , pi596 , pi597 , pi598 , pi599 ,
    pi600 , pi601 , pi602 , pi603 , pi604 , pi605 , pi606 ,
    pi607 , pi608 , pi609 , pi610 , pi611 , pi612 , pi613 ,
    pi614 , pi615 , pi616 , pi617 , pi618 , pi619 , pi620 ,
    pi621 , pi622 , pi623 , pi624 , pi625 , pi626 , pi627 ,
    pi628 , pi629 , pi630 , pi631 , pi632 , pi633 , pi634 ,
    pi635 , pi636 , pi637 , pi638 , pi639 , pi640 , pi641 ,
    pi642 , pi643 , pi644 , pi645 , pi646 , pi647 , pi648 ,
    pi649 , pi650 , pi651 , pi652 , pi653 , pi654 , pi655 ,
    pi656 , pi657 , pi658 , pi659 , pi660 , pi661 , pi662 ,
    pi663 , pi664 , pi665 , pi666 , pi667 , pi668 , pi669 ,
    pi670 , pi671 , pi672 , pi673 , pi674 , pi675 , pi676 ,
    pi677 , pi678 , pi679 , pi680 , pi681 , pi682 , pi683 ,
    pi684 , pi685 , pi686 , pi687 , pi688 , pi689 , pi690 ,
    pi691 , pi692 , pi693 , pi694 , pi695 , pi696 , pi697 ,
    pi698 , pi699 , pi700 , pi701 , pi702 , pi703 , pi704 ,
    pi705 , pi706 , pi707 , pi708 , pi709 , pi710 , pi711 ,
    pi712 , pi713 , pi714 , pi715 , pi716 , pi717 , pi718 ,
    pi719 , pi720 , pi721 , pi722 , pi723 , pi724 , pi725 ,
    pi726 , pi727 , pi728 , pi729 , pi730 , pi731 , pi732 ,
    pi733 , pi734 , pi735 , pi736 , pi737 , pi738 , pi739 ,
    pi740 , pi741 , pi742 , pi743 , pi744 , pi745 , pi746 ,
    pi747 , pi748 , pi749 , pi750 , pi751 , pi752 , pi753 ,
    pi754 , pi755 , pi756 , pi757 , pi758 , pi759 , pi760 ,
    pi761 , pi762 , pi763 , pi764 , pi765 , pi766 , pi767 ,
    pi768 , pi769 , pi770 , pi771 , pi772 , pi773 , pi774 ,
    pi775 , pi776 , pi777 , pi778 , pi779 , pi780 , pi781 ,
    pi782 , pi783 , pi784 , pi785 , pi786 , pi787 , pi788 ,
    pi789 , pi790 , pi791 , pi792 , pi793 , pi794 , pi795 ,
    pi796 , pi797 , pi798 , pi799 , pi800 , pi801 , pi802 ,
    pi803 , pi804 , pi805 , pi806 , pi807 , pi808 , pi809 ,
    pi810 , pi811 , pi812 , pi813 , pi814 , pi815 , pi816 ,
    pi817 , pi818 , pi819 , pi820 , pi821 , pi822 , pi823 ,
    pi824 , pi825 , pi826 , pi827 , pi828 , pi829 , pi830 ,
    pi831 , pi832 , pi833 , pi834 , pi835 , pi836 , pi837 ,
    pi838 , pi839 , pi840 , pi841 , pi842 , pi843 , pi844 ,
    pi845 , pi846 , pi847 , pi848 , pi849 , pi850 , pi851 ,
    pi852 , pi853 , pi854 , pi855 , pi856 , pi857 , pi858 ,
    pi859 , pi860 , pi861 , pi862 , pi863 , pi864 , pi865 ,
    pi866 , pi867 , pi868 , pi869 , pi870 , pi871 , pi872 ,
    pi873 , pi874 , pi875 , pi876 , pi877 , pi878 , pi879 ,
    pi880 , pi881 , pi882 , pi883 , pi884 , pi885 , pi886 ,
    pi887 , pi888 , pi889 , pi890 , pi891 , pi892 , pi893 ,
    pi894 , pi895 , pi896 , pi897 , pi898 , pi899 , pi900 ,
    pi901 , pi902 , pi903 , pi904 , pi905 , pi906 , pi907 ,
    pi908 , pi909 , pi910 , pi911 , pi912 , pi913 , pi914 ,
    pi915 , pi916 , pi917 , pi918 , pi919 , pi920 , pi921 ,
    pi922 , pi923 , pi924 , pi925 , pi926 , pi927 , pi928 ,
    pi929 , pi930 , pi931 , pi932 , pi933 , pi934 , pi935 ,
    pi936 , pi937 , pi938 , pi939 , pi940 , pi941 , pi942 ,
    pi943 , pi944 , pi945 , pi946 , pi947 , pi948 , pi949 ,
    pi950 , pi951 , pi952 , pi953 , pi954 , pi955 , pi956 ,
    pi957 , pi958 , pi959 , pi960 , pi961 , pi962 , pi963 ,
    pi964 , pi965 , pi966 , pi967 , pi968 , pi969 , pi970 ,
    pi971 , pi972 , pi973 , pi974 , pi975 , pi976 , pi977 ,
    pi978 , pi979 , pi980 , pi981 , pi982 , pi983 , pi984 ,
    pi985 , pi986 , pi987 , pi988 , pi989 , pi990 , pi991 ,
    pi992 , pi993 , pi994 , pi995 , pi996 , pi997 , pi998 ,
    pi999 , pi1000 ;
  output po0;
  wire n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182,
    n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302,
    n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422,
    n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434,
    n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464,
    n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482,
    n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494,
    n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542,
    n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572,
    n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602,
    n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614,
    n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632,
    n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674,
    n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692,
    n1693, n1694, n1695, n1696, n1697, n1698,
    n1699, n1700, n1701, n1702, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716,
    n1717, n1718, n1719, n1720, n1721, n1722,
    n1723, n1724, n1725, n1726, n1727, n1728,
    n1729, n1730, n1731, n1732, n1733, n1734,
    n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746,
    n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782,
    n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812,
    n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962,
    n1963, n1964, n1965, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986,
    n1987, n1988, n1989, n1990, n1991, n1992,
    n1993, n1994, n1995, n1996, n1997, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016,
    n2017, n2018, n2019, n2020, n2021, n2022,
    n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046,
    n2047, n2048, n2049, n2050, n2051, n2052,
    n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076,
    n2077, n2078, n2079, n2080, n2081, n2082,
    n2083, n2084, n2085, n2086, n2087, n2088,
    n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106,
    n2107, n2108, n2109, n2110, n2111, n2112,
    n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142,
    n2143, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202,
    n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232,
    n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2244,
    n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256,
    n2257, n2258, n2259, n2260, n2261, n2262,
    n2263, n2264, n2265, n2266, n2267, n2268,
    n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286,
    n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376,
    n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388,
    n2389, n2390, n2391, n2392, n2393, n2394,
    n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406,
    n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424,
    n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436,
    n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904,
    n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282,
    n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300,
    n3301, n3302, n3303, n3304, n3305, n3306,
    n3307, n3308, n3309, n3310, n3311, n3312,
    n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324,
    n3325, n3326, n3327, n3328, n3329, n3330,
    n3331, n3332, n3333, n3334, n3335, n3336,
    n3337, n3338, n3339, n3340, n3341, n3342,
    n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354,
    n3355, n3356, n3357, n3358, n3359, n3360,
    n3361, n3362, n3363, n3364, n3365, n3366,
    n3367, n3368, n3369, n3370, n3371, n3372,
    n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384,
    n3385, n3386, n3387, n3388, n3389, n3390,
    n3391, n3392, n3393, n3394, n3395, n3396,
    n3397, n3398, n3399, n3400, n3401, n3402,
    n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414,
    n3415, n3416, n3417, n3418, n3419, n3420,
    n3421, n3422, n3423, n3424, n3425, n3426,
    n3427, n3428, n3429, n3430, n3431, n3432,
    n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444,
    n3445, n3446, n3447, n3448, n3449, n3450,
    n3451, n3452, n3453, n3454, n3455, n3456,
    n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474,
    n3475, n3476, n3477, n3478, n3479, n3480,
    n3481, n3482, n3483, n3484, n3485, n3486,
    n3487, n3488, n3489, n3490, n3491, n3492,
    n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504,
    n3505, n3506, n3507, n3508, n3509, n3510,
    n3511, n3512, n3513, n3514, n3515, n3516,
    n3517, n3518, n3519, n3520, n3521, n3522,
    n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534,
    n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546,
    n3547, n3548, n3549, n3550, n3551, n3552,
    n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564,
    n3565, n3566, n3567, n3568, n3569, n3570,
    n3571, n3572, n3573, n3574, n3575, n3576,
    n3577, n3578, n3579, n3580, n3581, n3582,
    n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594,
    n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3603, n3604, n3605, n3606,
    n3607, n3608, n3609, n3610, n3611, n3612,
    n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624,
    n3625, n3626, n3627, n3628, n3629, n3630,
    n3631, n3632, n3633, n3634, n3635, n3636,
    n3637, n3638, n3639, n3640, n3641, n3642,
    n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654,
    n3655, n3656, n3657, n3658, n3659, n3660,
    n3661, n3662, n3663, n3664, n3665, n3666,
    n3667, n3668, n3669, n3670, n3671, n3672,
    n3673, n3674, n3675, n3676, n3677, n3678,
    n3679, n3680, n3681, n3682, n3683, n3684,
    n3685, n3686, n3687, n3688, n3689, n3690,
    n3691, n3692, n3693, n3694, n3695, n3696,
    n3697, n3698, n3699, n3700, n3701, n3702,
    n3703, n3704, n3705, n3706, n3707, n3708,
    n3709, n3710, n3711, n3712, n3713, n3714,
    n3715, n3716, n3717, n3718, n3719, n3720,
    n3721, n3722, n3723, n3724, n3725, n3726,
    n3727, n3728, n3729, n3730, n3731, n3732,
    n3733, n3734, n3735, n3736, n3737, n3738,
    n3739, n3740, n3741, n3742, n3743, n3744,
    n3745, n3746, n3747, n3748, n3749, n3750,
    n3751, n3752, n3753, n3754, n3755, n3756,
    n3757, n3758, n3759, n3760, n3761, n3762,
    n3763, n3764, n3765, n3766, n3767, n3768,
    n3769, n3770, n3771, n3772, n3773, n3774,
    n3775, n3776, n3777, n3778, n3779, n3780,
    n3781, n3782, n3783, n3784, n3785, n3786,
    n3787, n3788, n3789, n3790, n3791, n3792,
    n3793, n3794, n3795, n3796, n3797, n3798,
    n3799, n3800, n3801, n3802, n3803, n3804,
    n3805, n3806, n3807, n3808, n3809, n3810,
    n3811, n3812, n3813, n3814, n3815, n3816,
    n3817, n3818, n3819, n3820, n3821, n3822,
    n3823, n3824, n3825, n3826, n3827, n3828,
    n3829, n3830, n3831, n3832, n3833, n3834,
    n3835, n3836, n3837, n3838, n3839, n3840,
    n3841, n3842, n3843, n3844, n3845, n3846,
    n3847, n3848, n3849, n3850, n3851, n3852,
    n3853, n3854, n3855, n3856, n3857, n3858,
    n3859, n3860, n3861, n3862, n3863, n3864,
    n3865, n3866, n3867, n3868, n3869, n3870,
    n3871, n3872, n3873, n3874, n3875, n3876,
    n3877, n3878, n3879, n3880, n3881, n3882,
    n3883, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894,
    n3895, n3896, n3897, n3898, n3899, n3900,
    n3901, n3902, n3903, n3904, n3905, n3906,
    n3907, n3908, n3909, n3910, n3911, n3912,
    n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924,
    n3925, n3926, n3927, n3928, n3929, n3930,
    n3931, n3932, n3933, n3934, n3935, n3936,
    n3937, n3938, n3939, n3940, n3941, n3942,
    n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954,
    n3955, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966,
    n3967, n3968, n3969, n3970, n3971, n3972,
    n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990,
    n3991, n3992, n3993, n3994, n3995, n3996,
    n3997, n3998, n3999, n4000, n4001, n4002,
    n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014,
    n4015, n4016, n4017, n4018, n4019, n4020,
    n4021, n4022, n4023, n4024, n4025, n4026,
    n4027, n4028, n4029, n4030, n4031, n4032,
    n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044,
    n4045, n4046, n4047, n4048, n4049, n4050,
    n4051, n4052, n4053, n4054, n4055, n4056,
    n4057, n4058, n4059, n4060, n4061, n4062,
    n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074,
    n4075, n4076, n4077, n4078, n4079, n4080,
    n4081, n4082, n4083, n4084, n4085, n4086,
    n4087, n4088, n4089, n4090, n4091, n4092,
    n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4100, n4101, n4102, n4103, n4104,
    n4105, n4106, n4107, n4108, n4109, n4110,
    n4111, n4112, n4113, n4114, n4115, n4116,
    n4117, n4118, n4119, n4120, n4121, n4122,
    n4123, n4124, n4125, n4126, n4127, n4128,
    n4129, n4130, n4131, n4132, n4133, n4134,
    n4135, n4136, n4137, n4138, n4139, n4140,
    n4141, n4142, n4143, n4144, n4145, n4146,
    n4147, n4148, n4149, n4150, n4151, n4152,
    n4153, n4154, n4155, n4156, n4157, n4158,
    n4159, n4160, n4161, n4162, n4163, n4164,
    n4165, n4166, n4167, n4168, n4169, n4170,
    n4171, n4172, n4173, n4174, n4175, n4176,
    n4177, n4178, n4179, n4180, n4181, n4182,
    n4183, n4184, n4185, n4186, n4187, n4188,
    n4189, n4190, n4191, n4192, n4193, n4194,
    n4195, n4196, n4197, n4198, n4199, n4200,
    n4201, n4202, n4203, n4204, n4205, n4206,
    n4207, n4208, n4209, n4210, n4211, n4212,
    n4213, n4214, n4215, n4216, n4217, n4218,
    n4219, n4220, n4221, n4222, n4223, n4224,
    n4225, n4226, n4227, n4228, n4229, n4230,
    n4231, n4232, n4233, n4234, n4235, n4236,
    n4237, n4238, n4239, n4240, n4241, n4242,
    n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254,
    n4255, n4256, n4257, n4258, n4259, n4260,
    n4261, n4262, n4263, n4264, n4265, n4266,
    n4267, n4268, n4269, n4270, n4271, n4272,
    n4273, n4274, n4275, n4276, n4277, n4278,
    n4279, n4280, n4281, n4282, n4283, n4284,
    n4285, n4286, n4287, n4288, n4289, n4290,
    n4291, n4292, n4293, n4294, n4295, n4296,
    n4297, n4298, n4299, n4300, n4301, n4302,
    n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314,
    n4315, n4316, n4317, n4318, n4319, n4320,
    n4321, n4322, n4323, n4324, n4325, n4326,
    n4327, n4328, n4329, n4330, n4331, n4332,
    n4333, n4334, n4335, n4336, n4337, n4338,
    n4339, n4340, n4341, n4342, n4343, n4344,
    n4345, n4346, n4347, n4348, n4349, n4350,
    n4351, n4352, n4353, n4354, n4355, n4356,
    n4357, n4358, n4359, n4360, n4361, n4362,
    n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392,
    n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422,
    n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476,
    n4477, n4478, n4479, n4480, n4481, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596,
    n4597, n4598, n4599, n4600, n4601, n4602,
    n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626,
    n4627, n4628, n4629, n4630, n4631, n4632,
    n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644,
    n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4659, n4660, n4661, n4662,
    n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674,
    n4675, n4676, n4677, n4678, n4679, n4680,
    n4681, n4682, n4683, n4684, n4685, n4686,
    n4687, n4688, n4689, n4690, n4691, n4692,
    n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704,
    n4705, n4706, n4707, n4708, n4709, n4710,
    n4711, n4712, n4713, n4714, n4715, n4716,
    n4717, n4718, n4719, n4720, n4721, n4722,
    n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734,
    n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4752,
    n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764,
    n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776,
    n4777, n4778, n4779, n4780, n4781, n4782,
    n4783, n4784, n4785, n4786, n4787, n4788,
    n4789, n4790, n4791, n4792, n4793, n4794,
    n4795, n4796, n4797, n4798, n4799, n4800,
    n4801, n4802, n4803, n4804, n4805, n4806,
    n4807, n4808, n4809, n4810, n4811, n4812,
    n4813, n4814, n4815, n4816, n4817, n4818,
    n4819, n4820, n4821, n4822, n4823, n4824,
    n4825, n4826, n4827, n4828, n4829, n4830,
    n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842,
    n4843, n4844, n4845, n4846, n4847, n4848,
    n4849, n4850, n4851, n4852, n4853, n4854,
    n4855, n4856, n4857, n4858, n4859, n4860,
    n4861, n4862, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878,
    n4879, n4880, n4881, n4882, n4883, n4884,
    n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914,
    n4915, n4916, n4917, n4918, n4919, n4920,
    n4921, n4922, n4923, n4924, n4925, n4926,
    n4927, n4928, n4929, n4930, n4931, n4932,
    n4933, n4934, n4935, n4936, n4937, n4938,
    n4939, n4940, n4941, n4942, n4943, n4944,
    n4945, n4946, n4947, n4948, n4949, n4950,
    n4951, n4952, n4953, n4954, n4955, n4956,
    n4957, n4958, n4959, n4960, n4961, n4962,
    n4963, n4964, n4965, n4966, n4967, n4968,
    n4969, n4970, n4971, n4972, n4973, n4974,
    n4975, n4976, n4977, n4978, n4979, n4980,
    n4981, n4982, n4983, n4984, n4985, n4986,
    n4987, n4988, n4989, n4990, n4991, n4992,
    n4993, n4994, n4995, n4996, n4997, n4998,
    n4999, n5000, n5001, n5002, n5003, n5004,
    n5005, n5006, n5007, n5008, n5009, n5010,
    n5011, n5012, n5013, n5014, n5015, n5016,
    n5017, n5018, n5019, n5020, n5021, n5022,
    n5023, n5024, n5025, n5026, n5027, n5028,
    n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5037, n5038, n5039, n5040,
    n5041, n5042, n5043, n5044, n5045, n5046,
    n5047, n5048, n5049, n5050, n5051, n5052,
    n5053, n5054, n5055, n5056, n5057, n5058,
    n5059, n5060, n5061, n5062, n5063, n5064,
    n5065, n5066, n5067, n5068, n5069, n5070,
    n5071, n5072, n5073, n5074, n5075, n5076,
    n5077, n5078, n5079, n5080, n5081, n5082,
    n5083, n5084, n5085, n5086, n5087, n5088,
    n5089, n5090, n5091, n5092, n5093, n5094,
    n5095, n5096, n5097, n5098, n5099, n5100,
    n5101, n5102, n5103, n5104, n5105, n5106,
    n5107, n5108, n5109, n5110, n5111, n5112,
    n5113, n5114, n5115, n5116, n5117, n5118,
    n5119, n5120, n5121, n5122, n5123, n5124,
    n5125, n5126, n5127, n5128, n5129, n5130,
    n5131, n5132, n5133, n5134, n5135, n5136,
    n5137, n5138, n5139, n5140, n5141, n5142,
    n5143, n5144, n5145, n5146, n5147, n5148,
    n5149, n5150, n5151, n5152, n5153, n5154,
    n5155, n5156, n5157, n5158, n5159, n5160,
    n5161, n5162, n5163, n5164, n5165, n5166,
    n5167, n5168, n5169, n5170, n5171, n5172,
    n5173, n5174, n5175, n5176, n5177, n5178,
    n5179, n5180, n5181, n5182, n5183, n5184,
    n5185, n5186, n5187, n5188, n5189, n5190,
    n5191, n5192, n5193, n5194, n5195, n5196,
    n5197, n5198, n5199, n5200, n5201, n5202,
    n5203, n5204, n5205, n5206, n5207, n5208,
    n5209, n5210, n5211, n5212, n5213, n5214,
    n5215, n5216, n5217, n5218, n5219, n5220,
    n5221, n5222, n5223, n5224, n5225, n5226,
    n5227, n5228, n5229, n5230, n5231, n5232,
    n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5244,
    n5245, n5246, n5247, n5248, n5249, n5250,
    n5251, n5252, n5253, n5254, n5255, n5256,
    n5257, n5258, n5259, n5260, n5261, n5262,
    n5263, n5264, n5265, n5266, n5267, n5268,
    n5269, n5270, n5271, n5272, n5273, n5274,
    n5275, n5276, n5277, n5278, n5279, n5280,
    n5281, n5282, n5283, n5284, n5285, n5286,
    n5287, n5288, n5289, n5290, n5291, n5292,
    n5293, n5294, n5295, n5296, n5297, n5298,
    n5299, n5300, n5301, n5302, n5303, n5304,
    n5305, n5306, n5307, n5308, n5309, n5310,
    n5311, n5312, n5313, n5314, n5315, n5316,
    n5317, n5318, n5319, n5320, n5321, n5322,
    n5323, n5324, n5325, n5326, n5327, n5328,
    n5329, n5330, n5331, n5332, n5333, n5334,
    n5335, n5336, n5337, n5338, n5339, n5340,
    n5341, n5342, n5343, n5344, n5345, n5346,
    n5347, n5348, n5349, n5350, n5351, n5352,
    n5353, n5354, n5355, n5356, n5357, n5358,
    n5359, n5360, n5361, n5362, n5363, n5364,
    n5365, n5366, n5367, n5368, n5369, n5370,
    n5371, n5372, n5373, n5374, n5375, n5376,
    n5377, n5378, n5379, n5380, n5381, n5382,
    n5383, n5384, n5385, n5386, n5387, n5388,
    n5389, n5390, n5391, n5392, n5393, n5394,
    n5395, n5396, n5397, n5398, n5399, n5400,
    n5401, n5402, n5403, n5404, n5405, n5406,
    n5407, n5408, n5409, n5410, n5411, n5412,
    n5413, n5414, n5415, n5416, n5417, n5418,
    n5419, n5420, n5421, n5422, n5423, n5424,
    n5425, n5426, n5427, n5428, n5429, n5430,
    n5431, n5432, n5433, n5434, n5435, n5436,
    n5437, n5438, n5439, n5440, n5441, n5442,
    n5443, n5444, n5445, n5446, n5447, n5448,
    n5449, n5450, n5451, n5452, n5453, n5454,
    n5455, n5456, n5457, n5458, n5459, n5460,
    n5461, n5462, n5463, n5464, n5465, n5466,
    n5467, n5468, n5469, n5470, n5471, n5472,
    n5473, n5474, n5475, n5476, n5477, n5478,
    n5479, n5480, n5481, n5482, n5483, n5484,
    n5485, n5486, n5487, n5488, n5489, n5490,
    n5491, n5492, n5493, n5494, n5495, n5496,
    n5497, n5498, n5499, n5500, n5501, n5502,
    n5503, n5504, n5505, n5506, n5507, n5508,
    n5509, n5510, n5511, n5512, n5513, n5514,
    n5515, n5516, n5517, n5518, n5519, n5520,
    n5521, n5522, n5523, n5524, n5525, n5526,
    n5527, n5528, n5529, n5530, n5531, n5532,
    n5533, n5534, n5535, n5536, n5537, n5538,
    n5539, n5540, n5541, n5542, n5543, n5544,
    n5545, n5546, n5547, n5548, n5549, n5550,
    n5551, n5552, n5553, n5554, n5555, n5556,
    n5557, n5558, n5559, n5560, n5561, n5562,
    n5563, n5564, n5565, n5566, n5567, n5568,
    n5569, n5570, n5571, n5572, n5573, n5574,
    n5575, n5576, n5577, n5578, n5579, n5580,
    n5581, n5582, n5583, n5584, n5585, n5586,
    n5587, n5588, n5589, n5590, n5591, n5592,
    n5593, n5594, n5595, n5596, n5597, n5598,
    n5599, n5600, n5601, n5602, n5603, n5604,
    n5605, n5606, n5607, n5608, n5609, n5610,
    n5611, n5612, n5613, n5614, n5615, n5616,
    n5617, n5618, n5619, n5620, n5621, n5622,
    n5623, n5624, n5625, n5626, n5627, n5628,
    n5629, n5630, n5631, n5632, n5633, n5634,
    n5635, n5636, n5637, n5638, n5639, n5640,
    n5641, n5642, n5643, n5644, n5645, n5646,
    n5647, n5648, n5649, n5650, n5651, n5652,
    n5653, n5654, n5655, n5656, n5657, n5658,
    n5659, n5660, n5661, n5662, n5663, n5664,
    n5665, n5666, n5667, n5668, n5669, n5670,
    n5671, n5672, n5673, n5674, n5675, n5676,
    n5677, n5678, n5679, n5680, n5681, n5682,
    n5683, n5684, n5685, n5686, n5687, n5688,
    n5689, n5690, n5691, n5692, n5693, n5694,
    n5695, n5696, n5697, n5698, n5699, n5700,
    n5701, n5702, n5703, n5704, n5705, n5706,
    n5707, n5708, n5709, n5710, n5711, n5712,
    n5713, n5714, n5715, n5716, n5717, n5718,
    n5719, n5720, n5721, n5722, n5723, n5724,
    n5725, n5726, n5727, n5728, n5729, n5730,
    n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742,
    n5743, n5744, n5745, n5746, n5747, n5748,
    n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760,
    n5761, n5762, n5763, n5764, n5765, n5766,
    n5767, n5768, n5769, n5770, n5771, n5772,
    n5773, n5774, n5775, n5776, n5777, n5778,
    n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790,
    n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802,
    n5803, n5804, n5805, n5806, n5807, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814,
    n5815, n5816, n5817, n5818, n5819, n5820,
    n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5830, n5831, n5832,
    n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844,
    n5845, n5846, n5847, n5848, n5849, n5850,
    n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874,
    n5875, n5876, n5877, n5878, n5879, n5880,
    n5881, n5882, n5883, n5884, n5885, n5886,
    n5887, n5888, n5889, n5890, n5891, n5892,
    n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904,
    n5905, n5906, n5907, n5908, n5909, n5910,
    n5911, n5912, n5913, n5914, n5915, n5916,
    n5917, n5918, n5919, n5920, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934,
    n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946,
    n5947, n5948, n5949, n5950, n5951, n5952,
    n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964,
    n5965, n5966, n5967, n5968, n5969, n5970,
    n5971, n5972, n5973, n5974, n5975, n5976,
    n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994,
    n5995, n5996, n5997, n5998, n5999, n6000,
    n6001, n6002, n6003, n6004, n6005, n6006,
    n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6022, n6023, n6024,
    n6025, n6026, n6027, n6028, n6029, n6030,
    n6031, n6032, n6033, n6034, n6035, n6036,
    n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060,
    n6061, n6062, n6063, n6064, n6065, n6066,
    n6067, n6068, n6069, n6070, n6071, n6072,
    n6073, n6074, n6075, n6076, n6077, n6078,
    n6079, n6080, n6081, n6082, n6083, n6084,
    n6085, n6086, n6087, n6088, n6089, n6090,
    n6091, n6092, n6093, n6094, n6095, n6096,
    n6097, n6098, n6099, n6100, n6101, n6102,
    n6103, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114,
    n6115, n6116, n6117, n6118, n6119, n6120,
    n6121, n6122, n6123, n6124, n6125, n6126,
    n6127, n6128, n6129, n6130, n6131, n6132,
    n6133, n6134, n6135, n6136, n6137, n6138,
    n6139, n6140, n6141, n6142, n6143, n6144,
    n6145, n6146, n6147, n6148, n6149, n6150,
    n6151, n6152, n6153, n6154, n6155, n6156,
    n6157, n6158, n6159, n6160, n6161, n6162,
    n6163, n6164, n6165, n6166, n6167, n6168,
    n6169, n6170, n6171, n6172, n6173, n6174,
    n6175, n6176, n6177, n6178, n6179, n6180,
    n6181, n6182, n6183, n6184, n6185, n6186,
    n6187, n6188, n6189, n6190, n6191, n6192,
    n6193, n6194, n6195, n6196, n6197, n6198,
    n6199, n6200, n6201, n6202, n6203, n6204,
    n6205, n6206, n6207, n6208, n6209, n6210,
    n6211, n6212, n6213, n6214, n6215, n6216,
    n6217, n6218, n6219, n6220, n6221, n6222,
    n6223, n6224, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6233, n6234,
    n6235, n6236, n6237, n6238, n6239, n6240,
    n6241, n6242, n6243, n6244, n6245, n6246,
    n6247, n6248, n6249, n6250, n6251, n6252,
    n6253, n6254, n6255, n6256, n6257, n6258,
    n6259, n6260, n6261, n6262, n6263, n6264,
    n6265, n6266, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6274, n6275, n6276,
    n6277, n6278, n6279, n6280, n6281, n6282,
    n6283, n6284, n6285, n6286, n6287, n6288,
    n6289, n6290, n6291, n6292, n6293, n6294,
    n6295, n6296, n6297, n6298, n6299, n6300,
    n6301, n6302, n6303, n6304, n6305, n6306,
    n6307, n6308, n6309, n6310, n6311, n6312,
    n6313, n6314, n6315, n6316, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372,
    n6373, n6374, n6375, n6376, n6377, n6378,
    n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462,
    n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546,
    n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558,
    n6559, n6560, n6561, n6562, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570,
    n6571, n6572, n6573, n6574, n6575, n6576,
    n6577, n6578, n6579, n6580, n6581, n6582,
    n6583, n6584, n6585, n6586, n6587, n6588,
    n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600,
    n6601, n6602, n6603, n6604, n6605, n6606,
    n6607, n6608, n6609, n6610, n6611, n6612,
    n6613, n6614, n6615, n6616, n6617, n6618,
    n6619, n6620, n6621, n6622, n6623, n6624,
    n6625, n6626, n6627, n6628, n6629, n6630,
    n6631, n6632, n6633, n6634, n6635, n6636,
    n6637, n6638, n6639, n6640, n6641, n6642,
    n6643, n6644, n6645, n6646, n6647, n6648,
    n6649, n6650, n6651, n6652, n6653, n6654,
    n6655, n6656, n6657, n6658, n6659, n6660,
    n6661, n6662, n6663, n6664, n6665, n6666,
    n6667, n6668, n6669, n6670, n6671, n6672,
    n6673, n6674, n6675, n6676, n6677, n6678,
    n6679, n6680, n6681, n6682, n6683, n6684,
    n6685, n6686, n6687, n6688, n6689, n6690,
    n6691, n6692, n6693, n6694, n6695, n6696,
    n6697, n6698, n6699, n6700, n6701, n6702,
    n6703, n6704, n6705, n6706, n6707, n6708,
    n6709, n6710, n6711, n6712, n6713, n6714,
    n6715, n6716, n6717, n6718, n6719, n6720,
    n6721, n6722, n6723, n6724, n6725, n6726,
    n6727, n6728, n6729, n6730, n6731, n6732,
    n6733, n6734, n6735, n6736, n6737, n6738,
    n6739, n6740, n6741, n6742, n6743, n6744,
    n6745, n6746, n6747, n6748, n6749, n6750,
    n6751, n6752, n6753, n6754, n6755, n6756,
    n6757, n6758, n6759, n6760, n6761, n6762,
    n6763, n6764, n6765, n6766, n6767, n6768,
    n6769, n6770, n6771, n6772, n6773, n6774,
    n6775, n6776, n6777, n6778, n6779, n6780,
    n6781, n6782, n6783, n6784, n6785, n6786,
    n6787, n6788, n6789, n6790, n6791, n6792,
    n6793, n6794, n6795, n6796, n6797, n6798,
    n6799, n6800, n6801, n6802, n6803, n6804,
    n6805, n6806, n6807, n6808, n6809, n6810,
    n6811, n6812, n6813, n6814, n6815, n6816,
    n6817, n6818, n6819, n6820, n6821, n6822,
    n6823, n6824, n6825, n6826, n6827, n6828,
    n6829, n6830, n6831, n6832, n6833, n6834,
    n6835, n6836, n6837, n6838, n6839, n6840,
    n6841, n6842, n6843, n6844, n6845, n6846,
    n6847, n6848, n6849, n6850, n6851, n6852,
    n6853, n6854, n6855, n6856, n6857, n6858,
    n6859, n6860, n6861, n6862, n6863, n6864,
    n6865, n6866, n6867, n6868, n6869, n6870,
    n6871, n6872, n6873, n6874, n6875, n6876,
    n6877, n6878, n6879, n6880, n6881, n6882,
    n6883, n6884, n6885, n6886, n6887, n6888,
    n6889, n6890, n6891, n6892, n6893, n6894,
    n6895, n6896, n6897, n6898, n6899, n6900,
    n6901, n6902, n6903, n6904, n6905, n6906,
    n6907, n6908, n6909, n6910, n6911, n6912,
    n6913, n6914, n6915, n6916, n6917, n6918,
    n6919, n6920, n6921, n6922, n6923, n6924,
    n6925, n6926, n6927, n6928, n6929, n6930,
    n6931, n6932, n6933, n6934, n6935, n6936,
    n6937, n6938, n6939, n6940, n6941, n6942,
    n6943, n6944, n6945, n6946, n6947, n6948,
    n6949, n6950, n6951, n6952, n6953, n6954,
    n6955, n6956, n6957, n6958, n6959, n6960,
    n6961, n6962, n6963, n6964, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972,
    n6973, n6974, n6975, n6976, n6977, n6978,
    n6979, n6980, n6981, n6982, n6983, n6984,
    n6985, n6986, n6987, n6988, n6989, n6990,
    n6991, n6992, n6993, n6994, n6995, n6996,
    n6997, n6998, n6999, n7000, n7001, n7002,
    n7003, n7004, n7005, n7006, n7007, n7008,
    n7009, n7010, n7011, n7012, n7013, n7014,
    n7015, n7016, n7017, n7018, n7019, n7020,
    n7021, n7022, n7023, n7024, n7025, n7026,
    n7027, n7028, n7029, n7030, n7031, n7032,
    n7033, n7034, n7035, n7036, n7037, n7038,
    n7039, n7040, n7041, n7042, n7043, n7044,
    n7045, n7046, n7047, n7048, n7049, n7050,
    n7051, n7052, n7053, n7054, n7055, n7056,
    n7057, n7058, n7059, n7060, n7061, n7062,
    n7063, n7064, n7065, n7066, n7067, n7068,
    n7069, n7070, n7071, n7072, n7073, n7074,
    n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092,
    n7093, n7094, n7095, n7096, n7097, n7098,
    n7099, n7100, n7101, n7102, n7103, n7104,
    n7105, n7106, n7107, n7108, n7109, n7110,
    n7111, n7112, n7113, n7114, n7115, n7116,
    n7117, n7118, n7119, n7120, n7121, n7122,
    n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7133, n7134,
    n7135, n7136, n7137, n7138, n7139, n7140,
    n7141, n7142, n7143, n7144, n7145, n7146,
    n7147, n7148, n7149, n7150, n7151, n7152,
    n7153, n7154, n7155, n7156, n7157, n7158,
    n7159, n7160, n7161, n7162, n7163, n7164,
    n7165, n7166, n7167, n7168, n7169, n7170,
    n7171, n7172, n7173, n7174, n7175, n7176,
    n7177, n7178, n7179, n7180, n7181, n7182,
    n7183, n7184, n7185, n7186, n7187, n7188,
    n7189, n7190, n7191, n7192, n7193, n7194,
    n7195, n7196, n7197, n7198, n7199, n7200,
    n7201, n7202, n7203, n7204, n7205, n7206,
    n7207, n7208, n7209, n7210, n7211, n7212,
    n7213, n7214, n7215, n7216, n7217, n7218,
    n7219, n7220, n7221, n7222, n7223, n7224,
    n7225, n7226, n7227, n7228, n7229, n7230,
    n7231, n7232, n7233, n7234, n7235, n7236,
    n7237, n7238, n7239, n7240, n7241, n7242,
    n7243, n7244, n7245, n7246, n7247, n7248,
    n7249, n7250, n7251, n7252, n7253, n7254,
    n7255, n7256, n7257, n7258, n7259, n7260,
    n7261, n7262, n7263, n7264, n7265, n7266,
    n7267, n7268, n7269, n7270, n7271, n7272,
    n7273, n7274, n7275, n7276, n7277, n7278,
    n7279, n7280, n7281, n7282, n7283, n7284,
    n7285, n7286, n7287, n7288, n7289, n7290,
    n7291, n7292, n7293, n7294, n7295, n7296,
    n7297, n7298, n7299, n7300, n7301, n7302,
    n7303, n7304, n7305, n7306, n7307, n7308,
    n7309, n7310, n7311, n7312, n7313, n7314,
    n7315, n7316, n7317, n7318, n7319, n7320,
    n7321, n7322, n7323, n7324, n7325, n7326,
    n7327, n7328, n7329, n7330, n7331, n7332,
    n7333, n7334, n7335, n7336, n7337, n7338,
    n7339, n7340, n7341, n7342, n7343, n7344,
    n7345, n7346, n7347, n7348, n7349, n7350,
    n7351, n7352, n7353, n7354, n7355, n7356,
    n7357, n7358, n7359, n7360, n7361, n7362,
    n7363, n7364, n7365, n7366, n7367, n7368,
    n7369, n7370, n7371, n7372, n7373, n7374,
    n7375, n7376, n7377, n7378, n7379, n7380,
    n7381, n7382, n7383, n7384, n7385, n7386,
    n7387, n7388, n7389, n7390, n7391, n7392,
    n7393, n7394, n7395, n7396, n7397, n7398,
    n7399, n7400, n7401, n7402, n7403, n7404,
    n7405, n7406, n7407, n7408, n7409, n7410,
    n7411, n7412, n7413, n7414, n7415, n7416,
    n7417, n7418, n7419, n7420, n7421, n7422,
    n7423, n7424, n7425, n7426, n7427, n7428,
    n7429, n7430, n7431, n7432, n7433, n7434,
    n7435, n7436, n7437, n7438, n7439, n7440,
    n7441, n7442, n7443, n7444, n7445, n7446,
    n7447, n7448, n7449, n7450, n7451, n7452,
    n7453, n7454, n7455, n7456, n7457, n7458,
    n7459, n7460, n7461, n7462, n7463, n7464,
    n7465, n7466, n7467, n7468, n7469, n7470,
    n7471, n7472, n7473, n7474, n7475, n7476,
    n7477, n7478, n7479, n7480, n7481, n7482,
    n7483, n7484, n7485, n7486, n7487, n7488,
    n7489, n7490, n7491, n7492, n7493, n7494,
    n7495, n7496, n7497, n7498, n7499, n7500,
    n7501, n7502, n7503, n7504, n7505, n7506,
    n7507, n7508, n7509, n7510, n7511, n7512,
    n7513, n7514, n7515, n7516, n7517, n7518,
    n7519, n7520, n7521, n7522, n7523, n7524,
    n7525, n7526, n7527, n7528, n7529, n7530,
    n7531, n7532, n7533, n7534, n7535, n7536,
    n7537, n7538, n7539, n7540, n7541, n7542,
    n7543, n7544, n7545, n7546, n7547, n7548,
    n7549, n7550, n7551, n7552, n7553, n7554,
    n7555, n7556, n7557, n7558, n7559, n7560,
    n7561, n7562, n7563, n7564, n7565, n7566,
    n7567, n7568, n7569, n7570, n7571, n7572,
    n7573, n7574, n7575, n7576, n7577, n7578,
    n7579, n7580, n7581, n7582, n7583, n7584,
    n7585, n7586, n7587, n7588, n7589, n7590,
    n7591, n7592, n7593, n7594, n7595, n7596,
    n7597, n7598, n7599, n7600, n7601, n7602,
    n7603, n7604, n7605, n7606, n7607, n7608,
    n7609, n7610, n7611, n7612, n7613, n7614,
    n7615, n7616, n7617, n7618, n7619, n7620,
    n7621, n7622, n7623, n7624, n7625, n7626,
    n7627, n7628, n7629, n7630, n7631, n7632,
    n7633, n7634, n7635, n7636, n7637, n7638,
    n7639, n7640, n7641, n7642, n7643, n7644,
    n7645, n7646, n7647, n7648, n7649, n7650,
    n7651, n7652, n7653, n7654, n7655, n7656,
    n7657, n7658, n7659, n7660, n7661, n7662,
    n7663, n7664, n7665, n7666, n7667, n7668,
    n7669, n7670, n7671, n7672, n7673, n7674,
    n7675, n7676, n7677, n7678, n7679, n7680,
    n7681, n7682, n7683, n7684, n7685, n7686,
    n7687, n7688, n7689, n7690, n7691, n7692,
    n7693, n7694, n7695, n7696, n7697, n7698,
    n7699, n7700, n7701, n7702, n7703, n7704,
    n7705, n7706, n7707, n7708, n7709, n7710,
    n7711, n7712, n7713, n7714, n7715, n7716,
    n7717, n7718, n7719, n7720, n7721, n7722,
    n7723, n7724, n7725, n7726, n7727, n7728,
    n7729, n7730, n7731, n7732, n7733, n7734,
    n7735, n7736, n7737, n7738, n7739, n7740,
    n7741, n7742, n7743, n7744, n7745, n7746,
    n7747, n7748, n7749, n7750, n7751, n7752,
    n7753, n7754, n7755, n7756, n7757, n7758,
    n7759, n7760, n7761, n7762, n7763, n7764,
    n7765, n7766, n7767, n7768, n7769, n7770,
    n7771, n7772, n7773, n7774, n7775, n7776,
    n7777, n7778, n7779, n7780, n7781, n7782,
    n7783, n7784, n7785, n7786, n7787, n7788,
    n7789, n7790, n7791, n7792, n7793, n7794,
    n7795, n7796, n7797, n7798, n7799, n7800,
    n7801, n7802, n7803, n7804, n7805, n7806,
    n7807, n7808, n7809, n7810, n7811, n7812,
    n7813, n7814, n7815, n7816, n7817, n7818,
    n7819, n7820, n7821, n7822, n7823, n7824,
    n7825, n7826, n7827, n7828, n7829, n7830,
    n7831, n7832, n7833, n7834, n7835, n7836,
    n7837, n7838, n7839, n7840, n7841, n7842,
    n7843, n7844, n7845, n7846, n7847, n7848,
    n7849, n7850, n7851, n7852, n7853, n7854,
    n7855, n7856, n7857, n7858, n7859, n7860,
    n7861, n7862, n7863, n7864, n7865, n7866,
    n7867, n7868, n7869, n7870, n7871, n7872,
    n7873, n7874, n7875, n7876, n7877, n7878,
    n7879, n7880, n7881, n7882, n7883, n7884,
    n7885, n7886, n7887, n7888, n7889, n7890,
    n7891, n7892, n7893, n7894, n7895, n7896,
    n7897, n7898, n7899, n7900, n7901, n7902,
    n7903, n7904, n7905, n7906, n7907, n7908,
    n7909, n7910, n7911, n7912, n7913, n7914,
    n7915, n7916, n7917, n7918, n7919, n7920,
    n7921, n7922, n7923, n7924, n7925, n7926,
    n7927, n7928, n7929, n7930, n7931, n7932,
    n7933, n7934, n7935, n7936, n7937, n7938,
    n7939, n7940, n7941, n7942, n7943, n7944,
    n7945, n7946, n7947, n7948, n7949, n7950,
    n7951, n7952, n7953, n7954, n7955, n7956,
    n7957, n7958, n7959, n7960, n7961, n7962,
    n7963, n7964, n7965, n7966, n7967, n7968,
    n7969, n7970, n7971, n7972, n7973, n7974,
    n7975, n7976, n7977, n7978, n7979, n7980,
    n7981, n7982, n7983, n7984, n7985, n7986,
    n7987, n7988, n7989, n7990, n7991, n7992,
    n7993, n7994, n7995, n7996, n7997, n7998,
    n7999, n8000, n8001, n8002, n8003, n8004,
    n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016,
    n8017, n8018, n8019, n8020, n8021, n8022,
    n8023, n8024, n8025, n8026, n8027, n8028,
    n8029, n8030, n8031, n8032, n8033, n8034,
    n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046,
    n8047, n8048, n8049, n8050, n8051, n8052,
    n8053, n8054, n8055, n8056, n8057, n8058,
    n8059, n8060, n8061, n8062, n8063, n8064,
    n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076,
    n8077, n8078, n8079, n8080, n8081, n8082,
    n8083, n8084, n8085, n8086, n8087, n8088,
    n8089, n8090, n8091, n8092, n8093, n8094,
    n8095, n8096, n8097, n8098, n8099, n8100,
    n8101, n8102, n8103, n8104, n8105, n8106,
    n8107, n8108, n8109, n8110, n8111, n8112,
    n8113, n8114, n8115, n8116, n8117, n8118,
    n8119, n8120, n8121, n8122, n8123, n8124,
    n8125, n8126, n8127, n8128, n8129, n8130,
    n8131, n8132, n8133, n8134, n8135, n8136,
    n8137, n8138, n8139, n8140, n8141, n8142,
    n8143, n8144, n8145, n8146, n8147, n8148,
    n8149, n8150, n8151, n8152, n8153, n8154,
    n8155, n8156, n8157, n8158, n8159, n8160,
    n8161, n8162, n8163, n8164, n8165, n8166,
    n8167, n8168, n8169, n8170, n8171, n8172,
    n8173, n8174, n8175, n8176, n8177, n8178,
    n8179, n8180, n8181, n8182, n8183, n8184,
    n8185, n8186, n8187, n8188, n8189, n8190,
    n8191, n8192, n8193, n8194, n8195, n8196,
    n8197, n8198, n8199, n8200, n8201, n8202,
    n8203, n8204, n8205, n8206, n8207, n8208,
    n8209, n8210, n8211, n8212, n8213, n8214,
    n8215, n8216, n8217, n8218, n8219, n8220,
    n8221, n8222, n8223, n8224, n8225, n8226,
    n8227, n8228, n8229, n8230, n8231, n8232,
    n8233, n8234, n8235, n8236, n8237, n8238,
    n8239, n8240, n8241, n8242, n8243, n8244,
    n8245, n8246, n8247, n8248, n8249, n8250,
    n8251, n8252, n8253, n8254, n8255, n8256,
    n8257, n8258, n8259, n8260, n8261, n8262,
    n8263, n8264, n8265, n8266, n8267, n8268,
    n8269, n8270, n8271, n8272, n8273, n8274,
    n8275, n8276, n8277, n8278, n8279, n8280,
    n8281, n8282, n8283, n8284, n8285, n8286,
    n8287, n8288, n8289, n8290, n8291, n8292,
    n8293, n8294, n8295, n8296, n8297, n8298,
    n8299, n8300, n8301, n8302, n8303, n8304,
    n8305, n8306, n8307, n8308, n8309, n8310,
    n8311, n8312, n8313, n8314, n8315, n8316,
    n8317, n8318, n8319, n8320, n8321, n8322,
    n8323, n8324, n8325, n8326, n8327, n8328,
    n8329, n8330, n8331, n8332, n8333, n8334,
    n8335, n8336, n8337, n8338, n8339, n8340,
    n8341, n8342, n8343, n8344, n8345, n8346,
    n8347, n8348, n8349, n8350, n8351, n8352,
    n8353, n8354, n8355, n8356, n8357, n8358,
    n8359, n8360, n8361, n8362, n8363, n8364,
    n8365, n8366, n8367, n8368, n8369, n8370,
    n8371, n8372, n8373, n8374, n8375, n8376,
    n8377, n8378, n8379, n8380, n8381, n8382,
    n8383, n8384, n8385, n8386, n8387, n8388,
    n8389, n8390, n8391, n8392, n8393, n8394,
    n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8403, n8404, n8405, n8406,
    n8407, n8408, n8409, n8410, n8411, n8412,
    n8413, n8414, n8415, n8416, n8417, n8418,
    n8419, n8420, n8421, n8422, n8423, n8424,
    n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8434, n8435, n8436,
    n8437, n8438, n8439, n8440, n8441, n8442,
    n8443, n8444, n8445, n8446, n8447, n8448,
    n8449, n8450, n8451, n8452, n8453, n8454,
    n8455, n8456, n8457, n8458, n8459, n8460,
    n8461, n8462, n8463, n8464, n8465, n8466,
    n8467, n8468, n8469, n8470, n8471, n8472,
    n8473, n8474, n8475, n8476, n8477, n8478,
    n8479, n8480, n8481, n8482, n8483, n8484,
    n8485, n8486, n8487, n8488, n8489, n8490,
    n8491, n8492, n8493, n8494, n8495, n8496,
    n8497, n8498, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508,
    n8509, n8510, n8511, n8512, n8513, n8514,
    n8515, n8516, n8517, n8518, n8519, n8520,
    n8521, n8522, n8523, n8524, n8525, n8526,
    n8527, n8528, n8529, n8530, n8531, n8532,
    n8533, n8534, n8535, n8536, n8537, n8538,
    n8539, n8540, n8541, n8542, n8543, n8544,
    n8545, n8546, n8547, n8548, n8549, n8550,
    n8551, n8552, n8553, n8554, n8555, n8556,
    n8557, n8558, n8559, n8560, n8561, n8562,
    n8563, n8564, n8565, n8566, n8567, n8568,
    n8569, n8570, n8571, n8572, n8573, n8574,
    n8575, n8576, n8577, n8578, n8579, n8580,
    n8581, n8582, n8583, n8584, n8585, n8586,
    n8587, n8588, n8589, n8590, n8591, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598,
    n8599, n8600, n8601, n8602, n8603, n8604,
    n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8613, n8614, n8615, n8616,
    n8617, n8618, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8631, n8632, n8633, n8634,
    n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646,
    n8647, n8648, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658,
    n8659, n8660, n8661, n8662, n8663, n8664,
    n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676,
    n8677, n8678, n8679, n8680, n8681, n8682,
    n8683, n8684, n8685, n8686, n8687, n8688,
    n8689, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706,
    n8707, n8708, n8709, n8710, n8711, n8712,
    n8713, n8714, n8715, n8716, n8717, n8718,
    n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736,
    n8737, n8738, n8739, n8740, n8741, n8742,
    n8743, n8744, n8745, n8746, n8747, n8748,
    n8749, n8750, n8751, n8752, n8753, n8754,
    n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766,
    n8767, n8768, n8769, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778,
    n8779, n8780, n8781, n8782, n8783, n8784,
    n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796,
    n8797, n8798, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808,
    n8809, n8810, n8811, n8812, n8813, n8814,
    n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826,
    n8827, n8828, n8829, n8830, n8831, n8832,
    n8833, n8834, n8835, n8836, n8837, n8838,
    n8839, n8840, n8841, n8842, n8843, n8844,
    n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856,
    n8857, n8858, n8859, n8860, n8861, n8862,
    n8863, n8864, n8865, n8866, n8867, n8868,
    n8869, n8870, n8871, n8872, n8873, n8874,
    n8875, n8876, n8877, n8878, n8879, n8880,
    n8881, n8882, n8883, n8884, n8885, n8886,
    n8887, n8888, n8889, n8890, n8891, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898,
    n8899, n8900, n8901, n8902, n8903, n8904,
    n8905, n8906, n8907, n8908, n8909, n8910,
    n8911, n8912, n8913, n8914, n8915, n8916,
    n8917, n8918, n8919, n8920, n8921, n8922,
    n8923, n8924, n8925, n8926, n8927, n8928,
    n8929, n8930, n8931, n8932, n8933, n8934,
    n8935, n8936, n8937, n8938, n8939, n8940,
    n8941, n8942, n8943, n8944, n8945, n8946,
    n8947, n8948, n8949, n8950, n8951, n8952,
    n8953, n8954, n8955, n8956, n8957, n8958,
    n8959, n8960, n8961, n8962, n8963, n8964,
    n8965, n8966, n8967, n8968, n8969, n8970,
    n8971, n8972, n8973, n8974, n8975, n8976,
    n8977, n8978, n8979, n8980, n8981, n8982,
    n8983, n8984, n8985, n8986, n8987, n8988,
    n8989, n8990, n8991, n8992, n8993, n8994,
    n8995, n8996, n8997, n8998, n8999, n9000,
    n9001, n9002, n9003, n9004, n9005, n9006,
    n9007, n9008, n9009, n9010, n9011, n9012,
    n9013, n9014, n9015, n9016, n9017, n9018,
    n9019, n9020, n9021, n9022, n9023, n9024,
    n9025, n9026, n9027, n9028, n9029, n9030,
    n9031, n9032, n9033, n9034, n9035, n9036,
    n9037, n9038, n9039, n9040, n9041, n9042,
    n9043, n9044, n9045, n9046, n9047, n9048,
    n9049, n9050, n9051, n9052, n9053, n9054,
    n9055, n9056, n9057, n9058, n9059, n9060,
    n9061, n9062, n9063, n9064, n9065, n9066,
    n9067, n9068, n9069, n9070, n9071, n9072,
    n9073, n9074, n9075, n9076, n9077, n9078,
    n9079, n9080, n9081, n9082, n9083, n9084,
    n9085, n9086, n9087, n9088, n9089, n9090,
    n9091, n9092, n9093, n9094, n9095, n9096,
    n9097, n9098, n9099, n9100, n9101, n9102,
    n9103, n9104, n9105, n9106, n9107, n9108,
    n9109, n9110, n9111, n9112, n9113, n9114,
    n9115, n9116, n9117, n9118, n9119, n9120,
    n9121, n9122, n9123, n9124, n9125, n9126,
    n9127, n9128, n9129, n9130, n9131, n9132,
    n9133, n9134, n9135, n9136, n9137, n9138,
    n9139, n9140, n9141, n9142, n9143, n9144,
    n9145, n9146, n9147, n9148, n9149, n9150,
    n9151, n9152, n9153, n9154, n9155, n9156,
    n9157, n9158, n9159, n9160, n9161, n9162,
    n9163, n9164, n9165, n9166, n9167, n9168,
    n9169, n9170, n9171, n9172, n9173, n9174,
    n9175, n9176, n9177, n9178, n9179, n9180,
    n9181, n9182, n9183, n9184, n9185, n9186,
    n9187, n9188, n9189, n9190, n9191, n9192,
    n9193, n9194, n9195, n9196, n9197, n9198,
    n9199, n9200, n9201, n9202, n9203, n9204,
    n9205, n9206, n9207, n9208, n9209, n9210,
    n9211, n9212, n9213, n9214, n9215, n9216,
    n9217, n9218, n9219, n9220, n9221, n9222,
    n9223, n9224, n9225, n9226, n9227, n9228,
    n9229, n9230, n9231, n9232, n9233, n9234,
    n9235, n9236, n9237, n9238, n9239, n9240,
    n9241, n9242, n9243, n9244, n9245, n9246,
    n9247, n9248, n9249, n9250, n9251, n9252,
    n9253, n9254, n9255, n9256, n9257, n9258,
    n9259, n9260, n9261, n9262, n9263, n9264,
    n9265, n9266, n9267, n9268, n9269, n9270,
    n9271, n9272, n9273, n9274, n9275, n9276,
    n9277, n9278, n9279, n9280, n9281, n9282,
    n9283, n9284, n9285, n9286, n9287, n9288,
    n9289, n9290, n9291, n9292, n9293, n9294,
    n9295, n9296, n9297, n9298, n9299, n9300,
    n9301, n9302, n9303, n9304, n9305, n9306,
    n9307, n9308, n9309, n9310, n9311, n9312,
    n9313, n9314, n9315, n9316, n9317, n9318,
    n9319, n9320, n9321, n9322, n9323, n9324,
    n9325, n9326, n9327, n9328, n9329, n9330,
    n9331, n9332, n9333, n9334, n9335, n9336,
    n9337, n9338, n9339, n9340, n9341, n9342,
    n9343, n9344, n9345, n9346, n9347, n9348,
    n9349, n9350, n9351, n9352, n9353, n9354,
    n9355, n9356, n9357, n9358, n9359, n9360,
    n9361, n9362, n9363, n9364, n9365, n9366,
    n9367, n9368, n9369, n9370, n9371, n9372,
    n9373, n9374, n9375, n9376, n9377, n9378,
    n9379, n9380, n9381, n9382, n9383, n9384,
    n9385, n9386, n9387, n9388, n9389, n9390,
    n9391, n9392, n9393, n9394, n9395, n9396,
    n9397, n9398, n9399, n9400, n9401, n9402,
    n9403, n9404, n9405, n9406, n9407, n9408,
    n9409, n9410, n9411, n9412, n9413, n9414,
    n9415, n9416, n9417, n9418, n9419, n9420,
    n9421, n9422, n9423, n9424, n9425, n9426,
    n9427, n9428, n9429, n9430, n9431, n9432,
    n9433, n9434, n9435, n9436, n9437, n9438,
    n9439, n9440, n9441, n9442, n9443, n9444,
    n9445, n9446, n9447, n9448, n9449, n9450,
    n9451, n9452, n9453, n9454, n9455, n9456,
    n9457, n9458, n9459, n9460, n9461, n9462,
    n9463, n9464, n9465, n9466, n9467, n9468,
    n9469, n9470, n9471, n9472, n9473, n9474,
    n9475, n9476, n9477, n9478, n9479, n9480,
    n9481, n9482, n9483, n9484, n9485, n9486,
    n9487, n9488, n9489, n9490, n9491, n9492,
    n9493, n9494, n9495, n9496, n9497, n9498,
    n9499, n9500, n9501, n9502, n9503, n9504,
    n9505, n9506, n9507, n9508, n9509, n9510,
    n9511, n9512, n9513, n9514, n9515, n9516,
    n9517, n9518, n9519, n9520, n9521, n9522,
    n9523, n9524, n9525, n9526, n9527, n9528,
    n9529, n9530, n9531, n9532, n9533, n9534,
    n9535, n9536, n9537, n9538, n9539, n9540,
    n9541, n9542, n9543, n9544, n9545, n9546,
    n9547, n9548, n9549, n9550, n9551, n9552,
    n9553, n9554, n9555, n9556, n9557, n9558,
    n9559, n9560, n9561, n9562, n9563, n9564,
    n9565, n9566, n9567, n9568, n9569, n9570,
    n9571, n9572, n9573, n9574, n9575, n9576,
    n9577, n9578, n9579, n9580, n9581, n9582,
    n9583, n9584, n9585, n9586, n9587, n9588,
    n9589, n9590, n9591, n9592, n9593, n9594,
    n9595, n9596, n9597, n9598, n9599, n9600,
    n9601, n9602, n9603, n9604, n9605, n9606,
    n9607, n9608, n9609, n9610, n9611, n9612,
    n9613, n9614, n9615, n9616, n9617, n9618,
    n9619, n9620, n9621, n9622, n9623, n9624,
    n9625, n9626, n9627, n9628, n9629, n9630,
    n9631, n9632, n9633, n9634, n9635, n9636,
    n9637, n9638, n9639, n9640, n9641, n9642,
    n9643, n9644, n9645, n9646, n9647, n9648,
    n9649, n9650, n9651, n9652, n9653, n9654,
    n9655, n9656, n9657, n9658, n9659, n9660,
    n9661, n9662, n9663, n9664, n9665, n9666,
    n9667, n9668, n9669, n9670, n9671, n9672,
    n9673, n9674, n9675, n9676, n9677, n9678,
    n9679, n9680, n9681, n9682, n9683, n9684,
    n9685, n9686, n9687, n9688, n9689, n9690,
    n9691, n9692, n9693, n9694, n9695, n9696,
    n9697, n9698, n9699, n9700, n9701, n9702,
    n9703, n9704, n9705, n9706, n9707, n9708,
    n9709, n9710, n9711, n9712, n9713, n9714,
    n9715, n9716, n9717, n9718, n9719, n9720,
    n9721, n9722, n9723, n9724, n9725, n9726,
    n9727, n9728, n9729, n9730, n9731, n9732,
    n9733, n9734, n9735, n9736, n9737, n9738,
    n9739, n9740, n9741, n9742, n9743, n9744,
    n9745, n9746, n9747, n9748, n9749, n9750,
    n9751, n9752, n9753, n9754, n9755, n9756,
    n9757, n9758, n9759, n9760, n9761, n9762,
    n9763, n9764, n9765, n9766, n9767, n9768,
    n9769, n9770, n9771, n9772, n9773, n9774,
    n9775, n9776, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786,
    n9787, n9788, n9789, n9790, n9791, n9792,
    n9793, n9794, n9795, n9796, n9797, n9798,
    n9799, n9800, n9801, n9802, n9803, n9804,
    n9805, n9806, n9807, n9808, n9809, n9810,
    n9811, n9812, n9813, n9814, n9815, n9816,
    n9817, n9818, n9819, n9820, n9821, n9822,
    n9823, n9824, n9825, n9826, n9827, n9828,
    n9829, n9830, n9831, n9832, n9833, n9834,
    n9835, n9836, n9837, n9838, n9839, n9840,
    n9841, n9842, n9843, n9844, n9845, n9846,
    n9847, n9848, n9849, n9850, n9851, n9852,
    n9853, n9854, n9855, n9856, n9857, n9858,
    n9859, n9860, n9861, n9862, n9863, n9864,
    n9865, n9866, n9867, n9868, n9869, n9870,
    n9871, n9872, n9873, n9874, n9875, n9876,
    n9877, n9878, n9879, n9880, n9881, n9882,
    n9883, n9884, n9885, n9886, n9887, n9888,
    n9889, n9890, n9891, n9892, n9893, n9894,
    n9895, n9896, n9897, n9898, n9899, n9900,
    n9901, n9902, n9903, n9904, n9905, n9906,
    n9907, n9908, n9909, n9910, n9911, n9912,
    n9913, n9914, n9915, n9916, n9917, n9918,
    n9919, n9920, n9921, n9922, n9923, n9924,
    n9925, n9926, n9927, n9928, n9929, n9930,
    n9931, n9932, n9933, n9934, n9935, n9936,
    n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948,
    n9949, n9950, n9951, n9952, n9953, n9954,
    n9955, n9956, n9957, n9958, n9959, n9960,
    n9961, n9962, n9963, n9964, n9965, n9966,
    n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9990,
    n9991, n9992, n9993, n9994, n9995, n9996,
    n9997, n9998, n9999, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026,
    n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044,
    n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062,
    n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074,
    n10075, n10076, n10077, n10078, n10079, n10080,
    n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092,
    n10093, n10094, n10095, n10096, n10097, n10098,
    n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116,
    n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134,
    n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146,
    n10147, n10148, n10149, n10150, n10151, n10152,
    n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170,
    n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188,
    n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200,
    n10201, n10202, n10203, n10204, n10205, n10206,
    n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218,
    n10219, n10220, n10221, n10222, n10223, n10224,
    n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236,
    n10237, n10238, n10239, n10240, n10241, n10242,
    n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254,
    n10255, n10256, n10257, n10258, n10259, n10260,
    n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272,
    n10273, n10274, n10275, n10276, n10277, n10278,
    n10279, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290,
    n10291, n10292, n10293, n10294, n10295, n10296,
    n10297, n10298, n10299, n10300, n10301, n10302,
    n10303, n10304, n10305, n10306, n10307, n10308,
    n10309, n10310, n10311, n10312, n10313, n10314,
    n10315, n10316, n10317, n10318, n10319, n10320,
    n10321, n10322, n10323, n10324, n10325, n10326,
    n10327, n10328, n10329, n10330, n10331, n10332,
    n10333, n10334, n10335, n10336, n10337, n10338,
    n10339, n10340, n10341, n10342, n10343, n10344,
    n10345, n10346, n10347, n10348, n10349, n10350,
    n10351, n10352, n10353, n10354, n10355, n10356,
    n10357, n10358, n10359, n10360, n10361, n10362,
    n10363, n10364, n10365, n10366, n10367, n10368,
    n10369, n10370, n10371, n10372, n10373, n10374,
    n10375, n10376, n10377, n10378, n10379, n10380,
    n10381, n10382, n10383, n10384, n10385, n10386,
    n10387, n10388, n10389, n10390, n10391, n10392,
    n10393, n10394, n10395, n10396, n10397, n10398,
    n10399, n10400, n10401, n10402, n10403, n10404,
    n10405, n10406, n10407, n10408, n10409, n10410,
    n10411, n10412, n10413, n10414, n10415, n10416,
    n10417, n10418, n10419, n10420, n10421, n10422,
    n10423, n10424, n10425, n10426, n10427, n10428,
    n10429, n10430, n10431, n10432, n10433, n10434,
    n10435, n10436, n10437, n10438, n10439, n10440,
    n10441, n10442, n10443, n10444, n10445, n10446,
    n10447, n10448, n10449, n10450, n10451, n10452,
    n10453, n10454, n10455, n10456, n10457, n10458,
    n10459, n10460, n10461, n10462, n10463, n10464,
    n10465, n10466, n10467, n10468, n10469, n10470,
    n10471, n10472, n10473, n10474, n10475, n10476,
    n10477, n10478, n10479, n10480, n10481, n10482,
    n10483, n10484, n10485, n10486, n10487, n10488,
    n10489, n10490, n10491, n10492, n10493, n10494,
    n10495, n10496, n10497, n10498, n10499, n10500,
    n10501, n10502, n10503, n10504, n10505, n10506,
    n10507, n10508, n10509, n10510, n10511, n10512,
    n10513, n10514, n10515, n10516, n10517, n10518,
    n10519, n10520, n10521, n10522, n10523, n10524,
    n10525, n10526, n10527, n10528, n10529, n10530,
    n10531, n10532, n10533, n10534, n10535, n10536,
    n10537, n10538, n10539, n10540, n10541, n10542,
    n10543, n10544, n10545, n10546, n10547, n10548,
    n10549, n10550, n10551, n10552, n10553, n10554,
    n10555, n10556, n10557, n10558, n10559, n10560,
    n10561, n10562, n10563, n10564, n10565, n10566,
    n10567, n10568, n10569, n10570, n10571, n10572,
    n10573, n10574, n10575, n10576, n10577, n10578,
    n10579, n10580, n10581, n10582, n10583, n10584,
    n10585, n10586, n10587, n10588, n10589, n10590,
    n10591, n10592, n10593, n10594, n10595, n10596,
    n10597, n10598, n10599, n10600, n10601, n10602,
    n10603, n10604, n10605, n10606, n10607, n10608,
    n10609, n10610, n10611, n10612, n10613, n10614,
    n10615, n10616, n10617, n10618, n10619, n10620,
    n10621, n10622, n10623, n10624, n10625, n10626,
    n10627, n10628, n10629, n10630, n10631, n10632,
    n10633, n10634, n10635, n10636, n10637, n10638,
    n10639, n10640, n10641, n10642, n10643, n10644,
    n10645, n10646, n10647, n10648, n10649, n10650,
    n10651, n10652, n10653, n10654, n10655, n10656,
    n10657, n10658, n10659, n10660, n10661, n10662,
    n10663, n10664, n10665, n10666, n10667, n10668,
    n10669, n10670, n10671, n10672, n10673, n10674,
    n10675, n10676, n10677, n10678, n10679, n10680,
    n10681, n10682, n10683, n10684, n10685, n10686,
    n10687, n10688, n10689, n10690, n10691, n10692,
    n10693, n10694, n10695, n10696, n10697, n10698,
    n10699, n10700, n10701, n10702, n10703, n10704,
    n10705, n10706, n10707, n10708, n10709, n10710,
    n10711, n10712, n10713, n10714, n10715, n10716,
    n10717, n10718, n10719, n10720, n10721, n10722,
    n10723, n10724, n10725, n10726, n10727, n10728,
    n10729, n10730, n10731, n10732, n10733, n10734,
    n10735, n10736, n10737, n10738, n10739, n10740,
    n10741, n10742, n10743, n10744, n10745, n10746,
    n10747, n10748, n10749, n10750, n10751, n10752,
    n10753, n10754, n10755, n10756, n10757, n10758,
    n10759, n10760, n10761, n10762, n10763, n10764,
    n10765, n10766, n10767, n10768, n10769, n10770,
    n10771, n10772, n10773, n10774, n10775, n10776,
    n10777, n10778, n10779, n10780, n10781, n10782,
    n10783, n10784, n10785, n10786, n10787, n10788,
    n10789, n10790, n10791, n10792, n10793, n10794,
    n10795, n10796, n10797, n10798, n10799, n10800,
    n10801, n10802, n10803, n10804, n10805, n10806,
    n10807, n10808, n10809, n10810, n10811, n10812,
    n10813, n10814, n10815, n10816, n10817, n10818,
    n10819, n10820, n10821, n10822, n10823, n10824,
    n10825, n10826, n10827, n10828, n10829, n10830,
    n10831, n10832, n10833, n10834, n10835, n10836,
    n10837, n10838, n10839, n10840, n10841, n10842,
    n10843, n10844, n10845, n10846, n10847, n10848,
    n10849, n10850, n10851, n10852, n10853, n10854,
    n10855, n10856, n10857, n10858, n10859, n10860,
    n10861, n10862, n10863, n10864, n10865, n10866,
    n10867, n10868, n10869, n10870, n10871, n10872,
    n10873, n10874, n10875, n10876, n10877, n10878,
    n10879, n10880, n10881, n10882, n10883, n10884,
    n10885, n10886, n10887, n10888, n10889, n10890,
    n10891, n10892, n10893, n10894, n10895, n10896,
    n10897, n10898, n10899, n10900, n10901, n10902,
    n10903, n10904, n10905, n10906, n10907, n10908,
    n10909, n10910, n10911, n10912, n10913, n10914,
    n10915, n10916, n10917, n10918, n10919, n10920,
    n10921, n10922, n10923, n10924, n10925, n10926,
    n10927, n10928, n10929, n10930, n10931, n10932,
    n10933, n10934, n10935, n10936, n10937, n10938,
    n10939, n10940, n10941, n10942, n10943, n10944,
    n10945, n10946, n10947, n10948, n10949, n10950,
    n10951, n10952, n10953, n10954, n10955, n10956,
    n10957, n10958, n10959, n10960, n10961, n10962,
    n10963, n10964, n10965, n10966, n10967, n10968,
    n10969, n10970, n10971, n10972, n10973, n10974,
    n10975, n10976, n10977, n10978, n10979, n10980,
    n10981, n10982, n10983, n10984, n10985, n10986,
    n10987, n10988, n10989, n10990, n10991, n10992,
    n10993, n10994, n10995, n10996, n10997, n10998,
    n10999, n11000, n11001, n11002, n11003, n11004,
    n11005, n11006, n11007, n11008, n11009, n11010,
    n11011, n11012, n11013, n11014, n11015, n11016,
    n11017, n11018, n11019, n11020, n11021, n11022,
    n11023, n11024, n11025, n11026, n11027, n11028,
    n11029, n11030, n11031, n11032, n11033, n11034,
    n11035, n11036, n11037, n11038, n11039, n11040,
    n11041, n11042, n11043, n11044, n11045, n11046,
    n11047, n11048, n11049, n11050, n11051, n11052,
    n11053, n11054, n11055, n11056, n11057, n11058,
    n11059, n11060, n11061, n11062, n11063, n11064,
    n11065, n11066, n11067, n11068, n11069, n11070,
    n11071, n11072, n11073, n11074, n11075, n11076,
    n11077, n11078, n11079, n11080, n11081, n11082,
    n11083, n11084, n11085, n11086, n11087, n11088,
    n11089, n11090, n11091, n11092, n11093, n11094,
    n11095, n11096, n11097, n11098, n11099, n11100,
    n11101, n11102, n11103, n11104, n11105, n11106,
    n11107, n11108, n11109, n11110, n11111, n11112,
    n11113, n11114, n11115, n11116, n11117, n11118,
    n11119, n11120, n11121, n11122, n11123, n11124,
    n11125, n11126, n11127, n11128, n11129, n11130,
    n11131, n11132, n11133, n11134, n11135, n11136,
    n11137, n11138, n11139, n11140, n11141, n11142,
    n11143, n11144, n11145, n11146, n11147, n11148,
    n11149, n11150, n11151, n11152, n11153, n11154,
    n11155, n11156;
  assign n1003 = pi67  & ~pi68 ;
  assign n1004 = ~pi67  & pi68 ;
  assign n1005 = ~n1003 & ~n1004;
  assign n1006 = ~pi69  & ~n1005;
  assign n1007 = pi69  & n1005;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = pi70  & ~pi71 ;
  assign n1010 = ~pi70  & pi71 ;
  assign n1011 = ~n1009 & ~n1010;
  assign n1012 = ~pi72  & ~n1011;
  assign n1013 = pi72  & n1011;
  assign n1014 = ~n1012 & ~n1013;
  assign n1015 = ~n1008 & ~n1014;
  assign n1016 = pi70  & pi71 ;
  assign n1017 = pi72  & ~n1011;
  assign n1018 = ~n1016 & ~n1017;
  assign n1019 = pi67  & pi68 ;
  assign n1020 = pi69  & ~n1005;
  assign n1021 = ~n1019 & ~n1020;
  assign n1022 = n1018 & ~n1021;
  assign n1023 = ~n1018 & n1021;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = n1015 & ~n1024;
  assign n1026 = ~n1018 & ~n1021;
  assign n1027 = ~n1025 & ~n1026;
  assign n1028 = pi76  & pi77 ;
  assign n1029 = pi76  & ~pi77 ;
  assign n1030 = ~pi76  & pi77 ;
  assign n1031 = ~n1029 & ~n1030;
  assign n1032 = pi78  & ~n1031;
  assign n1033 = ~n1028 & ~n1032;
  assign n1034 = pi73  & pi74 ;
  assign n1035 = pi73  & ~pi74 ;
  assign n1036 = ~pi73  & pi74 ;
  assign n1037 = ~n1035 & ~n1036;
  assign n1038 = pi75  & ~n1037;
  assign n1039 = ~n1034 & ~n1038;
  assign n1040 = ~n1033 & n1039;
  assign n1041 = n1033 & ~n1039;
  assign n1042 = ~n1040 & ~n1041;
  assign n1043 = ~pi75  & ~n1037;
  assign n1044 = pi75  & n1037;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = ~pi78  & ~n1031;
  assign n1047 = pi78  & n1031;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = ~n1045 & ~n1048;
  assign n1050 = ~n1042 & n1049;
  assign n1051 = ~n1033 & ~n1039;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = n1015 & n1024;
  assign n1054 = ~n1015 & ~n1024;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = n1042 & n1049;
  assign n1057 = ~n1042 & ~n1049;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = ~n1052 & ~n1058;
  assign n1060 = ~n1027 & ~n1055;
  assign n1061 = ~n1008 & n1014;
  assign n1062 = n1008 & ~n1014;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = ~n1045 & n1048;
  assign n1065 = n1045 & ~n1048;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = ~n1063 & ~n1066;
  assign n1068 = ~n1059 & n1067;
  assign n1069 = ~n1060 & n1068;
  assign n1070 = n1058 & ~n1069;
  assign n1071 = ~n1055 & ~n1070;
  assign n1072 = n1058 & n1069;
  assign n1073 = n1069 & ~n1072;
  assign n1074 = ~n1071 & ~n1073;
  assign n1075 = n1052 & n1074;
  assign n1076 = ~n1027 & ~n1075;
  assign n1077 = ~n1052 & ~n1074;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = pi55  & ~pi56 ;
  assign n1080 = ~pi55  & pi56 ;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = ~pi57  & ~n1081;
  assign n1083 = pi57  & n1081;
  assign n1084 = ~n1082 & ~n1083;
  assign n1085 = pi58  & ~pi59 ;
  assign n1086 = ~pi58  & pi59 ;
  assign n1087 = ~n1085 & ~n1086;
  assign n1088 = ~pi60  & ~n1087;
  assign n1089 = pi60  & n1087;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = ~n1084 & ~n1090;
  assign n1092 = pi58  & pi59 ;
  assign n1093 = pi60  & ~n1087;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = pi55  & pi56 ;
  assign n1096 = pi57  & ~n1081;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = n1094 & ~n1097;
  assign n1099 = ~n1094 & n1097;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = n1091 & ~n1100;
  assign n1102 = ~n1094 & ~n1097;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = pi64  & pi65 ;
  assign n1105 = pi64  & ~pi65 ;
  assign n1106 = ~pi64  & pi65 ;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = pi66  & ~n1107;
  assign n1109 = ~n1104 & ~n1108;
  assign n1110 = pi61  & pi62 ;
  assign n1111 = pi61  & ~pi62 ;
  assign n1112 = ~pi61  & pi62 ;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = pi63  & ~n1113;
  assign n1115 = ~n1110 & ~n1114;
  assign n1116 = ~n1109 & n1115;
  assign n1117 = n1109 & ~n1115;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = ~pi63  & ~n1113;
  assign n1120 = pi63  & n1113;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122 = ~pi66  & ~n1107;
  assign n1123 = pi66  & n1107;
  assign n1124 = ~n1122 & ~n1123;
  assign n1125 = ~n1121 & ~n1124;
  assign n1126 = ~n1118 & n1125;
  assign n1127 = ~n1109 & ~n1115;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = n1091 & n1100;
  assign n1130 = ~n1091 & ~n1100;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = n1118 & n1125;
  assign n1133 = ~n1118 & ~n1125;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = ~n1128 & ~n1134;
  assign n1136 = ~n1103 & ~n1131;
  assign n1137 = ~n1084 & n1090;
  assign n1138 = n1084 & ~n1090;
  assign n1139 = ~n1137 & ~n1138;
  assign n1140 = ~n1121 & n1124;
  assign n1141 = n1121 & ~n1124;
  assign n1142 = ~n1140 & ~n1141;
  assign n1143 = ~n1139 & ~n1142;
  assign n1144 = ~n1135 & n1143;
  assign n1145 = ~n1136 & n1144;
  assign n1146 = n1134 & ~n1145;
  assign n1147 = ~n1131 & ~n1146;
  assign n1148 = ~n1134 & n1145;
  assign n1149 = ~n1147 & ~n1148;
  assign n1150 = n1128 & n1149;
  assign n1151 = ~n1103 & ~n1150;
  assign n1152 = ~n1128 & ~n1149;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = n1078 & n1153;
  assign n1155 = ~n1103 & n1128;
  assign n1156 = n1103 & ~n1128;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~n1149 & ~n1157;
  assign n1159 = n1149 & n1157;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = ~n1027 & n1052;
  assign n1162 = n1027 & ~n1052;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = ~n1074 & ~n1163;
  assign n1165 = n1074 & n1163;
  assign n1166 = ~n1164 & ~n1165;
  assign n1167 = n1160 & n1166;
  assign n1168 = ~n1063 & n1066;
  assign n1169 = n1063 & ~n1066;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = ~n1139 & n1142;
  assign n1172 = n1139 & ~n1142;
  assign n1173 = ~n1171 & ~n1172;
  assign n1174 = ~n1170 & ~n1173;
  assign n1175 = ~n1058 & ~n1069;
  assign n1176 = ~n1072 & ~n1175;
  assign n1177 = ~n1055 & n1176;
  assign n1178 = n1055 & ~n1176;
  assign n1179 = ~n1177 & ~n1178;
  assign n1180 = n1174 & ~n1179;
  assign n1181 = ~n1146 & ~n1148;
  assign n1182 = n1131 & n1181;
  assign n1183 = ~n1131 & ~n1181;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = ~n1174 & n1179;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = ~n1180 & ~n1186;
  assign n1188 = ~n1160 & ~n1166;
  assign n1189 = ~n1167 & ~n1188;
  assign n1190 = ~n1187 & n1189;
  assign n1191 = ~n1167 & ~n1190;
  assign n1192 = ~n1154 & ~n1191;
  assign n1193 = ~n1078 & ~n1153;
  assign n1194 = ~n1192 & ~n1193;
  assign n1195 = pi43  & ~pi44 ;
  assign n1196 = ~pi43  & pi44 ;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = ~pi45  & ~n1197;
  assign n1199 = pi45  & n1197;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = pi46  & ~pi47 ;
  assign n1202 = ~pi46  & pi47 ;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = ~pi48  & ~n1203;
  assign n1205 = pi48  & n1203;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = ~n1200 & n1206;
  assign n1208 = n1200 & ~n1206;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = pi49  & ~pi50 ;
  assign n1211 = ~pi49  & pi50 ;
  assign n1212 = ~n1210 & ~n1211;
  assign n1213 = ~pi51  & ~n1212;
  assign n1214 = pi51  & n1212;
  assign n1215 = ~n1213 & ~n1214;
  assign n1216 = pi52  & ~pi53 ;
  assign n1217 = ~pi52  & pi53 ;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = ~pi54  & ~n1218;
  assign n1220 = pi54  & n1218;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = ~n1215 & n1221;
  assign n1223 = n1215 & ~n1221;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = ~n1209 & n1224;
  assign n1226 = n1209 & ~n1224;
  assign n1227 = ~n1225 & ~n1226;
  assign n1228 = ~pi37  & pi38 ;
  assign n1229 = pi37  & ~pi38 ;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = ~pi39  & ~n1230;
  assign n1232 = pi39  & n1230;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = ~pi40  & pi41 ;
  assign n1235 = pi40  & ~pi41 ;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = ~pi42  & ~n1236;
  assign n1238 = pi42  & n1236;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = ~n1233 & n1239;
  assign n1241 = n1233 & ~n1239;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = ~pi31  & pi32 ;
  assign n1244 = pi31  & ~pi32 ;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = ~pi33  & ~n1245;
  assign n1247 = pi33  & n1245;
  assign n1248 = ~n1246 & ~n1247;
  assign n1249 = ~pi34  & pi35 ;
  assign n1250 = pi34  & ~pi35 ;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = ~pi36  & ~n1251;
  assign n1253 = pi36  & n1251;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = ~n1248 & n1254;
  assign n1256 = n1248 & ~n1254;
  assign n1257 = ~n1255 & ~n1256;
  assign n1258 = n1242 & ~n1257;
  assign n1259 = ~n1242 & n1257;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = ~n1227 & ~n1260;
  assign n1262 = ~n1200 & ~n1206;
  assign n1263 = pi46  & pi47 ;
  assign n1264 = pi48  & ~n1203;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = pi43  & pi44 ;
  assign n1267 = pi45  & ~n1197;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = n1265 & ~n1268;
  assign n1270 = ~n1265 & n1268;
  assign n1271 = ~n1269 & ~n1270;
  assign n1272 = n1262 & n1271;
  assign n1273 = ~n1262 & ~n1271;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = pi52  & pi53 ;
  assign n1276 = pi54  & ~n1218;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = pi49  & pi50 ;
  assign n1279 = pi51  & ~n1212;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = ~n1277 & n1280;
  assign n1282 = n1277 & ~n1280;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = ~n1215 & ~n1221;
  assign n1285 = n1283 & n1284;
  assign n1286 = ~n1283 & ~n1284;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = ~n1283 & n1284;
  assign n1289 = ~n1277 & ~n1280;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = ~n1287 & ~n1290;
  assign n1292 = n1262 & ~n1271;
  assign n1293 = ~n1265 & ~n1268;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = ~n1274 & ~n1294;
  assign n1296 = ~n1209 & ~n1224;
  assign n1297 = ~n1291 & n1296;
  assign n1298 = ~n1295 & n1297;
  assign n1299 = ~n1287 & ~n1298;
  assign n1300 = n1287 & n1298;
  assign n1301 = ~n1299 & ~n1300;
  assign n1302 = ~n1274 & n1301;
  assign n1303 = n1274 & ~n1301;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = n1261 & ~n1304;
  assign n1306 = pi34  & pi35 ;
  assign n1307 = pi36  & ~n1251;
  assign n1308 = ~n1306 & ~n1307;
  assign n1309 = pi31  & pi32 ;
  assign n1310 = pi33  & ~n1245;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = ~n1308 & n1311;
  assign n1313 = n1308 & ~n1311;
  assign n1314 = ~n1312 & ~n1313;
  assign n1315 = ~n1248 & ~n1254;
  assign n1316 = n1314 & n1315;
  assign n1317 = ~n1314 & ~n1315;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = pi40  & pi41 ;
  assign n1320 = pi42  & ~n1236;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = pi37  & pi38 ;
  assign n1323 = pi39  & ~n1230;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = ~n1321 & n1324;
  assign n1326 = n1321 & ~n1324;
  assign n1327 = ~n1325 & ~n1326;
  assign n1328 = ~n1233 & ~n1239;
  assign n1329 = n1327 & n1328;
  assign n1330 = ~n1327 & ~n1328;
  assign n1331 = ~n1329 & ~n1330;
  assign n1332 = ~n1327 & n1328;
  assign n1333 = ~n1321 & ~n1324;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = ~n1331 & ~n1334;
  assign n1336 = ~n1314 & n1315;
  assign n1337 = ~n1308 & ~n1311;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = ~n1318 & ~n1338;
  assign n1340 = ~n1242 & ~n1257;
  assign n1341 = ~n1335 & n1340;
  assign n1342 = ~n1339 & n1341;
  assign n1343 = n1331 & ~n1342;
  assign n1344 = ~n1331 & n1342;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = n1318 & n1345;
  assign n1347 = ~n1318 & ~n1345;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = ~n1261 & n1304;
  assign n1350 = ~n1348 & ~n1349;
  assign n1351 = ~n1305 & ~n1350;
  assign n1352 = ~n1318 & ~n1343;
  assign n1353 = ~n1344 & ~n1352;
  assign n1354 = n1334 & ~n1338;
  assign n1355 = ~n1334 & n1338;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = ~n1353 & ~n1356;
  assign n1358 = n1353 & n1356;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = n1287 & ~n1298;
  assign n1361 = ~n1274 & ~n1360;
  assign n1362 = n1298 & ~n1300;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = n1290 & ~n1294;
  assign n1365 = ~n1290 & n1294;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~n1363 & ~n1366;
  assign n1368 = n1363 & n1366;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = ~n1359 & ~n1369;
  assign n1371 = ~n1351 & ~n1370;
  assign n1372 = n1359 & n1369;
  assign n1373 = ~n1371 & ~n1372;
  assign n1374 = n1290 & n1363;
  assign n1375 = ~n1294 & ~n1374;
  assign n1376 = ~n1290 & ~n1363;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = n1334 & n1353;
  assign n1379 = ~n1338 & ~n1378;
  assign n1380 = ~n1334 & ~n1353;
  assign n1381 = ~n1379 & ~n1380;
  assign n1382 = n1377 & n1381;
  assign n1383 = ~n1373 & ~n1382;
  assign n1384 = ~n1377 & ~n1381;
  assign n1385 = ~n1383 & ~n1384;
  assign n1386 = ~n1194 & ~n1385;
  assign n1387 = ~n1154 & ~n1193;
  assign n1388 = ~n1191 & n1387;
  assign n1389 = n1191 & ~n1387;
  assign n1390 = ~n1388 & ~n1389;
  assign n1391 = n1377 & ~n1381;
  assign n1392 = ~n1377 & n1381;
  assign n1393 = ~n1372 & ~n1391;
  assign n1394 = ~n1392 & n1393;
  assign n1395 = ~n1371 & n1394;
  assign n1396 = n1383 & ~n1384;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = n1390 & n1397;
  assign n1399 = ~n1170 & n1173;
  assign n1400 = n1170 & ~n1173;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = ~n1227 & n1260;
  assign n1403 = n1227 & ~n1260;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = ~n1401 & ~n1404;
  assign n1406 = ~n1180 & ~n1185;
  assign n1407 = ~n1184 & ~n1406;
  assign n1408 = n1184 & n1406;
  assign n1409 = ~n1407 & ~n1408;
  assign n1410 = n1405 & ~n1409;
  assign n1411 = ~n1305 & ~n1349;
  assign n1412 = n1348 & n1411;
  assign n1413 = ~n1348 & ~n1411;
  assign n1414 = ~n1412 & ~n1413;
  assign n1415 = ~n1405 & n1409;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = ~n1410 & ~n1416;
  assign n1418 = ~n1370 & ~n1372;
  assign n1419 = ~n1351 & n1418;
  assign n1420 = n1351 & ~n1418;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = n1187 & ~n1189;
  assign n1423 = ~n1190 & ~n1422;
  assign n1424 = ~n1421 & ~n1423;
  assign n1425 = ~n1417 & ~n1424;
  assign n1426 = n1421 & n1423;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = ~n1390 & ~n1397;
  assign n1429 = ~n1427 & ~n1428;
  assign n1430 = ~n1398 & ~n1429;
  assign n1431 = n1194 & n1385;
  assign n1432 = ~n1386 & ~n1431;
  assign n1433 = ~n1430 & n1432;
  assign n1434 = ~n1386 & ~n1433;
  assign n1435 = pi994  & pi995 ;
  assign n1436 = ~pi994  & pi995 ;
  assign n1437 = pi994  & ~pi995 ;
  assign n1438 = ~n1436 & ~n1437;
  assign n1439 = pi996  & ~n1438;
  assign n1440 = ~n1435 & ~n1439;
  assign n1441 = pi991  & pi992 ;
  assign n1442 = ~pi991  & pi992 ;
  assign n1443 = pi991  & ~pi992 ;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = pi993  & ~n1444;
  assign n1446 = ~n1441 & ~n1445;
  assign n1447 = ~n1440 & n1446;
  assign n1448 = n1440 & ~n1446;
  assign n1449 = ~n1447 & ~n1448;
  assign n1450 = ~pi993  & ~n1444;
  assign n1451 = pi993  & n1444;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = ~pi996  & ~n1438;
  assign n1454 = pi996  & n1438;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = ~n1452 & ~n1455;
  assign n1457 = ~n1449 & n1456;
  assign n1458 = ~n1440 & ~n1446;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = ~n1452 & n1455;
  assign n1461 = n1452 & ~n1455;
  assign n1462 = ~n1460 & ~n1461;
  assign n1463 = n1449 & n1456;
  assign n1464 = ~n1449 & ~n1456;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = ~n1462 & ~n1465;
  assign n1467 = ~n1459 & ~n1466;
  assign n1468 = pi3  & pi4 ;
  assign n1469 = pi3  & ~pi4 ;
  assign n1470 = ~pi3  & pi4 ;
  assign n1471 = ~n1469 & ~n1470;
  assign n1472 = pi5  & ~n1471;
  assign n1473 = ~n1468 & ~n1472;
  assign n1474 = pi0  & pi1 ;
  assign n1475 = ~pi0  & pi1 ;
  assign n1476 = pi0  & ~pi1 ;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = pi2  & ~n1477;
  assign n1479 = ~n1474 & ~n1478;
  assign n1480 = ~n1473 & n1479;
  assign n1481 = n1473 & ~n1479;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = ~pi5  & ~n1471;
  assign n1484 = pi5  & n1471;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = ~pi2  & ~n1477;
  assign n1487 = pi2  & n1477;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = ~pi6  & ~n1488;
  assign n1490 = pi6  & n1488;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = ~n1485 & ~n1491;
  assign n1493 = pi6  & ~n1488;
  assign n1494 = ~n1492 & ~n1493;
  assign n1495 = ~n1482 & ~n1494;
  assign n1496 = ~n1473 & ~n1479;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = n1482 & n1494;
  assign n1499 = ~n1495 & ~n1498;
  assign n1500 = ~pi997  & pi998 ;
  assign n1501 = pi997  & ~pi998 ;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = ~pi999  & ~n1502;
  assign n1504 = pi999  & n1502;
  assign n1505 = ~n1503 & ~n1504;
  assign n1506 = n1485 & ~n1491;
  assign n1507 = ~n1485 & n1491;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = ~n1505 & ~n1508;
  assign n1510 = ~n1499 & ~n1509;
  assign n1511 = pi997  & pi998 ;
  assign n1512 = pi999  & ~n1502;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = n1499 & n1509;
  assign n1515 = ~n1510 & ~n1514;
  assign n1516 = n1513 & n1515;
  assign n1517 = ~n1510 & ~n1516;
  assign n1518 = n1497 & n1517;
  assign n1519 = ~n1497 & ~n1517;
  assign n1520 = ~n1518 & ~n1519;
  assign n1521 = n1505 & ~n1508;
  assign n1522 = ~n1505 & n1508;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = ~n1462 & ~n1523;
  assign n1525 = ~n1513 & ~n1515;
  assign n1526 = ~n1516 & ~n1525;
  assign n1527 = ~n1524 & n1526;
  assign n1528 = n1524 & ~n1526;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = n1465 & n1529;
  assign n1531 = ~n1527 & ~n1530;
  assign n1532 = n1520 & ~n1531;
  assign n1533 = n1467 & ~n1532;
  assign n1534 = ~n1497 & n1517;
  assign n1535 = n1533 & n1534;
  assign n1536 = pi19  & ~pi20 ;
  assign n1537 = ~pi19  & pi20 ;
  assign n1538 = ~n1536 & ~n1537;
  assign n1539 = ~pi21  & ~n1538;
  assign n1540 = pi21  & n1538;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = pi22  & ~pi23 ;
  assign n1543 = ~pi22  & pi23 ;
  assign n1544 = ~n1542 & ~n1543;
  assign n1545 = ~pi24  & ~n1544;
  assign n1546 = pi24  & n1544;
  assign n1547 = ~n1545 & ~n1546;
  assign n1548 = ~n1541 & ~n1547;
  assign n1549 = pi22  & pi23 ;
  assign n1550 = pi24  & ~n1544;
  assign n1551 = ~n1549 & ~n1550;
  assign n1552 = pi19  & pi20 ;
  assign n1553 = pi21  & ~n1538;
  assign n1554 = ~n1552 & ~n1553;
  assign n1555 = n1551 & ~n1554;
  assign n1556 = ~n1551 & n1554;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = n1548 & ~n1557;
  assign n1559 = ~n1551 & ~n1554;
  assign n1560 = ~n1558 & ~n1559;
  assign n1561 = pi28  & pi29 ;
  assign n1562 = pi28  & ~pi29 ;
  assign n1563 = ~pi28  & pi29 ;
  assign n1564 = ~n1562 & ~n1563;
  assign n1565 = pi30  & ~n1564;
  assign n1566 = ~n1561 & ~n1565;
  assign n1567 = pi25  & pi26 ;
  assign n1568 = pi25  & ~pi26 ;
  assign n1569 = ~pi25  & pi26 ;
  assign n1570 = ~n1568 & ~n1569;
  assign n1571 = pi27  & ~n1570;
  assign n1572 = ~n1567 & ~n1571;
  assign n1573 = ~n1566 & n1572;
  assign n1574 = n1566 & ~n1572;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = ~pi27  & ~n1570;
  assign n1577 = pi27  & n1570;
  assign n1578 = ~n1576 & ~n1577;
  assign n1579 = ~pi30  & ~n1564;
  assign n1580 = pi30  & n1564;
  assign n1581 = ~n1579 & ~n1580;
  assign n1582 = ~n1578 & ~n1581;
  assign n1583 = ~n1575 & n1582;
  assign n1584 = ~n1566 & ~n1572;
  assign n1585 = ~n1583 & ~n1584;
  assign n1586 = n1575 & n1582;
  assign n1587 = ~n1575 & ~n1582;
  assign n1588 = ~n1586 & ~n1587;
  assign n1589 = ~n1585 & ~n1588;
  assign n1590 = n1548 & n1557;
  assign n1591 = ~n1548 & ~n1557;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = ~n1560 & ~n1592;
  assign n1594 = ~n1541 & n1547;
  assign n1595 = n1541 & ~n1547;
  assign n1596 = ~n1594 & ~n1595;
  assign n1597 = ~n1578 & n1581;
  assign n1598 = n1578 & ~n1581;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = ~n1596 & ~n1599;
  assign n1601 = ~n1589 & n1600;
  assign n1602 = ~n1593 & n1601;
  assign n1603 = ~n1588 & n1602;
  assign n1604 = n1588 & ~n1602;
  assign n1605 = ~n1592 & ~n1604;
  assign n1606 = ~n1603 & ~n1605;
  assign n1607 = n1585 & n1606;
  assign n1608 = ~n1560 & ~n1607;
  assign n1609 = ~n1585 & ~n1606;
  assign n1610 = ~n1608 & ~n1609;
  assign n1611 = pi7  & ~pi8 ;
  assign n1612 = ~pi7  & pi8 ;
  assign n1613 = ~n1611 & ~n1612;
  assign n1614 = ~pi9  & ~n1613;
  assign n1615 = pi9  & n1613;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = pi10  & ~pi11 ;
  assign n1618 = ~pi10  & pi11 ;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = ~pi12  & ~n1619;
  assign n1621 = pi12  & n1619;
  assign n1622 = ~n1620 & ~n1621;
  assign n1623 = ~n1616 & ~n1622;
  assign n1624 = pi10  & pi11 ;
  assign n1625 = pi12  & ~n1619;
  assign n1626 = ~n1624 & ~n1625;
  assign n1627 = pi7  & pi8 ;
  assign n1628 = pi9  & ~n1613;
  assign n1629 = ~n1627 & ~n1628;
  assign n1630 = n1626 & ~n1629;
  assign n1631 = ~n1626 & n1629;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = n1623 & ~n1632;
  assign n1634 = ~n1626 & ~n1629;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = pi16  & pi17 ;
  assign n1637 = pi16  & ~pi17 ;
  assign n1638 = ~pi16  & pi17 ;
  assign n1639 = ~n1637 & ~n1638;
  assign n1640 = pi18  & ~n1639;
  assign n1641 = ~n1636 & ~n1640;
  assign n1642 = pi13  & pi14 ;
  assign n1643 = pi13  & ~pi14 ;
  assign n1644 = ~pi13  & pi14 ;
  assign n1645 = ~n1643 & ~n1644;
  assign n1646 = pi15  & ~n1645;
  assign n1647 = ~n1642 & ~n1646;
  assign n1648 = ~n1641 & n1647;
  assign n1649 = n1641 & ~n1647;
  assign n1650 = ~n1648 & ~n1649;
  assign n1651 = ~pi15  & ~n1645;
  assign n1652 = pi15  & n1645;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = ~pi18  & ~n1639;
  assign n1655 = pi18  & n1639;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = ~n1653 & ~n1656;
  assign n1658 = ~n1650 & n1657;
  assign n1659 = ~n1641 & ~n1647;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = n1650 & n1657;
  assign n1662 = ~n1650 & ~n1657;
  assign n1663 = ~n1661 & ~n1662;
  assign n1664 = ~n1660 & ~n1663;
  assign n1665 = n1623 & n1632;
  assign n1666 = ~n1623 & ~n1632;
  assign n1667 = ~n1665 & ~n1666;
  assign n1668 = ~n1635 & ~n1667;
  assign n1669 = ~n1616 & n1622;
  assign n1670 = n1616 & ~n1622;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = ~n1653 & n1656;
  assign n1673 = n1653 & ~n1656;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675 = ~n1671 & ~n1674;
  assign n1676 = ~n1664 & n1675;
  assign n1677 = ~n1668 & n1676;
  assign n1678 = ~n1663 & n1677;
  assign n1679 = n1663 & ~n1677;
  assign n1680 = ~n1667 & ~n1679;
  assign n1681 = ~n1678 & ~n1680;
  assign n1682 = n1660 & n1681;
  assign n1683 = ~n1635 & ~n1682;
  assign n1684 = ~n1660 & ~n1681;
  assign n1685 = ~n1683 & ~n1684;
  assign n1686 = n1610 & n1685;
  assign n1687 = ~n1635 & n1660;
  assign n1688 = n1635 & ~n1660;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = ~n1681 & ~n1689;
  assign n1691 = n1681 & n1689;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = ~n1560 & n1585;
  assign n1694 = n1560 & ~n1585;
  assign n1695 = ~n1693 & ~n1694;
  assign n1696 = ~n1606 & ~n1695;
  assign n1697 = n1606 & n1695;
  assign n1698 = ~n1696 & ~n1697;
  assign n1699 = n1692 & n1698;
  assign n1700 = ~n1596 & n1599;
  assign n1701 = n1596 & ~n1599;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n1671 & n1674;
  assign n1704 = n1671 & ~n1674;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = ~n1702 & ~n1705;
  assign n1707 = ~n1603 & ~n1604;
  assign n1708 = ~n1592 & ~n1707;
  assign n1709 = n1592 & n1707;
  assign n1710 = ~n1708 & ~n1709;
  assign n1711 = n1706 & ~n1710;
  assign n1712 = ~n1678 & ~n1679;
  assign n1713 = n1667 & n1712;
  assign n1714 = ~n1667 & ~n1712;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = ~n1706 & n1710;
  assign n1717 = ~n1715 & ~n1716;
  assign n1718 = ~n1711 & ~n1717;
  assign n1719 = ~n1692 & ~n1698;
  assign n1720 = ~n1699 & ~n1719;
  assign n1721 = ~n1718 & n1720;
  assign n1722 = ~n1699 & ~n1721;
  assign n1723 = ~n1686 & ~n1722;
  assign n1724 = ~n1610 & ~n1685;
  assign n1725 = ~n1723 & ~n1724;
  assign n1726 = n1535 & ~n1725;
  assign n1727 = ~n1535 & n1725;
  assign n1728 = ~n1726 & ~n1727;
  assign n1729 = ~n1520 & n1531;
  assign n1730 = ~n1534 & ~n1729;
  assign n1731 = ~n1533 & n1730;
  assign n1732 = ~n1535 & ~n1731;
  assign n1733 = ~n1686 & ~n1724;
  assign n1734 = ~n1722 & n1733;
  assign n1735 = n1722 & ~n1733;
  assign n1736 = ~n1734 & ~n1735;
  assign n1737 = n1732 & n1736;
  assign n1738 = ~n1702 & n1705;
  assign n1739 = n1702 & ~n1705;
  assign n1740 = ~n1738 & ~n1739;
  assign n1741 = ~n1462 & n1523;
  assign n1742 = n1462 & ~n1523;
  assign n1743 = ~n1741 & ~n1742;
  assign n1744 = ~n1740 & ~n1743;
  assign n1745 = ~n1711 & ~n1716;
  assign n1746 = ~n1715 & ~n1745;
  assign n1747 = n1715 & n1745;
  assign n1748 = ~n1746 & ~n1747;
  assign n1749 = n1744 & ~n1748;
  assign n1750 = ~n1465 & ~n1529;
  assign n1751 = ~n1530 & ~n1750;
  assign n1752 = ~n1744 & n1748;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = ~n1749 & ~n1753;
  assign n1755 = ~n1467 & ~n1520;
  assign n1756 = n1467 & n1520;
  assign n1757 = ~n1755 & ~n1756;
  assign n1758 = n1531 & ~n1757;
  assign n1759 = ~n1531 & n1757;
  assign n1760 = ~n1758 & ~n1759;
  assign n1761 = n1718 & ~n1720;
  assign n1762 = ~n1721 & ~n1761;
  assign n1763 = ~n1760 & ~n1762;
  assign n1764 = ~n1754 & ~n1763;
  assign n1765 = n1760 & n1762;
  assign n1766 = ~n1764 & ~n1765;
  assign n1767 = ~n1732 & ~n1736;
  assign n1768 = ~n1737 & ~n1767;
  assign n1769 = ~n1766 & n1768;
  assign n1770 = ~n1737 & ~n1769;
  assign n1771 = n1728 & ~n1770;
  assign n1772 = ~n1726 & ~n1771;
  assign n1773 = n1434 & n1772;
  assign n1774 = ~n1434 & ~n1772;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = ~n1728 & n1770;
  assign n1777 = ~n1771 & ~n1776;
  assign n1778 = n1430 & ~n1432;
  assign n1779 = ~n1433 & ~n1778;
  assign n1780 = n1777 & n1779;
  assign n1781 = ~n1763 & ~n1765;
  assign n1782 = ~n1754 & n1781;
  assign n1783 = n1754 & ~n1781;
  assign n1784 = ~n1782 & ~n1783;
  assign n1785 = ~n1424 & ~n1426;
  assign n1786 = ~n1417 & n1785;
  assign n1787 = n1417 & ~n1785;
  assign n1788 = ~n1786 & ~n1787;
  assign n1789 = n1784 & n1788;
  assign n1790 = ~n1401 & n1404;
  assign n1791 = n1401 & ~n1404;
  assign n1792 = ~n1790 & ~n1791;
  assign n1793 = ~n1740 & n1743;
  assign n1794 = n1740 & ~n1743;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = ~n1792 & ~n1795;
  assign n1797 = ~n1410 & ~n1415;
  assign n1798 = ~n1414 & ~n1797;
  assign n1799 = n1414 & n1797;
  assign n1800 = ~n1798 & ~n1799;
  assign n1801 = n1796 & ~n1800;
  assign n1802 = ~n1749 & ~n1752;
  assign n1803 = n1751 & n1802;
  assign n1804 = ~n1751 & ~n1802;
  assign n1805 = ~n1803 & ~n1804;
  assign n1806 = ~n1796 & n1800;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = ~n1801 & ~n1807;
  assign n1809 = ~n1784 & ~n1788;
  assign n1810 = ~n1789 & ~n1809;
  assign n1811 = ~n1808 & n1810;
  assign n1812 = ~n1789 & ~n1811;
  assign n1813 = ~n1398 & ~n1428;
  assign n1814 = ~n1427 & n1813;
  assign n1815 = n1427 & ~n1813;
  assign n1816 = ~n1814 & ~n1815;
  assign n1817 = n1766 & ~n1768;
  assign n1818 = ~n1769 & ~n1817;
  assign n1819 = ~n1816 & ~n1818;
  assign n1820 = ~n1812 & ~n1819;
  assign n1821 = n1816 & n1818;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = ~n1777 & ~n1779;
  assign n1824 = ~n1780 & ~n1823;
  assign n1825 = ~n1822 & n1824;
  assign n1826 = ~n1780 & ~n1825;
  assign n1827 = n1775 & ~n1826;
  assign n1828 = ~n1775 & n1826;
  assign n1829 = ~n1827 & ~n1828;
  assign n1830 = pi979  & ~pi980 ;
  assign n1831 = ~pi979  & pi980 ;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = ~pi981  & ~n1832;
  assign n1834 = pi981  & n1832;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = pi982  & ~pi983 ;
  assign n1837 = ~pi982  & pi983 ;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = ~pi984  & ~n1838;
  assign n1840 = pi984  & n1838;
  assign n1841 = ~n1839 & ~n1840;
  assign n1842 = ~n1835 & ~n1841;
  assign n1843 = pi982  & pi983 ;
  assign n1844 = pi984  & ~n1838;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = pi979  & pi980 ;
  assign n1847 = pi981  & ~n1832;
  assign n1848 = ~n1846 & ~n1847;
  assign n1849 = n1845 & ~n1848;
  assign n1850 = ~n1845 & n1848;
  assign n1851 = ~n1849 & ~n1850;
  assign n1852 = n1842 & ~n1851;
  assign n1853 = ~n1845 & ~n1848;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = pi988  & pi989 ;
  assign n1856 = pi988  & ~pi989 ;
  assign n1857 = ~pi988  & pi989 ;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = pi990  & ~n1858;
  assign n1860 = ~n1855 & ~n1859;
  assign n1861 = pi985  & pi986 ;
  assign n1862 = pi985  & ~pi986 ;
  assign n1863 = ~pi985  & pi986 ;
  assign n1864 = ~n1862 & ~n1863;
  assign n1865 = pi987  & ~n1864;
  assign n1866 = ~n1861 & ~n1865;
  assign n1867 = ~n1860 & n1866;
  assign n1868 = n1860 & ~n1866;
  assign n1869 = ~n1867 & ~n1868;
  assign n1870 = ~pi987  & ~n1864;
  assign n1871 = pi987  & n1864;
  assign n1872 = ~n1870 & ~n1871;
  assign n1873 = ~pi990  & ~n1858;
  assign n1874 = pi990  & n1858;
  assign n1875 = ~n1873 & ~n1874;
  assign n1876 = ~n1872 & ~n1875;
  assign n1877 = ~n1869 & n1876;
  assign n1878 = ~n1860 & ~n1866;
  assign n1879 = ~n1877 & ~n1878;
  assign n1880 = n1869 & n1876;
  assign n1881 = ~n1869 & ~n1876;
  assign n1882 = ~n1880 & ~n1881;
  assign n1883 = ~n1879 & ~n1882;
  assign n1884 = n1842 & n1851;
  assign n1885 = ~n1842 & ~n1851;
  assign n1886 = ~n1884 & ~n1885;
  assign n1887 = ~n1854 & ~n1886;
  assign n1888 = ~n1835 & n1841;
  assign n1889 = n1835 & ~n1841;
  assign n1890 = ~n1888 & ~n1889;
  assign n1891 = ~n1872 & n1875;
  assign n1892 = n1872 & ~n1875;
  assign n1893 = ~n1891 & ~n1892;
  assign n1894 = ~n1890 & ~n1893;
  assign n1895 = ~n1883 & n1894;
  assign n1896 = ~n1887 & n1895;
  assign n1897 = n1882 & ~n1896;
  assign n1898 = ~n1882 & n1896;
  assign n1899 = ~n1897 & ~n1898;
  assign n1900 = n1886 & n1899;
  assign n1901 = ~n1897 & ~n1900;
  assign n1902 = n1879 & ~n1901;
  assign n1903 = ~n1854 & ~n1902;
  assign n1904 = ~n1879 & n1901;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = pi967  & ~pi968 ;
  assign n1907 = ~pi967  & pi968 ;
  assign n1908 = ~n1906 & ~n1907;
  assign n1909 = ~pi969  & ~n1908;
  assign n1910 = pi969  & n1908;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = pi970  & ~pi971 ;
  assign n1913 = ~pi970  & pi971 ;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = ~pi972  & ~n1914;
  assign n1916 = pi972  & n1914;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = ~n1911 & ~n1917;
  assign n1919 = pi970  & pi971 ;
  assign n1920 = pi972  & ~n1914;
  assign n1921 = ~n1919 & ~n1920;
  assign n1922 = pi967  & pi968 ;
  assign n1923 = pi969  & ~n1908;
  assign n1924 = ~n1922 & ~n1923;
  assign n1925 = n1921 & ~n1924;
  assign n1926 = ~n1921 & n1924;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = n1918 & ~n1927;
  assign n1929 = ~n1921 & ~n1924;
  assign n1930 = ~n1928 & ~n1929;
  assign n1931 = pi976  & pi977 ;
  assign n1932 = pi976  & ~pi977 ;
  assign n1933 = ~pi976  & pi977 ;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = pi978  & ~n1934;
  assign n1936 = ~n1931 & ~n1935;
  assign n1937 = pi973  & pi974 ;
  assign n1938 = pi973  & ~pi974 ;
  assign n1939 = ~pi973  & pi974 ;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = pi975  & ~n1940;
  assign n1942 = ~n1937 & ~n1941;
  assign n1943 = ~n1936 & n1942;
  assign n1944 = n1936 & ~n1942;
  assign n1945 = ~n1943 & ~n1944;
  assign n1946 = ~pi975  & ~n1940;
  assign n1947 = pi975  & n1940;
  assign n1948 = ~n1946 & ~n1947;
  assign n1949 = ~pi978  & ~n1934;
  assign n1950 = pi978  & n1934;
  assign n1951 = ~n1949 & ~n1950;
  assign n1952 = ~n1948 & ~n1951;
  assign n1953 = ~n1945 & n1952;
  assign n1954 = ~n1936 & ~n1942;
  assign n1955 = ~n1953 & ~n1954;
  assign n1956 = n1945 & n1952;
  assign n1957 = ~n1945 & ~n1952;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = ~n1955 & ~n1958;
  assign n1960 = n1918 & n1927;
  assign n1961 = ~n1918 & ~n1927;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = ~n1930 & ~n1962;
  assign n1964 = ~n1911 & n1917;
  assign n1965 = n1911 & ~n1917;
  assign n1966 = ~n1964 & ~n1965;
  assign n1967 = ~n1948 & n1951;
  assign n1968 = n1948 & ~n1951;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = ~n1966 & ~n1969;
  assign n1971 = ~n1959 & n1970;
  assign n1972 = ~n1963 & n1971;
  assign n1973 = n1958 & ~n1972;
  assign n1974 = ~n1958 & n1972;
  assign n1975 = ~n1973 & ~n1974;
  assign n1976 = n1962 & n1975;
  assign n1977 = ~n1973 & ~n1976;
  assign n1978 = n1955 & ~n1977;
  assign n1979 = ~n1930 & ~n1978;
  assign n1980 = ~n1955 & n1977;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = n1905 & n1981;
  assign n1983 = ~n1930 & n1955;
  assign n1984 = n1930 & ~n1955;
  assign n1985 = ~n1983 & ~n1984;
  assign n1986 = n1977 & ~n1985;
  assign n1987 = ~n1977 & n1985;
  assign n1988 = ~n1986 & ~n1987;
  assign n1989 = ~n1854 & n1879;
  assign n1990 = n1854 & ~n1879;
  assign n1991 = ~n1989 & ~n1990;
  assign n1992 = n1901 & ~n1991;
  assign n1993 = ~n1901 & n1991;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = n1988 & n1994;
  assign n1996 = ~n1890 & n1893;
  assign n1997 = n1890 & ~n1893;
  assign n1998 = ~n1996 & ~n1997;
  assign n1999 = ~n1966 & n1969;
  assign n2000 = n1966 & ~n1969;
  assign n2001 = ~n1999 & ~n2000;
  assign n2002 = ~n1998 & ~n2001;
  assign n2003 = ~n1886 & ~n1899;
  assign n2004 = ~n1900 & ~n2003;
  assign n2005 = ~n2002 & n2004;
  assign n2006 = ~n1962 & ~n1975;
  assign n2007 = ~n1976 & ~n2006;
  assign n2008 = ~n2002 & ~n2004;
  assign n2009 = n2004 & ~n2005;
  assign n2010 = ~n2008 & ~n2009;
  assign n2011 = n2007 & ~n2010;
  assign n2012 = ~n2005 & ~n2011;
  assign n2013 = ~n1988 & ~n1994;
  assign n2014 = ~n1995 & ~n2013;
  assign n2015 = n2012 & n2014;
  assign n2016 = ~n1995 & ~n2015;
  assign n2017 = ~n1982 & ~n2016;
  assign n2018 = ~n1905 & ~n1981;
  assign n2019 = ~n2017 & ~n2018;
  assign n2020 = pi958  & pi959 ;
  assign n2021 = ~pi958  & pi959 ;
  assign n2022 = pi958  & ~pi959 ;
  assign n2023 = ~n2021 & ~n2022;
  assign n2024 = pi960  & ~n2023;
  assign n2025 = ~n2020 & ~n2024;
  assign n2026 = pi955  & pi956 ;
  assign n2027 = ~pi955  & pi956 ;
  assign n2028 = pi955  & ~pi956 ;
  assign n2029 = ~n2027 & ~n2028;
  assign n2030 = pi957  & ~n2029;
  assign n2031 = ~n2026 & ~n2030;
  assign n2032 = ~n2025 & n2031;
  assign n2033 = n2025 & ~n2031;
  assign n2034 = ~n2032 & ~n2033;
  assign n2035 = ~pi957  & ~n2029;
  assign n2036 = pi957  & n2029;
  assign n2037 = ~n2035 & ~n2036;
  assign n2038 = ~pi960  & ~n2023;
  assign n2039 = pi960  & n2023;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = ~n2037 & ~n2040;
  assign n2042 = ~n2034 & n2041;
  assign n2043 = ~n2025 & ~n2031;
  assign n2044 = ~n2042 & ~n2043;
  assign n2045 = pi964  & pi965 ;
  assign n2046 = ~pi964  & pi965 ;
  assign n2047 = pi964  & ~pi965 ;
  assign n2048 = ~n2046 & ~n2047;
  assign n2049 = pi966  & ~n2048;
  assign n2050 = ~n2045 & ~n2049;
  assign n2051 = pi961  & pi962 ;
  assign n2052 = ~pi961  & pi962 ;
  assign n2053 = pi961  & ~pi962 ;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = pi963  & ~n2054;
  assign n2056 = ~n2051 & ~n2055;
  assign n2057 = ~n2050 & n2056;
  assign n2058 = n2050 & ~n2056;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = ~pi963  & ~n2054;
  assign n2061 = pi963  & n2054;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = ~pi966  & ~n2048;
  assign n2064 = pi966  & n2048;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = ~n2062 & ~n2065;
  assign n2067 = ~n2059 & n2066;
  assign n2068 = ~n2050 & ~n2056;
  assign n2069 = ~n2067 & ~n2068;
  assign n2070 = n2059 & n2066;
  assign n2071 = ~n2059 & ~n2066;
  assign n2072 = ~n2070 & ~n2071;
  assign n2073 = n2034 & n2041;
  assign n2074 = ~n2034 & ~n2041;
  assign n2075 = ~n2073 & ~n2074;
  assign n2076 = ~n2044 & ~n2075;
  assign n2077 = ~n2069 & ~n2072;
  assign n2078 = ~n2062 & n2065;
  assign n2079 = n2062 & ~n2065;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = ~n2037 & n2040;
  assign n2082 = n2037 & ~n2040;
  assign n2083 = ~n2081 & ~n2082;
  assign n2084 = ~n2080 & ~n2083;
  assign n2085 = ~n2076 & n2084;
  assign n2086 = ~n2077 & n2085;
  assign n2087 = n2072 & ~n2086;
  assign n2088 = ~n2072 & n2086;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = n2075 & n2089;
  assign n2091 = ~n2087 & ~n2090;
  assign n2092 = n2069 & ~n2091;
  assign n2093 = ~n2044 & ~n2092;
  assign n2094 = ~n2069 & n2091;
  assign n2095 = ~n2093 & ~n2094;
  assign n2096 = pi946  & pi947 ;
  assign n2097 = ~pi946  & pi947 ;
  assign n2098 = pi946  & ~pi947 ;
  assign n2099 = ~n2097 & ~n2098;
  assign n2100 = pi948  & ~n2099;
  assign n2101 = ~n2096 & ~n2100;
  assign n2102 = pi943  & pi944 ;
  assign n2103 = ~pi943  & pi944 ;
  assign n2104 = pi943  & ~pi944 ;
  assign n2105 = ~n2103 & ~n2104;
  assign n2106 = pi945  & ~n2105;
  assign n2107 = ~n2102 & ~n2106;
  assign n2108 = ~n2101 & n2107;
  assign n2109 = n2101 & ~n2107;
  assign n2110 = ~n2108 & ~n2109;
  assign n2111 = ~pi945  & ~n2105;
  assign n2112 = pi945  & n2105;
  assign n2113 = ~n2111 & ~n2112;
  assign n2114 = ~pi948  & ~n2099;
  assign n2115 = pi948  & n2099;
  assign n2116 = ~n2114 & ~n2115;
  assign n2117 = ~n2113 & ~n2116;
  assign n2118 = ~n2110 & n2117;
  assign n2119 = ~n2101 & ~n2107;
  assign n2120 = ~n2118 & ~n2119;
  assign n2121 = pi952  & pi953 ;
  assign n2122 = ~pi952  & pi953 ;
  assign n2123 = pi952  & ~pi953 ;
  assign n2124 = ~n2122 & ~n2123;
  assign n2125 = pi954  & ~n2124;
  assign n2126 = ~n2121 & ~n2125;
  assign n2127 = pi949  & pi950 ;
  assign n2128 = ~pi949  & pi950 ;
  assign n2129 = pi949  & ~pi950 ;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = pi951  & ~n2130;
  assign n2132 = ~n2127 & ~n2131;
  assign n2133 = ~n2126 & n2132;
  assign n2134 = n2126 & ~n2132;
  assign n2135 = ~n2133 & ~n2134;
  assign n2136 = ~pi951  & ~n2130;
  assign n2137 = pi951  & n2130;
  assign n2138 = ~n2136 & ~n2137;
  assign n2139 = ~pi954  & ~n2124;
  assign n2140 = pi954  & n2124;
  assign n2141 = ~n2139 & ~n2140;
  assign n2142 = ~n2138 & ~n2141;
  assign n2143 = ~n2135 & n2142;
  assign n2144 = ~n2126 & ~n2132;
  assign n2145 = ~n2143 & ~n2144;
  assign n2146 = n2135 & n2142;
  assign n2147 = ~n2135 & ~n2142;
  assign n2148 = ~n2146 & ~n2147;
  assign n2149 = n2110 & n2117;
  assign n2150 = ~n2110 & ~n2117;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = ~n2120 & ~n2151;
  assign n2153 = ~n2145 & ~n2148;
  assign n2154 = ~n2138 & n2141;
  assign n2155 = n2138 & ~n2141;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = ~n2113 & n2116;
  assign n2158 = n2113 & ~n2116;
  assign n2159 = ~n2157 & ~n2158;
  assign n2160 = ~n2156 & ~n2159;
  assign n2161 = ~n2152 & n2160;
  assign n2162 = ~n2153 & n2161;
  assign n2163 = n2148 & ~n2162;
  assign n2164 = ~n2148 & n2162;
  assign n2165 = ~n2163 & ~n2164;
  assign n2166 = n2151 & n2165;
  assign n2167 = ~n2163 & ~n2166;
  assign n2168 = n2145 & ~n2167;
  assign n2169 = ~n2120 & ~n2168;
  assign n2170 = ~n2145 & n2167;
  assign n2171 = ~n2169 & ~n2170;
  assign n2172 = n2095 & n2171;
  assign n2173 = ~n2120 & n2145;
  assign n2174 = n2120 & ~n2145;
  assign n2175 = ~n2173 & ~n2174;
  assign n2176 = n2167 & ~n2175;
  assign n2177 = ~n2167 & n2175;
  assign n2178 = ~n2176 & ~n2177;
  assign n2179 = ~n2044 & n2069;
  assign n2180 = n2044 & ~n2069;
  assign n2181 = ~n2179 & ~n2180;
  assign n2182 = n2091 & ~n2181;
  assign n2183 = ~n2091 & n2181;
  assign n2184 = ~n2182 & ~n2183;
  assign n2185 = n2178 & n2184;
  assign n2186 = n2080 & ~n2083;
  assign n2187 = ~n2080 & n2083;
  assign n2188 = ~n2186 & ~n2187;
  assign n2189 = n2156 & ~n2159;
  assign n2190 = ~n2156 & n2159;
  assign n2191 = ~n2189 & ~n2190;
  assign n2192 = ~n2188 & ~n2191;
  assign n2193 = ~n2075 & ~n2089;
  assign n2194 = ~n2090 & ~n2193;
  assign n2195 = ~n2192 & n2194;
  assign n2196 = ~n2151 & ~n2165;
  assign n2197 = ~n2166 & ~n2196;
  assign n2198 = n2192 & ~n2194;
  assign n2199 = ~n2195 & ~n2198;
  assign n2200 = n2197 & n2199;
  assign n2201 = ~n2195 & ~n2200;
  assign n2202 = ~n2178 & ~n2184;
  assign n2203 = ~n2185 & ~n2202;
  assign n2204 = n2201 & n2203;
  assign n2205 = ~n2185 & ~n2204;
  assign n2206 = ~n2172 & ~n2205;
  assign n2207 = ~n2095 & ~n2171;
  assign n2208 = ~n2206 & ~n2207;
  assign n2209 = ~n2019 & ~n2208;
  assign n2210 = n2019 & n2208;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = ~n1982 & ~n2018;
  assign n2213 = ~n2016 & n2212;
  assign n2214 = n2016 & ~n2212;
  assign n2215 = ~n2213 & ~n2214;
  assign n2216 = ~n2172 & ~n2207;
  assign n2217 = ~n2205 & n2216;
  assign n2218 = n2205 & ~n2216;
  assign n2219 = ~n2217 & ~n2218;
  assign n2220 = n2215 & n2219;
  assign n2221 = ~n2201 & ~n2203;
  assign n2222 = ~n2204 & ~n2221;
  assign n2223 = ~n2012 & ~n2014;
  assign n2224 = ~n2015 & ~n2223;
  assign n2225 = n2222 & n2224;
  assign n2226 = ~n2222 & ~n2224;
  assign n2227 = ~n2225 & ~n2226;
  assign n2228 = ~n1998 & n2001;
  assign n2229 = n1998 & ~n2001;
  assign n2230 = ~n2228 & ~n2229;
  assign n2231 = ~n2188 & n2191;
  assign n2232 = n2188 & ~n2191;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = ~n2230 & ~n2233;
  assign n2235 = ~n2007 & n2010;
  assign n2236 = ~n2011 & ~n2235;
  assign n2237 = ~n2234 & n2236;
  assign n2238 = ~n2197 & ~n2199;
  assign n2239 = ~n2200 & ~n2238;
  assign n2240 = n2234 & ~n2236;
  assign n2241 = ~n2237 & ~n2240;
  assign n2242 = n2239 & n2241;
  assign n2243 = ~n2237 & ~n2242;
  assign n2244 = n2227 & n2243;
  assign n2245 = ~n2225 & ~n2244;
  assign n2246 = ~n2215 & ~n2219;
  assign n2247 = ~n2220 & ~n2246;
  assign n2248 = ~n2245 & n2247;
  assign n2249 = ~n2220 & ~n2248;
  assign n2250 = n2211 & ~n2249;
  assign n2251 = ~n2209 & ~n2250;
  assign n2252 = n1829 & ~n2251;
  assign n2253 = ~n2211 & n2249;
  assign n2254 = ~n2250 & ~n2253;
  assign n2255 = n1822 & ~n1824;
  assign n2256 = ~n1825 & ~n2255;
  assign n2257 = n2254 & n2256;
  assign n2258 = ~n2227 & ~n2243;
  assign n2259 = ~n2244 & ~n2258;
  assign n2260 = n1808 & ~n1810;
  assign n2261 = ~n1811 & ~n2260;
  assign n2262 = n2259 & n2261;
  assign n2263 = ~n1792 & n1795;
  assign n2264 = n1792 & ~n1795;
  assign n2265 = ~n2263 & ~n2264;
  assign n2266 = ~n2230 & n2233;
  assign n2267 = n2230 & ~n2233;
  assign n2268 = ~n2266 & ~n2267;
  assign n2269 = ~n2265 & ~n2268;
  assign n2270 = ~n1801 & ~n1806;
  assign n2271 = n1805 & n2270;
  assign n2272 = ~n1805 & ~n2270;
  assign n2273 = ~n2271 & ~n2272;
  assign n2274 = n2269 & ~n2273;
  assign n2275 = ~n2239 & ~n2241;
  assign n2276 = ~n2242 & ~n2275;
  assign n2277 = ~n2269 & n2273;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = ~n2274 & ~n2278;
  assign n2280 = ~n2259 & ~n2261;
  assign n2281 = ~n2262 & ~n2280;
  assign n2282 = ~n2279 & n2281;
  assign n2283 = ~n2262 & ~n2282;
  assign n2284 = ~n1819 & ~n1821;
  assign n2285 = ~n1812 & n2284;
  assign n2286 = n1812 & ~n2284;
  assign n2287 = ~n2285 & ~n2286;
  assign n2288 = n2245 & ~n2247;
  assign n2289 = ~n2248 & ~n2288;
  assign n2290 = ~n2287 & ~n2289;
  assign n2291 = ~n2283 & ~n2290;
  assign n2292 = ~n2285 & n2289;
  assign n2293 = ~n2286 & n2292;
  assign n2294 = ~n2291 & ~n2293;
  assign n2295 = ~n2254 & ~n2256;
  assign n2296 = ~n2257 & ~n2295;
  assign n2297 = ~n2294 & n2296;
  assign n2298 = ~n2257 & ~n2297;
  assign n2299 = ~n1829 & n2251;
  assign n2300 = ~n2252 & ~n2299;
  assign n2301 = ~n2298 & n2300;
  assign n2302 = ~n2252 & ~n2301;
  assign n2303 = ~n1774 & ~n1827;
  assign n2304 = ~n2302 & ~n2303;
  assign n2305 = ~n2302 & n2303;
  assign n2306 = n2302 & ~n2303;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = pi934  & pi935 ;
  assign n2309 = ~pi934  & pi935 ;
  assign n2310 = pi934  & ~pi935 ;
  assign n2311 = ~n2309 & ~n2310;
  assign n2312 = pi936  & ~n2311;
  assign n2313 = ~n2308 & ~n2312;
  assign n2314 = pi931  & pi932 ;
  assign n2315 = ~pi931  & pi932 ;
  assign n2316 = pi931  & ~pi932 ;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = pi933  & ~n2317;
  assign n2319 = ~n2314 & ~n2318;
  assign n2320 = ~n2313 & n2319;
  assign n2321 = n2313 & ~n2319;
  assign n2322 = ~n2320 & ~n2321;
  assign n2323 = ~pi933  & ~n2317;
  assign n2324 = pi933  & n2317;
  assign n2325 = ~n2323 & ~n2324;
  assign n2326 = ~pi936  & ~n2311;
  assign n2327 = pi936  & n2311;
  assign n2328 = ~n2326 & ~n2327;
  assign n2329 = ~n2325 & ~n2328;
  assign n2330 = ~n2322 & n2329;
  assign n2331 = ~n2313 & ~n2319;
  assign n2332 = ~n2330 & ~n2331;
  assign n2333 = pi940  & pi941 ;
  assign n2334 = ~pi940  & pi941 ;
  assign n2335 = pi940  & ~pi941 ;
  assign n2336 = ~n2334 & ~n2335;
  assign n2337 = pi942  & ~n2336;
  assign n2338 = ~n2333 & ~n2337;
  assign n2339 = pi937  & pi938 ;
  assign n2340 = ~pi937  & pi938 ;
  assign n2341 = pi937  & ~pi938 ;
  assign n2342 = ~n2340 & ~n2341;
  assign n2343 = pi939  & ~n2342;
  assign n2344 = ~n2339 & ~n2343;
  assign n2345 = ~n2338 & n2344;
  assign n2346 = n2338 & ~n2344;
  assign n2347 = ~n2345 & ~n2346;
  assign n2348 = ~pi939  & ~n2342;
  assign n2349 = pi939  & n2342;
  assign n2350 = ~n2348 & ~n2349;
  assign n2351 = ~pi942  & ~n2336;
  assign n2352 = pi942  & n2336;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = ~n2350 & ~n2353;
  assign n2355 = ~n2347 & n2354;
  assign n2356 = ~n2338 & ~n2344;
  assign n2357 = ~n2355 & ~n2356;
  assign n2358 = n2347 & n2354;
  assign n2359 = ~n2347 & ~n2354;
  assign n2360 = ~n2358 & ~n2359;
  assign n2361 = n2322 & n2329;
  assign n2362 = ~n2322 & ~n2329;
  assign n2363 = ~n2361 & ~n2362;
  assign n2364 = ~n2332 & ~n2363;
  assign n2365 = ~n2357 & ~n2360;
  assign n2366 = ~n2350 & n2353;
  assign n2367 = n2350 & ~n2353;
  assign n2368 = ~n2366 & ~n2367;
  assign n2369 = ~n2325 & n2328;
  assign n2370 = n2325 & ~n2328;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = ~n2368 & ~n2371;
  assign n2373 = ~n2364 & n2372;
  assign n2374 = ~n2365 & n2373;
  assign n2375 = n2360 & ~n2374;
  assign n2376 = ~n2360 & n2374;
  assign n2377 = ~n2375 & ~n2376;
  assign n2378 = n2363 & n2377;
  assign n2379 = ~n2375 & ~n2378;
  assign n2380 = n2357 & ~n2379;
  assign n2381 = ~n2332 & ~n2380;
  assign n2382 = ~n2357 & n2379;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = pi922  & pi923 ;
  assign n2385 = ~pi922  & pi923 ;
  assign n2386 = pi922  & ~pi923 ;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = pi924  & ~n2387;
  assign n2389 = ~n2384 & ~n2388;
  assign n2390 = pi919  & pi920 ;
  assign n2391 = ~pi919  & pi920 ;
  assign n2392 = pi919  & ~pi920 ;
  assign n2393 = ~n2391 & ~n2392;
  assign n2394 = pi921  & ~n2393;
  assign n2395 = ~n2390 & ~n2394;
  assign n2396 = ~n2389 & n2395;
  assign n2397 = n2389 & ~n2395;
  assign n2398 = ~n2396 & ~n2397;
  assign n2399 = ~pi921  & ~n2393;
  assign n2400 = pi921  & n2393;
  assign n2401 = ~n2399 & ~n2400;
  assign n2402 = ~pi924  & ~n2387;
  assign n2403 = pi924  & n2387;
  assign n2404 = ~n2402 & ~n2403;
  assign n2405 = ~n2401 & ~n2404;
  assign n2406 = ~n2398 & n2405;
  assign n2407 = ~n2389 & ~n2395;
  assign n2408 = ~n2406 & ~n2407;
  assign n2409 = pi928  & pi929 ;
  assign n2410 = ~pi928  & pi929 ;
  assign n2411 = pi928  & ~pi929 ;
  assign n2412 = ~n2410 & ~n2411;
  assign n2413 = pi930  & ~n2412;
  assign n2414 = ~n2409 & ~n2413;
  assign n2415 = pi925  & pi926 ;
  assign n2416 = ~pi925  & pi926 ;
  assign n2417 = pi925  & ~pi926 ;
  assign n2418 = ~n2416 & ~n2417;
  assign n2419 = pi927  & ~n2418;
  assign n2420 = ~n2415 & ~n2419;
  assign n2421 = ~n2414 & n2420;
  assign n2422 = n2414 & ~n2420;
  assign n2423 = ~n2421 & ~n2422;
  assign n2424 = ~pi927  & ~n2418;
  assign n2425 = pi927  & n2418;
  assign n2426 = ~n2424 & ~n2425;
  assign n2427 = ~pi930  & ~n2412;
  assign n2428 = pi930  & n2412;
  assign n2429 = ~n2427 & ~n2428;
  assign n2430 = ~n2426 & ~n2429;
  assign n2431 = ~n2423 & n2430;
  assign n2432 = ~n2414 & ~n2420;
  assign n2433 = ~n2431 & ~n2432;
  assign n2434 = n2423 & n2430;
  assign n2435 = ~n2423 & ~n2430;
  assign n2436 = ~n2434 & ~n2435;
  assign n2437 = n2398 & n2405;
  assign n2438 = ~n2398 & ~n2405;
  assign n2439 = ~n2437 & ~n2438;
  assign n2440 = ~n2408 & ~n2439;
  assign n2441 = ~n2433 & ~n2436;
  assign n2442 = ~n2426 & n2429;
  assign n2443 = n2426 & ~n2429;
  assign n2444 = ~n2442 & ~n2443;
  assign n2445 = ~n2401 & n2404;
  assign n2446 = n2401 & ~n2404;
  assign n2447 = ~n2445 & ~n2446;
  assign n2448 = ~n2444 & ~n2447;
  assign n2449 = ~n2440 & n2448;
  assign n2450 = ~n2441 & n2449;
  assign n2451 = n2436 & ~n2450;
  assign n2452 = ~n2436 & n2450;
  assign n2453 = ~n2451 & ~n2452;
  assign n2454 = n2439 & n2453;
  assign n2455 = ~n2451 & ~n2454;
  assign n2456 = n2433 & ~n2455;
  assign n2457 = ~n2408 & ~n2456;
  assign n2458 = ~n2433 & n2455;
  assign n2459 = ~n2457 & ~n2458;
  assign n2460 = n2383 & n2459;
  assign n2461 = ~n2408 & n2433;
  assign n2462 = n2408 & ~n2433;
  assign n2463 = ~n2461 & ~n2462;
  assign n2464 = n2455 & ~n2463;
  assign n2465 = ~n2455 & n2463;
  assign n2466 = ~n2464 & ~n2465;
  assign n2467 = ~n2332 & n2357;
  assign n2468 = n2332 & ~n2357;
  assign n2469 = ~n2467 & ~n2468;
  assign n2470 = n2379 & ~n2469;
  assign n2471 = ~n2379 & n2469;
  assign n2472 = ~n2470 & ~n2471;
  assign n2473 = n2466 & n2472;
  assign n2474 = n2368 & ~n2371;
  assign n2475 = ~n2368 & n2371;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = n2444 & ~n2447;
  assign n2478 = ~n2444 & n2447;
  assign n2479 = ~n2477 & ~n2478;
  assign n2480 = ~n2476 & ~n2479;
  assign n2481 = ~n2363 & ~n2377;
  assign n2482 = ~n2378 & ~n2481;
  assign n2483 = ~n2480 & n2482;
  assign n2484 = ~n2439 & ~n2453;
  assign n2485 = ~n2454 & ~n2484;
  assign n2486 = ~n2480 & ~n2482;
  assign n2487 = n2482 & ~n2483;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = n2485 & ~n2488;
  assign n2490 = ~n2483 & ~n2489;
  assign n2491 = ~n2466 & ~n2472;
  assign n2492 = ~n2473 & ~n2491;
  assign n2493 = n2490 & n2492;
  assign n2494 = ~n2473 & ~n2493;
  assign n2495 = ~n2460 & ~n2494;
  assign n2496 = ~n2383 & ~n2459;
  assign n2497 = ~n2495 & ~n2496;
  assign n2498 = pi910  & pi911 ;
  assign n2499 = ~pi910  & pi911 ;
  assign n2500 = pi910  & ~pi911 ;
  assign n2501 = ~n2499 & ~n2500;
  assign n2502 = pi912  & ~n2501;
  assign n2503 = ~n2498 & ~n2502;
  assign n2504 = pi907  & pi908 ;
  assign n2505 = ~pi907  & pi908 ;
  assign n2506 = pi907  & ~pi908 ;
  assign n2507 = ~n2505 & ~n2506;
  assign n2508 = pi909  & ~n2507;
  assign n2509 = ~n2504 & ~n2508;
  assign n2510 = ~n2503 & n2509;
  assign n2511 = n2503 & ~n2509;
  assign n2512 = ~n2510 & ~n2511;
  assign n2513 = ~pi909  & ~n2507;
  assign n2514 = pi909  & n2507;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = ~pi912  & ~n2501;
  assign n2517 = pi912  & n2501;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = ~n2515 & ~n2518;
  assign n2520 = ~n2512 & n2519;
  assign n2521 = ~n2503 & ~n2509;
  assign n2522 = ~n2520 & ~n2521;
  assign n2523 = pi916  & pi917 ;
  assign n2524 = ~pi916  & pi917 ;
  assign n2525 = pi916  & ~pi917 ;
  assign n2526 = ~n2524 & ~n2525;
  assign n2527 = pi918  & ~n2526;
  assign n2528 = ~n2523 & ~n2527;
  assign n2529 = pi913  & pi914 ;
  assign n2530 = ~pi913  & pi914 ;
  assign n2531 = pi913  & ~pi914 ;
  assign n2532 = ~n2530 & ~n2531;
  assign n2533 = pi915  & ~n2532;
  assign n2534 = ~n2529 & ~n2533;
  assign n2535 = ~n2528 & n2534;
  assign n2536 = n2528 & ~n2534;
  assign n2537 = ~n2535 & ~n2536;
  assign n2538 = ~pi915  & ~n2532;
  assign n2539 = pi915  & n2532;
  assign n2540 = ~n2538 & ~n2539;
  assign n2541 = ~pi918  & ~n2526;
  assign n2542 = pi918  & n2526;
  assign n2543 = ~n2541 & ~n2542;
  assign n2544 = ~n2540 & ~n2543;
  assign n2545 = ~n2537 & n2544;
  assign n2546 = ~n2528 & ~n2534;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = n2537 & n2544;
  assign n2549 = ~n2537 & ~n2544;
  assign n2550 = ~n2548 & ~n2549;
  assign n2551 = n2512 & n2519;
  assign n2552 = ~n2512 & ~n2519;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = ~n2522 & ~n2553;
  assign n2555 = ~n2547 & ~n2550;
  assign n2556 = ~n2540 & n2543;
  assign n2557 = n2540 & ~n2543;
  assign n2558 = ~n2556 & ~n2557;
  assign n2559 = ~n2515 & n2518;
  assign n2560 = n2515 & ~n2518;
  assign n2561 = ~n2559 & ~n2560;
  assign n2562 = ~n2558 & ~n2561;
  assign n2563 = ~n2554 & n2562;
  assign n2564 = ~n2555 & n2563;
  assign n2565 = n2550 & ~n2564;
  assign n2566 = ~n2550 & n2564;
  assign n2567 = ~n2565 & ~n2566;
  assign n2568 = n2553 & n2567;
  assign n2569 = ~n2565 & ~n2568;
  assign n2570 = n2547 & ~n2569;
  assign n2571 = ~n2522 & ~n2570;
  assign n2572 = ~n2547 & n2569;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = pi898  & pi899 ;
  assign n2575 = ~pi898  & pi899 ;
  assign n2576 = pi898  & ~pi899 ;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = pi900  & ~n2577;
  assign n2579 = ~n2574 & ~n2578;
  assign n2580 = pi895  & pi896 ;
  assign n2581 = ~pi895  & pi896 ;
  assign n2582 = pi895  & ~pi896 ;
  assign n2583 = ~n2581 & ~n2582;
  assign n2584 = pi897  & ~n2583;
  assign n2585 = ~n2580 & ~n2584;
  assign n2586 = ~n2579 & n2585;
  assign n2587 = n2579 & ~n2585;
  assign n2588 = ~n2586 & ~n2587;
  assign n2589 = ~pi897  & ~n2583;
  assign n2590 = pi897  & n2583;
  assign n2591 = ~n2589 & ~n2590;
  assign n2592 = ~pi900  & ~n2577;
  assign n2593 = pi900  & n2577;
  assign n2594 = ~n2592 & ~n2593;
  assign n2595 = ~n2591 & ~n2594;
  assign n2596 = ~n2588 & n2595;
  assign n2597 = ~n2579 & ~n2585;
  assign n2598 = ~n2596 & ~n2597;
  assign n2599 = pi904  & pi905 ;
  assign n2600 = ~pi904  & pi905 ;
  assign n2601 = pi904  & ~pi905 ;
  assign n2602 = ~n2600 & ~n2601;
  assign n2603 = pi906  & ~n2602;
  assign n2604 = ~n2599 & ~n2603;
  assign n2605 = pi901  & pi902 ;
  assign n2606 = ~pi901  & pi902 ;
  assign n2607 = pi901  & ~pi902 ;
  assign n2608 = ~n2606 & ~n2607;
  assign n2609 = pi903  & ~n2608;
  assign n2610 = ~n2605 & ~n2609;
  assign n2611 = ~n2604 & n2610;
  assign n2612 = n2604 & ~n2610;
  assign n2613 = ~n2611 & ~n2612;
  assign n2614 = ~pi903  & ~n2608;
  assign n2615 = pi903  & n2608;
  assign n2616 = ~n2614 & ~n2615;
  assign n2617 = ~pi906  & ~n2602;
  assign n2618 = pi906  & n2602;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = ~n2616 & ~n2619;
  assign n2621 = ~n2613 & n2620;
  assign n2622 = ~n2604 & ~n2610;
  assign n2623 = ~n2621 & ~n2622;
  assign n2624 = n2613 & n2620;
  assign n2625 = ~n2613 & ~n2620;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = n2588 & n2595;
  assign n2628 = ~n2588 & ~n2595;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = ~n2598 & ~n2629;
  assign n2631 = ~n2623 & ~n2626;
  assign n2632 = ~n2616 & n2619;
  assign n2633 = n2616 & ~n2619;
  assign n2634 = ~n2632 & ~n2633;
  assign n2635 = ~n2591 & n2594;
  assign n2636 = n2591 & ~n2594;
  assign n2637 = ~n2635 & ~n2636;
  assign n2638 = ~n2634 & ~n2637;
  assign n2639 = ~n2630 & n2638;
  assign n2640 = ~n2631 & n2639;
  assign n2641 = n2626 & ~n2640;
  assign n2642 = ~n2626 & n2640;
  assign n2643 = ~n2641 & ~n2642;
  assign n2644 = n2629 & n2643;
  assign n2645 = ~n2641 & ~n2644;
  assign n2646 = n2623 & ~n2645;
  assign n2647 = ~n2598 & ~n2646;
  assign n2648 = ~n2623 & n2645;
  assign n2649 = ~n2647 & ~n2648;
  assign n2650 = n2573 & n2649;
  assign n2651 = ~n2598 & n2623;
  assign n2652 = n2598 & ~n2623;
  assign n2653 = ~n2651 & ~n2652;
  assign n2654 = n2645 & ~n2653;
  assign n2655 = ~n2645 & n2653;
  assign n2656 = ~n2654 & ~n2655;
  assign n2657 = ~n2522 & n2547;
  assign n2658 = n2522 & ~n2547;
  assign n2659 = ~n2657 & ~n2658;
  assign n2660 = n2569 & ~n2659;
  assign n2661 = ~n2569 & n2659;
  assign n2662 = ~n2660 & ~n2661;
  assign n2663 = n2656 & n2662;
  assign n2664 = n2558 & ~n2561;
  assign n2665 = ~n2558 & n2561;
  assign n2666 = ~n2664 & ~n2665;
  assign n2667 = n2634 & ~n2637;
  assign n2668 = ~n2634 & n2637;
  assign n2669 = ~n2667 & ~n2668;
  assign n2670 = ~n2666 & ~n2669;
  assign n2671 = ~n2553 & ~n2567;
  assign n2672 = ~n2568 & ~n2671;
  assign n2673 = ~n2670 & n2672;
  assign n2674 = ~n2629 & ~n2643;
  assign n2675 = ~n2644 & ~n2674;
  assign n2676 = n2670 & ~n2672;
  assign n2677 = ~n2673 & ~n2676;
  assign n2678 = n2675 & n2677;
  assign n2679 = ~n2673 & ~n2678;
  assign n2680 = ~n2656 & ~n2662;
  assign n2681 = ~n2663 & ~n2680;
  assign n2682 = n2679 & n2681;
  assign n2683 = ~n2663 & ~n2682;
  assign n2684 = ~n2650 & ~n2683;
  assign n2685 = ~n2573 & ~n2649;
  assign n2686 = ~n2684 & ~n2685;
  assign n2687 = ~n2497 & ~n2686;
  assign n2688 = n2497 & n2686;
  assign n2689 = ~n2687 & ~n2688;
  assign n2690 = ~n2460 & ~n2496;
  assign n2691 = ~n2494 & n2690;
  assign n2692 = n2494 & ~n2690;
  assign n2693 = ~n2691 & ~n2692;
  assign n2694 = ~n2650 & ~n2685;
  assign n2695 = ~n2683 & n2694;
  assign n2696 = n2683 & ~n2694;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = n2693 & n2697;
  assign n2699 = ~n2679 & ~n2681;
  assign n2700 = ~n2682 & ~n2699;
  assign n2701 = ~n2490 & ~n2492;
  assign n2702 = ~n2493 & ~n2701;
  assign n2703 = n2700 & n2702;
  assign n2704 = ~n2700 & ~n2702;
  assign n2705 = ~n2703 & ~n2704;
  assign n2706 = ~n2476 & n2479;
  assign n2707 = n2476 & ~n2479;
  assign n2708 = ~n2706 & ~n2707;
  assign n2709 = ~n2666 & n2669;
  assign n2710 = n2666 & ~n2669;
  assign n2711 = ~n2709 & ~n2710;
  assign n2712 = ~n2708 & ~n2711;
  assign n2713 = ~n2485 & n2488;
  assign n2714 = ~n2489 & ~n2713;
  assign n2715 = ~n2712 & n2714;
  assign n2716 = ~n2675 & ~n2677;
  assign n2717 = ~n2678 & ~n2716;
  assign n2718 = n2712 & ~n2714;
  assign n2719 = ~n2715 & ~n2718;
  assign n2720 = n2717 & n2719;
  assign n2721 = ~n2715 & ~n2720;
  assign n2722 = n2705 & n2721;
  assign n2723 = ~n2703 & ~n2722;
  assign n2724 = ~n2693 & ~n2697;
  assign n2725 = ~n2698 & ~n2724;
  assign n2726 = ~n2723 & n2725;
  assign n2727 = ~n2698 & ~n2726;
  assign n2728 = n2689 & ~n2727;
  assign n2729 = ~n2687 & ~n2728;
  assign n2730 = pi886  & pi887 ;
  assign n2731 = ~pi886  & pi887 ;
  assign n2732 = pi886  & ~pi887 ;
  assign n2733 = ~n2731 & ~n2732;
  assign n2734 = pi888  & ~n2733;
  assign n2735 = ~n2730 & ~n2734;
  assign n2736 = pi883  & pi884 ;
  assign n2737 = ~pi883  & pi884 ;
  assign n2738 = pi883  & ~pi884 ;
  assign n2739 = ~n2737 & ~n2738;
  assign n2740 = pi885  & ~n2739;
  assign n2741 = ~n2736 & ~n2740;
  assign n2742 = ~n2735 & n2741;
  assign n2743 = n2735 & ~n2741;
  assign n2744 = ~n2742 & ~n2743;
  assign n2745 = ~pi885  & ~n2739;
  assign n2746 = pi885  & n2739;
  assign n2747 = ~n2745 & ~n2746;
  assign n2748 = ~pi888  & ~n2733;
  assign n2749 = pi888  & n2733;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = ~n2747 & ~n2750;
  assign n2752 = ~n2744 & n2751;
  assign n2753 = ~n2735 & ~n2741;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = pi892  & pi893 ;
  assign n2756 = ~pi892  & pi893 ;
  assign n2757 = pi892  & ~pi893 ;
  assign n2758 = ~n2756 & ~n2757;
  assign n2759 = pi894  & ~n2758;
  assign n2760 = ~n2755 & ~n2759;
  assign n2761 = pi889  & pi890 ;
  assign n2762 = ~pi889  & pi890 ;
  assign n2763 = pi889  & ~pi890 ;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = pi891  & ~n2764;
  assign n2766 = ~n2761 & ~n2765;
  assign n2767 = ~n2760 & n2766;
  assign n2768 = n2760 & ~n2766;
  assign n2769 = ~n2767 & ~n2768;
  assign n2770 = ~pi891  & ~n2764;
  assign n2771 = pi891  & n2764;
  assign n2772 = ~n2770 & ~n2771;
  assign n2773 = ~pi894  & ~n2758;
  assign n2774 = pi894  & n2758;
  assign n2775 = ~n2773 & ~n2774;
  assign n2776 = ~n2772 & ~n2775;
  assign n2777 = ~n2769 & n2776;
  assign n2778 = ~n2760 & ~n2766;
  assign n2779 = ~n2777 & ~n2778;
  assign n2780 = n2769 & n2776;
  assign n2781 = ~n2769 & ~n2776;
  assign n2782 = ~n2780 & ~n2781;
  assign n2783 = n2744 & n2751;
  assign n2784 = ~n2744 & ~n2751;
  assign n2785 = ~n2783 & ~n2784;
  assign n2786 = ~n2754 & ~n2785;
  assign n2787 = ~n2779 & ~n2782;
  assign n2788 = ~n2772 & n2775;
  assign n2789 = n2772 & ~n2775;
  assign n2790 = ~n2788 & ~n2789;
  assign n2791 = ~n2747 & n2750;
  assign n2792 = n2747 & ~n2750;
  assign n2793 = ~n2791 & ~n2792;
  assign n2794 = ~n2790 & ~n2793;
  assign n2795 = ~n2786 & n2794;
  assign n2796 = ~n2787 & n2795;
  assign n2797 = n2782 & ~n2796;
  assign n2798 = ~n2782 & n2796;
  assign n2799 = ~n2797 & ~n2798;
  assign n2800 = n2785 & n2799;
  assign n2801 = ~n2797 & ~n2800;
  assign n2802 = n2779 & ~n2801;
  assign n2803 = ~n2754 & ~n2802;
  assign n2804 = ~n2779 & n2801;
  assign n2805 = ~n2803 & ~n2804;
  assign n2806 = pi874  & pi875 ;
  assign n2807 = ~pi874  & pi875 ;
  assign n2808 = pi874  & ~pi875 ;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = pi876  & ~n2809;
  assign n2811 = ~n2806 & ~n2810;
  assign n2812 = pi871  & pi872 ;
  assign n2813 = ~pi871  & pi872 ;
  assign n2814 = pi871  & ~pi872 ;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = pi873  & ~n2815;
  assign n2817 = ~n2812 & ~n2816;
  assign n2818 = ~n2811 & n2817;
  assign n2819 = n2811 & ~n2817;
  assign n2820 = ~n2818 & ~n2819;
  assign n2821 = ~pi873  & ~n2815;
  assign n2822 = pi873  & n2815;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = ~pi876  & ~n2809;
  assign n2825 = pi876  & n2809;
  assign n2826 = ~n2824 & ~n2825;
  assign n2827 = ~n2823 & ~n2826;
  assign n2828 = ~n2820 & n2827;
  assign n2829 = ~n2811 & ~n2817;
  assign n2830 = ~n2828 & ~n2829;
  assign n2831 = pi880  & pi881 ;
  assign n2832 = ~pi880  & pi881 ;
  assign n2833 = pi880  & ~pi881 ;
  assign n2834 = ~n2832 & ~n2833;
  assign n2835 = pi882  & ~n2834;
  assign n2836 = ~n2831 & ~n2835;
  assign n2837 = pi877  & pi878 ;
  assign n2838 = ~pi877  & pi878 ;
  assign n2839 = pi877  & ~pi878 ;
  assign n2840 = ~n2838 & ~n2839;
  assign n2841 = pi879  & ~n2840;
  assign n2842 = ~n2837 & ~n2841;
  assign n2843 = ~n2836 & n2842;
  assign n2844 = n2836 & ~n2842;
  assign n2845 = ~n2843 & ~n2844;
  assign n2846 = ~pi879  & ~n2840;
  assign n2847 = pi879  & n2840;
  assign n2848 = ~n2846 & ~n2847;
  assign n2849 = ~pi882  & ~n2834;
  assign n2850 = pi882  & n2834;
  assign n2851 = ~n2849 & ~n2850;
  assign n2852 = ~n2848 & ~n2851;
  assign n2853 = ~n2845 & n2852;
  assign n2854 = ~n2836 & ~n2842;
  assign n2855 = ~n2853 & ~n2854;
  assign n2856 = n2845 & n2852;
  assign n2857 = ~n2845 & ~n2852;
  assign n2858 = ~n2856 & ~n2857;
  assign n2859 = n2820 & n2827;
  assign n2860 = ~n2820 & ~n2827;
  assign n2861 = ~n2859 & ~n2860;
  assign n2862 = ~n2830 & ~n2861;
  assign n2863 = ~n2855 & ~n2858;
  assign n2864 = ~n2848 & n2851;
  assign n2865 = n2848 & ~n2851;
  assign n2866 = ~n2864 & ~n2865;
  assign n2867 = ~n2823 & n2826;
  assign n2868 = n2823 & ~n2826;
  assign n2869 = ~n2867 & ~n2868;
  assign n2870 = ~n2866 & ~n2869;
  assign n2871 = ~n2862 & n2870;
  assign n2872 = ~n2863 & n2871;
  assign n2873 = n2858 & ~n2872;
  assign n2874 = ~n2858 & n2872;
  assign n2875 = ~n2873 & ~n2874;
  assign n2876 = n2861 & n2875;
  assign n2877 = ~n2873 & ~n2876;
  assign n2878 = n2855 & ~n2877;
  assign n2879 = ~n2830 & ~n2878;
  assign n2880 = ~n2855 & n2877;
  assign n2881 = ~n2879 & ~n2880;
  assign n2882 = n2805 & n2881;
  assign n2883 = ~n2830 & n2855;
  assign n2884 = n2830 & ~n2855;
  assign n2885 = ~n2883 & ~n2884;
  assign n2886 = n2877 & ~n2885;
  assign n2887 = ~n2877 & n2885;
  assign n2888 = ~n2886 & ~n2887;
  assign n2889 = ~n2754 & n2779;
  assign n2890 = n2754 & ~n2779;
  assign n2891 = ~n2889 & ~n2890;
  assign n2892 = n2801 & ~n2891;
  assign n2893 = ~n2801 & n2891;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = n2888 & n2894;
  assign n2896 = n2790 & ~n2793;
  assign n2897 = ~n2790 & n2793;
  assign n2898 = ~n2896 & ~n2897;
  assign n2899 = n2866 & ~n2869;
  assign n2900 = ~n2866 & n2869;
  assign n2901 = ~n2899 & ~n2900;
  assign n2902 = ~n2898 & ~n2901;
  assign n2903 = ~n2785 & ~n2799;
  assign n2904 = ~n2800 & ~n2903;
  assign n2905 = ~n2902 & n2904;
  assign n2906 = ~n2861 & ~n2875;
  assign n2907 = ~n2876 & ~n2906;
  assign n2908 = ~n2902 & ~n2904;
  assign n2909 = n2904 & ~n2905;
  assign n2910 = ~n2908 & ~n2909;
  assign n2911 = n2907 & ~n2910;
  assign n2912 = ~n2905 & ~n2911;
  assign n2913 = ~n2888 & ~n2894;
  assign n2914 = ~n2895 & ~n2913;
  assign n2915 = n2912 & n2914;
  assign n2916 = ~n2895 & ~n2915;
  assign n2917 = ~n2882 & ~n2916;
  assign n2918 = ~n2805 & ~n2881;
  assign n2919 = ~n2917 & ~n2918;
  assign n2920 = pi862  & pi863 ;
  assign n2921 = ~pi862  & pi863 ;
  assign n2922 = pi862  & ~pi863 ;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = pi864  & ~n2923;
  assign n2925 = ~n2920 & ~n2924;
  assign n2926 = pi859  & pi860 ;
  assign n2927 = ~pi859  & pi860 ;
  assign n2928 = pi859  & ~pi860 ;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = pi861  & ~n2929;
  assign n2931 = ~n2926 & ~n2930;
  assign n2932 = ~n2925 & n2931;
  assign n2933 = n2925 & ~n2931;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = ~pi861  & ~n2929;
  assign n2936 = pi861  & n2929;
  assign n2937 = ~n2935 & ~n2936;
  assign n2938 = ~pi864  & ~n2923;
  assign n2939 = pi864  & n2923;
  assign n2940 = ~n2938 & ~n2939;
  assign n2941 = ~n2937 & ~n2940;
  assign n2942 = ~n2934 & n2941;
  assign n2943 = ~n2925 & ~n2931;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = pi868  & pi869 ;
  assign n2946 = ~pi868  & pi869 ;
  assign n2947 = pi868  & ~pi869 ;
  assign n2948 = ~n2946 & ~n2947;
  assign n2949 = pi870  & ~n2948;
  assign n2950 = ~n2945 & ~n2949;
  assign n2951 = pi865  & pi866 ;
  assign n2952 = ~pi865  & pi866 ;
  assign n2953 = pi865  & ~pi866 ;
  assign n2954 = ~n2952 & ~n2953;
  assign n2955 = pi867  & ~n2954;
  assign n2956 = ~n2951 & ~n2955;
  assign n2957 = ~n2950 & n2956;
  assign n2958 = n2950 & ~n2956;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = ~pi867  & ~n2954;
  assign n2961 = pi867  & n2954;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = ~pi870  & ~n2948;
  assign n2964 = pi870  & n2948;
  assign n2965 = ~n2963 & ~n2964;
  assign n2966 = ~n2962 & ~n2965;
  assign n2967 = ~n2959 & n2966;
  assign n2968 = ~n2950 & ~n2956;
  assign n2969 = ~n2967 & ~n2968;
  assign n2970 = n2959 & n2966;
  assign n2971 = ~n2959 & ~n2966;
  assign n2972 = ~n2970 & ~n2971;
  assign n2973 = n2934 & n2941;
  assign n2974 = ~n2934 & ~n2941;
  assign n2975 = ~n2973 & ~n2974;
  assign n2976 = ~n2944 & ~n2975;
  assign n2977 = ~n2969 & ~n2972;
  assign n2978 = ~n2962 & n2965;
  assign n2979 = n2962 & ~n2965;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = ~n2937 & n2940;
  assign n2982 = n2937 & ~n2940;
  assign n2983 = ~n2981 & ~n2982;
  assign n2984 = ~n2980 & ~n2983;
  assign n2985 = ~n2976 & n2984;
  assign n2986 = ~n2977 & n2985;
  assign n2987 = n2972 & ~n2986;
  assign n2988 = ~n2972 & n2986;
  assign n2989 = ~n2987 & ~n2988;
  assign n2990 = n2975 & n2989;
  assign n2991 = ~n2987 & ~n2990;
  assign n2992 = n2969 & ~n2991;
  assign n2993 = ~n2944 & ~n2992;
  assign n2994 = ~n2969 & n2991;
  assign n2995 = ~n2993 & ~n2994;
  assign n2996 = pi850  & pi851 ;
  assign n2997 = ~pi850  & pi851 ;
  assign n2998 = pi850  & ~pi851 ;
  assign n2999 = ~n2997 & ~n2998;
  assign n3000 = pi852  & ~n2999;
  assign n3001 = ~n2996 & ~n3000;
  assign n3002 = pi847  & pi848 ;
  assign n3003 = ~pi847  & pi848 ;
  assign n3004 = pi847  & ~pi848 ;
  assign n3005 = ~n3003 & ~n3004;
  assign n3006 = pi849  & ~n3005;
  assign n3007 = ~n3002 & ~n3006;
  assign n3008 = ~n3001 & n3007;
  assign n3009 = n3001 & ~n3007;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = ~pi849  & ~n3005;
  assign n3012 = pi849  & n3005;
  assign n3013 = ~n3011 & ~n3012;
  assign n3014 = ~pi852  & ~n2999;
  assign n3015 = pi852  & n2999;
  assign n3016 = ~n3014 & ~n3015;
  assign n3017 = ~n3013 & ~n3016;
  assign n3018 = ~n3010 & n3017;
  assign n3019 = ~n3001 & ~n3007;
  assign n3020 = ~n3018 & ~n3019;
  assign n3021 = pi856  & pi857 ;
  assign n3022 = ~pi856  & pi857 ;
  assign n3023 = pi856  & ~pi857 ;
  assign n3024 = ~n3022 & ~n3023;
  assign n3025 = pi858  & ~n3024;
  assign n3026 = ~n3021 & ~n3025;
  assign n3027 = pi853  & pi854 ;
  assign n3028 = ~pi853  & pi854 ;
  assign n3029 = pi853  & ~pi854 ;
  assign n3030 = ~n3028 & ~n3029;
  assign n3031 = pi855  & ~n3030;
  assign n3032 = ~n3027 & ~n3031;
  assign n3033 = ~n3026 & n3032;
  assign n3034 = n3026 & ~n3032;
  assign n3035 = ~n3033 & ~n3034;
  assign n3036 = ~pi855  & ~n3030;
  assign n3037 = pi855  & n3030;
  assign n3038 = ~n3036 & ~n3037;
  assign n3039 = ~pi858  & ~n3024;
  assign n3040 = pi858  & n3024;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042 = ~n3038 & ~n3041;
  assign n3043 = ~n3035 & n3042;
  assign n3044 = ~n3026 & ~n3032;
  assign n3045 = ~n3043 & ~n3044;
  assign n3046 = n3035 & n3042;
  assign n3047 = ~n3035 & ~n3042;
  assign n3048 = ~n3046 & ~n3047;
  assign n3049 = n3010 & n3017;
  assign n3050 = ~n3010 & ~n3017;
  assign n3051 = ~n3049 & ~n3050;
  assign n3052 = ~n3020 & ~n3051;
  assign n3053 = ~n3045 & ~n3048;
  assign n3054 = ~n3038 & n3041;
  assign n3055 = n3038 & ~n3041;
  assign n3056 = ~n3054 & ~n3055;
  assign n3057 = ~n3013 & n3016;
  assign n3058 = n3013 & ~n3016;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = ~n3056 & ~n3059;
  assign n3061 = ~n3052 & n3060;
  assign n3062 = ~n3053 & n3061;
  assign n3063 = n3048 & ~n3062;
  assign n3064 = ~n3048 & n3062;
  assign n3065 = ~n3063 & ~n3064;
  assign n3066 = n3051 & n3065;
  assign n3067 = ~n3063 & ~n3066;
  assign n3068 = n3045 & ~n3067;
  assign n3069 = ~n3020 & ~n3068;
  assign n3070 = ~n3045 & n3067;
  assign n3071 = ~n3069 & ~n3070;
  assign n3072 = n2995 & n3071;
  assign n3073 = ~n3020 & n3045;
  assign n3074 = n3020 & ~n3045;
  assign n3075 = ~n3073 & ~n3074;
  assign n3076 = n3067 & ~n3075;
  assign n3077 = ~n3067 & n3075;
  assign n3078 = ~n3076 & ~n3077;
  assign n3079 = ~n2944 & n2969;
  assign n3080 = n2944 & ~n2969;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = n2991 & ~n3081;
  assign n3083 = ~n2991 & n3081;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = n3078 & n3084;
  assign n3086 = n2980 & ~n2983;
  assign n3087 = ~n2980 & n2983;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = n3056 & ~n3059;
  assign n3090 = ~n3056 & n3059;
  assign n3091 = ~n3089 & ~n3090;
  assign n3092 = ~n3088 & ~n3091;
  assign n3093 = ~n2975 & ~n2989;
  assign n3094 = ~n2990 & ~n3093;
  assign n3095 = ~n3092 & n3094;
  assign n3096 = ~n3051 & ~n3065;
  assign n3097 = ~n3066 & ~n3096;
  assign n3098 = n3092 & ~n3094;
  assign n3099 = ~n3095 & ~n3098;
  assign n3100 = n3097 & n3099;
  assign n3101 = ~n3095 & ~n3100;
  assign n3102 = ~n3078 & ~n3084;
  assign n3103 = ~n3085 & ~n3102;
  assign n3104 = n3101 & n3103;
  assign n3105 = ~n3085 & ~n3104;
  assign n3106 = ~n3072 & ~n3105;
  assign n3107 = ~n2995 & ~n3071;
  assign n3108 = ~n3106 & ~n3107;
  assign n3109 = ~n2919 & ~n3108;
  assign n3110 = n2919 & n3108;
  assign n3111 = ~n3109 & ~n3110;
  assign n3112 = ~n2882 & ~n2918;
  assign n3113 = ~n2916 & n3112;
  assign n3114 = n2916 & ~n3112;
  assign n3115 = ~n3113 & ~n3114;
  assign n3116 = ~n3072 & ~n3107;
  assign n3117 = ~n3105 & n3116;
  assign n3118 = n3105 & ~n3116;
  assign n3119 = ~n3117 & ~n3118;
  assign n3120 = n3115 & n3119;
  assign n3121 = ~n3101 & ~n3103;
  assign n3122 = ~n3104 & ~n3121;
  assign n3123 = ~n2912 & ~n2914;
  assign n3124 = ~n2915 & ~n3123;
  assign n3125 = n3122 & n3124;
  assign n3126 = ~n3122 & ~n3124;
  assign n3127 = ~n3125 & ~n3126;
  assign n3128 = ~n2898 & n2901;
  assign n3129 = n2898 & ~n2901;
  assign n3130 = ~n3128 & ~n3129;
  assign n3131 = ~n3088 & n3091;
  assign n3132 = n3088 & ~n3091;
  assign n3133 = ~n3131 & ~n3132;
  assign n3134 = ~n3130 & ~n3133;
  assign n3135 = ~n2907 & n2910;
  assign n3136 = ~n2911 & ~n3135;
  assign n3137 = ~n3134 & n3136;
  assign n3138 = ~n3097 & ~n3099;
  assign n3139 = ~n3100 & ~n3138;
  assign n3140 = n3134 & ~n3136;
  assign n3141 = ~n3137 & ~n3140;
  assign n3142 = n3139 & n3141;
  assign n3143 = ~n3137 & ~n3142;
  assign n3144 = n3127 & n3143;
  assign n3145 = ~n3125 & ~n3144;
  assign n3146 = ~n3115 & ~n3119;
  assign n3147 = ~n3120 & ~n3146;
  assign n3148 = ~n3145 & n3147;
  assign n3149 = ~n3120 & ~n3148;
  assign n3150 = n3111 & ~n3149;
  assign n3151 = ~n3109 & ~n3150;
  assign n3152 = ~n2729 & ~n3151;
  assign n3153 = n2729 & n3151;
  assign n3154 = ~n3152 & ~n3153;
  assign n3155 = ~n3111 & n3149;
  assign n3156 = ~n3150 & ~n3155;
  assign n3157 = ~n2689 & n2727;
  assign n3158 = ~n2728 & ~n3157;
  assign n3159 = n3156 & n3158;
  assign n3160 = n2723 & ~n2725;
  assign n3161 = ~n2726 & ~n3160;
  assign n3162 = n3145 & ~n3147;
  assign n3163 = ~n3148 & ~n3162;
  assign n3164 = n3161 & n3163;
  assign n3165 = ~n3161 & ~n3163;
  assign n3166 = ~n3164 & ~n3165;
  assign n3167 = ~n3127 & ~n3143;
  assign n3168 = ~n3144 & ~n3167;
  assign n3169 = ~n2705 & ~n2721;
  assign n3170 = ~n2722 & ~n3169;
  assign n3171 = n3168 & n3170;
  assign n3172 = ~n2708 & n2711;
  assign n3173 = n2708 & ~n2711;
  assign n3174 = ~n3172 & ~n3173;
  assign n3175 = ~n3130 & n3133;
  assign n3176 = n3130 & ~n3133;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = ~n3174 & ~n3177;
  assign n3179 = ~n2717 & ~n2719;
  assign n3180 = ~n2720 & ~n3179;
  assign n3181 = ~n3178 & n3180;
  assign n3182 = ~n3139 & ~n3141;
  assign n3183 = ~n3142 & ~n3182;
  assign n3184 = n3178 & ~n3180;
  assign n3185 = ~n3181 & ~n3184;
  assign n3186 = n3183 & n3185;
  assign n3187 = ~n3181 & ~n3186;
  assign n3188 = ~n3168 & ~n3170;
  assign n3189 = ~n3171 & ~n3188;
  assign n3190 = n3187 & n3189;
  assign n3191 = ~n3171 & ~n3190;
  assign n3192 = n3166 & ~n3191;
  assign n3193 = ~n3164 & ~n3192;
  assign n3194 = ~n3156 & ~n3158;
  assign n3195 = ~n3159 & ~n3194;
  assign n3196 = ~n3193 & n3195;
  assign n3197 = ~n3159 & ~n3196;
  assign n3198 = n3154 & ~n3197;
  assign n3199 = ~n3152 & ~n3198;
  assign n3200 = ~n2307 & ~n3199;
  assign n3201 = n2298 & ~n2300;
  assign n3202 = ~n2301 & ~n3201;
  assign n3203 = ~n3154 & n3197;
  assign n3204 = ~n3198 & ~n3203;
  assign n3205 = n3202 & n3204;
  assign n3206 = n3193 & ~n3195;
  assign n3207 = ~n3196 & ~n3206;
  assign n3208 = n2294 & ~n2296;
  assign n3209 = ~n2297 & ~n3208;
  assign n3210 = n3207 & n3209;
  assign n3211 = ~n3187 & ~n3189;
  assign n3212 = ~n3190 & ~n3211;
  assign n3213 = n2279 & ~n2281;
  assign n3214 = ~n2282 & ~n3213;
  assign n3215 = n3212 & n3214;
  assign n3216 = ~n2265 & n2268;
  assign n3217 = n2265 & ~n2268;
  assign n3218 = ~n3216 & ~n3217;
  assign n3219 = ~n3174 & n3177;
  assign n3220 = n3174 & ~n3177;
  assign n3221 = ~n3219 & ~n3220;
  assign n3222 = ~n3218 & ~n3221;
  assign n3223 = ~n2274 & ~n2277;
  assign n3224 = n2276 & n3223;
  assign n3225 = ~n2276 & ~n3223;
  assign n3226 = ~n3224 & ~n3225;
  assign n3227 = n3222 & ~n3226;
  assign n3228 = ~n3183 & ~n3185;
  assign n3229 = ~n3186 & ~n3228;
  assign n3230 = ~n3222 & n3226;
  assign n3231 = ~n3229 & ~n3230;
  assign n3232 = ~n3227 & ~n3231;
  assign n3233 = ~n3212 & ~n3214;
  assign n3234 = ~n3215 & ~n3233;
  assign n3235 = ~n3232 & n3234;
  assign n3236 = ~n3215 & ~n3235;
  assign n3237 = ~n2290 & ~n2293;
  assign n3238 = ~n2283 & n3237;
  assign n3239 = n2283 & ~n3237;
  assign n3240 = ~n3238 & ~n3239;
  assign n3241 = ~n3166 & n3191;
  assign n3242 = ~n3192 & ~n3241;
  assign n3243 = ~n3240 & ~n3242;
  assign n3244 = ~n3236 & ~n3243;
  assign n3245 = n3240 & n3242;
  assign n3246 = ~n3244 & ~n3245;
  assign n3247 = ~n3207 & ~n3209;
  assign n3248 = ~n3210 & ~n3247;
  assign n3249 = ~n3246 & n3248;
  assign n3250 = ~n3210 & ~n3249;
  assign n3251 = ~n3202 & ~n3204;
  assign n3252 = ~n3205 & ~n3251;
  assign n3253 = ~n3250 & n3252;
  assign n3254 = ~n3205 & ~n3253;
  assign n3255 = n2307 & n3199;
  assign n3256 = ~n3200 & ~n3255;
  assign n3257 = ~n3254 & n3256;
  assign n3258 = ~n3200 & ~n3257;
  assign n3259 = n2304 & ~n3258;
  assign n3260 = pi451  & ~pi452 ;
  assign n3261 = ~pi451  & pi452 ;
  assign n3262 = ~n3260 & ~n3261;
  assign n3263 = ~pi453  & ~n3262;
  assign n3264 = pi453  & n3262;
  assign n3265 = ~n3263 & ~n3264;
  assign n3266 = pi454  & ~pi455 ;
  assign n3267 = ~pi454  & pi455 ;
  assign n3268 = ~n3266 & ~n3267;
  assign n3269 = ~pi456  & ~n3268;
  assign n3270 = pi456  & n3268;
  assign n3271 = ~n3269 & ~n3270;
  assign n3272 = ~n3265 & ~n3271;
  assign n3273 = pi454  & pi455 ;
  assign n3274 = pi456  & ~n3268;
  assign n3275 = ~n3273 & ~n3274;
  assign n3276 = pi451  & pi452 ;
  assign n3277 = pi453  & ~n3262;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = n3275 & ~n3278;
  assign n3280 = ~n3275 & n3278;
  assign n3281 = ~n3279 & ~n3280;
  assign n3282 = n3272 & ~n3281;
  assign n3283 = ~n3275 & ~n3278;
  assign n3284 = ~n3282 & ~n3283;
  assign n3285 = pi460  & pi461 ;
  assign n3286 = pi460  & ~pi461 ;
  assign n3287 = ~pi460  & pi461 ;
  assign n3288 = ~n3286 & ~n3287;
  assign n3289 = pi462  & ~n3288;
  assign n3290 = ~n3285 & ~n3289;
  assign n3291 = pi457  & pi458 ;
  assign n3292 = pi457  & ~pi458 ;
  assign n3293 = ~pi457  & pi458 ;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = pi459  & ~n3294;
  assign n3296 = ~n3291 & ~n3295;
  assign n3297 = ~n3290 & n3296;
  assign n3298 = n3290 & ~n3296;
  assign n3299 = ~n3297 & ~n3298;
  assign n3300 = ~pi459  & ~n3294;
  assign n3301 = pi459  & n3294;
  assign n3302 = ~n3300 & ~n3301;
  assign n3303 = ~pi462  & ~n3288;
  assign n3304 = pi462  & n3288;
  assign n3305 = ~n3303 & ~n3304;
  assign n3306 = ~n3302 & ~n3305;
  assign n3307 = ~n3299 & n3306;
  assign n3308 = ~n3290 & ~n3296;
  assign n3309 = ~n3307 & ~n3308;
  assign n3310 = n3272 & n3281;
  assign n3311 = ~n3272 & ~n3281;
  assign n3312 = ~n3310 & ~n3311;
  assign n3313 = n3299 & n3306;
  assign n3314 = ~n3299 & ~n3306;
  assign n3315 = ~n3313 & ~n3314;
  assign n3316 = ~n3309 & ~n3315;
  assign n3317 = ~n3284 & ~n3312;
  assign n3318 = ~n3265 & n3271;
  assign n3319 = n3265 & ~n3271;
  assign n3320 = ~n3318 & ~n3319;
  assign n3321 = ~n3302 & n3305;
  assign n3322 = n3302 & ~n3305;
  assign n3323 = ~n3321 & ~n3322;
  assign n3324 = ~n3320 & ~n3323;
  assign n3325 = ~n3316 & n3324;
  assign n3326 = ~n3317 & n3325;
  assign n3327 = n3315 & ~n3326;
  assign n3328 = ~n3312 & ~n3327;
  assign n3329 = n3315 & n3326;
  assign n3330 = n3326 & ~n3329;
  assign n3331 = ~n3328 & ~n3330;
  assign n3332 = n3309 & n3331;
  assign n3333 = ~n3284 & ~n3332;
  assign n3334 = ~n3309 & ~n3331;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = pi439  & ~pi440 ;
  assign n3337 = ~pi439  & pi440 ;
  assign n3338 = ~n3336 & ~n3337;
  assign n3339 = ~pi441  & ~n3338;
  assign n3340 = pi441  & n3338;
  assign n3341 = ~n3339 & ~n3340;
  assign n3342 = pi442  & ~pi443 ;
  assign n3343 = ~pi442  & pi443 ;
  assign n3344 = ~n3342 & ~n3343;
  assign n3345 = ~pi444  & ~n3344;
  assign n3346 = pi444  & n3344;
  assign n3347 = ~n3345 & ~n3346;
  assign n3348 = ~n3341 & ~n3347;
  assign n3349 = pi442  & pi443 ;
  assign n3350 = pi444  & ~n3344;
  assign n3351 = ~n3349 & ~n3350;
  assign n3352 = pi439  & pi440 ;
  assign n3353 = pi441  & ~n3338;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355 = n3351 & ~n3354;
  assign n3356 = ~n3351 & n3354;
  assign n3357 = ~n3355 & ~n3356;
  assign n3358 = n3348 & ~n3357;
  assign n3359 = ~n3351 & ~n3354;
  assign n3360 = ~n3358 & ~n3359;
  assign n3361 = pi448  & pi449 ;
  assign n3362 = pi448  & ~pi449 ;
  assign n3363 = ~pi448  & pi449 ;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = pi450  & ~n3364;
  assign n3366 = ~n3361 & ~n3365;
  assign n3367 = pi445  & pi446 ;
  assign n3368 = pi445  & ~pi446 ;
  assign n3369 = ~pi445  & pi446 ;
  assign n3370 = ~n3368 & ~n3369;
  assign n3371 = pi447  & ~n3370;
  assign n3372 = ~n3367 & ~n3371;
  assign n3373 = ~n3366 & n3372;
  assign n3374 = n3366 & ~n3372;
  assign n3375 = ~n3373 & ~n3374;
  assign n3376 = ~pi447  & ~n3370;
  assign n3377 = pi447  & n3370;
  assign n3378 = ~n3376 & ~n3377;
  assign n3379 = ~pi450  & ~n3364;
  assign n3380 = pi450  & n3364;
  assign n3381 = ~n3379 & ~n3380;
  assign n3382 = ~n3378 & ~n3381;
  assign n3383 = ~n3375 & n3382;
  assign n3384 = ~n3366 & ~n3372;
  assign n3385 = ~n3383 & ~n3384;
  assign n3386 = n3348 & n3357;
  assign n3387 = ~n3348 & ~n3357;
  assign n3388 = ~n3386 & ~n3387;
  assign n3389 = n3375 & n3382;
  assign n3390 = ~n3375 & ~n3382;
  assign n3391 = ~n3389 & ~n3390;
  assign n3392 = ~n3385 & ~n3391;
  assign n3393 = ~n3360 & ~n3388;
  assign n3394 = ~n3341 & n3347;
  assign n3395 = n3341 & ~n3347;
  assign n3396 = ~n3394 & ~n3395;
  assign n3397 = ~n3378 & n3381;
  assign n3398 = n3378 & ~n3381;
  assign n3399 = ~n3397 & ~n3398;
  assign n3400 = ~n3396 & ~n3399;
  assign n3401 = ~n3392 & n3400;
  assign n3402 = ~n3393 & n3401;
  assign n3403 = n3391 & ~n3402;
  assign n3404 = ~n3388 & ~n3403;
  assign n3405 = ~n3391 & n3402;
  assign n3406 = ~n3404 & ~n3405;
  assign n3407 = n3385 & n3406;
  assign n3408 = ~n3360 & ~n3407;
  assign n3409 = ~n3385 & ~n3406;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = n3335 & n3410;
  assign n3412 = ~n3360 & n3385;
  assign n3413 = n3360 & ~n3385;
  assign n3414 = ~n3412 & ~n3413;
  assign n3415 = ~n3406 & ~n3414;
  assign n3416 = n3406 & n3414;
  assign n3417 = ~n3415 & ~n3416;
  assign n3418 = ~n3284 & n3309;
  assign n3419 = n3284 & ~n3309;
  assign n3420 = ~n3418 & ~n3419;
  assign n3421 = ~n3331 & ~n3420;
  assign n3422 = n3331 & n3420;
  assign n3423 = ~n3421 & ~n3422;
  assign n3424 = n3417 & n3423;
  assign n3425 = ~n3320 & n3323;
  assign n3426 = n3320 & ~n3323;
  assign n3427 = ~n3425 & ~n3426;
  assign n3428 = ~n3396 & n3399;
  assign n3429 = n3396 & ~n3399;
  assign n3430 = ~n3428 & ~n3429;
  assign n3431 = ~n3427 & ~n3430;
  assign n3432 = ~n3315 & ~n3326;
  assign n3433 = ~n3329 & ~n3432;
  assign n3434 = ~n3312 & n3433;
  assign n3435 = n3312 & ~n3433;
  assign n3436 = ~n3434 & ~n3435;
  assign n3437 = n3431 & ~n3436;
  assign n3438 = ~n3403 & ~n3405;
  assign n3439 = n3388 & n3438;
  assign n3440 = ~n3388 & ~n3438;
  assign n3441 = ~n3439 & ~n3440;
  assign n3442 = ~n3431 & n3436;
  assign n3443 = ~n3441 & ~n3442;
  assign n3444 = ~n3437 & ~n3443;
  assign n3445 = ~n3417 & ~n3423;
  assign n3446 = ~n3424 & ~n3445;
  assign n3447 = ~n3444 & n3446;
  assign n3448 = ~n3424 & ~n3447;
  assign n3449 = ~n3411 & ~n3448;
  assign n3450 = ~n3335 & ~n3410;
  assign n3451 = ~n3449 & ~n3450;
  assign n3452 = pi418  & pi419 ;
  assign n3453 = ~pi418  & pi419 ;
  assign n3454 = pi418  & ~pi419 ;
  assign n3455 = ~n3453 & ~n3454;
  assign n3456 = pi420  & ~n3455;
  assign n3457 = ~n3452 & ~n3456;
  assign n3458 = pi415  & pi416 ;
  assign n3459 = ~pi415  & pi416 ;
  assign n3460 = pi415  & ~pi416 ;
  assign n3461 = ~n3459 & ~n3460;
  assign n3462 = pi417  & ~n3461;
  assign n3463 = ~n3458 & ~n3462;
  assign n3464 = ~n3457 & n3463;
  assign n3465 = n3457 & ~n3463;
  assign n3466 = ~n3464 & ~n3465;
  assign n3467 = ~pi417  & ~n3461;
  assign n3468 = pi417  & n3461;
  assign n3469 = ~n3467 & ~n3468;
  assign n3470 = ~pi420  & ~n3455;
  assign n3471 = pi420  & n3455;
  assign n3472 = ~n3470 & ~n3471;
  assign n3473 = ~n3469 & ~n3472;
  assign n3474 = n3466 & n3473;
  assign n3475 = ~n3466 & ~n3473;
  assign n3476 = ~n3474 & ~n3475;
  assign n3477 = pi424  & pi425 ;
  assign n3478 = ~pi424  & pi425 ;
  assign n3479 = pi424  & ~pi425 ;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = pi426  & ~n3480;
  assign n3482 = ~n3477 & ~n3481;
  assign n3483 = pi421  & pi422 ;
  assign n3484 = ~pi421  & pi422 ;
  assign n3485 = pi421  & ~pi422 ;
  assign n3486 = ~n3484 & ~n3485;
  assign n3487 = pi423  & ~n3486;
  assign n3488 = ~n3483 & ~n3487;
  assign n3489 = ~n3482 & n3488;
  assign n3490 = n3482 & ~n3488;
  assign n3491 = ~n3489 & ~n3490;
  assign n3492 = ~pi423  & ~n3486;
  assign n3493 = pi423  & n3486;
  assign n3494 = ~n3492 & ~n3493;
  assign n3495 = ~pi426  & ~n3480;
  assign n3496 = pi426  & n3480;
  assign n3497 = ~n3495 & ~n3496;
  assign n3498 = ~n3494 & ~n3497;
  assign n3499 = n3491 & n3498;
  assign n3500 = ~n3491 & ~n3498;
  assign n3501 = ~n3499 & ~n3500;
  assign n3502 = ~n3491 & n3498;
  assign n3503 = ~n3482 & ~n3488;
  assign n3504 = ~n3502 & ~n3503;
  assign n3505 = ~n3501 & ~n3504;
  assign n3506 = ~n3466 & n3473;
  assign n3507 = ~n3457 & ~n3463;
  assign n3508 = ~n3506 & ~n3507;
  assign n3509 = ~n3476 & ~n3508;
  assign n3510 = ~n3494 & n3497;
  assign n3511 = n3494 & ~n3497;
  assign n3512 = ~n3510 & ~n3511;
  assign n3513 = ~n3469 & n3472;
  assign n3514 = n3469 & ~n3472;
  assign n3515 = ~n3513 & ~n3514;
  assign n3516 = ~n3512 & ~n3515;
  assign n3517 = ~n3505 & n3516;
  assign n3518 = ~n3509 & n3517;
  assign n3519 = n3501 & ~n3518;
  assign n3520 = ~n3476 & ~n3519;
  assign n3521 = ~n3501 & n3518;
  assign n3522 = ~n3520 & ~n3521;
  assign n3523 = n3504 & ~n3508;
  assign n3524 = ~n3504 & n3508;
  assign n3525 = ~n3523 & ~n3524;
  assign n3526 = ~n3522 & ~n3525;
  assign n3527 = n3522 & n3525;
  assign n3528 = ~n3526 & ~n3527;
  assign n3529 = pi427  & ~pi428 ;
  assign n3530 = ~pi427  & pi428 ;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = ~pi429  & ~n3531;
  assign n3533 = pi429  & n3531;
  assign n3534 = ~n3532 & ~n3533;
  assign n3535 = pi430  & ~pi431 ;
  assign n3536 = ~pi430  & pi431 ;
  assign n3537 = ~n3535 & ~n3536;
  assign n3538 = ~pi432  & ~n3537;
  assign n3539 = pi432  & n3537;
  assign n3540 = ~n3538 & ~n3539;
  assign n3541 = ~n3534 & ~n3540;
  assign n3542 = pi430  & pi431 ;
  assign n3543 = pi432  & ~n3537;
  assign n3544 = ~n3542 & ~n3543;
  assign n3545 = pi427  & pi428 ;
  assign n3546 = pi429  & ~n3531;
  assign n3547 = ~n3545 & ~n3546;
  assign n3548 = n3544 & ~n3547;
  assign n3549 = ~n3544 & n3547;
  assign n3550 = ~n3548 & ~n3549;
  assign n3551 = n3541 & n3550;
  assign n3552 = ~n3541 & ~n3550;
  assign n3553 = ~n3551 & ~n3552;
  assign n3554 = pi436  & pi437 ;
  assign n3555 = pi436  & ~pi437 ;
  assign n3556 = ~pi436  & pi437 ;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = pi438  & ~n3557;
  assign n3559 = ~n3554 & ~n3558;
  assign n3560 = pi433  & pi434 ;
  assign n3561 = pi433  & ~pi434 ;
  assign n3562 = ~pi433  & pi434 ;
  assign n3563 = ~n3561 & ~n3562;
  assign n3564 = pi435  & ~n3563;
  assign n3565 = ~n3560 & ~n3564;
  assign n3566 = ~n3559 & n3565;
  assign n3567 = n3559 & ~n3565;
  assign n3568 = ~n3566 & ~n3567;
  assign n3569 = ~pi435  & ~n3563;
  assign n3570 = pi435  & n3563;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = ~pi438  & ~n3557;
  assign n3573 = pi438  & n3557;
  assign n3574 = ~n3572 & ~n3573;
  assign n3575 = ~n3571 & ~n3574;
  assign n3576 = n3568 & n3575;
  assign n3577 = ~n3568 & ~n3575;
  assign n3578 = ~n3576 & ~n3577;
  assign n3579 = ~n3568 & n3575;
  assign n3580 = ~n3559 & ~n3565;
  assign n3581 = ~n3579 & ~n3580;
  assign n3582 = ~n3578 & ~n3581;
  assign n3583 = n3541 & ~n3550;
  assign n3584 = ~n3544 & ~n3547;
  assign n3585 = ~n3583 & ~n3584;
  assign n3586 = ~n3553 & ~n3585;
  assign n3587 = ~n3534 & n3540;
  assign n3588 = n3534 & ~n3540;
  assign n3589 = ~n3587 & ~n3588;
  assign n3590 = ~n3571 & n3574;
  assign n3591 = n3571 & ~n3574;
  assign n3592 = ~n3590 & ~n3591;
  assign n3593 = ~n3589 & ~n3592;
  assign n3594 = ~n3582 & n3593;
  assign n3595 = ~n3586 & n3594;
  assign n3596 = n3578 & ~n3595;
  assign n3597 = ~n3553 & ~n3596;
  assign n3598 = n3578 & n3595;
  assign n3599 = n3595 & ~n3598;
  assign n3600 = ~n3597 & ~n3599;
  assign n3601 = n3581 & ~n3585;
  assign n3602 = ~n3581 & n3585;
  assign n3603 = ~n3601 & ~n3602;
  assign n3604 = ~n3600 & ~n3603;
  assign n3605 = n3600 & n3603;
  assign n3606 = ~n3604 & ~n3605;
  assign n3607 = n3528 & n3606;
  assign n3608 = ~n3589 & n3592;
  assign n3609 = n3589 & ~n3592;
  assign n3610 = ~n3608 & ~n3609;
  assign n3611 = n3512 & ~n3515;
  assign n3612 = ~n3512 & n3515;
  assign n3613 = ~n3611 & ~n3612;
  assign n3614 = ~n3610 & ~n3613;
  assign n3615 = ~n3578 & ~n3595;
  assign n3616 = ~n3598 & ~n3615;
  assign n3617 = ~n3553 & n3616;
  assign n3618 = n3553 & ~n3616;
  assign n3619 = ~n3617 & ~n3618;
  assign n3620 = n3614 & ~n3619;
  assign n3621 = ~n3519 & ~n3521;
  assign n3622 = n3476 & n3621;
  assign n3623 = ~n3476 & ~n3621;
  assign n3624 = ~n3622 & ~n3623;
  assign n3625 = ~n3614 & n3619;
  assign n3626 = ~n3624 & ~n3625;
  assign n3627 = ~n3620 & ~n3626;
  assign n3628 = ~n3528 & ~n3606;
  assign n3629 = ~n3627 & ~n3628;
  assign n3630 = ~n3607 & ~n3629;
  assign n3631 = n3581 & n3600;
  assign n3632 = ~n3585 & ~n3631;
  assign n3633 = ~n3581 & ~n3600;
  assign n3634 = ~n3632 & ~n3633;
  assign n3635 = n3504 & n3522;
  assign n3636 = ~n3508 & ~n3635;
  assign n3637 = ~n3504 & ~n3522;
  assign n3638 = ~n3636 & ~n3637;
  assign n3639 = n3634 & n3638;
  assign n3640 = ~n3630 & ~n3639;
  assign n3641 = ~n3634 & ~n3638;
  assign n3642 = ~n3640 & ~n3641;
  assign n3643 = ~n3451 & ~n3642;
  assign n3644 = ~n3427 & n3430;
  assign n3645 = n3427 & ~n3430;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = ~n3610 & n3613;
  assign n3648 = n3610 & ~n3613;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650 = ~n3646 & ~n3649;
  assign n3651 = ~n3437 & ~n3442;
  assign n3652 = ~n3441 & ~n3651;
  assign n3653 = n3441 & n3651;
  assign n3654 = ~n3652 & ~n3653;
  assign n3655 = n3650 & ~n3654;
  assign n3656 = ~n3620 & ~n3625;
  assign n3657 = n3624 & n3656;
  assign n3658 = ~n3624 & ~n3656;
  assign n3659 = ~n3657 & ~n3658;
  assign n3660 = ~n3650 & n3654;
  assign n3661 = ~n3659 & ~n3660;
  assign n3662 = ~n3655 & ~n3661;
  assign n3663 = ~n3607 & ~n3628;
  assign n3664 = ~n3627 & n3663;
  assign n3665 = n3627 & ~n3663;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = n3444 & ~n3446;
  assign n3668 = ~n3447 & ~n3667;
  assign n3669 = ~n3666 & ~n3668;
  assign n3670 = ~n3662 & ~n3669;
  assign n3671 = n3666 & n3668;
  assign n3672 = ~n3670 & ~n3671;
  assign n3673 = ~n3411 & ~n3450;
  assign n3674 = ~n3448 & n3673;
  assign n3675 = n3448 & ~n3673;
  assign n3676 = ~n3674 & ~n3675;
  assign n3677 = n3634 & ~n3638;
  assign n3678 = ~n3634 & n3638;
  assign n3679 = ~n3607 & ~n3677;
  assign n3680 = ~n3678 & n3679;
  assign n3681 = ~n3629 & n3680;
  assign n3682 = n3640 & ~n3641;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = ~n3676 & ~n3683;
  assign n3685 = ~n3672 & ~n3684;
  assign n3686 = n3676 & n3683;
  assign n3687 = ~n3685 & ~n3686;
  assign n3688 = n3451 & n3642;
  assign n3689 = ~n3643 & ~n3688;
  assign n3690 = ~n3687 & n3689;
  assign n3691 = ~n3643 & ~n3690;
  assign n3692 = pi403  & ~pi404 ;
  assign n3693 = ~pi403  & pi404 ;
  assign n3694 = ~n3692 & ~n3693;
  assign n3695 = ~pi405  & ~n3694;
  assign n3696 = pi405  & n3694;
  assign n3697 = ~n3695 & ~n3696;
  assign n3698 = pi406  & ~pi407 ;
  assign n3699 = ~pi406  & pi407 ;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = ~pi408  & ~n3700;
  assign n3702 = pi408  & n3700;
  assign n3703 = ~n3701 & ~n3702;
  assign n3704 = ~n3697 & ~n3703;
  assign n3705 = pi406  & pi407 ;
  assign n3706 = pi408  & ~n3700;
  assign n3707 = ~n3705 & ~n3706;
  assign n3708 = pi403  & pi404 ;
  assign n3709 = pi405  & ~n3694;
  assign n3710 = ~n3708 & ~n3709;
  assign n3711 = n3707 & ~n3710;
  assign n3712 = ~n3707 & n3710;
  assign n3713 = ~n3711 & ~n3712;
  assign n3714 = n3704 & ~n3713;
  assign n3715 = ~n3707 & ~n3710;
  assign n3716 = ~n3714 & ~n3715;
  assign n3717 = pi412  & pi413 ;
  assign n3718 = pi412  & ~pi413 ;
  assign n3719 = ~pi412  & pi413 ;
  assign n3720 = ~n3718 & ~n3719;
  assign n3721 = pi414  & ~n3720;
  assign n3722 = ~n3717 & ~n3721;
  assign n3723 = pi409  & pi410 ;
  assign n3724 = pi409  & ~pi410 ;
  assign n3725 = ~pi409  & pi410 ;
  assign n3726 = ~n3724 & ~n3725;
  assign n3727 = pi411  & ~n3726;
  assign n3728 = ~n3723 & ~n3727;
  assign n3729 = ~n3722 & n3728;
  assign n3730 = n3722 & ~n3728;
  assign n3731 = ~n3729 & ~n3730;
  assign n3732 = ~pi411  & ~n3726;
  assign n3733 = pi411  & n3726;
  assign n3734 = ~n3732 & ~n3733;
  assign n3735 = ~pi414  & ~n3720;
  assign n3736 = pi414  & n3720;
  assign n3737 = ~n3735 & ~n3736;
  assign n3738 = ~n3734 & ~n3737;
  assign n3739 = ~n3731 & n3738;
  assign n3740 = ~n3722 & ~n3728;
  assign n3741 = ~n3739 & ~n3740;
  assign n3742 = n3704 & n3713;
  assign n3743 = ~n3704 & ~n3713;
  assign n3744 = ~n3742 & ~n3743;
  assign n3745 = n3731 & n3738;
  assign n3746 = ~n3731 & ~n3738;
  assign n3747 = ~n3745 & ~n3746;
  assign n3748 = ~n3741 & ~n3747;
  assign n3749 = ~n3716 & ~n3744;
  assign n3750 = ~n3697 & n3703;
  assign n3751 = n3697 & ~n3703;
  assign n3752 = ~n3750 & ~n3751;
  assign n3753 = ~n3734 & n3737;
  assign n3754 = n3734 & ~n3737;
  assign n3755 = ~n3753 & ~n3754;
  assign n3756 = ~n3752 & ~n3755;
  assign n3757 = ~n3748 & n3756;
  assign n3758 = ~n3749 & n3757;
  assign n3759 = n3747 & ~n3758;
  assign n3760 = ~n3744 & ~n3759;
  assign n3761 = n3747 & n3758;
  assign n3762 = n3758 & ~n3761;
  assign n3763 = ~n3760 & ~n3762;
  assign n3764 = n3741 & n3763;
  assign n3765 = ~n3716 & ~n3764;
  assign n3766 = ~n3741 & ~n3763;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = pi391  & ~pi392 ;
  assign n3769 = ~pi391  & pi392 ;
  assign n3770 = ~n3768 & ~n3769;
  assign n3771 = ~pi393  & ~n3770;
  assign n3772 = pi393  & n3770;
  assign n3773 = ~n3771 & ~n3772;
  assign n3774 = pi394  & ~pi395 ;
  assign n3775 = ~pi394  & pi395 ;
  assign n3776 = ~n3774 & ~n3775;
  assign n3777 = ~pi396  & ~n3776;
  assign n3778 = pi396  & n3776;
  assign n3779 = ~n3777 & ~n3778;
  assign n3780 = ~n3773 & ~n3779;
  assign n3781 = pi394  & pi395 ;
  assign n3782 = pi396  & ~n3776;
  assign n3783 = ~n3781 & ~n3782;
  assign n3784 = pi391  & pi392 ;
  assign n3785 = pi393  & ~n3770;
  assign n3786 = ~n3784 & ~n3785;
  assign n3787 = n3783 & ~n3786;
  assign n3788 = ~n3783 & n3786;
  assign n3789 = ~n3787 & ~n3788;
  assign n3790 = n3780 & ~n3789;
  assign n3791 = ~n3783 & ~n3786;
  assign n3792 = ~n3790 & ~n3791;
  assign n3793 = pi400  & pi401 ;
  assign n3794 = pi400  & ~pi401 ;
  assign n3795 = ~pi400  & pi401 ;
  assign n3796 = ~n3794 & ~n3795;
  assign n3797 = pi402  & ~n3796;
  assign n3798 = ~n3793 & ~n3797;
  assign n3799 = pi397  & pi398 ;
  assign n3800 = pi397  & ~pi398 ;
  assign n3801 = ~pi397  & pi398 ;
  assign n3802 = ~n3800 & ~n3801;
  assign n3803 = pi399  & ~n3802;
  assign n3804 = ~n3799 & ~n3803;
  assign n3805 = ~n3798 & n3804;
  assign n3806 = n3798 & ~n3804;
  assign n3807 = ~n3805 & ~n3806;
  assign n3808 = ~pi399  & ~n3802;
  assign n3809 = pi399  & n3802;
  assign n3810 = ~n3808 & ~n3809;
  assign n3811 = ~pi402  & ~n3796;
  assign n3812 = pi402  & n3796;
  assign n3813 = ~n3811 & ~n3812;
  assign n3814 = ~n3810 & ~n3813;
  assign n3815 = ~n3807 & n3814;
  assign n3816 = ~n3798 & ~n3804;
  assign n3817 = ~n3815 & ~n3816;
  assign n3818 = n3780 & n3789;
  assign n3819 = ~n3780 & ~n3789;
  assign n3820 = ~n3818 & ~n3819;
  assign n3821 = n3807 & n3814;
  assign n3822 = ~n3807 & ~n3814;
  assign n3823 = ~n3821 & ~n3822;
  assign n3824 = ~n3817 & ~n3823;
  assign n3825 = ~n3792 & ~n3820;
  assign n3826 = ~n3773 & n3779;
  assign n3827 = n3773 & ~n3779;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = ~n3810 & n3813;
  assign n3830 = n3810 & ~n3813;
  assign n3831 = ~n3829 & ~n3830;
  assign n3832 = ~n3828 & ~n3831;
  assign n3833 = ~n3824 & n3832;
  assign n3834 = ~n3825 & n3833;
  assign n3835 = n3823 & ~n3834;
  assign n3836 = ~n3820 & ~n3835;
  assign n3837 = ~n3823 & n3834;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = n3817 & n3838;
  assign n3840 = ~n3792 & ~n3839;
  assign n3841 = ~n3817 & ~n3838;
  assign n3842 = ~n3840 & ~n3841;
  assign n3843 = n3767 & n3842;
  assign n3844 = ~n3792 & n3817;
  assign n3845 = n3792 & ~n3817;
  assign n3846 = ~n3844 & ~n3845;
  assign n3847 = ~n3838 & ~n3846;
  assign n3848 = n3838 & n3846;
  assign n3849 = ~n3847 & ~n3848;
  assign n3850 = ~n3716 & n3741;
  assign n3851 = n3716 & ~n3741;
  assign n3852 = ~n3850 & ~n3851;
  assign n3853 = ~n3763 & ~n3852;
  assign n3854 = n3763 & n3852;
  assign n3855 = ~n3853 & ~n3854;
  assign n3856 = n3849 & n3855;
  assign n3857 = ~n3752 & n3755;
  assign n3858 = n3752 & ~n3755;
  assign n3859 = ~n3857 & ~n3858;
  assign n3860 = ~n3828 & n3831;
  assign n3861 = n3828 & ~n3831;
  assign n3862 = ~n3860 & ~n3861;
  assign n3863 = ~n3859 & ~n3862;
  assign n3864 = ~n3747 & ~n3758;
  assign n3865 = ~n3761 & ~n3864;
  assign n3866 = ~n3744 & n3865;
  assign n3867 = n3744 & ~n3865;
  assign n3868 = ~n3866 & ~n3867;
  assign n3869 = n3863 & ~n3868;
  assign n3870 = ~n3835 & ~n3837;
  assign n3871 = n3820 & n3870;
  assign n3872 = ~n3820 & ~n3870;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = ~n3863 & n3868;
  assign n3875 = ~n3873 & ~n3874;
  assign n3876 = ~n3869 & ~n3875;
  assign n3877 = ~n3849 & ~n3855;
  assign n3878 = ~n3856 & ~n3877;
  assign n3879 = ~n3876 & n3878;
  assign n3880 = ~n3856 & ~n3879;
  assign n3881 = ~n3843 & ~n3880;
  assign n3882 = ~n3767 & ~n3842;
  assign n3883 = ~n3881 & ~n3882;
  assign n3884 = ~pi385  & pi386 ;
  assign n3885 = pi385  & ~pi386 ;
  assign n3886 = ~n3884 & ~n3885;
  assign n3887 = ~pi387  & ~n3886;
  assign n3888 = pi387  & n3886;
  assign n3889 = ~n3887 & ~n3888;
  assign n3890 = ~pi388  & pi389 ;
  assign n3891 = pi388  & ~pi389 ;
  assign n3892 = ~n3890 & ~n3891;
  assign n3893 = ~pi390  & ~n3892;
  assign n3894 = pi390  & n3892;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = ~n3889 & n3895;
  assign n3897 = n3889 & ~n3895;
  assign n3898 = ~n3896 & ~n3897;
  assign n3899 = ~pi379  & pi380 ;
  assign n3900 = pi379  & ~pi380 ;
  assign n3901 = ~n3899 & ~n3900;
  assign n3902 = ~pi381  & ~n3901;
  assign n3903 = pi381  & n3901;
  assign n3904 = ~n3902 & ~n3903;
  assign n3905 = ~pi382  & pi383 ;
  assign n3906 = pi382  & ~pi383 ;
  assign n3907 = ~n3905 & ~n3906;
  assign n3908 = ~pi384  & ~n3907;
  assign n3909 = pi384  & n3907;
  assign n3910 = ~n3908 & ~n3909;
  assign n3911 = ~n3904 & n3910;
  assign n3912 = n3904 & ~n3910;
  assign n3913 = ~n3911 & ~n3912;
  assign n3914 = n3898 & ~n3913;
  assign n3915 = ~n3898 & n3913;
  assign n3916 = ~n3914 & ~n3915;
  assign n3917 = ~pi373  & pi374 ;
  assign n3918 = pi373  & ~pi374 ;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = ~pi375  & ~n3919;
  assign n3921 = pi375  & n3919;
  assign n3922 = ~n3920 & ~n3921;
  assign n3923 = ~pi376  & pi377 ;
  assign n3924 = pi376  & ~pi377 ;
  assign n3925 = ~n3923 & ~n3924;
  assign n3926 = ~pi378  & ~n3925;
  assign n3927 = pi378  & n3925;
  assign n3928 = ~n3926 & ~n3927;
  assign n3929 = ~n3922 & n3928;
  assign n3930 = n3922 & ~n3928;
  assign n3931 = ~n3929 & ~n3930;
  assign n3932 = ~pi367  & pi368 ;
  assign n3933 = pi367  & ~pi368 ;
  assign n3934 = ~n3932 & ~n3933;
  assign n3935 = ~pi369  & ~n3934;
  assign n3936 = pi369  & n3934;
  assign n3937 = ~n3935 & ~n3936;
  assign n3938 = ~pi370  & pi371 ;
  assign n3939 = pi370  & ~pi371 ;
  assign n3940 = ~n3938 & ~n3939;
  assign n3941 = ~pi372  & ~n3940;
  assign n3942 = pi372  & n3940;
  assign n3943 = ~n3941 & ~n3942;
  assign n3944 = ~n3937 & n3943;
  assign n3945 = n3937 & ~n3943;
  assign n3946 = ~n3944 & ~n3945;
  assign n3947 = n3931 & ~n3946;
  assign n3948 = ~n3931 & n3946;
  assign n3949 = ~n3947 & ~n3948;
  assign n3950 = ~n3916 & ~n3949;
  assign n3951 = pi382  & pi383 ;
  assign n3952 = pi384  & ~n3907;
  assign n3953 = ~n3951 & ~n3952;
  assign n3954 = pi379  & pi380 ;
  assign n3955 = pi381  & ~n3901;
  assign n3956 = ~n3954 & ~n3955;
  assign n3957 = ~n3953 & n3956;
  assign n3958 = n3953 & ~n3956;
  assign n3959 = ~n3957 & ~n3958;
  assign n3960 = ~n3904 & ~n3910;
  assign n3961 = n3959 & n3960;
  assign n3962 = ~n3959 & ~n3960;
  assign n3963 = ~n3961 & ~n3962;
  assign n3964 = pi388  & pi389 ;
  assign n3965 = pi390  & ~n3892;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = pi385  & pi386 ;
  assign n3968 = pi387  & ~n3886;
  assign n3969 = ~n3967 & ~n3968;
  assign n3970 = ~n3966 & n3969;
  assign n3971 = n3966 & ~n3969;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = ~n3889 & ~n3895;
  assign n3974 = n3972 & n3973;
  assign n3975 = ~n3972 & ~n3973;
  assign n3976 = ~n3974 & ~n3975;
  assign n3977 = ~n3972 & n3973;
  assign n3978 = ~n3966 & ~n3969;
  assign n3979 = ~n3977 & ~n3978;
  assign n3980 = ~n3976 & ~n3979;
  assign n3981 = ~n3959 & n3960;
  assign n3982 = ~n3953 & ~n3956;
  assign n3983 = ~n3981 & ~n3982;
  assign n3984 = ~n3963 & ~n3983;
  assign n3985 = ~n3898 & ~n3913;
  assign n3986 = ~n3980 & n3985;
  assign n3987 = ~n3984 & n3986;
  assign n3988 = n3976 & ~n3987;
  assign n3989 = ~n3976 & n3987;
  assign n3990 = ~n3988 & ~n3989;
  assign n3991 = ~n3963 & ~n3990;
  assign n3992 = n3963 & n3990;
  assign n3993 = ~n3991 & ~n3992;
  assign n3994 = n3950 & ~n3993;
  assign n3995 = pi370  & pi371 ;
  assign n3996 = pi372  & ~n3940;
  assign n3997 = ~n3995 & ~n3996;
  assign n3998 = pi367  & pi368 ;
  assign n3999 = pi369  & ~n3934;
  assign n4000 = ~n3998 & ~n3999;
  assign n4001 = ~n3997 & n4000;
  assign n4002 = n3997 & ~n4000;
  assign n4003 = ~n4001 & ~n4002;
  assign n4004 = ~n3937 & ~n3943;
  assign n4005 = n4003 & n4004;
  assign n4006 = ~n4003 & ~n4004;
  assign n4007 = ~n4005 & ~n4006;
  assign n4008 = pi376  & pi377 ;
  assign n4009 = pi378  & ~n3925;
  assign n4010 = ~n4008 & ~n4009;
  assign n4011 = pi373  & pi374 ;
  assign n4012 = pi375  & ~n3919;
  assign n4013 = ~n4011 & ~n4012;
  assign n4014 = ~n4010 & n4013;
  assign n4015 = n4010 & ~n4013;
  assign n4016 = ~n4014 & ~n4015;
  assign n4017 = ~n3922 & ~n3928;
  assign n4018 = n4016 & n4017;
  assign n4019 = ~n4016 & ~n4017;
  assign n4020 = ~n4018 & ~n4019;
  assign n4021 = ~n4016 & n4017;
  assign n4022 = ~n4010 & ~n4013;
  assign n4023 = ~n4021 & ~n4022;
  assign n4024 = ~n4020 & ~n4023;
  assign n4025 = ~n4003 & n4004;
  assign n4026 = ~n3997 & ~n4000;
  assign n4027 = ~n4025 & ~n4026;
  assign n4028 = ~n4007 & ~n4027;
  assign n4029 = ~n3931 & ~n3946;
  assign n4030 = ~n4024 & n4029;
  assign n4031 = ~n4028 & n4030;
  assign n4032 = n4020 & ~n4031;
  assign n4033 = ~n4020 & n4031;
  assign n4034 = ~n4032 & ~n4033;
  assign n4035 = n4007 & n4034;
  assign n4036 = ~n4007 & ~n4034;
  assign n4037 = ~n4035 & ~n4036;
  assign n4038 = ~n3950 & n3993;
  assign n4039 = ~n4037 & ~n4038;
  assign n4040 = ~n3994 & ~n4039;
  assign n4041 = ~n4007 & ~n4032;
  assign n4042 = ~n4033 & ~n4041;
  assign n4043 = n4023 & ~n4027;
  assign n4044 = ~n4023 & n4027;
  assign n4045 = ~n4043 & ~n4044;
  assign n4046 = ~n4042 & ~n4045;
  assign n4047 = n4042 & n4045;
  assign n4048 = ~n4046 & ~n4047;
  assign n4049 = ~n3963 & ~n3988;
  assign n4050 = ~n3989 & ~n4049;
  assign n4051 = n3979 & ~n3983;
  assign n4052 = ~n3979 & n3983;
  assign n4053 = ~n4051 & ~n4052;
  assign n4054 = ~n4050 & ~n4053;
  assign n4055 = n4050 & n4053;
  assign n4056 = ~n4054 & ~n4055;
  assign n4057 = ~n4048 & ~n4056;
  assign n4058 = ~n4040 & ~n4057;
  assign n4059 = n4048 & n4056;
  assign n4060 = ~n4058 & ~n4059;
  assign n4061 = n3979 & n4050;
  assign n4062 = ~n3983 & ~n4061;
  assign n4063 = ~n3979 & ~n4050;
  assign n4064 = ~n4062 & ~n4063;
  assign n4065 = n4023 & n4042;
  assign n4066 = ~n4027 & ~n4065;
  assign n4067 = ~n4023 & ~n4042;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = n4064 & n4068;
  assign n4070 = ~n4060 & ~n4069;
  assign n4071 = ~n4064 & ~n4068;
  assign n4072 = ~n4070 & ~n4071;
  assign n4073 = ~n3883 & ~n4072;
  assign n4074 = ~n4057 & ~n4059;
  assign n4075 = ~n4040 & n4074;
  assign n4076 = n4040 & ~n4074;
  assign n4077 = ~n4075 & ~n4076;
  assign n4078 = n3876 & ~n3878;
  assign n4079 = ~n3879 & ~n4078;
  assign n4080 = n4077 & n4079;
  assign n4081 = ~n3859 & n3862;
  assign n4082 = n3859 & ~n3862;
  assign n4083 = ~n4081 & ~n4082;
  assign n4084 = ~n3916 & n3949;
  assign n4085 = n3916 & ~n3949;
  assign n4086 = ~n4084 & ~n4085;
  assign n4087 = ~n4083 & ~n4086;
  assign n4088 = ~n3869 & ~n3874;
  assign n4089 = ~n3873 & ~n4088;
  assign n4090 = n3873 & n4088;
  assign n4091 = ~n4089 & ~n4090;
  assign n4092 = n4087 & ~n4091;
  assign n4093 = ~n3994 & ~n4038;
  assign n4094 = n4037 & n4093;
  assign n4095 = ~n4037 & ~n4093;
  assign n4096 = ~n4094 & ~n4095;
  assign n4097 = ~n4087 & n4091;
  assign n4098 = ~n4096 & ~n4097;
  assign n4099 = ~n4092 & ~n4098;
  assign n4100 = ~n4077 & ~n4079;
  assign n4101 = ~n4080 & ~n4100;
  assign n4102 = ~n4099 & n4101;
  assign n4103 = ~n4080 & ~n4102;
  assign n4104 = ~n3843 & ~n3882;
  assign n4105 = ~n3880 & n4104;
  assign n4106 = n3880 & ~n4104;
  assign n4107 = ~n4105 & ~n4106;
  assign n4108 = n4064 & ~n4068;
  assign n4109 = ~n4064 & n4068;
  assign n4110 = ~n4059 & ~n4108;
  assign n4111 = ~n4109 & n4110;
  assign n4112 = ~n4058 & n4111;
  assign n4113 = n4070 & ~n4071;
  assign n4114 = ~n4112 & ~n4113;
  assign n4115 = ~n4107 & ~n4114;
  assign n4116 = ~n4103 & ~n4115;
  assign n4117 = n4107 & n4114;
  assign n4118 = ~n4116 & ~n4117;
  assign n4119 = n3883 & n4072;
  assign n4120 = ~n4073 & ~n4119;
  assign n4121 = ~n4118 & n4120;
  assign n4122 = ~n4073 & ~n4121;
  assign n4123 = ~n3691 & ~n4122;
  assign n4124 = n3691 & n4122;
  assign n4125 = ~n4123 & ~n4124;
  assign n4126 = n4118 & ~n4120;
  assign n4127 = ~n4121 & ~n4126;
  assign n4128 = n3687 & ~n3689;
  assign n4129 = ~n3690 & ~n4128;
  assign n4130 = n4127 & n4129;
  assign n4131 = n4099 & ~n4101;
  assign n4132 = ~n4102 & ~n4131;
  assign n4133 = ~n3669 & ~n3671;
  assign n4134 = ~n3662 & n4133;
  assign n4135 = n3662 & ~n4133;
  assign n4136 = ~n4134 & ~n4135;
  assign n4137 = n4132 & n4136;
  assign n4138 = ~n3646 & n3649;
  assign n4139 = n3646 & ~n3649;
  assign n4140 = ~n4138 & ~n4139;
  assign n4141 = ~n4083 & n4086;
  assign n4142 = n4083 & ~n4086;
  assign n4143 = ~n4141 & ~n4142;
  assign n4144 = ~n4140 & ~n4143;
  assign n4145 = ~n3655 & ~n3660;
  assign n4146 = ~n3659 & ~n4145;
  assign n4147 = n3659 & n4145;
  assign n4148 = ~n4146 & ~n4147;
  assign n4149 = n4144 & ~n4148;
  assign n4150 = ~n4092 & ~n4097;
  assign n4151 = n4096 & n4150;
  assign n4152 = ~n4096 & ~n4150;
  assign n4153 = ~n4151 & ~n4152;
  assign n4154 = ~n4144 & n4148;
  assign n4155 = ~n4153 & ~n4154;
  assign n4156 = ~n4149 & ~n4155;
  assign n4157 = ~n4132 & ~n4136;
  assign n4158 = ~n4137 & ~n4157;
  assign n4159 = ~n4156 & n4158;
  assign n4160 = ~n4137 & ~n4159;
  assign n4161 = ~n3684 & ~n3686;
  assign n4162 = ~n3672 & n4161;
  assign n4163 = n3672 & ~n4161;
  assign n4164 = ~n4162 & ~n4163;
  assign n4165 = ~n4115 & ~n4117;
  assign n4166 = ~n4103 & n4165;
  assign n4167 = n4103 & ~n4165;
  assign n4168 = ~n4166 & ~n4167;
  assign n4169 = ~n4164 & ~n4168;
  assign n4170 = ~n4160 & ~n4169;
  assign n4171 = n4164 & n4168;
  assign n4172 = ~n4170 & ~n4171;
  assign n4173 = ~n4127 & ~n4129;
  assign n4174 = ~n4130 & ~n4173;
  assign n4175 = ~n4172 & n4174;
  assign n4176 = ~n4130 & ~n4175;
  assign n4177 = n4125 & ~n4176;
  assign n4178 = ~n4123 & ~n4177;
  assign n4179 = pi355  & ~pi356 ;
  assign n4180 = ~pi355  & pi356 ;
  assign n4181 = ~n4179 & ~n4180;
  assign n4182 = ~pi357  & ~n4181;
  assign n4183 = pi357  & n4181;
  assign n4184 = ~n4182 & ~n4183;
  assign n4185 = pi358  & ~pi359 ;
  assign n4186 = ~pi358  & pi359 ;
  assign n4187 = ~n4185 & ~n4186;
  assign n4188 = ~pi360  & ~n4187;
  assign n4189 = pi360  & n4187;
  assign n4190 = ~n4188 & ~n4189;
  assign n4191 = ~n4184 & ~n4190;
  assign n4192 = pi358  & pi359 ;
  assign n4193 = pi360  & ~n4187;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = pi355  & pi356 ;
  assign n4196 = pi357  & ~n4181;
  assign n4197 = ~n4195 & ~n4196;
  assign n4198 = n4194 & ~n4197;
  assign n4199 = ~n4194 & n4197;
  assign n4200 = ~n4198 & ~n4199;
  assign n4201 = n4191 & ~n4200;
  assign n4202 = ~n4194 & ~n4197;
  assign n4203 = ~n4201 & ~n4202;
  assign n4204 = pi364  & pi365 ;
  assign n4205 = pi364  & ~pi365 ;
  assign n4206 = ~pi364  & pi365 ;
  assign n4207 = ~n4205 & ~n4206;
  assign n4208 = pi366  & ~n4207;
  assign n4209 = ~n4204 & ~n4208;
  assign n4210 = pi361  & pi362 ;
  assign n4211 = pi361  & ~pi362 ;
  assign n4212 = ~pi361  & pi362 ;
  assign n4213 = ~n4211 & ~n4212;
  assign n4214 = pi363  & ~n4213;
  assign n4215 = ~n4210 & ~n4214;
  assign n4216 = ~n4209 & n4215;
  assign n4217 = n4209 & ~n4215;
  assign n4218 = ~n4216 & ~n4217;
  assign n4219 = ~pi363  & ~n4213;
  assign n4220 = pi363  & n4213;
  assign n4221 = ~n4219 & ~n4220;
  assign n4222 = ~pi366  & ~n4207;
  assign n4223 = pi366  & n4207;
  assign n4224 = ~n4222 & ~n4223;
  assign n4225 = ~n4221 & ~n4224;
  assign n4226 = ~n4218 & n4225;
  assign n4227 = ~n4209 & ~n4215;
  assign n4228 = ~n4226 & ~n4227;
  assign n4229 = n4191 & n4200;
  assign n4230 = ~n4191 & ~n4200;
  assign n4231 = ~n4229 & ~n4230;
  assign n4232 = n4218 & n4225;
  assign n4233 = ~n4218 & ~n4225;
  assign n4234 = ~n4232 & ~n4233;
  assign n4235 = ~n4228 & ~n4234;
  assign n4236 = ~n4203 & ~n4231;
  assign n4237 = ~n4184 & n4190;
  assign n4238 = n4184 & ~n4190;
  assign n4239 = ~n4237 & ~n4238;
  assign n4240 = ~n4221 & n4224;
  assign n4241 = n4221 & ~n4224;
  assign n4242 = ~n4240 & ~n4241;
  assign n4243 = ~n4239 & ~n4242;
  assign n4244 = ~n4235 & n4243;
  assign n4245 = ~n4236 & n4244;
  assign n4246 = n4234 & ~n4245;
  assign n4247 = ~n4231 & ~n4246;
  assign n4248 = n4234 & n4245;
  assign n4249 = n4245 & ~n4248;
  assign n4250 = ~n4247 & ~n4249;
  assign n4251 = n4228 & n4250;
  assign n4252 = ~n4203 & ~n4251;
  assign n4253 = ~n4228 & ~n4250;
  assign n4254 = ~n4252 & ~n4253;
  assign n4255 = pi343  & ~pi344 ;
  assign n4256 = ~pi343  & pi344 ;
  assign n4257 = ~n4255 & ~n4256;
  assign n4258 = ~pi345  & ~n4257;
  assign n4259 = pi345  & n4257;
  assign n4260 = ~n4258 & ~n4259;
  assign n4261 = pi346  & ~pi347 ;
  assign n4262 = ~pi346  & pi347 ;
  assign n4263 = ~n4261 & ~n4262;
  assign n4264 = ~pi348  & ~n4263;
  assign n4265 = pi348  & n4263;
  assign n4266 = ~n4264 & ~n4265;
  assign n4267 = ~n4260 & ~n4266;
  assign n4268 = pi346  & pi347 ;
  assign n4269 = pi348  & ~n4263;
  assign n4270 = ~n4268 & ~n4269;
  assign n4271 = pi343  & pi344 ;
  assign n4272 = pi345  & ~n4257;
  assign n4273 = ~n4271 & ~n4272;
  assign n4274 = n4270 & ~n4273;
  assign n4275 = ~n4270 & n4273;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = n4267 & ~n4276;
  assign n4278 = ~n4270 & ~n4273;
  assign n4279 = ~n4277 & ~n4278;
  assign n4280 = pi352  & pi353 ;
  assign n4281 = pi352  & ~pi353 ;
  assign n4282 = ~pi352  & pi353 ;
  assign n4283 = ~n4281 & ~n4282;
  assign n4284 = pi354  & ~n4283;
  assign n4285 = ~n4280 & ~n4284;
  assign n4286 = pi349  & pi350 ;
  assign n4287 = pi349  & ~pi350 ;
  assign n4288 = ~pi349  & pi350 ;
  assign n4289 = ~n4287 & ~n4288;
  assign n4290 = pi351  & ~n4289;
  assign n4291 = ~n4286 & ~n4290;
  assign n4292 = ~n4285 & n4291;
  assign n4293 = n4285 & ~n4291;
  assign n4294 = ~n4292 & ~n4293;
  assign n4295 = ~pi351  & ~n4289;
  assign n4296 = pi351  & n4289;
  assign n4297 = ~n4295 & ~n4296;
  assign n4298 = ~pi354  & ~n4283;
  assign n4299 = pi354  & n4283;
  assign n4300 = ~n4298 & ~n4299;
  assign n4301 = ~n4297 & ~n4300;
  assign n4302 = ~n4294 & n4301;
  assign n4303 = ~n4285 & ~n4291;
  assign n4304 = ~n4302 & ~n4303;
  assign n4305 = n4267 & n4276;
  assign n4306 = ~n4267 & ~n4276;
  assign n4307 = ~n4305 & ~n4306;
  assign n4308 = n4294 & n4301;
  assign n4309 = ~n4294 & ~n4301;
  assign n4310 = ~n4308 & ~n4309;
  assign n4311 = ~n4304 & ~n4310;
  assign n4312 = ~n4279 & ~n4307;
  assign n4313 = ~n4260 & n4266;
  assign n4314 = n4260 & ~n4266;
  assign n4315 = ~n4313 & ~n4314;
  assign n4316 = ~n4297 & n4300;
  assign n4317 = n4297 & ~n4300;
  assign n4318 = ~n4316 & ~n4317;
  assign n4319 = ~n4315 & ~n4318;
  assign n4320 = ~n4311 & n4319;
  assign n4321 = ~n4312 & n4320;
  assign n4322 = n4310 & ~n4321;
  assign n4323 = ~n4307 & ~n4322;
  assign n4324 = ~n4310 & n4321;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = n4304 & n4325;
  assign n4327 = ~n4279 & ~n4326;
  assign n4328 = ~n4304 & ~n4325;
  assign n4329 = ~n4327 & ~n4328;
  assign n4330 = n4254 & n4329;
  assign n4331 = ~n4279 & n4304;
  assign n4332 = n4279 & ~n4304;
  assign n4333 = ~n4331 & ~n4332;
  assign n4334 = ~n4325 & ~n4333;
  assign n4335 = n4325 & n4333;
  assign n4336 = ~n4334 & ~n4335;
  assign n4337 = ~n4203 & n4228;
  assign n4338 = n4203 & ~n4228;
  assign n4339 = ~n4337 & ~n4338;
  assign n4340 = ~n4250 & ~n4339;
  assign n4341 = n4250 & n4339;
  assign n4342 = ~n4340 & ~n4341;
  assign n4343 = n4336 & n4342;
  assign n4344 = ~n4239 & n4242;
  assign n4345 = n4239 & ~n4242;
  assign n4346 = ~n4344 & ~n4345;
  assign n4347 = ~n4315 & n4318;
  assign n4348 = n4315 & ~n4318;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = ~n4346 & ~n4349;
  assign n4351 = ~n4234 & ~n4245;
  assign n4352 = ~n4248 & ~n4351;
  assign n4353 = ~n4231 & n4352;
  assign n4354 = n4231 & ~n4352;
  assign n4355 = ~n4353 & ~n4354;
  assign n4356 = n4350 & ~n4355;
  assign n4357 = ~n4322 & ~n4324;
  assign n4358 = n4307 & n4357;
  assign n4359 = ~n4307 & ~n4357;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = ~n4350 & n4355;
  assign n4362 = ~n4360 & ~n4361;
  assign n4363 = ~n4356 & ~n4362;
  assign n4364 = ~n4336 & ~n4342;
  assign n4365 = ~n4343 & ~n4364;
  assign n4366 = ~n4363 & n4365;
  assign n4367 = ~n4343 & ~n4366;
  assign n4368 = ~n4330 & ~n4367;
  assign n4369 = ~n4254 & ~n4329;
  assign n4370 = ~n4368 & ~n4369;
  assign n4371 = pi322  & pi323 ;
  assign n4372 = ~pi322  & pi323 ;
  assign n4373 = pi322  & ~pi323 ;
  assign n4374 = ~n4372 & ~n4373;
  assign n4375 = pi324  & ~n4374;
  assign n4376 = ~n4371 & ~n4375;
  assign n4377 = pi319  & pi320 ;
  assign n4378 = ~pi319  & pi320 ;
  assign n4379 = pi319  & ~pi320 ;
  assign n4380 = ~n4378 & ~n4379;
  assign n4381 = pi321  & ~n4380;
  assign n4382 = ~n4377 & ~n4381;
  assign n4383 = ~n4376 & n4382;
  assign n4384 = n4376 & ~n4382;
  assign n4385 = ~n4383 & ~n4384;
  assign n4386 = ~pi321  & ~n4380;
  assign n4387 = pi321  & n4380;
  assign n4388 = ~n4386 & ~n4387;
  assign n4389 = ~pi324  & ~n4374;
  assign n4390 = pi324  & n4374;
  assign n4391 = ~n4389 & ~n4390;
  assign n4392 = ~n4388 & ~n4391;
  assign n4393 = n4385 & n4392;
  assign n4394 = ~n4385 & ~n4392;
  assign n4395 = ~n4393 & ~n4394;
  assign n4396 = pi328  & pi329 ;
  assign n4397 = ~pi328  & pi329 ;
  assign n4398 = pi328  & ~pi329 ;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = pi330  & ~n4399;
  assign n4401 = ~n4396 & ~n4400;
  assign n4402 = pi325  & pi326 ;
  assign n4403 = ~pi325  & pi326 ;
  assign n4404 = pi325  & ~pi326 ;
  assign n4405 = ~n4403 & ~n4404;
  assign n4406 = pi327  & ~n4405;
  assign n4407 = ~n4402 & ~n4406;
  assign n4408 = ~n4401 & n4407;
  assign n4409 = n4401 & ~n4407;
  assign n4410 = ~n4408 & ~n4409;
  assign n4411 = ~pi327  & ~n4405;
  assign n4412 = pi327  & n4405;
  assign n4413 = ~n4411 & ~n4412;
  assign n4414 = ~pi330  & ~n4399;
  assign n4415 = pi330  & n4399;
  assign n4416 = ~n4414 & ~n4415;
  assign n4417 = ~n4413 & ~n4416;
  assign n4418 = n4410 & n4417;
  assign n4419 = ~n4410 & ~n4417;
  assign n4420 = ~n4418 & ~n4419;
  assign n4421 = ~n4410 & n4417;
  assign n4422 = ~n4401 & ~n4407;
  assign n4423 = ~n4421 & ~n4422;
  assign n4424 = ~n4420 & ~n4423;
  assign n4425 = ~n4385 & n4392;
  assign n4426 = ~n4376 & ~n4382;
  assign n4427 = ~n4425 & ~n4426;
  assign n4428 = ~n4395 & ~n4427;
  assign n4429 = ~n4413 & n4416;
  assign n4430 = n4413 & ~n4416;
  assign n4431 = ~n4429 & ~n4430;
  assign n4432 = ~n4388 & n4391;
  assign n4433 = n4388 & ~n4391;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = ~n4431 & ~n4434;
  assign n4436 = ~n4424 & n4435;
  assign n4437 = ~n4428 & n4436;
  assign n4438 = n4420 & ~n4437;
  assign n4439 = ~n4395 & ~n4438;
  assign n4440 = ~n4420 & n4437;
  assign n4441 = ~n4439 & ~n4440;
  assign n4442 = n4423 & ~n4427;
  assign n4443 = ~n4423 & n4427;
  assign n4444 = ~n4442 & ~n4443;
  assign n4445 = ~n4441 & ~n4444;
  assign n4446 = n4441 & n4444;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = pi331  & ~pi332 ;
  assign n4449 = ~pi331  & pi332 ;
  assign n4450 = ~n4448 & ~n4449;
  assign n4451 = ~pi333  & ~n4450;
  assign n4452 = pi333  & n4450;
  assign n4453 = ~n4451 & ~n4452;
  assign n4454 = pi334  & ~pi335 ;
  assign n4455 = ~pi334  & pi335 ;
  assign n4456 = ~n4454 & ~n4455;
  assign n4457 = ~pi336  & ~n4456;
  assign n4458 = pi336  & n4456;
  assign n4459 = ~n4457 & ~n4458;
  assign n4460 = ~n4453 & ~n4459;
  assign n4461 = pi334  & pi335 ;
  assign n4462 = pi336  & ~n4456;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = pi331  & pi332 ;
  assign n4465 = pi333  & ~n4450;
  assign n4466 = ~n4464 & ~n4465;
  assign n4467 = n4463 & ~n4466;
  assign n4468 = ~n4463 & n4466;
  assign n4469 = ~n4467 & ~n4468;
  assign n4470 = n4460 & n4469;
  assign n4471 = ~n4460 & ~n4469;
  assign n4472 = ~n4470 & ~n4471;
  assign n4473 = pi340  & pi341 ;
  assign n4474 = pi340  & ~pi341 ;
  assign n4475 = ~pi340  & pi341 ;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = pi342  & ~n4476;
  assign n4478 = ~n4473 & ~n4477;
  assign n4479 = pi337  & pi338 ;
  assign n4480 = pi337  & ~pi338 ;
  assign n4481 = ~pi337  & pi338 ;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = pi339  & ~n4482;
  assign n4484 = ~n4479 & ~n4483;
  assign n4485 = ~n4478 & n4484;
  assign n4486 = n4478 & ~n4484;
  assign n4487 = ~n4485 & ~n4486;
  assign n4488 = ~pi339  & ~n4482;
  assign n4489 = pi339  & n4482;
  assign n4490 = ~n4488 & ~n4489;
  assign n4491 = ~pi342  & ~n4476;
  assign n4492 = pi342  & n4476;
  assign n4493 = ~n4491 & ~n4492;
  assign n4494 = ~n4490 & ~n4493;
  assign n4495 = n4487 & n4494;
  assign n4496 = ~n4487 & ~n4494;
  assign n4497 = ~n4495 & ~n4496;
  assign n4498 = ~n4487 & n4494;
  assign n4499 = ~n4478 & ~n4484;
  assign n4500 = ~n4498 & ~n4499;
  assign n4501 = ~n4497 & ~n4500;
  assign n4502 = n4460 & ~n4469;
  assign n4503 = ~n4463 & ~n4466;
  assign n4504 = ~n4502 & ~n4503;
  assign n4505 = ~n4472 & ~n4504;
  assign n4506 = ~n4453 & n4459;
  assign n4507 = n4453 & ~n4459;
  assign n4508 = ~n4506 & ~n4507;
  assign n4509 = ~n4490 & n4493;
  assign n4510 = n4490 & ~n4493;
  assign n4511 = ~n4509 & ~n4510;
  assign n4512 = ~n4508 & ~n4511;
  assign n4513 = ~n4501 & n4512;
  assign n4514 = ~n4505 & n4513;
  assign n4515 = n4497 & ~n4514;
  assign n4516 = ~n4472 & ~n4515;
  assign n4517 = n4497 & n4514;
  assign n4518 = n4514 & ~n4517;
  assign n4519 = ~n4516 & ~n4518;
  assign n4520 = n4500 & ~n4504;
  assign n4521 = ~n4500 & n4504;
  assign n4522 = ~n4520 & ~n4521;
  assign n4523 = ~n4519 & ~n4522;
  assign n4524 = n4519 & n4522;
  assign n4525 = ~n4523 & ~n4524;
  assign n4526 = n4447 & n4525;
  assign n4527 = ~n4508 & n4511;
  assign n4528 = n4508 & ~n4511;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = n4431 & ~n4434;
  assign n4531 = ~n4431 & n4434;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = ~n4529 & ~n4532;
  assign n4534 = ~n4497 & ~n4514;
  assign n4535 = ~n4517 & ~n4534;
  assign n4536 = ~n4472 & n4535;
  assign n4537 = n4472 & ~n4535;
  assign n4538 = ~n4536 & ~n4537;
  assign n4539 = n4533 & ~n4538;
  assign n4540 = ~n4438 & ~n4440;
  assign n4541 = n4395 & n4540;
  assign n4542 = ~n4395 & ~n4540;
  assign n4543 = ~n4541 & ~n4542;
  assign n4544 = ~n4533 & n4538;
  assign n4545 = ~n4543 & ~n4544;
  assign n4546 = ~n4539 & ~n4545;
  assign n4547 = ~n4447 & ~n4525;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = ~n4526 & ~n4548;
  assign n4550 = n4500 & n4519;
  assign n4551 = ~n4504 & ~n4550;
  assign n4552 = ~n4500 & ~n4519;
  assign n4553 = ~n4551 & ~n4552;
  assign n4554 = n4423 & n4441;
  assign n4555 = ~n4427 & ~n4554;
  assign n4556 = ~n4423 & ~n4441;
  assign n4557 = ~n4555 & ~n4556;
  assign n4558 = n4553 & n4557;
  assign n4559 = ~n4549 & ~n4558;
  assign n4560 = ~n4553 & ~n4557;
  assign n4561 = ~n4559 & ~n4560;
  assign n4562 = ~n4370 & ~n4561;
  assign n4563 = ~n4346 & n4349;
  assign n4564 = n4346 & ~n4349;
  assign n4565 = ~n4563 & ~n4564;
  assign n4566 = ~n4529 & n4532;
  assign n4567 = n4529 & ~n4532;
  assign n4568 = ~n4566 & ~n4567;
  assign n4569 = ~n4565 & ~n4568;
  assign n4570 = ~n4356 & ~n4361;
  assign n4571 = ~n4360 & ~n4570;
  assign n4572 = n4360 & n4570;
  assign n4573 = ~n4571 & ~n4572;
  assign n4574 = n4569 & ~n4573;
  assign n4575 = ~n4539 & ~n4544;
  assign n4576 = n4543 & n4575;
  assign n4577 = ~n4543 & ~n4575;
  assign n4578 = ~n4576 & ~n4577;
  assign n4579 = ~n4569 & n4573;
  assign n4580 = ~n4578 & ~n4579;
  assign n4581 = ~n4574 & ~n4580;
  assign n4582 = ~n4526 & ~n4547;
  assign n4583 = ~n4546 & n4582;
  assign n4584 = n4546 & ~n4582;
  assign n4585 = ~n4583 & ~n4584;
  assign n4586 = n4363 & ~n4365;
  assign n4587 = ~n4366 & ~n4586;
  assign n4588 = ~n4585 & ~n4587;
  assign n4589 = ~n4581 & ~n4588;
  assign n4590 = n4585 & n4587;
  assign n4591 = ~n4589 & ~n4590;
  assign n4592 = ~n4330 & ~n4369;
  assign n4593 = ~n4367 & n4592;
  assign n4594 = n4367 & ~n4592;
  assign n4595 = ~n4593 & ~n4594;
  assign n4596 = n4553 & ~n4557;
  assign n4597 = ~n4553 & n4557;
  assign n4598 = ~n4526 & ~n4596;
  assign n4599 = ~n4597 & n4598;
  assign n4600 = ~n4548 & n4599;
  assign n4601 = n4559 & ~n4560;
  assign n4602 = ~n4600 & ~n4601;
  assign n4603 = ~n4595 & ~n4602;
  assign n4604 = ~n4591 & ~n4603;
  assign n4605 = n4595 & n4602;
  assign n4606 = ~n4604 & ~n4605;
  assign n4607 = n4370 & n4561;
  assign n4608 = ~n4562 & ~n4607;
  assign n4609 = ~n4606 & n4608;
  assign n4610 = ~n4562 & ~n4609;
  assign n4611 = pi310  & pi311 ;
  assign n4612 = ~pi310  & pi311 ;
  assign n4613 = pi310  & ~pi311 ;
  assign n4614 = ~n4612 & ~n4613;
  assign n4615 = pi312  & ~n4614;
  assign n4616 = ~n4611 & ~n4615;
  assign n4617 = pi307  & pi308 ;
  assign n4618 = ~pi307  & pi308 ;
  assign n4619 = pi307  & ~pi308 ;
  assign n4620 = ~n4618 & ~n4619;
  assign n4621 = pi309  & ~n4620;
  assign n4622 = ~n4617 & ~n4621;
  assign n4623 = ~n4616 & n4622;
  assign n4624 = n4616 & ~n4622;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = ~pi309  & ~n4620;
  assign n4627 = pi309  & n4620;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = ~pi312  & ~n4614;
  assign n4630 = pi312  & n4614;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = ~n4628 & ~n4631;
  assign n4633 = ~n4625 & n4632;
  assign n4634 = ~n4616 & ~n4622;
  assign n4635 = ~n4633 & ~n4634;
  assign n4636 = pi316  & pi317 ;
  assign n4637 = ~pi316  & pi317 ;
  assign n4638 = pi316  & ~pi317 ;
  assign n4639 = ~n4637 & ~n4638;
  assign n4640 = pi318  & ~n4639;
  assign n4641 = ~n4636 & ~n4640;
  assign n4642 = pi313  & pi314 ;
  assign n4643 = ~pi313  & pi314 ;
  assign n4644 = pi313  & ~pi314 ;
  assign n4645 = ~n4643 & ~n4644;
  assign n4646 = pi315  & ~n4645;
  assign n4647 = ~n4642 & ~n4646;
  assign n4648 = ~n4641 & n4647;
  assign n4649 = n4641 & ~n4647;
  assign n4650 = ~n4648 & ~n4649;
  assign n4651 = ~pi315  & ~n4645;
  assign n4652 = pi315  & n4645;
  assign n4653 = ~n4651 & ~n4652;
  assign n4654 = ~pi318  & ~n4639;
  assign n4655 = pi318  & n4639;
  assign n4656 = ~n4654 & ~n4655;
  assign n4657 = ~n4653 & ~n4656;
  assign n4658 = ~n4650 & n4657;
  assign n4659 = ~n4641 & ~n4647;
  assign n4660 = ~n4658 & ~n4659;
  assign n4661 = n4650 & n4657;
  assign n4662 = ~n4650 & ~n4657;
  assign n4663 = ~n4661 & ~n4662;
  assign n4664 = ~n4660 & ~n4663;
  assign n4665 = n4625 & n4632;
  assign n4666 = ~n4625 & ~n4632;
  assign n4667 = ~n4665 & ~n4666;
  assign n4668 = ~n4635 & ~n4667;
  assign n4669 = ~n4653 & n4656;
  assign n4670 = n4653 & ~n4656;
  assign n4671 = ~n4669 & ~n4670;
  assign n4672 = ~n4628 & n4631;
  assign n4673 = n4628 & ~n4631;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = ~n4671 & ~n4674;
  assign n4676 = ~n4664 & n4675;
  assign n4677 = ~n4668 & n4676;
  assign n4678 = ~n4663 & n4677;
  assign n4679 = n4663 & ~n4677;
  assign n4680 = ~n4667 & ~n4679;
  assign n4681 = ~n4678 & ~n4680;
  assign n4682 = n4660 & n4681;
  assign n4683 = ~n4635 & ~n4682;
  assign n4684 = ~n4660 & ~n4681;
  assign n4685 = ~n4683 & ~n4684;
  assign n4686 = pi298  & pi299 ;
  assign n4687 = ~pi298  & pi299 ;
  assign n4688 = pi298  & ~pi299 ;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = pi300  & ~n4689;
  assign n4691 = ~n4686 & ~n4690;
  assign n4692 = pi295  & pi296 ;
  assign n4693 = ~pi295  & pi296 ;
  assign n4694 = pi295  & ~pi296 ;
  assign n4695 = ~n4693 & ~n4694;
  assign n4696 = pi297  & ~n4695;
  assign n4697 = ~n4692 & ~n4696;
  assign n4698 = ~n4691 & n4697;
  assign n4699 = n4691 & ~n4697;
  assign n4700 = ~n4698 & ~n4699;
  assign n4701 = ~pi297  & ~n4695;
  assign n4702 = pi297  & n4695;
  assign n4703 = ~n4701 & ~n4702;
  assign n4704 = ~pi300  & ~n4689;
  assign n4705 = pi300  & n4689;
  assign n4706 = ~n4704 & ~n4705;
  assign n4707 = ~n4703 & ~n4706;
  assign n4708 = ~n4700 & n4707;
  assign n4709 = ~n4691 & ~n4697;
  assign n4710 = ~n4708 & ~n4709;
  assign n4711 = pi304  & pi305 ;
  assign n4712 = ~pi304  & pi305 ;
  assign n4713 = pi304  & ~pi305 ;
  assign n4714 = ~n4712 & ~n4713;
  assign n4715 = pi306  & ~n4714;
  assign n4716 = ~n4711 & ~n4715;
  assign n4717 = pi301  & pi302 ;
  assign n4718 = ~pi301  & pi302 ;
  assign n4719 = pi301  & ~pi302 ;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = pi303  & ~n4720;
  assign n4722 = ~n4717 & ~n4721;
  assign n4723 = ~n4716 & n4722;
  assign n4724 = n4716 & ~n4722;
  assign n4725 = ~n4723 & ~n4724;
  assign n4726 = ~pi303  & ~n4720;
  assign n4727 = pi303  & n4720;
  assign n4728 = ~n4726 & ~n4727;
  assign n4729 = ~pi306  & ~n4714;
  assign n4730 = pi306  & n4714;
  assign n4731 = ~n4729 & ~n4730;
  assign n4732 = ~n4728 & ~n4731;
  assign n4733 = ~n4725 & n4732;
  assign n4734 = ~n4716 & ~n4722;
  assign n4735 = ~n4733 & ~n4734;
  assign n4736 = n4725 & n4732;
  assign n4737 = ~n4725 & ~n4732;
  assign n4738 = ~n4736 & ~n4737;
  assign n4739 = ~n4735 & ~n4738;
  assign n4740 = n4700 & n4707;
  assign n4741 = ~n4700 & ~n4707;
  assign n4742 = ~n4740 & ~n4741;
  assign n4743 = ~n4710 & ~n4742;
  assign n4744 = ~n4728 & n4731;
  assign n4745 = n4728 & ~n4731;
  assign n4746 = ~n4744 & ~n4745;
  assign n4747 = ~n4703 & n4706;
  assign n4748 = n4703 & ~n4706;
  assign n4749 = ~n4747 & ~n4748;
  assign n4750 = ~n4746 & ~n4749;
  assign n4751 = ~n4739 & n4750;
  assign n4752 = ~n4743 & n4751;
  assign n4753 = ~n4738 & n4752;
  assign n4754 = n4738 & ~n4752;
  assign n4755 = ~n4742 & ~n4754;
  assign n4756 = ~n4753 & ~n4755;
  assign n4757 = n4735 & n4756;
  assign n4758 = ~n4710 & ~n4757;
  assign n4759 = ~n4735 & ~n4756;
  assign n4760 = ~n4758 & ~n4759;
  assign n4761 = n4685 & n4760;
  assign n4762 = ~n4710 & n4735;
  assign n4763 = n4710 & ~n4735;
  assign n4764 = ~n4762 & ~n4763;
  assign n4765 = ~n4756 & ~n4764;
  assign n4766 = n4756 & n4764;
  assign n4767 = ~n4765 & ~n4766;
  assign n4768 = ~n4635 & n4660;
  assign n4769 = n4635 & ~n4660;
  assign n4770 = ~n4768 & ~n4769;
  assign n4771 = ~n4681 & ~n4770;
  assign n4772 = n4681 & n4770;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = n4767 & n4773;
  assign n4775 = n4671 & ~n4674;
  assign n4776 = ~n4671 & n4674;
  assign n4777 = ~n4775 & ~n4776;
  assign n4778 = n4746 & ~n4749;
  assign n4779 = ~n4746 & n4749;
  assign n4780 = ~n4778 & ~n4779;
  assign n4781 = ~n4777 & ~n4780;
  assign n4782 = ~n4678 & ~n4679;
  assign n4783 = ~n4667 & ~n4782;
  assign n4784 = n4667 & n4782;
  assign n4785 = ~n4783 & ~n4784;
  assign n4786 = n4781 & ~n4785;
  assign n4787 = ~n4753 & ~n4754;
  assign n4788 = n4742 & n4787;
  assign n4789 = ~n4742 & ~n4787;
  assign n4790 = ~n4788 & ~n4789;
  assign n4791 = ~n4781 & n4785;
  assign n4792 = ~n4790 & ~n4791;
  assign n4793 = ~n4786 & ~n4792;
  assign n4794 = ~n4767 & ~n4773;
  assign n4795 = ~n4774 & ~n4794;
  assign n4796 = ~n4793 & n4795;
  assign n4797 = ~n4774 & ~n4796;
  assign n4798 = ~n4761 & ~n4797;
  assign n4799 = ~n4685 & ~n4760;
  assign n4800 = ~n4798 & ~n4799;
  assign n4801 = ~pi289  & pi290 ;
  assign n4802 = pi289  & ~pi290 ;
  assign n4803 = ~n4801 & ~n4802;
  assign n4804 = ~pi291  & ~n4803;
  assign n4805 = pi291  & n4803;
  assign n4806 = ~n4804 & ~n4805;
  assign n4807 = ~pi292  & pi293 ;
  assign n4808 = pi292  & ~pi293 ;
  assign n4809 = ~n4807 & ~n4808;
  assign n4810 = ~pi294  & ~n4809;
  assign n4811 = pi294  & n4809;
  assign n4812 = ~n4810 & ~n4811;
  assign n4813 = ~n4806 & n4812;
  assign n4814 = n4806 & ~n4812;
  assign n4815 = ~n4813 & ~n4814;
  assign n4816 = ~pi283  & pi284 ;
  assign n4817 = pi283  & ~pi284 ;
  assign n4818 = ~n4816 & ~n4817;
  assign n4819 = ~pi285  & ~n4818;
  assign n4820 = pi285  & n4818;
  assign n4821 = ~n4819 & ~n4820;
  assign n4822 = ~pi286  & pi287 ;
  assign n4823 = pi286  & ~pi287 ;
  assign n4824 = ~n4822 & ~n4823;
  assign n4825 = ~pi288  & ~n4824;
  assign n4826 = pi288  & n4824;
  assign n4827 = ~n4825 & ~n4826;
  assign n4828 = ~n4821 & n4827;
  assign n4829 = n4821 & ~n4827;
  assign n4830 = ~n4828 & ~n4829;
  assign n4831 = n4815 & ~n4830;
  assign n4832 = ~n4815 & n4830;
  assign n4833 = ~n4831 & ~n4832;
  assign n4834 = ~pi277  & pi278 ;
  assign n4835 = pi277  & ~pi278 ;
  assign n4836 = ~n4834 & ~n4835;
  assign n4837 = ~pi279  & ~n4836;
  assign n4838 = pi279  & n4836;
  assign n4839 = ~n4837 & ~n4838;
  assign n4840 = ~pi280  & pi281 ;
  assign n4841 = pi280  & ~pi281 ;
  assign n4842 = ~n4840 & ~n4841;
  assign n4843 = ~pi282  & ~n4842;
  assign n4844 = pi282  & n4842;
  assign n4845 = ~n4843 & ~n4844;
  assign n4846 = ~n4839 & n4845;
  assign n4847 = n4839 & ~n4845;
  assign n4848 = ~n4846 & ~n4847;
  assign n4849 = ~pi271  & pi272 ;
  assign n4850 = pi271  & ~pi272 ;
  assign n4851 = ~n4849 & ~n4850;
  assign n4852 = ~pi273  & ~n4851;
  assign n4853 = pi273  & n4851;
  assign n4854 = ~n4852 & ~n4853;
  assign n4855 = ~pi274  & pi275 ;
  assign n4856 = pi274  & ~pi275 ;
  assign n4857 = ~n4855 & ~n4856;
  assign n4858 = ~pi276  & ~n4857;
  assign n4859 = pi276  & n4857;
  assign n4860 = ~n4858 & ~n4859;
  assign n4861 = ~n4854 & n4860;
  assign n4862 = n4854 & ~n4860;
  assign n4863 = ~n4861 & ~n4862;
  assign n4864 = n4848 & ~n4863;
  assign n4865 = ~n4848 & n4863;
  assign n4866 = ~n4864 & ~n4865;
  assign n4867 = ~n4833 & ~n4866;
  assign n4868 = pi286  & pi287 ;
  assign n4869 = pi288  & ~n4824;
  assign n4870 = ~n4868 & ~n4869;
  assign n4871 = pi283  & pi284 ;
  assign n4872 = pi285  & ~n4818;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = ~n4870 & n4873;
  assign n4875 = n4870 & ~n4873;
  assign n4876 = ~n4874 & ~n4875;
  assign n4877 = ~n4821 & ~n4827;
  assign n4878 = n4876 & n4877;
  assign n4879 = ~n4876 & ~n4877;
  assign n4880 = ~n4878 & ~n4879;
  assign n4881 = pi292  & pi293 ;
  assign n4882 = pi294  & ~n4809;
  assign n4883 = ~n4881 & ~n4882;
  assign n4884 = pi289  & pi290 ;
  assign n4885 = pi291  & ~n4803;
  assign n4886 = ~n4884 & ~n4885;
  assign n4887 = ~n4883 & n4886;
  assign n4888 = n4883 & ~n4886;
  assign n4889 = ~n4887 & ~n4888;
  assign n4890 = ~n4806 & ~n4812;
  assign n4891 = n4889 & n4890;
  assign n4892 = ~n4889 & ~n4890;
  assign n4893 = ~n4891 & ~n4892;
  assign n4894 = ~n4889 & n4890;
  assign n4895 = ~n4883 & ~n4886;
  assign n4896 = ~n4894 & ~n4895;
  assign n4897 = ~n4893 & ~n4896;
  assign n4898 = ~n4876 & n4877;
  assign n4899 = ~n4870 & ~n4873;
  assign n4900 = ~n4898 & ~n4899;
  assign n4901 = ~n4880 & ~n4900;
  assign n4902 = ~n4815 & ~n4830;
  assign n4903 = ~n4897 & n4902;
  assign n4904 = ~n4901 & n4903;
  assign n4905 = n4893 & ~n4904;
  assign n4906 = ~n4893 & n4904;
  assign n4907 = ~n4905 & ~n4906;
  assign n4908 = ~n4880 & ~n4907;
  assign n4909 = n4880 & n4907;
  assign n4910 = ~n4908 & ~n4909;
  assign n4911 = n4867 & ~n4910;
  assign n4912 = pi274  & pi275 ;
  assign n4913 = pi276  & ~n4857;
  assign n4914 = ~n4912 & ~n4913;
  assign n4915 = pi271  & pi272 ;
  assign n4916 = pi273  & ~n4851;
  assign n4917 = ~n4915 & ~n4916;
  assign n4918 = ~n4914 & n4917;
  assign n4919 = n4914 & ~n4917;
  assign n4920 = ~n4918 & ~n4919;
  assign n4921 = ~n4854 & ~n4860;
  assign n4922 = n4920 & n4921;
  assign n4923 = ~n4920 & ~n4921;
  assign n4924 = ~n4922 & ~n4923;
  assign n4925 = pi280  & pi281 ;
  assign n4926 = pi282  & ~n4842;
  assign n4927 = ~n4925 & ~n4926;
  assign n4928 = pi277  & pi278 ;
  assign n4929 = pi279  & ~n4836;
  assign n4930 = ~n4928 & ~n4929;
  assign n4931 = ~n4927 & n4930;
  assign n4932 = n4927 & ~n4930;
  assign n4933 = ~n4931 & ~n4932;
  assign n4934 = ~n4839 & ~n4845;
  assign n4935 = n4933 & n4934;
  assign n4936 = ~n4933 & ~n4934;
  assign n4937 = ~n4935 & ~n4936;
  assign n4938 = ~n4933 & n4934;
  assign n4939 = ~n4927 & ~n4930;
  assign n4940 = ~n4938 & ~n4939;
  assign n4941 = ~n4937 & ~n4940;
  assign n4942 = ~n4920 & n4921;
  assign n4943 = ~n4914 & ~n4917;
  assign n4944 = ~n4942 & ~n4943;
  assign n4945 = ~n4924 & ~n4944;
  assign n4946 = ~n4848 & ~n4863;
  assign n4947 = ~n4941 & n4946;
  assign n4948 = ~n4945 & n4947;
  assign n4949 = n4937 & ~n4948;
  assign n4950 = ~n4937 & n4948;
  assign n4951 = ~n4949 & ~n4950;
  assign n4952 = n4924 & n4951;
  assign n4953 = ~n4924 & ~n4951;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = ~n4867 & n4910;
  assign n4956 = ~n4954 & ~n4955;
  assign n4957 = ~n4911 & ~n4956;
  assign n4958 = ~n4924 & ~n4949;
  assign n4959 = ~n4950 & ~n4958;
  assign n4960 = n4940 & ~n4944;
  assign n4961 = ~n4940 & n4944;
  assign n4962 = ~n4960 & ~n4961;
  assign n4963 = ~n4959 & ~n4962;
  assign n4964 = n4959 & n4962;
  assign n4965 = ~n4963 & ~n4964;
  assign n4966 = ~n4880 & ~n4905;
  assign n4967 = ~n4906 & ~n4966;
  assign n4968 = n4896 & ~n4900;
  assign n4969 = ~n4896 & n4900;
  assign n4970 = ~n4968 & ~n4969;
  assign n4971 = ~n4967 & ~n4970;
  assign n4972 = n4967 & n4970;
  assign n4973 = ~n4971 & ~n4972;
  assign n4974 = ~n4965 & ~n4973;
  assign n4975 = ~n4957 & ~n4974;
  assign n4976 = n4965 & n4973;
  assign n4977 = ~n4975 & ~n4976;
  assign n4978 = n4896 & n4967;
  assign n4979 = ~n4900 & ~n4978;
  assign n4980 = ~n4896 & ~n4967;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = n4940 & n4959;
  assign n4983 = ~n4944 & ~n4982;
  assign n4984 = ~n4940 & ~n4959;
  assign n4985 = ~n4983 & ~n4984;
  assign n4986 = n4981 & n4985;
  assign n4987 = ~n4977 & ~n4986;
  assign n4988 = ~n4981 & ~n4985;
  assign n4989 = ~n4987 & ~n4988;
  assign n4990 = ~n4800 & ~n4989;
  assign n4991 = ~n4974 & ~n4976;
  assign n4992 = ~n4957 & n4991;
  assign n4993 = n4957 & ~n4991;
  assign n4994 = ~n4992 & ~n4993;
  assign n4995 = n4793 & ~n4795;
  assign n4996 = ~n4796 & ~n4995;
  assign n4997 = n4994 & n4996;
  assign n4998 = ~n4777 & n4780;
  assign n4999 = n4777 & ~n4780;
  assign n5000 = ~n4998 & ~n4999;
  assign n5001 = ~n4833 & n4866;
  assign n5002 = n4833 & ~n4866;
  assign n5003 = ~n5001 & ~n5002;
  assign n5004 = ~n5000 & ~n5003;
  assign n5005 = ~n4786 & ~n4791;
  assign n5006 = ~n4790 & ~n5005;
  assign n5007 = n4790 & n5005;
  assign n5008 = ~n5006 & ~n5007;
  assign n5009 = n5004 & ~n5008;
  assign n5010 = ~n4911 & ~n4955;
  assign n5011 = n4954 & n5010;
  assign n5012 = ~n4954 & ~n5010;
  assign n5013 = ~n5011 & ~n5012;
  assign n5014 = ~n5004 & n5008;
  assign n5015 = ~n5013 & ~n5014;
  assign n5016 = ~n5009 & ~n5015;
  assign n5017 = ~n4994 & ~n4996;
  assign n5018 = ~n4997 & ~n5017;
  assign n5019 = ~n5016 & n5018;
  assign n5020 = ~n4997 & ~n5019;
  assign n5021 = ~n4761 & ~n4799;
  assign n5022 = ~n4797 & n5021;
  assign n5023 = n4797 & ~n5021;
  assign n5024 = ~n5022 & ~n5023;
  assign n5025 = n4981 & ~n4985;
  assign n5026 = ~n4981 & n4985;
  assign n5027 = ~n4976 & ~n5025;
  assign n5028 = ~n5026 & n5027;
  assign n5029 = ~n4975 & n5028;
  assign n5030 = n4987 & ~n4988;
  assign n5031 = ~n5029 & ~n5030;
  assign n5032 = ~n5024 & ~n5031;
  assign n5033 = ~n5020 & ~n5032;
  assign n5034 = n5024 & n5031;
  assign n5035 = ~n5033 & ~n5034;
  assign n5036 = n4800 & n4989;
  assign n5037 = ~n4990 & ~n5036;
  assign n5038 = ~n5035 & n5037;
  assign n5039 = ~n4990 & ~n5038;
  assign n5040 = ~n4610 & ~n5039;
  assign n5041 = n4610 & n5039;
  assign n5042 = ~n5040 & ~n5041;
  assign n5043 = n5035 & ~n5037;
  assign n5044 = ~n5038 & ~n5043;
  assign n5045 = n4606 & ~n4608;
  assign n5046 = ~n4609 & ~n5045;
  assign n5047 = n5044 & n5046;
  assign n5048 = n5016 & ~n5018;
  assign n5049 = ~n5019 & ~n5048;
  assign n5050 = ~n4588 & ~n4590;
  assign n5051 = ~n4581 & n5050;
  assign n5052 = n4581 & ~n5050;
  assign n5053 = ~n5051 & ~n5052;
  assign n5054 = n5049 & n5053;
  assign n5055 = ~n4565 & n4568;
  assign n5056 = n4565 & ~n4568;
  assign n5057 = ~n5055 & ~n5056;
  assign n5058 = ~n5000 & n5003;
  assign n5059 = n5000 & ~n5003;
  assign n5060 = ~n5058 & ~n5059;
  assign n5061 = ~n5057 & ~n5060;
  assign n5062 = ~n4574 & ~n4579;
  assign n5063 = ~n4578 & ~n5062;
  assign n5064 = n4578 & n5062;
  assign n5065 = ~n5063 & ~n5064;
  assign n5066 = n5061 & ~n5065;
  assign n5067 = ~n5009 & ~n5014;
  assign n5068 = n5013 & n5067;
  assign n5069 = ~n5013 & ~n5067;
  assign n5070 = ~n5068 & ~n5069;
  assign n5071 = ~n5061 & n5065;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = ~n5066 & ~n5072;
  assign n5074 = ~n5049 & ~n5053;
  assign n5075 = ~n5054 & ~n5074;
  assign n5076 = ~n5073 & n5075;
  assign n5077 = ~n5054 & ~n5076;
  assign n5078 = ~n4603 & ~n4605;
  assign n5079 = ~n4591 & n5078;
  assign n5080 = n4591 & ~n5078;
  assign n5081 = ~n5079 & ~n5080;
  assign n5082 = ~n5032 & ~n5034;
  assign n5083 = ~n5020 & n5082;
  assign n5084 = n5020 & ~n5082;
  assign n5085 = ~n5083 & ~n5084;
  assign n5086 = ~n5081 & ~n5085;
  assign n5087 = ~n5077 & ~n5086;
  assign n5088 = n5081 & n5085;
  assign n5089 = ~n5087 & ~n5088;
  assign n5090 = ~n5044 & ~n5046;
  assign n5091 = ~n5047 & ~n5090;
  assign n5092 = ~n5089 & n5091;
  assign n5093 = ~n5047 & ~n5092;
  assign n5094 = n5042 & ~n5093;
  assign n5095 = ~n5040 & ~n5094;
  assign n5096 = ~n4178 & ~n5095;
  assign n5097 = n4178 & n5095;
  assign n5098 = ~n5096 & ~n5097;
  assign n5099 = ~n4125 & n4176;
  assign n5100 = ~n4177 & ~n5099;
  assign n5101 = ~n5042 & n5093;
  assign n5102 = ~n5094 & ~n5101;
  assign n5103 = n5100 & n5102;
  assign n5104 = ~n4169 & ~n4171;
  assign n5105 = ~n4160 & n5104;
  assign n5106 = n4160 & ~n5104;
  assign n5107 = ~n5105 & ~n5106;
  assign n5108 = ~n5086 & ~n5088;
  assign n5109 = ~n5077 & n5108;
  assign n5110 = n5077 & ~n5108;
  assign n5111 = ~n5109 & ~n5110;
  assign n5112 = n5107 & n5111;
  assign n5113 = ~n4140 & n4143;
  assign n5114 = n4140 & ~n4143;
  assign n5115 = ~n5113 & ~n5114;
  assign n5116 = ~n5057 & n5060;
  assign n5117 = n5057 & ~n5060;
  assign n5118 = ~n5116 & ~n5117;
  assign n5119 = ~n5115 & ~n5118;
  assign n5120 = ~n4149 & ~n4154;
  assign n5121 = n4153 & n5120;
  assign n5122 = ~n4153 & ~n5120;
  assign n5123 = ~n5121 & ~n5122;
  assign n5124 = n5119 & ~n5123;
  assign n5125 = ~n5066 & ~n5071;
  assign n5126 = n5070 & n5125;
  assign n5127 = ~n5070 & ~n5125;
  assign n5128 = ~n5126 & ~n5127;
  assign n5129 = ~n5119 & n5123;
  assign n5130 = ~n5128 & ~n5129;
  assign n5131 = ~n5124 & ~n5130;
  assign n5132 = n5073 & ~n5075;
  assign n5133 = ~n5076 & ~n5132;
  assign n5134 = n4156 & ~n4158;
  assign n5135 = ~n4159 & ~n5134;
  assign n5136 = ~n5133 & ~n5135;
  assign n5137 = ~n5131 & ~n5136;
  assign n5138 = n5133 & n5135;
  assign n5139 = ~n5137 & ~n5138;
  assign n5140 = ~n5107 & ~n5111;
  assign n5141 = ~n5139 & ~n5140;
  assign n5142 = ~n5112 & ~n5141;
  assign n5143 = n5089 & ~n5091;
  assign n5144 = ~n5092 & ~n5143;
  assign n5145 = n4172 & ~n4174;
  assign n5146 = ~n4175 & ~n5145;
  assign n5147 = ~n5144 & ~n5146;
  assign n5148 = ~n5142 & ~n5147;
  assign n5149 = n5144 & n5146;
  assign n5150 = ~n5148 & ~n5149;
  assign n5151 = ~n5100 & ~n5102;
  assign n5152 = ~n5103 & ~n5151;
  assign n5153 = ~n5150 & n5152;
  assign n5154 = ~n5103 & ~n5153;
  assign n5155 = n5098 & ~n5154;
  assign n5156 = ~n5096 & ~n5155;
  assign n5157 = pi259  & ~pi260 ;
  assign n5158 = ~pi259  & pi260 ;
  assign n5159 = ~n5157 & ~n5158;
  assign n5160 = ~pi261  & ~n5159;
  assign n5161 = pi261  & n5159;
  assign n5162 = ~n5160 & ~n5161;
  assign n5163 = pi262  & ~pi263 ;
  assign n5164 = ~pi262  & pi263 ;
  assign n5165 = ~n5163 & ~n5164;
  assign n5166 = ~pi264  & ~n5165;
  assign n5167 = pi264  & n5165;
  assign n5168 = ~n5166 & ~n5167;
  assign n5169 = ~n5162 & ~n5168;
  assign n5170 = pi262  & pi263 ;
  assign n5171 = pi264  & ~n5165;
  assign n5172 = ~n5170 & ~n5171;
  assign n5173 = pi259  & pi260 ;
  assign n5174 = pi261  & ~n5159;
  assign n5175 = ~n5173 & ~n5174;
  assign n5176 = n5172 & ~n5175;
  assign n5177 = ~n5172 & n5175;
  assign n5178 = ~n5176 & ~n5177;
  assign n5179 = n5169 & ~n5178;
  assign n5180 = ~n5172 & ~n5175;
  assign n5181 = ~n5179 & ~n5180;
  assign n5182 = pi268  & pi269 ;
  assign n5183 = pi268  & ~pi269 ;
  assign n5184 = ~pi268  & pi269 ;
  assign n5185 = ~n5183 & ~n5184;
  assign n5186 = pi270  & ~n5185;
  assign n5187 = ~n5182 & ~n5186;
  assign n5188 = pi265  & pi266 ;
  assign n5189 = pi265  & ~pi266 ;
  assign n5190 = ~pi265  & pi266 ;
  assign n5191 = ~n5189 & ~n5190;
  assign n5192 = pi267  & ~n5191;
  assign n5193 = ~n5188 & ~n5192;
  assign n5194 = ~n5187 & n5193;
  assign n5195 = n5187 & ~n5193;
  assign n5196 = ~n5194 & ~n5195;
  assign n5197 = ~pi267  & ~n5191;
  assign n5198 = pi267  & n5191;
  assign n5199 = ~n5197 & ~n5198;
  assign n5200 = ~pi270  & ~n5185;
  assign n5201 = pi270  & n5185;
  assign n5202 = ~n5200 & ~n5201;
  assign n5203 = ~n5199 & ~n5202;
  assign n5204 = ~n5196 & n5203;
  assign n5205 = ~n5187 & ~n5193;
  assign n5206 = ~n5204 & ~n5205;
  assign n5207 = n5169 & n5178;
  assign n5208 = ~n5169 & ~n5178;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = n5196 & n5203;
  assign n5211 = ~n5196 & ~n5203;
  assign n5212 = ~n5210 & ~n5211;
  assign n5213 = ~n5206 & ~n5212;
  assign n5214 = ~n5181 & ~n5209;
  assign n5215 = ~n5162 & n5168;
  assign n5216 = n5162 & ~n5168;
  assign n5217 = ~n5215 & ~n5216;
  assign n5218 = ~n5199 & n5202;
  assign n5219 = n5199 & ~n5202;
  assign n5220 = ~n5218 & ~n5219;
  assign n5221 = ~n5217 & ~n5220;
  assign n5222 = ~n5213 & n5221;
  assign n5223 = ~n5214 & n5222;
  assign n5224 = n5212 & ~n5223;
  assign n5225 = ~n5209 & ~n5224;
  assign n5226 = n5212 & n5223;
  assign n5227 = n5223 & ~n5226;
  assign n5228 = ~n5225 & ~n5227;
  assign n5229 = n5206 & n5228;
  assign n5230 = ~n5181 & ~n5229;
  assign n5231 = ~n5206 & ~n5228;
  assign n5232 = ~n5230 & ~n5231;
  assign n5233 = pi247  & ~pi248 ;
  assign n5234 = ~pi247  & pi248 ;
  assign n5235 = ~n5233 & ~n5234;
  assign n5236 = ~pi249  & ~n5235;
  assign n5237 = pi249  & n5235;
  assign n5238 = ~n5236 & ~n5237;
  assign n5239 = pi250  & ~pi251 ;
  assign n5240 = ~pi250  & pi251 ;
  assign n5241 = ~n5239 & ~n5240;
  assign n5242 = ~pi252  & ~n5241;
  assign n5243 = pi252  & n5241;
  assign n5244 = ~n5242 & ~n5243;
  assign n5245 = ~n5238 & ~n5244;
  assign n5246 = pi250  & pi251 ;
  assign n5247 = pi252  & ~n5241;
  assign n5248 = ~n5246 & ~n5247;
  assign n5249 = pi247  & pi248 ;
  assign n5250 = pi249  & ~n5235;
  assign n5251 = ~n5249 & ~n5250;
  assign n5252 = n5248 & ~n5251;
  assign n5253 = ~n5248 & n5251;
  assign n5254 = ~n5252 & ~n5253;
  assign n5255 = n5245 & ~n5254;
  assign n5256 = ~n5248 & ~n5251;
  assign n5257 = ~n5255 & ~n5256;
  assign n5258 = pi256  & pi257 ;
  assign n5259 = pi256  & ~pi257 ;
  assign n5260 = ~pi256  & pi257 ;
  assign n5261 = ~n5259 & ~n5260;
  assign n5262 = pi258  & ~n5261;
  assign n5263 = ~n5258 & ~n5262;
  assign n5264 = pi253  & pi254 ;
  assign n5265 = pi253  & ~pi254 ;
  assign n5266 = ~pi253  & pi254 ;
  assign n5267 = ~n5265 & ~n5266;
  assign n5268 = pi255  & ~n5267;
  assign n5269 = ~n5264 & ~n5268;
  assign n5270 = ~n5263 & n5269;
  assign n5271 = n5263 & ~n5269;
  assign n5272 = ~n5270 & ~n5271;
  assign n5273 = ~pi255  & ~n5267;
  assign n5274 = pi255  & n5267;
  assign n5275 = ~n5273 & ~n5274;
  assign n5276 = ~pi258  & ~n5261;
  assign n5277 = pi258  & n5261;
  assign n5278 = ~n5276 & ~n5277;
  assign n5279 = ~n5275 & ~n5278;
  assign n5280 = ~n5272 & n5279;
  assign n5281 = ~n5263 & ~n5269;
  assign n5282 = ~n5280 & ~n5281;
  assign n5283 = n5245 & n5254;
  assign n5284 = ~n5245 & ~n5254;
  assign n5285 = ~n5283 & ~n5284;
  assign n5286 = n5272 & n5279;
  assign n5287 = ~n5272 & ~n5279;
  assign n5288 = ~n5286 & ~n5287;
  assign n5289 = ~n5282 & ~n5288;
  assign n5290 = ~n5257 & ~n5285;
  assign n5291 = ~n5238 & n5244;
  assign n5292 = n5238 & ~n5244;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = ~n5275 & n5278;
  assign n5295 = n5275 & ~n5278;
  assign n5296 = ~n5294 & ~n5295;
  assign n5297 = ~n5293 & ~n5296;
  assign n5298 = ~n5289 & n5297;
  assign n5299 = ~n5290 & n5298;
  assign n5300 = n5288 & ~n5299;
  assign n5301 = ~n5285 & ~n5300;
  assign n5302 = ~n5288 & n5299;
  assign n5303 = ~n5301 & ~n5302;
  assign n5304 = n5282 & n5303;
  assign n5305 = ~n5257 & ~n5304;
  assign n5306 = ~n5282 & ~n5303;
  assign n5307 = ~n5305 & ~n5306;
  assign n5308 = n5232 & n5307;
  assign n5309 = ~n5257 & n5282;
  assign n5310 = n5257 & ~n5282;
  assign n5311 = ~n5309 & ~n5310;
  assign n5312 = ~n5303 & ~n5311;
  assign n5313 = n5303 & n5311;
  assign n5314 = ~n5312 & ~n5313;
  assign n5315 = ~n5181 & n5206;
  assign n5316 = n5181 & ~n5206;
  assign n5317 = ~n5315 & ~n5316;
  assign n5318 = ~n5228 & ~n5317;
  assign n5319 = n5228 & n5317;
  assign n5320 = ~n5318 & ~n5319;
  assign n5321 = n5314 & n5320;
  assign n5322 = ~n5217 & n5220;
  assign n5323 = n5217 & ~n5220;
  assign n5324 = ~n5322 & ~n5323;
  assign n5325 = ~n5293 & n5296;
  assign n5326 = n5293 & ~n5296;
  assign n5327 = ~n5325 & ~n5326;
  assign n5328 = ~n5324 & ~n5327;
  assign n5329 = ~n5212 & ~n5223;
  assign n5330 = ~n5226 & ~n5329;
  assign n5331 = ~n5209 & n5330;
  assign n5332 = n5209 & ~n5330;
  assign n5333 = ~n5331 & ~n5332;
  assign n5334 = n5328 & ~n5333;
  assign n5335 = ~n5300 & ~n5302;
  assign n5336 = n5285 & n5335;
  assign n5337 = ~n5285 & ~n5335;
  assign n5338 = ~n5336 & ~n5337;
  assign n5339 = ~n5328 & n5333;
  assign n5340 = ~n5338 & ~n5339;
  assign n5341 = ~n5334 & ~n5340;
  assign n5342 = ~n5314 & ~n5320;
  assign n5343 = ~n5321 & ~n5342;
  assign n5344 = ~n5341 & n5343;
  assign n5345 = ~n5321 & ~n5344;
  assign n5346 = ~n5308 & ~n5345;
  assign n5347 = ~n5232 & ~n5307;
  assign n5348 = ~n5346 & ~n5347;
  assign n5349 = pi226  & pi227 ;
  assign n5350 = ~pi226  & pi227 ;
  assign n5351 = pi226  & ~pi227 ;
  assign n5352 = ~n5350 & ~n5351;
  assign n5353 = pi228  & ~n5352;
  assign n5354 = ~n5349 & ~n5353;
  assign n5355 = pi223  & pi224 ;
  assign n5356 = ~pi223  & pi224 ;
  assign n5357 = pi223  & ~pi224 ;
  assign n5358 = ~n5356 & ~n5357;
  assign n5359 = pi225  & ~n5358;
  assign n5360 = ~n5355 & ~n5359;
  assign n5361 = ~n5354 & n5360;
  assign n5362 = n5354 & ~n5360;
  assign n5363 = ~n5361 & ~n5362;
  assign n5364 = ~pi225  & ~n5358;
  assign n5365 = pi225  & n5358;
  assign n5366 = ~n5364 & ~n5365;
  assign n5367 = ~pi228  & ~n5352;
  assign n5368 = pi228  & n5352;
  assign n5369 = ~n5367 & ~n5368;
  assign n5370 = ~n5366 & ~n5369;
  assign n5371 = n5363 & n5370;
  assign n5372 = ~n5363 & ~n5370;
  assign n5373 = ~n5371 & ~n5372;
  assign n5374 = pi232  & pi233 ;
  assign n5375 = ~pi232  & pi233 ;
  assign n5376 = pi232  & ~pi233 ;
  assign n5377 = ~n5375 & ~n5376;
  assign n5378 = pi234  & ~n5377;
  assign n5379 = ~n5374 & ~n5378;
  assign n5380 = pi229  & pi230 ;
  assign n5381 = ~pi229  & pi230 ;
  assign n5382 = pi229  & ~pi230 ;
  assign n5383 = ~n5381 & ~n5382;
  assign n5384 = pi231  & ~n5383;
  assign n5385 = ~n5380 & ~n5384;
  assign n5386 = ~n5379 & n5385;
  assign n5387 = n5379 & ~n5385;
  assign n5388 = ~n5386 & ~n5387;
  assign n5389 = ~pi231  & ~n5383;
  assign n5390 = pi231  & n5383;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = ~pi234  & ~n5377;
  assign n5393 = pi234  & n5377;
  assign n5394 = ~n5392 & ~n5393;
  assign n5395 = ~n5391 & ~n5394;
  assign n5396 = n5388 & n5395;
  assign n5397 = ~n5388 & ~n5395;
  assign n5398 = ~n5396 & ~n5397;
  assign n5399 = ~n5388 & n5395;
  assign n5400 = ~n5379 & ~n5385;
  assign n5401 = ~n5399 & ~n5400;
  assign n5402 = ~n5398 & ~n5401;
  assign n5403 = ~n5363 & n5370;
  assign n5404 = ~n5354 & ~n5360;
  assign n5405 = ~n5403 & ~n5404;
  assign n5406 = ~n5373 & ~n5405;
  assign n5407 = ~n5391 & n5394;
  assign n5408 = n5391 & ~n5394;
  assign n5409 = ~n5407 & ~n5408;
  assign n5410 = ~n5366 & n5369;
  assign n5411 = n5366 & ~n5369;
  assign n5412 = ~n5410 & ~n5411;
  assign n5413 = ~n5409 & ~n5412;
  assign n5414 = ~n5402 & n5413;
  assign n5415 = ~n5406 & n5414;
  assign n5416 = n5398 & ~n5415;
  assign n5417 = ~n5373 & ~n5416;
  assign n5418 = ~n5398 & n5415;
  assign n5419 = ~n5417 & ~n5418;
  assign n5420 = n5401 & ~n5405;
  assign n5421 = ~n5401 & n5405;
  assign n5422 = ~n5420 & ~n5421;
  assign n5423 = ~n5419 & ~n5422;
  assign n5424 = n5419 & n5422;
  assign n5425 = ~n5423 & ~n5424;
  assign n5426 = pi235  & ~pi236 ;
  assign n5427 = ~pi235  & pi236 ;
  assign n5428 = ~n5426 & ~n5427;
  assign n5429 = ~pi237  & ~n5428;
  assign n5430 = pi237  & n5428;
  assign n5431 = ~n5429 & ~n5430;
  assign n5432 = pi238  & ~pi239 ;
  assign n5433 = ~pi238  & pi239 ;
  assign n5434 = ~n5432 & ~n5433;
  assign n5435 = ~pi240  & ~n5434;
  assign n5436 = pi240  & n5434;
  assign n5437 = ~n5435 & ~n5436;
  assign n5438 = ~n5431 & ~n5437;
  assign n5439 = pi238  & pi239 ;
  assign n5440 = pi240  & ~n5434;
  assign n5441 = ~n5439 & ~n5440;
  assign n5442 = pi235  & pi236 ;
  assign n5443 = pi237  & ~n5428;
  assign n5444 = ~n5442 & ~n5443;
  assign n5445 = n5441 & ~n5444;
  assign n5446 = ~n5441 & n5444;
  assign n5447 = ~n5445 & ~n5446;
  assign n5448 = n5438 & n5447;
  assign n5449 = ~n5438 & ~n5447;
  assign n5450 = ~n5448 & ~n5449;
  assign n5451 = pi244  & pi245 ;
  assign n5452 = pi244  & ~pi245 ;
  assign n5453 = ~pi244  & pi245 ;
  assign n5454 = ~n5452 & ~n5453;
  assign n5455 = pi246  & ~n5454;
  assign n5456 = ~n5451 & ~n5455;
  assign n5457 = pi241  & pi242 ;
  assign n5458 = pi241  & ~pi242 ;
  assign n5459 = ~pi241  & pi242 ;
  assign n5460 = ~n5458 & ~n5459;
  assign n5461 = pi243  & ~n5460;
  assign n5462 = ~n5457 & ~n5461;
  assign n5463 = ~n5456 & n5462;
  assign n5464 = n5456 & ~n5462;
  assign n5465 = ~n5463 & ~n5464;
  assign n5466 = ~pi243  & ~n5460;
  assign n5467 = pi243  & n5460;
  assign n5468 = ~n5466 & ~n5467;
  assign n5469 = ~pi246  & ~n5454;
  assign n5470 = pi246  & n5454;
  assign n5471 = ~n5469 & ~n5470;
  assign n5472 = ~n5468 & ~n5471;
  assign n5473 = n5465 & n5472;
  assign n5474 = ~n5465 & ~n5472;
  assign n5475 = ~n5473 & ~n5474;
  assign n5476 = ~n5465 & n5472;
  assign n5477 = ~n5456 & ~n5462;
  assign n5478 = ~n5476 & ~n5477;
  assign n5479 = ~n5475 & ~n5478;
  assign n5480 = n5438 & ~n5447;
  assign n5481 = ~n5441 & ~n5444;
  assign n5482 = ~n5480 & ~n5481;
  assign n5483 = ~n5450 & ~n5482;
  assign n5484 = ~n5431 & n5437;
  assign n5485 = n5431 & ~n5437;
  assign n5486 = ~n5484 & ~n5485;
  assign n5487 = ~n5468 & n5471;
  assign n5488 = n5468 & ~n5471;
  assign n5489 = ~n5487 & ~n5488;
  assign n5490 = ~n5486 & ~n5489;
  assign n5491 = ~n5479 & n5490;
  assign n5492 = ~n5483 & n5491;
  assign n5493 = n5475 & ~n5492;
  assign n5494 = ~n5450 & ~n5493;
  assign n5495 = n5475 & n5492;
  assign n5496 = n5492 & ~n5495;
  assign n5497 = ~n5494 & ~n5496;
  assign n5498 = n5478 & ~n5482;
  assign n5499 = ~n5478 & n5482;
  assign n5500 = ~n5498 & ~n5499;
  assign n5501 = ~n5497 & ~n5500;
  assign n5502 = n5497 & n5500;
  assign n5503 = ~n5501 & ~n5502;
  assign n5504 = n5425 & n5503;
  assign n5505 = ~n5486 & n5489;
  assign n5506 = n5486 & ~n5489;
  assign n5507 = ~n5505 & ~n5506;
  assign n5508 = n5409 & ~n5412;
  assign n5509 = ~n5409 & n5412;
  assign n5510 = ~n5508 & ~n5509;
  assign n5511 = ~n5507 & ~n5510;
  assign n5512 = ~n5475 & ~n5492;
  assign n5513 = ~n5495 & ~n5512;
  assign n5514 = ~n5450 & n5513;
  assign n5515 = n5450 & ~n5513;
  assign n5516 = ~n5514 & ~n5515;
  assign n5517 = n5511 & ~n5516;
  assign n5518 = ~n5416 & ~n5418;
  assign n5519 = n5373 & n5518;
  assign n5520 = ~n5373 & ~n5518;
  assign n5521 = ~n5519 & ~n5520;
  assign n5522 = ~n5511 & n5516;
  assign n5523 = ~n5521 & ~n5522;
  assign n5524 = ~n5517 & ~n5523;
  assign n5525 = ~n5425 & ~n5503;
  assign n5526 = ~n5524 & ~n5525;
  assign n5527 = ~n5504 & ~n5526;
  assign n5528 = n5478 & n5497;
  assign n5529 = ~n5482 & ~n5528;
  assign n5530 = ~n5478 & ~n5497;
  assign n5531 = ~n5529 & ~n5530;
  assign n5532 = n5401 & n5419;
  assign n5533 = ~n5405 & ~n5532;
  assign n5534 = ~n5401 & ~n5419;
  assign n5535 = ~n5533 & ~n5534;
  assign n5536 = n5531 & n5535;
  assign n5537 = ~n5527 & ~n5536;
  assign n5538 = ~n5531 & ~n5535;
  assign n5539 = ~n5537 & ~n5538;
  assign n5540 = ~n5348 & ~n5539;
  assign n5541 = ~n5324 & n5327;
  assign n5542 = n5324 & ~n5327;
  assign n5543 = ~n5541 & ~n5542;
  assign n5544 = ~n5507 & n5510;
  assign n5545 = n5507 & ~n5510;
  assign n5546 = ~n5544 & ~n5545;
  assign n5547 = ~n5543 & ~n5546;
  assign n5548 = ~n5334 & ~n5339;
  assign n5549 = ~n5338 & ~n5548;
  assign n5550 = n5338 & n5548;
  assign n5551 = ~n5549 & ~n5550;
  assign n5552 = n5547 & ~n5551;
  assign n5553 = ~n5517 & ~n5522;
  assign n5554 = n5521 & n5553;
  assign n5555 = ~n5521 & ~n5553;
  assign n5556 = ~n5554 & ~n5555;
  assign n5557 = ~n5547 & n5551;
  assign n5558 = ~n5556 & ~n5557;
  assign n5559 = ~n5552 & ~n5558;
  assign n5560 = ~n5504 & ~n5525;
  assign n5561 = ~n5524 & n5560;
  assign n5562 = n5524 & ~n5560;
  assign n5563 = ~n5561 & ~n5562;
  assign n5564 = n5341 & ~n5343;
  assign n5565 = ~n5344 & ~n5564;
  assign n5566 = ~n5563 & ~n5565;
  assign n5567 = ~n5559 & ~n5566;
  assign n5568 = n5563 & n5565;
  assign n5569 = ~n5567 & ~n5568;
  assign n5570 = ~n5308 & ~n5347;
  assign n5571 = ~n5345 & n5570;
  assign n5572 = n5345 & ~n5570;
  assign n5573 = ~n5571 & ~n5572;
  assign n5574 = n5531 & ~n5535;
  assign n5575 = ~n5531 & n5535;
  assign n5576 = ~n5504 & ~n5574;
  assign n5577 = ~n5575 & n5576;
  assign n5578 = ~n5526 & n5577;
  assign n5579 = n5537 & ~n5538;
  assign n5580 = ~n5578 & ~n5579;
  assign n5581 = ~n5573 & ~n5580;
  assign n5582 = ~n5569 & ~n5581;
  assign n5583 = n5573 & n5580;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = n5348 & n5539;
  assign n5586 = ~n5540 & ~n5585;
  assign n5587 = ~n5584 & n5586;
  assign n5588 = ~n5540 & ~n5587;
  assign n5589 = pi211  & ~pi212 ;
  assign n5590 = ~pi211  & pi212 ;
  assign n5591 = ~n5589 & ~n5590;
  assign n5592 = ~pi213  & ~n5591;
  assign n5593 = pi213  & n5591;
  assign n5594 = ~n5592 & ~n5593;
  assign n5595 = pi214  & ~pi215 ;
  assign n5596 = ~pi214  & pi215 ;
  assign n5597 = ~n5595 & ~n5596;
  assign n5598 = ~pi216  & ~n5597;
  assign n5599 = pi216  & n5597;
  assign n5600 = ~n5598 & ~n5599;
  assign n5601 = ~n5594 & ~n5600;
  assign n5602 = pi214  & pi215 ;
  assign n5603 = pi216  & ~n5597;
  assign n5604 = ~n5602 & ~n5603;
  assign n5605 = pi211  & pi212 ;
  assign n5606 = pi213  & ~n5591;
  assign n5607 = ~n5605 & ~n5606;
  assign n5608 = n5604 & ~n5607;
  assign n5609 = ~n5604 & n5607;
  assign n5610 = ~n5608 & ~n5609;
  assign n5611 = n5601 & ~n5610;
  assign n5612 = ~n5604 & ~n5607;
  assign n5613 = ~n5611 & ~n5612;
  assign n5614 = pi220  & pi221 ;
  assign n5615 = pi220  & ~pi221 ;
  assign n5616 = ~pi220  & pi221 ;
  assign n5617 = ~n5615 & ~n5616;
  assign n5618 = pi222  & ~n5617;
  assign n5619 = ~n5614 & ~n5618;
  assign n5620 = pi217  & pi218 ;
  assign n5621 = pi217  & ~pi218 ;
  assign n5622 = ~pi217  & pi218 ;
  assign n5623 = ~n5621 & ~n5622;
  assign n5624 = pi219  & ~n5623;
  assign n5625 = ~n5620 & ~n5624;
  assign n5626 = ~n5619 & n5625;
  assign n5627 = n5619 & ~n5625;
  assign n5628 = ~n5626 & ~n5627;
  assign n5629 = ~pi219  & ~n5623;
  assign n5630 = pi219  & n5623;
  assign n5631 = ~n5629 & ~n5630;
  assign n5632 = ~pi222  & ~n5617;
  assign n5633 = pi222  & n5617;
  assign n5634 = ~n5632 & ~n5633;
  assign n5635 = ~n5631 & ~n5634;
  assign n5636 = ~n5628 & n5635;
  assign n5637 = ~n5619 & ~n5625;
  assign n5638 = ~n5636 & ~n5637;
  assign n5639 = n5601 & n5610;
  assign n5640 = ~n5601 & ~n5610;
  assign n5641 = ~n5639 & ~n5640;
  assign n5642 = n5628 & n5635;
  assign n5643 = ~n5628 & ~n5635;
  assign n5644 = ~n5642 & ~n5643;
  assign n5645 = ~n5638 & ~n5644;
  assign n5646 = ~n5613 & ~n5641;
  assign n5647 = ~n5594 & n5600;
  assign n5648 = n5594 & ~n5600;
  assign n5649 = ~n5647 & ~n5648;
  assign n5650 = ~n5631 & n5634;
  assign n5651 = n5631 & ~n5634;
  assign n5652 = ~n5650 & ~n5651;
  assign n5653 = ~n5649 & ~n5652;
  assign n5654 = ~n5645 & n5653;
  assign n5655 = ~n5646 & n5654;
  assign n5656 = n5644 & ~n5655;
  assign n5657 = ~n5641 & ~n5656;
  assign n5658 = n5644 & n5655;
  assign n5659 = n5655 & ~n5658;
  assign n5660 = ~n5657 & ~n5659;
  assign n5661 = n5638 & n5660;
  assign n5662 = ~n5613 & ~n5661;
  assign n5663 = ~n5638 & ~n5660;
  assign n5664 = ~n5662 & ~n5663;
  assign n5665 = pi199  & ~pi200 ;
  assign n5666 = ~pi199  & pi200 ;
  assign n5667 = ~n5665 & ~n5666;
  assign n5668 = ~pi201  & ~n5667;
  assign n5669 = pi201  & n5667;
  assign n5670 = ~n5668 & ~n5669;
  assign n5671 = pi202  & ~pi203 ;
  assign n5672 = ~pi202  & pi203 ;
  assign n5673 = ~n5671 & ~n5672;
  assign n5674 = ~pi204  & ~n5673;
  assign n5675 = pi204  & n5673;
  assign n5676 = ~n5674 & ~n5675;
  assign n5677 = ~n5670 & ~n5676;
  assign n5678 = pi202  & pi203 ;
  assign n5679 = pi204  & ~n5673;
  assign n5680 = ~n5678 & ~n5679;
  assign n5681 = pi199  & pi200 ;
  assign n5682 = pi201  & ~n5667;
  assign n5683 = ~n5681 & ~n5682;
  assign n5684 = n5680 & ~n5683;
  assign n5685 = ~n5680 & n5683;
  assign n5686 = ~n5684 & ~n5685;
  assign n5687 = n5677 & ~n5686;
  assign n5688 = ~n5680 & ~n5683;
  assign n5689 = ~n5687 & ~n5688;
  assign n5690 = pi208  & pi209 ;
  assign n5691 = pi208  & ~pi209 ;
  assign n5692 = ~pi208  & pi209 ;
  assign n5693 = ~n5691 & ~n5692;
  assign n5694 = pi210  & ~n5693;
  assign n5695 = ~n5690 & ~n5694;
  assign n5696 = pi205  & pi206 ;
  assign n5697 = pi205  & ~pi206 ;
  assign n5698 = ~pi205  & pi206 ;
  assign n5699 = ~n5697 & ~n5698;
  assign n5700 = pi207  & ~n5699;
  assign n5701 = ~n5696 & ~n5700;
  assign n5702 = ~n5695 & n5701;
  assign n5703 = n5695 & ~n5701;
  assign n5704 = ~n5702 & ~n5703;
  assign n5705 = ~pi207  & ~n5699;
  assign n5706 = pi207  & n5699;
  assign n5707 = ~n5705 & ~n5706;
  assign n5708 = ~pi210  & ~n5693;
  assign n5709 = pi210  & n5693;
  assign n5710 = ~n5708 & ~n5709;
  assign n5711 = ~n5707 & ~n5710;
  assign n5712 = ~n5704 & n5711;
  assign n5713 = ~n5695 & ~n5701;
  assign n5714 = ~n5712 & ~n5713;
  assign n5715 = n5677 & n5686;
  assign n5716 = ~n5677 & ~n5686;
  assign n5717 = ~n5715 & ~n5716;
  assign n5718 = n5704 & n5711;
  assign n5719 = ~n5704 & ~n5711;
  assign n5720 = ~n5718 & ~n5719;
  assign n5721 = ~n5714 & ~n5720;
  assign n5722 = ~n5689 & ~n5717;
  assign n5723 = ~n5670 & n5676;
  assign n5724 = n5670 & ~n5676;
  assign n5725 = ~n5723 & ~n5724;
  assign n5726 = ~n5707 & n5710;
  assign n5727 = n5707 & ~n5710;
  assign n5728 = ~n5726 & ~n5727;
  assign n5729 = ~n5725 & ~n5728;
  assign n5730 = ~n5721 & n5729;
  assign n5731 = ~n5722 & n5730;
  assign n5732 = n5720 & ~n5731;
  assign n5733 = ~n5717 & ~n5732;
  assign n5734 = ~n5720 & n5731;
  assign n5735 = ~n5733 & ~n5734;
  assign n5736 = n5714 & n5735;
  assign n5737 = ~n5689 & ~n5736;
  assign n5738 = ~n5714 & ~n5735;
  assign n5739 = ~n5737 & ~n5738;
  assign n5740 = n5664 & n5739;
  assign n5741 = ~n5689 & n5714;
  assign n5742 = n5689 & ~n5714;
  assign n5743 = ~n5741 & ~n5742;
  assign n5744 = ~n5735 & ~n5743;
  assign n5745 = n5735 & n5743;
  assign n5746 = ~n5744 & ~n5745;
  assign n5747 = ~n5613 & n5638;
  assign n5748 = n5613 & ~n5638;
  assign n5749 = ~n5747 & ~n5748;
  assign n5750 = ~n5660 & ~n5749;
  assign n5751 = n5660 & n5749;
  assign n5752 = ~n5750 & ~n5751;
  assign n5753 = n5746 & n5752;
  assign n5754 = ~n5649 & n5652;
  assign n5755 = n5649 & ~n5652;
  assign n5756 = ~n5754 & ~n5755;
  assign n5757 = ~n5725 & n5728;
  assign n5758 = n5725 & ~n5728;
  assign n5759 = ~n5757 & ~n5758;
  assign n5760 = ~n5756 & ~n5759;
  assign n5761 = ~n5644 & ~n5655;
  assign n5762 = ~n5658 & ~n5761;
  assign n5763 = ~n5641 & n5762;
  assign n5764 = n5641 & ~n5762;
  assign n5765 = ~n5763 & ~n5764;
  assign n5766 = n5760 & ~n5765;
  assign n5767 = ~n5732 & ~n5734;
  assign n5768 = n5717 & n5767;
  assign n5769 = ~n5717 & ~n5767;
  assign n5770 = ~n5768 & ~n5769;
  assign n5771 = ~n5760 & n5765;
  assign n5772 = ~n5770 & ~n5771;
  assign n5773 = ~n5766 & ~n5772;
  assign n5774 = ~n5746 & ~n5752;
  assign n5775 = ~n5753 & ~n5774;
  assign n5776 = ~n5773 & n5775;
  assign n5777 = ~n5753 & ~n5776;
  assign n5778 = ~n5740 & ~n5777;
  assign n5779 = ~n5664 & ~n5739;
  assign n5780 = ~n5778 & ~n5779;
  assign n5781 = ~pi193  & pi194 ;
  assign n5782 = pi193  & ~pi194 ;
  assign n5783 = ~n5781 & ~n5782;
  assign n5784 = ~pi195  & ~n5783;
  assign n5785 = pi195  & n5783;
  assign n5786 = ~n5784 & ~n5785;
  assign n5787 = ~pi196  & pi197 ;
  assign n5788 = pi196  & ~pi197 ;
  assign n5789 = ~n5787 & ~n5788;
  assign n5790 = ~pi198  & ~n5789;
  assign n5791 = pi198  & n5789;
  assign n5792 = ~n5790 & ~n5791;
  assign n5793 = ~n5786 & n5792;
  assign n5794 = n5786 & ~n5792;
  assign n5795 = ~n5793 & ~n5794;
  assign n5796 = ~pi187  & pi188 ;
  assign n5797 = pi187  & ~pi188 ;
  assign n5798 = ~n5796 & ~n5797;
  assign n5799 = ~pi189  & ~n5798;
  assign n5800 = pi189  & n5798;
  assign n5801 = ~n5799 & ~n5800;
  assign n5802 = ~pi190  & pi191 ;
  assign n5803 = pi190  & ~pi191 ;
  assign n5804 = ~n5802 & ~n5803;
  assign n5805 = ~pi192  & ~n5804;
  assign n5806 = pi192  & n5804;
  assign n5807 = ~n5805 & ~n5806;
  assign n5808 = ~n5801 & n5807;
  assign n5809 = n5801 & ~n5807;
  assign n5810 = ~n5808 & ~n5809;
  assign n5811 = n5795 & ~n5810;
  assign n5812 = ~n5795 & n5810;
  assign n5813 = ~n5811 & ~n5812;
  assign n5814 = ~pi181  & pi182 ;
  assign n5815 = pi181  & ~pi182 ;
  assign n5816 = ~n5814 & ~n5815;
  assign n5817 = ~pi183  & ~n5816;
  assign n5818 = pi183  & n5816;
  assign n5819 = ~n5817 & ~n5818;
  assign n5820 = ~pi184  & pi185 ;
  assign n5821 = pi184  & ~pi185 ;
  assign n5822 = ~n5820 & ~n5821;
  assign n5823 = ~pi186  & ~n5822;
  assign n5824 = pi186  & n5822;
  assign n5825 = ~n5823 & ~n5824;
  assign n5826 = ~n5819 & n5825;
  assign n5827 = n5819 & ~n5825;
  assign n5828 = ~n5826 & ~n5827;
  assign n5829 = ~pi175  & pi176 ;
  assign n5830 = pi175  & ~pi176 ;
  assign n5831 = ~n5829 & ~n5830;
  assign n5832 = ~pi177  & ~n5831;
  assign n5833 = pi177  & n5831;
  assign n5834 = ~n5832 & ~n5833;
  assign n5835 = ~pi178  & pi179 ;
  assign n5836 = pi178  & ~pi179 ;
  assign n5837 = ~n5835 & ~n5836;
  assign n5838 = ~pi180  & ~n5837;
  assign n5839 = pi180  & n5837;
  assign n5840 = ~n5838 & ~n5839;
  assign n5841 = ~n5834 & n5840;
  assign n5842 = n5834 & ~n5840;
  assign n5843 = ~n5841 & ~n5842;
  assign n5844 = n5828 & ~n5843;
  assign n5845 = ~n5828 & n5843;
  assign n5846 = ~n5844 & ~n5845;
  assign n5847 = ~n5813 & ~n5846;
  assign n5848 = pi190  & pi191 ;
  assign n5849 = pi192  & ~n5804;
  assign n5850 = ~n5848 & ~n5849;
  assign n5851 = pi187  & pi188 ;
  assign n5852 = pi189  & ~n5798;
  assign n5853 = ~n5851 & ~n5852;
  assign n5854 = ~n5850 & n5853;
  assign n5855 = n5850 & ~n5853;
  assign n5856 = ~n5854 & ~n5855;
  assign n5857 = ~n5801 & ~n5807;
  assign n5858 = n5856 & n5857;
  assign n5859 = ~n5856 & ~n5857;
  assign n5860 = ~n5858 & ~n5859;
  assign n5861 = pi196  & pi197 ;
  assign n5862 = pi198  & ~n5789;
  assign n5863 = ~n5861 & ~n5862;
  assign n5864 = pi193  & pi194 ;
  assign n5865 = pi195  & ~n5783;
  assign n5866 = ~n5864 & ~n5865;
  assign n5867 = ~n5863 & n5866;
  assign n5868 = n5863 & ~n5866;
  assign n5869 = ~n5867 & ~n5868;
  assign n5870 = ~n5786 & ~n5792;
  assign n5871 = n5869 & n5870;
  assign n5872 = ~n5869 & ~n5870;
  assign n5873 = ~n5871 & ~n5872;
  assign n5874 = ~n5869 & n5870;
  assign n5875 = ~n5863 & ~n5866;
  assign n5876 = ~n5874 & ~n5875;
  assign n5877 = ~n5873 & ~n5876;
  assign n5878 = ~n5856 & n5857;
  assign n5879 = ~n5850 & ~n5853;
  assign n5880 = ~n5878 & ~n5879;
  assign n5881 = ~n5860 & ~n5880;
  assign n5882 = ~n5795 & ~n5810;
  assign n5883 = ~n5877 & n5882;
  assign n5884 = ~n5881 & n5883;
  assign n5885 = n5873 & ~n5884;
  assign n5886 = ~n5873 & n5884;
  assign n5887 = ~n5885 & ~n5886;
  assign n5888 = ~n5860 & ~n5887;
  assign n5889 = n5860 & n5887;
  assign n5890 = ~n5888 & ~n5889;
  assign n5891 = n5847 & ~n5890;
  assign n5892 = pi178  & pi179 ;
  assign n5893 = pi180  & ~n5837;
  assign n5894 = ~n5892 & ~n5893;
  assign n5895 = pi175  & pi176 ;
  assign n5896 = pi177  & ~n5831;
  assign n5897 = ~n5895 & ~n5896;
  assign n5898 = ~n5894 & n5897;
  assign n5899 = n5894 & ~n5897;
  assign n5900 = ~n5898 & ~n5899;
  assign n5901 = ~n5834 & ~n5840;
  assign n5902 = n5900 & n5901;
  assign n5903 = ~n5900 & ~n5901;
  assign n5904 = ~n5902 & ~n5903;
  assign n5905 = pi184  & pi185 ;
  assign n5906 = pi186  & ~n5822;
  assign n5907 = ~n5905 & ~n5906;
  assign n5908 = pi181  & pi182 ;
  assign n5909 = pi183  & ~n5816;
  assign n5910 = ~n5908 & ~n5909;
  assign n5911 = ~n5907 & n5910;
  assign n5912 = n5907 & ~n5910;
  assign n5913 = ~n5911 & ~n5912;
  assign n5914 = ~n5819 & ~n5825;
  assign n5915 = n5913 & n5914;
  assign n5916 = ~n5913 & ~n5914;
  assign n5917 = ~n5915 & ~n5916;
  assign n5918 = ~n5913 & n5914;
  assign n5919 = ~n5907 & ~n5910;
  assign n5920 = ~n5918 & ~n5919;
  assign n5921 = ~n5917 & ~n5920;
  assign n5922 = ~n5900 & n5901;
  assign n5923 = ~n5894 & ~n5897;
  assign n5924 = ~n5922 & ~n5923;
  assign n5925 = ~n5904 & ~n5924;
  assign n5926 = ~n5828 & ~n5843;
  assign n5927 = ~n5921 & n5926;
  assign n5928 = ~n5925 & n5927;
  assign n5929 = n5917 & ~n5928;
  assign n5930 = ~n5917 & n5928;
  assign n5931 = ~n5929 & ~n5930;
  assign n5932 = n5904 & n5931;
  assign n5933 = ~n5904 & ~n5931;
  assign n5934 = ~n5932 & ~n5933;
  assign n5935 = ~n5847 & n5890;
  assign n5936 = ~n5934 & ~n5935;
  assign n5937 = ~n5891 & ~n5936;
  assign n5938 = ~n5904 & ~n5929;
  assign n5939 = ~n5930 & ~n5938;
  assign n5940 = n5920 & ~n5924;
  assign n5941 = ~n5920 & n5924;
  assign n5942 = ~n5940 & ~n5941;
  assign n5943 = ~n5939 & ~n5942;
  assign n5944 = n5939 & n5942;
  assign n5945 = ~n5943 & ~n5944;
  assign n5946 = ~n5860 & ~n5885;
  assign n5947 = ~n5886 & ~n5946;
  assign n5948 = n5876 & ~n5880;
  assign n5949 = ~n5876 & n5880;
  assign n5950 = ~n5948 & ~n5949;
  assign n5951 = ~n5947 & ~n5950;
  assign n5952 = n5947 & n5950;
  assign n5953 = ~n5951 & ~n5952;
  assign n5954 = ~n5945 & ~n5953;
  assign n5955 = ~n5937 & ~n5954;
  assign n5956 = n5945 & n5953;
  assign n5957 = ~n5955 & ~n5956;
  assign n5958 = n5876 & n5947;
  assign n5959 = ~n5880 & ~n5958;
  assign n5960 = ~n5876 & ~n5947;
  assign n5961 = ~n5959 & ~n5960;
  assign n5962 = n5920 & n5939;
  assign n5963 = ~n5924 & ~n5962;
  assign n5964 = ~n5920 & ~n5939;
  assign n5965 = ~n5963 & ~n5964;
  assign n5966 = n5961 & n5965;
  assign n5967 = ~n5957 & ~n5966;
  assign n5968 = ~n5961 & ~n5965;
  assign n5969 = ~n5967 & ~n5968;
  assign n5970 = ~n5780 & ~n5969;
  assign n5971 = ~n5954 & ~n5956;
  assign n5972 = ~n5937 & n5971;
  assign n5973 = n5937 & ~n5971;
  assign n5974 = ~n5972 & ~n5973;
  assign n5975 = n5773 & ~n5775;
  assign n5976 = ~n5776 & ~n5975;
  assign n5977 = n5974 & n5976;
  assign n5978 = ~n5756 & n5759;
  assign n5979 = n5756 & ~n5759;
  assign n5980 = ~n5978 & ~n5979;
  assign n5981 = ~n5813 & n5846;
  assign n5982 = n5813 & ~n5846;
  assign n5983 = ~n5981 & ~n5982;
  assign n5984 = ~n5980 & ~n5983;
  assign n5985 = ~n5766 & ~n5771;
  assign n5986 = ~n5770 & ~n5985;
  assign n5987 = n5770 & n5985;
  assign n5988 = ~n5986 & ~n5987;
  assign n5989 = n5984 & ~n5988;
  assign n5990 = ~n5891 & ~n5935;
  assign n5991 = n5934 & n5990;
  assign n5992 = ~n5934 & ~n5990;
  assign n5993 = ~n5991 & ~n5992;
  assign n5994 = ~n5984 & n5988;
  assign n5995 = ~n5993 & ~n5994;
  assign n5996 = ~n5989 & ~n5995;
  assign n5997 = ~n5974 & ~n5976;
  assign n5998 = ~n5977 & ~n5997;
  assign n5999 = ~n5996 & n5998;
  assign n6000 = ~n5977 & ~n5999;
  assign n6001 = ~n5740 & ~n5779;
  assign n6002 = ~n5777 & n6001;
  assign n6003 = n5777 & ~n6001;
  assign n6004 = ~n6002 & ~n6003;
  assign n6005 = n5961 & ~n5965;
  assign n6006 = ~n5961 & n5965;
  assign n6007 = ~n5956 & ~n6005;
  assign n6008 = ~n6006 & n6007;
  assign n6009 = ~n5955 & n6008;
  assign n6010 = n5967 & ~n5968;
  assign n6011 = ~n6009 & ~n6010;
  assign n6012 = ~n6004 & ~n6011;
  assign n6013 = ~n6000 & ~n6012;
  assign n6014 = n6004 & n6011;
  assign n6015 = ~n6013 & ~n6014;
  assign n6016 = n5780 & n5969;
  assign n6017 = ~n5970 & ~n6016;
  assign n6018 = ~n6015 & n6017;
  assign n6019 = ~n5970 & ~n6018;
  assign n6020 = ~n5588 & ~n6019;
  assign n6021 = n5588 & n6019;
  assign n6022 = ~n6020 & ~n6021;
  assign n6023 = n6015 & ~n6017;
  assign n6024 = ~n6018 & ~n6023;
  assign n6025 = n5584 & ~n5586;
  assign n6026 = ~n5587 & ~n6025;
  assign n6027 = n6024 & n6026;
  assign n6028 = n5996 & ~n5998;
  assign n6029 = ~n5999 & ~n6028;
  assign n6030 = ~n5566 & ~n5568;
  assign n6031 = ~n5559 & n6030;
  assign n6032 = n5559 & ~n6030;
  assign n6033 = ~n6031 & ~n6032;
  assign n6034 = n6029 & n6033;
  assign n6035 = ~n5543 & n5546;
  assign n6036 = n5543 & ~n5546;
  assign n6037 = ~n6035 & ~n6036;
  assign n6038 = ~n5980 & n5983;
  assign n6039 = n5980 & ~n5983;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = ~n6037 & ~n6040;
  assign n6042 = ~n5552 & ~n5557;
  assign n6043 = ~n5556 & ~n6042;
  assign n6044 = n5556 & n6042;
  assign n6045 = ~n6043 & ~n6044;
  assign n6046 = n6041 & ~n6045;
  assign n6047 = ~n5989 & ~n5994;
  assign n6048 = n5993 & n6047;
  assign n6049 = ~n5993 & ~n6047;
  assign n6050 = ~n6048 & ~n6049;
  assign n6051 = ~n6041 & n6045;
  assign n6052 = ~n6050 & ~n6051;
  assign n6053 = ~n6046 & ~n6052;
  assign n6054 = ~n6029 & ~n6033;
  assign n6055 = ~n6034 & ~n6054;
  assign n6056 = ~n6053 & n6055;
  assign n6057 = ~n6034 & ~n6056;
  assign n6058 = ~n5581 & ~n5583;
  assign n6059 = ~n5569 & n6058;
  assign n6060 = n5569 & ~n6058;
  assign n6061 = ~n6059 & ~n6060;
  assign n6062 = ~n6012 & ~n6014;
  assign n6063 = ~n6000 & n6062;
  assign n6064 = n6000 & ~n6062;
  assign n6065 = ~n6063 & ~n6064;
  assign n6066 = ~n6061 & ~n6065;
  assign n6067 = ~n6057 & ~n6066;
  assign n6068 = n6061 & n6065;
  assign n6069 = ~n6067 & ~n6068;
  assign n6070 = ~n6024 & ~n6026;
  assign n6071 = ~n6027 & ~n6070;
  assign n6072 = ~n6069 & n6071;
  assign n6073 = ~n6027 & ~n6072;
  assign n6074 = n6022 & ~n6073;
  assign n6075 = ~n6020 & ~n6074;
  assign n6076 = pi166  & pi167 ;
  assign n6077 = ~pi166  & pi167 ;
  assign n6078 = pi166  & ~pi167 ;
  assign n6079 = ~n6077 & ~n6078;
  assign n6080 = pi168  & ~n6079;
  assign n6081 = ~n6076 & ~n6080;
  assign n6082 = pi163  & pi164 ;
  assign n6083 = ~pi163  & pi164 ;
  assign n6084 = pi163  & ~pi164 ;
  assign n6085 = ~n6083 & ~n6084;
  assign n6086 = pi165  & ~n6085;
  assign n6087 = ~n6082 & ~n6086;
  assign n6088 = ~n6081 & n6087;
  assign n6089 = n6081 & ~n6087;
  assign n6090 = ~n6088 & ~n6089;
  assign n6091 = ~pi165  & ~n6085;
  assign n6092 = pi165  & n6085;
  assign n6093 = ~n6091 & ~n6092;
  assign n6094 = ~pi168  & ~n6079;
  assign n6095 = pi168  & n6079;
  assign n6096 = ~n6094 & ~n6095;
  assign n6097 = ~n6093 & ~n6096;
  assign n6098 = ~n6090 & n6097;
  assign n6099 = ~n6081 & ~n6087;
  assign n6100 = ~n6098 & ~n6099;
  assign n6101 = pi172  & pi173 ;
  assign n6102 = ~pi172  & pi173 ;
  assign n6103 = pi172  & ~pi173 ;
  assign n6104 = ~n6102 & ~n6103;
  assign n6105 = pi174  & ~n6104;
  assign n6106 = ~n6101 & ~n6105;
  assign n6107 = pi169  & pi170 ;
  assign n6108 = ~pi169  & pi170 ;
  assign n6109 = pi169  & ~pi170 ;
  assign n6110 = ~n6108 & ~n6109;
  assign n6111 = pi171  & ~n6110;
  assign n6112 = ~n6107 & ~n6111;
  assign n6113 = ~n6106 & n6112;
  assign n6114 = n6106 & ~n6112;
  assign n6115 = ~n6113 & ~n6114;
  assign n6116 = ~pi171  & ~n6110;
  assign n6117 = pi171  & n6110;
  assign n6118 = ~n6116 & ~n6117;
  assign n6119 = ~pi174  & ~n6104;
  assign n6120 = pi174  & n6104;
  assign n6121 = ~n6119 & ~n6120;
  assign n6122 = ~n6118 & ~n6121;
  assign n6123 = ~n6115 & n6122;
  assign n6124 = ~n6106 & ~n6112;
  assign n6125 = ~n6123 & ~n6124;
  assign n6126 = n6115 & n6122;
  assign n6127 = ~n6115 & ~n6122;
  assign n6128 = ~n6126 & ~n6127;
  assign n6129 = ~n6125 & ~n6128;
  assign n6130 = n6090 & n6097;
  assign n6131 = ~n6090 & ~n6097;
  assign n6132 = ~n6130 & ~n6131;
  assign n6133 = ~n6100 & ~n6132;
  assign n6134 = ~n6118 & n6121;
  assign n6135 = n6118 & ~n6121;
  assign n6136 = ~n6134 & ~n6135;
  assign n6137 = ~n6093 & n6096;
  assign n6138 = n6093 & ~n6096;
  assign n6139 = ~n6137 & ~n6138;
  assign n6140 = ~n6136 & ~n6139;
  assign n6141 = ~n6129 & n6140;
  assign n6142 = ~n6133 & n6141;
  assign n6143 = ~n6128 & n6142;
  assign n6144 = n6128 & ~n6142;
  assign n6145 = ~n6132 & ~n6144;
  assign n6146 = ~n6143 & ~n6145;
  assign n6147 = n6125 & n6146;
  assign n6148 = ~n6100 & ~n6147;
  assign n6149 = ~n6125 & ~n6146;
  assign n6150 = ~n6148 & ~n6149;
  assign n6151 = pi154  & pi155 ;
  assign n6152 = ~pi154  & pi155 ;
  assign n6153 = pi154  & ~pi155 ;
  assign n6154 = ~n6152 & ~n6153;
  assign n6155 = pi156  & ~n6154;
  assign n6156 = ~n6151 & ~n6155;
  assign n6157 = pi151  & pi152 ;
  assign n6158 = ~pi151  & pi152 ;
  assign n6159 = pi151  & ~pi152 ;
  assign n6160 = ~n6158 & ~n6159;
  assign n6161 = pi153  & ~n6160;
  assign n6162 = ~n6157 & ~n6161;
  assign n6163 = ~n6156 & n6162;
  assign n6164 = n6156 & ~n6162;
  assign n6165 = ~n6163 & ~n6164;
  assign n6166 = ~pi153  & ~n6160;
  assign n6167 = pi153  & n6160;
  assign n6168 = ~n6166 & ~n6167;
  assign n6169 = ~pi156  & ~n6154;
  assign n6170 = pi156  & n6154;
  assign n6171 = ~n6169 & ~n6170;
  assign n6172 = ~n6168 & ~n6171;
  assign n6173 = ~n6165 & n6172;
  assign n6174 = ~n6156 & ~n6162;
  assign n6175 = ~n6173 & ~n6174;
  assign n6176 = pi160  & pi161 ;
  assign n6177 = ~pi160  & pi161 ;
  assign n6178 = pi160  & ~pi161 ;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = pi162  & ~n6179;
  assign n6181 = ~n6176 & ~n6180;
  assign n6182 = pi157  & pi158 ;
  assign n6183 = ~pi157  & pi158 ;
  assign n6184 = pi157  & ~pi158 ;
  assign n6185 = ~n6183 & ~n6184;
  assign n6186 = pi159  & ~n6185;
  assign n6187 = ~n6182 & ~n6186;
  assign n6188 = ~n6181 & n6187;
  assign n6189 = n6181 & ~n6187;
  assign n6190 = ~n6188 & ~n6189;
  assign n6191 = ~pi159  & ~n6185;
  assign n6192 = pi159  & n6185;
  assign n6193 = ~n6191 & ~n6192;
  assign n6194 = ~pi162  & ~n6179;
  assign n6195 = pi162  & n6179;
  assign n6196 = ~n6194 & ~n6195;
  assign n6197 = ~n6193 & ~n6196;
  assign n6198 = ~n6190 & n6197;
  assign n6199 = ~n6181 & ~n6187;
  assign n6200 = ~n6198 & ~n6199;
  assign n6201 = n6190 & n6197;
  assign n6202 = ~n6190 & ~n6197;
  assign n6203 = ~n6201 & ~n6202;
  assign n6204 = ~n6200 & ~n6203;
  assign n6205 = n6165 & n6172;
  assign n6206 = ~n6165 & ~n6172;
  assign n6207 = ~n6205 & ~n6206;
  assign n6208 = ~n6175 & ~n6207;
  assign n6209 = ~n6193 & n6196;
  assign n6210 = n6193 & ~n6196;
  assign n6211 = ~n6209 & ~n6210;
  assign n6212 = ~n6168 & n6171;
  assign n6213 = n6168 & ~n6171;
  assign n6214 = ~n6212 & ~n6213;
  assign n6215 = ~n6211 & ~n6214;
  assign n6216 = ~n6204 & n6215;
  assign n6217 = ~n6208 & n6216;
  assign n6218 = ~n6203 & n6217;
  assign n6219 = n6203 & ~n6217;
  assign n6220 = ~n6207 & ~n6219;
  assign n6221 = ~n6218 & ~n6220;
  assign n6222 = n6200 & n6221;
  assign n6223 = ~n6175 & ~n6222;
  assign n6224 = ~n6200 & ~n6221;
  assign n6225 = ~n6223 & ~n6224;
  assign n6226 = n6150 & n6225;
  assign n6227 = ~n6175 & n6200;
  assign n6228 = n6175 & ~n6200;
  assign n6229 = ~n6227 & ~n6228;
  assign n6230 = ~n6221 & ~n6229;
  assign n6231 = n6221 & n6229;
  assign n6232 = ~n6230 & ~n6231;
  assign n6233 = ~n6100 & n6125;
  assign n6234 = n6100 & ~n6125;
  assign n6235 = ~n6233 & ~n6234;
  assign n6236 = ~n6146 & ~n6235;
  assign n6237 = n6146 & n6235;
  assign n6238 = ~n6236 & ~n6237;
  assign n6239 = n6232 & n6238;
  assign n6240 = n6136 & ~n6139;
  assign n6241 = ~n6136 & n6139;
  assign n6242 = ~n6240 & ~n6241;
  assign n6243 = n6211 & ~n6214;
  assign n6244 = ~n6211 & n6214;
  assign n6245 = ~n6243 & ~n6244;
  assign n6246 = ~n6242 & ~n6245;
  assign n6247 = ~n6143 & ~n6144;
  assign n6248 = ~n6132 & ~n6247;
  assign n6249 = n6132 & n6247;
  assign n6250 = ~n6248 & ~n6249;
  assign n6251 = n6246 & ~n6250;
  assign n6252 = ~n6218 & ~n6219;
  assign n6253 = n6207 & n6252;
  assign n6254 = ~n6207 & ~n6252;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~n6246 & n6250;
  assign n6257 = ~n6255 & ~n6256;
  assign n6258 = ~n6251 & ~n6257;
  assign n6259 = ~n6232 & ~n6238;
  assign n6260 = ~n6239 & ~n6259;
  assign n6261 = ~n6258 & n6260;
  assign n6262 = ~n6239 & ~n6261;
  assign n6263 = ~n6226 & ~n6262;
  assign n6264 = ~n6150 & ~n6225;
  assign n6265 = ~n6263 & ~n6264;
  assign n6266 = ~pi145  & pi146 ;
  assign n6267 = pi145  & ~pi146 ;
  assign n6268 = ~n6266 & ~n6267;
  assign n6269 = ~pi147  & ~n6268;
  assign n6270 = pi147  & n6268;
  assign n6271 = ~n6269 & ~n6270;
  assign n6272 = ~pi148  & pi149 ;
  assign n6273 = pi148  & ~pi149 ;
  assign n6274 = ~n6272 & ~n6273;
  assign n6275 = ~pi150  & ~n6274;
  assign n6276 = pi150  & n6274;
  assign n6277 = ~n6275 & ~n6276;
  assign n6278 = ~n6271 & n6277;
  assign n6279 = n6271 & ~n6277;
  assign n6280 = ~n6278 & ~n6279;
  assign n6281 = ~pi139  & pi140 ;
  assign n6282 = pi139  & ~pi140 ;
  assign n6283 = ~n6281 & ~n6282;
  assign n6284 = ~pi141  & ~n6283;
  assign n6285 = pi141  & n6283;
  assign n6286 = ~n6284 & ~n6285;
  assign n6287 = ~pi142  & pi143 ;
  assign n6288 = pi142  & ~pi143 ;
  assign n6289 = ~n6287 & ~n6288;
  assign n6290 = ~pi144  & ~n6289;
  assign n6291 = pi144  & n6289;
  assign n6292 = ~n6290 & ~n6291;
  assign n6293 = ~n6286 & n6292;
  assign n6294 = n6286 & ~n6292;
  assign n6295 = ~n6293 & ~n6294;
  assign n6296 = n6280 & ~n6295;
  assign n6297 = ~n6280 & n6295;
  assign n6298 = ~n6296 & ~n6297;
  assign n6299 = ~pi133  & pi134 ;
  assign n6300 = pi133  & ~pi134 ;
  assign n6301 = ~n6299 & ~n6300;
  assign n6302 = ~pi135  & ~n6301;
  assign n6303 = pi135  & n6301;
  assign n6304 = ~n6302 & ~n6303;
  assign n6305 = ~pi136  & pi137 ;
  assign n6306 = pi136  & ~pi137 ;
  assign n6307 = ~n6305 & ~n6306;
  assign n6308 = ~pi138  & ~n6307;
  assign n6309 = pi138  & n6307;
  assign n6310 = ~n6308 & ~n6309;
  assign n6311 = ~n6304 & n6310;
  assign n6312 = n6304 & ~n6310;
  assign n6313 = ~n6311 & ~n6312;
  assign n6314 = ~pi127  & pi128 ;
  assign n6315 = pi127  & ~pi128 ;
  assign n6316 = ~n6314 & ~n6315;
  assign n6317 = ~pi129  & ~n6316;
  assign n6318 = pi129  & n6316;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = ~pi130  & pi131 ;
  assign n6321 = pi130  & ~pi131 ;
  assign n6322 = ~n6320 & ~n6321;
  assign n6323 = ~pi132  & ~n6322;
  assign n6324 = pi132  & n6322;
  assign n6325 = ~n6323 & ~n6324;
  assign n6326 = ~n6319 & n6325;
  assign n6327 = n6319 & ~n6325;
  assign n6328 = ~n6326 & ~n6327;
  assign n6329 = n6313 & ~n6328;
  assign n6330 = ~n6313 & n6328;
  assign n6331 = ~n6329 & ~n6330;
  assign n6332 = ~n6298 & ~n6331;
  assign n6333 = pi142  & pi143 ;
  assign n6334 = pi144  & ~n6289;
  assign n6335 = ~n6333 & ~n6334;
  assign n6336 = pi139  & pi140 ;
  assign n6337 = pi141  & ~n6283;
  assign n6338 = ~n6336 & ~n6337;
  assign n6339 = ~n6335 & n6338;
  assign n6340 = n6335 & ~n6338;
  assign n6341 = ~n6339 & ~n6340;
  assign n6342 = ~n6286 & ~n6292;
  assign n6343 = n6341 & n6342;
  assign n6344 = ~n6341 & ~n6342;
  assign n6345 = ~n6343 & ~n6344;
  assign n6346 = pi148  & pi149 ;
  assign n6347 = pi150  & ~n6274;
  assign n6348 = ~n6346 & ~n6347;
  assign n6349 = pi145  & pi146 ;
  assign n6350 = pi147  & ~n6268;
  assign n6351 = ~n6349 & ~n6350;
  assign n6352 = ~n6348 & n6351;
  assign n6353 = n6348 & ~n6351;
  assign n6354 = ~n6352 & ~n6353;
  assign n6355 = ~n6271 & ~n6277;
  assign n6356 = n6354 & n6355;
  assign n6357 = ~n6354 & ~n6355;
  assign n6358 = ~n6356 & ~n6357;
  assign n6359 = ~n6354 & n6355;
  assign n6360 = ~n6348 & ~n6351;
  assign n6361 = ~n6359 & ~n6360;
  assign n6362 = ~n6358 & ~n6361;
  assign n6363 = ~n6341 & n6342;
  assign n6364 = ~n6335 & ~n6338;
  assign n6365 = ~n6363 & ~n6364;
  assign n6366 = ~n6345 & ~n6365;
  assign n6367 = ~n6280 & ~n6295;
  assign n6368 = ~n6362 & n6367;
  assign n6369 = ~n6366 & n6368;
  assign n6370 = n6358 & ~n6369;
  assign n6371 = ~n6358 & n6369;
  assign n6372 = ~n6370 & ~n6371;
  assign n6373 = ~n6345 & ~n6372;
  assign n6374 = n6345 & n6372;
  assign n6375 = ~n6373 & ~n6374;
  assign n6376 = n6332 & ~n6375;
  assign n6377 = pi130  & pi131 ;
  assign n6378 = pi132  & ~n6322;
  assign n6379 = ~n6377 & ~n6378;
  assign n6380 = pi127  & pi128 ;
  assign n6381 = pi129  & ~n6316;
  assign n6382 = ~n6380 & ~n6381;
  assign n6383 = ~n6379 & n6382;
  assign n6384 = n6379 & ~n6382;
  assign n6385 = ~n6383 & ~n6384;
  assign n6386 = ~n6319 & ~n6325;
  assign n6387 = n6385 & n6386;
  assign n6388 = ~n6385 & ~n6386;
  assign n6389 = ~n6387 & ~n6388;
  assign n6390 = pi136  & pi137 ;
  assign n6391 = pi138  & ~n6307;
  assign n6392 = ~n6390 & ~n6391;
  assign n6393 = pi133  & pi134 ;
  assign n6394 = pi135  & ~n6301;
  assign n6395 = ~n6393 & ~n6394;
  assign n6396 = ~n6392 & n6395;
  assign n6397 = n6392 & ~n6395;
  assign n6398 = ~n6396 & ~n6397;
  assign n6399 = ~n6304 & ~n6310;
  assign n6400 = n6398 & n6399;
  assign n6401 = ~n6398 & ~n6399;
  assign n6402 = ~n6400 & ~n6401;
  assign n6403 = ~n6398 & n6399;
  assign n6404 = ~n6392 & ~n6395;
  assign n6405 = ~n6403 & ~n6404;
  assign n6406 = ~n6402 & ~n6405;
  assign n6407 = ~n6385 & n6386;
  assign n6408 = ~n6379 & ~n6382;
  assign n6409 = ~n6407 & ~n6408;
  assign n6410 = ~n6389 & ~n6409;
  assign n6411 = ~n6313 & ~n6328;
  assign n6412 = ~n6406 & n6411;
  assign n6413 = ~n6410 & n6412;
  assign n6414 = n6402 & ~n6413;
  assign n6415 = ~n6402 & n6413;
  assign n6416 = ~n6414 & ~n6415;
  assign n6417 = n6389 & n6416;
  assign n6418 = ~n6389 & ~n6416;
  assign n6419 = ~n6417 & ~n6418;
  assign n6420 = ~n6332 & n6375;
  assign n6421 = ~n6419 & ~n6420;
  assign n6422 = ~n6376 & ~n6421;
  assign n6423 = ~n6389 & ~n6414;
  assign n6424 = ~n6415 & ~n6423;
  assign n6425 = n6405 & ~n6409;
  assign n6426 = ~n6405 & n6409;
  assign n6427 = ~n6425 & ~n6426;
  assign n6428 = ~n6424 & ~n6427;
  assign n6429 = n6424 & n6427;
  assign n6430 = ~n6428 & ~n6429;
  assign n6431 = ~n6345 & ~n6370;
  assign n6432 = ~n6371 & ~n6431;
  assign n6433 = n6361 & ~n6365;
  assign n6434 = ~n6361 & n6365;
  assign n6435 = ~n6433 & ~n6434;
  assign n6436 = ~n6432 & ~n6435;
  assign n6437 = n6432 & n6435;
  assign n6438 = ~n6436 & ~n6437;
  assign n6439 = ~n6430 & ~n6438;
  assign n6440 = ~n6422 & ~n6439;
  assign n6441 = n6430 & n6438;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = n6361 & n6432;
  assign n6444 = ~n6365 & ~n6443;
  assign n6445 = ~n6361 & ~n6432;
  assign n6446 = ~n6444 & ~n6445;
  assign n6447 = n6405 & n6424;
  assign n6448 = ~n6409 & ~n6447;
  assign n6449 = ~n6405 & ~n6424;
  assign n6450 = ~n6448 & ~n6449;
  assign n6451 = n6446 & n6450;
  assign n6452 = ~n6442 & ~n6451;
  assign n6453 = ~n6446 & ~n6450;
  assign n6454 = ~n6452 & ~n6453;
  assign n6455 = ~n6265 & ~n6454;
  assign n6456 = ~n6439 & ~n6441;
  assign n6457 = ~n6422 & n6456;
  assign n6458 = n6422 & ~n6456;
  assign n6459 = ~n6457 & ~n6458;
  assign n6460 = n6258 & ~n6260;
  assign n6461 = ~n6261 & ~n6460;
  assign n6462 = n6459 & n6461;
  assign n6463 = ~n6242 & n6245;
  assign n6464 = n6242 & ~n6245;
  assign n6465 = ~n6463 & ~n6464;
  assign n6466 = ~n6298 & n6331;
  assign n6467 = n6298 & ~n6331;
  assign n6468 = ~n6466 & ~n6467;
  assign n6469 = ~n6465 & ~n6468;
  assign n6470 = ~n6251 & ~n6256;
  assign n6471 = ~n6255 & ~n6470;
  assign n6472 = n6255 & n6470;
  assign n6473 = ~n6471 & ~n6472;
  assign n6474 = n6469 & ~n6473;
  assign n6475 = ~n6376 & ~n6420;
  assign n6476 = n6419 & n6475;
  assign n6477 = ~n6419 & ~n6475;
  assign n6478 = ~n6476 & ~n6477;
  assign n6479 = ~n6469 & n6473;
  assign n6480 = ~n6478 & ~n6479;
  assign n6481 = ~n6474 & ~n6480;
  assign n6482 = ~n6459 & ~n6461;
  assign n6483 = ~n6462 & ~n6482;
  assign n6484 = ~n6481 & n6483;
  assign n6485 = ~n6462 & ~n6484;
  assign n6486 = ~n6226 & ~n6264;
  assign n6487 = ~n6262 & n6486;
  assign n6488 = n6262 & ~n6486;
  assign n6489 = ~n6487 & ~n6488;
  assign n6490 = n6446 & ~n6450;
  assign n6491 = ~n6446 & n6450;
  assign n6492 = ~n6441 & ~n6490;
  assign n6493 = ~n6491 & n6492;
  assign n6494 = ~n6440 & n6493;
  assign n6495 = n6452 & ~n6453;
  assign n6496 = ~n6494 & ~n6495;
  assign n6497 = ~n6489 & ~n6496;
  assign n6498 = ~n6485 & ~n6497;
  assign n6499 = n6489 & n6496;
  assign n6500 = ~n6498 & ~n6499;
  assign n6501 = n6265 & n6454;
  assign n6502 = ~n6455 & ~n6501;
  assign n6503 = ~n6500 & n6502;
  assign n6504 = ~n6455 & ~n6503;
  assign n6505 = pi118  & pi119 ;
  assign n6506 = ~pi118  & pi119 ;
  assign n6507 = pi118  & ~pi119 ;
  assign n6508 = ~n6506 & ~n6507;
  assign n6509 = pi120  & ~n6508;
  assign n6510 = ~n6505 & ~n6509;
  assign n6511 = pi115  & pi116 ;
  assign n6512 = ~pi115  & pi116 ;
  assign n6513 = pi115  & ~pi116 ;
  assign n6514 = ~n6512 & ~n6513;
  assign n6515 = pi117  & ~n6514;
  assign n6516 = ~n6511 & ~n6515;
  assign n6517 = ~n6510 & n6516;
  assign n6518 = n6510 & ~n6516;
  assign n6519 = ~n6517 & ~n6518;
  assign n6520 = ~pi117  & ~n6514;
  assign n6521 = pi117  & n6514;
  assign n6522 = ~n6520 & ~n6521;
  assign n6523 = ~pi120  & ~n6508;
  assign n6524 = pi120  & n6508;
  assign n6525 = ~n6523 & ~n6524;
  assign n6526 = ~n6522 & ~n6525;
  assign n6527 = ~n6519 & n6526;
  assign n6528 = ~n6510 & ~n6516;
  assign n6529 = ~n6527 & ~n6528;
  assign n6530 = pi124  & pi125 ;
  assign n6531 = ~pi124  & pi125 ;
  assign n6532 = pi124  & ~pi125 ;
  assign n6533 = ~n6531 & ~n6532;
  assign n6534 = pi126  & ~n6533;
  assign n6535 = ~n6530 & ~n6534;
  assign n6536 = pi121  & pi122 ;
  assign n6537 = ~pi121  & pi122 ;
  assign n6538 = pi121  & ~pi122 ;
  assign n6539 = ~n6537 & ~n6538;
  assign n6540 = pi123  & ~n6539;
  assign n6541 = ~n6536 & ~n6540;
  assign n6542 = ~n6535 & n6541;
  assign n6543 = n6535 & ~n6541;
  assign n6544 = ~n6542 & ~n6543;
  assign n6545 = ~pi123  & ~n6539;
  assign n6546 = pi123  & n6539;
  assign n6547 = ~n6545 & ~n6546;
  assign n6548 = ~pi126  & ~n6533;
  assign n6549 = pi126  & n6533;
  assign n6550 = ~n6548 & ~n6549;
  assign n6551 = ~n6547 & ~n6550;
  assign n6552 = ~n6544 & n6551;
  assign n6553 = ~n6535 & ~n6541;
  assign n6554 = ~n6552 & ~n6553;
  assign n6555 = n6544 & n6551;
  assign n6556 = ~n6544 & ~n6551;
  assign n6557 = ~n6555 & ~n6556;
  assign n6558 = ~n6554 & ~n6557;
  assign n6559 = n6519 & n6526;
  assign n6560 = ~n6519 & ~n6526;
  assign n6561 = ~n6559 & ~n6560;
  assign n6562 = ~n6529 & ~n6561;
  assign n6563 = ~n6547 & n6550;
  assign n6564 = n6547 & ~n6550;
  assign n6565 = ~n6563 & ~n6564;
  assign n6566 = ~n6522 & n6525;
  assign n6567 = n6522 & ~n6525;
  assign n6568 = ~n6566 & ~n6567;
  assign n6569 = ~n6565 & ~n6568;
  assign n6570 = ~n6558 & n6569;
  assign n6571 = ~n6562 & n6570;
  assign n6572 = ~n6557 & n6571;
  assign n6573 = n6557 & ~n6571;
  assign n6574 = ~n6561 & ~n6573;
  assign n6575 = ~n6572 & ~n6574;
  assign n6576 = n6554 & n6575;
  assign n6577 = ~n6529 & ~n6576;
  assign n6578 = ~n6554 & ~n6575;
  assign n6579 = ~n6577 & ~n6578;
  assign n6580 = pi106  & pi107 ;
  assign n6581 = ~pi106  & pi107 ;
  assign n6582 = pi106  & ~pi107 ;
  assign n6583 = ~n6581 & ~n6582;
  assign n6584 = pi108  & ~n6583;
  assign n6585 = ~n6580 & ~n6584;
  assign n6586 = pi103  & pi104 ;
  assign n6587 = ~pi103  & pi104 ;
  assign n6588 = pi103  & ~pi104 ;
  assign n6589 = ~n6587 & ~n6588;
  assign n6590 = pi105  & ~n6589;
  assign n6591 = ~n6586 & ~n6590;
  assign n6592 = ~n6585 & n6591;
  assign n6593 = n6585 & ~n6591;
  assign n6594 = ~n6592 & ~n6593;
  assign n6595 = ~pi105  & ~n6589;
  assign n6596 = pi105  & n6589;
  assign n6597 = ~n6595 & ~n6596;
  assign n6598 = ~pi108  & ~n6583;
  assign n6599 = pi108  & n6583;
  assign n6600 = ~n6598 & ~n6599;
  assign n6601 = ~n6597 & ~n6600;
  assign n6602 = ~n6594 & n6601;
  assign n6603 = ~n6585 & ~n6591;
  assign n6604 = ~n6602 & ~n6603;
  assign n6605 = pi112  & pi113 ;
  assign n6606 = ~pi112  & pi113 ;
  assign n6607 = pi112  & ~pi113 ;
  assign n6608 = ~n6606 & ~n6607;
  assign n6609 = pi114  & ~n6608;
  assign n6610 = ~n6605 & ~n6609;
  assign n6611 = pi109  & pi110 ;
  assign n6612 = ~pi109  & pi110 ;
  assign n6613 = pi109  & ~pi110 ;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = pi111  & ~n6614;
  assign n6616 = ~n6611 & ~n6615;
  assign n6617 = ~n6610 & n6616;
  assign n6618 = n6610 & ~n6616;
  assign n6619 = ~n6617 & ~n6618;
  assign n6620 = ~pi111  & ~n6614;
  assign n6621 = pi111  & n6614;
  assign n6622 = ~n6620 & ~n6621;
  assign n6623 = ~pi114  & ~n6608;
  assign n6624 = pi114  & n6608;
  assign n6625 = ~n6623 & ~n6624;
  assign n6626 = ~n6622 & ~n6625;
  assign n6627 = ~n6619 & n6626;
  assign n6628 = ~n6610 & ~n6616;
  assign n6629 = ~n6627 & ~n6628;
  assign n6630 = n6619 & n6626;
  assign n6631 = ~n6619 & ~n6626;
  assign n6632 = ~n6630 & ~n6631;
  assign n6633 = ~n6629 & ~n6632;
  assign n6634 = n6594 & n6601;
  assign n6635 = ~n6594 & ~n6601;
  assign n6636 = ~n6634 & ~n6635;
  assign n6637 = ~n6604 & ~n6636;
  assign n6638 = ~n6622 & n6625;
  assign n6639 = n6622 & ~n6625;
  assign n6640 = ~n6638 & ~n6639;
  assign n6641 = ~n6597 & n6600;
  assign n6642 = n6597 & ~n6600;
  assign n6643 = ~n6641 & ~n6642;
  assign n6644 = ~n6640 & ~n6643;
  assign n6645 = ~n6633 & n6644;
  assign n6646 = ~n6637 & n6645;
  assign n6647 = ~n6632 & n6646;
  assign n6648 = n6632 & ~n6646;
  assign n6649 = ~n6636 & ~n6648;
  assign n6650 = ~n6647 & ~n6649;
  assign n6651 = n6629 & n6650;
  assign n6652 = ~n6604 & ~n6651;
  assign n6653 = ~n6629 & ~n6650;
  assign n6654 = ~n6652 & ~n6653;
  assign n6655 = n6579 & n6654;
  assign n6656 = ~n6604 & n6629;
  assign n6657 = n6604 & ~n6629;
  assign n6658 = ~n6656 & ~n6657;
  assign n6659 = ~n6650 & ~n6658;
  assign n6660 = n6650 & n6658;
  assign n6661 = ~n6659 & ~n6660;
  assign n6662 = ~n6529 & n6554;
  assign n6663 = n6529 & ~n6554;
  assign n6664 = ~n6662 & ~n6663;
  assign n6665 = ~n6575 & ~n6664;
  assign n6666 = n6575 & n6664;
  assign n6667 = ~n6665 & ~n6666;
  assign n6668 = n6661 & n6667;
  assign n6669 = n6565 & ~n6568;
  assign n6670 = ~n6565 & n6568;
  assign n6671 = ~n6669 & ~n6670;
  assign n6672 = n6640 & ~n6643;
  assign n6673 = ~n6640 & n6643;
  assign n6674 = ~n6672 & ~n6673;
  assign n6675 = ~n6671 & ~n6674;
  assign n6676 = ~n6572 & ~n6573;
  assign n6677 = ~n6561 & ~n6676;
  assign n6678 = n6561 & n6676;
  assign n6679 = ~n6677 & ~n6678;
  assign n6680 = n6675 & ~n6679;
  assign n6681 = ~n6647 & ~n6648;
  assign n6682 = n6636 & n6681;
  assign n6683 = ~n6636 & ~n6681;
  assign n6684 = ~n6682 & ~n6683;
  assign n6685 = ~n6675 & n6679;
  assign n6686 = ~n6684 & ~n6685;
  assign n6687 = ~n6680 & ~n6686;
  assign n6688 = ~n6661 & ~n6667;
  assign n6689 = ~n6668 & ~n6688;
  assign n6690 = ~n6687 & n6689;
  assign n6691 = ~n6668 & ~n6690;
  assign n6692 = ~n6655 & ~n6691;
  assign n6693 = ~n6579 & ~n6654;
  assign n6694 = ~n6692 & ~n6693;
  assign n6695 = ~pi97  & pi98 ;
  assign n6696 = pi97  & ~pi98 ;
  assign n6697 = ~n6695 & ~n6696;
  assign n6698 = ~pi99  & ~n6697;
  assign n6699 = pi99  & n6697;
  assign n6700 = ~n6698 & ~n6699;
  assign n6701 = ~pi100  & pi101 ;
  assign n6702 = pi100  & ~pi101 ;
  assign n6703 = ~n6701 & ~n6702;
  assign n6704 = ~pi102  & ~n6703;
  assign n6705 = pi102  & n6703;
  assign n6706 = ~n6704 & ~n6705;
  assign n6707 = ~n6700 & n6706;
  assign n6708 = n6700 & ~n6706;
  assign n6709 = ~n6707 & ~n6708;
  assign n6710 = ~pi91  & pi92 ;
  assign n6711 = pi91  & ~pi92 ;
  assign n6712 = ~n6710 & ~n6711;
  assign n6713 = ~pi93  & ~n6712;
  assign n6714 = pi93  & n6712;
  assign n6715 = ~n6713 & ~n6714;
  assign n6716 = ~pi94  & pi95 ;
  assign n6717 = pi94  & ~pi95 ;
  assign n6718 = ~n6716 & ~n6717;
  assign n6719 = ~pi96  & ~n6718;
  assign n6720 = pi96  & n6718;
  assign n6721 = ~n6719 & ~n6720;
  assign n6722 = ~n6715 & n6721;
  assign n6723 = n6715 & ~n6721;
  assign n6724 = ~n6722 & ~n6723;
  assign n6725 = n6709 & ~n6724;
  assign n6726 = ~n6709 & n6724;
  assign n6727 = ~n6725 & ~n6726;
  assign n6728 = ~pi85  & pi86 ;
  assign n6729 = pi85  & ~pi86 ;
  assign n6730 = ~n6728 & ~n6729;
  assign n6731 = ~pi87  & ~n6730;
  assign n6732 = pi87  & n6730;
  assign n6733 = ~n6731 & ~n6732;
  assign n6734 = ~pi88  & pi89 ;
  assign n6735 = pi88  & ~pi89 ;
  assign n6736 = ~n6734 & ~n6735;
  assign n6737 = ~pi90  & ~n6736;
  assign n6738 = pi90  & n6736;
  assign n6739 = ~n6737 & ~n6738;
  assign n6740 = ~n6733 & n6739;
  assign n6741 = n6733 & ~n6739;
  assign n6742 = ~n6740 & ~n6741;
  assign n6743 = ~pi79  & pi80 ;
  assign n6744 = pi79  & ~pi80 ;
  assign n6745 = ~n6743 & ~n6744;
  assign n6746 = ~pi81  & ~n6745;
  assign n6747 = pi81  & n6745;
  assign n6748 = ~n6746 & ~n6747;
  assign n6749 = ~pi82  & pi83 ;
  assign n6750 = pi82  & ~pi83 ;
  assign n6751 = ~n6749 & ~n6750;
  assign n6752 = ~pi84  & ~n6751;
  assign n6753 = pi84  & n6751;
  assign n6754 = ~n6752 & ~n6753;
  assign n6755 = ~n6748 & n6754;
  assign n6756 = n6748 & ~n6754;
  assign n6757 = ~n6755 & ~n6756;
  assign n6758 = n6742 & ~n6757;
  assign n6759 = ~n6742 & n6757;
  assign n6760 = ~n6758 & ~n6759;
  assign n6761 = ~n6727 & ~n6760;
  assign n6762 = pi94  & pi95 ;
  assign n6763 = pi96  & ~n6718;
  assign n6764 = ~n6762 & ~n6763;
  assign n6765 = pi91  & pi92 ;
  assign n6766 = pi93  & ~n6712;
  assign n6767 = ~n6765 & ~n6766;
  assign n6768 = ~n6764 & n6767;
  assign n6769 = n6764 & ~n6767;
  assign n6770 = ~n6768 & ~n6769;
  assign n6771 = ~n6715 & ~n6721;
  assign n6772 = n6770 & n6771;
  assign n6773 = ~n6770 & ~n6771;
  assign n6774 = ~n6772 & ~n6773;
  assign n6775 = pi100  & pi101 ;
  assign n6776 = pi102  & ~n6703;
  assign n6777 = ~n6775 & ~n6776;
  assign n6778 = pi97  & pi98 ;
  assign n6779 = pi99  & ~n6697;
  assign n6780 = ~n6778 & ~n6779;
  assign n6781 = ~n6777 & n6780;
  assign n6782 = n6777 & ~n6780;
  assign n6783 = ~n6781 & ~n6782;
  assign n6784 = ~n6700 & ~n6706;
  assign n6785 = n6783 & n6784;
  assign n6786 = ~n6783 & ~n6784;
  assign n6787 = ~n6785 & ~n6786;
  assign n6788 = ~n6783 & n6784;
  assign n6789 = ~n6777 & ~n6780;
  assign n6790 = ~n6788 & ~n6789;
  assign n6791 = ~n6787 & ~n6790;
  assign n6792 = ~n6770 & n6771;
  assign n6793 = ~n6764 & ~n6767;
  assign n6794 = ~n6792 & ~n6793;
  assign n6795 = ~n6774 & ~n6794;
  assign n6796 = ~n6709 & ~n6724;
  assign n6797 = ~n6791 & n6796;
  assign n6798 = ~n6795 & n6797;
  assign n6799 = n6787 & ~n6798;
  assign n6800 = ~n6787 & n6798;
  assign n6801 = ~n6799 & ~n6800;
  assign n6802 = ~n6774 & ~n6801;
  assign n6803 = n6774 & n6801;
  assign n6804 = ~n6802 & ~n6803;
  assign n6805 = n6761 & ~n6804;
  assign n6806 = pi82  & pi83 ;
  assign n6807 = pi84  & ~n6751;
  assign n6808 = ~n6806 & ~n6807;
  assign n6809 = pi79  & pi80 ;
  assign n6810 = pi81  & ~n6745;
  assign n6811 = ~n6809 & ~n6810;
  assign n6812 = ~n6808 & n6811;
  assign n6813 = n6808 & ~n6811;
  assign n6814 = ~n6812 & ~n6813;
  assign n6815 = ~n6748 & ~n6754;
  assign n6816 = n6814 & n6815;
  assign n6817 = ~n6814 & ~n6815;
  assign n6818 = ~n6816 & ~n6817;
  assign n6819 = pi88  & pi89 ;
  assign n6820 = pi90  & ~n6736;
  assign n6821 = ~n6819 & ~n6820;
  assign n6822 = pi85  & pi86 ;
  assign n6823 = pi87  & ~n6730;
  assign n6824 = ~n6822 & ~n6823;
  assign n6825 = ~n6821 & n6824;
  assign n6826 = n6821 & ~n6824;
  assign n6827 = ~n6825 & ~n6826;
  assign n6828 = ~n6733 & ~n6739;
  assign n6829 = n6827 & n6828;
  assign n6830 = ~n6827 & ~n6828;
  assign n6831 = ~n6829 & ~n6830;
  assign n6832 = ~n6827 & n6828;
  assign n6833 = ~n6821 & ~n6824;
  assign n6834 = ~n6832 & ~n6833;
  assign n6835 = ~n6831 & ~n6834;
  assign n6836 = ~n6814 & n6815;
  assign n6837 = ~n6808 & ~n6811;
  assign n6838 = ~n6836 & ~n6837;
  assign n6839 = ~n6818 & ~n6838;
  assign n6840 = ~n6742 & ~n6757;
  assign n6841 = ~n6835 & n6840;
  assign n6842 = ~n6839 & n6841;
  assign n6843 = n6831 & ~n6842;
  assign n6844 = ~n6831 & n6842;
  assign n6845 = ~n6843 & ~n6844;
  assign n6846 = n6818 & n6845;
  assign n6847 = ~n6818 & ~n6845;
  assign n6848 = ~n6846 & ~n6847;
  assign n6849 = ~n6761 & n6804;
  assign n6850 = ~n6848 & ~n6849;
  assign n6851 = ~n6805 & ~n6850;
  assign n6852 = ~n6818 & ~n6843;
  assign n6853 = ~n6844 & ~n6852;
  assign n6854 = n6834 & ~n6838;
  assign n6855 = ~n6834 & n6838;
  assign n6856 = ~n6854 & ~n6855;
  assign n6857 = ~n6853 & ~n6856;
  assign n6858 = n6853 & n6856;
  assign n6859 = ~n6857 & ~n6858;
  assign n6860 = ~n6774 & ~n6799;
  assign n6861 = ~n6800 & ~n6860;
  assign n6862 = n6790 & ~n6794;
  assign n6863 = ~n6790 & n6794;
  assign n6864 = ~n6862 & ~n6863;
  assign n6865 = ~n6861 & ~n6864;
  assign n6866 = n6861 & n6864;
  assign n6867 = ~n6865 & ~n6866;
  assign n6868 = ~n6859 & ~n6867;
  assign n6869 = ~n6851 & ~n6868;
  assign n6870 = n6859 & n6867;
  assign n6871 = ~n6869 & ~n6870;
  assign n6872 = n6790 & n6861;
  assign n6873 = ~n6794 & ~n6872;
  assign n6874 = ~n6790 & ~n6861;
  assign n6875 = ~n6873 & ~n6874;
  assign n6876 = n6834 & n6853;
  assign n6877 = ~n6838 & ~n6876;
  assign n6878 = ~n6834 & ~n6853;
  assign n6879 = ~n6877 & ~n6878;
  assign n6880 = n6875 & n6879;
  assign n6881 = ~n6871 & ~n6880;
  assign n6882 = ~n6875 & ~n6879;
  assign n6883 = ~n6881 & ~n6882;
  assign n6884 = ~n6694 & ~n6883;
  assign n6885 = ~n6868 & ~n6870;
  assign n6886 = ~n6851 & n6885;
  assign n6887 = n6851 & ~n6885;
  assign n6888 = ~n6886 & ~n6887;
  assign n6889 = n6687 & ~n6689;
  assign n6890 = ~n6690 & ~n6889;
  assign n6891 = n6888 & n6890;
  assign n6892 = ~n6671 & n6674;
  assign n6893 = n6671 & ~n6674;
  assign n6894 = ~n6892 & ~n6893;
  assign n6895 = ~n6727 & n6760;
  assign n6896 = n6727 & ~n6760;
  assign n6897 = ~n6895 & ~n6896;
  assign n6898 = ~n6894 & ~n6897;
  assign n6899 = ~n6680 & ~n6685;
  assign n6900 = ~n6684 & ~n6899;
  assign n6901 = n6684 & n6899;
  assign n6902 = ~n6900 & ~n6901;
  assign n6903 = n6898 & ~n6902;
  assign n6904 = ~n6805 & ~n6849;
  assign n6905 = n6848 & n6904;
  assign n6906 = ~n6848 & ~n6904;
  assign n6907 = ~n6905 & ~n6906;
  assign n6908 = ~n6898 & n6902;
  assign n6909 = ~n6907 & ~n6908;
  assign n6910 = ~n6903 & ~n6909;
  assign n6911 = ~n6888 & ~n6890;
  assign n6912 = ~n6891 & ~n6911;
  assign n6913 = ~n6910 & n6912;
  assign n6914 = ~n6891 & ~n6913;
  assign n6915 = ~n6655 & ~n6693;
  assign n6916 = ~n6691 & n6915;
  assign n6917 = n6691 & ~n6915;
  assign n6918 = ~n6916 & ~n6917;
  assign n6919 = n6875 & ~n6879;
  assign n6920 = ~n6875 & n6879;
  assign n6921 = ~n6870 & ~n6919;
  assign n6922 = ~n6920 & n6921;
  assign n6923 = ~n6869 & n6922;
  assign n6924 = n6881 & ~n6882;
  assign n6925 = ~n6923 & ~n6924;
  assign n6926 = ~n6918 & ~n6925;
  assign n6927 = ~n6914 & ~n6926;
  assign n6928 = n6918 & n6925;
  assign n6929 = ~n6927 & ~n6928;
  assign n6930 = n6694 & n6883;
  assign n6931 = ~n6884 & ~n6930;
  assign n6932 = ~n6929 & n6931;
  assign n6933 = ~n6884 & ~n6932;
  assign n6934 = ~n6504 & ~n6933;
  assign n6935 = n6504 & n6933;
  assign n6936 = ~n6934 & ~n6935;
  assign n6937 = n6929 & ~n6931;
  assign n6938 = ~n6932 & ~n6937;
  assign n6939 = n6500 & ~n6502;
  assign n6940 = ~n6503 & ~n6939;
  assign n6941 = n6938 & n6940;
  assign n6942 = ~n6465 & n6468;
  assign n6943 = n6465 & ~n6468;
  assign n6944 = ~n6942 & ~n6943;
  assign n6945 = ~n6894 & n6897;
  assign n6946 = n6894 & ~n6897;
  assign n6947 = ~n6945 & ~n6946;
  assign n6948 = ~n6944 & ~n6947;
  assign n6949 = ~n6474 & ~n6479;
  assign n6950 = ~n6478 & ~n6949;
  assign n6951 = n6478 & n6949;
  assign n6952 = ~n6950 & ~n6951;
  assign n6953 = n6948 & ~n6952;
  assign n6954 = ~n6903 & ~n6908;
  assign n6955 = n6907 & n6954;
  assign n6956 = ~n6907 & ~n6954;
  assign n6957 = ~n6955 & ~n6956;
  assign n6958 = ~n6948 & n6952;
  assign n6959 = ~n6957 & ~n6958;
  assign n6960 = ~n6953 & ~n6959;
  assign n6961 = n6910 & ~n6912;
  assign n6962 = ~n6913 & ~n6961;
  assign n6963 = n6481 & ~n6483;
  assign n6964 = ~n6484 & ~n6963;
  assign n6965 = ~n6962 & ~n6964;
  assign n6966 = ~n6960 & ~n6965;
  assign n6967 = n6962 & n6964;
  assign n6968 = ~n6966 & ~n6967;
  assign n6969 = ~n6497 & ~n6499;
  assign n6970 = ~n6485 & n6969;
  assign n6971 = n6485 & ~n6969;
  assign n6972 = ~n6970 & ~n6971;
  assign n6973 = ~n6926 & ~n6928;
  assign n6974 = ~n6914 & n6973;
  assign n6975 = n6914 & ~n6973;
  assign n6976 = ~n6974 & ~n6975;
  assign n6977 = ~n6972 & ~n6976;
  assign n6978 = ~n6968 & ~n6977;
  assign n6979 = n6972 & n6976;
  assign n6980 = ~n6978 & ~n6979;
  assign n6981 = ~n6938 & ~n6940;
  assign n6982 = ~n6941 & ~n6981;
  assign n6983 = ~n6980 & n6982;
  assign n6984 = ~n6941 & ~n6983;
  assign n6985 = n6936 & ~n6984;
  assign n6986 = ~n6934 & ~n6985;
  assign n6987 = ~n6075 & ~n6986;
  assign n6988 = n6075 & n6986;
  assign n6989 = ~n6987 & ~n6988;
  assign n6990 = ~n6022 & n6073;
  assign n6991 = ~n6074 & ~n6990;
  assign n6992 = ~n6936 & n6984;
  assign n6993 = ~n6985 & ~n6992;
  assign n6994 = n6991 & n6993;
  assign n6995 = ~n6066 & ~n6068;
  assign n6996 = ~n6057 & n6995;
  assign n6997 = n6057 & ~n6995;
  assign n6998 = ~n6996 & ~n6997;
  assign n6999 = ~n6977 & ~n6979;
  assign n7000 = ~n6968 & n6999;
  assign n7001 = n6968 & ~n6999;
  assign n7002 = ~n7000 & ~n7001;
  assign n7003 = n6998 & n7002;
  assign n7004 = ~n6965 & ~n6967;
  assign n7005 = ~n6960 & n7004;
  assign n7006 = n6960 & ~n7004;
  assign n7007 = ~n7005 & ~n7006;
  assign n7008 = n6053 & ~n6055;
  assign n7009 = ~n6056 & ~n7008;
  assign n7010 = n7007 & n7009;
  assign n7011 = ~n6037 & n6040;
  assign n7012 = n6037 & ~n6040;
  assign n7013 = ~n7011 & ~n7012;
  assign n7014 = ~n6944 & n6947;
  assign n7015 = n6944 & ~n6947;
  assign n7016 = ~n7014 & ~n7015;
  assign n7017 = ~n7013 & ~n7016;
  assign n7018 = ~n6046 & ~n6051;
  assign n7019 = n6050 & n7018;
  assign n7020 = ~n6050 & ~n7018;
  assign n7021 = ~n7019 & ~n7020;
  assign n7022 = n7017 & ~n7021;
  assign n7023 = ~n6953 & ~n6958;
  assign n7024 = n6957 & n7023;
  assign n7025 = ~n6957 & ~n7023;
  assign n7026 = ~n7024 & ~n7025;
  assign n7027 = ~n7017 & n7021;
  assign n7028 = ~n7026 & ~n7027;
  assign n7029 = ~n7022 & ~n7028;
  assign n7030 = ~n7007 & ~n7009;
  assign n7031 = ~n7010 & ~n7030;
  assign n7032 = ~n7029 & n7031;
  assign n7033 = ~n7010 & ~n7032;
  assign n7034 = ~n6998 & ~n7002;
  assign n7035 = ~n7033 & ~n7034;
  assign n7036 = ~n7003 & ~n7035;
  assign n7037 = n6980 & ~n6982;
  assign n7038 = ~n6983 & ~n7037;
  assign n7039 = n6069 & ~n6071;
  assign n7040 = ~n6072 & ~n7039;
  assign n7041 = ~n7038 & ~n7040;
  assign n7042 = ~n7036 & ~n7041;
  assign n7043 = n7038 & n7040;
  assign n7044 = ~n7042 & ~n7043;
  assign n7045 = ~n6991 & ~n6993;
  assign n7046 = ~n6994 & ~n7045;
  assign n7047 = ~n7044 & n7046;
  assign n7048 = ~n6994 & ~n7047;
  assign n7049 = n6989 & ~n7048;
  assign n7050 = ~n6987 & ~n7049;
  assign n7051 = ~n5156 & ~n7050;
  assign n7052 = n5156 & n7050;
  assign n7053 = ~n7051 & ~n7052;
  assign n7054 = ~n6989 & n7048;
  assign n7055 = ~n7049 & ~n7054;
  assign n7056 = ~n5098 & n5154;
  assign n7057 = ~n5155 & ~n7056;
  assign n7058 = n7055 & n7057;
  assign n7059 = ~n7041 & ~n7043;
  assign n7060 = ~n7036 & n7059;
  assign n7061 = n7036 & ~n7059;
  assign n7062 = ~n7060 & ~n7061;
  assign n7063 = ~n5147 & ~n5149;
  assign n7064 = ~n5142 & n7063;
  assign n7065 = n5142 & ~n7063;
  assign n7066 = ~n7064 & ~n7065;
  assign n7067 = n7062 & n7066;
  assign n7068 = n7029 & ~n7031;
  assign n7069 = ~n7032 & ~n7068;
  assign n7070 = ~n5136 & ~n5138;
  assign n7071 = ~n5131 & n7070;
  assign n7072 = n5131 & ~n7070;
  assign n7073 = ~n7071 & ~n7072;
  assign n7074 = n7069 & n7073;
  assign n7075 = ~n5115 & n5118;
  assign n7076 = n5115 & ~n5118;
  assign n7077 = ~n7075 & ~n7076;
  assign n7078 = ~n7013 & n7016;
  assign n7079 = n7013 & ~n7016;
  assign n7080 = ~n7078 & ~n7079;
  assign n7081 = ~n7077 & ~n7080;
  assign n7082 = ~n5124 & ~n5129;
  assign n7083 = n5128 & n7082;
  assign n7084 = ~n5128 & ~n7082;
  assign n7085 = ~n7083 & ~n7084;
  assign n7086 = n7081 & ~n7085;
  assign n7087 = ~n7022 & ~n7027;
  assign n7088 = n7026 & n7087;
  assign n7089 = ~n7026 & ~n7087;
  assign n7090 = ~n7088 & ~n7089;
  assign n7091 = ~n7081 & n7085;
  assign n7092 = ~n7090 & ~n7091;
  assign n7093 = ~n7086 & ~n7092;
  assign n7094 = ~n7069 & ~n7073;
  assign n7095 = ~n7074 & ~n7094;
  assign n7096 = ~n7093 & n7095;
  assign n7097 = ~n7074 & ~n7096;
  assign n7098 = ~n5112 & ~n5140;
  assign n7099 = ~n5139 & n7098;
  assign n7100 = n5139 & ~n7098;
  assign n7101 = ~n7099 & ~n7100;
  assign n7102 = ~n7003 & ~n7034;
  assign n7103 = ~n7033 & n7102;
  assign n7104 = n7033 & ~n7102;
  assign n7105 = ~n7103 & ~n7104;
  assign n7106 = ~n7101 & ~n7105;
  assign n7107 = ~n7097 & ~n7106;
  assign n7108 = n7101 & n7105;
  assign n7109 = ~n7107 & ~n7108;
  assign n7110 = ~n7062 & ~n7066;
  assign n7111 = ~n7067 & ~n7110;
  assign n7112 = ~n7109 & n7111;
  assign n7113 = ~n7067 & ~n7112;
  assign n7114 = n5150 & ~n5152;
  assign n7115 = ~n5153 & ~n7114;
  assign n7116 = n7044 & ~n7046;
  assign n7117 = ~n7047 & ~n7116;
  assign n7118 = ~n7115 & ~n7117;
  assign n7119 = ~n7113 & ~n7118;
  assign n7120 = n7115 & n7117;
  assign n7121 = ~n7119 & ~n7120;
  assign n7122 = ~n7055 & ~n7057;
  assign n7123 = ~n7058 & ~n7122;
  assign n7124 = ~n7121 & n7123;
  assign n7125 = ~n7058 & ~n7124;
  assign n7126 = n7053 & ~n7125;
  assign n7127 = ~n7051 & ~n7126;
  assign n7128 = n3259 & ~n7127;
  assign n7129 = ~n3259 & n7127;
  assign n7130 = ~n7128 & ~n7129;
  assign n7131 = ~n2304 & n3258;
  assign n7132 = ~n3259 & ~n7131;
  assign n7133 = ~n7053 & n7125;
  assign n7134 = ~n7126 & ~n7133;
  assign n7135 = n7132 & n7134;
  assign n7136 = ~n7118 & ~n7120;
  assign n7137 = ~n7113 & n7136;
  assign n7138 = n7113 & ~n7136;
  assign n7139 = ~n7137 & ~n7138;
  assign n7140 = n3250 & ~n3252;
  assign n7141 = ~n3253 & ~n7140;
  assign n7142 = n7139 & n7141;
  assign n7143 = ~n7106 & ~n7108;
  assign n7144 = ~n7097 & n7143;
  assign n7145 = n7097 & ~n7143;
  assign n7146 = ~n7144 & ~n7145;
  assign n7147 = ~n3243 & ~n3245;
  assign n7148 = ~n3236 & n7147;
  assign n7149 = n3236 & ~n7147;
  assign n7150 = ~n7148 & ~n7149;
  assign n7151 = n7146 & n7150;
  assign n7152 = ~n7077 & n7080;
  assign n7153 = n7077 & ~n7080;
  assign n7154 = ~n7152 & ~n7153;
  assign n7155 = ~n3218 & n3221;
  assign n7156 = n3218 & ~n3221;
  assign n7157 = ~n7155 & ~n7156;
  assign n7158 = ~n7154 & ~n7157;
  assign n7159 = ~n7086 & ~n7091;
  assign n7160 = ~n7090 & ~n7159;
  assign n7161 = n7090 & n7159;
  assign n7162 = ~n7160 & ~n7161;
  assign n7163 = n7158 & ~n7162;
  assign n7164 = ~n3227 & ~n3230;
  assign n7165 = n3229 & n7164;
  assign n7166 = ~n3229 & ~n7164;
  assign n7167 = ~n7165 & ~n7166;
  assign n7168 = ~n7158 & n7162;
  assign n7169 = ~n7167 & ~n7168;
  assign n7170 = ~n7163 & ~n7169;
  assign n7171 = n3232 & ~n3234;
  assign n7172 = ~n3235 & ~n7171;
  assign n7173 = n7093 & ~n7095;
  assign n7174 = ~n7096 & ~n7173;
  assign n7175 = ~n7172 & ~n7174;
  assign n7176 = ~n7170 & ~n7175;
  assign n7177 = n7172 & n7174;
  assign n7178 = ~n7176 & ~n7177;
  assign n7179 = ~n7146 & ~n7150;
  assign n7180 = ~n7178 & ~n7179;
  assign n7181 = ~n7151 & ~n7180;
  assign n7182 = n3246 & ~n3248;
  assign n7183 = ~n3249 & ~n7182;
  assign n7184 = n7109 & ~n7111;
  assign n7185 = ~n7112 & ~n7184;
  assign n7186 = ~n7183 & ~n7185;
  assign n7187 = ~n7181 & ~n7186;
  assign n7188 = n7183 & n7185;
  assign n7189 = ~n7187 & ~n7188;
  assign n7190 = ~n7139 & ~n7141;
  assign n7191 = ~n7142 & ~n7190;
  assign n7192 = ~n7189 & n7191;
  assign n7193 = ~n7142 & ~n7192;
  assign n7194 = n3254 & ~n3256;
  assign n7195 = ~n3257 & ~n7194;
  assign n7196 = n7121 & ~n7123;
  assign n7197 = ~n7124 & ~n7196;
  assign n7198 = ~n7195 & ~n7197;
  assign n7199 = ~n7193 & ~n7198;
  assign n7200 = n7195 & n7197;
  assign n7201 = ~n7199 & ~n7200;
  assign n7202 = ~n7132 & ~n7134;
  assign n7203 = ~n7135 & ~n7202;
  assign n7204 = ~n7201 & n7203;
  assign n7205 = ~n7135 & ~n7204;
  assign n7206 = n7130 & ~n7205;
  assign n7207 = ~n7128 & ~n7206;
  assign n7208 = ~n7130 & n7205;
  assign n7209 = ~n7206 & ~n7208;
  assign n7210 = pi835  & ~pi836 ;
  assign n7211 = ~pi835  & pi836 ;
  assign n7212 = ~n7210 & ~n7211;
  assign n7213 = ~pi837  & ~n7212;
  assign n7214 = pi837  & n7212;
  assign n7215 = ~n7213 & ~n7214;
  assign n7216 = pi838  & ~pi839 ;
  assign n7217 = ~pi838  & pi839 ;
  assign n7218 = ~n7216 & ~n7217;
  assign n7219 = ~pi840  & ~n7218;
  assign n7220 = pi840  & n7218;
  assign n7221 = ~n7219 & ~n7220;
  assign n7222 = ~n7215 & ~n7221;
  assign n7223 = pi838  & pi839 ;
  assign n7224 = pi840  & ~n7218;
  assign n7225 = ~n7223 & ~n7224;
  assign n7226 = pi835  & pi836 ;
  assign n7227 = pi837  & ~n7212;
  assign n7228 = ~n7226 & ~n7227;
  assign n7229 = n7225 & ~n7228;
  assign n7230 = ~n7225 & n7228;
  assign n7231 = ~n7229 & ~n7230;
  assign n7232 = n7222 & ~n7231;
  assign n7233 = ~n7225 & ~n7228;
  assign n7234 = ~n7232 & ~n7233;
  assign n7235 = pi844  & pi845 ;
  assign n7236 = pi844  & ~pi845 ;
  assign n7237 = ~pi844  & pi845 ;
  assign n7238 = ~n7236 & ~n7237;
  assign n7239 = pi846  & ~n7238;
  assign n7240 = ~n7235 & ~n7239;
  assign n7241 = pi841  & pi842 ;
  assign n7242 = pi841  & ~pi842 ;
  assign n7243 = ~pi841  & pi842 ;
  assign n7244 = ~n7242 & ~n7243;
  assign n7245 = pi843  & ~n7244;
  assign n7246 = ~n7241 & ~n7245;
  assign n7247 = ~n7240 & n7246;
  assign n7248 = n7240 & ~n7246;
  assign n7249 = ~n7247 & ~n7248;
  assign n7250 = ~pi843  & ~n7244;
  assign n7251 = pi843  & n7244;
  assign n7252 = ~n7250 & ~n7251;
  assign n7253 = ~pi846  & ~n7238;
  assign n7254 = pi846  & n7238;
  assign n7255 = ~n7253 & ~n7254;
  assign n7256 = ~n7252 & ~n7255;
  assign n7257 = ~n7249 & n7256;
  assign n7258 = ~n7240 & ~n7246;
  assign n7259 = ~n7257 & ~n7258;
  assign n7260 = n7249 & n7256;
  assign n7261 = ~n7249 & ~n7256;
  assign n7262 = ~n7260 & ~n7261;
  assign n7263 = ~n7259 & ~n7262;
  assign n7264 = n7222 & n7231;
  assign n7265 = ~n7222 & ~n7231;
  assign n7266 = ~n7264 & ~n7265;
  assign n7267 = ~n7234 & ~n7266;
  assign n7268 = ~n7215 & n7221;
  assign n7269 = n7215 & ~n7221;
  assign n7270 = ~n7268 & ~n7269;
  assign n7271 = ~n7252 & n7255;
  assign n7272 = n7252 & ~n7255;
  assign n7273 = ~n7271 & ~n7272;
  assign n7274 = ~n7270 & ~n7273;
  assign n7275 = ~n7263 & n7274;
  assign n7276 = ~n7267 & n7275;
  assign n7277 = n7262 & ~n7276;
  assign n7278 = ~n7262 & n7276;
  assign n7279 = ~n7277 & ~n7278;
  assign n7280 = n7266 & n7279;
  assign n7281 = ~n7277 & ~n7280;
  assign n7282 = n7259 & ~n7281;
  assign n7283 = ~n7234 & ~n7282;
  assign n7284 = ~n7259 & n7281;
  assign n7285 = ~n7283 & ~n7284;
  assign n7286 = pi823  & ~pi824 ;
  assign n7287 = ~pi823  & pi824 ;
  assign n7288 = ~n7286 & ~n7287;
  assign n7289 = ~pi825  & ~n7288;
  assign n7290 = pi825  & n7288;
  assign n7291 = ~n7289 & ~n7290;
  assign n7292 = pi826  & ~pi827 ;
  assign n7293 = ~pi826  & pi827 ;
  assign n7294 = ~n7292 & ~n7293;
  assign n7295 = ~pi828  & ~n7294;
  assign n7296 = pi828  & n7294;
  assign n7297 = ~n7295 & ~n7296;
  assign n7298 = ~n7291 & ~n7297;
  assign n7299 = pi826  & pi827 ;
  assign n7300 = pi828  & ~n7294;
  assign n7301 = ~n7299 & ~n7300;
  assign n7302 = pi823  & pi824 ;
  assign n7303 = pi825  & ~n7288;
  assign n7304 = ~n7302 & ~n7303;
  assign n7305 = n7301 & ~n7304;
  assign n7306 = ~n7301 & n7304;
  assign n7307 = ~n7305 & ~n7306;
  assign n7308 = n7298 & ~n7307;
  assign n7309 = ~n7301 & ~n7304;
  assign n7310 = ~n7308 & ~n7309;
  assign n7311 = pi832  & pi833 ;
  assign n7312 = pi832  & ~pi833 ;
  assign n7313 = ~pi832  & pi833 ;
  assign n7314 = ~n7312 & ~n7313;
  assign n7315 = pi834  & ~n7314;
  assign n7316 = ~n7311 & ~n7315;
  assign n7317 = pi829  & pi830 ;
  assign n7318 = pi829  & ~pi830 ;
  assign n7319 = ~pi829  & pi830 ;
  assign n7320 = ~n7318 & ~n7319;
  assign n7321 = pi831  & ~n7320;
  assign n7322 = ~n7317 & ~n7321;
  assign n7323 = ~n7316 & n7322;
  assign n7324 = n7316 & ~n7322;
  assign n7325 = ~n7323 & ~n7324;
  assign n7326 = ~pi831  & ~n7320;
  assign n7327 = pi831  & n7320;
  assign n7328 = ~n7326 & ~n7327;
  assign n7329 = ~pi834  & ~n7314;
  assign n7330 = pi834  & n7314;
  assign n7331 = ~n7329 & ~n7330;
  assign n7332 = ~n7328 & ~n7331;
  assign n7333 = ~n7325 & n7332;
  assign n7334 = ~n7316 & ~n7322;
  assign n7335 = ~n7333 & ~n7334;
  assign n7336 = n7325 & n7332;
  assign n7337 = ~n7325 & ~n7332;
  assign n7338 = ~n7336 & ~n7337;
  assign n7339 = ~n7335 & ~n7338;
  assign n7340 = n7298 & n7307;
  assign n7341 = ~n7298 & ~n7307;
  assign n7342 = ~n7340 & ~n7341;
  assign n7343 = ~n7310 & ~n7342;
  assign n7344 = ~n7291 & n7297;
  assign n7345 = n7291 & ~n7297;
  assign n7346 = ~n7344 & ~n7345;
  assign n7347 = ~n7328 & n7331;
  assign n7348 = n7328 & ~n7331;
  assign n7349 = ~n7347 & ~n7348;
  assign n7350 = ~n7346 & ~n7349;
  assign n7351 = ~n7339 & n7350;
  assign n7352 = ~n7343 & n7351;
  assign n7353 = n7338 & ~n7352;
  assign n7354 = ~n7338 & n7352;
  assign n7355 = ~n7353 & ~n7354;
  assign n7356 = n7342 & n7355;
  assign n7357 = ~n7353 & ~n7356;
  assign n7358 = n7335 & ~n7357;
  assign n7359 = ~n7310 & ~n7358;
  assign n7360 = ~n7335 & n7357;
  assign n7361 = ~n7359 & ~n7360;
  assign n7362 = n7285 & n7361;
  assign n7363 = ~n7310 & n7335;
  assign n7364 = n7310 & ~n7335;
  assign n7365 = ~n7363 & ~n7364;
  assign n7366 = n7357 & ~n7365;
  assign n7367 = ~n7357 & n7365;
  assign n7368 = ~n7366 & ~n7367;
  assign n7369 = ~n7234 & n7259;
  assign n7370 = n7234 & ~n7259;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = n7281 & ~n7371;
  assign n7373 = ~n7281 & n7371;
  assign n7374 = ~n7372 & ~n7373;
  assign n7375 = n7368 & n7374;
  assign n7376 = ~n7270 & n7273;
  assign n7377 = n7270 & ~n7273;
  assign n7378 = ~n7376 & ~n7377;
  assign n7379 = ~n7346 & n7349;
  assign n7380 = n7346 & ~n7349;
  assign n7381 = ~n7379 & ~n7380;
  assign n7382 = ~n7378 & ~n7381;
  assign n7383 = ~n7266 & ~n7279;
  assign n7384 = ~n7280 & ~n7383;
  assign n7385 = ~n7382 & n7384;
  assign n7386 = ~n7342 & ~n7355;
  assign n7387 = ~n7356 & ~n7386;
  assign n7388 = ~n7382 & ~n7384;
  assign n7389 = n7384 & ~n7385;
  assign n7390 = ~n7388 & ~n7389;
  assign n7391 = n7387 & ~n7390;
  assign n7392 = ~n7385 & ~n7391;
  assign n7393 = ~n7368 & ~n7374;
  assign n7394 = ~n7375 & ~n7393;
  assign n7395 = n7392 & n7394;
  assign n7396 = ~n7375 & ~n7395;
  assign n7397 = ~n7362 & ~n7396;
  assign n7398 = ~n7285 & ~n7361;
  assign n7399 = ~n7397 & ~n7398;
  assign n7400 = pi811  & ~pi812 ;
  assign n7401 = ~pi811  & pi812 ;
  assign n7402 = ~n7400 & ~n7401;
  assign n7403 = ~pi813  & ~n7402;
  assign n7404 = pi813  & n7402;
  assign n7405 = ~n7403 & ~n7404;
  assign n7406 = pi814  & ~pi815 ;
  assign n7407 = ~pi814  & pi815 ;
  assign n7408 = ~n7406 & ~n7407;
  assign n7409 = ~pi816  & ~n7408;
  assign n7410 = pi816  & n7408;
  assign n7411 = ~n7409 & ~n7410;
  assign n7412 = ~n7405 & ~n7411;
  assign n7413 = pi814  & pi815 ;
  assign n7414 = pi816  & ~n7408;
  assign n7415 = ~n7413 & ~n7414;
  assign n7416 = pi811  & pi812 ;
  assign n7417 = pi813  & ~n7402;
  assign n7418 = ~n7416 & ~n7417;
  assign n7419 = n7415 & ~n7418;
  assign n7420 = ~n7415 & n7418;
  assign n7421 = ~n7419 & ~n7420;
  assign n7422 = n7412 & ~n7421;
  assign n7423 = ~n7415 & ~n7418;
  assign n7424 = ~n7422 & ~n7423;
  assign n7425 = pi820  & pi821 ;
  assign n7426 = pi820  & ~pi821 ;
  assign n7427 = ~pi820  & pi821 ;
  assign n7428 = ~n7426 & ~n7427;
  assign n7429 = pi822  & ~n7428;
  assign n7430 = ~n7425 & ~n7429;
  assign n7431 = pi817  & pi818 ;
  assign n7432 = pi817  & ~pi818 ;
  assign n7433 = ~pi817  & pi818 ;
  assign n7434 = ~n7432 & ~n7433;
  assign n7435 = pi819  & ~n7434;
  assign n7436 = ~n7431 & ~n7435;
  assign n7437 = ~n7430 & n7436;
  assign n7438 = n7430 & ~n7436;
  assign n7439 = ~n7437 & ~n7438;
  assign n7440 = ~pi819  & ~n7434;
  assign n7441 = pi819  & n7434;
  assign n7442 = ~n7440 & ~n7441;
  assign n7443 = ~pi822  & ~n7428;
  assign n7444 = pi822  & n7428;
  assign n7445 = ~n7443 & ~n7444;
  assign n7446 = ~n7442 & ~n7445;
  assign n7447 = ~n7439 & n7446;
  assign n7448 = ~n7430 & ~n7436;
  assign n7449 = ~n7447 & ~n7448;
  assign n7450 = n7439 & n7446;
  assign n7451 = ~n7439 & ~n7446;
  assign n7452 = ~n7450 & ~n7451;
  assign n7453 = ~n7449 & ~n7452;
  assign n7454 = n7412 & n7421;
  assign n7455 = ~n7412 & ~n7421;
  assign n7456 = ~n7454 & ~n7455;
  assign n7457 = ~n7424 & ~n7456;
  assign n7458 = ~n7405 & n7411;
  assign n7459 = n7405 & ~n7411;
  assign n7460 = ~n7458 & ~n7459;
  assign n7461 = ~n7442 & n7445;
  assign n7462 = n7442 & ~n7445;
  assign n7463 = ~n7461 & ~n7462;
  assign n7464 = ~n7460 & ~n7463;
  assign n7465 = ~n7453 & n7464;
  assign n7466 = ~n7457 & n7465;
  assign n7467 = n7452 & ~n7466;
  assign n7468 = ~n7452 & n7466;
  assign n7469 = ~n7467 & ~n7468;
  assign n7470 = n7456 & n7469;
  assign n7471 = ~n7467 & ~n7470;
  assign n7472 = n7449 & ~n7471;
  assign n7473 = ~n7424 & ~n7472;
  assign n7474 = ~n7449 & n7471;
  assign n7475 = ~n7473 & ~n7474;
  assign n7476 = pi802  & pi803 ;
  assign n7477 = ~pi802  & pi803 ;
  assign n7478 = pi802  & ~pi803 ;
  assign n7479 = ~n7477 & ~n7478;
  assign n7480 = pi804  & ~n7479;
  assign n7481 = ~n7476 & ~n7480;
  assign n7482 = pi799  & pi800 ;
  assign n7483 = ~pi799  & pi800 ;
  assign n7484 = pi799  & ~pi800 ;
  assign n7485 = ~n7483 & ~n7484;
  assign n7486 = pi801  & ~n7485;
  assign n7487 = ~n7482 & ~n7486;
  assign n7488 = ~n7481 & n7487;
  assign n7489 = n7481 & ~n7487;
  assign n7490 = ~n7488 & ~n7489;
  assign n7491 = ~pi801  & ~n7485;
  assign n7492 = pi801  & n7485;
  assign n7493 = ~n7491 & ~n7492;
  assign n7494 = ~pi804  & ~n7479;
  assign n7495 = pi804  & n7479;
  assign n7496 = ~n7494 & ~n7495;
  assign n7497 = ~n7493 & ~n7496;
  assign n7498 = ~n7490 & n7497;
  assign n7499 = ~n7481 & ~n7487;
  assign n7500 = ~n7498 & ~n7499;
  assign n7501 = pi808  & pi809 ;
  assign n7502 = ~pi808  & pi809 ;
  assign n7503 = pi808  & ~pi809 ;
  assign n7504 = ~n7502 & ~n7503;
  assign n7505 = pi810  & ~n7504;
  assign n7506 = ~n7501 & ~n7505;
  assign n7507 = pi805  & pi806 ;
  assign n7508 = ~pi805  & pi806 ;
  assign n7509 = pi805  & ~pi806 ;
  assign n7510 = ~n7508 & ~n7509;
  assign n7511 = pi807  & ~n7510;
  assign n7512 = ~n7507 & ~n7511;
  assign n7513 = ~n7506 & n7512;
  assign n7514 = n7506 & ~n7512;
  assign n7515 = ~n7513 & ~n7514;
  assign n7516 = ~pi807  & ~n7510;
  assign n7517 = pi807  & n7510;
  assign n7518 = ~n7516 & ~n7517;
  assign n7519 = ~pi810  & ~n7504;
  assign n7520 = pi810  & n7504;
  assign n7521 = ~n7519 & ~n7520;
  assign n7522 = ~n7518 & ~n7521;
  assign n7523 = ~n7515 & n7522;
  assign n7524 = ~n7506 & ~n7512;
  assign n7525 = ~n7523 & ~n7524;
  assign n7526 = n7515 & n7522;
  assign n7527 = ~n7515 & ~n7522;
  assign n7528 = ~n7526 & ~n7527;
  assign n7529 = n7490 & n7497;
  assign n7530 = ~n7490 & ~n7497;
  assign n7531 = ~n7529 & ~n7530;
  assign n7532 = ~n7500 & ~n7531;
  assign n7533 = ~n7525 & ~n7528;
  assign n7534 = ~n7518 & n7521;
  assign n7535 = n7518 & ~n7521;
  assign n7536 = ~n7534 & ~n7535;
  assign n7537 = ~n7493 & n7496;
  assign n7538 = n7493 & ~n7496;
  assign n7539 = ~n7537 & ~n7538;
  assign n7540 = ~n7536 & ~n7539;
  assign n7541 = ~n7532 & n7540;
  assign n7542 = ~n7533 & n7541;
  assign n7543 = n7528 & ~n7542;
  assign n7544 = ~n7528 & n7542;
  assign n7545 = ~n7543 & ~n7544;
  assign n7546 = n7531 & n7545;
  assign n7547 = ~n7543 & ~n7546;
  assign n7548 = n7525 & ~n7547;
  assign n7549 = ~n7500 & ~n7548;
  assign n7550 = ~n7525 & n7547;
  assign n7551 = ~n7549 & ~n7550;
  assign n7552 = n7475 & n7551;
  assign n7553 = ~n7500 & n7525;
  assign n7554 = n7500 & ~n7525;
  assign n7555 = ~n7553 & ~n7554;
  assign n7556 = n7547 & ~n7555;
  assign n7557 = ~n7547 & n7555;
  assign n7558 = ~n7556 & ~n7557;
  assign n7559 = ~n7424 & n7449;
  assign n7560 = n7424 & ~n7449;
  assign n7561 = ~n7559 & ~n7560;
  assign n7562 = n7471 & ~n7561;
  assign n7563 = ~n7471 & n7561;
  assign n7564 = ~n7562 & ~n7563;
  assign n7565 = n7558 & n7564;
  assign n7566 = ~n7460 & n7463;
  assign n7567 = n7460 & ~n7463;
  assign n7568 = ~n7566 & ~n7567;
  assign n7569 = n7536 & ~n7539;
  assign n7570 = ~n7536 & n7539;
  assign n7571 = ~n7569 & ~n7570;
  assign n7572 = ~n7568 & ~n7571;
  assign n7573 = ~n7456 & ~n7469;
  assign n7574 = ~n7470 & ~n7573;
  assign n7575 = ~n7572 & n7574;
  assign n7576 = ~n7531 & ~n7545;
  assign n7577 = ~n7546 & ~n7576;
  assign n7578 = n7572 & ~n7574;
  assign n7579 = ~n7575 & ~n7578;
  assign n7580 = n7577 & n7579;
  assign n7581 = ~n7575 & ~n7580;
  assign n7582 = ~n7558 & ~n7564;
  assign n7583 = ~n7565 & ~n7582;
  assign n7584 = n7581 & n7583;
  assign n7585 = ~n7565 & ~n7584;
  assign n7586 = ~n7552 & ~n7585;
  assign n7587 = ~n7475 & ~n7551;
  assign n7588 = ~n7586 & ~n7587;
  assign n7589 = ~n7399 & ~n7588;
  assign n7590 = n7399 & n7588;
  assign n7591 = ~n7589 & ~n7590;
  assign n7592 = ~n7362 & ~n7398;
  assign n7593 = ~n7396 & n7592;
  assign n7594 = n7396 & ~n7592;
  assign n7595 = ~n7593 & ~n7594;
  assign n7596 = ~n7552 & ~n7587;
  assign n7597 = ~n7585 & n7596;
  assign n7598 = n7585 & ~n7596;
  assign n7599 = ~n7597 & ~n7598;
  assign n7600 = n7595 & n7599;
  assign n7601 = ~n7581 & ~n7583;
  assign n7602 = ~n7584 & ~n7601;
  assign n7603 = ~n7392 & ~n7394;
  assign n7604 = ~n7395 & ~n7603;
  assign n7605 = n7602 & n7604;
  assign n7606 = ~n7602 & ~n7604;
  assign n7607 = ~n7605 & ~n7606;
  assign n7608 = ~n7378 & n7381;
  assign n7609 = n7378 & ~n7381;
  assign n7610 = ~n7608 & ~n7609;
  assign n7611 = ~n7568 & n7571;
  assign n7612 = n7568 & ~n7571;
  assign n7613 = ~n7611 & ~n7612;
  assign n7614 = ~n7610 & ~n7613;
  assign n7615 = ~n7387 & n7390;
  assign n7616 = ~n7391 & ~n7615;
  assign n7617 = ~n7614 & n7616;
  assign n7618 = ~n7577 & ~n7579;
  assign n7619 = ~n7580 & ~n7618;
  assign n7620 = n7614 & ~n7616;
  assign n7621 = ~n7617 & ~n7620;
  assign n7622 = n7619 & n7621;
  assign n7623 = ~n7617 & ~n7622;
  assign n7624 = n7607 & n7623;
  assign n7625 = ~n7605 & ~n7624;
  assign n7626 = ~n7595 & ~n7599;
  assign n7627 = ~n7600 & ~n7626;
  assign n7628 = ~n7625 & n7627;
  assign n7629 = ~n7600 & ~n7628;
  assign n7630 = n7591 & ~n7629;
  assign n7631 = ~n7589 & ~n7630;
  assign n7632 = pi787  & ~pi788 ;
  assign n7633 = ~pi787  & pi788 ;
  assign n7634 = ~n7632 & ~n7633;
  assign n7635 = ~pi789  & ~n7634;
  assign n7636 = pi789  & n7634;
  assign n7637 = ~n7635 & ~n7636;
  assign n7638 = pi790  & ~pi791 ;
  assign n7639 = ~pi790  & pi791 ;
  assign n7640 = ~n7638 & ~n7639;
  assign n7641 = ~pi792  & ~n7640;
  assign n7642 = pi792  & n7640;
  assign n7643 = ~n7641 & ~n7642;
  assign n7644 = ~n7637 & ~n7643;
  assign n7645 = pi790  & pi791 ;
  assign n7646 = pi792  & ~n7640;
  assign n7647 = ~n7645 & ~n7646;
  assign n7648 = pi787  & pi788 ;
  assign n7649 = pi789  & ~n7634;
  assign n7650 = ~n7648 & ~n7649;
  assign n7651 = n7647 & ~n7650;
  assign n7652 = ~n7647 & n7650;
  assign n7653 = ~n7651 & ~n7652;
  assign n7654 = n7644 & ~n7653;
  assign n7655 = ~n7647 & ~n7650;
  assign n7656 = ~n7654 & ~n7655;
  assign n7657 = pi796  & pi797 ;
  assign n7658 = pi796  & ~pi797 ;
  assign n7659 = ~pi796  & pi797 ;
  assign n7660 = ~n7658 & ~n7659;
  assign n7661 = pi798  & ~n7660;
  assign n7662 = ~n7657 & ~n7661;
  assign n7663 = pi793  & pi794 ;
  assign n7664 = pi793  & ~pi794 ;
  assign n7665 = ~pi793  & pi794 ;
  assign n7666 = ~n7664 & ~n7665;
  assign n7667 = pi795  & ~n7666;
  assign n7668 = ~n7663 & ~n7667;
  assign n7669 = ~n7662 & n7668;
  assign n7670 = n7662 & ~n7668;
  assign n7671 = ~n7669 & ~n7670;
  assign n7672 = ~pi795  & ~n7666;
  assign n7673 = pi795  & n7666;
  assign n7674 = ~n7672 & ~n7673;
  assign n7675 = ~pi798  & ~n7660;
  assign n7676 = pi798  & n7660;
  assign n7677 = ~n7675 & ~n7676;
  assign n7678 = ~n7674 & ~n7677;
  assign n7679 = ~n7671 & n7678;
  assign n7680 = ~n7662 & ~n7668;
  assign n7681 = ~n7679 & ~n7680;
  assign n7682 = n7671 & n7678;
  assign n7683 = ~n7671 & ~n7678;
  assign n7684 = ~n7682 & ~n7683;
  assign n7685 = ~n7681 & ~n7684;
  assign n7686 = n7644 & n7653;
  assign n7687 = ~n7644 & ~n7653;
  assign n7688 = ~n7686 & ~n7687;
  assign n7689 = ~n7656 & ~n7688;
  assign n7690 = ~n7637 & n7643;
  assign n7691 = n7637 & ~n7643;
  assign n7692 = ~n7690 & ~n7691;
  assign n7693 = ~n7674 & n7677;
  assign n7694 = n7674 & ~n7677;
  assign n7695 = ~n7693 & ~n7694;
  assign n7696 = ~n7692 & ~n7695;
  assign n7697 = ~n7685 & n7696;
  assign n7698 = ~n7689 & n7697;
  assign n7699 = n7684 & ~n7698;
  assign n7700 = ~n7684 & n7698;
  assign n7701 = ~n7699 & ~n7700;
  assign n7702 = n7688 & n7701;
  assign n7703 = ~n7699 & ~n7702;
  assign n7704 = n7681 & ~n7703;
  assign n7705 = ~n7656 & ~n7704;
  assign n7706 = ~n7681 & n7703;
  assign n7707 = ~n7705 & ~n7706;
  assign n7708 = pi775  & ~pi776 ;
  assign n7709 = ~pi775  & pi776 ;
  assign n7710 = ~n7708 & ~n7709;
  assign n7711 = ~pi777  & ~n7710;
  assign n7712 = pi777  & n7710;
  assign n7713 = ~n7711 & ~n7712;
  assign n7714 = pi778  & ~pi779 ;
  assign n7715 = ~pi778  & pi779 ;
  assign n7716 = ~n7714 & ~n7715;
  assign n7717 = ~pi780  & ~n7716;
  assign n7718 = pi780  & n7716;
  assign n7719 = ~n7717 & ~n7718;
  assign n7720 = ~n7713 & ~n7719;
  assign n7721 = pi778  & pi779 ;
  assign n7722 = pi780  & ~n7716;
  assign n7723 = ~n7721 & ~n7722;
  assign n7724 = pi775  & pi776 ;
  assign n7725 = pi777  & ~n7710;
  assign n7726 = ~n7724 & ~n7725;
  assign n7727 = n7723 & ~n7726;
  assign n7728 = ~n7723 & n7726;
  assign n7729 = ~n7727 & ~n7728;
  assign n7730 = n7720 & ~n7729;
  assign n7731 = ~n7723 & ~n7726;
  assign n7732 = ~n7730 & ~n7731;
  assign n7733 = pi784  & pi785 ;
  assign n7734 = pi784  & ~pi785 ;
  assign n7735 = ~pi784  & pi785 ;
  assign n7736 = ~n7734 & ~n7735;
  assign n7737 = pi786  & ~n7736;
  assign n7738 = ~n7733 & ~n7737;
  assign n7739 = pi781  & pi782 ;
  assign n7740 = pi781  & ~pi782 ;
  assign n7741 = ~pi781  & pi782 ;
  assign n7742 = ~n7740 & ~n7741;
  assign n7743 = pi783  & ~n7742;
  assign n7744 = ~n7739 & ~n7743;
  assign n7745 = ~n7738 & n7744;
  assign n7746 = n7738 & ~n7744;
  assign n7747 = ~n7745 & ~n7746;
  assign n7748 = ~pi783  & ~n7742;
  assign n7749 = pi783  & n7742;
  assign n7750 = ~n7748 & ~n7749;
  assign n7751 = ~pi786  & ~n7736;
  assign n7752 = pi786  & n7736;
  assign n7753 = ~n7751 & ~n7752;
  assign n7754 = ~n7750 & ~n7753;
  assign n7755 = ~n7747 & n7754;
  assign n7756 = ~n7738 & ~n7744;
  assign n7757 = ~n7755 & ~n7756;
  assign n7758 = n7747 & n7754;
  assign n7759 = ~n7747 & ~n7754;
  assign n7760 = ~n7758 & ~n7759;
  assign n7761 = ~n7757 & ~n7760;
  assign n7762 = n7720 & n7729;
  assign n7763 = ~n7720 & ~n7729;
  assign n7764 = ~n7762 & ~n7763;
  assign n7765 = ~n7732 & ~n7764;
  assign n7766 = ~n7713 & n7719;
  assign n7767 = n7713 & ~n7719;
  assign n7768 = ~n7766 & ~n7767;
  assign n7769 = ~n7750 & n7753;
  assign n7770 = n7750 & ~n7753;
  assign n7771 = ~n7769 & ~n7770;
  assign n7772 = ~n7768 & ~n7771;
  assign n7773 = ~n7761 & n7772;
  assign n7774 = ~n7765 & n7773;
  assign n7775 = n7760 & ~n7774;
  assign n7776 = ~n7760 & n7774;
  assign n7777 = ~n7775 & ~n7776;
  assign n7778 = n7764 & n7777;
  assign n7779 = ~n7775 & ~n7778;
  assign n7780 = n7757 & ~n7779;
  assign n7781 = ~n7732 & ~n7780;
  assign n7782 = ~n7757 & n7779;
  assign n7783 = ~n7781 & ~n7782;
  assign n7784 = n7707 & n7783;
  assign n7785 = ~n7732 & n7757;
  assign n7786 = n7732 & ~n7757;
  assign n7787 = ~n7785 & ~n7786;
  assign n7788 = n7779 & ~n7787;
  assign n7789 = ~n7779 & n7787;
  assign n7790 = ~n7788 & ~n7789;
  assign n7791 = ~n7656 & n7681;
  assign n7792 = n7656 & ~n7681;
  assign n7793 = ~n7791 & ~n7792;
  assign n7794 = n7703 & ~n7793;
  assign n7795 = ~n7703 & n7793;
  assign n7796 = ~n7794 & ~n7795;
  assign n7797 = n7790 & n7796;
  assign n7798 = ~n7692 & n7695;
  assign n7799 = n7692 & ~n7695;
  assign n7800 = ~n7798 & ~n7799;
  assign n7801 = ~n7768 & n7771;
  assign n7802 = n7768 & ~n7771;
  assign n7803 = ~n7801 & ~n7802;
  assign n7804 = ~n7800 & ~n7803;
  assign n7805 = ~n7688 & ~n7701;
  assign n7806 = ~n7702 & ~n7805;
  assign n7807 = ~n7804 & n7806;
  assign n7808 = ~n7764 & ~n7777;
  assign n7809 = ~n7778 & ~n7808;
  assign n7810 = ~n7804 & ~n7806;
  assign n7811 = n7806 & ~n7807;
  assign n7812 = ~n7810 & ~n7811;
  assign n7813 = n7809 & ~n7812;
  assign n7814 = ~n7807 & ~n7813;
  assign n7815 = ~n7790 & ~n7796;
  assign n7816 = ~n7797 & ~n7815;
  assign n7817 = n7814 & n7816;
  assign n7818 = ~n7797 & ~n7817;
  assign n7819 = ~n7784 & ~n7818;
  assign n7820 = ~n7707 & ~n7783;
  assign n7821 = ~n7819 & ~n7820;
  assign n7822 = pi766  & pi767 ;
  assign n7823 = ~pi766  & pi767 ;
  assign n7824 = pi766  & ~pi767 ;
  assign n7825 = ~n7823 & ~n7824;
  assign n7826 = pi768  & ~n7825;
  assign n7827 = ~n7822 & ~n7826;
  assign n7828 = pi763  & pi764 ;
  assign n7829 = ~pi763  & pi764 ;
  assign n7830 = pi763  & ~pi764 ;
  assign n7831 = ~n7829 & ~n7830;
  assign n7832 = pi765  & ~n7831;
  assign n7833 = ~n7828 & ~n7832;
  assign n7834 = ~n7827 & n7833;
  assign n7835 = n7827 & ~n7833;
  assign n7836 = ~n7834 & ~n7835;
  assign n7837 = ~pi765  & ~n7831;
  assign n7838 = pi765  & n7831;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = ~pi768  & ~n7825;
  assign n7841 = pi768  & n7825;
  assign n7842 = ~n7840 & ~n7841;
  assign n7843 = ~n7839 & ~n7842;
  assign n7844 = ~n7836 & n7843;
  assign n7845 = ~n7827 & ~n7833;
  assign n7846 = ~n7844 & ~n7845;
  assign n7847 = pi772  & pi773 ;
  assign n7848 = ~pi772  & pi773 ;
  assign n7849 = pi772  & ~pi773 ;
  assign n7850 = ~n7848 & ~n7849;
  assign n7851 = pi774  & ~n7850;
  assign n7852 = ~n7847 & ~n7851;
  assign n7853 = pi769  & pi770 ;
  assign n7854 = ~pi769  & pi770 ;
  assign n7855 = pi769  & ~pi770 ;
  assign n7856 = ~n7854 & ~n7855;
  assign n7857 = pi771  & ~n7856;
  assign n7858 = ~n7853 & ~n7857;
  assign n7859 = ~n7852 & n7858;
  assign n7860 = n7852 & ~n7858;
  assign n7861 = ~n7859 & ~n7860;
  assign n7862 = ~pi771  & ~n7856;
  assign n7863 = pi771  & n7856;
  assign n7864 = ~n7862 & ~n7863;
  assign n7865 = ~pi774  & ~n7850;
  assign n7866 = pi774  & n7850;
  assign n7867 = ~n7865 & ~n7866;
  assign n7868 = ~n7864 & ~n7867;
  assign n7869 = ~n7861 & n7868;
  assign n7870 = ~n7852 & ~n7858;
  assign n7871 = ~n7869 & ~n7870;
  assign n7872 = n7861 & n7868;
  assign n7873 = ~n7861 & ~n7868;
  assign n7874 = ~n7872 & ~n7873;
  assign n7875 = n7836 & n7843;
  assign n7876 = ~n7836 & ~n7843;
  assign n7877 = ~n7875 & ~n7876;
  assign n7878 = ~n7846 & ~n7877;
  assign n7879 = ~n7871 & ~n7874;
  assign n7880 = ~n7864 & n7867;
  assign n7881 = n7864 & ~n7867;
  assign n7882 = ~n7880 & ~n7881;
  assign n7883 = ~n7839 & n7842;
  assign n7884 = n7839 & ~n7842;
  assign n7885 = ~n7883 & ~n7884;
  assign n7886 = ~n7882 & ~n7885;
  assign n7887 = ~n7878 & n7886;
  assign n7888 = ~n7879 & n7887;
  assign n7889 = n7874 & ~n7888;
  assign n7890 = ~n7874 & n7888;
  assign n7891 = ~n7889 & ~n7890;
  assign n7892 = n7877 & n7891;
  assign n7893 = ~n7889 & ~n7892;
  assign n7894 = n7871 & ~n7893;
  assign n7895 = ~n7846 & ~n7894;
  assign n7896 = ~n7871 & n7893;
  assign n7897 = ~n7895 & ~n7896;
  assign n7898 = pi754  & pi755 ;
  assign n7899 = ~pi754  & pi755 ;
  assign n7900 = pi754  & ~pi755 ;
  assign n7901 = ~n7899 & ~n7900;
  assign n7902 = pi756  & ~n7901;
  assign n7903 = ~n7898 & ~n7902;
  assign n7904 = pi751  & pi752 ;
  assign n7905 = ~pi751  & pi752 ;
  assign n7906 = pi751  & ~pi752 ;
  assign n7907 = ~n7905 & ~n7906;
  assign n7908 = pi753  & ~n7907;
  assign n7909 = ~n7904 & ~n7908;
  assign n7910 = ~n7903 & n7909;
  assign n7911 = n7903 & ~n7909;
  assign n7912 = ~n7910 & ~n7911;
  assign n7913 = ~pi753  & ~n7907;
  assign n7914 = pi753  & n7907;
  assign n7915 = ~n7913 & ~n7914;
  assign n7916 = ~pi756  & ~n7901;
  assign n7917 = pi756  & n7901;
  assign n7918 = ~n7916 & ~n7917;
  assign n7919 = ~n7915 & ~n7918;
  assign n7920 = ~n7912 & n7919;
  assign n7921 = ~n7903 & ~n7909;
  assign n7922 = ~n7920 & ~n7921;
  assign n7923 = pi760  & pi761 ;
  assign n7924 = ~pi760  & pi761 ;
  assign n7925 = pi760  & ~pi761 ;
  assign n7926 = ~n7924 & ~n7925;
  assign n7927 = pi762  & ~n7926;
  assign n7928 = ~n7923 & ~n7927;
  assign n7929 = pi757  & pi758 ;
  assign n7930 = ~pi757  & pi758 ;
  assign n7931 = pi757  & ~pi758 ;
  assign n7932 = ~n7930 & ~n7931;
  assign n7933 = pi759  & ~n7932;
  assign n7934 = ~n7929 & ~n7933;
  assign n7935 = ~n7928 & n7934;
  assign n7936 = n7928 & ~n7934;
  assign n7937 = ~n7935 & ~n7936;
  assign n7938 = ~pi759  & ~n7932;
  assign n7939 = pi759  & n7932;
  assign n7940 = ~n7938 & ~n7939;
  assign n7941 = ~pi762  & ~n7926;
  assign n7942 = pi762  & n7926;
  assign n7943 = ~n7941 & ~n7942;
  assign n7944 = ~n7940 & ~n7943;
  assign n7945 = ~n7937 & n7944;
  assign n7946 = ~n7928 & ~n7934;
  assign n7947 = ~n7945 & ~n7946;
  assign n7948 = n7937 & n7944;
  assign n7949 = ~n7937 & ~n7944;
  assign n7950 = ~n7948 & ~n7949;
  assign n7951 = n7912 & n7919;
  assign n7952 = ~n7912 & ~n7919;
  assign n7953 = ~n7951 & ~n7952;
  assign n7954 = ~n7922 & ~n7953;
  assign n7955 = ~n7947 & ~n7950;
  assign n7956 = ~n7940 & n7943;
  assign n7957 = n7940 & ~n7943;
  assign n7958 = ~n7956 & ~n7957;
  assign n7959 = ~n7915 & n7918;
  assign n7960 = n7915 & ~n7918;
  assign n7961 = ~n7959 & ~n7960;
  assign n7962 = ~n7958 & ~n7961;
  assign n7963 = ~n7954 & n7962;
  assign n7964 = ~n7955 & n7963;
  assign n7965 = n7950 & ~n7964;
  assign n7966 = ~n7950 & n7964;
  assign n7967 = ~n7965 & ~n7966;
  assign n7968 = n7953 & n7967;
  assign n7969 = ~n7965 & ~n7968;
  assign n7970 = n7947 & ~n7969;
  assign n7971 = ~n7922 & ~n7970;
  assign n7972 = ~n7947 & n7969;
  assign n7973 = ~n7971 & ~n7972;
  assign n7974 = n7897 & n7973;
  assign n7975 = ~n7922 & n7947;
  assign n7976 = n7922 & ~n7947;
  assign n7977 = ~n7975 & ~n7976;
  assign n7978 = n7969 & ~n7977;
  assign n7979 = ~n7969 & n7977;
  assign n7980 = ~n7978 & ~n7979;
  assign n7981 = ~n7846 & n7871;
  assign n7982 = n7846 & ~n7871;
  assign n7983 = ~n7981 & ~n7982;
  assign n7984 = n7893 & ~n7983;
  assign n7985 = ~n7893 & n7983;
  assign n7986 = ~n7984 & ~n7985;
  assign n7987 = n7980 & n7986;
  assign n7988 = n7882 & ~n7885;
  assign n7989 = ~n7882 & n7885;
  assign n7990 = ~n7988 & ~n7989;
  assign n7991 = n7958 & ~n7961;
  assign n7992 = ~n7958 & n7961;
  assign n7993 = ~n7991 & ~n7992;
  assign n7994 = ~n7990 & ~n7993;
  assign n7995 = ~n7877 & ~n7891;
  assign n7996 = ~n7892 & ~n7995;
  assign n7997 = ~n7994 & n7996;
  assign n7998 = ~n7953 & ~n7967;
  assign n7999 = ~n7968 & ~n7998;
  assign n8000 = n7994 & ~n7996;
  assign n8001 = ~n7997 & ~n8000;
  assign n8002 = n7999 & n8001;
  assign n8003 = ~n7997 & ~n8002;
  assign n8004 = ~n7980 & ~n7986;
  assign n8005 = ~n7987 & ~n8004;
  assign n8006 = n8003 & n8005;
  assign n8007 = ~n7987 & ~n8006;
  assign n8008 = ~n7974 & ~n8007;
  assign n8009 = ~n7897 & ~n7973;
  assign n8010 = ~n8008 & ~n8009;
  assign n8011 = ~n7821 & ~n8010;
  assign n8012 = n7821 & n8010;
  assign n8013 = ~n8011 & ~n8012;
  assign n8014 = ~n7784 & ~n7820;
  assign n8015 = ~n7818 & n8014;
  assign n8016 = n7818 & ~n8014;
  assign n8017 = ~n8015 & ~n8016;
  assign n8018 = ~n7974 & ~n8009;
  assign n8019 = ~n8007 & n8018;
  assign n8020 = n8007 & ~n8018;
  assign n8021 = ~n8019 & ~n8020;
  assign n8022 = n8017 & n8021;
  assign n8023 = ~n8003 & ~n8005;
  assign n8024 = ~n8006 & ~n8023;
  assign n8025 = ~n7814 & ~n7816;
  assign n8026 = ~n7817 & ~n8025;
  assign n8027 = n8024 & n8026;
  assign n8028 = ~n8024 & ~n8026;
  assign n8029 = ~n8027 & ~n8028;
  assign n8030 = ~n7800 & n7803;
  assign n8031 = n7800 & ~n7803;
  assign n8032 = ~n8030 & ~n8031;
  assign n8033 = ~n7990 & n7993;
  assign n8034 = n7990 & ~n7993;
  assign n8035 = ~n8033 & ~n8034;
  assign n8036 = ~n8032 & ~n8035;
  assign n8037 = ~n7809 & n7812;
  assign n8038 = ~n7813 & ~n8037;
  assign n8039 = ~n8036 & n8038;
  assign n8040 = ~n7999 & ~n8001;
  assign n8041 = ~n8002 & ~n8040;
  assign n8042 = n8036 & ~n8038;
  assign n8043 = ~n8039 & ~n8042;
  assign n8044 = n8041 & n8043;
  assign n8045 = ~n8039 & ~n8044;
  assign n8046 = n8029 & n8045;
  assign n8047 = ~n8027 & ~n8046;
  assign n8048 = ~n8017 & ~n8021;
  assign n8049 = ~n8022 & ~n8048;
  assign n8050 = ~n8047 & n8049;
  assign n8051 = ~n8022 & ~n8050;
  assign n8052 = n8013 & ~n8051;
  assign n8053 = ~n8011 & ~n8052;
  assign n8054 = ~n7631 & ~n8053;
  assign n8055 = ~n8013 & n8051;
  assign n8056 = ~n8052 & ~n8055;
  assign n8057 = ~n7591 & n7629;
  assign n8058 = ~n7630 & ~n8057;
  assign n8059 = n8056 & n8058;
  assign n8060 = n7625 & ~n7627;
  assign n8061 = ~n7628 & ~n8060;
  assign n8062 = n8047 & ~n8049;
  assign n8063 = ~n8050 & ~n8062;
  assign n8064 = n8061 & n8063;
  assign n8065 = ~n8061 & ~n8063;
  assign n8066 = ~n8064 & ~n8065;
  assign n8067 = ~n8029 & ~n8045;
  assign n8068 = ~n8046 & ~n8067;
  assign n8069 = ~n7607 & ~n7623;
  assign n8070 = ~n7624 & ~n8069;
  assign n8071 = n8068 & n8070;
  assign n8072 = ~n8068 & ~n8070;
  assign n8073 = ~n8071 & ~n8072;
  assign n8074 = ~n7610 & n7613;
  assign n8075 = n7610 & ~n7613;
  assign n8076 = ~n8074 & ~n8075;
  assign n8077 = ~n8032 & n8035;
  assign n8078 = n8032 & ~n8035;
  assign n8079 = ~n8077 & ~n8078;
  assign n8080 = ~n8076 & ~n8079;
  assign n8081 = ~n7619 & ~n7621;
  assign n8082 = ~n7622 & ~n8081;
  assign n8083 = ~n8080 & n8082;
  assign n8084 = ~n8041 & ~n8043;
  assign n8085 = ~n8044 & ~n8084;
  assign n8086 = n8080 & ~n8082;
  assign n8087 = ~n8083 & ~n8086;
  assign n8088 = n8085 & n8087;
  assign n8089 = ~n8083 & ~n8088;
  assign n8090 = n8073 & n8089;
  assign n8091 = ~n8071 & ~n8090;
  assign n8092 = n8066 & ~n8091;
  assign n8093 = ~n8064 & ~n8092;
  assign n8094 = ~n8056 & ~n8058;
  assign n8095 = ~n8059 & ~n8094;
  assign n8096 = ~n8093 & n8095;
  assign n8097 = ~n8059 & ~n8096;
  assign n8098 = n7631 & n8053;
  assign n8099 = ~n8054 & ~n8098;
  assign n8100 = ~n8097 & n8099;
  assign n8101 = ~n8054 & ~n8100;
  assign n8102 = pi739  & ~pi740 ;
  assign n8103 = ~pi739  & pi740 ;
  assign n8104 = ~n8102 & ~n8103;
  assign n8105 = ~pi741  & ~n8104;
  assign n8106 = pi741  & n8104;
  assign n8107 = ~n8105 & ~n8106;
  assign n8108 = pi742  & ~pi743 ;
  assign n8109 = ~pi742  & pi743 ;
  assign n8110 = ~n8108 & ~n8109;
  assign n8111 = ~pi744  & ~n8110;
  assign n8112 = pi744  & n8110;
  assign n8113 = ~n8111 & ~n8112;
  assign n8114 = ~n8107 & ~n8113;
  assign n8115 = pi742  & pi743 ;
  assign n8116 = pi744  & ~n8110;
  assign n8117 = ~n8115 & ~n8116;
  assign n8118 = pi739  & pi740 ;
  assign n8119 = pi741  & ~n8104;
  assign n8120 = ~n8118 & ~n8119;
  assign n8121 = n8117 & ~n8120;
  assign n8122 = ~n8117 & n8120;
  assign n8123 = ~n8121 & ~n8122;
  assign n8124 = n8114 & ~n8123;
  assign n8125 = ~n8117 & ~n8120;
  assign n8126 = ~n8124 & ~n8125;
  assign n8127 = pi748  & pi749 ;
  assign n8128 = pi748  & ~pi749 ;
  assign n8129 = ~pi748  & pi749 ;
  assign n8130 = ~n8128 & ~n8129;
  assign n8131 = pi750  & ~n8130;
  assign n8132 = ~n8127 & ~n8131;
  assign n8133 = pi745  & pi746 ;
  assign n8134 = pi745  & ~pi746 ;
  assign n8135 = ~pi745  & pi746 ;
  assign n8136 = ~n8134 & ~n8135;
  assign n8137 = pi747  & ~n8136;
  assign n8138 = ~n8133 & ~n8137;
  assign n8139 = ~n8132 & n8138;
  assign n8140 = n8132 & ~n8138;
  assign n8141 = ~n8139 & ~n8140;
  assign n8142 = ~pi747  & ~n8136;
  assign n8143 = pi747  & n8136;
  assign n8144 = ~n8142 & ~n8143;
  assign n8145 = ~pi750  & ~n8130;
  assign n8146 = pi750  & n8130;
  assign n8147 = ~n8145 & ~n8146;
  assign n8148 = ~n8144 & ~n8147;
  assign n8149 = ~n8141 & n8148;
  assign n8150 = ~n8132 & ~n8138;
  assign n8151 = ~n8149 & ~n8150;
  assign n8152 = n8141 & n8148;
  assign n8153 = ~n8141 & ~n8148;
  assign n8154 = ~n8152 & ~n8153;
  assign n8155 = ~n8151 & ~n8154;
  assign n8156 = n8114 & n8123;
  assign n8157 = ~n8114 & ~n8123;
  assign n8158 = ~n8156 & ~n8157;
  assign n8159 = ~n8126 & ~n8158;
  assign n8160 = ~n8107 & n8113;
  assign n8161 = n8107 & ~n8113;
  assign n8162 = ~n8160 & ~n8161;
  assign n8163 = ~n8144 & n8147;
  assign n8164 = n8144 & ~n8147;
  assign n8165 = ~n8163 & ~n8164;
  assign n8166 = ~n8162 & ~n8165;
  assign n8167 = ~n8155 & n8166;
  assign n8168 = ~n8159 & n8167;
  assign n8169 = n8154 & ~n8168;
  assign n8170 = ~n8154 & n8168;
  assign n8171 = ~n8169 & ~n8170;
  assign n8172 = n8158 & n8171;
  assign n8173 = ~n8169 & ~n8172;
  assign n8174 = n8151 & ~n8173;
  assign n8175 = ~n8126 & ~n8174;
  assign n8176 = ~n8151 & n8173;
  assign n8177 = ~n8175 & ~n8176;
  assign n8178 = pi727  & ~pi728 ;
  assign n8179 = ~pi727  & pi728 ;
  assign n8180 = ~n8178 & ~n8179;
  assign n8181 = ~pi729  & ~n8180;
  assign n8182 = pi729  & n8180;
  assign n8183 = ~n8181 & ~n8182;
  assign n8184 = pi730  & ~pi731 ;
  assign n8185 = ~pi730  & pi731 ;
  assign n8186 = ~n8184 & ~n8185;
  assign n8187 = ~pi732  & ~n8186;
  assign n8188 = pi732  & n8186;
  assign n8189 = ~n8187 & ~n8188;
  assign n8190 = ~n8183 & ~n8189;
  assign n8191 = pi730  & pi731 ;
  assign n8192 = pi732  & ~n8186;
  assign n8193 = ~n8191 & ~n8192;
  assign n8194 = pi727  & pi728 ;
  assign n8195 = pi729  & ~n8180;
  assign n8196 = ~n8194 & ~n8195;
  assign n8197 = n8193 & ~n8196;
  assign n8198 = ~n8193 & n8196;
  assign n8199 = ~n8197 & ~n8198;
  assign n8200 = n8190 & ~n8199;
  assign n8201 = ~n8193 & ~n8196;
  assign n8202 = ~n8200 & ~n8201;
  assign n8203 = pi736  & pi737 ;
  assign n8204 = pi736  & ~pi737 ;
  assign n8205 = ~pi736  & pi737 ;
  assign n8206 = ~n8204 & ~n8205;
  assign n8207 = pi738  & ~n8206;
  assign n8208 = ~n8203 & ~n8207;
  assign n8209 = pi733  & pi734 ;
  assign n8210 = pi733  & ~pi734 ;
  assign n8211 = ~pi733  & pi734 ;
  assign n8212 = ~n8210 & ~n8211;
  assign n8213 = pi735  & ~n8212;
  assign n8214 = ~n8209 & ~n8213;
  assign n8215 = ~n8208 & n8214;
  assign n8216 = n8208 & ~n8214;
  assign n8217 = ~n8215 & ~n8216;
  assign n8218 = ~pi735  & ~n8212;
  assign n8219 = pi735  & n8212;
  assign n8220 = ~n8218 & ~n8219;
  assign n8221 = ~pi738  & ~n8206;
  assign n8222 = pi738  & n8206;
  assign n8223 = ~n8221 & ~n8222;
  assign n8224 = ~n8220 & ~n8223;
  assign n8225 = ~n8217 & n8224;
  assign n8226 = ~n8208 & ~n8214;
  assign n8227 = ~n8225 & ~n8226;
  assign n8228 = n8217 & n8224;
  assign n8229 = ~n8217 & ~n8224;
  assign n8230 = ~n8228 & ~n8229;
  assign n8231 = ~n8227 & ~n8230;
  assign n8232 = n8190 & n8199;
  assign n8233 = ~n8190 & ~n8199;
  assign n8234 = ~n8232 & ~n8233;
  assign n8235 = ~n8202 & ~n8234;
  assign n8236 = ~n8183 & n8189;
  assign n8237 = n8183 & ~n8189;
  assign n8238 = ~n8236 & ~n8237;
  assign n8239 = ~n8220 & n8223;
  assign n8240 = n8220 & ~n8223;
  assign n8241 = ~n8239 & ~n8240;
  assign n8242 = ~n8238 & ~n8241;
  assign n8243 = ~n8231 & n8242;
  assign n8244 = ~n8235 & n8243;
  assign n8245 = n8230 & ~n8244;
  assign n8246 = ~n8230 & n8244;
  assign n8247 = ~n8245 & ~n8246;
  assign n8248 = n8234 & n8247;
  assign n8249 = ~n8245 & ~n8248;
  assign n8250 = n8227 & ~n8249;
  assign n8251 = ~n8202 & ~n8250;
  assign n8252 = ~n8227 & n8249;
  assign n8253 = ~n8251 & ~n8252;
  assign n8254 = n8177 & n8253;
  assign n8255 = ~n8202 & n8227;
  assign n8256 = n8202 & ~n8227;
  assign n8257 = ~n8255 & ~n8256;
  assign n8258 = n8249 & ~n8257;
  assign n8259 = ~n8249 & n8257;
  assign n8260 = ~n8258 & ~n8259;
  assign n8261 = ~n8126 & n8151;
  assign n8262 = n8126 & ~n8151;
  assign n8263 = ~n8261 & ~n8262;
  assign n8264 = n8173 & ~n8263;
  assign n8265 = ~n8173 & n8263;
  assign n8266 = ~n8264 & ~n8265;
  assign n8267 = n8260 & n8266;
  assign n8268 = ~n8162 & n8165;
  assign n8269 = n8162 & ~n8165;
  assign n8270 = ~n8268 & ~n8269;
  assign n8271 = ~n8238 & n8241;
  assign n8272 = n8238 & ~n8241;
  assign n8273 = ~n8271 & ~n8272;
  assign n8274 = ~n8270 & ~n8273;
  assign n8275 = ~n8158 & ~n8171;
  assign n8276 = ~n8172 & ~n8275;
  assign n8277 = ~n8274 & n8276;
  assign n8278 = ~n8234 & ~n8247;
  assign n8279 = ~n8248 & ~n8278;
  assign n8280 = ~n8274 & ~n8276;
  assign n8281 = n8276 & ~n8277;
  assign n8282 = ~n8280 & ~n8281;
  assign n8283 = n8279 & ~n8282;
  assign n8284 = ~n8277 & ~n8283;
  assign n8285 = ~n8260 & ~n8266;
  assign n8286 = ~n8267 & ~n8285;
  assign n8287 = n8284 & n8286;
  assign n8288 = ~n8267 & ~n8287;
  assign n8289 = ~n8254 & ~n8288;
  assign n8290 = ~n8177 & ~n8253;
  assign n8291 = ~n8289 & ~n8290;
  assign n8292 = pi715  & ~pi716 ;
  assign n8293 = ~pi715  & pi716 ;
  assign n8294 = ~n8292 & ~n8293;
  assign n8295 = ~pi717  & ~n8294;
  assign n8296 = pi717  & n8294;
  assign n8297 = ~n8295 & ~n8296;
  assign n8298 = pi718  & ~pi719 ;
  assign n8299 = ~pi718  & pi719 ;
  assign n8300 = ~n8298 & ~n8299;
  assign n8301 = ~pi720  & ~n8300;
  assign n8302 = pi720  & n8300;
  assign n8303 = ~n8301 & ~n8302;
  assign n8304 = ~n8297 & ~n8303;
  assign n8305 = pi718  & pi719 ;
  assign n8306 = pi720  & ~n8300;
  assign n8307 = ~n8305 & ~n8306;
  assign n8308 = pi715  & pi716 ;
  assign n8309 = pi717  & ~n8294;
  assign n8310 = ~n8308 & ~n8309;
  assign n8311 = n8307 & ~n8310;
  assign n8312 = ~n8307 & n8310;
  assign n8313 = ~n8311 & ~n8312;
  assign n8314 = n8304 & ~n8313;
  assign n8315 = ~n8307 & ~n8310;
  assign n8316 = ~n8314 & ~n8315;
  assign n8317 = pi724  & pi725 ;
  assign n8318 = pi724  & ~pi725 ;
  assign n8319 = ~pi724  & pi725 ;
  assign n8320 = ~n8318 & ~n8319;
  assign n8321 = pi726  & ~n8320;
  assign n8322 = ~n8317 & ~n8321;
  assign n8323 = pi721  & pi722 ;
  assign n8324 = pi721  & ~pi722 ;
  assign n8325 = ~pi721  & pi722 ;
  assign n8326 = ~n8324 & ~n8325;
  assign n8327 = pi723  & ~n8326;
  assign n8328 = ~n8323 & ~n8327;
  assign n8329 = ~n8322 & n8328;
  assign n8330 = n8322 & ~n8328;
  assign n8331 = ~n8329 & ~n8330;
  assign n8332 = ~pi723  & ~n8326;
  assign n8333 = pi723  & n8326;
  assign n8334 = ~n8332 & ~n8333;
  assign n8335 = ~pi726  & ~n8320;
  assign n8336 = pi726  & n8320;
  assign n8337 = ~n8335 & ~n8336;
  assign n8338 = ~n8334 & ~n8337;
  assign n8339 = ~n8331 & n8338;
  assign n8340 = ~n8322 & ~n8328;
  assign n8341 = ~n8339 & ~n8340;
  assign n8342 = n8331 & n8338;
  assign n8343 = ~n8331 & ~n8338;
  assign n8344 = ~n8342 & ~n8343;
  assign n8345 = ~n8341 & ~n8344;
  assign n8346 = n8304 & n8313;
  assign n8347 = ~n8304 & ~n8313;
  assign n8348 = ~n8346 & ~n8347;
  assign n8349 = ~n8316 & ~n8348;
  assign n8350 = ~n8297 & n8303;
  assign n8351 = n8297 & ~n8303;
  assign n8352 = ~n8350 & ~n8351;
  assign n8353 = ~n8334 & n8337;
  assign n8354 = n8334 & ~n8337;
  assign n8355 = ~n8353 & ~n8354;
  assign n8356 = ~n8352 & ~n8355;
  assign n8357 = ~n8345 & n8356;
  assign n8358 = ~n8349 & n8357;
  assign n8359 = n8344 & ~n8358;
  assign n8360 = ~n8344 & n8358;
  assign n8361 = ~n8359 & ~n8360;
  assign n8362 = n8348 & n8361;
  assign n8363 = ~n8359 & ~n8362;
  assign n8364 = n8341 & ~n8363;
  assign n8365 = ~n8316 & ~n8364;
  assign n8366 = ~n8341 & n8363;
  assign n8367 = ~n8365 & ~n8366;
  assign n8368 = pi706  & pi707 ;
  assign n8369 = ~pi706  & pi707 ;
  assign n8370 = pi706  & ~pi707 ;
  assign n8371 = ~n8369 & ~n8370;
  assign n8372 = pi708  & ~n8371;
  assign n8373 = ~n8368 & ~n8372;
  assign n8374 = pi703  & pi704 ;
  assign n8375 = ~pi703  & pi704 ;
  assign n8376 = pi703  & ~pi704 ;
  assign n8377 = ~n8375 & ~n8376;
  assign n8378 = pi705  & ~n8377;
  assign n8379 = ~n8374 & ~n8378;
  assign n8380 = ~n8373 & n8379;
  assign n8381 = n8373 & ~n8379;
  assign n8382 = ~n8380 & ~n8381;
  assign n8383 = ~pi705  & ~n8377;
  assign n8384 = pi705  & n8377;
  assign n8385 = ~n8383 & ~n8384;
  assign n8386 = ~pi708  & ~n8371;
  assign n8387 = pi708  & n8371;
  assign n8388 = ~n8386 & ~n8387;
  assign n8389 = ~n8385 & ~n8388;
  assign n8390 = ~n8382 & n8389;
  assign n8391 = ~n8373 & ~n8379;
  assign n8392 = ~n8390 & ~n8391;
  assign n8393 = pi712  & pi713 ;
  assign n8394 = ~pi712  & pi713 ;
  assign n8395 = pi712  & ~pi713 ;
  assign n8396 = ~n8394 & ~n8395;
  assign n8397 = pi714  & ~n8396;
  assign n8398 = ~n8393 & ~n8397;
  assign n8399 = pi709  & pi710 ;
  assign n8400 = ~pi709  & pi710 ;
  assign n8401 = pi709  & ~pi710 ;
  assign n8402 = ~n8400 & ~n8401;
  assign n8403 = pi711  & ~n8402;
  assign n8404 = ~n8399 & ~n8403;
  assign n8405 = ~n8398 & n8404;
  assign n8406 = n8398 & ~n8404;
  assign n8407 = ~n8405 & ~n8406;
  assign n8408 = ~pi711  & ~n8402;
  assign n8409 = pi711  & n8402;
  assign n8410 = ~n8408 & ~n8409;
  assign n8411 = ~pi714  & ~n8396;
  assign n8412 = pi714  & n8396;
  assign n8413 = ~n8411 & ~n8412;
  assign n8414 = ~n8410 & ~n8413;
  assign n8415 = ~n8407 & n8414;
  assign n8416 = ~n8398 & ~n8404;
  assign n8417 = ~n8415 & ~n8416;
  assign n8418 = n8407 & n8414;
  assign n8419 = ~n8407 & ~n8414;
  assign n8420 = ~n8418 & ~n8419;
  assign n8421 = n8382 & n8389;
  assign n8422 = ~n8382 & ~n8389;
  assign n8423 = ~n8421 & ~n8422;
  assign n8424 = ~n8392 & ~n8423;
  assign n8425 = ~n8417 & ~n8420;
  assign n8426 = ~n8410 & n8413;
  assign n8427 = n8410 & ~n8413;
  assign n8428 = ~n8426 & ~n8427;
  assign n8429 = ~n8385 & n8388;
  assign n8430 = n8385 & ~n8388;
  assign n8431 = ~n8429 & ~n8430;
  assign n8432 = ~n8428 & ~n8431;
  assign n8433 = ~n8424 & n8432;
  assign n8434 = ~n8425 & n8433;
  assign n8435 = n8420 & ~n8434;
  assign n8436 = ~n8420 & n8434;
  assign n8437 = ~n8435 & ~n8436;
  assign n8438 = n8423 & n8437;
  assign n8439 = ~n8435 & ~n8438;
  assign n8440 = n8417 & ~n8439;
  assign n8441 = ~n8392 & ~n8440;
  assign n8442 = ~n8417 & n8439;
  assign n8443 = ~n8441 & ~n8442;
  assign n8444 = n8367 & n8443;
  assign n8445 = ~n8392 & n8417;
  assign n8446 = n8392 & ~n8417;
  assign n8447 = ~n8445 & ~n8446;
  assign n8448 = n8439 & ~n8447;
  assign n8449 = ~n8439 & n8447;
  assign n8450 = ~n8448 & ~n8449;
  assign n8451 = ~n8316 & n8341;
  assign n8452 = n8316 & ~n8341;
  assign n8453 = ~n8451 & ~n8452;
  assign n8454 = n8363 & ~n8453;
  assign n8455 = ~n8363 & n8453;
  assign n8456 = ~n8454 & ~n8455;
  assign n8457 = n8450 & n8456;
  assign n8458 = ~n8352 & n8355;
  assign n8459 = n8352 & ~n8355;
  assign n8460 = ~n8458 & ~n8459;
  assign n8461 = n8428 & ~n8431;
  assign n8462 = ~n8428 & n8431;
  assign n8463 = ~n8461 & ~n8462;
  assign n8464 = ~n8460 & ~n8463;
  assign n8465 = ~n8348 & ~n8361;
  assign n8466 = ~n8362 & ~n8465;
  assign n8467 = ~n8464 & n8466;
  assign n8468 = ~n8423 & ~n8437;
  assign n8469 = ~n8438 & ~n8468;
  assign n8470 = n8464 & ~n8466;
  assign n8471 = ~n8467 & ~n8470;
  assign n8472 = n8469 & n8471;
  assign n8473 = ~n8467 & ~n8472;
  assign n8474 = ~n8450 & ~n8456;
  assign n8475 = ~n8457 & ~n8474;
  assign n8476 = n8473 & n8475;
  assign n8477 = ~n8457 & ~n8476;
  assign n8478 = ~n8444 & ~n8477;
  assign n8479 = ~n8367 & ~n8443;
  assign n8480 = ~n8478 & ~n8479;
  assign n8481 = ~n8291 & ~n8480;
  assign n8482 = n8291 & n8480;
  assign n8483 = ~n8481 & ~n8482;
  assign n8484 = ~n8254 & ~n8290;
  assign n8485 = ~n8288 & n8484;
  assign n8486 = n8288 & ~n8484;
  assign n8487 = ~n8485 & ~n8486;
  assign n8488 = ~n8444 & ~n8479;
  assign n8489 = ~n8477 & n8488;
  assign n8490 = n8477 & ~n8488;
  assign n8491 = ~n8489 & ~n8490;
  assign n8492 = n8487 & n8491;
  assign n8493 = ~n8473 & ~n8475;
  assign n8494 = ~n8476 & ~n8493;
  assign n8495 = ~n8284 & ~n8286;
  assign n8496 = ~n8287 & ~n8495;
  assign n8497 = n8494 & n8496;
  assign n8498 = ~n8494 & ~n8496;
  assign n8499 = ~n8497 & ~n8498;
  assign n8500 = ~n8270 & n8273;
  assign n8501 = n8270 & ~n8273;
  assign n8502 = ~n8500 & ~n8501;
  assign n8503 = ~n8460 & n8463;
  assign n8504 = n8460 & ~n8463;
  assign n8505 = ~n8503 & ~n8504;
  assign n8506 = ~n8502 & ~n8505;
  assign n8507 = ~n8279 & n8282;
  assign n8508 = ~n8283 & ~n8507;
  assign n8509 = ~n8506 & n8508;
  assign n8510 = ~n8469 & ~n8471;
  assign n8511 = ~n8472 & ~n8510;
  assign n8512 = n8506 & ~n8508;
  assign n8513 = ~n8509 & ~n8512;
  assign n8514 = n8511 & n8513;
  assign n8515 = ~n8509 & ~n8514;
  assign n8516 = n8499 & n8515;
  assign n8517 = ~n8497 & ~n8516;
  assign n8518 = ~n8487 & ~n8491;
  assign n8519 = ~n8492 & ~n8518;
  assign n8520 = ~n8517 & n8519;
  assign n8521 = ~n8492 & ~n8520;
  assign n8522 = n8483 & ~n8521;
  assign n8523 = ~n8481 & ~n8522;
  assign n8524 = pi694  & pi695 ;
  assign n8525 = ~pi694  & pi695 ;
  assign n8526 = pi694  & ~pi695 ;
  assign n8527 = ~n8525 & ~n8526;
  assign n8528 = pi696  & ~n8527;
  assign n8529 = ~n8524 & ~n8528;
  assign n8530 = pi691  & pi692 ;
  assign n8531 = ~pi691  & pi692 ;
  assign n8532 = pi691  & ~pi692 ;
  assign n8533 = ~n8531 & ~n8532;
  assign n8534 = pi693  & ~n8533;
  assign n8535 = ~n8530 & ~n8534;
  assign n8536 = ~n8529 & n8535;
  assign n8537 = n8529 & ~n8535;
  assign n8538 = ~n8536 & ~n8537;
  assign n8539 = ~pi693  & ~n8533;
  assign n8540 = pi693  & n8533;
  assign n8541 = ~n8539 & ~n8540;
  assign n8542 = ~pi696  & ~n8527;
  assign n8543 = pi696  & n8527;
  assign n8544 = ~n8542 & ~n8543;
  assign n8545 = ~n8541 & ~n8544;
  assign n8546 = ~n8538 & n8545;
  assign n8547 = ~n8529 & ~n8535;
  assign n8548 = ~n8546 & ~n8547;
  assign n8549 = pi700  & pi701 ;
  assign n8550 = ~pi700  & pi701 ;
  assign n8551 = pi700  & ~pi701 ;
  assign n8552 = ~n8550 & ~n8551;
  assign n8553 = pi702  & ~n8552;
  assign n8554 = ~n8549 & ~n8553;
  assign n8555 = pi697  & pi698 ;
  assign n8556 = ~pi697  & pi698 ;
  assign n8557 = pi697  & ~pi698 ;
  assign n8558 = ~n8556 & ~n8557;
  assign n8559 = pi699  & ~n8558;
  assign n8560 = ~n8555 & ~n8559;
  assign n8561 = ~n8554 & n8560;
  assign n8562 = n8554 & ~n8560;
  assign n8563 = ~n8561 & ~n8562;
  assign n8564 = ~pi699  & ~n8558;
  assign n8565 = pi699  & n8558;
  assign n8566 = ~n8564 & ~n8565;
  assign n8567 = ~pi702  & ~n8552;
  assign n8568 = pi702  & n8552;
  assign n8569 = ~n8567 & ~n8568;
  assign n8570 = ~n8566 & ~n8569;
  assign n8571 = ~n8563 & n8570;
  assign n8572 = ~n8554 & ~n8560;
  assign n8573 = ~n8571 & ~n8572;
  assign n8574 = n8563 & n8570;
  assign n8575 = ~n8563 & ~n8570;
  assign n8576 = ~n8574 & ~n8575;
  assign n8577 = n8538 & n8545;
  assign n8578 = ~n8538 & ~n8545;
  assign n8579 = ~n8577 & ~n8578;
  assign n8580 = ~n8548 & ~n8579;
  assign n8581 = ~n8573 & ~n8576;
  assign n8582 = ~n8566 & n8569;
  assign n8583 = n8566 & ~n8569;
  assign n8584 = ~n8582 & ~n8583;
  assign n8585 = ~n8541 & n8544;
  assign n8586 = n8541 & ~n8544;
  assign n8587 = ~n8585 & ~n8586;
  assign n8588 = ~n8584 & ~n8587;
  assign n8589 = ~n8580 & n8588;
  assign n8590 = ~n8581 & n8589;
  assign n8591 = n8576 & ~n8590;
  assign n8592 = ~n8576 & n8590;
  assign n8593 = ~n8591 & ~n8592;
  assign n8594 = n8579 & n8593;
  assign n8595 = ~n8591 & ~n8594;
  assign n8596 = n8573 & ~n8595;
  assign n8597 = ~n8548 & ~n8596;
  assign n8598 = ~n8573 & n8595;
  assign n8599 = ~n8597 & ~n8598;
  assign n8600 = pi682  & pi683 ;
  assign n8601 = ~pi682  & pi683 ;
  assign n8602 = pi682  & ~pi683 ;
  assign n8603 = ~n8601 & ~n8602;
  assign n8604 = pi684  & ~n8603;
  assign n8605 = ~n8600 & ~n8604;
  assign n8606 = pi679  & pi680 ;
  assign n8607 = ~pi679  & pi680 ;
  assign n8608 = pi679  & ~pi680 ;
  assign n8609 = ~n8607 & ~n8608;
  assign n8610 = pi681  & ~n8609;
  assign n8611 = ~n8606 & ~n8610;
  assign n8612 = ~n8605 & n8611;
  assign n8613 = n8605 & ~n8611;
  assign n8614 = ~n8612 & ~n8613;
  assign n8615 = ~pi681  & ~n8609;
  assign n8616 = pi681  & n8609;
  assign n8617 = ~n8615 & ~n8616;
  assign n8618 = ~pi684  & ~n8603;
  assign n8619 = pi684  & n8603;
  assign n8620 = ~n8618 & ~n8619;
  assign n8621 = ~n8617 & ~n8620;
  assign n8622 = ~n8614 & n8621;
  assign n8623 = ~n8605 & ~n8611;
  assign n8624 = ~n8622 & ~n8623;
  assign n8625 = pi688  & pi689 ;
  assign n8626 = ~pi688  & pi689 ;
  assign n8627 = pi688  & ~pi689 ;
  assign n8628 = ~n8626 & ~n8627;
  assign n8629 = pi690  & ~n8628;
  assign n8630 = ~n8625 & ~n8629;
  assign n8631 = pi685  & pi686 ;
  assign n8632 = ~pi685  & pi686 ;
  assign n8633 = pi685  & ~pi686 ;
  assign n8634 = ~n8632 & ~n8633;
  assign n8635 = pi687  & ~n8634;
  assign n8636 = ~n8631 & ~n8635;
  assign n8637 = ~n8630 & n8636;
  assign n8638 = n8630 & ~n8636;
  assign n8639 = ~n8637 & ~n8638;
  assign n8640 = ~pi687  & ~n8634;
  assign n8641 = pi687  & n8634;
  assign n8642 = ~n8640 & ~n8641;
  assign n8643 = ~pi690  & ~n8628;
  assign n8644 = pi690  & n8628;
  assign n8645 = ~n8643 & ~n8644;
  assign n8646 = ~n8642 & ~n8645;
  assign n8647 = ~n8639 & n8646;
  assign n8648 = ~n8630 & ~n8636;
  assign n8649 = ~n8647 & ~n8648;
  assign n8650 = n8639 & n8646;
  assign n8651 = ~n8639 & ~n8646;
  assign n8652 = ~n8650 & ~n8651;
  assign n8653 = n8614 & n8621;
  assign n8654 = ~n8614 & ~n8621;
  assign n8655 = ~n8653 & ~n8654;
  assign n8656 = ~n8624 & ~n8655;
  assign n8657 = ~n8649 & ~n8652;
  assign n8658 = ~n8642 & n8645;
  assign n8659 = n8642 & ~n8645;
  assign n8660 = ~n8658 & ~n8659;
  assign n8661 = ~n8617 & n8620;
  assign n8662 = n8617 & ~n8620;
  assign n8663 = ~n8661 & ~n8662;
  assign n8664 = ~n8660 & ~n8663;
  assign n8665 = ~n8656 & n8664;
  assign n8666 = ~n8657 & n8665;
  assign n8667 = n8652 & ~n8666;
  assign n8668 = ~n8652 & n8666;
  assign n8669 = ~n8667 & ~n8668;
  assign n8670 = n8655 & n8669;
  assign n8671 = ~n8667 & ~n8670;
  assign n8672 = n8649 & ~n8671;
  assign n8673 = ~n8624 & ~n8672;
  assign n8674 = ~n8649 & n8671;
  assign n8675 = ~n8673 & ~n8674;
  assign n8676 = n8599 & n8675;
  assign n8677 = ~n8624 & n8649;
  assign n8678 = n8624 & ~n8649;
  assign n8679 = ~n8677 & ~n8678;
  assign n8680 = n8671 & ~n8679;
  assign n8681 = ~n8671 & n8679;
  assign n8682 = ~n8680 & ~n8681;
  assign n8683 = ~n8548 & n8573;
  assign n8684 = n8548 & ~n8573;
  assign n8685 = ~n8683 & ~n8684;
  assign n8686 = n8595 & ~n8685;
  assign n8687 = ~n8595 & n8685;
  assign n8688 = ~n8686 & ~n8687;
  assign n8689 = n8682 & n8688;
  assign n8690 = n8584 & ~n8587;
  assign n8691 = ~n8584 & n8587;
  assign n8692 = ~n8690 & ~n8691;
  assign n8693 = n8660 & ~n8663;
  assign n8694 = ~n8660 & n8663;
  assign n8695 = ~n8693 & ~n8694;
  assign n8696 = ~n8692 & ~n8695;
  assign n8697 = ~n8579 & ~n8593;
  assign n8698 = ~n8594 & ~n8697;
  assign n8699 = ~n8696 & n8698;
  assign n8700 = ~n8655 & ~n8669;
  assign n8701 = ~n8670 & ~n8700;
  assign n8702 = ~n8696 & ~n8698;
  assign n8703 = n8698 & ~n8699;
  assign n8704 = ~n8702 & ~n8703;
  assign n8705 = n8701 & ~n8704;
  assign n8706 = ~n8699 & ~n8705;
  assign n8707 = ~n8682 & ~n8688;
  assign n8708 = ~n8689 & ~n8707;
  assign n8709 = n8706 & n8708;
  assign n8710 = ~n8689 & ~n8709;
  assign n8711 = ~n8676 & ~n8710;
  assign n8712 = ~n8599 & ~n8675;
  assign n8713 = ~n8711 & ~n8712;
  assign n8714 = pi670  & pi671 ;
  assign n8715 = ~pi670  & pi671 ;
  assign n8716 = pi670  & ~pi671 ;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = pi672  & ~n8717;
  assign n8719 = ~n8714 & ~n8718;
  assign n8720 = pi667  & pi668 ;
  assign n8721 = ~pi667  & pi668 ;
  assign n8722 = pi667  & ~pi668 ;
  assign n8723 = ~n8721 & ~n8722;
  assign n8724 = pi669  & ~n8723;
  assign n8725 = ~n8720 & ~n8724;
  assign n8726 = ~n8719 & n8725;
  assign n8727 = n8719 & ~n8725;
  assign n8728 = ~n8726 & ~n8727;
  assign n8729 = ~pi669  & ~n8723;
  assign n8730 = pi669  & n8723;
  assign n8731 = ~n8729 & ~n8730;
  assign n8732 = ~pi672  & ~n8717;
  assign n8733 = pi672  & n8717;
  assign n8734 = ~n8732 & ~n8733;
  assign n8735 = ~n8731 & ~n8734;
  assign n8736 = ~n8728 & n8735;
  assign n8737 = ~n8719 & ~n8725;
  assign n8738 = ~n8736 & ~n8737;
  assign n8739 = pi676  & pi677 ;
  assign n8740 = ~pi676  & pi677 ;
  assign n8741 = pi676  & ~pi677 ;
  assign n8742 = ~n8740 & ~n8741;
  assign n8743 = pi678  & ~n8742;
  assign n8744 = ~n8739 & ~n8743;
  assign n8745 = pi673  & pi674 ;
  assign n8746 = ~pi673  & pi674 ;
  assign n8747 = pi673  & ~pi674 ;
  assign n8748 = ~n8746 & ~n8747;
  assign n8749 = pi675  & ~n8748;
  assign n8750 = ~n8745 & ~n8749;
  assign n8751 = ~n8744 & n8750;
  assign n8752 = n8744 & ~n8750;
  assign n8753 = ~n8751 & ~n8752;
  assign n8754 = ~pi675  & ~n8748;
  assign n8755 = pi675  & n8748;
  assign n8756 = ~n8754 & ~n8755;
  assign n8757 = ~pi678  & ~n8742;
  assign n8758 = pi678  & n8742;
  assign n8759 = ~n8757 & ~n8758;
  assign n8760 = ~n8756 & ~n8759;
  assign n8761 = ~n8753 & n8760;
  assign n8762 = ~n8744 & ~n8750;
  assign n8763 = ~n8761 & ~n8762;
  assign n8764 = n8753 & n8760;
  assign n8765 = ~n8753 & ~n8760;
  assign n8766 = ~n8764 & ~n8765;
  assign n8767 = n8728 & n8735;
  assign n8768 = ~n8728 & ~n8735;
  assign n8769 = ~n8767 & ~n8768;
  assign n8770 = ~n8738 & ~n8769;
  assign n8771 = ~n8763 & ~n8766;
  assign n8772 = ~n8756 & n8759;
  assign n8773 = n8756 & ~n8759;
  assign n8774 = ~n8772 & ~n8773;
  assign n8775 = ~n8731 & n8734;
  assign n8776 = n8731 & ~n8734;
  assign n8777 = ~n8775 & ~n8776;
  assign n8778 = ~n8774 & ~n8777;
  assign n8779 = ~n8770 & n8778;
  assign n8780 = ~n8771 & n8779;
  assign n8781 = n8766 & ~n8780;
  assign n8782 = ~n8766 & n8780;
  assign n8783 = ~n8781 & ~n8782;
  assign n8784 = n8769 & n8783;
  assign n8785 = ~n8781 & ~n8784;
  assign n8786 = n8763 & ~n8785;
  assign n8787 = ~n8738 & ~n8786;
  assign n8788 = ~n8763 & n8785;
  assign n8789 = ~n8787 & ~n8788;
  assign n8790 = pi658  & pi659 ;
  assign n8791 = ~pi658  & pi659 ;
  assign n8792 = pi658  & ~pi659 ;
  assign n8793 = ~n8791 & ~n8792;
  assign n8794 = pi660  & ~n8793;
  assign n8795 = ~n8790 & ~n8794;
  assign n8796 = pi655  & pi656 ;
  assign n8797 = ~pi655  & pi656 ;
  assign n8798 = pi655  & ~pi656 ;
  assign n8799 = ~n8797 & ~n8798;
  assign n8800 = pi657  & ~n8799;
  assign n8801 = ~n8796 & ~n8800;
  assign n8802 = ~n8795 & n8801;
  assign n8803 = n8795 & ~n8801;
  assign n8804 = ~n8802 & ~n8803;
  assign n8805 = ~pi657  & ~n8799;
  assign n8806 = pi657  & n8799;
  assign n8807 = ~n8805 & ~n8806;
  assign n8808 = ~pi660  & ~n8793;
  assign n8809 = pi660  & n8793;
  assign n8810 = ~n8808 & ~n8809;
  assign n8811 = ~n8807 & ~n8810;
  assign n8812 = ~n8804 & n8811;
  assign n8813 = ~n8795 & ~n8801;
  assign n8814 = ~n8812 & ~n8813;
  assign n8815 = pi664  & pi665 ;
  assign n8816 = ~pi664  & pi665 ;
  assign n8817 = pi664  & ~pi665 ;
  assign n8818 = ~n8816 & ~n8817;
  assign n8819 = pi666  & ~n8818;
  assign n8820 = ~n8815 & ~n8819;
  assign n8821 = pi661  & pi662 ;
  assign n8822 = ~pi661  & pi662 ;
  assign n8823 = pi661  & ~pi662 ;
  assign n8824 = ~n8822 & ~n8823;
  assign n8825 = pi663  & ~n8824;
  assign n8826 = ~n8821 & ~n8825;
  assign n8827 = ~n8820 & n8826;
  assign n8828 = n8820 & ~n8826;
  assign n8829 = ~n8827 & ~n8828;
  assign n8830 = ~pi663  & ~n8824;
  assign n8831 = pi663  & n8824;
  assign n8832 = ~n8830 & ~n8831;
  assign n8833 = ~pi666  & ~n8818;
  assign n8834 = pi666  & n8818;
  assign n8835 = ~n8833 & ~n8834;
  assign n8836 = ~n8832 & ~n8835;
  assign n8837 = ~n8829 & n8836;
  assign n8838 = ~n8820 & ~n8826;
  assign n8839 = ~n8837 & ~n8838;
  assign n8840 = n8829 & n8836;
  assign n8841 = ~n8829 & ~n8836;
  assign n8842 = ~n8840 & ~n8841;
  assign n8843 = n8804 & n8811;
  assign n8844 = ~n8804 & ~n8811;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = ~n8814 & ~n8845;
  assign n8847 = ~n8839 & ~n8842;
  assign n8848 = ~n8832 & n8835;
  assign n8849 = n8832 & ~n8835;
  assign n8850 = ~n8848 & ~n8849;
  assign n8851 = ~n8807 & n8810;
  assign n8852 = n8807 & ~n8810;
  assign n8853 = ~n8851 & ~n8852;
  assign n8854 = ~n8850 & ~n8853;
  assign n8855 = ~n8846 & n8854;
  assign n8856 = ~n8847 & n8855;
  assign n8857 = n8842 & ~n8856;
  assign n8858 = ~n8842 & n8856;
  assign n8859 = ~n8857 & ~n8858;
  assign n8860 = n8845 & n8859;
  assign n8861 = ~n8857 & ~n8860;
  assign n8862 = n8839 & ~n8861;
  assign n8863 = ~n8814 & ~n8862;
  assign n8864 = ~n8839 & n8861;
  assign n8865 = ~n8863 & ~n8864;
  assign n8866 = n8789 & n8865;
  assign n8867 = ~n8814 & n8839;
  assign n8868 = n8814 & ~n8839;
  assign n8869 = ~n8867 & ~n8868;
  assign n8870 = n8861 & ~n8869;
  assign n8871 = ~n8861 & n8869;
  assign n8872 = ~n8870 & ~n8871;
  assign n8873 = ~n8738 & n8763;
  assign n8874 = n8738 & ~n8763;
  assign n8875 = ~n8873 & ~n8874;
  assign n8876 = n8785 & ~n8875;
  assign n8877 = ~n8785 & n8875;
  assign n8878 = ~n8876 & ~n8877;
  assign n8879 = n8872 & n8878;
  assign n8880 = n8774 & ~n8777;
  assign n8881 = ~n8774 & n8777;
  assign n8882 = ~n8880 & ~n8881;
  assign n8883 = n8850 & ~n8853;
  assign n8884 = ~n8850 & n8853;
  assign n8885 = ~n8883 & ~n8884;
  assign n8886 = ~n8882 & ~n8885;
  assign n8887 = ~n8769 & ~n8783;
  assign n8888 = ~n8784 & ~n8887;
  assign n8889 = ~n8886 & n8888;
  assign n8890 = ~n8845 & ~n8859;
  assign n8891 = ~n8860 & ~n8890;
  assign n8892 = n8886 & ~n8888;
  assign n8893 = ~n8889 & ~n8892;
  assign n8894 = n8891 & n8893;
  assign n8895 = ~n8889 & ~n8894;
  assign n8896 = ~n8872 & ~n8878;
  assign n8897 = ~n8879 & ~n8896;
  assign n8898 = n8895 & n8897;
  assign n8899 = ~n8879 & ~n8898;
  assign n8900 = ~n8866 & ~n8899;
  assign n8901 = ~n8789 & ~n8865;
  assign n8902 = ~n8900 & ~n8901;
  assign n8903 = ~n8713 & ~n8902;
  assign n8904 = n8713 & n8902;
  assign n8905 = ~n8903 & ~n8904;
  assign n8906 = ~n8676 & ~n8712;
  assign n8907 = ~n8710 & n8906;
  assign n8908 = n8710 & ~n8906;
  assign n8909 = ~n8907 & ~n8908;
  assign n8910 = ~n8866 & ~n8901;
  assign n8911 = ~n8899 & n8910;
  assign n8912 = n8899 & ~n8910;
  assign n8913 = ~n8911 & ~n8912;
  assign n8914 = n8909 & n8913;
  assign n8915 = ~n8895 & ~n8897;
  assign n8916 = ~n8898 & ~n8915;
  assign n8917 = ~n8706 & ~n8708;
  assign n8918 = ~n8709 & ~n8917;
  assign n8919 = n8916 & n8918;
  assign n8920 = ~n8916 & ~n8918;
  assign n8921 = ~n8919 & ~n8920;
  assign n8922 = ~n8692 & n8695;
  assign n8923 = n8692 & ~n8695;
  assign n8924 = ~n8922 & ~n8923;
  assign n8925 = ~n8882 & n8885;
  assign n8926 = n8882 & ~n8885;
  assign n8927 = ~n8925 & ~n8926;
  assign n8928 = ~n8924 & ~n8927;
  assign n8929 = ~n8701 & n8704;
  assign n8930 = ~n8705 & ~n8929;
  assign n8931 = ~n8928 & n8930;
  assign n8932 = ~n8891 & ~n8893;
  assign n8933 = ~n8894 & ~n8932;
  assign n8934 = n8928 & ~n8930;
  assign n8935 = ~n8931 & ~n8934;
  assign n8936 = n8933 & n8935;
  assign n8937 = ~n8931 & ~n8936;
  assign n8938 = n8921 & n8937;
  assign n8939 = ~n8919 & ~n8938;
  assign n8940 = ~n8909 & ~n8913;
  assign n8941 = ~n8914 & ~n8940;
  assign n8942 = ~n8939 & n8941;
  assign n8943 = ~n8914 & ~n8942;
  assign n8944 = n8905 & ~n8943;
  assign n8945 = ~n8903 & ~n8944;
  assign n8946 = ~n8523 & ~n8945;
  assign n8947 = ~n8905 & n8943;
  assign n8948 = ~n8944 & ~n8947;
  assign n8949 = ~n8483 & n8521;
  assign n8950 = ~n8522 & ~n8949;
  assign n8951 = n8948 & n8950;
  assign n8952 = n8517 & ~n8519;
  assign n8953 = ~n8520 & ~n8952;
  assign n8954 = n8939 & ~n8941;
  assign n8955 = ~n8942 & ~n8954;
  assign n8956 = n8953 & n8955;
  assign n8957 = ~n8953 & ~n8955;
  assign n8958 = ~n8956 & ~n8957;
  assign n8959 = ~n8921 & ~n8937;
  assign n8960 = ~n8938 & ~n8959;
  assign n8961 = ~n8499 & ~n8515;
  assign n8962 = ~n8516 & ~n8961;
  assign n8963 = n8960 & n8962;
  assign n8964 = ~n8502 & n8505;
  assign n8965 = n8502 & ~n8505;
  assign n8966 = ~n8964 & ~n8965;
  assign n8967 = ~n8924 & n8927;
  assign n8968 = n8924 & ~n8927;
  assign n8969 = ~n8967 & ~n8968;
  assign n8970 = ~n8966 & ~n8969;
  assign n8971 = ~n8511 & ~n8513;
  assign n8972 = ~n8514 & ~n8971;
  assign n8973 = ~n8970 & n8972;
  assign n8974 = ~n8933 & ~n8935;
  assign n8975 = ~n8936 & ~n8974;
  assign n8976 = n8970 & ~n8972;
  assign n8977 = ~n8973 & ~n8976;
  assign n8978 = n8975 & n8977;
  assign n8979 = ~n8973 & ~n8978;
  assign n8980 = ~n8960 & ~n8962;
  assign n8981 = ~n8963 & ~n8980;
  assign n8982 = n8979 & n8981;
  assign n8983 = ~n8963 & ~n8982;
  assign n8984 = n8958 & ~n8983;
  assign n8985 = ~n8956 & ~n8984;
  assign n8986 = ~n8948 & ~n8950;
  assign n8987 = ~n8951 & ~n8986;
  assign n8988 = ~n8985 & n8987;
  assign n8989 = ~n8951 & ~n8988;
  assign n8990 = n8523 & n8945;
  assign n8991 = ~n8946 & ~n8990;
  assign n8992 = ~n8989 & n8991;
  assign n8993 = ~n8946 & ~n8992;
  assign n8994 = ~n8101 & ~n8993;
  assign n8995 = n8101 & n8993;
  assign n8996 = ~n8994 & ~n8995;
  assign n8997 = n8097 & ~n8099;
  assign n8998 = ~n8100 & ~n8997;
  assign n8999 = n8989 & ~n8991;
  assign n9000 = ~n8992 & ~n8999;
  assign n9001 = n8998 & n9000;
  assign n9002 = ~n8979 & ~n8981;
  assign n9003 = ~n8982 & ~n9002;
  assign n9004 = ~n8073 & ~n8089;
  assign n9005 = ~n8090 & ~n9004;
  assign n9006 = n9003 & n9005;
  assign n9007 = ~n8076 & n8079;
  assign n9008 = n8076 & ~n8079;
  assign n9009 = ~n9007 & ~n9008;
  assign n9010 = ~n8966 & n8969;
  assign n9011 = n8966 & ~n8969;
  assign n9012 = ~n9010 & ~n9011;
  assign n9013 = ~n9009 & ~n9012;
  assign n9014 = ~n8085 & ~n8087;
  assign n9015 = ~n8088 & ~n9014;
  assign n9016 = n9013 & ~n9015;
  assign n9017 = ~n8975 & ~n8977;
  assign n9018 = ~n8978 & ~n9017;
  assign n9019 = ~n9013 & n9015;
  assign n9020 = ~n9018 & ~n9019;
  assign n9021 = ~n9016 & ~n9020;
  assign n9022 = ~n9003 & ~n9005;
  assign n9023 = ~n9006 & ~n9022;
  assign n9024 = ~n9021 & n9023;
  assign n9025 = ~n9006 & ~n9024;
  assign n9026 = ~n8066 & n8091;
  assign n9027 = ~n8092 & ~n9026;
  assign n9028 = ~n8958 & n8983;
  assign n9029 = ~n8984 & ~n9028;
  assign n9030 = ~n9027 & ~n9029;
  assign n9031 = ~n9025 & ~n9030;
  assign n9032 = n9027 & n9029;
  assign n9033 = ~n9031 & ~n9032;
  assign n9034 = n8985 & ~n8987;
  assign n9035 = ~n8988 & ~n9034;
  assign n9036 = n8093 & ~n8095;
  assign n9037 = ~n8096 & ~n9036;
  assign n9038 = ~n9035 & ~n9037;
  assign n9039 = ~n9033 & ~n9038;
  assign n9040 = n9035 & n9037;
  assign n9041 = ~n9039 & ~n9040;
  assign n9042 = ~n8998 & ~n9000;
  assign n9043 = ~n9001 & ~n9042;
  assign n9044 = ~n9041 & n9043;
  assign n9045 = ~n9001 & ~n9044;
  assign n9046 = n8996 & ~n9045;
  assign n9047 = ~n8994 & ~n9046;
  assign n9048 = pi646  & pi647 ;
  assign n9049 = ~pi646  & pi647 ;
  assign n9050 = pi646  & ~pi647 ;
  assign n9051 = ~n9049 & ~n9050;
  assign n9052 = pi648  & ~n9051;
  assign n9053 = ~n9048 & ~n9052;
  assign n9054 = pi643  & pi644 ;
  assign n9055 = ~pi643  & pi644 ;
  assign n9056 = pi643  & ~pi644 ;
  assign n9057 = ~n9055 & ~n9056;
  assign n9058 = pi645  & ~n9057;
  assign n9059 = ~n9054 & ~n9058;
  assign n9060 = ~n9053 & n9059;
  assign n9061 = n9053 & ~n9059;
  assign n9062 = ~n9060 & ~n9061;
  assign n9063 = ~pi645  & ~n9057;
  assign n9064 = pi645  & n9057;
  assign n9065 = ~n9063 & ~n9064;
  assign n9066 = ~pi648  & ~n9051;
  assign n9067 = pi648  & n9051;
  assign n9068 = ~n9066 & ~n9067;
  assign n9069 = ~n9065 & ~n9068;
  assign n9070 = ~n9062 & n9069;
  assign n9071 = ~n9053 & ~n9059;
  assign n9072 = ~n9070 & ~n9071;
  assign n9073 = pi652  & pi653 ;
  assign n9074 = ~pi652  & pi653 ;
  assign n9075 = pi652  & ~pi653 ;
  assign n9076 = ~n9074 & ~n9075;
  assign n9077 = pi654  & ~n9076;
  assign n9078 = ~n9073 & ~n9077;
  assign n9079 = pi649  & pi650 ;
  assign n9080 = ~pi649  & pi650 ;
  assign n9081 = pi649  & ~pi650 ;
  assign n9082 = ~n9080 & ~n9081;
  assign n9083 = pi651  & ~n9082;
  assign n9084 = ~n9079 & ~n9083;
  assign n9085 = ~n9078 & n9084;
  assign n9086 = n9078 & ~n9084;
  assign n9087 = ~n9085 & ~n9086;
  assign n9088 = ~pi651  & ~n9082;
  assign n9089 = pi651  & n9082;
  assign n9090 = ~n9088 & ~n9089;
  assign n9091 = ~pi654  & ~n9076;
  assign n9092 = pi654  & n9076;
  assign n9093 = ~n9091 & ~n9092;
  assign n9094 = ~n9090 & ~n9093;
  assign n9095 = ~n9087 & n9094;
  assign n9096 = ~n9078 & ~n9084;
  assign n9097 = ~n9095 & ~n9096;
  assign n9098 = n9087 & n9094;
  assign n9099 = ~n9087 & ~n9094;
  assign n9100 = ~n9098 & ~n9099;
  assign n9101 = n9062 & n9069;
  assign n9102 = ~n9062 & ~n9069;
  assign n9103 = ~n9101 & ~n9102;
  assign n9104 = ~n9072 & ~n9103;
  assign n9105 = ~n9097 & ~n9100;
  assign n9106 = ~n9090 & n9093;
  assign n9107 = n9090 & ~n9093;
  assign n9108 = ~n9106 & ~n9107;
  assign n9109 = ~n9065 & n9068;
  assign n9110 = n9065 & ~n9068;
  assign n9111 = ~n9109 & ~n9110;
  assign n9112 = ~n9108 & ~n9111;
  assign n9113 = ~n9104 & n9112;
  assign n9114 = ~n9105 & n9113;
  assign n9115 = n9100 & ~n9114;
  assign n9116 = ~n9100 & n9114;
  assign n9117 = ~n9115 & ~n9116;
  assign n9118 = n9103 & n9117;
  assign n9119 = ~n9115 & ~n9118;
  assign n9120 = n9097 & ~n9119;
  assign n9121 = ~n9072 & ~n9120;
  assign n9122 = ~n9097 & n9119;
  assign n9123 = ~n9121 & ~n9122;
  assign n9124 = pi634  & pi635 ;
  assign n9125 = ~pi634  & pi635 ;
  assign n9126 = pi634  & ~pi635 ;
  assign n9127 = ~n9125 & ~n9126;
  assign n9128 = pi636  & ~n9127;
  assign n9129 = ~n9124 & ~n9128;
  assign n9130 = pi631  & pi632 ;
  assign n9131 = ~pi631  & pi632 ;
  assign n9132 = pi631  & ~pi632 ;
  assign n9133 = ~n9131 & ~n9132;
  assign n9134 = pi633  & ~n9133;
  assign n9135 = ~n9130 & ~n9134;
  assign n9136 = ~n9129 & n9135;
  assign n9137 = n9129 & ~n9135;
  assign n9138 = ~n9136 & ~n9137;
  assign n9139 = ~pi633  & ~n9133;
  assign n9140 = pi633  & n9133;
  assign n9141 = ~n9139 & ~n9140;
  assign n9142 = ~pi636  & ~n9127;
  assign n9143 = pi636  & n9127;
  assign n9144 = ~n9142 & ~n9143;
  assign n9145 = ~n9141 & ~n9144;
  assign n9146 = ~n9138 & n9145;
  assign n9147 = ~n9129 & ~n9135;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = pi640  & pi641 ;
  assign n9150 = ~pi640  & pi641 ;
  assign n9151 = pi640  & ~pi641 ;
  assign n9152 = ~n9150 & ~n9151;
  assign n9153 = pi642  & ~n9152;
  assign n9154 = ~n9149 & ~n9153;
  assign n9155 = pi637  & pi638 ;
  assign n9156 = ~pi637  & pi638 ;
  assign n9157 = pi637  & ~pi638 ;
  assign n9158 = ~n9156 & ~n9157;
  assign n9159 = pi639  & ~n9158;
  assign n9160 = ~n9155 & ~n9159;
  assign n9161 = ~n9154 & n9160;
  assign n9162 = n9154 & ~n9160;
  assign n9163 = ~n9161 & ~n9162;
  assign n9164 = ~pi639  & ~n9158;
  assign n9165 = pi639  & n9158;
  assign n9166 = ~n9164 & ~n9165;
  assign n9167 = ~pi642  & ~n9152;
  assign n9168 = pi642  & n9152;
  assign n9169 = ~n9167 & ~n9168;
  assign n9170 = ~n9166 & ~n9169;
  assign n9171 = ~n9163 & n9170;
  assign n9172 = ~n9154 & ~n9160;
  assign n9173 = ~n9171 & ~n9172;
  assign n9174 = n9163 & n9170;
  assign n9175 = ~n9163 & ~n9170;
  assign n9176 = ~n9174 & ~n9175;
  assign n9177 = n9138 & n9145;
  assign n9178 = ~n9138 & ~n9145;
  assign n9179 = ~n9177 & ~n9178;
  assign n9180 = ~n9148 & ~n9179;
  assign n9181 = ~n9173 & ~n9176;
  assign n9182 = ~n9166 & n9169;
  assign n9183 = n9166 & ~n9169;
  assign n9184 = ~n9182 & ~n9183;
  assign n9185 = ~n9141 & n9144;
  assign n9186 = n9141 & ~n9144;
  assign n9187 = ~n9185 & ~n9186;
  assign n9188 = ~n9184 & ~n9187;
  assign n9189 = ~n9180 & n9188;
  assign n9190 = ~n9181 & n9189;
  assign n9191 = n9176 & ~n9190;
  assign n9192 = ~n9176 & n9190;
  assign n9193 = ~n9191 & ~n9192;
  assign n9194 = n9179 & n9193;
  assign n9195 = ~n9191 & ~n9194;
  assign n9196 = n9173 & ~n9195;
  assign n9197 = ~n9148 & ~n9196;
  assign n9198 = ~n9173 & n9195;
  assign n9199 = ~n9197 & ~n9198;
  assign n9200 = n9123 & n9199;
  assign n9201 = ~n9148 & n9173;
  assign n9202 = n9148 & ~n9173;
  assign n9203 = ~n9201 & ~n9202;
  assign n9204 = n9195 & ~n9203;
  assign n9205 = ~n9195 & n9203;
  assign n9206 = ~n9204 & ~n9205;
  assign n9207 = ~n9072 & n9097;
  assign n9208 = n9072 & ~n9097;
  assign n9209 = ~n9207 & ~n9208;
  assign n9210 = n9119 & ~n9209;
  assign n9211 = ~n9119 & n9209;
  assign n9212 = ~n9210 & ~n9211;
  assign n9213 = n9206 & n9212;
  assign n9214 = n9108 & ~n9111;
  assign n9215 = ~n9108 & n9111;
  assign n9216 = ~n9214 & ~n9215;
  assign n9217 = n9184 & ~n9187;
  assign n9218 = ~n9184 & n9187;
  assign n9219 = ~n9217 & ~n9218;
  assign n9220 = ~n9216 & ~n9219;
  assign n9221 = ~n9103 & ~n9117;
  assign n9222 = ~n9118 & ~n9221;
  assign n9223 = ~n9220 & n9222;
  assign n9224 = ~n9179 & ~n9193;
  assign n9225 = ~n9194 & ~n9224;
  assign n9226 = ~n9220 & ~n9222;
  assign n9227 = n9222 & ~n9223;
  assign n9228 = ~n9226 & ~n9227;
  assign n9229 = n9225 & ~n9228;
  assign n9230 = ~n9223 & ~n9229;
  assign n9231 = ~n9206 & ~n9212;
  assign n9232 = ~n9213 & ~n9231;
  assign n9233 = n9230 & n9232;
  assign n9234 = ~n9213 & ~n9233;
  assign n9235 = ~n9200 & ~n9234;
  assign n9236 = ~n9123 & ~n9199;
  assign n9237 = ~n9235 & ~n9236;
  assign n9238 = pi622  & pi623 ;
  assign n9239 = ~pi622  & pi623 ;
  assign n9240 = pi622  & ~pi623 ;
  assign n9241 = ~n9239 & ~n9240;
  assign n9242 = pi624  & ~n9241;
  assign n9243 = ~n9238 & ~n9242;
  assign n9244 = pi619  & pi620 ;
  assign n9245 = ~pi619  & pi620 ;
  assign n9246 = pi619  & ~pi620 ;
  assign n9247 = ~n9245 & ~n9246;
  assign n9248 = pi621  & ~n9247;
  assign n9249 = ~n9244 & ~n9248;
  assign n9250 = ~n9243 & n9249;
  assign n9251 = n9243 & ~n9249;
  assign n9252 = ~n9250 & ~n9251;
  assign n9253 = ~pi621  & ~n9247;
  assign n9254 = pi621  & n9247;
  assign n9255 = ~n9253 & ~n9254;
  assign n9256 = ~pi624  & ~n9241;
  assign n9257 = pi624  & n9241;
  assign n9258 = ~n9256 & ~n9257;
  assign n9259 = ~n9255 & ~n9258;
  assign n9260 = ~n9252 & n9259;
  assign n9261 = ~n9243 & ~n9249;
  assign n9262 = ~n9260 & ~n9261;
  assign n9263 = pi628  & pi629 ;
  assign n9264 = ~pi628  & pi629 ;
  assign n9265 = pi628  & ~pi629 ;
  assign n9266 = ~n9264 & ~n9265;
  assign n9267 = pi630  & ~n9266;
  assign n9268 = ~n9263 & ~n9267;
  assign n9269 = pi625  & pi626 ;
  assign n9270 = ~pi625  & pi626 ;
  assign n9271 = pi625  & ~pi626 ;
  assign n9272 = ~n9270 & ~n9271;
  assign n9273 = pi627  & ~n9272;
  assign n9274 = ~n9269 & ~n9273;
  assign n9275 = ~n9268 & n9274;
  assign n9276 = n9268 & ~n9274;
  assign n9277 = ~n9275 & ~n9276;
  assign n9278 = ~pi627  & ~n9272;
  assign n9279 = pi627  & n9272;
  assign n9280 = ~n9278 & ~n9279;
  assign n9281 = ~pi630  & ~n9266;
  assign n9282 = pi630  & n9266;
  assign n9283 = ~n9281 & ~n9282;
  assign n9284 = ~n9280 & ~n9283;
  assign n9285 = ~n9277 & n9284;
  assign n9286 = ~n9268 & ~n9274;
  assign n9287 = ~n9285 & ~n9286;
  assign n9288 = n9277 & n9284;
  assign n9289 = ~n9277 & ~n9284;
  assign n9290 = ~n9288 & ~n9289;
  assign n9291 = n9252 & n9259;
  assign n9292 = ~n9252 & ~n9259;
  assign n9293 = ~n9291 & ~n9292;
  assign n9294 = ~n9262 & ~n9293;
  assign n9295 = ~n9287 & ~n9290;
  assign n9296 = ~n9280 & n9283;
  assign n9297 = n9280 & ~n9283;
  assign n9298 = ~n9296 & ~n9297;
  assign n9299 = ~n9255 & n9258;
  assign n9300 = n9255 & ~n9258;
  assign n9301 = ~n9299 & ~n9300;
  assign n9302 = ~n9298 & ~n9301;
  assign n9303 = ~n9294 & n9302;
  assign n9304 = ~n9295 & n9303;
  assign n9305 = n9290 & ~n9304;
  assign n9306 = ~n9290 & n9304;
  assign n9307 = ~n9305 & ~n9306;
  assign n9308 = n9293 & n9307;
  assign n9309 = ~n9305 & ~n9308;
  assign n9310 = n9287 & ~n9309;
  assign n9311 = ~n9262 & ~n9310;
  assign n9312 = ~n9287 & n9309;
  assign n9313 = ~n9311 & ~n9312;
  assign n9314 = pi610  & pi611 ;
  assign n9315 = ~pi610  & pi611 ;
  assign n9316 = pi610  & ~pi611 ;
  assign n9317 = ~n9315 & ~n9316;
  assign n9318 = pi612  & ~n9317;
  assign n9319 = ~n9314 & ~n9318;
  assign n9320 = pi607  & pi608 ;
  assign n9321 = ~pi607  & pi608 ;
  assign n9322 = pi607  & ~pi608 ;
  assign n9323 = ~n9321 & ~n9322;
  assign n9324 = pi609  & ~n9323;
  assign n9325 = ~n9320 & ~n9324;
  assign n9326 = ~n9319 & n9325;
  assign n9327 = n9319 & ~n9325;
  assign n9328 = ~n9326 & ~n9327;
  assign n9329 = ~pi609  & ~n9323;
  assign n9330 = pi609  & n9323;
  assign n9331 = ~n9329 & ~n9330;
  assign n9332 = ~pi612  & ~n9317;
  assign n9333 = pi612  & n9317;
  assign n9334 = ~n9332 & ~n9333;
  assign n9335 = ~n9331 & ~n9334;
  assign n9336 = ~n9328 & n9335;
  assign n9337 = ~n9319 & ~n9325;
  assign n9338 = ~n9336 & ~n9337;
  assign n9339 = pi616  & pi617 ;
  assign n9340 = ~pi616  & pi617 ;
  assign n9341 = pi616  & ~pi617 ;
  assign n9342 = ~n9340 & ~n9341;
  assign n9343 = pi618  & ~n9342;
  assign n9344 = ~n9339 & ~n9343;
  assign n9345 = pi613  & pi614 ;
  assign n9346 = ~pi613  & pi614 ;
  assign n9347 = pi613  & ~pi614 ;
  assign n9348 = ~n9346 & ~n9347;
  assign n9349 = pi615  & ~n9348;
  assign n9350 = ~n9345 & ~n9349;
  assign n9351 = ~n9344 & n9350;
  assign n9352 = n9344 & ~n9350;
  assign n9353 = ~n9351 & ~n9352;
  assign n9354 = ~pi615  & ~n9348;
  assign n9355 = pi615  & n9348;
  assign n9356 = ~n9354 & ~n9355;
  assign n9357 = ~pi618  & ~n9342;
  assign n9358 = pi618  & n9342;
  assign n9359 = ~n9357 & ~n9358;
  assign n9360 = ~n9356 & ~n9359;
  assign n9361 = ~n9353 & n9360;
  assign n9362 = ~n9344 & ~n9350;
  assign n9363 = ~n9361 & ~n9362;
  assign n9364 = n9353 & n9360;
  assign n9365 = ~n9353 & ~n9360;
  assign n9366 = ~n9364 & ~n9365;
  assign n9367 = n9328 & n9335;
  assign n9368 = ~n9328 & ~n9335;
  assign n9369 = ~n9367 & ~n9368;
  assign n9370 = ~n9338 & ~n9369;
  assign n9371 = ~n9363 & ~n9366;
  assign n9372 = ~n9356 & n9359;
  assign n9373 = n9356 & ~n9359;
  assign n9374 = ~n9372 & ~n9373;
  assign n9375 = ~n9331 & n9334;
  assign n9376 = n9331 & ~n9334;
  assign n9377 = ~n9375 & ~n9376;
  assign n9378 = ~n9374 & ~n9377;
  assign n9379 = ~n9370 & n9378;
  assign n9380 = ~n9371 & n9379;
  assign n9381 = n9366 & ~n9380;
  assign n9382 = ~n9366 & n9380;
  assign n9383 = ~n9381 & ~n9382;
  assign n9384 = n9369 & n9383;
  assign n9385 = ~n9381 & ~n9384;
  assign n9386 = n9363 & ~n9385;
  assign n9387 = ~n9338 & ~n9386;
  assign n9388 = ~n9363 & n9385;
  assign n9389 = ~n9387 & ~n9388;
  assign n9390 = n9313 & n9389;
  assign n9391 = ~n9338 & n9363;
  assign n9392 = n9338 & ~n9363;
  assign n9393 = ~n9391 & ~n9392;
  assign n9394 = n9385 & ~n9393;
  assign n9395 = ~n9385 & n9393;
  assign n9396 = ~n9394 & ~n9395;
  assign n9397 = ~n9262 & n9287;
  assign n9398 = n9262 & ~n9287;
  assign n9399 = ~n9397 & ~n9398;
  assign n9400 = n9309 & ~n9399;
  assign n9401 = ~n9309 & n9399;
  assign n9402 = ~n9400 & ~n9401;
  assign n9403 = n9396 & n9402;
  assign n9404 = n9298 & ~n9301;
  assign n9405 = ~n9298 & n9301;
  assign n9406 = ~n9404 & ~n9405;
  assign n9407 = n9374 & ~n9377;
  assign n9408 = ~n9374 & n9377;
  assign n9409 = ~n9407 & ~n9408;
  assign n9410 = ~n9406 & ~n9409;
  assign n9411 = ~n9293 & ~n9307;
  assign n9412 = ~n9308 & ~n9411;
  assign n9413 = ~n9410 & n9412;
  assign n9414 = ~n9369 & ~n9383;
  assign n9415 = ~n9384 & ~n9414;
  assign n9416 = n9410 & ~n9412;
  assign n9417 = ~n9413 & ~n9416;
  assign n9418 = n9415 & n9417;
  assign n9419 = ~n9413 & ~n9418;
  assign n9420 = ~n9396 & ~n9402;
  assign n9421 = ~n9403 & ~n9420;
  assign n9422 = n9419 & n9421;
  assign n9423 = ~n9403 & ~n9422;
  assign n9424 = ~n9390 & ~n9423;
  assign n9425 = ~n9313 & ~n9389;
  assign n9426 = ~n9424 & ~n9425;
  assign n9427 = ~n9237 & ~n9426;
  assign n9428 = n9237 & n9426;
  assign n9429 = ~n9427 & ~n9428;
  assign n9430 = ~n9200 & ~n9236;
  assign n9431 = ~n9234 & n9430;
  assign n9432 = n9234 & ~n9430;
  assign n9433 = ~n9431 & ~n9432;
  assign n9434 = ~n9390 & ~n9425;
  assign n9435 = ~n9423 & n9434;
  assign n9436 = n9423 & ~n9434;
  assign n9437 = ~n9435 & ~n9436;
  assign n9438 = n9433 & n9437;
  assign n9439 = ~n9419 & ~n9421;
  assign n9440 = ~n9422 & ~n9439;
  assign n9441 = ~n9230 & ~n9232;
  assign n9442 = ~n9233 & ~n9441;
  assign n9443 = n9440 & n9442;
  assign n9444 = ~n9440 & ~n9442;
  assign n9445 = ~n9443 & ~n9444;
  assign n9446 = ~n9216 & n9219;
  assign n9447 = n9216 & ~n9219;
  assign n9448 = ~n9446 & ~n9447;
  assign n9449 = ~n9406 & n9409;
  assign n9450 = n9406 & ~n9409;
  assign n9451 = ~n9449 & ~n9450;
  assign n9452 = ~n9448 & ~n9451;
  assign n9453 = ~n9225 & n9228;
  assign n9454 = ~n9229 & ~n9453;
  assign n9455 = ~n9452 & n9454;
  assign n9456 = ~n9415 & ~n9417;
  assign n9457 = ~n9418 & ~n9456;
  assign n9458 = n9452 & ~n9454;
  assign n9459 = ~n9455 & ~n9458;
  assign n9460 = n9457 & n9459;
  assign n9461 = ~n9455 & ~n9460;
  assign n9462 = n9445 & n9461;
  assign n9463 = ~n9443 & ~n9462;
  assign n9464 = ~n9433 & ~n9437;
  assign n9465 = ~n9438 & ~n9464;
  assign n9466 = ~n9463 & n9465;
  assign n9467 = ~n9438 & ~n9466;
  assign n9468 = n9429 & ~n9467;
  assign n9469 = ~n9427 & ~n9468;
  assign n9470 = pi598  & pi599 ;
  assign n9471 = ~pi598  & pi599 ;
  assign n9472 = pi598  & ~pi599 ;
  assign n9473 = ~n9471 & ~n9472;
  assign n9474 = pi600  & ~n9473;
  assign n9475 = ~n9470 & ~n9474;
  assign n9476 = pi595  & pi596 ;
  assign n9477 = ~pi595  & pi596 ;
  assign n9478 = pi595  & ~pi596 ;
  assign n9479 = ~n9477 & ~n9478;
  assign n9480 = pi597  & ~n9479;
  assign n9481 = ~n9476 & ~n9480;
  assign n9482 = ~n9475 & n9481;
  assign n9483 = n9475 & ~n9481;
  assign n9484 = ~n9482 & ~n9483;
  assign n9485 = ~pi597  & ~n9479;
  assign n9486 = pi597  & n9479;
  assign n9487 = ~n9485 & ~n9486;
  assign n9488 = ~pi600  & ~n9473;
  assign n9489 = pi600  & n9473;
  assign n9490 = ~n9488 & ~n9489;
  assign n9491 = ~n9487 & ~n9490;
  assign n9492 = ~n9484 & n9491;
  assign n9493 = ~n9475 & ~n9481;
  assign n9494 = ~n9492 & ~n9493;
  assign n9495 = pi604  & pi605 ;
  assign n9496 = ~pi604  & pi605 ;
  assign n9497 = pi604  & ~pi605 ;
  assign n9498 = ~n9496 & ~n9497;
  assign n9499 = pi606  & ~n9498;
  assign n9500 = ~n9495 & ~n9499;
  assign n9501 = pi601  & pi602 ;
  assign n9502 = ~pi601  & pi602 ;
  assign n9503 = pi601  & ~pi602 ;
  assign n9504 = ~n9502 & ~n9503;
  assign n9505 = pi603  & ~n9504;
  assign n9506 = ~n9501 & ~n9505;
  assign n9507 = ~n9500 & n9506;
  assign n9508 = n9500 & ~n9506;
  assign n9509 = ~n9507 & ~n9508;
  assign n9510 = ~pi603  & ~n9504;
  assign n9511 = pi603  & n9504;
  assign n9512 = ~n9510 & ~n9511;
  assign n9513 = ~pi606  & ~n9498;
  assign n9514 = pi606  & n9498;
  assign n9515 = ~n9513 & ~n9514;
  assign n9516 = ~n9512 & ~n9515;
  assign n9517 = ~n9509 & n9516;
  assign n9518 = ~n9500 & ~n9506;
  assign n9519 = ~n9517 & ~n9518;
  assign n9520 = n9509 & n9516;
  assign n9521 = ~n9509 & ~n9516;
  assign n9522 = ~n9520 & ~n9521;
  assign n9523 = n9484 & n9491;
  assign n9524 = ~n9484 & ~n9491;
  assign n9525 = ~n9523 & ~n9524;
  assign n9526 = ~n9494 & ~n9525;
  assign n9527 = ~n9519 & ~n9522;
  assign n9528 = ~n9512 & n9515;
  assign n9529 = n9512 & ~n9515;
  assign n9530 = ~n9528 & ~n9529;
  assign n9531 = ~n9487 & n9490;
  assign n9532 = n9487 & ~n9490;
  assign n9533 = ~n9531 & ~n9532;
  assign n9534 = ~n9530 & ~n9533;
  assign n9535 = ~n9526 & n9534;
  assign n9536 = ~n9527 & n9535;
  assign n9537 = n9522 & ~n9536;
  assign n9538 = ~n9522 & n9536;
  assign n9539 = ~n9537 & ~n9538;
  assign n9540 = n9525 & n9539;
  assign n9541 = ~n9537 & ~n9540;
  assign n9542 = n9519 & ~n9541;
  assign n9543 = ~n9494 & ~n9542;
  assign n9544 = ~n9519 & n9541;
  assign n9545 = ~n9543 & ~n9544;
  assign n9546 = pi586  & pi587 ;
  assign n9547 = ~pi586  & pi587 ;
  assign n9548 = pi586  & ~pi587 ;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = pi588  & ~n9549;
  assign n9551 = ~n9546 & ~n9550;
  assign n9552 = pi583  & pi584 ;
  assign n9553 = ~pi583  & pi584 ;
  assign n9554 = pi583  & ~pi584 ;
  assign n9555 = ~n9553 & ~n9554;
  assign n9556 = pi585  & ~n9555;
  assign n9557 = ~n9552 & ~n9556;
  assign n9558 = ~n9551 & n9557;
  assign n9559 = n9551 & ~n9557;
  assign n9560 = ~n9558 & ~n9559;
  assign n9561 = ~pi585  & ~n9555;
  assign n9562 = pi585  & n9555;
  assign n9563 = ~n9561 & ~n9562;
  assign n9564 = ~pi588  & ~n9549;
  assign n9565 = pi588  & n9549;
  assign n9566 = ~n9564 & ~n9565;
  assign n9567 = ~n9563 & ~n9566;
  assign n9568 = ~n9560 & n9567;
  assign n9569 = ~n9551 & ~n9557;
  assign n9570 = ~n9568 & ~n9569;
  assign n9571 = pi592  & pi593 ;
  assign n9572 = ~pi592  & pi593 ;
  assign n9573 = pi592  & ~pi593 ;
  assign n9574 = ~n9572 & ~n9573;
  assign n9575 = pi594  & ~n9574;
  assign n9576 = ~n9571 & ~n9575;
  assign n9577 = pi589  & pi590 ;
  assign n9578 = ~pi589  & pi590 ;
  assign n9579 = pi589  & ~pi590 ;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = pi591  & ~n9580;
  assign n9582 = ~n9577 & ~n9581;
  assign n9583 = ~n9576 & n9582;
  assign n9584 = n9576 & ~n9582;
  assign n9585 = ~n9583 & ~n9584;
  assign n9586 = ~pi591  & ~n9580;
  assign n9587 = pi591  & n9580;
  assign n9588 = ~n9586 & ~n9587;
  assign n9589 = ~pi594  & ~n9574;
  assign n9590 = pi594  & n9574;
  assign n9591 = ~n9589 & ~n9590;
  assign n9592 = ~n9588 & ~n9591;
  assign n9593 = ~n9585 & n9592;
  assign n9594 = ~n9576 & ~n9582;
  assign n9595 = ~n9593 & ~n9594;
  assign n9596 = n9585 & n9592;
  assign n9597 = ~n9585 & ~n9592;
  assign n9598 = ~n9596 & ~n9597;
  assign n9599 = n9560 & n9567;
  assign n9600 = ~n9560 & ~n9567;
  assign n9601 = ~n9599 & ~n9600;
  assign n9602 = ~n9570 & ~n9601;
  assign n9603 = ~n9595 & ~n9598;
  assign n9604 = ~n9588 & n9591;
  assign n9605 = n9588 & ~n9591;
  assign n9606 = ~n9604 & ~n9605;
  assign n9607 = ~n9563 & n9566;
  assign n9608 = n9563 & ~n9566;
  assign n9609 = ~n9607 & ~n9608;
  assign n9610 = ~n9606 & ~n9609;
  assign n9611 = ~n9602 & n9610;
  assign n9612 = ~n9603 & n9611;
  assign n9613 = n9598 & ~n9612;
  assign n9614 = ~n9598 & n9612;
  assign n9615 = ~n9613 & ~n9614;
  assign n9616 = n9601 & n9615;
  assign n9617 = ~n9613 & ~n9616;
  assign n9618 = n9595 & ~n9617;
  assign n9619 = ~n9570 & ~n9618;
  assign n9620 = ~n9595 & n9617;
  assign n9621 = ~n9619 & ~n9620;
  assign n9622 = n9545 & n9621;
  assign n9623 = ~n9570 & n9595;
  assign n9624 = n9570 & ~n9595;
  assign n9625 = ~n9623 & ~n9624;
  assign n9626 = n9617 & ~n9625;
  assign n9627 = ~n9617 & n9625;
  assign n9628 = ~n9626 & ~n9627;
  assign n9629 = ~n9494 & n9519;
  assign n9630 = n9494 & ~n9519;
  assign n9631 = ~n9629 & ~n9630;
  assign n9632 = n9541 & ~n9631;
  assign n9633 = ~n9541 & n9631;
  assign n9634 = ~n9632 & ~n9633;
  assign n9635 = n9628 & n9634;
  assign n9636 = n9530 & ~n9533;
  assign n9637 = ~n9530 & n9533;
  assign n9638 = ~n9636 & ~n9637;
  assign n9639 = n9606 & ~n9609;
  assign n9640 = ~n9606 & n9609;
  assign n9641 = ~n9639 & ~n9640;
  assign n9642 = ~n9638 & ~n9641;
  assign n9643 = ~n9525 & ~n9539;
  assign n9644 = ~n9540 & ~n9643;
  assign n9645 = ~n9642 & n9644;
  assign n9646 = ~n9601 & ~n9615;
  assign n9647 = ~n9616 & ~n9646;
  assign n9648 = ~n9642 & ~n9644;
  assign n9649 = n9644 & ~n9645;
  assign n9650 = ~n9648 & ~n9649;
  assign n9651 = n9647 & ~n9650;
  assign n9652 = ~n9645 & ~n9651;
  assign n9653 = ~n9628 & ~n9634;
  assign n9654 = ~n9635 & ~n9653;
  assign n9655 = n9652 & n9654;
  assign n9656 = ~n9635 & ~n9655;
  assign n9657 = ~n9622 & ~n9656;
  assign n9658 = ~n9545 & ~n9621;
  assign n9659 = ~n9657 & ~n9658;
  assign n9660 = pi574  & pi575 ;
  assign n9661 = ~pi574  & pi575 ;
  assign n9662 = pi574  & ~pi575 ;
  assign n9663 = ~n9661 & ~n9662;
  assign n9664 = pi576  & ~n9663;
  assign n9665 = ~n9660 & ~n9664;
  assign n9666 = pi571  & pi572 ;
  assign n9667 = ~pi571  & pi572 ;
  assign n9668 = pi571  & ~pi572 ;
  assign n9669 = ~n9667 & ~n9668;
  assign n9670 = pi573  & ~n9669;
  assign n9671 = ~n9666 & ~n9670;
  assign n9672 = ~n9665 & n9671;
  assign n9673 = n9665 & ~n9671;
  assign n9674 = ~n9672 & ~n9673;
  assign n9675 = ~pi573  & ~n9669;
  assign n9676 = pi573  & n9669;
  assign n9677 = ~n9675 & ~n9676;
  assign n9678 = ~pi576  & ~n9663;
  assign n9679 = pi576  & n9663;
  assign n9680 = ~n9678 & ~n9679;
  assign n9681 = ~n9677 & ~n9680;
  assign n9682 = ~n9674 & n9681;
  assign n9683 = ~n9665 & ~n9671;
  assign n9684 = ~n9682 & ~n9683;
  assign n9685 = pi580  & pi581 ;
  assign n9686 = ~pi580  & pi581 ;
  assign n9687 = pi580  & ~pi581 ;
  assign n9688 = ~n9686 & ~n9687;
  assign n9689 = pi582  & ~n9688;
  assign n9690 = ~n9685 & ~n9689;
  assign n9691 = pi577  & pi578 ;
  assign n9692 = ~pi577  & pi578 ;
  assign n9693 = pi577  & ~pi578 ;
  assign n9694 = ~n9692 & ~n9693;
  assign n9695 = pi579  & ~n9694;
  assign n9696 = ~n9691 & ~n9695;
  assign n9697 = ~n9690 & n9696;
  assign n9698 = n9690 & ~n9696;
  assign n9699 = ~n9697 & ~n9698;
  assign n9700 = ~pi579  & ~n9694;
  assign n9701 = pi579  & n9694;
  assign n9702 = ~n9700 & ~n9701;
  assign n9703 = ~pi582  & ~n9688;
  assign n9704 = pi582  & n9688;
  assign n9705 = ~n9703 & ~n9704;
  assign n9706 = ~n9702 & ~n9705;
  assign n9707 = ~n9699 & n9706;
  assign n9708 = ~n9690 & ~n9696;
  assign n9709 = ~n9707 & ~n9708;
  assign n9710 = n9699 & n9706;
  assign n9711 = ~n9699 & ~n9706;
  assign n9712 = ~n9710 & ~n9711;
  assign n9713 = n9674 & n9681;
  assign n9714 = ~n9674 & ~n9681;
  assign n9715 = ~n9713 & ~n9714;
  assign n9716 = ~n9684 & ~n9715;
  assign n9717 = ~n9709 & ~n9712;
  assign n9718 = ~n9702 & n9705;
  assign n9719 = n9702 & ~n9705;
  assign n9720 = ~n9718 & ~n9719;
  assign n9721 = ~n9677 & n9680;
  assign n9722 = n9677 & ~n9680;
  assign n9723 = ~n9721 & ~n9722;
  assign n9724 = ~n9720 & ~n9723;
  assign n9725 = ~n9716 & n9724;
  assign n9726 = ~n9717 & n9725;
  assign n9727 = n9712 & ~n9726;
  assign n9728 = ~n9712 & n9726;
  assign n9729 = ~n9727 & ~n9728;
  assign n9730 = n9715 & n9729;
  assign n9731 = ~n9727 & ~n9730;
  assign n9732 = n9709 & ~n9731;
  assign n9733 = ~n9684 & ~n9732;
  assign n9734 = ~n9709 & n9731;
  assign n9735 = ~n9733 & ~n9734;
  assign n9736 = pi562  & pi563 ;
  assign n9737 = ~pi562  & pi563 ;
  assign n9738 = pi562  & ~pi563 ;
  assign n9739 = ~n9737 & ~n9738;
  assign n9740 = pi564  & ~n9739;
  assign n9741 = ~n9736 & ~n9740;
  assign n9742 = pi559  & pi560 ;
  assign n9743 = ~pi559  & pi560 ;
  assign n9744 = pi559  & ~pi560 ;
  assign n9745 = ~n9743 & ~n9744;
  assign n9746 = pi561  & ~n9745;
  assign n9747 = ~n9742 & ~n9746;
  assign n9748 = ~n9741 & n9747;
  assign n9749 = n9741 & ~n9747;
  assign n9750 = ~n9748 & ~n9749;
  assign n9751 = ~pi561  & ~n9745;
  assign n9752 = pi561  & n9745;
  assign n9753 = ~n9751 & ~n9752;
  assign n9754 = ~pi564  & ~n9739;
  assign n9755 = pi564  & n9739;
  assign n9756 = ~n9754 & ~n9755;
  assign n9757 = ~n9753 & ~n9756;
  assign n9758 = ~n9750 & n9757;
  assign n9759 = ~n9741 & ~n9747;
  assign n9760 = ~n9758 & ~n9759;
  assign n9761 = pi568  & pi569 ;
  assign n9762 = ~pi568  & pi569 ;
  assign n9763 = pi568  & ~pi569 ;
  assign n9764 = ~n9762 & ~n9763;
  assign n9765 = pi570  & ~n9764;
  assign n9766 = ~n9761 & ~n9765;
  assign n9767 = pi565  & pi566 ;
  assign n9768 = ~pi565  & pi566 ;
  assign n9769 = pi565  & ~pi566 ;
  assign n9770 = ~n9768 & ~n9769;
  assign n9771 = pi567  & ~n9770;
  assign n9772 = ~n9767 & ~n9771;
  assign n9773 = ~n9766 & n9772;
  assign n9774 = n9766 & ~n9772;
  assign n9775 = ~n9773 & ~n9774;
  assign n9776 = ~pi567  & ~n9770;
  assign n9777 = pi567  & n9770;
  assign n9778 = ~n9776 & ~n9777;
  assign n9779 = ~pi570  & ~n9764;
  assign n9780 = pi570  & n9764;
  assign n9781 = ~n9779 & ~n9780;
  assign n9782 = ~n9778 & ~n9781;
  assign n9783 = ~n9775 & n9782;
  assign n9784 = ~n9766 & ~n9772;
  assign n9785 = ~n9783 & ~n9784;
  assign n9786 = n9775 & n9782;
  assign n9787 = ~n9775 & ~n9782;
  assign n9788 = ~n9786 & ~n9787;
  assign n9789 = n9750 & n9757;
  assign n9790 = ~n9750 & ~n9757;
  assign n9791 = ~n9789 & ~n9790;
  assign n9792 = ~n9760 & ~n9791;
  assign n9793 = ~n9785 & ~n9788;
  assign n9794 = ~n9778 & n9781;
  assign n9795 = n9778 & ~n9781;
  assign n9796 = ~n9794 & ~n9795;
  assign n9797 = ~n9753 & n9756;
  assign n9798 = n9753 & ~n9756;
  assign n9799 = ~n9797 & ~n9798;
  assign n9800 = ~n9796 & ~n9799;
  assign n9801 = ~n9792 & n9800;
  assign n9802 = ~n9793 & n9801;
  assign n9803 = n9788 & ~n9802;
  assign n9804 = ~n9788 & n9802;
  assign n9805 = ~n9803 & ~n9804;
  assign n9806 = n9791 & n9805;
  assign n9807 = ~n9803 & ~n9806;
  assign n9808 = n9785 & ~n9807;
  assign n9809 = ~n9760 & ~n9808;
  assign n9810 = ~n9785 & n9807;
  assign n9811 = ~n9809 & ~n9810;
  assign n9812 = n9735 & n9811;
  assign n9813 = ~n9760 & n9785;
  assign n9814 = n9760 & ~n9785;
  assign n9815 = ~n9813 & ~n9814;
  assign n9816 = n9807 & ~n9815;
  assign n9817 = ~n9807 & n9815;
  assign n9818 = ~n9816 & ~n9817;
  assign n9819 = ~n9684 & n9709;
  assign n9820 = n9684 & ~n9709;
  assign n9821 = ~n9819 & ~n9820;
  assign n9822 = n9731 & ~n9821;
  assign n9823 = ~n9731 & n9821;
  assign n9824 = ~n9822 & ~n9823;
  assign n9825 = n9818 & n9824;
  assign n9826 = n9720 & ~n9723;
  assign n9827 = ~n9720 & n9723;
  assign n9828 = ~n9826 & ~n9827;
  assign n9829 = n9796 & ~n9799;
  assign n9830 = ~n9796 & n9799;
  assign n9831 = ~n9829 & ~n9830;
  assign n9832 = ~n9828 & ~n9831;
  assign n9833 = ~n9715 & ~n9729;
  assign n9834 = ~n9730 & ~n9833;
  assign n9835 = ~n9832 & n9834;
  assign n9836 = ~n9791 & ~n9805;
  assign n9837 = ~n9806 & ~n9836;
  assign n9838 = n9832 & ~n9834;
  assign n9839 = ~n9835 & ~n9838;
  assign n9840 = n9837 & n9839;
  assign n9841 = ~n9835 & ~n9840;
  assign n9842 = ~n9818 & ~n9824;
  assign n9843 = ~n9825 & ~n9842;
  assign n9844 = n9841 & n9843;
  assign n9845 = ~n9825 & ~n9844;
  assign n9846 = ~n9812 & ~n9845;
  assign n9847 = ~n9735 & ~n9811;
  assign n9848 = ~n9846 & ~n9847;
  assign n9849 = ~n9659 & ~n9848;
  assign n9850 = n9659 & n9848;
  assign n9851 = ~n9849 & ~n9850;
  assign n9852 = ~n9622 & ~n9658;
  assign n9853 = ~n9656 & n9852;
  assign n9854 = n9656 & ~n9852;
  assign n9855 = ~n9853 & ~n9854;
  assign n9856 = ~n9812 & ~n9847;
  assign n9857 = ~n9845 & n9856;
  assign n9858 = n9845 & ~n9856;
  assign n9859 = ~n9857 & ~n9858;
  assign n9860 = n9855 & n9859;
  assign n9861 = ~n9841 & ~n9843;
  assign n9862 = ~n9844 & ~n9861;
  assign n9863 = ~n9652 & ~n9654;
  assign n9864 = ~n9655 & ~n9863;
  assign n9865 = n9862 & n9864;
  assign n9866 = ~n9862 & ~n9864;
  assign n9867 = ~n9865 & ~n9866;
  assign n9868 = ~n9638 & n9641;
  assign n9869 = n9638 & ~n9641;
  assign n9870 = ~n9868 & ~n9869;
  assign n9871 = ~n9828 & n9831;
  assign n9872 = n9828 & ~n9831;
  assign n9873 = ~n9871 & ~n9872;
  assign n9874 = ~n9870 & ~n9873;
  assign n9875 = ~n9647 & n9650;
  assign n9876 = ~n9651 & ~n9875;
  assign n9877 = ~n9874 & n9876;
  assign n9878 = ~n9837 & ~n9839;
  assign n9879 = ~n9840 & ~n9878;
  assign n9880 = n9874 & ~n9876;
  assign n9881 = ~n9877 & ~n9880;
  assign n9882 = n9879 & n9881;
  assign n9883 = ~n9877 & ~n9882;
  assign n9884 = n9867 & n9883;
  assign n9885 = ~n9865 & ~n9884;
  assign n9886 = ~n9855 & ~n9859;
  assign n9887 = ~n9860 & ~n9886;
  assign n9888 = ~n9885 & n9887;
  assign n9889 = ~n9860 & ~n9888;
  assign n9890 = n9851 & ~n9889;
  assign n9891 = ~n9849 & ~n9890;
  assign n9892 = ~n9469 & ~n9891;
  assign n9893 = ~n9851 & n9889;
  assign n9894 = ~n9890 & ~n9893;
  assign n9895 = ~n9429 & n9467;
  assign n9896 = ~n9468 & ~n9895;
  assign n9897 = n9894 & n9896;
  assign n9898 = n9463 & ~n9465;
  assign n9899 = ~n9466 & ~n9898;
  assign n9900 = n9885 & ~n9887;
  assign n9901 = ~n9888 & ~n9900;
  assign n9902 = n9899 & n9901;
  assign n9903 = ~n9899 & ~n9901;
  assign n9904 = ~n9902 & ~n9903;
  assign n9905 = ~n9867 & ~n9883;
  assign n9906 = ~n9884 & ~n9905;
  assign n9907 = ~n9445 & ~n9461;
  assign n9908 = ~n9462 & ~n9907;
  assign n9909 = n9906 & n9908;
  assign n9910 = ~n9906 & ~n9908;
  assign n9911 = ~n9909 & ~n9910;
  assign n9912 = ~n9448 & n9451;
  assign n9913 = n9448 & ~n9451;
  assign n9914 = ~n9912 & ~n9913;
  assign n9915 = ~n9870 & n9873;
  assign n9916 = n9870 & ~n9873;
  assign n9917 = ~n9915 & ~n9916;
  assign n9918 = ~n9914 & ~n9917;
  assign n9919 = ~n9457 & ~n9459;
  assign n9920 = ~n9460 & ~n9919;
  assign n9921 = ~n9918 & n9920;
  assign n9922 = ~n9879 & ~n9881;
  assign n9923 = ~n9882 & ~n9922;
  assign n9924 = n9918 & ~n9920;
  assign n9925 = ~n9921 & ~n9924;
  assign n9926 = n9923 & n9925;
  assign n9927 = ~n9921 & ~n9926;
  assign n9928 = n9911 & n9927;
  assign n9929 = ~n9909 & ~n9928;
  assign n9930 = n9904 & ~n9929;
  assign n9931 = ~n9902 & ~n9930;
  assign n9932 = ~n9894 & ~n9896;
  assign n9933 = ~n9897 & ~n9932;
  assign n9934 = ~n9931 & n9933;
  assign n9935 = ~n9897 & ~n9934;
  assign n9936 = n9469 & n9891;
  assign n9937 = ~n9892 & ~n9936;
  assign n9938 = ~n9935 & n9937;
  assign n9939 = ~n9892 & ~n9938;
  assign n9940 = pi550  & pi551 ;
  assign n9941 = ~pi550  & pi551 ;
  assign n9942 = pi550  & ~pi551 ;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = pi552  & ~n9943;
  assign n9945 = ~n9940 & ~n9944;
  assign n9946 = pi547  & pi548 ;
  assign n9947 = ~pi547  & pi548 ;
  assign n9948 = pi547  & ~pi548 ;
  assign n9949 = ~n9947 & ~n9948;
  assign n9950 = pi549  & ~n9949;
  assign n9951 = ~n9946 & ~n9950;
  assign n9952 = ~n9945 & n9951;
  assign n9953 = n9945 & ~n9951;
  assign n9954 = ~n9952 & ~n9953;
  assign n9955 = ~pi549  & ~n9949;
  assign n9956 = pi549  & n9949;
  assign n9957 = ~n9955 & ~n9956;
  assign n9958 = ~pi552  & ~n9943;
  assign n9959 = pi552  & n9943;
  assign n9960 = ~n9958 & ~n9959;
  assign n9961 = ~n9957 & ~n9960;
  assign n9962 = ~n9954 & n9961;
  assign n9963 = ~n9945 & ~n9951;
  assign n9964 = ~n9962 & ~n9963;
  assign n9965 = pi556  & pi557 ;
  assign n9966 = ~pi556  & pi557 ;
  assign n9967 = pi556  & ~pi557 ;
  assign n9968 = ~n9966 & ~n9967;
  assign n9969 = pi558  & ~n9968;
  assign n9970 = ~n9965 & ~n9969;
  assign n9971 = pi553  & pi554 ;
  assign n9972 = ~pi553  & pi554 ;
  assign n9973 = pi553  & ~pi554 ;
  assign n9974 = ~n9972 & ~n9973;
  assign n9975 = pi555  & ~n9974;
  assign n9976 = ~n9971 & ~n9975;
  assign n9977 = ~n9970 & n9976;
  assign n9978 = n9970 & ~n9976;
  assign n9979 = ~n9977 & ~n9978;
  assign n9980 = ~pi555  & ~n9974;
  assign n9981 = pi555  & n9974;
  assign n9982 = ~n9980 & ~n9981;
  assign n9983 = ~pi558  & ~n9968;
  assign n9984 = pi558  & n9968;
  assign n9985 = ~n9983 & ~n9984;
  assign n9986 = ~n9982 & ~n9985;
  assign n9987 = ~n9979 & n9986;
  assign n9988 = ~n9970 & ~n9976;
  assign n9989 = ~n9987 & ~n9988;
  assign n9990 = n9979 & n9986;
  assign n9991 = ~n9979 & ~n9986;
  assign n9992 = ~n9990 & ~n9991;
  assign n9993 = n9954 & n9961;
  assign n9994 = ~n9954 & ~n9961;
  assign n9995 = ~n9993 & ~n9994;
  assign n9996 = ~n9964 & ~n9995;
  assign n9997 = ~n9989 & ~n9992;
  assign n9998 = ~n9982 & n9985;
  assign n9999 = n9982 & ~n9985;
  assign n10000 = ~n9998 & ~n9999;
  assign n10001 = ~n9957 & n9960;
  assign n10002 = n9957 & ~n9960;
  assign n10003 = ~n10001 & ~n10002;
  assign n10004 = ~n10000 & ~n10003;
  assign n10005 = ~n9996 & n10004;
  assign n10006 = ~n9997 & n10005;
  assign n10007 = n9992 & ~n10006;
  assign n10008 = ~n9992 & n10006;
  assign n10009 = ~n10007 & ~n10008;
  assign n10010 = n9995 & n10009;
  assign n10011 = ~n10007 & ~n10010;
  assign n10012 = n9989 & ~n10011;
  assign n10013 = ~n9964 & ~n10012;
  assign n10014 = ~n9989 & n10011;
  assign n10015 = ~n10013 & ~n10014;
  assign n10016 = pi538  & pi539 ;
  assign n10017 = ~pi538  & pi539 ;
  assign n10018 = pi538  & ~pi539 ;
  assign n10019 = ~n10017 & ~n10018;
  assign n10020 = pi540  & ~n10019;
  assign n10021 = ~n10016 & ~n10020;
  assign n10022 = pi535  & pi536 ;
  assign n10023 = ~pi535  & pi536 ;
  assign n10024 = pi535  & ~pi536 ;
  assign n10025 = ~n10023 & ~n10024;
  assign n10026 = pi537  & ~n10025;
  assign n10027 = ~n10022 & ~n10026;
  assign n10028 = ~n10021 & n10027;
  assign n10029 = n10021 & ~n10027;
  assign n10030 = ~n10028 & ~n10029;
  assign n10031 = ~pi537  & ~n10025;
  assign n10032 = pi537  & n10025;
  assign n10033 = ~n10031 & ~n10032;
  assign n10034 = ~pi540  & ~n10019;
  assign n10035 = pi540  & n10019;
  assign n10036 = ~n10034 & ~n10035;
  assign n10037 = ~n10033 & ~n10036;
  assign n10038 = ~n10030 & n10037;
  assign n10039 = ~n10021 & ~n10027;
  assign n10040 = ~n10038 & ~n10039;
  assign n10041 = pi544  & pi545 ;
  assign n10042 = ~pi544  & pi545 ;
  assign n10043 = pi544  & ~pi545 ;
  assign n10044 = ~n10042 & ~n10043;
  assign n10045 = pi546  & ~n10044;
  assign n10046 = ~n10041 & ~n10045;
  assign n10047 = pi541  & pi542 ;
  assign n10048 = ~pi541  & pi542 ;
  assign n10049 = pi541  & ~pi542 ;
  assign n10050 = ~n10048 & ~n10049;
  assign n10051 = pi543  & ~n10050;
  assign n10052 = ~n10047 & ~n10051;
  assign n10053 = ~n10046 & n10052;
  assign n10054 = n10046 & ~n10052;
  assign n10055 = ~n10053 & ~n10054;
  assign n10056 = ~pi543  & ~n10050;
  assign n10057 = pi543  & n10050;
  assign n10058 = ~n10056 & ~n10057;
  assign n10059 = ~pi546  & ~n10044;
  assign n10060 = pi546  & n10044;
  assign n10061 = ~n10059 & ~n10060;
  assign n10062 = ~n10058 & ~n10061;
  assign n10063 = ~n10055 & n10062;
  assign n10064 = ~n10046 & ~n10052;
  assign n10065 = ~n10063 & ~n10064;
  assign n10066 = n10055 & n10062;
  assign n10067 = ~n10055 & ~n10062;
  assign n10068 = ~n10066 & ~n10067;
  assign n10069 = n10030 & n10037;
  assign n10070 = ~n10030 & ~n10037;
  assign n10071 = ~n10069 & ~n10070;
  assign n10072 = ~n10040 & ~n10071;
  assign n10073 = ~n10065 & ~n10068;
  assign n10074 = ~n10058 & n10061;
  assign n10075 = n10058 & ~n10061;
  assign n10076 = ~n10074 & ~n10075;
  assign n10077 = ~n10033 & n10036;
  assign n10078 = n10033 & ~n10036;
  assign n10079 = ~n10077 & ~n10078;
  assign n10080 = ~n10076 & ~n10079;
  assign n10081 = ~n10072 & n10080;
  assign n10082 = ~n10073 & n10081;
  assign n10083 = n10068 & ~n10082;
  assign n10084 = ~n10068 & n10082;
  assign n10085 = ~n10083 & ~n10084;
  assign n10086 = n10071 & n10085;
  assign n10087 = ~n10083 & ~n10086;
  assign n10088 = n10065 & ~n10087;
  assign n10089 = ~n10040 & ~n10088;
  assign n10090 = ~n10065 & n10087;
  assign n10091 = ~n10089 & ~n10090;
  assign n10092 = n10015 & n10091;
  assign n10093 = ~n10040 & n10065;
  assign n10094 = n10040 & ~n10065;
  assign n10095 = ~n10093 & ~n10094;
  assign n10096 = n10087 & ~n10095;
  assign n10097 = ~n10087 & n10095;
  assign n10098 = ~n10096 & ~n10097;
  assign n10099 = ~n9964 & n9989;
  assign n10100 = n9964 & ~n9989;
  assign n10101 = ~n10099 & ~n10100;
  assign n10102 = n10011 & ~n10101;
  assign n10103 = ~n10011 & n10101;
  assign n10104 = ~n10102 & ~n10103;
  assign n10105 = n10098 & n10104;
  assign n10106 = n10000 & ~n10003;
  assign n10107 = ~n10000 & n10003;
  assign n10108 = ~n10106 & ~n10107;
  assign n10109 = n10076 & ~n10079;
  assign n10110 = ~n10076 & n10079;
  assign n10111 = ~n10109 & ~n10110;
  assign n10112 = ~n10108 & ~n10111;
  assign n10113 = ~n9995 & ~n10009;
  assign n10114 = ~n10010 & ~n10113;
  assign n10115 = ~n10112 & n10114;
  assign n10116 = ~n10071 & ~n10085;
  assign n10117 = ~n10086 & ~n10116;
  assign n10118 = ~n10112 & ~n10114;
  assign n10119 = n10114 & ~n10115;
  assign n10120 = ~n10118 & ~n10119;
  assign n10121 = n10117 & ~n10120;
  assign n10122 = ~n10115 & ~n10121;
  assign n10123 = ~n10098 & ~n10104;
  assign n10124 = ~n10105 & ~n10123;
  assign n10125 = n10122 & n10124;
  assign n10126 = ~n10105 & ~n10125;
  assign n10127 = ~n10092 & ~n10126;
  assign n10128 = ~n10015 & ~n10091;
  assign n10129 = ~n10127 & ~n10128;
  assign n10130 = pi526  & pi527 ;
  assign n10131 = ~pi526  & pi527 ;
  assign n10132 = pi526  & ~pi527 ;
  assign n10133 = ~n10131 & ~n10132;
  assign n10134 = pi528  & ~n10133;
  assign n10135 = ~n10130 & ~n10134;
  assign n10136 = pi523  & pi524 ;
  assign n10137 = ~pi523  & pi524 ;
  assign n10138 = pi523  & ~pi524 ;
  assign n10139 = ~n10137 & ~n10138;
  assign n10140 = pi525  & ~n10139;
  assign n10141 = ~n10136 & ~n10140;
  assign n10142 = ~n10135 & n10141;
  assign n10143 = n10135 & ~n10141;
  assign n10144 = ~n10142 & ~n10143;
  assign n10145 = ~pi525  & ~n10139;
  assign n10146 = pi525  & n10139;
  assign n10147 = ~n10145 & ~n10146;
  assign n10148 = ~pi528  & ~n10133;
  assign n10149 = pi528  & n10133;
  assign n10150 = ~n10148 & ~n10149;
  assign n10151 = ~n10147 & ~n10150;
  assign n10152 = ~n10144 & n10151;
  assign n10153 = ~n10135 & ~n10141;
  assign n10154 = ~n10152 & ~n10153;
  assign n10155 = pi532  & pi533 ;
  assign n10156 = ~pi532  & pi533 ;
  assign n10157 = pi532  & ~pi533 ;
  assign n10158 = ~n10156 & ~n10157;
  assign n10159 = pi534  & ~n10158;
  assign n10160 = ~n10155 & ~n10159;
  assign n10161 = pi529  & pi530 ;
  assign n10162 = ~pi529  & pi530 ;
  assign n10163 = pi529  & ~pi530 ;
  assign n10164 = ~n10162 & ~n10163;
  assign n10165 = pi531  & ~n10164;
  assign n10166 = ~n10161 & ~n10165;
  assign n10167 = ~n10160 & n10166;
  assign n10168 = n10160 & ~n10166;
  assign n10169 = ~n10167 & ~n10168;
  assign n10170 = ~pi531  & ~n10164;
  assign n10171 = pi531  & n10164;
  assign n10172 = ~n10170 & ~n10171;
  assign n10173 = ~pi534  & ~n10158;
  assign n10174 = pi534  & n10158;
  assign n10175 = ~n10173 & ~n10174;
  assign n10176 = ~n10172 & ~n10175;
  assign n10177 = ~n10169 & n10176;
  assign n10178 = ~n10160 & ~n10166;
  assign n10179 = ~n10177 & ~n10178;
  assign n10180 = n10169 & n10176;
  assign n10181 = ~n10169 & ~n10176;
  assign n10182 = ~n10180 & ~n10181;
  assign n10183 = n10144 & n10151;
  assign n10184 = ~n10144 & ~n10151;
  assign n10185 = ~n10183 & ~n10184;
  assign n10186 = ~n10154 & ~n10185;
  assign n10187 = ~n10179 & ~n10182;
  assign n10188 = ~n10172 & n10175;
  assign n10189 = n10172 & ~n10175;
  assign n10190 = ~n10188 & ~n10189;
  assign n10191 = ~n10147 & n10150;
  assign n10192 = n10147 & ~n10150;
  assign n10193 = ~n10191 & ~n10192;
  assign n10194 = ~n10190 & ~n10193;
  assign n10195 = ~n10186 & n10194;
  assign n10196 = ~n10187 & n10195;
  assign n10197 = n10182 & ~n10196;
  assign n10198 = ~n10182 & n10196;
  assign n10199 = ~n10197 & ~n10198;
  assign n10200 = n10185 & n10199;
  assign n10201 = ~n10197 & ~n10200;
  assign n10202 = n10179 & ~n10201;
  assign n10203 = ~n10154 & ~n10202;
  assign n10204 = ~n10179 & n10201;
  assign n10205 = ~n10203 & ~n10204;
  assign n10206 = pi514  & pi515 ;
  assign n10207 = ~pi514  & pi515 ;
  assign n10208 = pi514  & ~pi515 ;
  assign n10209 = ~n10207 & ~n10208;
  assign n10210 = pi516  & ~n10209;
  assign n10211 = ~n10206 & ~n10210;
  assign n10212 = pi511  & pi512 ;
  assign n10213 = ~pi511  & pi512 ;
  assign n10214 = pi511  & ~pi512 ;
  assign n10215 = ~n10213 & ~n10214;
  assign n10216 = pi513  & ~n10215;
  assign n10217 = ~n10212 & ~n10216;
  assign n10218 = ~n10211 & n10217;
  assign n10219 = n10211 & ~n10217;
  assign n10220 = ~n10218 & ~n10219;
  assign n10221 = ~pi513  & ~n10215;
  assign n10222 = pi513  & n10215;
  assign n10223 = ~n10221 & ~n10222;
  assign n10224 = ~pi516  & ~n10209;
  assign n10225 = pi516  & n10209;
  assign n10226 = ~n10224 & ~n10225;
  assign n10227 = ~n10223 & ~n10226;
  assign n10228 = ~n10220 & n10227;
  assign n10229 = ~n10211 & ~n10217;
  assign n10230 = ~n10228 & ~n10229;
  assign n10231 = pi520  & pi521 ;
  assign n10232 = ~pi520  & pi521 ;
  assign n10233 = pi520  & ~pi521 ;
  assign n10234 = ~n10232 & ~n10233;
  assign n10235 = pi522  & ~n10234;
  assign n10236 = ~n10231 & ~n10235;
  assign n10237 = pi517  & pi518 ;
  assign n10238 = ~pi517  & pi518 ;
  assign n10239 = pi517  & ~pi518 ;
  assign n10240 = ~n10238 & ~n10239;
  assign n10241 = pi519  & ~n10240;
  assign n10242 = ~n10237 & ~n10241;
  assign n10243 = ~n10236 & n10242;
  assign n10244 = n10236 & ~n10242;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = ~pi519  & ~n10240;
  assign n10247 = pi519  & n10240;
  assign n10248 = ~n10246 & ~n10247;
  assign n10249 = ~pi522  & ~n10234;
  assign n10250 = pi522  & n10234;
  assign n10251 = ~n10249 & ~n10250;
  assign n10252 = ~n10248 & ~n10251;
  assign n10253 = ~n10245 & n10252;
  assign n10254 = ~n10236 & ~n10242;
  assign n10255 = ~n10253 & ~n10254;
  assign n10256 = n10245 & n10252;
  assign n10257 = ~n10245 & ~n10252;
  assign n10258 = ~n10256 & ~n10257;
  assign n10259 = n10220 & n10227;
  assign n10260 = ~n10220 & ~n10227;
  assign n10261 = ~n10259 & ~n10260;
  assign n10262 = ~n10230 & ~n10261;
  assign n10263 = ~n10255 & ~n10258;
  assign n10264 = ~n10248 & n10251;
  assign n10265 = n10248 & ~n10251;
  assign n10266 = ~n10264 & ~n10265;
  assign n10267 = ~n10223 & n10226;
  assign n10268 = n10223 & ~n10226;
  assign n10269 = ~n10267 & ~n10268;
  assign n10270 = ~n10266 & ~n10269;
  assign n10271 = ~n10262 & n10270;
  assign n10272 = ~n10263 & n10271;
  assign n10273 = n10258 & ~n10272;
  assign n10274 = ~n10258 & n10272;
  assign n10275 = ~n10273 & ~n10274;
  assign n10276 = n10261 & n10275;
  assign n10277 = ~n10273 & ~n10276;
  assign n10278 = n10255 & ~n10277;
  assign n10279 = ~n10230 & ~n10278;
  assign n10280 = ~n10255 & n10277;
  assign n10281 = ~n10279 & ~n10280;
  assign n10282 = n10205 & n10281;
  assign n10283 = ~n10230 & n10255;
  assign n10284 = n10230 & ~n10255;
  assign n10285 = ~n10283 & ~n10284;
  assign n10286 = n10277 & ~n10285;
  assign n10287 = ~n10277 & n10285;
  assign n10288 = ~n10286 & ~n10287;
  assign n10289 = ~n10154 & n10179;
  assign n10290 = n10154 & ~n10179;
  assign n10291 = ~n10289 & ~n10290;
  assign n10292 = n10201 & ~n10291;
  assign n10293 = ~n10201 & n10291;
  assign n10294 = ~n10292 & ~n10293;
  assign n10295 = n10288 & n10294;
  assign n10296 = n10190 & ~n10193;
  assign n10297 = ~n10190 & n10193;
  assign n10298 = ~n10296 & ~n10297;
  assign n10299 = n10266 & ~n10269;
  assign n10300 = ~n10266 & n10269;
  assign n10301 = ~n10299 & ~n10300;
  assign n10302 = ~n10298 & ~n10301;
  assign n10303 = ~n10185 & ~n10199;
  assign n10304 = ~n10200 & ~n10303;
  assign n10305 = ~n10302 & n10304;
  assign n10306 = ~n10261 & ~n10275;
  assign n10307 = ~n10276 & ~n10306;
  assign n10308 = n10302 & ~n10304;
  assign n10309 = ~n10305 & ~n10308;
  assign n10310 = n10307 & n10309;
  assign n10311 = ~n10305 & ~n10310;
  assign n10312 = ~n10288 & ~n10294;
  assign n10313 = ~n10295 & ~n10312;
  assign n10314 = n10311 & n10313;
  assign n10315 = ~n10295 & ~n10314;
  assign n10316 = ~n10282 & ~n10315;
  assign n10317 = ~n10205 & ~n10281;
  assign n10318 = ~n10316 & ~n10317;
  assign n10319 = ~n10129 & ~n10318;
  assign n10320 = n10129 & n10318;
  assign n10321 = ~n10319 & ~n10320;
  assign n10322 = ~n10092 & ~n10128;
  assign n10323 = ~n10126 & n10322;
  assign n10324 = n10126 & ~n10322;
  assign n10325 = ~n10323 & ~n10324;
  assign n10326 = ~n10282 & ~n10317;
  assign n10327 = ~n10315 & n10326;
  assign n10328 = n10315 & ~n10326;
  assign n10329 = ~n10327 & ~n10328;
  assign n10330 = n10325 & n10329;
  assign n10331 = ~n10311 & ~n10313;
  assign n10332 = ~n10314 & ~n10331;
  assign n10333 = ~n10122 & ~n10124;
  assign n10334 = ~n10125 & ~n10333;
  assign n10335 = n10332 & n10334;
  assign n10336 = ~n10332 & ~n10334;
  assign n10337 = ~n10335 & ~n10336;
  assign n10338 = ~n10108 & n10111;
  assign n10339 = n10108 & ~n10111;
  assign n10340 = ~n10338 & ~n10339;
  assign n10341 = ~n10298 & n10301;
  assign n10342 = n10298 & ~n10301;
  assign n10343 = ~n10341 & ~n10342;
  assign n10344 = ~n10340 & ~n10343;
  assign n10345 = ~n10117 & n10120;
  assign n10346 = ~n10121 & ~n10345;
  assign n10347 = ~n10344 & n10346;
  assign n10348 = ~n10307 & ~n10309;
  assign n10349 = ~n10310 & ~n10348;
  assign n10350 = n10344 & ~n10346;
  assign n10351 = ~n10347 & ~n10350;
  assign n10352 = n10349 & n10351;
  assign n10353 = ~n10347 & ~n10352;
  assign n10354 = n10337 & n10353;
  assign n10355 = ~n10335 & ~n10354;
  assign n10356 = ~n10325 & ~n10329;
  assign n10357 = ~n10330 & ~n10356;
  assign n10358 = ~n10355 & n10357;
  assign n10359 = ~n10330 & ~n10358;
  assign n10360 = n10321 & ~n10359;
  assign n10361 = ~n10319 & ~n10360;
  assign n10362 = pi502  & pi503 ;
  assign n10363 = ~pi502  & pi503 ;
  assign n10364 = pi502  & ~pi503 ;
  assign n10365 = ~n10363 & ~n10364;
  assign n10366 = pi504  & ~n10365;
  assign n10367 = ~n10362 & ~n10366;
  assign n10368 = pi499  & pi500 ;
  assign n10369 = ~pi499  & pi500 ;
  assign n10370 = pi499  & ~pi500 ;
  assign n10371 = ~n10369 & ~n10370;
  assign n10372 = pi501  & ~n10371;
  assign n10373 = ~n10368 & ~n10372;
  assign n10374 = ~n10367 & n10373;
  assign n10375 = n10367 & ~n10373;
  assign n10376 = ~n10374 & ~n10375;
  assign n10377 = ~pi501  & ~n10371;
  assign n10378 = pi501  & n10371;
  assign n10379 = ~n10377 & ~n10378;
  assign n10380 = ~pi504  & ~n10365;
  assign n10381 = pi504  & n10365;
  assign n10382 = ~n10380 & ~n10381;
  assign n10383 = ~n10379 & ~n10382;
  assign n10384 = ~n10376 & n10383;
  assign n10385 = ~n10367 & ~n10373;
  assign n10386 = ~n10384 & ~n10385;
  assign n10387 = pi508  & pi509 ;
  assign n10388 = ~pi508  & pi509 ;
  assign n10389 = pi508  & ~pi509 ;
  assign n10390 = ~n10388 & ~n10389;
  assign n10391 = pi510  & ~n10390;
  assign n10392 = ~n10387 & ~n10391;
  assign n10393 = pi505  & pi506 ;
  assign n10394 = ~pi505  & pi506 ;
  assign n10395 = pi505  & ~pi506 ;
  assign n10396 = ~n10394 & ~n10395;
  assign n10397 = pi507  & ~n10396;
  assign n10398 = ~n10393 & ~n10397;
  assign n10399 = ~n10392 & n10398;
  assign n10400 = n10392 & ~n10398;
  assign n10401 = ~n10399 & ~n10400;
  assign n10402 = ~pi507  & ~n10396;
  assign n10403 = pi507  & n10396;
  assign n10404 = ~n10402 & ~n10403;
  assign n10405 = ~pi510  & ~n10390;
  assign n10406 = pi510  & n10390;
  assign n10407 = ~n10405 & ~n10406;
  assign n10408 = ~n10404 & ~n10407;
  assign n10409 = ~n10401 & n10408;
  assign n10410 = ~n10392 & ~n10398;
  assign n10411 = ~n10409 & ~n10410;
  assign n10412 = n10401 & n10408;
  assign n10413 = ~n10401 & ~n10408;
  assign n10414 = ~n10412 & ~n10413;
  assign n10415 = n10376 & n10383;
  assign n10416 = ~n10376 & ~n10383;
  assign n10417 = ~n10415 & ~n10416;
  assign n10418 = ~n10386 & ~n10417;
  assign n10419 = ~n10411 & ~n10414;
  assign n10420 = ~n10404 & n10407;
  assign n10421 = n10404 & ~n10407;
  assign n10422 = ~n10420 & ~n10421;
  assign n10423 = ~n10379 & n10382;
  assign n10424 = n10379 & ~n10382;
  assign n10425 = ~n10423 & ~n10424;
  assign n10426 = ~n10422 & ~n10425;
  assign n10427 = ~n10418 & n10426;
  assign n10428 = ~n10419 & n10427;
  assign n10429 = n10414 & ~n10428;
  assign n10430 = ~n10414 & n10428;
  assign n10431 = ~n10429 & ~n10430;
  assign n10432 = n10417 & n10431;
  assign n10433 = ~n10429 & ~n10432;
  assign n10434 = n10411 & ~n10433;
  assign n10435 = ~n10386 & ~n10434;
  assign n10436 = ~n10411 & n10433;
  assign n10437 = ~n10435 & ~n10436;
  assign n10438 = pi490  & pi491 ;
  assign n10439 = ~pi490  & pi491 ;
  assign n10440 = pi490  & ~pi491 ;
  assign n10441 = ~n10439 & ~n10440;
  assign n10442 = pi492  & ~n10441;
  assign n10443 = ~n10438 & ~n10442;
  assign n10444 = pi487  & pi488 ;
  assign n10445 = ~pi487  & pi488 ;
  assign n10446 = pi487  & ~pi488 ;
  assign n10447 = ~n10445 & ~n10446;
  assign n10448 = pi489  & ~n10447;
  assign n10449 = ~n10444 & ~n10448;
  assign n10450 = ~n10443 & n10449;
  assign n10451 = n10443 & ~n10449;
  assign n10452 = ~n10450 & ~n10451;
  assign n10453 = ~pi489  & ~n10447;
  assign n10454 = pi489  & n10447;
  assign n10455 = ~n10453 & ~n10454;
  assign n10456 = ~pi492  & ~n10441;
  assign n10457 = pi492  & n10441;
  assign n10458 = ~n10456 & ~n10457;
  assign n10459 = ~n10455 & ~n10458;
  assign n10460 = ~n10452 & n10459;
  assign n10461 = ~n10443 & ~n10449;
  assign n10462 = ~n10460 & ~n10461;
  assign n10463 = pi496  & pi497 ;
  assign n10464 = ~pi496  & pi497 ;
  assign n10465 = pi496  & ~pi497 ;
  assign n10466 = ~n10464 & ~n10465;
  assign n10467 = pi498  & ~n10466;
  assign n10468 = ~n10463 & ~n10467;
  assign n10469 = pi493  & pi494 ;
  assign n10470 = ~pi493  & pi494 ;
  assign n10471 = pi493  & ~pi494 ;
  assign n10472 = ~n10470 & ~n10471;
  assign n10473 = pi495  & ~n10472;
  assign n10474 = ~n10469 & ~n10473;
  assign n10475 = ~n10468 & n10474;
  assign n10476 = n10468 & ~n10474;
  assign n10477 = ~n10475 & ~n10476;
  assign n10478 = ~pi495  & ~n10472;
  assign n10479 = pi495  & n10472;
  assign n10480 = ~n10478 & ~n10479;
  assign n10481 = ~pi498  & ~n10466;
  assign n10482 = pi498  & n10466;
  assign n10483 = ~n10481 & ~n10482;
  assign n10484 = ~n10480 & ~n10483;
  assign n10485 = ~n10477 & n10484;
  assign n10486 = ~n10468 & ~n10474;
  assign n10487 = ~n10485 & ~n10486;
  assign n10488 = n10477 & n10484;
  assign n10489 = ~n10477 & ~n10484;
  assign n10490 = ~n10488 & ~n10489;
  assign n10491 = n10452 & n10459;
  assign n10492 = ~n10452 & ~n10459;
  assign n10493 = ~n10491 & ~n10492;
  assign n10494 = ~n10462 & ~n10493;
  assign n10495 = ~n10487 & ~n10490;
  assign n10496 = ~n10480 & n10483;
  assign n10497 = n10480 & ~n10483;
  assign n10498 = ~n10496 & ~n10497;
  assign n10499 = ~n10455 & n10458;
  assign n10500 = n10455 & ~n10458;
  assign n10501 = ~n10499 & ~n10500;
  assign n10502 = ~n10498 & ~n10501;
  assign n10503 = ~n10494 & n10502;
  assign n10504 = ~n10495 & n10503;
  assign n10505 = n10490 & ~n10504;
  assign n10506 = ~n10490 & n10504;
  assign n10507 = ~n10505 & ~n10506;
  assign n10508 = n10493 & n10507;
  assign n10509 = ~n10505 & ~n10508;
  assign n10510 = n10487 & ~n10509;
  assign n10511 = ~n10462 & ~n10510;
  assign n10512 = ~n10487 & n10509;
  assign n10513 = ~n10511 & ~n10512;
  assign n10514 = n10437 & n10513;
  assign n10515 = ~n10462 & n10487;
  assign n10516 = n10462 & ~n10487;
  assign n10517 = ~n10515 & ~n10516;
  assign n10518 = n10509 & ~n10517;
  assign n10519 = ~n10509 & n10517;
  assign n10520 = ~n10518 & ~n10519;
  assign n10521 = ~n10386 & n10411;
  assign n10522 = n10386 & ~n10411;
  assign n10523 = ~n10521 & ~n10522;
  assign n10524 = n10433 & ~n10523;
  assign n10525 = ~n10433 & n10523;
  assign n10526 = ~n10524 & ~n10525;
  assign n10527 = n10520 & n10526;
  assign n10528 = n10422 & ~n10425;
  assign n10529 = ~n10422 & n10425;
  assign n10530 = ~n10528 & ~n10529;
  assign n10531 = n10498 & ~n10501;
  assign n10532 = ~n10498 & n10501;
  assign n10533 = ~n10531 & ~n10532;
  assign n10534 = ~n10530 & ~n10533;
  assign n10535 = ~n10417 & ~n10431;
  assign n10536 = ~n10432 & ~n10535;
  assign n10537 = ~n10534 & n10536;
  assign n10538 = ~n10493 & ~n10507;
  assign n10539 = ~n10508 & ~n10538;
  assign n10540 = ~n10534 & ~n10536;
  assign n10541 = n10536 & ~n10537;
  assign n10542 = ~n10540 & ~n10541;
  assign n10543 = n10539 & ~n10542;
  assign n10544 = ~n10537 & ~n10543;
  assign n10545 = ~n10520 & ~n10526;
  assign n10546 = ~n10527 & ~n10545;
  assign n10547 = n10544 & n10546;
  assign n10548 = ~n10527 & ~n10547;
  assign n10549 = ~n10514 & ~n10548;
  assign n10550 = ~n10437 & ~n10513;
  assign n10551 = ~n10549 & ~n10550;
  assign n10552 = pi478  & pi479 ;
  assign n10553 = ~pi478  & pi479 ;
  assign n10554 = pi478  & ~pi479 ;
  assign n10555 = ~n10553 & ~n10554;
  assign n10556 = pi480  & ~n10555;
  assign n10557 = ~n10552 & ~n10556;
  assign n10558 = pi475  & pi476 ;
  assign n10559 = ~pi475  & pi476 ;
  assign n10560 = pi475  & ~pi476 ;
  assign n10561 = ~n10559 & ~n10560;
  assign n10562 = pi477  & ~n10561;
  assign n10563 = ~n10558 & ~n10562;
  assign n10564 = ~n10557 & n10563;
  assign n10565 = n10557 & ~n10563;
  assign n10566 = ~n10564 & ~n10565;
  assign n10567 = ~pi477  & ~n10561;
  assign n10568 = pi477  & n10561;
  assign n10569 = ~n10567 & ~n10568;
  assign n10570 = ~pi480  & ~n10555;
  assign n10571 = pi480  & n10555;
  assign n10572 = ~n10570 & ~n10571;
  assign n10573 = ~n10569 & ~n10572;
  assign n10574 = ~n10566 & n10573;
  assign n10575 = ~n10557 & ~n10563;
  assign n10576 = ~n10574 & ~n10575;
  assign n10577 = pi484  & pi485 ;
  assign n10578 = ~pi484  & pi485 ;
  assign n10579 = pi484  & ~pi485 ;
  assign n10580 = ~n10578 & ~n10579;
  assign n10581 = pi486  & ~n10580;
  assign n10582 = ~n10577 & ~n10581;
  assign n10583 = pi481  & pi482 ;
  assign n10584 = ~pi481  & pi482 ;
  assign n10585 = pi481  & ~pi482 ;
  assign n10586 = ~n10584 & ~n10585;
  assign n10587 = pi483  & ~n10586;
  assign n10588 = ~n10583 & ~n10587;
  assign n10589 = ~n10582 & n10588;
  assign n10590 = n10582 & ~n10588;
  assign n10591 = ~n10589 & ~n10590;
  assign n10592 = ~pi483  & ~n10586;
  assign n10593 = pi483  & n10586;
  assign n10594 = ~n10592 & ~n10593;
  assign n10595 = ~pi486  & ~n10580;
  assign n10596 = pi486  & n10580;
  assign n10597 = ~n10595 & ~n10596;
  assign n10598 = ~n10594 & ~n10597;
  assign n10599 = ~n10591 & n10598;
  assign n10600 = ~n10582 & ~n10588;
  assign n10601 = ~n10599 & ~n10600;
  assign n10602 = n10591 & n10598;
  assign n10603 = ~n10591 & ~n10598;
  assign n10604 = ~n10602 & ~n10603;
  assign n10605 = n10566 & n10573;
  assign n10606 = ~n10566 & ~n10573;
  assign n10607 = ~n10605 & ~n10606;
  assign n10608 = ~n10576 & ~n10607;
  assign n10609 = ~n10601 & ~n10604;
  assign n10610 = ~n10594 & n10597;
  assign n10611 = n10594 & ~n10597;
  assign n10612 = ~n10610 & ~n10611;
  assign n10613 = ~n10569 & n10572;
  assign n10614 = n10569 & ~n10572;
  assign n10615 = ~n10613 & ~n10614;
  assign n10616 = ~n10612 & ~n10615;
  assign n10617 = ~n10608 & n10616;
  assign n10618 = ~n10609 & n10617;
  assign n10619 = n10604 & ~n10618;
  assign n10620 = ~n10604 & n10618;
  assign n10621 = ~n10619 & ~n10620;
  assign n10622 = n10607 & n10621;
  assign n10623 = ~n10619 & ~n10622;
  assign n10624 = n10601 & ~n10623;
  assign n10625 = ~n10576 & ~n10624;
  assign n10626 = ~n10601 & n10623;
  assign n10627 = ~n10625 & ~n10626;
  assign n10628 = ~pi466  & pi467 ;
  assign n10629 = pi466  & ~pi467 ;
  assign n10630 = ~n10628 & ~n10629;
  assign n10631 = ~pi468  & ~n10630;
  assign n10632 = pi468  & n10630;
  assign n10633 = ~n10631 & ~n10632;
  assign n10634 = ~pi463  & pi464 ;
  assign n10635 = pi463  & ~pi464 ;
  assign n10636 = ~n10634 & ~n10635;
  assign n10637 = ~pi465  & ~n10636;
  assign n10638 = pi465  & n10636;
  assign n10639 = ~n10637 & ~n10638;
  assign n10640 = ~n10633 & ~n10639;
  assign n10641 = pi466  & pi467 ;
  assign n10642 = pi468  & ~n10630;
  assign n10643 = ~n10641 & ~n10642;
  assign n10644 = pi463  & pi464 ;
  assign n10645 = pi465  & ~n10636;
  assign n10646 = ~n10644 & ~n10645;
  assign n10647 = n10643 & ~n10646;
  assign n10648 = ~n10643 & n10646;
  assign n10649 = ~n10647 & ~n10648;
  assign n10650 = n10640 & ~n10649;
  assign n10651 = ~n10643 & ~n10646;
  assign n10652 = ~n10650 & ~n10651;
  assign n10653 = pi472  & pi473 ;
  assign n10654 = ~pi472  & pi473 ;
  assign n10655 = pi472  & ~pi473 ;
  assign n10656 = ~n10654 & ~n10655;
  assign n10657 = pi474  & ~n10656;
  assign n10658 = ~n10653 & ~n10657;
  assign n10659 = pi469  & pi470 ;
  assign n10660 = ~pi469  & pi470 ;
  assign n10661 = pi469  & ~pi470 ;
  assign n10662 = ~n10660 & ~n10661;
  assign n10663 = pi471  & ~n10662;
  assign n10664 = ~n10659 & ~n10663;
  assign n10665 = ~n10658 & n10664;
  assign n10666 = n10658 & ~n10664;
  assign n10667 = ~n10665 & ~n10666;
  assign n10668 = ~pi471  & ~n10662;
  assign n10669 = pi471  & n10662;
  assign n10670 = ~n10668 & ~n10669;
  assign n10671 = ~pi474  & ~n10656;
  assign n10672 = pi474  & n10656;
  assign n10673 = ~n10671 & ~n10672;
  assign n10674 = ~n10670 & ~n10673;
  assign n10675 = ~n10667 & n10674;
  assign n10676 = ~n10658 & ~n10664;
  assign n10677 = ~n10675 & ~n10676;
  assign n10678 = n10667 & n10674;
  assign n10679 = ~n10667 & ~n10674;
  assign n10680 = ~n10678 & ~n10679;
  assign n10681 = n10640 & n10649;
  assign n10682 = ~n10640 & ~n10649;
  assign n10683 = ~n10681 & ~n10682;
  assign n10684 = ~n10652 & ~n10683;
  assign n10685 = ~n10677 & ~n10680;
  assign n10686 = ~n10670 & n10673;
  assign n10687 = n10670 & ~n10673;
  assign n10688 = ~n10686 & ~n10687;
  assign n10689 = ~n10633 & n10639;
  assign n10690 = n10633 & ~n10639;
  assign n10691 = ~n10689 & ~n10690;
  assign n10692 = ~n10688 & ~n10691;
  assign n10693 = ~n10684 & n10692;
  assign n10694 = ~n10685 & n10693;
  assign n10695 = n10680 & ~n10694;
  assign n10696 = ~n10680 & n10694;
  assign n10697 = ~n10695 & ~n10696;
  assign n10698 = n10683 & n10697;
  assign n10699 = ~n10695 & ~n10698;
  assign n10700 = n10677 & ~n10699;
  assign n10701 = ~n10652 & ~n10700;
  assign n10702 = ~n10677 & n10699;
  assign n10703 = ~n10701 & ~n10702;
  assign n10704 = n10627 & n10703;
  assign n10705 = ~n10652 & n10677;
  assign n10706 = n10652 & ~n10677;
  assign n10707 = ~n10705 & ~n10706;
  assign n10708 = n10699 & ~n10707;
  assign n10709 = ~n10699 & n10707;
  assign n10710 = ~n10708 & ~n10709;
  assign n10711 = ~n10576 & n10601;
  assign n10712 = n10576 & ~n10601;
  assign n10713 = ~n10711 & ~n10712;
  assign n10714 = n10623 & ~n10713;
  assign n10715 = ~n10623 & n10713;
  assign n10716 = ~n10714 & ~n10715;
  assign n10717 = n10710 & n10716;
  assign n10718 = n10688 & ~n10691;
  assign n10719 = ~n10688 & n10691;
  assign n10720 = ~n10718 & ~n10719;
  assign n10721 = n10612 & ~n10615;
  assign n10722 = ~n10612 & n10615;
  assign n10723 = ~n10721 & ~n10722;
  assign n10724 = ~n10720 & ~n10723;
  assign n10725 = ~n10607 & ~n10621;
  assign n10726 = ~n10622 & ~n10725;
  assign n10727 = ~n10724 & n10726;
  assign n10728 = ~n10683 & ~n10697;
  assign n10729 = ~n10698 & ~n10728;
  assign n10730 = n10724 & ~n10726;
  assign n10731 = ~n10727 & ~n10730;
  assign n10732 = n10729 & n10731;
  assign n10733 = ~n10727 & ~n10732;
  assign n10734 = ~n10710 & ~n10716;
  assign n10735 = ~n10717 & ~n10734;
  assign n10736 = n10733 & n10735;
  assign n10737 = ~n10717 & ~n10736;
  assign n10738 = ~n10704 & ~n10737;
  assign n10739 = ~n10627 & ~n10703;
  assign n10740 = ~n10738 & ~n10739;
  assign n10741 = ~n10551 & ~n10740;
  assign n10742 = n10551 & n10740;
  assign n10743 = ~n10741 & ~n10742;
  assign n10744 = ~n10514 & ~n10550;
  assign n10745 = ~n10548 & n10744;
  assign n10746 = n10548 & ~n10744;
  assign n10747 = ~n10745 & ~n10746;
  assign n10748 = ~n10704 & ~n10739;
  assign n10749 = ~n10737 & n10748;
  assign n10750 = n10737 & ~n10748;
  assign n10751 = ~n10749 & ~n10750;
  assign n10752 = n10747 & n10751;
  assign n10753 = ~n10733 & ~n10735;
  assign n10754 = ~n10736 & ~n10753;
  assign n10755 = ~n10544 & ~n10546;
  assign n10756 = ~n10547 & ~n10755;
  assign n10757 = n10754 & n10756;
  assign n10758 = ~n10754 & ~n10756;
  assign n10759 = ~n10757 & ~n10758;
  assign n10760 = ~n10720 & n10723;
  assign n10761 = n10720 & ~n10723;
  assign n10762 = ~n10760 & ~n10761;
  assign n10763 = ~n10530 & n10533;
  assign n10764 = n10530 & ~n10533;
  assign n10765 = ~n10763 & ~n10764;
  assign n10766 = ~n10762 & ~n10765;
  assign n10767 = ~n10539 & n10542;
  assign n10768 = ~n10543 & ~n10767;
  assign n10769 = ~n10766 & n10768;
  assign n10770 = ~n10729 & ~n10731;
  assign n10771 = ~n10732 & ~n10770;
  assign n10772 = n10766 & ~n10768;
  assign n10773 = ~n10769 & ~n10772;
  assign n10774 = n10771 & n10773;
  assign n10775 = ~n10769 & ~n10774;
  assign n10776 = n10759 & n10775;
  assign n10777 = ~n10757 & ~n10776;
  assign n10778 = ~n10747 & ~n10751;
  assign n10779 = ~n10752 & ~n10778;
  assign n10780 = ~n10777 & n10779;
  assign n10781 = ~n10752 & ~n10780;
  assign n10782 = n10743 & ~n10781;
  assign n10783 = ~n10741 & ~n10782;
  assign n10784 = ~n10361 & ~n10783;
  assign n10785 = ~n10743 & n10781;
  assign n10786 = ~n10782 & ~n10785;
  assign n10787 = ~n10321 & n10359;
  assign n10788 = ~n10360 & ~n10787;
  assign n10789 = n10786 & n10788;
  assign n10790 = n10355 & ~n10357;
  assign n10791 = ~n10358 & ~n10790;
  assign n10792 = n10777 & ~n10779;
  assign n10793 = ~n10780 & ~n10792;
  assign n10794 = n10791 & n10793;
  assign n10795 = ~n10791 & ~n10793;
  assign n10796 = ~n10794 & ~n10795;
  assign n10797 = ~n10759 & ~n10775;
  assign n10798 = ~n10776 & ~n10797;
  assign n10799 = ~n10337 & ~n10353;
  assign n10800 = ~n10354 & ~n10799;
  assign n10801 = n10798 & n10800;
  assign n10802 = ~n10762 & n10765;
  assign n10803 = n10762 & ~n10765;
  assign n10804 = ~n10802 & ~n10803;
  assign n10805 = ~n10340 & n10343;
  assign n10806 = n10340 & ~n10343;
  assign n10807 = ~n10805 & ~n10806;
  assign n10808 = ~n10804 & ~n10807;
  assign n10809 = ~n10349 & ~n10351;
  assign n10810 = ~n10352 & ~n10809;
  assign n10811 = ~n10808 & n10810;
  assign n10812 = ~n10771 & ~n10773;
  assign n10813 = ~n10774 & ~n10812;
  assign n10814 = n10808 & ~n10810;
  assign n10815 = ~n10811 & ~n10814;
  assign n10816 = n10813 & n10815;
  assign n10817 = ~n10811 & ~n10816;
  assign n10818 = ~n10798 & ~n10800;
  assign n10819 = ~n10801 & ~n10818;
  assign n10820 = n10817 & n10819;
  assign n10821 = ~n10801 & ~n10820;
  assign n10822 = n10796 & ~n10821;
  assign n10823 = ~n10794 & ~n10822;
  assign n10824 = ~n10786 & ~n10788;
  assign n10825 = ~n10789 & ~n10824;
  assign n10826 = ~n10823 & n10825;
  assign n10827 = ~n10789 & ~n10826;
  assign n10828 = n10361 & n10783;
  assign n10829 = ~n10784 & ~n10828;
  assign n10830 = ~n10827 & n10829;
  assign n10831 = ~n10784 & ~n10830;
  assign n10832 = ~n9939 & ~n10831;
  assign n10833 = n9939 & n10831;
  assign n10834 = ~n10832 & ~n10833;
  assign n10835 = n9935 & ~n9937;
  assign n10836 = ~n9938 & ~n10835;
  assign n10837 = n10827 & ~n10829;
  assign n10838 = ~n10830 & ~n10837;
  assign n10839 = n10836 & n10838;
  assign n10840 = ~n10817 & ~n10819;
  assign n10841 = ~n10820 & ~n10840;
  assign n10842 = ~n9911 & ~n9927;
  assign n10843 = ~n9928 & ~n10842;
  assign n10844 = n10841 & n10843;
  assign n10845 = ~n10841 & ~n10843;
  assign n10846 = ~n10844 & ~n10845;
  assign n10847 = ~n10804 & n10807;
  assign n10848 = n10804 & ~n10807;
  assign n10849 = ~n10847 & ~n10848;
  assign n10850 = ~n9914 & n9917;
  assign n10851 = n9914 & ~n9917;
  assign n10852 = ~n10850 & ~n10851;
  assign n10853 = ~n10849 & ~n10852;
  assign n10854 = ~n9923 & ~n9925;
  assign n10855 = ~n9926 & ~n10854;
  assign n10856 = ~n10853 & n10855;
  assign n10857 = ~n10813 & ~n10815;
  assign n10858 = ~n10816 & ~n10857;
  assign n10859 = n10853 & ~n10855;
  assign n10860 = ~n10856 & ~n10859;
  assign n10861 = n10858 & n10860;
  assign n10862 = ~n10856 & ~n10861;
  assign n10863 = n10846 & n10862;
  assign n10864 = ~n10844 & ~n10863;
  assign n10865 = ~n9904 & n9929;
  assign n10866 = ~n9930 & ~n10865;
  assign n10867 = ~n10796 & n10821;
  assign n10868 = ~n10822 & ~n10867;
  assign n10869 = ~n10866 & ~n10868;
  assign n10870 = ~n10864 & ~n10869;
  assign n10871 = n10866 & n10868;
  assign n10872 = ~n10870 & ~n10871;
  assign n10873 = n10823 & ~n10825;
  assign n10874 = ~n10826 & ~n10873;
  assign n10875 = n9931 & ~n9933;
  assign n10876 = ~n9934 & ~n10875;
  assign n10877 = ~n10874 & ~n10876;
  assign n10878 = ~n10872 & ~n10877;
  assign n10879 = n10874 & n10876;
  assign n10880 = ~n10878 & ~n10879;
  assign n10881 = ~n10836 & ~n10838;
  assign n10882 = ~n10839 & ~n10881;
  assign n10883 = ~n10880 & n10882;
  assign n10884 = ~n10839 & ~n10883;
  assign n10885 = n10834 & ~n10884;
  assign n10886 = ~n10832 & ~n10885;
  assign n10887 = ~n9047 & ~n10886;
  assign n10888 = n9047 & n10886;
  assign n10889 = ~n10887 & ~n10888;
  assign n10890 = ~n10834 & n10884;
  assign n10891 = ~n10885 & ~n10890;
  assign n10892 = ~n8996 & n9045;
  assign n10893 = ~n9046 & ~n10892;
  assign n10894 = n10891 & n10893;
  assign n10895 = n9041 & ~n9043;
  assign n10896 = ~n9044 & ~n10895;
  assign n10897 = n10880 & ~n10882;
  assign n10898 = ~n10883 & ~n10897;
  assign n10899 = n10896 & n10898;
  assign n10900 = ~n10877 & ~n10879;
  assign n10901 = ~n10872 & n10900;
  assign n10902 = n10872 & ~n10900;
  assign n10903 = ~n10901 & ~n10902;
  assign n10904 = ~n9038 & ~n9040;
  assign n10905 = ~n9033 & n10904;
  assign n10906 = n9033 & ~n10904;
  assign n10907 = ~n10905 & ~n10906;
  assign n10908 = n10903 & n10907;
  assign n10909 = ~n9030 & ~n9032;
  assign n10910 = ~n9025 & n10909;
  assign n10911 = n9025 & ~n10909;
  assign n10912 = ~n10910 & ~n10911;
  assign n10913 = ~n10869 & ~n10871;
  assign n10914 = ~n10864 & n10913;
  assign n10915 = n10864 & ~n10913;
  assign n10916 = ~n10914 & ~n10915;
  assign n10917 = n10912 & n10916;
  assign n10918 = ~n10912 & ~n10916;
  assign n10919 = ~n10917 & ~n10918;
  assign n10920 = ~n10846 & ~n10862;
  assign n10921 = ~n10863 & ~n10920;
  assign n10922 = n9021 & ~n9023;
  assign n10923 = ~n9024 & ~n10922;
  assign n10924 = n10921 & n10923;
  assign n10925 = ~n10849 & n10852;
  assign n10926 = n10849 & ~n10852;
  assign n10927 = ~n10925 & ~n10926;
  assign n10928 = ~n9009 & n9012;
  assign n10929 = n9009 & ~n9012;
  assign n10930 = ~n10928 & ~n10929;
  assign n10931 = ~n10927 & ~n10930;
  assign n10932 = ~n9016 & ~n9019;
  assign n10933 = ~n9018 & ~n10932;
  assign n10934 = n9018 & n10932;
  assign n10935 = ~n10933 & ~n10934;
  assign n10936 = ~n10931 & n10935;
  assign n10937 = ~n10858 & ~n10860;
  assign n10938 = ~n10861 & ~n10937;
  assign n10939 = n10931 & ~n10935;
  assign n10940 = ~n10936 & ~n10939;
  assign n10941 = n10938 & n10940;
  assign n10942 = ~n10936 & ~n10941;
  assign n10943 = ~n10921 & ~n10923;
  assign n10944 = ~n10924 & ~n10943;
  assign n10945 = n10942 & n10944;
  assign n10946 = ~n10924 & ~n10945;
  assign n10947 = n10919 & ~n10946;
  assign n10948 = ~n10917 & ~n10947;
  assign n10949 = ~n10903 & ~n10907;
  assign n10950 = ~n10908 & ~n10949;
  assign n10951 = ~n10948 & n10950;
  assign n10952 = ~n10908 & ~n10951;
  assign n10953 = ~n10896 & ~n10898;
  assign n10954 = ~n10899 & ~n10953;
  assign n10955 = ~n10952 & n10954;
  assign n10956 = ~n10899 & ~n10955;
  assign n10957 = ~n10891 & ~n10893;
  assign n10958 = ~n10894 & ~n10957;
  assign n10959 = ~n10956 & n10958;
  assign n10960 = ~n10894 & ~n10959;
  assign n10961 = n10889 & ~n10960;
  assign n10962 = ~n10887 & ~n10961;
  assign n10963 = n7209 & ~n10962;
  assign n10964 = ~n7209 & n10962;
  assign n10965 = ~n10963 & ~n10964;
  assign n10966 = n7201 & ~n7203;
  assign n10967 = ~n7204 & ~n10966;
  assign n10968 = ~n10889 & n10960;
  assign n10969 = ~n10961 & ~n10968;
  assign n10970 = n10967 & n10969;
  assign n10971 = ~n10967 & ~n10969;
  assign n10972 = ~n10970 & ~n10971;
  assign n10973 = ~n7198 & ~n7200;
  assign n10974 = ~n7193 & n10973;
  assign n10975 = n7193 & ~n10973;
  assign n10976 = ~n10974 & ~n10975;
  assign n10977 = n10956 & ~n10958;
  assign n10978 = ~n10959 & ~n10977;
  assign n10979 = n10976 & n10978;
  assign n10980 = ~n10976 & ~n10978;
  assign n10981 = ~n10979 & ~n10980;
  assign n10982 = n7189 & ~n7191;
  assign n10983 = ~n7192 & ~n10982;
  assign n10984 = n10952 & ~n10954;
  assign n10985 = ~n10955 & ~n10984;
  assign n10986 = n10983 & n10985;
  assign n10987 = ~n7186 & ~n7188;
  assign n10988 = ~n7181 & n10987;
  assign n10989 = n7181 & ~n10987;
  assign n10990 = ~n10988 & ~n10989;
  assign n10991 = n10948 & ~n10950;
  assign n10992 = ~n10951 & ~n10991;
  assign n10993 = n10990 & n10992;
  assign n10994 = ~n7151 & ~n7179;
  assign n10995 = ~n7178 & n10994;
  assign n10996 = n7178 & ~n10994;
  assign n10997 = ~n10995 & ~n10996;
  assign n10998 = ~n10919 & n10946;
  assign n10999 = ~n10947 & ~n10998;
  assign n11000 = ~n10997 & ~n10999;
  assign n11001 = ~n7175 & ~n7177;
  assign n11002 = ~n7170 & n11001;
  assign n11003 = n7170 & ~n11001;
  assign n11004 = ~n11002 & ~n11003;
  assign n11005 = ~n10942 & ~n10944;
  assign n11006 = ~n10945 & ~n11005;
  assign n11007 = n11004 & n11006;
  assign n11008 = ~n10938 & ~n10940;
  assign n11009 = ~n10941 & ~n11008;
  assign n11010 = ~n10927 & n10930;
  assign n11011 = n10927 & ~n10930;
  assign n11012 = ~n11010 & ~n11011;
  assign n11013 = ~n7154 & n7157;
  assign n11014 = n7154 & ~n7157;
  assign n11015 = ~n11013 & ~n11014;
  assign n11016 = ~n11012 & ~n11015;
  assign n11017 = ~n7163 & ~n7168;
  assign n11018 = ~n7167 & ~n11017;
  assign n11019 = n7167 & n11017;
  assign n11020 = ~n11018 & ~n11019;
  assign n11021 = ~n11016 & n11020;
  assign n11022 = ~n11009 & ~n11021;
  assign n11023 = n11016 & ~n11020;
  assign n11024 = ~n11022 & ~n11023;
  assign n11025 = ~n11004 & ~n11006;
  assign n11026 = ~n11007 & ~n11025;
  assign n11027 = ~n11024 & n11026;
  assign n11028 = ~n11007 & ~n11027;
  assign n11029 = ~n11000 & ~n11028;
  assign n11030 = n10997 & n10999;
  assign n11031 = ~n11029 & ~n11030;
  assign n11032 = ~n10990 & ~n10992;
  assign n11033 = ~n10993 & ~n11032;
  assign n11034 = ~n11031 & n11033;
  assign n11035 = ~n10993 & ~n11034;
  assign n11036 = ~n10983 & ~n10985;
  assign n11037 = ~n10986 & ~n11036;
  assign n11038 = ~n11035 & n11037;
  assign n11039 = ~n10986 & ~n11038;
  assign n11040 = n10981 & ~n11039;
  assign n11041 = ~n10979 & ~n11040;
  assign n11042 = n10972 & ~n11041;
  assign n11043 = ~n10970 & ~n11042;
  assign n11044 = n10965 & ~n11043;
  assign n11045 = ~n10963 & ~n11044;
  assign n11046 = n7207 & ~n11045;
  assign n11047 = ~n7207 & n11045;
  assign n11048 = ~n11046 & ~n11047;
  assign n11049 = ~n11000 & ~n11030;
  assign n11050 = n11028 & ~n11049;
  assign n11051 = ~n11028 & n11049;
  assign n11052 = ~n11050 & ~n11051;
  assign n11053 = n11024 & ~n11026;
  assign n11054 = ~n11027 & ~n11053;
  assign n11055 = n11012 & ~n11015;
  assign n11056 = ~n11012 & n11015;
  assign n11057 = ~n11055 & ~n11056;
  assign n11058 = pi1000  & ~n11057;
  assign n11059 = ~n11021 & ~n11023;
  assign n11060 = n11009 & n11059;
  assign n11061 = ~n11009 & ~n11059;
  assign n11062 = ~n11060 & ~n11061;
  assign n11063 = n11058 & ~n11062;
  assign n11064 = n11054 & n11063;
  assign n11065 = n11052 & n11064;
  assign n11066 = n11031 & ~n11033;
  assign n11067 = ~n11034 & ~n11066;
  assign n11068 = n11065 & n11067;
  assign n11069 = n11035 & ~n11037;
  assign n11070 = ~n11038 & ~n11069;
  assign n11071 = n11068 & n11070;
  assign n11072 = ~n10981 & n11039;
  assign n11073 = ~n11040 & ~n11072;
  assign n11074 = n11071 & n11073;
  assign n11075 = ~n10972 & n11041;
  assign n11076 = ~n11042 & ~n11075;
  assign n11077 = n11074 & n11076;
  assign n11078 = ~n10965 & n11043;
  assign n11079 = ~n11044 & ~n11078;
  assign n11080 = n11077 & n11079;
  assign n11081 = n11048 & n11080;
  assign n11082 = ~n11048 & ~n11080;
  assign n11083 = ~n11081 & ~n11082;
  assign n11084 = ~n11054 & ~n11063;
  assign n11085 = ~n11064 & ~n11084;
  assign n11086 = ~n11058 & ~n11062;
  assign n11087 = n11058 & n11062;
  assign n11088 = ~n11086 & ~n11087;
  assign n11089 = ~n11085 & n11088;
  assign n11090 = ~n11052 & ~n11064;
  assign n11091 = ~n11065 & ~n11090;
  assign n11092 = ~n11089 & n11091;
  assign n11093 = ~n11065 & ~n11067;
  assign n11094 = ~n11068 & ~n11093;
  assign n11095 = ~n11092 & ~n11094;
  assign n11096 = ~n11068 & ~n11070;
  assign n11097 = ~n11071 & ~n11096;
  assign n11098 = ~n11095 & n11097;
  assign n11099 = ~n11071 & ~n11073;
  assign n11100 = ~n11074 & ~n11099;
  assign n11101 = n11098 & n11100;
  assign n11102 = ~n11074 & ~n11076;
  assign n11103 = ~n11077 & ~n11102;
  assign n11104 = n11101 & n11103;
  assign n11105 = ~n11077 & ~n11079;
  assign n11106 = ~n11080 & ~n11105;
  assign n11107 = n11104 & n11106;
  assign n11108 = ~n11083 & n11107;
  assign n11109 = ~n7207 & ~n11045;
  assign n11110 = n11080 & ~n11081;
  assign n11111 = ~n11109 & ~n11110;
  assign n11112 = ~n11108 & n11111;
  assign n11113 = n11089 & ~n11091;
  assign n11114 = ~n11092 & ~n11113;
  assign n11115 = ~pi1000  & ~n11057;
  assign n11116 = pi1000  & n11057;
  assign n11117 = ~n11115 & ~n11116;
  assign n11118 = n11085 & ~n11088;
  assign n11119 = ~n11089 & ~n11118;
  assign n11120 = n11117 & n11119;
  assign n11121 = n11085 & ~n11120;
  assign n11122 = ~n11117 & ~n11119;
  assign n11123 = ~n11121 & ~n11122;
  assign n11124 = ~n11114 & n11123;
  assign n11125 = n11091 & ~n11124;
  assign n11126 = n11114 & ~n11123;
  assign n11127 = ~n11125 & ~n11126;
  assign n11128 = ~n11092 & ~n11127;
  assign n11129 = n11092 & n11094;
  assign n11130 = n11095 & ~n11097;
  assign n11131 = ~n11098 & ~n11130;
  assign n11132 = ~n11129 & ~n11131;
  assign n11133 = ~n11128 & n11132;
  assign n11134 = n11097 & ~n11133;
  assign n11135 = ~n11128 & ~n11129;
  assign n11136 = n11131 & ~n11135;
  assign n11137 = ~n11134 & ~n11136;
  assign n11138 = n11098 & ~n11137;
  assign n11139 = ~n11098 & n11100;
  assign n11140 = ~n11101 & ~n11103;
  assign n11141 = ~n11104 & ~n11140;
  assign n11142 = ~n11139 & ~n11141;
  assign n11143 = ~n11138 & n11142;
  assign n11144 = n11103 & ~n11143;
  assign n11145 = ~n11138 & ~n11139;
  assign n11146 = n11141 & ~n11145;
  assign n11147 = ~n11144 & ~n11146;
  assign n11148 = n11104 & ~n11107;
  assign n11149 = ~n11147 & n11148;
  assign n11150 = n11107 & n11143;
  assign n11151 = n11106 & ~n11150;
  assign n11152 = ~n11149 & ~n11151;
  assign n11153 = n11107 & ~n11108;
  assign n11154 = ~n11152 & n11153;
  assign n11155 = n11083 & ~n11154;
  assign n11156 = n11112 & ~n11155;
  assign po0 = ~n11112 | n11156;
endmodule
