module mem_ctrl ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17,
    pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26,
    pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44,
    pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53,
    pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62,
    pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80,
    pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107,
    pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116,
    pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125,
    pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134,
    pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143,
    pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152,
    pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161,
    pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170,
    pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197,
    pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206,
    pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215,
    pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224,
    pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233,
    pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242,
    pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251,
    pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260,
    pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287,
    pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296,
    pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305,
    pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314,
    pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323,
    pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332,
    pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341,
    pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350,
    pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377,
    pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386,
    pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395,
    pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404,
    pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413,
    pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422,
    pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431,
    pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440,
    pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467,
    pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476,
    pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485,
    pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494,
    pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503,
    pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, pi512,
    pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520, pi521,
    pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529, pi530,
    pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539,
    pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548,
    pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557,
    pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566,
    pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574, pi575,
    pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583, pi584,
    pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592, pi593,
    pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601, pi602,
    pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610, pi611,
    pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619, pi620,
    pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629,
    pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638,
    pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647,
    pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656,
    pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664, pi665,
    pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673, pi674,
    pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682, pi683,
    pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691, pi692,
    pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700, pi701,
    pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709, pi710,
    pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719,
    pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728,
    pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737,
    pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746,
    pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754, pi755,
    pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763, pi764,
    pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772, pi773,
    pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781, pi782,
    pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790, pi791,
    pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799, pi800,
    pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808, pi809,
    pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818,
    pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827,
    pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835, pi836,
    pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844, pi845,
    pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853, pi854,
    pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862, pi863,
    pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871, pi872,
    pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880, pi881,
    pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889, pi890,
    pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898, pi899,
    pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907, pi908,
    pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916, pi917,
    pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925, pi926,
    pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934, pi935,
    pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943, pi944,
    pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952, pi953,
    pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961, pi962,
    pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970, pi971,
    pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979, pi980,
    pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988, pi989,
    pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997, pi998,
    pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0, po1, po2, po3, po4, po5, po6, po7, po8,
    po9, po10, po11, po12, po13, po14, po15, po16, po17,
    po18, po19, po20, po21, po22, po23, po24, po25, po26,
    po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44,
    po45, po46, po47, po48, po49, po50, po51, po52, po53,
    po54, po55, po56, po57, po58, po59, po60, po61, po62,
    po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80,
    po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98,
    po99, po100, po101, po102, po103, po104, po105, po106, po107,
    po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125,
    po126, po127, po128, po129, po130, po131, po132, po133, po134,
    po135, po136, po137, po138, po139, po140, po141, po142, po143,
    po144, po145, po146, po147, po148, po149, po150, po151, po152,
    po153, po154, po155, po156, po157, po158, po159, po160, po161,
    po162, po163, po164, po165, po166, po167, po168, po169, po170,
    po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188,
    po189, po190, po191, po192, po193, po194, po195, po196, po197,
    po198, po199, po200, po201, po202, po203, po204, po205, po206,
    po207, po208, po209, po210, po211, po212, po213, po214, po215,
    po216, po217, po218, po219, po220, po221, po222, po223, po224,
    po225, po226, po227, po228, po229, po230, po231, po232, po233,
    po234, po235, po236, po237, po238, po239, po240, po241, po242,
    po243, po244, po245, po246, po247, po248, po249, po250, po251,
    po252, po253, po254, po255, po256, po257, po258, po259, po260,
    po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278,
    po279, po280, po281, po282, po283, po284, po285, po286, po287,
    po288, po289, po290, po291, po292, po293, po294, po295, po296,
    po297, po298, po299, po300, po301, po302, po303, po304, po305,
    po306, po307, po308, po309, po310, po311, po312, po313, po314,
    po315, po316, po317, po318, po319, po320, po321, po322, po323,
    po324, po325, po326, po327, po328, po329, po330, po331, po332,
    po333, po334, po335, po336, po337, po338, po339, po340, po341,
    po342, po343, po344, po345, po346, po347, po348, po349, po350,
    po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368,
    po369, po370, po371, po372, po373, po374, po375, po376, po377,
    po378, po379, po380, po381, po382, po383, po384, po385, po386,
    po387, po388, po389, po390, po391, po392, po393, po394, po395,
    po396, po397, po398, po399, po400, po401, po402, po403, po404,
    po405, po406, po407, po408, po409, po410, po411, po412, po413,
    po414, po415, po416, po417, po418, po419, po420, po421, po422,
    po423, po424, po425, po426, po427, po428, po429, po430, po431,
    po432, po433, po434, po435, po436, po437, po438, po439, po440,
    po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458,
    po459, po460, po461, po462, po463, po464, po465, po466, po467,
    po468, po469, po470, po471, po472, po473, po474, po475, po476,
    po477, po478, po479, po480, po481, po482, po483, po484, po485,
    po486, po487, po488, po489, po490, po491, po492, po493, po494,
    po495, po496, po497, po498, po499, po500, po501, po502, po503,
    po504, po505, po506, po507, po508, po509, po510, po511, po512,
    po513, po514, po515, po516, po517, po518, po519, po520, po521,
    po522, po523, po524, po525, po526, po527, po528, po529, po530,
    po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548,
    po549, po550, po551, po552, po553, po554, po555, po556, po557,
    po558, po559, po560, po561, po562, po563, po564, po565, po566,
    po567, po568, po569, po570, po571, po572, po573, po574, po575,
    po576, po577, po578, po579, po580, po581, po582, po583, po584,
    po585, po586, po587, po588, po589, po590, po591, po592, po593,
    po594, po595, po596, po597, po598, po599, po600, po601, po602,
    po603, po604, po605, po606, po607, po608, po609, po610, po611,
    po612, po613, po614, po615, po616, po617, po618, po619, po620,
    po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638,
    po639, po640, po641, po642, po643, po644, po645, po646, po647,
    po648, po649, po650, po651, po652, po653, po654, po655, po656,
    po657, po658, po659, po660, po661, po662, po663, po664, po665,
    po666, po667, po668, po669, po670, po671, po672, po673, po674,
    po675, po676, po677, po678, po679, po680, po681, po682, po683,
    po684, po685, po686, po687, po688, po689, po690, po691, po692,
    po693, po694, po695, po696, po697, po698, po699, po700, po701,
    po702, po703, po704, po705, po706, po707, po708, po709, po710,
    po711, po712, po713, po714, po715, po716, po717, po718, po719,
    po720, po721, po722, po723, po724, po725, po726, po727, po728,
    po729, po730, po731, po732, po733, po734, po735, po736, po737,
    po738, po739, po740, po741, po742, po743, po744, po745, po746,
    po747, po748, po749, po750, po751, po752, po753, po754, po755,
    po756, po757, po758, po759, po760, po761, po762, po763, po764,
    po765, po766, po767, po768, po769, po770, po771, po772, po773,
    po774, po775, po776, po777, po778, po779, po780, po781, po782,
    po783, po784, po785, po786, po787, po788, po789, po790, po791,
    po792, po793, po794, po795, po796, po797, po798, po799, po800,
    po801, po802, po803, po804, po805, po806, po807, po808, po809,
    po810, po811, po812, po813, po814, po815, po816, po817, po818,
    po819, po820, po821, po822, po823, po824, po825, po826, po827,
    po828, po829, po830, po831, po832, po833, po834, po835, po836,
    po837, po838, po839, po840, po841, po842, po843, po844, po845,
    po846, po847, po848, po849, po850, po851, po852, po853, po854,
    po855, po856, po857, po858, po859, po860, po861, po862, po863,
    po864, po865, po866, po867, po868, po869, po870, po871, po872,
    po873, po874, po875, po876, po877, po878, po879, po880, po881,
    po882, po883, po884, po885, po886, po887, po888, po889, po890,
    po891, po892, po893, po894, po895, po896, po897, po898, po899,
    po900, po901, po902, po903, po904, po905, po906, po907, po908,
    po909, po910, po911, po912, po913, po914, po915, po916, po917,
    po918, po919, po920, po921, po922, po923, po924, po925, po926,
    po927, po928, po929, po930, po931, po932, po933, po934, po935,
    po936, po937, po938, po939, po940, po941, po942, po943, po944,
    po945, po946, po947, po948, po949, po950, po951, po952, po953,
    po954, po955, po956, po957, po958, po959, po960, po961, po962,
    po963, po964, po965, po966, po967, po968, po969, po970, po971,
    po972, po973, po974, po975, po976, po977, po978, po979, po980,
    po981, po982, po983, po984, po985, po986, po987, po988, po989,
    po990, po991, po992, po993, po994, po995, po996, po997, po998,
    po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7,
    pi8, pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16,
    pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25,
    pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34,
    pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43,
    pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52,
    pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61,
    pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70,
    pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97,
    pi98, pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106,
    pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115,
    pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124,
    pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133,
    pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142,
    pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151,
    pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160,
    pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187,
    pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196,
    pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205,
    pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214,
    pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223,
    pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232,
    pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241,
    pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250,
    pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277,
    pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286,
    pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295,
    pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304,
    pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313,
    pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322,
    pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331,
    pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340,
    pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367,
    pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376,
    pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385,
    pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394,
    pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403,
    pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412,
    pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421,
    pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430,
    pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457,
    pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466,
    pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475,
    pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484,
    pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493,
    pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502,
    pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511,
    pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520,
    pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529,
    pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538,
    pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547,
    pi548, pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556,
    pi557, pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565,
    pi566, pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574,
    pi575, pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583,
    pi584, pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592,
    pi593, pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601,
    pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610,
    pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619,
    pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628,
    pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637,
    pi638, pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646,
    pi647, pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655,
    pi656, pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664,
    pi665, pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673,
    pi674, pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682,
    pi683, pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691,
    pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700,
    pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709,
    pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718,
    pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727,
    pi728, pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736,
    pi737, pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745,
    pi746, pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754,
    pi755, pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763,
    pi764, pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772,
    pi773, pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781,
    pi782, pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790,
    pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799,
    pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808,
    pi809, pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817,
    pi818, pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826,
    pi827, pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835,
    pi836, pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844,
    pi845, pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853,
    pi854, pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862,
    pi863, pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871,
    pi872, pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880,
    pi881, pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889,
    pi890, pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898,
    pi899, pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907,
    pi908, pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916,
    pi917, pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925,
    pi926, pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934,
    pi935, pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943,
    pi944, pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952,
    pi953, pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961,
    pi962, pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970,
    pi971, pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979,
    pi980, pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988,
    pi989, pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997,
    pi998, pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0, po1, po2, po3, po4, po5, po6, po7,
    po8, po9, po10, po11, po12, po13, po14, po15, po16,
    po17, po18, po19, po20, po21, po22, po23, po24, po25,
    po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43,
    po44, po45, po46, po47, po48, po49, po50, po51, po52,
    po53, po54, po55, po56, po57, po58, po59, po60, po61,
    po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88,
    po89, po90, po91, po92, po93, po94, po95, po96, po97,
    po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115,
    po116, po117, po118, po119, po120, po121, po122, po123, po124,
    po125, po126, po127, po128, po129, po130, po131, po132, po133,
    po134, po135, po136, po137, po138, po139, po140, po141, po142,
    po143, po144, po145, po146, po147, po148, po149, po150, po151,
    po152, po153, po154, po155, po156, po157, po158, po159, po160,
    po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178,
    po179, po180, po181, po182, po183, po184, po185, po186, po187,
    po188, po189, po190, po191, po192, po193, po194, po195, po196,
    po197, po198, po199, po200, po201, po202, po203, po204, po205,
    po206, po207, po208, po209, po210, po211, po212, po213, po214,
    po215, po216, po217, po218, po219, po220, po221, po222, po223,
    po224, po225, po226, po227, po228, po229, po230, po231, po232,
    po233, po234, po235, po236, po237, po238, po239, po240, po241,
    po242, po243, po244, po245, po246, po247, po248, po249, po250,
    po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268,
    po269, po270, po271, po272, po273, po274, po275, po276, po277,
    po278, po279, po280, po281, po282, po283, po284, po285, po286,
    po287, po288, po289, po290, po291, po292, po293, po294, po295,
    po296, po297, po298, po299, po300, po301, po302, po303, po304,
    po305, po306, po307, po308, po309, po310, po311, po312, po313,
    po314, po315, po316, po317, po318, po319, po320, po321, po322,
    po323, po324, po325, po326, po327, po328, po329, po330, po331,
    po332, po333, po334, po335, po336, po337, po338, po339, po340,
    po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358,
    po359, po360, po361, po362, po363, po364, po365, po366, po367,
    po368, po369, po370, po371, po372, po373, po374, po375, po376,
    po377, po378, po379, po380, po381, po382, po383, po384, po385,
    po386, po387, po388, po389, po390, po391, po392, po393, po394,
    po395, po396, po397, po398, po399, po400, po401, po402, po403,
    po404, po405, po406, po407, po408, po409, po410, po411, po412,
    po413, po414, po415, po416, po417, po418, po419, po420, po421,
    po422, po423, po424, po425, po426, po427, po428, po429, po430,
    po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448,
    po449, po450, po451, po452, po453, po454, po455, po456, po457,
    po458, po459, po460, po461, po462, po463, po464, po465, po466,
    po467, po468, po469, po470, po471, po472, po473, po474, po475,
    po476, po477, po478, po479, po480, po481, po482, po483, po484,
    po485, po486, po487, po488, po489, po490, po491, po492, po493,
    po494, po495, po496, po497, po498, po499, po500, po501, po502,
    po503, po504, po505, po506, po507, po508, po509, po510, po511,
    po512, po513, po514, po515, po516, po517, po518, po519, po520,
    po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538,
    po539, po540, po541, po542, po543, po544, po545, po546, po547,
    po548, po549, po550, po551, po552, po553, po554, po555, po556,
    po557, po558, po559, po560, po561, po562, po563, po564, po565,
    po566, po567, po568, po569, po570, po571, po572, po573, po574,
    po575, po576, po577, po578, po579, po580, po581, po582, po583,
    po584, po585, po586, po587, po588, po589, po590, po591, po592,
    po593, po594, po595, po596, po597, po598, po599, po600, po601,
    po602, po603, po604, po605, po606, po607, po608, po609, po610,
    po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628,
    po629, po630, po631, po632, po633, po634, po635, po636, po637,
    po638, po639, po640, po641, po642, po643, po644, po645, po646,
    po647, po648, po649, po650, po651, po652, po653, po654, po655,
    po656, po657, po658, po659, po660, po661, po662, po663, po664,
    po665, po666, po667, po668, po669, po670, po671, po672, po673,
    po674, po675, po676, po677, po678, po679, po680, po681, po682,
    po683, po684, po685, po686, po687, po688, po689, po690, po691,
    po692, po693, po694, po695, po696, po697, po698, po699, po700,
    po701, po702, po703, po704, po705, po706, po707, po708, po709,
    po710, po711, po712, po713, po714, po715, po716, po717, po718,
    po719, po720, po721, po722, po723, po724, po725, po726, po727,
    po728, po729, po730, po731, po732, po733, po734, po735, po736,
    po737, po738, po739, po740, po741, po742, po743, po744, po745,
    po746, po747, po748, po749, po750, po751, po752, po753, po754,
    po755, po756, po757, po758, po759, po760, po761, po762, po763,
    po764, po765, po766, po767, po768, po769, po770, po771, po772,
    po773, po774, po775, po776, po777, po778, po779, po780, po781,
    po782, po783, po784, po785, po786, po787, po788, po789, po790,
    po791, po792, po793, po794, po795, po796, po797, po798, po799,
    po800, po801, po802, po803, po804, po805, po806, po807, po808,
    po809, po810, po811, po812, po813, po814, po815, po816, po817,
    po818, po819, po820, po821, po822, po823, po824, po825, po826,
    po827, po828, po829, po830, po831, po832, po833, po834, po835,
    po836, po837, po838, po839, po840, po841, po842, po843, po844,
    po845, po846, po847, po848, po849, po850, po851, po852, po853,
    po854, po855, po856, po857, po858, po859, po860, po861, po862,
    po863, po864, po865, po866, po867, po868, po869, po870, po871,
    po872, po873, po874, po875, po876, po877, po878, po879, po880,
    po881, po882, po883, po884, po885, po886, po887, po888, po889,
    po890, po891, po892, po893, po894, po895, po896, po897, po898,
    po899, po900, po901, po902, po903, po904, po905, po906, po907,
    po908, po909, po910, po911, po912, po913, po914, po915, po916,
    po917, po918, po919, po920, po921, po922, po923, po924, po925,
    po926, po927, po928, po929, po930, po931, po932, po933, po934,
    po935, po936, po937, po938, po939, po940, po941, po942, po943,
    po944, po945, po946, po947, po948, po949, po950, po951, po952,
    po953, po954, po955, po956, po957, po958, po959, po960, po961,
    po962, po963, po964, po965, po966, po967, po968, po969, po970,
    po971, po972, po973, po974, po975, po976, po977, po978, po979,
    po980, po981, po982, po983, po984, po985, po986, po987, po988,
    po989, po990, po991, po992, po993, po994, po995, po996, po997,
    po998, po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671,
    n2672, n2673, n2674, n2675, n2676, n2677,
    n2678, n2679, n2680, n2681, n2682, n2683,
    n2684, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695,
    n2696, n2697, n2698, n2699, n2700, n2701,
    n2702, n2703, n2704, n2705, n2706, n2707,
    n2708, n2709, n2710, n2711, n2712, n2713,
    n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731,
    n2732, n2733, n2734, n2735, n2736, n2737,
    n2738, n2739, n2740, n2741, n2742, n2743,
    n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761,
    n2762, n2763, n2764, n2765, n2766, n2767,
    n2768, n2769, n2770, n2771, n2772, n2773,
    n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791,
    n2792, n2793, n2794, n2795, n2796, n2797,
    n2798, n2799, n2800, n2801, n2802, n2803,
    n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821,
    n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851,
    n2852, n2853, n2854, n2855, n2856, n2857,
    n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2878, n2879, n2880, n2881,
    n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893,
    n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905,
    n2906, n2907, n2908, n2909, n2910, n2911,
    n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2940, n2941,
    n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953,
    n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971,
    n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001,
    n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013,
    n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031,
    n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055,
    n3056, n3057, n3058, n3059, n3060, n3061,
    n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085,
    n3086, n3087, n3088, n3089, n3090, n3091,
    n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109,
    n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3117, n3118, n3119, n3120, n3121,
    n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151,
    n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3174, n3175,
    n3176, n3177, n3178, n3179, n3180, n3181,
    n3182, n3183, n3184, n3185, n3186, n3187,
    n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211,
    n3212, n3213, n3214, n3215, n3216, n3217,
    n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241,
    n3242, n3243, n3244, n3245, n3246, n3247,
    n3248, n3249, n3250, n3251, n3252, n3253,
    n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265,
    n3266, n3267, n3268, n3269, n3270, n3271,
    n3272, n3273, n3274, n3275, n3276, n3277,
    n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535,
    n3536, n3537, n3538, n3539, n3540, n3541,
    n3542, n3543, n3544, n3545, n3546, n3547,
    n3548, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565,
    n3566, n3567, n3568, n3569, n3570, n3571,
    n3572, n3573, n3574, n3575, n3576, n3577,
    n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601,
    n3602, n3603, n3604, n3605, n3606, n3607,
    n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631,
    n3632, n3633, n3634, n3635, n3636, n3637,
    n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661,
    n3662, n3663, n3664, n3665, n3666, n3667,
    n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691,
    n3692, n3693, n3694, n3695, n3696, n3697,
    n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721,
    n3722, n3723, n3724, n3725, n3726, n3727,
    n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751,
    n3752, n3753, n3754, n3755, n3756, n3757,
    n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775,
    n3776, n3777, n3778, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787,
    n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805,
    n3806, n3807, n3808, n3809, n3810, n3811,
    n3812, n3813, n3814, n3815, n3816, n3817,
    n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835,
    n3836, n3837, n3838, n3839, n3840, n3841,
    n3842, n3843, n3844, n3845, n3846, n3847,
    n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865,
    n3866, n3867, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877,
    n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901,
    n3902, n3903, n3904, n3905, n3906, n3907,
    n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931,
    n3932, n3933, n3934, n3935, n3936, n3937,
    n3938, n3939, n3940, n3941, n3942, n3943,
    n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961,
    n3962, n3963, n3964, n3965, n3966, n3967,
    n3968, n3969, n3970, n3971, n3972, n3973,
    n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985,
    n3986, n3987, n3988, n3989, n3990, n3991,
    n3992, n3993, n3994, n3995, n3996, n3997,
    n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027,
    n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057,
    n4058, n4059, n4060, n4061, n4062, n4063,
    n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4083, n4084, n4085, n4086, n4087,
    n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4095, n4096, n4097, n4098, n4099,
    n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117,
    n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141,
    n4142, n4143, n4144, n4145, n4146, n4147,
    n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171,
    n4172, n4173, n4174, n4175, n4176, n4177,
    n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188, n4189,
    n4190, n4191, n4192, n4193, n4194, n4195,
    n4196, n4197, n4198, n4199, n4200, n4201,
    n4202, n4203, n4204, n4205, n4206, n4207,
    n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219,
    n4220, n4221, n4222, n4223, n4224, n4225,
    n4226, n4227, n4228, n4229, n4230, n4231,
    n4232, n4233, n4234, n4235, n4236, n4237,
    n4238, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249,
    n4250, n4251, n4252, n4253, n4254, n4255,
    n4256, n4257, n4258, n4259, n4260, n4261,
    n4262, n4263, n4264, n4265, n4266, n4267,
    n4268, n4269, n4270, n4271, n4272, n4273,
    n4274, n4275, n4276, n4277, n4278, n4279,
    n4280, n4281, n4282, n4283, n4284, n4285,
    n4286, n4287, n4288, n4289, n4290, n4291,
    n4292, n4293, n4294, n4295, n4296, n4297,
    n4298, n4299, n4300, n4301, n4302, n4303,
    n4304, n4305, n4306, n4307, n4308, n4309,
    n4310, n4311, n4312, n4313, n4314, n4315,
    n4316, n4317, n4318, n4319, n4320, n4321,
    n4322, n4323, n4324, n4325, n4326, n4327,
    n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339,
    n4340, n4341, n4342, n4343, n4344, n4345,
    n4346, n4347, n4348, n4349, n4350, n4351,
    n4352, n4353, n4354, n4355, n4356, n4357,
    n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4368, n4369,
    n4370, n4371, n4372, n4373, n4374, n4375,
    n4376, n4377, n4378, n4379, n4380, n4381,
    n4382, n4383, n4384, n4385, n4386, n4387,
    n4388, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4396, n4397, n4398, n4399,
    n4400, n4401, n4402, n4403, n4404, n4405,
    n4406, n4407, n4408, n4409, n4410, n4411,
    n4412, n4413, n4414, n4415, n4416, n4417,
    n4418, n4419, n4420, n4421, n4422, n4423,
    n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4432, n4433, n4434, n4435,
    n4436, n4437, n4438, n4439, n4440, n4441,
    n4442, n4443, n4444, n4445, n4446, n4447,
    n4448, n4449, n4450, n4451, n4452, n4453,
    n4454, n4455, n4456, n4457, n4458, n4459,
    n4460, n4461, n4462, n4463, n4464, n4465,
    n4466, n4467, n4468, n4469, n4470, n4471,
    n4472, n4473, n4474, n4475, n4476, n4477,
    n4478, n4479, n4480, n4481, n4482, n4483,
    n4484, n4485, n4486, n4487, n4488, n4489,
    n4490, n4491, n4492, n4493, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501,
    n4502, n4503, n4504, n4505, n4506, n4507,
    n4508, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525,
    n4526, n4527, n4528, n4529, n4530, n4531,
    n4532, n4533, n4534, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747,
    n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837,
    n4838, n4839, n4840, n4841, n4842, n4843,
    n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861,
    n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873,
    n4874, n4875, n4876, n4877, n4878, n4879,
    n4880, n4881, n4882, n4883, n4884, n4885,
    n4886, n4887, n4888, n4889, n4890, n4891,
    n4892, n4893, n4894, n4895, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101,
    n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5122, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131,
    n5132, n5133, n5134, n5135, n5136, n5137,
    n5138, n5139, n5140, n5141, n5142, n5143,
    n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161,
    n5162, n5163, n5164, n5165, n5166, n5167,
    n5168, n5169, n5170, n5171, n5172, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179,
    n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191,
    n5192, n5193, n5194, n5195, n5196, n5197,
    n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5205, n5206, n5207, n5208, n5209,
    n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221,
    n5222, n5223, n5224, n5225, n5226, n5227,
    n5228, n5229, n5230, n5231, n5232, n5233,
    n5234, n5235, n5236, n5237, n5238, n5239,
    n5240, n5241, n5242, n5243, n5244, n5245,
    n5246, n5247, n5248, n5249, n5250, n5251,
    n5252, n5253, n5254, n5255, n5256, n5257,
    n5258, n5259, n5260, n5261, n5262, n5263,
    n5264, n5265, n5266, n5267, n5268, n5269,
    n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281,
    n5282, n5283, n5284, n5285, n5286, n5287,
    n5288, n5289, n5290, n5291, n5292, n5293,
    n5294, n5295, n5296, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305,
    n5306, n5307, n5308, n5309, n5310, n5311,
    n5312, n5313, n5314, n5315, n5316, n5317,
    n5318, n5319, n5320, n5321, n5322, n5323,
    n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5333, n5334, n5335,
    n5336, n5337, n5338, n5339, n5340, n5341,
    n5342, n5343, n5344, n5345, n5346, n5347,
    n5348, n5349, n5350, n5351, n5352, n5353,
    n5354, n5355, n5356, n5357, n5358, n5359,
    n5360, n5361, n5362, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371,
    n5372, n5373, n5374, n5375, n5376, n5377,
    n5378, n5379, n5380, n5381, n5382, n5383,
    n5384, n5385, n5386, n5387, n5388, n5389,
    n5390, n5391, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401,
    n5402, n5403, n5404, n5405, n5406, n5407,
    n5408, n5409, n5410, n5411, n5412, n5413,
    n5414, n5415, n5416, n5417, n5418, n5419,
    n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431,
    n5432, n5433, n5434, n5435, n5436, n5437,
    n5438, n5439, n5440, n5441, n5442, n5443,
    n5444, n5445, n5446, n5447, n5448, n5449,
    n5450, n5451, n5452, n5453, n5454, n5455,
    n5456, n5457, n5458, n5459, n5460, n5461,
    n5462, n5463, n5464, n5465, n5466, n5467,
    n5468, n5469, n5470, n5471, n5472, n5473,
    n5474, n5475, n5476, n5477, n5478, n5479,
    n5480, n5481, n5482, n5483, n5484, n5485,
    n5486, n5487, n5488, n5489, n5490, n5491,
    n5492, n5493, n5494, n5495, n5496, n5497,
    n5498, n5499, n5500, n5501, n5502, n5503,
    n5504, n5505, n5506, n5507, n5508, n5509,
    n5510, n5511, n5512, n5513, n5514, n5515,
    n5516, n5517, n5518, n5519, n5520, n5521,
    n5522, n5523, n5524, n5525, n5526, n5527,
    n5528, n5529, n5530, n5531, n5532, n5533,
    n5534, n5535, n5536, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551,
    n5552, n5553, n5554, n5555, n5556, n5557,
    n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581,
    n5582, n5583, n5584, n5585, n5586, n5587,
    n5588, n5589, n5590, n5591, n5592, n5593,
    n5594, n5595, n5596, n5597, n5598, n5599,
    n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611,
    n5612, n5613, n5614, n5615, n5616, n5617,
    n5618, n5619, n5620, n5621, n5622, n5623,
    n5624, n5625, n5626, n5627, n5628, n5629,
    n5630, n5631, n5632, n5633, n5634, n5635,
    n5636, n5637, n5638, n5639, n5640, n5641,
    n5642, n5643, n5644, n5645, n5646, n5647,
    n5648, n5649, n5650, n5651, n5652, n5653,
    n5654, n5655, n5656, n5657, n5658, n5659,
    n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5667, n5668, n5669, n5670, n5671,
    n5672, n5673, n5674, n5675, n5676, n5677,
    n5678, n5679, n5680, n5681, n5682, n5683,
    n5684, n5685, n5686, n5687, n5688, n5689,
    n5690, n5691, n5692, n5693, n5694, n5695,
    n5696, n5697, n5698, n5699, n5700, n5701,
    n5702, n5703, n5704, n5705, n5706, n5707,
    n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5715, n5716, n5717, n5718, n5719,
    n5720, n5721, n5722, n5723, n5724, n5725,
    n5726, n5727, n5728, n5729, n5730, n5731,
    n5732, n5733, n5734, n5735, n5736, n5737,
    n5738, n5739, n5740, n5741, n5742, n5743,
    n5744, n5745, n5746, n5747, n5748, n5749,
    n5750, n5751, n5752, n5753, n5754, n5755,
    n5756, n5757, n5758, n5759, n5760, n5761,
    n5762, n5763, n5764, n5765, n5766, n5767,
    n5768, n5769, n5770, n5771, n5772, n5773,
    n5774, n5775, n5776, n5777, n5778, n5779,
    n5780, n5781, n5782, n5783, n5784, n5785,
    n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5794, n5795, n5796, n5797,
    n5798, n5799, n5800, n5801, n5802, n5803,
    n5804, n5805, n5806, n5807, n5808, n5809,
    n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5817, n5818, n5819, n5820, n5821,
    n5822, n5823, n5824, n5825, n5826, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833,
    n5834, n5835, n5836, n5837, n5838, n5839,
    n5840, n5841, n5842, n5843, n5844, n5845,
    n5846, n5847, n5848, n5849, n5850, n5851,
    n5852, n5853, n5854, n5855, n5856, n5857,
    n5858, n5859, n5860, n5861, n5862, n5863,
    n5864, n5865, n5866, n5867, n5868, n5869,
    n5870, n5871, n5872, n5873, n5874, n5875,
    n5876, n5877, n5878, n5879, n5880, n5881,
    n5882, n5883, n5884, n5885, n5886, n5887,
    n5888, n5889, n5890, n5891, n5892, n5893,
    n5894, n5895, n5896, n5897, n5898, n5899,
    n5900, n5901, n5902, n5903, n5904, n5905,
    n5906, n5907, n5908, n5909, n5910, n5911,
    n5912, n5913, n5914, n5915, n5916, n5917,
    n5918, n5919, n5920, n5921, n5922, n5923,
    n5924, n5925, n5926, n5927, n5928, n5929,
    n5930, n5931, n5932, n5933, n5934, n5935,
    n5936, n5937, n5938, n5939, n5940, n5941,
    n5942, n5943, n5944, n5945, n5946, n5947,
    n5948, n5949, n5950, n5951, n5952, n5953,
    n5954, n5955, n5956, n5957, n5958, n5959,
    n5960, n5961, n5962, n5963, n5964, n5965,
    n5966, n5967, n5968, n5969, n5970, n5971,
    n5972, n5973, n5974, n5975, n5976, n5977,
    n5978, n5979, n5980, n5981, n5982, n5983,
    n5984, n5985, n5986, n5987, n5988, n5989,
    n5990, n5991, n5992, n5993, n5994, n5995,
    n5996, n5997, n5998, n5999, n6000, n6001,
    n6002, n6003, n6004, n6005, n6006, n6007,
    n6008, n6009, n6010, n6011, n6012, n6013,
    n6014, n6015, n6016, n6017, n6018, n6019,
    n6020, n6021, n6022, n6023, n6024, n6025,
    n6026, n6027, n6028, n6029, n6030, n6031,
    n6032, n6033, n6034, n6035, n6036, n6037,
    n6038, n6039, n6040, n6041, n6042, n6043,
    n6044, n6045, n6046, n6047, n6048, n6049,
    n6050, n6051, n6052, n6053, n6054, n6055,
    n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067,
    n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079,
    n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097,
    n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6126, n6127,
    n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145,
    n6146, n6147, n6148, n6149, n6150, n6151,
    n6152, n6153, n6154, n6155, n6156, n6157,
    n6158, n6159, n6160, n6161, n6162, n6163,
    n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175,
    n6176, n6177, n6178, n6179, n6180, n6181,
    n6182, n6183, n6184, n6185, n6186, n6187,
    n6188, n6189, n6190, n6191, n6192, n6193,
    n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6202, n6203, n6204, n6205,
    n6206, n6207, n6208, n6209, n6210, n6211,
    n6212, n6213, n6214, n6215, n6216, n6217,
    n6218, n6219, n6220, n6221, n6222, n6223,
    n6224, n6225, n6226, n6227, n6228, n6229,
    n6230, n6231, n6232, n6233, n6234, n6235,
    n6236, n6237, n6238, n6239, n6240, n6241,
    n6242, n6243, n6244, n6245, n6246, n6247,
    n6248, n6249, n6250, n6251, n6252, n6253,
    n6254, n6255, n6256, n6257, n6258, n6259,
    n6260, n6261, n6262, n6263, n6264, n6265,
    n6266, n6267, n6268, n6269, n6270, n6271,
    n6272, n6273, n6274, n6275, n6276, n6277,
    n6278, n6279, n6280, n6281, n6282, n6283,
    n6284, n6285, n6286, n6287, n6288, n6289,
    n6290, n6291, n6292, n6293, n6294, n6295,
    n6296, n6297, n6298, n6299, n6300, n6301,
    n6302, n6303, n6305, n6306, n6307, n6308,
    n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326,
    n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6360, n6361, n6362,
    n6363, n6364, n6365, n6366, n6367, n6368,
    n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386,
    n6387, n6388, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398,
    n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6416, n6417,
    n6418, n6419, n6420, n6421, n6422, n6423,
    n6424, n6425, n6426, n6427, n6428, n6429,
    n6430, n6431, n6432, n6433, n6434, n6435,
    n6436, n6437, n6438, n6439, n6440, n6441,
    n6442, n6443, n6444, n6445, n6446, n6447,
    n6448, n6449, n6450, n6451, n6452, n6453,
    n6454, n6455, n6456, n6457, n6458, n6459,
    n6460, n6461, n6462, n6463, n6464, n6465,
    n6466, n6467, n6468, n6469, n6470, n6471,
    n6472, n6473, n6474, n6475, n6476, n6477,
    n6478, n6479, n6480, n6481, n6482, n6483,
    n6484, n6485, n6486, n6487, n6488, n6489,
    n6490, n6491, n6492, n6493, n6494, n6495,
    n6496, n6497, n6498, n6499, n6500, n6501,
    n6502, n6503, n6504, n6505, n6506, n6507,
    n6508, n6509, n6510, n6511, n6512, n6513,
    n6514, n6515, n6516, n6517, n6518, n6519,
    n6520, n6521, n6522, n6523, n6524, n6525,
    n6526, n6527, n6528, n6529, n6530, n6531,
    n6532, n6533, n6534, n6535, n6536, n6537,
    n6538, n6539, n6540, n6541, n6542, n6543,
    n6544, n6545, n6546, n6547, n6548, n6549,
    n6550, n6551, n6552, n6553, n6554, n6555,
    n6556, n6557, n6558, n6559, n6560, n6561,
    n6562, n6563, n6564, n6565, n6566, n6567,
    n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579,
    n6580, n6581, n6582, n6583, n6584, n6585,
    n6586, n6587, n6588, n6589, n6590, n6591,
    n6592, n6593, n6594, n6595, n6596, n6597,
    n6598, n6599, n6600, n6601, n6602, n6603,
    n6604, n6605, n6606, n6607, n6608, n6609,
    n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621,
    n6622, n6623, n6624, n6625, n6626, n6627,
    n6628, n6629, n6630, n6631, n6632, n6633,
    n6634, n6635, n6636, n6637, n6638, n6639,
    n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651,
    n6652, n6653, n6654, n6655, n6656, n6657,
    n6658, n6659, n6660, n6661, n6662, n6663,
    n6664, n6665, n6666, n6667, n6668, n6669,
    n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6680, n6681,
    n6682, n6683, n6684, n6685, n6686, n6687,
    n6688, n6689, n6690, n6691, n6692, n6693,
    n6694, n6695, n6696, n6697, n6698, n6699,
    n6700, n6701, n6702, n6703, n6704, n6705,
    n6706, n6707, n6708, n6709, n6710, n6711,
    n6712, n6713, n6714, n6715, n6716, n6717,
    n6718, n6719, n6720, n6721, n6722, n6723,
    n6724, n6725, n6726, n6727, n6728, n6729,
    n6730, n6731, n6732, n6733, n6734, n6735,
    n6736, n6737, n6738, n6739, n6740, n6741,
    n6742, n6743, n6744, n6745, n6746, n6747,
    n6748, n6749, n6750, n6751, n6752, n6753,
    n6754, n6755, n6756, n6757, n6758, n6759,
    n6760, n6761, n6762, n6763, n6764, n6765,
    n6766, n6767, n6768, n6769, n6770, n6771,
    n6772, n6773, n6774, n6775, n6776, n6777,
    n6778, n6779, n6780, n6781, n6782, n6783,
    n6784, n6785, n6786, n6787, n6788, n6789,
    n6790, n6791, n6792, n6793, n6794, n6795,
    n6796, n6797, n6798, n6799, n6800, n6801,
    n6802, n6803, n6804, n6805, n6806, n6807,
    n6808, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831,
    n6832, n6833, n6834, n6835, n6836, n6837,
    n6838, n6839, n6840, n6841, n6842, n6843,
    n6844, n6845, n6846, n6847, n6848, n6849,
    n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861,
    n6862, n6863, n6864, n6865, n6866, n6867,
    n6868, n6869, n6870, n6871, n6872, n6873,
    n6874, n6875, n6876, n6877, n6878, n6879,
    n6880, n6881, n6882, n6883, n6884, n6885,
    n6886, n6887, n6888, n6889, n6890, n6891,
    n6892, n6893, n6894, n6895, n6896, n6897,
    n6898, n6899, n6900, n6901, n6902, n6903,
    n6904, n6905, n6906, n6907, n6908, n6909,
    n6910, n6911, n6912, n6913, n6914, n6915,
    n6916, n6917, n6918, n6919, n6920, n6921,
    n6922, n6923, n6924, n6925, n6926, n6927,
    n6928, n6929, n6930, n6931, n6932, n6933,
    n6934, n6935, n6936, n6937, n6938, n6939,
    n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951,
    n6952, n6953, n6954, n6955, n6956, n6957,
    n6958, n6959, n6960, n6961, n6962, n6963,
    n6964, n6965, n6966, n6967, n6968, n6969,
    n6970, n6971, n6972, n6973, n6974, n6975,
    n6976, n6977, n6978, n6979, n6980, n6981,
    n6982, n6983, n6984, n6985, n6986, n6987,
    n6988, n6989, n6990, n6991, n6992, n6993,
    n6994, n6995, n6996, n6997, n6998, n6999,
    n7000, n7001, n7002, n7003, n7004, n7005,
    n7006, n7007, n7008, n7009, n7010, n7011,
    n7012, n7013, n7014, n7015, n7016, n7017,
    n7018, n7019, n7020, n7021, n7022, n7023,
    n7024, n7025, n7026, n7027, n7028, n7029,
    n7030, n7031, n7032, n7033, n7034, n7035,
    n7036, n7037, n7038, n7039, n7040, n7041,
    n7042, n7043, n7044, n7045, n7046, n7047,
    n7048, n7049, n7050, n7051, n7052, n7053,
    n7054, n7055, n7056, n7057, n7058, n7059,
    n7060, n7061, n7062, n7063, n7064, n7065,
    n7066, n7067, n7068, n7069, n7070, n7071,
    n7072, n7073, n7074, n7075, n7076, n7077,
    n7078, n7079, n7080, n7081, n7082, n7083,
    n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095,
    n7096, n7097, n7098, n7099, n7100, n7101,
    n7102, n7103, n7104, n7105, n7106, n7107,
    n7108, n7109, n7110, n7111, n7112, n7113,
    n7114, n7115, n7116, n7117, n7118, n7119,
    n7120, n7121, n7122, n7123, n7124, n7125,
    n7126, n7127, n7128, n7129, n7130, n7131,
    n7132, n7133, n7134, n7135, n7136, n7137,
    n7138, n7139, n7140, n7141, n7142, n7143,
    n7144, n7145, n7146, n7147, n7148, n7149,
    n7150, n7151, n7152, n7153, n7154, n7155,
    n7156, n7157, n7158, n7159, n7160, n7161,
    n7162, n7163, n7164, n7165, n7166, n7167,
    n7168, n7169, n7170, n7171, n7172, n7173,
    n7174, n7175, n7176, n7177, n7178, n7179,
    n7180, n7181, n7182, n7183, n7184, n7185,
    n7186, n7187, n7188, n7189, n7190, n7191,
    n7192, n7193, n7194, n7195, n7196, n7197,
    n7198, n7199, n7200, n7201, n7202, n7203,
    n7204, n7205, n7206, n7207, n7208, n7209,
    n7210, n7211, n7212, n7213, n7214, n7215,
    n7216, n7217, n7218, n7219, n7220, n7221,
    n7222, n7223, n7224, n7225, n7226, n7227,
    n7228, n7229, n7230, n7231, n7232, n7233,
    n7234, n7235, n7236, n7237, n7238, n7239,
    n7240, n7241, n7242, n7243, n7244, n7245,
    n7246, n7247, n7248, n7249, n7250, n7251,
    n7252, n7253, n7254, n7255, n7256, n7257,
    n7258, n7259, n7260, n7261, n7262, n7263,
    n7264, n7265, n7266, n7267, n7268, n7269,
    n7270, n7271, n7272, n7273, n7274, n7275,
    n7276, n7277, n7278, n7279, n7280, n7281,
    n7282, n7283, n7284, n7285, n7286, n7287,
    n7288, n7289, n7290, n7291, n7292, n7293,
    n7294, n7295, n7296, n7297, n7298, n7299,
    n7300, n7301, n7302, n7303, n7304, n7305,
    n7306, n7307, n7308, n7309, n7310, n7311,
    n7312, n7313, n7314, n7315, n7316, n7317,
    n7318, n7319, n7320, n7321, n7322, n7323,
    n7324, n7325, n7326, n7327, n7328, n7329,
    n7330, n7331, n7332, n7333, n7334, n7335,
    n7336, n7337, n7338, n7339, n7340, n7341,
    n7342, n7343, n7344, n7345, n7346, n7347,
    n7348, n7349, n7350, n7351, n7352, n7353,
    n7354, n7355, n7356, n7357, n7358, n7359,
    n7360, n7361, n7362, n7363, n7364, n7365,
    n7366, n7367, n7368, n7369, n7370, n7371,
    n7372, n7373, n7374, n7375, n7376, n7377,
    n7378, n7379, n7380, n7381, n7382, n7383,
    n7384, n7385, n7386, n7387, n7388, n7389,
    n7390, n7391, n7392, n7393, n7394, n7395,
    n7396, n7397, n7398, n7399, n7400, n7401,
    n7402, n7403, n7404, n7405, n7406, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431,
    n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443,
    n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7461,
    n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473,
    n7474, n7475, n7476, n7477, n7478, n7479,
    n7480, n7481, n7482, n7483, n7484, n7485,
    n7486, n7487, n7488, n7489, n7490, n7491,
    n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503,
    n7504, n7505, n7506, n7507, n7508, n7509,
    n7510, n7511, n7512, n7513, n7514, n7515,
    n7516, n7517, n7518, n7519, n7520, n7521,
    n7522, n7523, n7524, n7525, n7526, n7527,
    n7528, n7529, n7530, n7531, n7532, n7533,
    n7534, n7535, n7536, n7537, n7538, n7539,
    n7540, n7541, n7542, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551,
    n7552, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563,
    n7564, n7565, n7566, n7567, n7568, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581,
    n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611,
    n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653,
    n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683,
    n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713,
    n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7721, n7722, n7723, n7724, n7725,
    n7726, n7727, n7728, n7729, n7730, n7731,
    n7732, n7733, n7734, n7735, n7736, n7737,
    n7738, n7739, n7740, n7741, n7742, n7743,
    n7744, n7745, n7746, n7747, n7748, n7749,
    n7750, n7751, n7752, n7753, n7754, n7755,
    n7756, n7757, n7758, n7759, n7760, n7761,
    n7762, n7763, n7764, n7765, n7766, n7767,
    n7768, n7769, n7770, n7771, n7772, n7773,
    n7774, n7775, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785,
    n7786, n7787, n7788, n7789, n7790, n7791,
    n7792, n7793, n7794, n7795, n7796, n7797,
    n7798, n7799, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821,
    n7822, n7823, n7824, n7825, n7826, n7827,
    n7828, n7829, n7830, n7831, n7832, n7833,
    n7834, n7835, n7836, n7837, n7838, n7839,
    n7840, n7841, n7842, n7843, n7844, n7845,
    n7846, n7847, n7848, n7849, n7850, n7851,
    n7852, n7853, n7854, n7855, n7856, n7857,
    n7858, n7859, n7860, n7861, n7862, n7863,
    n7864, n7865, n7866, n7867, n7868, n7869,
    n7870, n7871, n7872, n7873, n7874, n7875,
    n7876, n7877, n7878, n7879, n7880, n7881,
    n7882, n7883, n7884, n7885, n7886, n7887,
    n7888, n7889, n7890, n7891, n7892, n7893,
    n7894, n7895, n7896, n7897, n7898, n7899,
    n7900, n7901, n7902, n7903, n7904, n7905,
    n7906, n7907, n7908, n7909, n7910, n7911,
    n7912, n7913, n7914, n7915, n7916, n7917,
    n7918, n7919, n7920, n7921, n7922, n7923,
    n7924, n7925, n7926, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935,
    n7936, n7937, n7938, n7939, n7940, n7941,
    n7942, n7943, n7944, n7945, n7946, n7947,
    n7948, n7949, n7950, n7951, n7952, n7953,
    n7954, n7955, n7956, n7957, n7958, n7959,
    n7960, n7961, n7962, n7963, n7964, n7965,
    n7966, n7967, n7968, n7969, n7970, n7971,
    n7972, n7973, n7974, n7975, n7976, n7977,
    n7978, n7979, n7980, n7981, n7982, n7983,
    n7984, n7985, n7986, n7987, n7988, n7989,
    n7990, n7991, n7992, n7993, n7994, n7995,
    n7996, n7997, n7998, n7999, n8000, n8001,
    n8002, n8003, n8004, n8005, n8006, n8007,
    n8008, n8009, n8010, n8011, n8012, n8013,
    n8014, n8015, n8016, n8017, n8018, n8019,
    n8020, n8021, n8022, n8023, n8024, n8025,
    n8026, n8027, n8028, n8029, n8030, n8031,
    n8032, n8033, n8034, n8035, n8036, n8037,
    n8038, n8039, n8040, n8041, n8042, n8043,
    n8044, n8045, n8046, n8047, n8048, n8049,
    n8050, n8051, n8052, n8053, n8054, n8055,
    n8056, n8057, n8058, n8059, n8060, n8061,
    n8062, n8063, n8064, n8065, n8066, n8067,
    n8068, n8069, n8070, n8071, n8072, n8073,
    n8074, n8075, n8076, n8077, n8078, n8079,
    n8080, n8081, n8082, n8083, n8084, n8085,
    n8086, n8087, n8088, n8089, n8090, n8091,
    n8092, n8093, n8094, n8095, n8096, n8097,
    n8098, n8099, n8100, n8101, n8102, n8103,
    n8104, n8105, n8106, n8107, n8108, n8109,
    n8110, n8111, n8112, n8113, n8114, n8115,
    n8116, n8117, n8118, n8119, n8120, n8121,
    n8122, n8123, n8124, n8125, n8126, n8127,
    n8128, n8129, n8130, n8131, n8132, n8133,
    n8134, n8135, n8136, n8137, n8138, n8139,
    n8140, n8141, n8142, n8143, n8144, n8145,
    n8146, n8147, n8148, n8149, n8150, n8151,
    n8152, n8153, n8154, n8155, n8156, n8157,
    n8158, n8159, n8160, n8161, n8162, n8163,
    n8164, n8165, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176,
    n8177, n8178, n8179, n8180, n8181, n8182,
    n8183, n8184, n8185, n8186, n8187, n8188,
    n8189, n8190, n8191, n8192, n8193, n8194,
    n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206,
    n8207, n8208, n8209, n8210, n8211, n8212,
    n8213, n8214, n8215, n8216, n8217, n8218,
    n8219, n8220, n8221, n8222, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236,
    n8237, n8238, n8239, n8240, n8241, n8242,
    n8243, n8244, n8245, n8246, n8247, n8248,
    n8249, n8250, n8251, n8252, n8253, n8254,
    n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266,
    n8267, n8268, n8269, n8270, n8271, n8272,
    n8273, n8274, n8275, n8276, n8277, n8278,
    n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296,
    n8297, n8298, n8299, n8300, n8301, n8302,
    n8303, n8304, n8305, n8306, n8307, n8308,
    n8309, n8310, n8311, n8312, n8313, n8314,
    n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326,
    n8327, n8328, n8329, n8330, n8331, n8332,
    n8333, n8334, n8335, n8336, n8337, n8338,
    n8339, n8340, n8341, n8342, n8343, n8344,
    n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356,
    n8357, n8358, n8359, n8360, n8361, n8362,
    n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8370, n8371, n8372, n8373, n8374,
    n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386,
    n8387, n8388, n8389, n8390, n8391, n8392,
    n8393, n8394, n8395, n8396, n8397, n8398,
    n8399, n8400, n8401, n8402, n8403, n8404,
    n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8414, n8415, n8416,
    n8417, n8418, n8419, n8420, n8421, n8422,
    n8423, n8424, n8425, n8426, n8427, n8428,
    n8429, n8430, n8431, n8432, n8433, n8434,
    n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446,
    n8447, n8448, n8449, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8463, n8464,
    n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476,
    n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494,
    n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8505, n8506,
    n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518,
    n8519, n8520, n8521, n8522, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530,
    n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548,
    n8549, n8550, n8551, n8552, n8553, n8554,
    n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8564, n8565, n8566,
    n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590,
    n8591, n8592, n8593, n8594, n8595, n8596,
    n8597, n8598, n8599, n8600, n8601, n8602,
    n8603, n8604, n8605, n8606, n8607, n8608,
    n8609, n8610, n8611, n8612, n8613, n8614,
    n8615, n8616, n8617, n8618, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626,
    n8627, n8628, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8636, n8637, n8638,
    n8639, n8640, n8641, n8642, n8643, n8644,
    n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656,
    n8657, n8658, n8659, n8660, n8661, n8662,
    n8663, n8664, n8665, n8666, n8667, n8668,
    n8669, n8670, n8671, n8672, n8673, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686,
    n8687, n8688, n8689, n8690, n8691, n8692,
    n8693, n8694, n8695, n8696, n8697, n8698,
    n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722,
    n8723, n8724, n8725, n8726, n8727, n8728,
    n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746,
    n8747, n8748, n8749, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8757, n8758,
    n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776,
    n8777, n8778, n8780, n8781, n8782, n8783,
    n8784, n8785, n8786, n8787, n8788, n8789,
    n8790, n8791, n8792, n8793, n8794, n8795,
    n8796, n8797, n8798, n8799, n8800, n8801,
    n8802, n8803, n8804, n8805, n8806, n8807,
    n8808, n8809, n8810, n8811, n8812, n8813,
    n8814, n8815, n8816, n8817, n8818, n8819,
    n8820, n8821, n8822, n8823, n8824, n8825,
    n8826, n8827, n8828, n8829, n8830, n8831,
    n8832, n8833, n8834, n8835, n8836, n8837,
    n8838, n8839, n8840, n8841, n8842, n8843,
    n8844, n8845, n8846, n8847, n8848, n8849,
    n8850, n8851, n8852, n8853, n8854, n8855,
    n8856, n8857, n8858, n8859, n8860, n8861,
    n8862, n8863, n8864, n8865, n8866, n8867,
    n8868, n8869, n8870, n8871, n8872, n8873,
    n8874, n8875, n8876, n8877, n8878, n8879,
    n8880, n8881, n8882, n8883, n8884, n8885,
    n8886, n8887, n8888, n8889, n8890, n8891,
    n8892, n8893, n8894, n8895, n8896, n8897,
    n8898, n8899, n8900, n8901, n8902, n8903,
    n8904, n8905, n8906, n8907, n8908, n8909,
    n8910, n8911, n8912, n8913, n8914, n8915,
    n8916, n8917, n8918, n8919, n8920, n8921,
    n8922, n8923, n8924, n8925, n8926, n8927,
    n8928, n8929, n8930, n8931, n8932, n8933,
    n8934, n8935, n8936, n8937, n8938, n8939,
    n8940, n8941, n8942, n8943, n8944, n8945,
    n8946, n8947, n8948, n8949, n8950, n8951,
    n8952, n8953, n8954, n8955, n8956, n8957,
    n8958, n8959, n8960, n8961, n8962, n8963,
    n8964, n8965, n8966, n8967, n8968, n8969,
    n8970, n8971, n8972, n8973, n8974, n8975,
    n8976, n8977, n8978, n8979, n8980, n8981,
    n8982, n8983, n8984, n8985, n8986, n8987,
    n8988, n8989, n8990, n8991, n8992, n8993,
    n8994, n8995, n8996, n8997, n8998, n8999,
    n9000, n9001, n9002, n9003, n9004, n9005,
    n9006, n9007, n9008, n9009, n9010, n9011,
    n9012, n9013, n9014, n9015, n9016, n9017,
    n9018, n9019, n9020, n9021, n9022, n9023,
    n9024, n9025, n9026, n9027, n9028, n9029,
    n9030, n9031, n9032, n9033, n9034, n9035,
    n9036, n9037, n9038, n9039, n9040, n9041,
    n9042, n9043, n9044, n9045, n9046, n9047,
    n9048, n9049, n9050, n9051, n9052, n9053,
    n9054, n9055, n9056, n9057, n9058, n9059,
    n9060, n9061, n9062, n9063, n9064, n9065,
    n9066, n9067, n9068, n9069, n9070, n9071,
    n9072, n9073, n9074, n9075, n9076, n9077,
    n9078, n9079, n9080, n9081, n9082, n9083,
    n9084, n9085, n9086, n9087, n9088, n9089,
    n9090, n9091, n9092, n9093, n9094, n9095,
    n9096, n9097, n9098, n9099, n9100, n9101,
    n9102, n9103, n9104, n9105, n9106, n9107,
    n9108, n9109, n9110, n9111, n9112, n9113,
    n9114, n9115, n9116, n9117, n9118, n9119,
    n9120, n9121, n9122, n9123, n9124, n9125,
    n9126, n9127, n9128, n9129, n9130, n9131,
    n9132, n9133, n9134, n9135, n9136, n9137,
    n9138, n9139, n9140, n9141, n9142, n9143,
    n9144, n9145, n9146, n9147, n9148, n9149,
    n9150, n9151, n9152, n9153, n9154, n9155,
    n9156, n9157, n9158, n9159, n9160, n9161,
    n9162, n9163, n9164, n9165, n9166, n9167,
    n9168, n9169, n9170, n9171, n9172, n9173,
    n9174, n9175, n9176, n9177, n9178, n9179,
    n9180, n9181, n9182, n9183, n9184, n9185,
    n9186, n9187, n9188, n9189, n9190, n9191,
    n9192, n9193, n9194, n9195, n9196, n9197,
    n9198, n9199, n9200, n9201, n9202, n9203,
    n9204, n9205, n9206, n9207, n9208, n9209,
    n9210, n9211, n9212, n9213, n9214, n9215,
    n9216, n9217, n9218, n9219, n9220, n9221,
    n9222, n9223, n9224, n9225, n9226, n9227,
    n9228, n9229, n9230, n9231, n9232, n9233,
    n9234, n9235, n9236, n9237, n9238, n9239,
    n9240, n9241, n9242, n9243, n9244, n9245,
    n9246, n9247, n9248, n9249, n9250, n9251,
    n9252, n9253, n9254, n9255, n9256, n9257,
    n9258, n9259, n9260, n9261, n9262, n9263,
    n9264, n9265, n9266, n9267, n9268, n9269,
    n9270, n9271, n9272, n9273, n9274, n9275,
    n9276, n9277, n9278, n9279, n9280, n9281,
    n9282, n9283, n9284, n9285, n9286, n9287,
    n9288, n9289, n9290, n9291, n9292, n9293,
    n9294, n9295, n9296, n9297, n9298, n9299,
    n9300, n9301, n9302, n9303, n9304, n9305,
    n9306, n9307, n9308, n9309, n9310, n9311,
    n9312, n9313, n9314, n9315, n9316, n9317,
    n9318, n9319, n9320, n9321, n9322, n9323,
    n9324, n9325, n9326, n9327, n9328, n9329,
    n9330, n9331, n9332, n9333, n9334, n9335,
    n9336, n9337, n9338, n9339, n9340, n9341,
    n9342, n9343, n9344, n9345, n9346, n9347,
    n9348, n9349, n9350, n9351, n9352, n9353,
    n9354, n9355, n9356, n9357, n9358, n9359,
    n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9370, n9371,
    n9372, n9373, n9374, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9382, n9383,
    n9384, n9385, n9386, n9387, n9388, n9389,
    n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401,
    n9402, n9403, n9404, n9405, n9406, n9407,
    n9408, n9409, n9410, n9411, n9412, n9413,
    n9414, n9415, n9416, n9417, n9418, n9419,
    n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431,
    n9432, n9433, n9434, n9435, n9436, n9437,
    n9438, n9439, n9440, n9441, n9442, n9443,
    n9444, n9445, n9446, n9447, n9448, n9449,
    n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461,
    n9462, n9463, n9464, n9465, n9466, n9467,
    n9468, n9469, n9470, n9471, n9472, n9473,
    n9474, n9475, n9476, n9477, n9478, n9479,
    n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491,
    n9492, n9493, n9494, n9495, n9496, n9497,
    n9498, n9499, n9500, n9501, n9502, n9503,
    n9504, n9505, n9506, n9507, n9508, n9509,
    n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521,
    n9522, n9523, n9524, n9525, n9526, n9527,
    n9528, n9529, n9530, n9531, n9532, n9533,
    n9534, n9535, n9536, n9537, n9538, n9539,
    n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9547, n9548, n9549, n9550, n9551,
    n9552, n9553, n9554, n9555, n9556, n9557,
    n9558, n9559, n9560, n9561, n9562, n9563,
    n9564, n9565, n9566, n9567, n9568, n9569,
    n9570, n9571, n9572, n9573, n9574, n9575,
    n9576, n9577, n9578, n9579, n9580, n9581,
    n9582, n9583, n9584, n9585, n9586, n9587,
    n9588, n9589, n9590, n9591, n9592, n9593,
    n9594, n9595, n9596, n9597, n9598, n9599,
    n9600, n9601, n9602, n9603, n9604, n9605,
    n9606, n9607, n9608, n9609, n9610, n9611,
    n9612, n9613, n9614, n9615, n9616, n9617,
    n9618, n9619, n9620, n9621, n9622, n9623,
    n9624, n9625, n9626, n9627, n9628, n9629,
    n9630, n9631, n9632, n9633, n9634, n9635,
    n9636, n9637, n9638, n9639, n9640, n9641,
    n9642, n9643, n9644, n9645, n9646, n9647,
    n9648, n9649, n9650, n9651, n9652, n9653,
    n9654, n9655, n9656, n9657, n9658, n9659,
    n9660, n9661, n9662, n9663, n9664, n9665,
    n9666, n9667, n9668, n9669, n9670, n9671,
    n9672, n9673, n9674, n9675, n9676, n9677,
    n9678, n9679, n9680, n9681, n9682, n9683,
    n9684, n9685, n9686, n9687, n9688, n9689,
    n9690, n9691, n9692, n9693, n9694, n9695,
    n9696, n9697, n9698, n9699, n9700, n9701,
    n9702, n9703, n9704, n9705, n9706, n9707,
    n9708, n9709, n9710, n9711, n9712, n9713,
    n9714, n9715, n9716, n9717, n9718, n9719,
    n9720, n9721, n9722, n9723, n9724, n9725,
    n9726, n9727, n9728, n9729, n9730, n9731,
    n9732, n9733, n9734, n9735, n9736, n9737,
    n9738, n9739, n9740, n9741, n9742, n9743,
    n9744, n9745, n9746, n9747, n9748, n9749,
    n9750, n9751, n9752, n9753, n9754, n9755,
    n9756, n9757, n9758, n9759, n9760, n9761,
    n9762, n9763, n9764, n9765, n9766, n9767,
    n9768, n9769, n9770, n9771, n9772, n9773,
    n9774, n9775, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786,
    n9787, n9788, n9789, n9790, n9791, n9792,
    n9793, n9794, n9795, n9796, n9797, n9798,
    n9799, n9800, n9801, n9802, n9803, n9804,
    n9805, n9806, n9807, n9808, n9809, n9810,
    n9811, n9812, n9813, n9814, n9815, n9816,
    n9817, n9818, n9819, n9820, n9821, n9822,
    n9823, n9824, n9825, n9826, n9827, n9828,
    n9829, n9830, n9831, n9832, n9833, n9834,
    n9835, n9836, n9837, n9838, n9839, n9840,
    n9841, n9842, n9843, n9844, n9845, n9846,
    n9847, n9848, n9849, n9850, n9851, n9852,
    n9853, n9854, n9855, n9856, n9857, n9858,
    n9859, n9860, n9861, n9862, n9863, n9864,
    n9865, n9866, n9867, n9868, n9869, n9870,
    n9871, n9872, n9873, n9874, n9875, n9876,
    n9877, n9878, n9879, n9880, n9881, n9882,
    n9883, n9884, n9885, n9886, n9887, n9888,
    n9889, n9890, n9891, n9892, n9893, n9894,
    n9895, n9896, n9897, n9898, n9899, n9900,
    n9901, n9902, n9903, n9904, n9905, n9906,
    n9907, n9908, n9909, n9910, n9911, n9912,
    n9913, n9914, n9915, n9916, n9917, n9918,
    n9919, n9920, n9921, n9922, n9923, n9924,
    n9925, n9926, n9927, n9928, n9929, n9930,
    n9931, n9932, n9933, n9934, n9935, n9936,
    n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948,
    n9949, n9950, n9951, n9952, n9953, n9954,
    n9955, n9956, n9957, n9958, n9959, n9960,
    n9961, n9962, n9963, n9964, n9965, n9966,
    n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9990,
    n9991, n9992, n9993, n9994, n9995, n9996,
    n9997, n9998, n9999, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026,
    n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044,
    n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062,
    n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074,
    n10075, n10076, n10077, n10078, n10079, n10080,
    n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092,
    n10093, n10094, n10095, n10096, n10097, n10098,
    n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116,
    n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134,
    n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146,
    n10147, n10148, n10149, n10150, n10151, n10152,
    n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170,
    n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188,
    n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200,
    n10201, n10202, n10203, n10204, n10205, n10206,
    n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218,
    n10219, n10220, n10221, n10222, n10223, n10224,
    n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236,
    n10237, n10238, n10239, n10240, n10241, n10242,
    n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254,
    n10255, n10256, n10257, n10258, n10259, n10260,
    n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272,
    n10273, n10274, n10275, n10276, n10277, n10278,
    n10279, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290,
    n10291, n10292, n10293, n10294, n10295, n10296,
    n10297, n10298, n10299, n10300, n10301, n10302,
    n10303, n10304, n10305, n10306, n10307, n10308,
    n10309, n10310, n10311, n10312, n10313, n10314,
    n10315, n10316, n10317, n10318, n10319, n10320,
    n10321, n10322, n10323, n10324, n10325, n10326,
    n10327, n10328, n10329, n10330, n10331, n10332,
    n10333, n10334, n10335, n10336, n10337, n10338,
    n10339, n10340, n10341, n10342, n10343, n10344,
    n10345, n10346, n10347, n10348, n10349, n10350,
    n10351, n10352, n10353, n10354, n10355, n10356,
    n10357, n10358, n10359, n10360, n10361, n10363,
    n10364, n10365, n10366, n10367, n10368, n10369,
    n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381,
    n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10395, n10396, n10397, n10398, n10399,
    n10400, n10401, n10402, n10403, n10404, n10405,
    n10406, n10407, n10408, n10409, n10410, n10411,
    n10412, n10413, n10414, n10415, n10416, n10417,
    n10418, n10419, n10420, n10421, n10422, n10423,
    n10424, n10425, n10426, n10427, n10428, n10429,
    n10430, n10431, n10432, n10433, n10434, n10435,
    n10436, n10437, n10438, n10439, n10440, n10441,
    n10442, n10443, n10444, n10445, n10446, n10447,
    n10448, n10449, n10450, n10451, n10452, n10453,
    n10454, n10455, n10456, n10457, n10458, n10459,
    n10460, n10461, n10462, n10463, n10464, n10465,
    n10466, n10467, n10468, n10469, n10470, n10471,
    n10472, n10473, n10474, n10475, n10476, n10477,
    n10478, n10479, n10480, n10481, n10482, n10483,
    n10484, n10485, n10486, n10487, n10488, n10489,
    n10490, n10491, n10492, n10493, n10494, n10495,
    n10496, n10497, n10498, n10499, n10500, n10501,
    n10502, n10503, n10504, n10505, n10506, n10507,
    n10508, n10509, n10510, n10511, n10512, n10513,
    n10514, n10515, n10516, n10517, n10518, n10519,
    n10520, n10521, n10522, n10523, n10524, n10525,
    n10526, n10527, n10528, n10529, n10530, n10531,
    n10532, n10533, n10534, n10535, n10536, n10537,
    n10538, n10539, n10540, n10541, n10542, n10543,
    n10544, n10545, n10546, n10547, n10548, n10549,
    n10550, n10551, n10552, n10553, n10554, n10555,
    n10556, n10557, n10558, n10559, n10560, n10561,
    n10562, n10563, n10564, n10565, n10566, n10567,
    n10568, n10569, n10570, n10571, n10572, n10573,
    n10574, n10575, n10576, n10577, n10578, n10579,
    n10580, n10581, n10582, n10583, n10584, n10585,
    n10586, n10587, n10588, n10589, n10590, n10591,
    n10592, n10593, n10594, n10595, n10596, n10597,
    n10598, n10599, n10600, n10601, n10602, n10603,
    n10604, n10605, n10606, n10607, n10608, n10609,
    n10610, n10611, n10612, n10613, n10614, n10615,
    n10616, n10617, n10618, n10619, n10620, n10621,
    n10622, n10623, n10624, n10625, n10626, n10627,
    n10628, n10629, n10630, n10631, n10632, n10633,
    n10634, n10635, n10636, n10637, n10638, n10639,
    n10640, n10641, n10642, n10643, n10644, n10645,
    n10646, n10647, n10648, n10649, n10650, n10651,
    n10652, n10653, n10654, n10655, n10656, n10657,
    n10658, n10659, n10660, n10661, n10662, n10663,
    n10664, n10665, n10666, n10667, n10668, n10669,
    n10670, n10671, n10672, n10673, n10674, n10675,
    n10676, n10677, n10678, n10679, n10680, n10681,
    n10682, n10683, n10684, n10685, n10686, n10687,
    n10688, n10689, n10690, n10691, n10692, n10693,
    n10694, n10695, n10696, n10697, n10698, n10699,
    n10700, n10701, n10702, n10703, n10704, n10705,
    n10706, n10707, n10708, n10709, n10710, n10711,
    n10712, n10713, n10714, n10715, n10716, n10717,
    n10718, n10719, n10720, n10721, n10722, n10723,
    n10724, n10725, n10726, n10727, n10728, n10729,
    n10730, n10731, n10732, n10733, n10734, n10735,
    n10736, n10737, n10738, n10739, n10740, n10741,
    n10742, n10743, n10744, n10745, n10746, n10747,
    n10748, n10749, n10750, n10751, n10752, n10753,
    n10754, n10755, n10756, n10757, n10758, n10759,
    n10760, n10761, n10762, n10763, n10764, n10765,
    n10766, n10767, n10768, n10769, n10770, n10771,
    n10772, n10773, n10774, n10775, n10776, n10777,
    n10778, n10779, n10780, n10781, n10782, n10783,
    n10784, n10785, n10786, n10787, n10788, n10789,
    n10790, n10791, n10792, n10793, n10794, n10795,
    n10796, n10797, n10798, n10799, n10800, n10801,
    n10802, n10803, n10804, n10805, n10806, n10807,
    n10808, n10809, n10810, n10811, n10812, n10813,
    n10814, n10815, n10816, n10817, n10818, n10819,
    n10820, n10821, n10822, n10823, n10824, n10825,
    n10826, n10827, n10828, n10829, n10830, n10831,
    n10832, n10833, n10834, n10835, n10836, n10837,
    n10838, n10839, n10840, n10841, n10842, n10843,
    n10844, n10845, n10846, n10847, n10848, n10849,
    n10850, n10851, n10852, n10853, n10854, n10855,
    n10856, n10857, n10858, n10859, n10860, n10861,
    n10862, n10863, n10864, n10865, n10866, n10867,
    n10868, n10869, n10870, n10871, n10872, n10873,
    n10874, n10875, n10876, n10877, n10878, n10879,
    n10880, n10881, n10882, n10883, n10884, n10885,
    n10886, n10887, n10888, n10889, n10890, n10891,
    n10892, n10893, n10894, n10895, n10896, n10897,
    n10898, n10899, n10900, n10901, n10902, n10903,
    n10904, n10905, n10906, n10907, n10908, n10909,
    n10910, n10911, n10912, n10913, n10914, n10915,
    n10916, n10917, n10918, n10919, n10920, n10921,
    n10922, n10923, n10924, n10925, n10926, n10927,
    n10928, n10929, n10930, n10931, n10932, n10933,
    n10934, n10935, n10936, n10937, n10938, n10939,
    n10940, n10941, n10942, n10943, n10944, n10945,
    n10946, n10947, n10948, n10949, n10950, n10951,
    n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10960, n10961, n10962, n10963, n10964,
    n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10981, n10982,
    n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994,
    n10995, n10996, n10997, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012,
    n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030,
    n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048,
    n11049, n11050, n11051, n11052, n11053, n11054,
    n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066,
    n11067, n11068, n11069, n11070, n11071, n11072,
    n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084,
    n11085, n11086, n11087, n11088, n11089, n11090,
    n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102,
    n11103, n11104, n11105, n11106, n11107, n11108,
    n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120,
    n11121, n11122, n11123, n11124, n11125, n11126,
    n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138,
    n11139, n11140, n11141, n11142, n11143, n11144,
    n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11152, n11153, n11154, n11155, n11156,
    n11157, n11158, n11159, n11160, n11161, n11162,
    n11163, n11164, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174,
    n11175, n11176, n11177, n11178, n11179, n11180,
    n11181, n11182, n11183, n11184, n11185, n11186,
    n11187, n11188, n11189, n11190, n11191, n11192,
    n11193, n11194, n11195, n11196, n11197, n11198,
    n11199, n11200, n11201, n11202, n11203, n11204,
    n11205, n11206, n11207, n11208, n11209, n11210,
    n11211, n11212, n11213, n11214, n11215, n11216,
    n11217, n11218, n11219, n11220, n11221, n11222,
    n11223, n11224, n11225, n11226, n11227, n11228,
    n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240,
    n11241, n11242, n11243, n11244, n11245, n11246,
    n11247, n11248, n11249, n11250, n11251, n11252,
    n11253, n11254, n11255, n11256, n11257, n11258,
    n11259, n11260, n11261, n11262, n11263, n11264,
    n11265, n11266, n11267, n11268, n11269, n11270,
    n11271, n11272, n11273, n11274, n11275, n11276,
    n11277, n11278, n11279, n11280, n11281, n11282,
    n11283, n11284, n11285, n11286, n11287, n11288,
    n11289, n11290, n11291, n11292, n11293, n11294,
    n11295, n11296, n11297, n11298, n11299, n11300,
    n11301, n11302, n11303, n11304, n11305, n11306,
    n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318,
    n11319, n11320, n11321, n11322, n11323, n11324,
    n11325, n11326, n11327, n11328, n11329, n11330,
    n11331, n11332, n11333, n11334, n11335, n11336,
    n11337, n11338, n11339, n11340, n11341, n11342,
    n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11350, n11351, n11352, n11353, n11354,
    n11355, n11356, n11357, n11358, n11359, n11360,
    n11361, n11362, n11363, n11364, n11365, n11366,
    n11367, n11368, n11369, n11370, n11371, n11372,
    n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11386, n11387, n11388, n11389, n11390,
    n11391, n11392, n11393, n11394, n11395, n11396,
    n11397, n11398, n11399, n11400, n11401, n11402,
    n11403, n11404, n11405, n11406, n11407, n11408,
    n11409, n11410, n11411, n11412, n11413, n11414,
    n11415, n11416, n11417, n11418, n11419, n11420,
    n11421, n11422, n11423, n11424, n11425, n11426,
    n11427, n11428, n11429, n11430, n11431, n11432,
    n11433, n11434, n11435, n11436, n11437, n11438,
    n11439, n11440, n11441, n11442, n11443, n11444,
    n11445, n11446, n11447, n11448, n11449, n11450,
    n11451, n11452, n11453, n11454, n11455, n11456,
    n11457, n11458, n11459, n11460, n11461, n11462,
    n11463, n11464, n11465, n11466, n11467, n11468,
    n11469, n11470, n11471, n11472, n11473, n11474,
    n11475, n11476, n11477, n11478, n11479, n11480,
    n11481, n11482, n11483, n11484, n11485, n11486,
    n11487, n11488, n11489, n11490, n11491, n11492,
    n11493, n11494, n11495, n11496, n11497, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504,
    n11505, n11506, n11507, n11508, n11509, n11510,
    n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11520, n11521, n11522, n11523,
    n11524, n11525, n11526, n11527, n11528, n11529,
    n11530, n11531, n11532, n11533, n11534, n11535,
    n11536, n11537, n11538, n11539, n11540, n11541,
    n11542, n11543, n11544, n11545, n11546, n11547,
    n11548, n11549, n11550, n11551, n11552, n11553,
    n11554, n11555, n11556, n11557, n11558, n11559,
    n11560, n11561, n11562, n11563, n11564, n11565,
    n11566, n11567, n11568, n11569, n11570, n11571,
    n11572, n11573, n11574, n11575, n11576, n11577,
    n11578, n11579, n11580, n11581, n11582, n11583,
    n11584, n11585, n11586, n11587, n11588, n11589,
    n11590, n11591, n11592, n11593, n11594, n11595,
    n11596, n11597, n11598, n11599, n11600, n11601,
    n11602, n11603, n11604, n11605, n11606, n11607,
    n11608, n11609, n11610, n11611, n11612, n11613,
    n11614, n11615, n11616, n11617, n11618, n11619,
    n11620, n11621, n11622, n11623, n11624, n11625,
    n11626, n11627, n11628, n11629, n11630, n11631,
    n11632, n11633, n11634, n11635, n11636, n11637,
    n11638, n11639, n11640, n11641, n11642, n11643,
    n11644, n11645, n11646, n11647, n11648, n11649,
    n11650, n11651, n11652, n11653, n11654, n11655,
    n11656, n11657, n11658, n11659, n11660, n11661,
    n11662, n11663, n11664, n11665, n11666, n11667,
    n11668, n11669, n11670, n11671, n11672, n11673,
    n11674, n11675, n11676, n11677, n11678, n11679,
    n11680, n11681, n11682, n11683, n11684, n11685,
    n11686, n11687, n11688, n11689, n11690, n11691,
    n11692, n11693, n11694, n11695, n11696, n11697,
    n11698, n11699, n11700, n11701, n11702, n11703,
    n11704, n11705, n11706, n11707, n11708, n11709,
    n11710, n11711, n11712, n11713, n11714, n11715,
    n11716, n11717, n11718, n11719, n11720, n11721,
    n11722, n11723, n11724, n11725, n11726, n11727,
    n11728, n11729, n11730, n11731, n11732, n11733,
    n11734, n11735, n11736, n11737, n11738, n11739,
    n11740, n11741, n11742, n11743, n11744, n11745,
    n11746, n11747, n11748, n11749, n11750, n11751,
    n11752, n11753, n11754, n11755, n11756, n11757,
    n11758, n11759, n11760, n11761, n11762, n11763,
    n11764, n11765, n11766, n11767, n11768, n11769,
    n11770, n11771, n11772, n11773, n11774, n11775,
    n11776, n11777, n11778, n11779, n11780, n11781,
    n11782, n11783, n11784, n11785, n11786, n11787,
    n11788, n11789, n11790, n11791, n11792, n11793,
    n11794, n11795, n11796, n11797, n11798, n11799,
    n11800, n11801, n11802, n11803, n11804, n11805,
    n11806, n11807, n11808, n11809, n11810, n11811,
    n11812, n11813, n11814, n11815, n11816, n11817,
    n11818, n11819, n11820, n11821, n11822, n11823,
    n11824, n11825, n11826, n11827, n11828, n11829,
    n11830, n11831, n11832, n11833, n11834, n11835,
    n11836, n11837, n11838, n11839, n11840, n11841,
    n11842, n11843, n11844, n11845, n11846, n11847,
    n11848, n11849, n11850, n11851, n11852, n11853,
    n11854, n11855, n11856, n11857, n11858, n11859,
    n11860, n11861, n11862, n11863, n11864, n11865,
    n11866, n11867, n11868, n11869, n11870, n11871,
    n11872, n11873, n11874, n11875, n11876, n11877,
    n11878, n11879, n11880, n11881, n11882, n11883,
    n11884, n11885, n11886, n11887, n11888, n11889,
    n11890, n11891, n11892, n11893, n11894, n11895,
    n11896, n11897, n11898, n11899, n11900, n11901,
    n11902, n11903, n11904, n11905, n11906, n11907,
    n11908, n11909, n11910, n11911, n11912, n11913,
    n11914, n11915, n11916, n11917, n11918, n11919,
    n11920, n11921, n11922, n11923, n11924, n11925,
    n11926, n11927, n11928, n11929, n11930, n11931,
    n11932, n11933, n11934, n11935, n11936, n11937,
    n11938, n11939, n11940, n11941, n11942, n11943,
    n11944, n11945, n11946, n11947, n11948, n11949,
    n11950, n11951, n11952, n11953, n11954, n11955,
    n11956, n11957, n11958, n11959, n11960, n11961,
    n11962, n11963, n11964, n11965, n11966, n11967,
    n11968, n11969, n11970, n11971, n11972, n11973,
    n11974, n11975, n11976, n11977, n11978, n11979,
    n11980, n11981, n11982, n11983, n11984, n11985,
    n11986, n11987, n11988, n11989, n11990, n11991,
    n11992, n11993, n11994, n11995, n11996, n11997,
    n11998, n11999, n12000, n12001, n12002, n12003,
    n12004, n12005, n12006, n12007, n12008, n12009,
    n12010, n12011, n12012, n12013, n12014, n12015,
    n12016, n12017, n12018, n12019, n12020, n12021,
    n12022, n12023, n12024, n12025, n12026, n12027,
    n12028, n12029, n12030, n12031, n12032, n12033,
    n12034, n12035, n12036, n12037, n12038, n12039,
    n12040, n12041, n12042, n12043, n12044, n12045,
    n12046, n12047, n12048, n12049, n12050, n12051,
    n12052, n12053, n12054, n12055, n12056, n12057,
    n12058, n12059, n12060, n12061, n12062, n12063,
    n12064, n12065, n12066, n12067, n12068, n12069,
    n12070, n12071, n12073, n12074, n12075, n12076,
    n12077, n12078, n12079, n12080, n12081, n12082,
    n12083, n12084, n12085, n12086, n12087, n12088,
    n12089, n12090, n12091, n12092, n12093, n12094,
    n12095, n12096, n12097, n12098, n12099, n12100,
    n12101, n12102, n12103, n12104, n12105, n12106,
    n12107, n12108, n12109, n12110, n12111, n12112,
    n12113, n12114, n12115, n12116, n12117, n12118,
    n12119, n12120, n12121, n12122, n12123, n12124,
    n12125, n12126, n12127, n12128, n12129, n12130,
    n12131, n12132, n12133, n12134, n12135, n12136,
    n12137, n12138, n12139, n12140, n12141, n12142,
    n12143, n12144, n12145, n12146, n12147, n12148,
    n12149, n12150, n12151, n12152, n12153, n12154,
    n12155, n12156, n12157, n12158, n12159, n12160,
    n12161, n12162, n12163, n12164, n12165, n12166,
    n12167, n12168, n12169, n12170, n12171, n12172,
    n12173, n12174, n12175, n12176, n12177, n12178,
    n12179, n12180, n12181, n12182, n12183, n12184,
    n12185, n12186, n12187, n12188, n12189, n12190,
    n12191, n12192, n12193, n12194, n12195, n12196,
    n12197, n12198, n12199, n12200, n12201, n12202,
    n12203, n12204, n12205, n12206, n12207, n12208,
    n12209, n12210, n12211, n12212, n12213, n12214,
    n12215, n12216, n12217, n12218, n12219, n12220,
    n12221, n12222, n12223, n12224, n12225, n12226,
    n12227, n12228, n12229, n12230, n12231, n12232,
    n12233, n12234, n12235, n12236, n12237, n12238,
    n12239, n12240, n12241, n12242, n12243, n12244,
    n12245, n12246, n12247, n12248, n12249, n12250,
    n12251, n12252, n12253, n12254, n12255, n12256,
    n12257, n12258, n12259, n12260, n12261, n12262,
    n12263, n12264, n12265, n12266, n12267, n12268,
    n12269, n12270, n12271, n12272, n12273, n12274,
    n12275, n12276, n12277, n12278, n12279, n12280,
    n12281, n12282, n12283, n12284, n12285, n12286,
    n12287, n12288, n12289, n12290, n12291, n12292,
    n12293, n12294, n12295, n12296, n12297, n12298,
    n12299, n12300, n12301, n12302, n12303, n12304,
    n12305, n12306, n12307, n12308, n12309, n12310,
    n12311, n12312, n12313, n12314, n12315, n12316,
    n12317, n12318, n12319, n12320, n12321, n12322,
    n12323, n12324, n12325, n12326, n12327, n12328,
    n12329, n12330, n12331, n12332, n12333, n12334,
    n12335, n12336, n12337, n12338, n12339, n12340,
    n12341, n12342, n12343, n12344, n12345, n12346,
    n12347, n12348, n12349, n12350, n12351, n12352,
    n12353, n12354, n12355, n12356, n12357, n12358,
    n12359, n12360, n12361, n12362, n12363, n12364,
    n12365, n12366, n12367, n12368, n12369, n12370,
    n12371, n12372, n12373, n12374, n12375, n12376,
    n12377, n12378, n12379, n12380, n12381, n12382,
    n12383, n12384, n12385, n12386, n12387, n12388,
    n12389, n12390, n12391, n12392, n12393, n12394,
    n12395, n12396, n12397, n12398, n12399, n12400,
    n12401, n12402, n12403, n12404, n12405, n12406,
    n12407, n12408, n12409, n12410, n12411, n12412,
    n12413, n12414, n12415, n12416, n12417, n12418,
    n12419, n12420, n12421, n12422, n12423, n12424,
    n12425, n12426, n12427, n12428, n12429, n12430,
    n12431, n12432, n12433, n12434, n12435, n12436,
    n12437, n12438, n12439, n12440, n12441, n12442,
    n12443, n12444, n12445, n12446, n12447, n12448,
    n12449, n12450, n12451, n12452, n12453, n12454,
    n12455, n12456, n12457, n12458, n12459, n12460,
    n12461, n12462, n12463, n12464, n12465, n12466,
    n12467, n12468, n12469, n12470, n12471, n12472,
    n12473, n12474, n12475, n12476, n12477, n12478,
    n12479, n12480, n12481, n12482, n12483, n12484,
    n12485, n12486, n12487, n12488, n12489, n12490,
    n12491, n12492, n12493, n12494, n12495, n12496,
    n12497, n12498, n12499, n12500, n12501, n12502,
    n12503, n12504, n12505, n12506, n12507, n12508,
    n12509, n12510, n12511, n12512, n12513, n12514,
    n12515, n12516, n12517, n12518, n12519, n12520,
    n12521, n12522, n12523, n12524, n12525, n12526,
    n12527, n12528, n12529, n12530, n12531, n12532,
    n12533, n12534, n12535, n12536, n12537, n12538,
    n12539, n12540, n12541, n12542, n12543, n12544,
    n12545, n12546, n12547, n12548, n12549, n12550,
    n12551, n12552, n12553, n12554, n12555, n12556,
    n12557, n12558, n12559, n12560, n12561, n12562,
    n12563, n12564, n12565, n12566, n12567, n12568,
    n12569, n12570, n12571, n12572, n12573, n12574,
    n12575, n12576, n12577, n12578, n12579, n12580,
    n12581, n12582, n12583, n12584, n12585, n12586,
    n12587, n12588, n12589, n12590, n12591, n12592,
    n12593, n12594, n12595, n12596, n12597, n12598,
    n12599, n12600, n12601, n12602, n12603, n12604,
    n12605, n12606, n12607, n12608, n12609, n12610,
    n12611, n12612, n12613, n12614, n12615, n12616,
    n12617, n12618, n12619, n12620, n12621, n12622,
    n12623, n12624, n12625, n12626, n12628, n12629,
    n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641,
    n12642, n12643, n12644, n12645, n12646, n12647,
    n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659,
    n12660, n12661, n12662, n12663, n12664, n12665,
    n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677,
    n12678, n12679, n12680, n12681, n12682, n12683,
    n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12691, n12692, n12693, n12694, n12695,
    n12696, n12697, n12698, n12699, n12700, n12701,
    n12702, n12703, n12704, n12705, n12706, n12707,
    n12708, n12709, n12710, n12711, n12712, n12713,
    n12714, n12715, n12716, n12717, n12718, n12719,
    n12720, n12721, n12722, n12723, n12724, n12725,
    n12726, n12727, n12728, n12729, n12730, n12731,
    n12732, n12733, n12734, n12735, n12736, n12737,
    n12738, n12739, n12740, n12741, n12742, n12743,
    n12744, n12745, n12746, n12747, n12748, n12749,
    n12750, n12751, n12752, n12753, n12754, n12755,
    n12756, n12757, n12758, n12759, n12760, n12761,
    n12762, n12763, n12764, n12765, n12766, n12767,
    n12768, n12769, n12770, n12771, n12772, n12773,
    n12774, n12775, n12776, n12777, n12778, n12779,
    n12780, n12781, n12782, n12783, n12784, n12785,
    n12786, n12787, n12788, n12789, n12790, n12791,
    n12792, n12793, n12794, n12795, n12796, n12797,
    n12798, n12799, n12800, n12801, n12802, n12803,
    n12804, n12805, n12806, n12807, n12808, n12809,
    n12810, n12811, n12812, n12813, n12814, n12815,
    n12816, n12817, n12818, n12819, n12820, n12821,
    n12822, n12823, n12824, n12825, n12826, n12827,
    n12828, n12829, n12830, n12831, n12832, n12833,
    n12834, n12835, n12836, n12837, n12838, n12839,
    n12840, n12841, n12842, n12843, n12844, n12845,
    n12846, n12847, n12848, n12849, n12850, n12851,
    n12852, n12853, n12854, n12855, n12856, n12857,
    n12858, n12859, n12860, n12861, n12862, n12863,
    n12864, n12865, n12866, n12867, n12868, n12869,
    n12870, n12871, n12872, n12873, n12874, n12875,
    n12876, n12877, n12878, n12879, n12880, n12881,
    n12882, n12883, n12884, n12885, n12886, n12887,
    n12888, n12889, n12890, n12891, n12892, n12893,
    n12894, n12895, n12896, n12897, n12898, n12899,
    n12900, n12901, n12902, n12903, n12904, n12905,
    n12906, n12907, n12908, n12909, n12910, n12911,
    n12912, n12913, n12914, n12915, n12916, n12917,
    n12918, n12919, n12920, n12921, n12922, n12923,
    n12924, n12925, n12926, n12927, n12928, n12929,
    n12930, n12931, n12932, n12933, n12934, n12935,
    n12936, n12937, n12938, n12939, n12940, n12941,
    n12942, n12943, n12944, n12945, n12946, n12947,
    n12948, n12949, n12950, n12951, n12952, n12953,
    n12954, n12955, n12956, n12957, n12958, n12959,
    n12960, n12961, n12962, n12963, n12964, n12965,
    n12966, n12967, n12968, n12969, n12970, n12971,
    n12972, n12973, n12974, n12975, n12976, n12977,
    n12978, n12979, n12980, n12981, n12982, n12983,
    n12984, n12985, n12986, n12987, n12988, n12989,
    n12990, n12991, n12992, n12993, n12994, n12995,
    n12996, n12997, n12998, n12999, n13000, n13001,
    n13002, n13003, n13004, n13005, n13006, n13007,
    n13008, n13009, n13010, n13011, n13012, n13013,
    n13014, n13015, n13016, n13017, n13018, n13019,
    n13020, n13021, n13022, n13023, n13024, n13025,
    n13026, n13027, n13028, n13029, n13030, n13031,
    n13032, n13033, n13034, n13035, n13036, n13037,
    n13038, n13039, n13040, n13041, n13042, n13043,
    n13044, n13045, n13046, n13047, n13048, n13049,
    n13050, n13051, n13052, n13053, n13054, n13055,
    n13056, n13057, n13058, n13059, n13060, n13061,
    n13062, n13063, n13064, n13065, n13066, n13067,
    n13068, n13069, n13070, n13071, n13072, n13073,
    n13074, n13075, n13076, n13077, n13078, n13079,
    n13080, n13081, n13082, n13083, n13084, n13085,
    n13086, n13087, n13088, n13089, n13090, n13091,
    n13092, n13093, n13094, n13095, n13096, n13097,
    n13098, n13099, n13100, n13101, n13102, n13103,
    n13104, n13105, n13106, n13107, n13108, n13109,
    n13110, n13111, n13112, n13113, n13114, n13115,
    n13116, n13117, n13118, n13119, n13120, n13121,
    n13122, n13123, n13124, n13125, n13126, n13127,
    n13128, n13129, n13130, n13131, n13132, n13133,
    n13134, n13135, n13136, n13137, n13138, n13139,
    n13140, n13141, n13142, n13143, n13144, n13145,
    n13146, n13147, n13148, n13149, n13150, n13151,
    n13152, n13153, n13154, n13155, n13156, n13157,
    n13158, n13159, n13160, n13161, n13162, n13163,
    n13164, n13165, n13166, n13167, n13168, n13169,
    n13170, n13171, n13172, n13173, n13174, n13175,
    n13176, n13177, n13179, n13180, n13181, n13182,
    n13183, n13184, n13185, n13186, n13187, n13188,
    n13189, n13190, n13191, n13192, n13193, n13194,
    n13195, n13196, n13197, n13198, n13199, n13200,
    n13201, n13202, n13203, n13204, n13205, n13206,
    n13207, n13208, n13209, n13210, n13211, n13212,
    n13213, n13214, n13215, n13216, n13217, n13218,
    n13219, n13220, n13221, n13222, n13223, n13224,
    n13225, n13226, n13227, n13228, n13229, n13230,
    n13231, n13232, n13233, n13234, n13235, n13236,
    n13237, n13238, n13239, n13240, n13241, n13242,
    n13243, n13244, n13245, n13246, n13247, n13248,
    n13249, n13250, n13251, n13252, n13253, n13254,
    n13255, n13256, n13257, n13258, n13259, n13260,
    n13261, n13262, n13263, n13264, n13265, n13266,
    n13267, n13268, n13269, n13270, n13271, n13272,
    n13273, n13274, n13275, n13276, n13277, n13278,
    n13279, n13280, n13281, n13282, n13283, n13284,
    n13285, n13286, n13287, n13288, n13289, n13290,
    n13291, n13292, n13293, n13294, n13295, n13296,
    n13297, n13298, n13299, n13300, n13301, n13302,
    n13303, n13304, n13305, n13306, n13307, n13308,
    n13309, n13310, n13311, n13312, n13313, n13314,
    n13315, n13316, n13317, n13318, n13319, n13320,
    n13321, n13322, n13323, n13324, n13325, n13326,
    n13327, n13328, n13329, n13330, n13331, n13332,
    n13333, n13334, n13335, n13336, n13337, n13338,
    n13339, n13340, n13341, n13342, n13343, n13344,
    n13345, n13346, n13347, n13348, n13349, n13350,
    n13351, n13352, n13353, n13354, n13355, n13356,
    n13357, n13358, n13359, n13360, n13361, n13362,
    n13363, n13364, n13365, n13366, n13367, n13368,
    n13369, n13370, n13371, n13372, n13373, n13374,
    n13375, n13376, n13377, n13378, n13379, n13380,
    n13381, n13382, n13383, n13384, n13385, n13386,
    n13387, n13388, n13389, n13390, n13391, n13392,
    n13393, n13394, n13395, n13396, n13397, n13398,
    n13399, n13400, n13401, n13402, n13403, n13404,
    n13405, n13406, n13407, n13408, n13409, n13410,
    n13411, n13412, n13413, n13414, n13415, n13416,
    n13417, n13418, n13419, n13420, n13421, n13422,
    n13423, n13424, n13425, n13426, n13427, n13428,
    n13429, n13430, n13431, n13432, n13433, n13434,
    n13435, n13436, n13437, n13438, n13439, n13440,
    n13441, n13442, n13443, n13444, n13445, n13446,
    n13447, n13448, n13449, n13450, n13451, n13452,
    n13453, n13454, n13455, n13456, n13457, n13458,
    n13459, n13460, n13461, n13462, n13463, n13464,
    n13465, n13466, n13467, n13468, n13469, n13470,
    n13471, n13472, n13473, n13474, n13475, n13476,
    n13477, n13478, n13479, n13480, n13481, n13482,
    n13483, n13484, n13485, n13486, n13487, n13488,
    n13489, n13490, n13491, n13492, n13493, n13494,
    n13495, n13496, n13497, n13498, n13499, n13500,
    n13501, n13502, n13503, n13504, n13505, n13506,
    n13507, n13508, n13509, n13510, n13511, n13512,
    n13513, n13514, n13515, n13516, n13517, n13518,
    n13519, n13520, n13521, n13522, n13523, n13524,
    n13525, n13526, n13527, n13528, n13529, n13530,
    n13531, n13532, n13533, n13534, n13535, n13536,
    n13537, n13538, n13539, n13540, n13541, n13542,
    n13543, n13544, n13545, n13546, n13547, n13548,
    n13549, n13550, n13551, n13552, n13553, n13554,
    n13555, n13556, n13557, n13558, n13559, n13560,
    n13561, n13562, n13563, n13564, n13565, n13566,
    n13567, n13568, n13569, n13570, n13571, n13572,
    n13573, n13574, n13575, n13576, n13577, n13578,
    n13579, n13580, n13581, n13582, n13583, n13584,
    n13585, n13586, n13587, n13588, n13589, n13590,
    n13591, n13592, n13593, n13594, n13595, n13596,
    n13597, n13598, n13599, n13600, n13601, n13602,
    n13603, n13604, n13605, n13606, n13607, n13608,
    n13609, n13610, n13611, n13612, n13613, n13614,
    n13615, n13616, n13617, n13618, n13619, n13620,
    n13621, n13622, n13623, n13624, n13625, n13626,
    n13627, n13628, n13629, n13630, n13631, n13632,
    n13633, n13634, n13635, n13636, n13637, n13638,
    n13639, n13640, n13641, n13642, n13643, n13644,
    n13645, n13646, n13647, n13648, n13649, n13650,
    n13651, n13652, n13653, n13654, n13655, n13656,
    n13657, n13658, n13659, n13660, n13661, n13662,
    n13663, n13664, n13665, n13666, n13667, n13668,
    n13669, n13670, n13671, n13672, n13673, n13674,
    n13675, n13676, n13677, n13678, n13679, n13680,
    n13681, n13682, n13683, n13684, n13685, n13686,
    n13687, n13688, n13689, n13690, n13691, n13692,
    n13693, n13694, n13695, n13696, n13697, n13698,
    n13699, n13700, n13702, n13703, n13704, n13705,
    n13706, n13707, n13708, n13709, n13710, n13711,
    n13712, n13713, n13714, n13715, n13716, n13717,
    n13718, n13719, n13720, n13721, n13722, n13723,
    n13724, n13725, n13726, n13727, n13728, n13729,
    n13730, n13731, n13732, n13733, n13734, n13735,
    n13736, n13737, n13738, n13739, n13740, n13741,
    n13742, n13743, n13744, n13745, n13746, n13747,
    n13748, n13749, n13750, n13751, n13752, n13753,
    n13754, n13755, n13756, n13757, n13758, n13759,
    n13760, n13761, n13762, n13763, n13764, n13765,
    n13766, n13767, n13768, n13769, n13770, n13771,
    n13772, n13773, n13774, n13775, n13776, n13777,
    n13778, n13779, n13780, n13781, n13782, n13783,
    n13784, n13785, n13786, n13787, n13788, n13789,
    n13790, n13791, n13792, n13793, n13794, n13795,
    n13796, n13797, n13798, n13799, n13800, n13801,
    n13802, n13803, n13804, n13805, n13806, n13807,
    n13808, n13809, n13810, n13811, n13812, n13813,
    n13814, n13815, n13816, n13817, n13818, n13819,
    n13820, n13821, n13822, n13823, n13824, n13825,
    n13826, n13827, n13828, n13829, n13830, n13831,
    n13832, n13833, n13834, n13835, n13836, n13837,
    n13838, n13839, n13840, n13841, n13842, n13843,
    n13844, n13845, n13846, n13847, n13848, n13849,
    n13850, n13851, n13852, n13853, n13854, n13855,
    n13856, n13857, n13858, n13859, n13860, n13861,
    n13862, n13863, n13864, n13865, n13866, n13867,
    n13868, n13869, n13870, n13871, n13872, n13873,
    n13874, n13875, n13876, n13877, n13878, n13879,
    n13880, n13881, n13882, n13883, n13884, n13885,
    n13886, n13887, n13888, n13889, n13890, n13891,
    n13892, n13893, n13894, n13895, n13896, n13897,
    n13898, n13899, n13900, n13901, n13902, n13903,
    n13904, n13905, n13906, n13907, n13908, n13909,
    n13910, n13911, n13912, n13913, n13914, n13915,
    n13916, n13917, n13918, n13919, n13920, n13921,
    n13922, n13923, n13924, n13925, n13926, n13927,
    n13928, n13929, n13930, n13931, n13932, n13933,
    n13934, n13935, n13936, n13937, n13938, n13939,
    n13940, n13941, n13942, n13943, n13944, n13945,
    n13946, n13947, n13948, n13949, n13950, n13951,
    n13952, n13953, n13954, n13955, n13956, n13957,
    n13958, n13959, n13960, n13961, n13962, n13963,
    n13964, n13965, n13966, n13967, n13968, n13969,
    n13970, n13971, n13972, n13973, n13974, n13975,
    n13976, n13977, n13978, n13979, n13980, n13981,
    n13982, n13983, n13984, n13985, n13986, n13987,
    n13988, n13989, n13990, n13991, n13992, n13993,
    n13994, n13995, n13996, n13997, n13998, n13999,
    n14000, n14001, n14002, n14003, n14004, n14005,
    n14006, n14007, n14008, n14009, n14010, n14011,
    n14012, n14013, n14014, n14015, n14016, n14017,
    n14018, n14019, n14020, n14021, n14022, n14023,
    n14024, n14025, n14026, n14027, n14028, n14029,
    n14030, n14031, n14032, n14033, n14034, n14035,
    n14036, n14037, n14038, n14039, n14040, n14041,
    n14042, n14043, n14044, n14045, n14046, n14047,
    n14048, n14049, n14050, n14051, n14052, n14053,
    n14054, n14055, n14056, n14057, n14058, n14059,
    n14060, n14061, n14062, n14063, n14064, n14065,
    n14066, n14067, n14068, n14069, n14070, n14071,
    n14072, n14073, n14074, n14075, n14076, n14077,
    n14078, n14079, n14080, n14081, n14082, n14083,
    n14084, n14085, n14086, n14087, n14088, n14089,
    n14090, n14091, n14092, n14093, n14094, n14095,
    n14096, n14097, n14098, n14099, n14100, n14101,
    n14102, n14103, n14104, n14105, n14106, n14107,
    n14108, n14109, n14110, n14111, n14112, n14113,
    n14114, n14115, n14116, n14117, n14118, n14119,
    n14120, n14121, n14122, n14123, n14124, n14125,
    n14126, n14127, n14128, n14129, n14130, n14131,
    n14132, n14133, n14134, n14135, n14136, n14137,
    n14138, n14139, n14140, n14141, n14142, n14143,
    n14144, n14145, n14146, n14147, n14148, n14149,
    n14150, n14151, n14152, n14153, n14154, n14155,
    n14156, n14157, n14158, n14159, n14160, n14161,
    n14162, n14163, n14164, n14165, n14166, n14167,
    n14168, n14169, n14170, n14171, n14172, n14173,
    n14174, n14175, n14176, n14177, n14178, n14179,
    n14180, n14181, n14182, n14183, n14184, n14185,
    n14186, n14187, n14188, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197,
    n14198, n14199, n14200, n14201, n14202, n14203,
    n14204, n14205, n14206, n14207, n14208, n14209,
    n14210, n14211, n14212, n14213, n14214, n14215,
    n14216, n14217, n14218, n14219, n14220, n14221,
    n14222, n14223, n14224, n14225, n14226, n14227,
    n14228, n14229, n14230, n14231, n14232, n14233,
    n14234, n14235, n14236, n14237, n14238, n14239,
    n14240, n14241, n14242, n14243, n14244, n14245,
    n14246, n14247, n14248, n14249, n14250, n14251,
    n14252, n14253, n14254, n14255, n14256, n14257,
    n14258, n14259, n14260, n14261, n14262, n14263,
    n14264, n14265, n14266, n14267, n14268, n14269,
    n14270, n14271, n14272, n14273, n14274, n14275,
    n14276, n14277, n14278, n14279, n14280, n14281,
    n14282, n14283, n14284, n14285, n14286, n14287,
    n14288, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14329, n14330,
    n14331, n14332, n14333, n14334, n14335, n14336,
    n14337, n14338, n14339, n14340, n14341, n14342,
    n14343, n14344, n14345, n14346, n14347, n14348,
    n14349, n14350, n14351, n14352, n14353, n14354,
    n14355, n14356, n14357, n14358, n14359, n14360,
    n14361, n14362, n14363, n14364, n14365, n14366,
    n14367, n14368, n14369, n14370, n14371, n14372,
    n14373, n14374, n14375, n14376, n14377, n14378,
    n14379, n14380, n14381, n14382, n14383, n14384,
    n14385, n14386, n14387, n14388, n14389, n14390,
    n14391, n14392, n14393, n14394, n14395, n14396,
    n14397, n14398, n14399, n14400, n14401, n14402,
    n14403, n14404, n14405, n14406, n14407, n14408,
    n14409, n14410, n14411, n14412, n14413, n14414,
    n14415, n14416, n14417, n14418, n14419, n14420,
    n14421, n14422, n14423, n14424, n14425, n14426,
    n14427, n14428, n14429, n14430, n14431, n14432,
    n14433, n14434, n14435, n14436, n14437, n14438,
    n14439, n14440, n14441, n14442, n14443, n14444,
    n14445, n14446, n14447, n14448, n14449, n14450,
    n14451, n14452, n14453, n14454, n14455, n14456,
    n14457, n14458, n14459, n14460, n14461, n14462,
    n14463, n14464, n14465, n14466, n14467, n14468,
    n14469, n14470, n14471, n14472, n14473, n14474,
    n14475, n14476, n14477, n14478, n14479, n14480,
    n14481, n14482, n14483, n14484, n14485, n14486,
    n14487, n14488, n14489, n14490, n14491, n14492,
    n14493, n14494, n14495, n14496, n14497, n14498,
    n14499, n14500, n14501, n14502, n14503, n14504,
    n14505, n14506, n14507, n14508, n14509, n14510,
    n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522,
    n14523, n14524, n14525, n14526, n14527, n14528,
    n14529, n14530, n14531, n14532, n14533, n14534,
    n14535, n14536, n14537, n14538, n14539, n14540,
    n14541, n14542, n14543, n14544, n14545, n14546,
    n14547, n14548, n14549, n14550, n14551, n14552,
    n14553, n14554, n14555, n14556, n14557, n14558,
    n14559, n14560, n14561, n14562, n14563, n14564,
    n14565, n14566, n14567, n14568, n14569, n14570,
    n14571, n14572, n14573, n14574, n14575, n14576,
    n14577, n14578, n14579, n14580, n14581, n14582,
    n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594,
    n14595, n14596, n14597, n14598, n14599, n14600,
    n14601, n14602, n14603, n14604, n14605, n14606,
    n14607, n14608, n14609, n14610, n14611, n14612,
    n14613, n14614, n14615, n14616, n14617, n14618,
    n14619, n14620, n14621, n14622, n14623, n14624,
    n14625, n14626, n14627, n14628, n14629, n14630,
    n14631, n14632, n14633, n14634, n14635, n14636,
    n14637, n14638, n14639, n14640, n14641, n14642,
    n14643, n14644, n14645, n14646, n14647, n14648,
    n14649, n14650, n14651, n14652, n14653, n14654,
    n14655, n14656, n14657, n14658, n14659, n14660,
    n14661, n14662, n14663, n14664, n14665, n14666,
    n14667, n14668, n14669, n14670, n14671, n14672,
    n14673, n14674, n14675, n14676, n14677, n14678,
    n14679, n14680, n14681, n14682, n14683, n14684,
    n14685, n14686, n14687, n14688, n14689, n14690,
    n14691, n14692, n14693, n14694, n14695, n14696,
    n14697, n14698, n14699, n14700, n14701, n14702,
    n14703, n14704, n14705, n14706, n14707, n14708,
    n14709, n14710, n14711, n14712, n14713, n14714,
    n14715, n14716, n14717, n14718, n14719, n14720,
    n14721, n14722, n14723, n14724, n14725, n14726,
    n14727, n14728, n14729, n14730, n14731, n14732,
    n14733, n14734, n14735, n14736, n14737, n14738,
    n14739, n14740, n14741, n14742, n14743, n14744,
    n14745, n14746, n14747, n14748, n14749, n14750,
    n14751, n14752, n14753, n14754, n14755, n14756,
    n14757, n14758, n14759, n14760, n14761, n14762,
    n14763, n14764, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780,
    n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816,
    n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828,
    n14830, n14831, n14832, n14833, n14834, n14835,
    n14836, n14837, n14838, n14839, n14840, n14841,
    n14842, n14843, n14844, n14845, n14846, n14847,
    n14848, n14849, n14850, n14851, n14852, n14853,
    n14854, n14855, n14856, n14857, n14858, n14859,
    n14860, n14861, n14862, n14863, n14864, n14865,
    n14866, n14867, n14868, n14869, n14870, n14871,
    n14872, n14873, n14874, n14875, n14876, n14877,
    n14878, n14879, n14880, n14881, n14882, n14883,
    n14884, n14885, n14886, n14887, n14888, n14889,
    n14890, n14891, n14892, n14893, n14894, n14895,
    n14896, n14897, n14898, n14899, n14900, n14901,
    n14902, n14903, n14904, n14905, n14906, n14907,
    n14908, n14909, n14910, n14911, n14912, n14913,
    n14914, n14915, n14916, n14917, n14918, n14919,
    n14920, n14921, n14922, n14923, n14924, n14925,
    n14926, n14927, n14928, n14929, n14930, n14931,
    n14932, n14933, n14934, n14935, n14936, n14937,
    n14938, n14939, n14940, n14941, n14942, n14943,
    n14944, n14945, n14946, n14947, n14948, n14949,
    n14950, n14951, n14952, n14953, n14954, n14955,
    n14956, n14957, n14958, n14959, n14960, n14961,
    n14962, n14963, n14964, n14965, n14966, n14967,
    n14968, n14969, n14970, n14971, n14972, n14973,
    n14974, n14975, n14976, n14977, n14978, n14979,
    n14980, n14981, n14982, n14983, n14984, n14985,
    n14986, n14987, n14988, n14989, n14990, n14991,
    n14992, n14993, n14994, n14995, n14996, n14997,
    n14998, n14999, n15000, n15001, n15002, n15003,
    n15004, n15005, n15006, n15007, n15008, n15009,
    n15010, n15011, n15012, n15013, n15014, n15015,
    n15016, n15017, n15018, n15019, n15020, n15021,
    n15022, n15023, n15024, n15025, n15026, n15027,
    n15028, n15029, n15030, n15031, n15032, n15033,
    n15034, n15035, n15036, n15037, n15038, n15039,
    n15040, n15041, n15042, n15043, n15044, n15045,
    n15046, n15047, n15048, n15049, n15050, n15051,
    n15052, n15053, n15054, n15055, n15056, n15057,
    n15058, n15059, n15060, n15061, n15062, n15063,
    n15064, n15065, n15066, n15067, n15068, n15069,
    n15070, n15071, n15072, n15073, n15074, n15075,
    n15076, n15077, n15078, n15079, n15080, n15081,
    n15082, n15083, n15084, n15085, n15086, n15087,
    n15088, n15089, n15090, n15091, n15092, n15093,
    n15094, n15095, n15096, n15097, n15098, n15099,
    n15100, n15101, n15102, n15103, n15104, n15105,
    n15106, n15107, n15108, n15109, n15110, n15111,
    n15112, n15113, n15114, n15115, n15116, n15117,
    n15118, n15119, n15120, n15121, n15122, n15123,
    n15124, n15125, n15126, n15127, n15128, n15129,
    n15130, n15131, n15132, n15133, n15134, n15135,
    n15136, n15137, n15138, n15139, n15140, n15141,
    n15142, n15143, n15144, n15145, n15146, n15147,
    n15148, n15149, n15150, n15151, n15152, n15153,
    n15154, n15155, n15156, n15157, n15158, n15159,
    n15160, n15161, n15162, n15163, n15164, n15165,
    n15166, n15167, n15168, n15169, n15170, n15171,
    n15172, n15173, n15174, n15175, n15176, n15177,
    n15178, n15179, n15180, n15181, n15182, n15183,
    n15184, n15185, n15186, n15187, n15188, n15189,
    n15190, n15191, n15192, n15193, n15194, n15195,
    n15196, n15197, n15198, n15199, n15200, n15201,
    n15202, n15203, n15204, n15205, n15206, n15207,
    n15208, n15209, n15210, n15211, n15212, n15213,
    n15214, n15215, n15216, n15217, n15218, n15219,
    n15220, n15221, n15222, n15223, n15224, n15225,
    n15226, n15227, n15228, n15229, n15230, n15231,
    n15232, n15233, n15234, n15235, n15236, n15237,
    n15238, n15239, n15240, n15241, n15242, n15243,
    n15244, n15245, n15246, n15247, n15248, n15249,
    n15250, n15251, n15252, n15253, n15254, n15255,
    n15256, n15257, n15258, n15259, n15260, n15261,
    n15262, n15263, n15264, n15265, n15266, n15267,
    n15268, n15269, n15270, n15271, n15272, n15273,
    n15274, n15275, n15276, n15277, n15278, n15279,
    n15280, n15281, n15282, n15283, n15284, n15285,
    n15286, n15287, n15288, n15289, n15290, n15291,
    n15292, n15293, n15294, n15295, n15296, n15297,
    n15298, n15299, n15300, n15301, n15302, n15303,
    n15304, n15305, n15306, n15307, n15308, n15309,
    n15310, n15311, n15312, n15313, n15314, n15315,
    n15316, n15317, n15318, n15319, n15320, n15321,
    n15322, n15323, n15324, n15325, n15326, n15327,
    n15328, n15329, n15330, n15331, n15332, n15333,
    n15334, n15335, n15336, n15337, n15338, n15339,
    n15340, n15341, n15342, n15343, n15344, n15345,
    n15346, n15347, n15348, n15349, n15350, n15351,
    n15352, n15353, n15354, n15355, n15356, n15357,
    n15358, n15359, n15360, n15361, n15362, n15363,
    n15364, n15365, n15366, n15367, n15368, n15369,
    n15370, n15371, n15372, n15373, n15374, n15375,
    n15376, n15377, n15378, n15379, n15380, n15381,
    n15382, n15383, n15384, n15385, n15386, n15387,
    n15388, n15389, n15390, n15391, n15392, n15393,
    n15394, n15395, n15396, n15397, n15398, n15399,
    n15400, n15401, n15402, n15403, n15404, n15405,
    n15406, n15407, n15408, n15409, n15410, n15411,
    n15412, n15413, n15414, n15415, n15416, n15417,
    n15418, n15419, n15420, n15421, n15422, n15423,
    n15424, n15425, n15426, n15427, n15428, n15429,
    n15431, n15432, n15433, n15434, n15435, n15436,
    n15437, n15438, n15439, n15440, n15441, n15442,
    n15443, n15444, n15445, n15446, n15447, n15448,
    n15449, n15450, n15451, n15452, n15453, n15454,
    n15455, n15456, n15457, n15458, n15459, n15460,
    n15461, n15462, n15463, n15464, n15465, n15466,
    n15467, n15468, n15469, n15470, n15471, n15472,
    n15473, n15474, n15475, n15476, n15477, n15478,
    n15479, n15480, n15481, n15482, n15483, n15484,
    n15485, n15486, n15487, n15488, n15489, n15490,
    n15491, n15492, n15493, n15494, n15495, n15496,
    n15497, n15498, n15499, n15500, n15501, n15502,
    n15503, n15504, n15505, n15506, n15507, n15508,
    n15509, n15510, n15511, n15512, n15513, n15514,
    n15515, n15516, n15517, n15518, n15519, n15520,
    n15521, n15522, n15523, n15524, n15525, n15526,
    n15527, n15528, n15529, n15530, n15531, n15532,
    n15533, n15534, n15535, n15536, n15537, n15538,
    n15539, n15540, n15541, n15542, n15543, n15544,
    n15545, n15546, n15547, n15548, n15549, n15550,
    n15551, n15552, n15553, n15554, n15555, n15556,
    n15557, n15558, n15559, n15560, n15561, n15562,
    n15563, n15564, n15565, n15566, n15567, n15568,
    n15569, n15570, n15571, n15572, n15573, n15574,
    n15575, n15576, n15577, n15578, n15579, n15580,
    n15581, n15582, n15583, n15584, n15585, n15586,
    n15587, n15588, n15589, n15590, n15591, n15592,
    n15593, n15594, n15595, n15596, n15597, n15598,
    n15599, n15600, n15601, n15602, n15603, n15604,
    n15605, n15606, n15607, n15608, n15609, n15610,
    n15611, n15612, n15613, n15614, n15615, n15616,
    n15617, n15618, n15619, n15620, n15621, n15622,
    n15623, n15624, n15625, n15626, n15627, n15628,
    n15629, n15630, n15631, n15632, n15633, n15634,
    n15635, n15636, n15637, n15638, n15639, n15640,
    n15641, n15642, n15643, n15644, n15645, n15646,
    n15647, n15648, n15649, n15650, n15651, n15652,
    n15653, n15654, n15655, n15656, n15657, n15658,
    n15659, n15660, n15661, n15662, n15663, n15664,
    n15665, n15666, n15667, n15668, n15669, n15670,
    n15671, n15672, n15673, n15674, n15675, n15676,
    n15677, n15678, n15679, n15680, n15681, n15682,
    n15683, n15684, n15685, n15686, n15687, n15688,
    n15689, n15690, n15691, n15692, n15693, n15694,
    n15695, n15696, n15697, n15698, n15699, n15700,
    n15701, n15702, n15703, n15704, n15705, n15706,
    n15707, n15708, n15709, n15710, n15711, n15712,
    n15713, n15714, n15715, n15716, n15717, n15718,
    n15719, n15720, n15721, n15722, n15723, n15724,
    n15725, n15726, n15727, n15728, n15729, n15730,
    n15731, n15732, n15733, n15734, n15735, n15736,
    n15737, n15738, n15739, n15740, n15741, n15742,
    n15743, n15744, n15745, n15746, n15747, n15748,
    n15749, n15750, n15751, n15752, n15753, n15754,
    n15755, n15756, n15757, n15758, n15759, n15760,
    n15761, n15762, n15763, n15764, n15765, n15766,
    n15767, n15768, n15769, n15770, n15771, n15772,
    n15773, n15774, n15775, n15776, n15777, n15778,
    n15779, n15780, n15781, n15782, n15783, n15784,
    n15785, n15786, n15787, n15788, n15789, n15790,
    n15791, n15792, n15793, n15794, n15795, n15796,
    n15797, n15798, n15799, n15800, n15801, n15802,
    n15803, n15804, n15805, n15806, n15807, n15808,
    n15809, n15810, n15811, n15812, n15813, n15814,
    n15815, n15816, n15817, n15818, n15819, n15820,
    n15821, n15822, n15823, n15824, n15825, n15826,
    n15827, n15828, n15829, n15830, n15831, n15832,
    n15833, n15834, n15835, n15836, n15837, n15838,
    n15839, n15840, n15841, n15842, n15843, n15844,
    n15845, n15846, n15847, n15848, n15849, n15850,
    n15851, n15852, n15853, n15854, n15855, n15856,
    n15857, n15858, n15859, n15860, n15861, n15862,
    n15863, n15864, n15865, n15866, n15867, n15868,
    n15869, n15870, n15871, n15872, n15873, n15874,
    n15875, n15876, n15877, n15878, n15879, n15880,
    n15881, n15882, n15883, n15884, n15885, n15886,
    n15887, n15888, n15889, n15890, n15891, n15892,
    n15893, n15894, n15895, n15896, n15897, n15898,
    n15899, n15900, n15901, n15902, n15903, n15904,
    n15905, n15906, n15907, n15908, n15909, n15910,
    n15911, n15912, n15913, n15914, n15915, n15916,
    n15917, n15918, n15919, n15920, n15921, n15922,
    n15923, n15924, n15925, n15926, n15927, n15928,
    n15929, n15930, n15931, n15932, n15933, n15934,
    n15935, n15936, n15937, n15938, n15939, n15940,
    n15941, n15942, n15943, n15944, n15945, n15946,
    n15947, n15948, n15949, n15950, n15951, n15952,
    n15953, n15954, n15955, n15956, n15957, n15958,
    n15959, n15960, n15961, n15962, n15963, n15964,
    n15965, n15966, n15967, n15968, n15969, n15970,
    n15972, n15973, n15974, n15975, n15976, n15977,
    n15978, n15979, n15980, n15981, n15982, n15983,
    n15984, n15985, n15986, n15987, n15988, n15989,
    n15990, n15991, n15992, n15993, n15994, n15995,
    n15996, n15997, n15998, n15999, n16000, n16001,
    n16002, n16003, n16004, n16005, n16006, n16007,
    n16008, n16009, n16010, n16011, n16012, n16013,
    n16014, n16015, n16016, n16017, n16018, n16019,
    n16020, n16021, n16022, n16023, n16024, n16025,
    n16026, n16027, n16028, n16029, n16030, n16031,
    n16032, n16033, n16034, n16035, n16036, n16037,
    n16038, n16039, n16040, n16041, n16042, n16043,
    n16044, n16045, n16046, n16047, n16048, n16049,
    n16050, n16051, n16052, n16053, n16054, n16055,
    n16056, n16057, n16058, n16059, n16060, n16061,
    n16062, n16063, n16064, n16065, n16066, n16067,
    n16068, n16069, n16070, n16071, n16072, n16073,
    n16074, n16075, n16076, n16077, n16078, n16079,
    n16080, n16081, n16082, n16083, n16084, n16085,
    n16086, n16087, n16088, n16089, n16090, n16091,
    n16092, n16093, n16094, n16095, n16096, n16097,
    n16098, n16099, n16100, n16101, n16102, n16103,
    n16104, n16105, n16106, n16107, n16108, n16109,
    n16110, n16111, n16112, n16113, n16114, n16115,
    n16116, n16117, n16118, n16119, n16120, n16121,
    n16122, n16123, n16124, n16125, n16126, n16127,
    n16128, n16129, n16130, n16131, n16132, n16133,
    n16134, n16135, n16136, n16137, n16138, n16139,
    n16140, n16141, n16142, n16143, n16144, n16145,
    n16146, n16147, n16148, n16149, n16150, n16151,
    n16152, n16153, n16154, n16155, n16156, n16157,
    n16158, n16159, n16160, n16161, n16162, n16163,
    n16164, n16165, n16166, n16167, n16168, n16169,
    n16170, n16171, n16172, n16173, n16174, n16175,
    n16176, n16177, n16178, n16179, n16180, n16181,
    n16182, n16183, n16184, n16185, n16186, n16187,
    n16188, n16189, n16190, n16191, n16192, n16193,
    n16194, n16195, n16196, n16197, n16198, n16199,
    n16200, n16201, n16202, n16203, n16204, n16205,
    n16206, n16207, n16208, n16209, n16210, n16211,
    n16212, n16213, n16214, n16215, n16216, n16217,
    n16218, n16219, n16220, n16221, n16222, n16223,
    n16224, n16225, n16226, n16227, n16228, n16229,
    n16230, n16231, n16232, n16233, n16234, n16235,
    n16236, n16237, n16238, n16239, n16240, n16241,
    n16242, n16243, n16244, n16245, n16246, n16247,
    n16248, n16249, n16250, n16251, n16252, n16253,
    n16254, n16255, n16256, n16257, n16258, n16259,
    n16260, n16261, n16262, n16263, n16264, n16265,
    n16266, n16267, n16268, n16269, n16270, n16271,
    n16272, n16273, n16274, n16275, n16276, n16277,
    n16278, n16279, n16280, n16281, n16282, n16283,
    n16284, n16285, n16286, n16287, n16288, n16289,
    n16290, n16291, n16292, n16293, n16294, n16295,
    n16296, n16297, n16298, n16299, n16300, n16301,
    n16302, n16303, n16304, n16305, n16306, n16307,
    n16308, n16309, n16310, n16311, n16312, n16313,
    n16314, n16315, n16316, n16317, n16318, n16319,
    n16320, n16321, n16322, n16323, n16324, n16325,
    n16326, n16327, n16328, n16329, n16330, n16331,
    n16332, n16333, n16334, n16335, n16336, n16337,
    n16338, n16339, n16340, n16341, n16342, n16343,
    n16344, n16345, n16346, n16347, n16348, n16349,
    n16350, n16351, n16352, n16353, n16354, n16355,
    n16356, n16357, n16358, n16359, n16360, n16361,
    n16362, n16363, n16364, n16365, n16366, n16367,
    n16368, n16369, n16370, n16371, n16372, n16373,
    n16374, n16375, n16376, n16377, n16378, n16379,
    n16380, n16381, n16382, n16383, n16384, n16385,
    n16386, n16387, n16388, n16389, n16390, n16391,
    n16392, n16393, n16394, n16395, n16396, n16397,
    n16398, n16399, n16400, n16401, n16402, n16403,
    n16404, n16405, n16406, n16407, n16408, n16409,
    n16410, n16411, n16412, n16413, n16414, n16415,
    n16416, n16417, n16418, n16419, n16420, n16421,
    n16422, n16423, n16424, n16425, n16426, n16427,
    n16428, n16429, n16430, n16431, n16432, n16433,
    n16434, n16435, n16436, n16437, n16438, n16439,
    n16440, n16441, n16442, n16443, n16444, n16445,
    n16446, n16447, n16448, n16449, n16450, n16451,
    n16452, n16453, n16454, n16455, n16456, n16457,
    n16458, n16459, n16460, n16461, n16462, n16463,
    n16464, n16465, n16466, n16467, n16468, n16469,
    n16470, n16471, n16472, n16473, n16474, n16475,
    n16476, n16477, n16478, n16479, n16480, n16481,
    n16482, n16483, n16484, n16485, n16486, n16487,
    n16488, n16489, n16490, n16491, n16492, n16493,
    n16494, n16495, n16496, n16497, n16498, n16499,
    n16500, n16501, n16502, n16503, n16504, n16505,
    n16506, n16507, n16508, n16509, n16510, n16511,
    n16513, n16514, n16515, n16516, n16517, n16518,
    n16519, n16520, n16521, n16522, n16523, n16524,
    n16525, n16526, n16527, n16528, n16529, n16530,
    n16531, n16532, n16533, n16534, n16535, n16536,
    n16537, n16538, n16539, n16540, n16541, n16542,
    n16543, n16544, n16545, n16546, n16547, n16548,
    n16549, n16550, n16551, n16552, n16553, n16554,
    n16555, n16556, n16557, n16558, n16559, n16560,
    n16561, n16562, n16563, n16564, n16565, n16566,
    n16567, n16568, n16569, n16570, n16571, n16572,
    n16573, n16574, n16575, n16576, n16577, n16578,
    n16579, n16580, n16581, n16582, n16583, n16584,
    n16585, n16586, n16587, n16588, n16589, n16590,
    n16591, n16592, n16593, n16594, n16595, n16596,
    n16597, n16598, n16599, n16600, n16601, n16602,
    n16603, n16604, n16605, n16606, n16607, n16608,
    n16609, n16610, n16611, n16612, n16613, n16614,
    n16615, n16616, n16617, n16618, n16619, n16620,
    n16621, n16622, n16623, n16624, n16625, n16626,
    n16627, n16628, n16629, n16630, n16631, n16632,
    n16633, n16634, n16635, n16636, n16637, n16638,
    n16639, n16640, n16641, n16642, n16643, n16644,
    n16645, n16646, n16647, n16648, n16649, n16650,
    n16651, n16652, n16653, n16654, n16655, n16656,
    n16657, n16658, n16659, n16660, n16661, n16662,
    n16663, n16664, n16665, n16666, n16667, n16668,
    n16669, n16670, n16671, n16672, n16673, n16674,
    n16675, n16676, n16677, n16678, n16679, n16680,
    n16681, n16682, n16683, n16684, n16685, n16686,
    n16687, n16688, n16689, n16690, n16691, n16692,
    n16693, n16694, n16695, n16696, n16697, n16698,
    n16699, n16700, n16701, n16702, n16703, n16704,
    n16705, n16706, n16707, n16708, n16709, n16710,
    n16711, n16712, n16713, n16714, n16715, n16716,
    n16717, n16718, n16719, n16720, n16721, n16722,
    n16723, n16724, n16725, n16726, n16727, n16728,
    n16729, n16730, n16731, n16732, n16733, n16734,
    n16735, n16736, n16737, n16738, n16739, n16740,
    n16741, n16742, n16743, n16744, n16745, n16746,
    n16747, n16748, n16749, n16750, n16751, n16752,
    n16753, n16754, n16755, n16756, n16757, n16758,
    n16759, n16760, n16761, n16762, n16763, n16764,
    n16765, n16766, n16767, n16768, n16769, n16770,
    n16771, n16772, n16773, n16774, n16775, n16776,
    n16777, n16778, n16779, n16780, n16781, n16782,
    n16783, n16784, n16785, n16786, n16787, n16788,
    n16789, n16790, n16791, n16792, n16793, n16794,
    n16795, n16796, n16797, n16798, n16799, n16800,
    n16801, n16802, n16803, n16804, n16805, n16806,
    n16807, n16808, n16809, n16810, n16811, n16812,
    n16813, n16814, n16815, n16816, n16817, n16818,
    n16819, n16820, n16821, n16822, n16823, n16824,
    n16825, n16826, n16827, n16828, n16829, n16830,
    n16831, n16832, n16833, n16834, n16835, n16836,
    n16837, n16838, n16839, n16840, n16841, n16842,
    n16843, n16844, n16845, n16846, n16847, n16848,
    n16849, n16850, n16851, n16852, n16853, n16854,
    n16855, n16856, n16857, n16858, n16859, n16860,
    n16861, n16862, n16863, n16864, n16865, n16866,
    n16867, n16868, n16869, n16870, n16871, n16872,
    n16873, n16874, n16875, n16876, n16877, n16878,
    n16879, n16880, n16881, n16882, n16883, n16884,
    n16885, n16886, n16887, n16888, n16889, n16890,
    n16891, n16892, n16893, n16894, n16895, n16896,
    n16897, n16898, n16899, n16900, n16901, n16902,
    n16903, n16904, n16905, n16906, n16907, n16908,
    n16909, n16910, n16911, n16912, n16913, n16914,
    n16915, n16916, n16917, n16918, n16919, n16920,
    n16921, n16922, n16923, n16924, n16925, n16926,
    n16927, n16928, n16929, n16930, n16931, n16932,
    n16933, n16934, n16935, n16936, n16937, n16938,
    n16939, n16940, n16941, n16942, n16943, n16944,
    n16945, n16946, n16947, n16948, n16949, n16950,
    n16951, n16952, n16953, n16954, n16955, n16956,
    n16957, n16958, n16959, n16960, n16961, n16962,
    n16963, n16964, n16965, n16966, n16967, n16968,
    n16969, n16970, n16971, n16972, n16973, n16974,
    n16975, n16976, n16977, n16978, n16979, n16980,
    n16981, n16982, n16983, n16984, n16985, n16986,
    n16987, n16988, n16989, n16990, n16991, n16992,
    n16993, n16994, n16995, n16996, n16997, n16998,
    n16999, n17000, n17001, n17002, n17003, n17004,
    n17005, n17006, n17007, n17008, n17009, n17010,
    n17011, n17012, n17013, n17014, n17015, n17016,
    n17017, n17018, n17019, n17020, n17021, n17022,
    n17023, n17024, n17025, n17026, n17027, n17028,
    n17029, n17030, n17031, n17032, n17033, n17034,
    n17035, n17036, n17037, n17038, n17039, n17040,
    n17041, n17042, n17043, n17044, n17045, n17046,
    n17047, n17048, n17049, n17050, n17051, n17053,
    n17054, n17055, n17056, n17057, n17058, n17059,
    n17060, n17061, n17062, n17063, n17064, n17065,
    n17066, n17067, n17068, n17069, n17070, n17071,
    n17072, n17073, n17074, n17075, n17076, n17077,
    n17078, n17079, n17080, n17081, n17082, n17083,
    n17084, n17085, n17086, n17087, n17088, n17089,
    n17090, n17091, n17092, n17093, n17094, n17095,
    n17096, n17097, n17098, n17099, n17100, n17101,
    n17102, n17103, n17104, n17105, n17106, n17107,
    n17108, n17109, n17110, n17111, n17112, n17113,
    n17114, n17115, n17116, n17117, n17118, n17119,
    n17120, n17121, n17122, n17123, n17124, n17125,
    n17126, n17127, n17128, n17129, n17130, n17131,
    n17132, n17133, n17134, n17135, n17136, n17137,
    n17138, n17139, n17140, n17141, n17142, n17143,
    n17144, n17145, n17146, n17147, n17148, n17149,
    n17150, n17151, n17152, n17153, n17154, n17155,
    n17156, n17157, n17158, n17159, n17160, n17161,
    n17162, n17163, n17164, n17165, n17166, n17167,
    n17168, n17169, n17170, n17171, n17172, n17173,
    n17174, n17175, n17176, n17177, n17178, n17179,
    n17180, n17181, n17182, n17183, n17184, n17185,
    n17186, n17187, n17188, n17189, n17190, n17191,
    n17192, n17193, n17194, n17195, n17196, n17197,
    n17198, n17199, n17200, n17201, n17202, n17203,
    n17204, n17205, n17206, n17207, n17208, n17209,
    n17210, n17211, n17212, n17213, n17214, n17215,
    n17216, n17217, n17218, n17219, n17220, n17221,
    n17222, n17223, n17224, n17225, n17226, n17227,
    n17228, n17229, n17230, n17231, n17232, n17233,
    n17234, n17235, n17236, n17237, n17238, n17239,
    n17240, n17241, n17242, n17243, n17244, n17245,
    n17246, n17247, n17248, n17249, n17250, n17251,
    n17252, n17253, n17254, n17255, n17256, n17257,
    n17258, n17259, n17260, n17261, n17262, n17263,
    n17264, n17265, n17266, n17267, n17268, n17269,
    n17270, n17271, n17272, n17273, n17274, n17275,
    n17276, n17277, n17278, n17279, n17280, n17281,
    n17282, n17283, n17284, n17285, n17286, n17287,
    n17288, n17289, n17290, n17291, n17292, n17293,
    n17294, n17295, n17296, n17297, n17298, n17299,
    n17300, n17301, n17302, n17303, n17304, n17305,
    n17306, n17307, n17308, n17309, n17310, n17311,
    n17312, n17313, n17314, n17315, n17316, n17317,
    n17318, n17319, n17320, n17321, n17322, n17323,
    n17324, n17325, n17326, n17327, n17328, n17329,
    n17330, n17331, n17332, n17333, n17334, n17335,
    n17336, n17337, n17338, n17339, n17340, n17341,
    n17342, n17343, n17344, n17345, n17346, n17347,
    n17348, n17349, n17350, n17351, n17352, n17353,
    n17354, n17355, n17356, n17357, n17358, n17359,
    n17360, n17361, n17362, n17363, n17364, n17365,
    n17366, n17367, n17368, n17369, n17370, n17371,
    n17372, n17373, n17374, n17375, n17376, n17377,
    n17378, n17379, n17380, n17381, n17382, n17383,
    n17384, n17385, n17386, n17387, n17388, n17389,
    n17390, n17391, n17392, n17393, n17394, n17395,
    n17396, n17397, n17398, n17399, n17400, n17401,
    n17402, n17403, n17404, n17405, n17406, n17407,
    n17408, n17409, n17410, n17411, n17412, n17413,
    n17414, n17415, n17416, n17417, n17418, n17419,
    n17420, n17421, n17422, n17423, n17424, n17425,
    n17426, n17427, n17428, n17429, n17430, n17431,
    n17432, n17433, n17434, n17435, n17436, n17437,
    n17438, n17439, n17440, n17441, n17442, n17443,
    n17444, n17445, n17446, n17447, n17448, n17449,
    n17450, n17451, n17452, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461,
    n17462, n17463, n17464, n17465, n17466, n17467,
    n17468, n17469, n17470, n17471, n17472, n17473,
    n17474, n17475, n17476, n17477, n17478, n17479,
    n17480, n17481, n17482, n17483, n17484, n17485,
    n17486, n17487, n17488, n17489, n17490, n17491,
    n17492, n17493, n17494, n17495, n17496, n17497,
    n17498, n17499, n17500, n17501, n17502, n17503,
    n17504, n17505, n17506, n17507, n17508, n17509,
    n17510, n17511, n17512, n17513, n17514, n17515,
    n17516, n17517, n17518, n17519, n17520, n17521,
    n17522, n17523, n17524, n17525, n17526, n17527,
    n17528, n17529, n17530, n17531, n17532, n17533,
    n17534, n17535, n17536, n17537, n17538, n17539,
    n17540, n17541, n17542, n17543, n17544, n17545,
    n17546, n17547, n17548, n17549, n17550, n17551,
    n17552, n17553, n17554, n17555, n17556, n17557,
    n17558, n17559, n17560, n17561, n17562, n17563,
    n17564, n17565, n17566, n17567, n17568, n17569,
    n17570, n17571, n17572, n17573, n17574, n17575,
    n17576, n17577, n17578, n17579, n17580, n17581,
    n17582, n17583, n17584, n17585, n17586, n17587,
    n17588, n17589, n17590, n17591, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600,
    n17601, n17602, n17603, n17604, n17605, n17606,
    n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618,
    n17619, n17620, n17621, n17622, n17623, n17624,
    n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636,
    n17637, n17638, n17639, n17640, n17641, n17642,
    n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654,
    n17655, n17656, n17657, n17658, n17659, n17660,
    n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672,
    n17673, n17674, n17675, n17676, n17677, n17678,
    n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690,
    n17691, n17692, n17693, n17694, n17695, n17696,
    n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708,
    n17709, n17710, n17711, n17712, n17713, n17714,
    n17715, n17716, n17717, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726,
    n17727, n17728, n17729, n17730, n17731, n17732,
    n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744,
    n17745, n17746, n17747, n17748, n17749, n17750,
    n17751, n17752, n17753, n17754, n17755, n17756,
    n17757, n17758, n17759, n17760, n17761, n17762,
    n17763, n17764, n17765, n17766, n17767, n17768,
    n17769, n17770, n17771, n17772, n17773, n17774,
    n17775, n17776, n17777, n17778, n17779, n17780,
    n17781, n17782, n17783, n17784, n17785, n17786,
    n17787, n17788, n17789, n17790, n17791, n17792,
    n17793, n17794, n17795, n17796, n17797, n17798,
    n17799, n17800, n17801, n17802, n17803, n17804,
    n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17813, n17814, n17815, n17816,
    n17817, n17818, n17819, n17820, n17821, n17822,
    n17823, n17824, n17825, n17826, n17827, n17828,
    n17829, n17830, n17831, n17832, n17833, n17834,
    n17835, n17836, n17837, n17838, n17839, n17840,
    n17841, n17842, n17843, n17844, n17845, n17846,
    n17847, n17848, n17849, n17850, n17851, n17852,
    n17853, n17854, n17855, n17856, n17857, n17858,
    n17859, n17860, n17861, n17862, n17863, n17864,
    n17865, n17866, n17867, n17868, n17869, n17870,
    n17871, n17872, n17873, n17874, n17875, n17876,
    n17877, n17878, n17879, n17880, n17881, n17882,
    n17883, n17884, n17885, n17886, n17887, n17888,
    n17889, n17890, n17891, n17892, n17893, n17894,
    n17895, n17896, n17897, n17898, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906,
    n17907, n17908, n17909, n17910, n17911, n17912,
    n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17921, n17922, n17923, n17924,
    n17925, n17926, n17927, n17928, n17929, n17930,
    n17931, n17932, n17933, n17934, n17935, n17936,
    n17937, n17938, n17939, n17940, n17941, n17942,
    n17943, n17944, n17945, n17946, n17947, n17948,
    n17949, n17950, n17951, n17952, n17953, n17954,
    n17955, n17956, n17957, n17958, n17959, n17960,
    n17961, n17962, n17963, n17964, n17965, n17966,
    n17967, n17968, n17969, n17970, n17971, n17972,
    n17973, n17974, n17975, n17976, n17977, n17978,
    n17979, n17980, n17981, n17982, n17983, n17984,
    n17985, n17986, n17987, n17988, n17989, n17990,
    n17991, n17992, n17993, n17994, n17995, n17996,
    n17997, n17998, n17999, n18000, n18001, n18002,
    n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014,
    n18015, n18016, n18017, n18018, n18019, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032,
    n18033, n18034, n18035, n18036, n18037, n18038,
    n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050,
    n18051, n18052, n18053, n18054, n18055, n18056,
    n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068,
    n18069, n18070, n18071, n18072, n18073, n18074,
    n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086,
    n18087, n18088, n18089, n18090, n18091, n18092,
    n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104,
    n18105, n18106, n18107, n18108, n18109, n18110,
    n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122,
    n18123, n18124, n18125, n18126, n18127, n18128,
    n18129, n18130, n18131, n18133, n18134, n18135,
    n18136, n18137, n18138, n18139, n18140, n18141,
    n18142, n18143, n18144, n18145, n18146, n18147,
    n18148, n18149, n18150, n18151, n18152, n18153,
    n18154, n18155, n18156, n18157, n18158, n18159,
    n18160, n18161, n18162, n18163, n18164, n18165,
    n18166, n18167, n18168, n18169, n18170, n18171,
    n18172, n18173, n18174, n18175, n18176, n18177,
    n18178, n18179, n18180, n18181, n18182, n18183,
    n18184, n18185, n18186, n18187, n18188, n18189,
    n18190, n18191, n18192, n18193, n18194, n18195,
    n18196, n18197, n18198, n18199, n18200, n18201,
    n18202, n18203, n18204, n18205, n18206, n18207,
    n18208, n18209, n18210, n18211, n18212, n18213,
    n18214, n18215, n18216, n18217, n18218, n18219,
    n18220, n18221, n18222, n18223, n18224, n18225,
    n18226, n18227, n18228, n18229, n18230, n18231,
    n18232, n18233, n18234, n18235, n18236, n18237,
    n18238, n18239, n18240, n18241, n18242, n18243,
    n18244, n18245, n18246, n18247, n18248, n18249,
    n18250, n18251, n18252, n18253, n18254, n18255,
    n18256, n18257, n18258, n18259, n18260, n18261,
    n18262, n18263, n18264, n18265, n18266, n18267,
    n18268, n18269, n18270, n18271, n18272, n18273,
    n18274, n18275, n18276, n18277, n18278, n18279,
    n18280, n18281, n18282, n18283, n18284, n18285,
    n18286, n18287, n18288, n18289, n18290, n18291,
    n18292, n18293, n18294, n18295, n18296, n18297,
    n18298, n18299, n18300, n18301, n18302, n18303,
    n18304, n18305, n18306, n18307, n18308, n18309,
    n18310, n18311, n18312, n18313, n18314, n18315,
    n18316, n18317, n18318, n18319, n18320, n18321,
    n18322, n18323, n18324, n18325, n18326, n18327,
    n18328, n18329, n18330, n18331, n18332, n18333,
    n18334, n18335, n18336, n18337, n18338, n18339,
    n18340, n18341, n18342, n18343, n18344, n18345,
    n18346, n18347, n18348, n18349, n18350, n18351,
    n18352, n18353, n18354, n18355, n18356, n18357,
    n18358, n18359, n18360, n18361, n18362, n18363,
    n18364, n18365, n18366, n18367, n18368, n18369,
    n18370, n18371, n18372, n18373, n18374, n18375,
    n18376, n18377, n18378, n18379, n18380, n18381,
    n18382, n18383, n18384, n18385, n18386, n18387,
    n18388, n18389, n18390, n18391, n18392, n18393,
    n18394, n18395, n18396, n18397, n18398, n18399,
    n18400, n18401, n18402, n18403, n18404, n18405,
    n18406, n18407, n18408, n18409, n18410, n18411,
    n18412, n18413, n18414, n18415, n18416, n18417,
    n18418, n18419, n18420, n18421, n18422, n18423,
    n18424, n18425, n18426, n18427, n18428, n18429,
    n18430, n18431, n18432, n18433, n18434, n18435,
    n18436, n18437, n18438, n18439, n18440, n18441,
    n18442, n18443, n18444, n18445, n18446, n18447,
    n18448, n18449, n18450, n18451, n18452, n18453,
    n18454, n18455, n18456, n18457, n18458, n18459,
    n18460, n18461, n18462, n18463, n18464, n18465,
    n18466, n18467, n18468, n18469, n18470, n18471,
    n18472, n18473, n18474, n18475, n18476, n18477,
    n18478, n18479, n18480, n18481, n18482, n18483,
    n18484, n18485, n18486, n18487, n18488, n18489,
    n18490, n18491, n18492, n18493, n18494, n18495,
    n18496, n18497, n18498, n18499, n18500, n18501,
    n18502, n18503, n18504, n18505, n18506, n18507,
    n18508, n18509, n18510, n18511, n18512, n18513,
    n18514, n18515, n18516, n18517, n18518, n18519,
    n18520, n18521, n18522, n18523, n18524, n18525,
    n18526, n18527, n18528, n18529, n18530, n18531,
    n18532, n18533, n18534, n18535, n18536, n18537,
    n18538, n18539, n18540, n18541, n18542, n18543,
    n18544, n18545, n18546, n18547, n18548, n18549,
    n18550, n18551, n18552, n18553, n18554, n18555,
    n18556, n18557, n18558, n18559, n18560, n18561,
    n18562, n18563, n18564, n18565, n18566, n18567,
    n18568, n18569, n18570, n18571, n18572, n18573,
    n18574, n18575, n18576, n18577, n18578, n18579,
    n18580, n18581, n18582, n18583, n18584, n18585,
    n18586, n18587, n18588, n18589, n18590, n18591,
    n18592, n18593, n18594, n18595, n18596, n18597,
    n18598, n18599, n18600, n18601, n18602, n18603,
    n18604, n18605, n18606, n18607, n18608, n18609,
    n18610, n18611, n18612, n18613, n18614, n18615,
    n18616, n18617, n18618, n18619, n18620, n18621,
    n18622, n18623, n18624, n18625, n18626, n18627,
    n18628, n18629, n18630, n18631, n18632, n18633,
    n18634, n18635, n18636, n18637, n18638, n18639,
    n18640, n18641, n18642, n18643, n18644, n18645,
    n18646, n18647, n18648, n18649, n18650, n18651,
    n18652, n18653, n18654, n18655, n18656, n18657,
    n18658, n18659, n18660, n18661, n18662, n18663,
    n18664, n18665, n18666, n18667, n18668, n18669,
    n18670, n18671, n18672, n18674, n18675, n18676,
    n18677, n18678, n18679, n18680, n18681, n18682,
    n18683, n18684, n18685, n18686, n18687, n18688,
    n18689, n18690, n18691, n18692, n18693, n18694,
    n18695, n18696, n18697, n18698, n18699, n18700,
    n18701, n18702, n18703, n18704, n18705, n18706,
    n18707, n18708, n18709, n18710, n18711, n18712,
    n18713, n18714, n18715, n18716, n18717, n18718,
    n18719, n18720, n18721, n18722, n18723, n18724,
    n18725, n18726, n18727, n18728, n18729, n18730,
    n18731, n18732, n18733, n18734, n18735, n18736,
    n18737, n18738, n18739, n18740, n18741, n18742,
    n18743, n18744, n18745, n18746, n18747, n18748,
    n18749, n18750, n18751, n18752, n18753, n18754,
    n18755, n18756, n18757, n18758, n18759, n18760,
    n18761, n18762, n18763, n18764, n18765, n18766,
    n18767, n18768, n18769, n18770, n18771, n18772,
    n18773, n18774, n18775, n18776, n18777, n18778,
    n18779, n18780, n18781, n18782, n18783, n18784,
    n18785, n18786, n18787, n18788, n18789, n18790,
    n18791, n18792, n18793, n18794, n18795, n18796,
    n18797, n18798, n18799, n18800, n18801, n18802,
    n18803, n18804, n18805, n18806, n18807, n18808,
    n18809, n18810, n18811, n18812, n18813, n18814,
    n18815, n18816, n18817, n18818, n18819, n18820,
    n18821, n18822, n18823, n18824, n18825, n18826,
    n18827, n18828, n18829, n18830, n18831, n18832,
    n18833, n18834, n18835, n18836, n18837, n18838,
    n18839, n18840, n18841, n18842, n18843, n18844,
    n18845, n18846, n18847, n18848, n18849, n18850,
    n18851, n18852, n18853, n18854, n18855, n18856,
    n18857, n18858, n18859, n18860, n18861, n18862,
    n18863, n18864, n18865, n18866, n18867, n18868,
    n18869, n18870, n18871, n18872, n18873, n18874,
    n18875, n18876, n18877, n18878, n18879, n18880,
    n18881, n18882, n18883, n18884, n18885, n18886,
    n18887, n18888, n18889, n18890, n18891, n18892,
    n18893, n18894, n18895, n18896, n18897, n18898,
    n18899, n18900, n18901, n18902, n18903, n18904,
    n18905, n18906, n18907, n18908, n18909, n18910,
    n18911, n18912, n18913, n18914, n18915, n18916,
    n18917, n18918, n18919, n18920, n18921, n18922,
    n18923, n18924, n18925, n18926, n18927, n18928,
    n18929, n18930, n18931, n18932, n18933, n18934,
    n18935, n18936, n18937, n18938, n18939, n18940,
    n18941, n18942, n18943, n18944, n18945, n18946,
    n18947, n18948, n18949, n18950, n18951, n18952,
    n18953, n18954, n18955, n18956, n18957, n18958,
    n18959, n18960, n18961, n18962, n18963, n18964,
    n18965, n18966, n18967, n18968, n18969, n18970,
    n18971, n18972, n18973, n18974, n18975, n18976,
    n18977, n18978, n18979, n18980, n18981, n18982,
    n18983, n18984, n18985, n18986, n18987, n18988,
    n18989, n18990, n18991, n18992, n18993, n18994,
    n18995, n18996, n18997, n18998, n18999, n19000,
    n19001, n19002, n19003, n19004, n19005, n19006,
    n19007, n19008, n19009, n19010, n19011, n19012,
    n19013, n19014, n19015, n19016, n19017, n19018,
    n19019, n19020, n19021, n19022, n19023, n19024,
    n19025, n19026, n19027, n19028, n19029, n19030,
    n19031, n19032, n19033, n19034, n19035, n19036,
    n19037, n19038, n19039, n19040, n19041, n19042,
    n19043, n19044, n19045, n19046, n19047, n19048,
    n19049, n19050, n19051, n19052, n19053, n19054,
    n19055, n19056, n19057, n19058, n19059, n19060,
    n19061, n19062, n19063, n19064, n19065, n19066,
    n19067, n19068, n19069, n19070, n19071, n19072,
    n19073, n19074, n19075, n19076, n19077, n19078,
    n19079, n19080, n19081, n19082, n19083, n19084,
    n19085, n19086, n19087, n19088, n19089, n19090,
    n19091, n19092, n19093, n19094, n19095, n19096,
    n19097, n19098, n19099, n19100, n19101, n19102,
    n19103, n19104, n19105, n19106, n19107, n19108,
    n19109, n19110, n19111, n19112, n19113, n19114,
    n19115, n19116, n19117, n19118, n19119, n19120,
    n19121, n19122, n19123, n19124, n19125, n19126,
    n19127, n19128, n19129, n19130, n19131, n19132,
    n19133, n19134, n19135, n19136, n19137, n19138,
    n19139, n19140, n19141, n19142, n19143, n19144,
    n19145, n19146, n19147, n19148, n19149, n19150,
    n19151, n19152, n19153, n19154, n19155, n19156,
    n19157, n19158, n19159, n19160, n19161, n19162,
    n19163, n19164, n19165, n19166, n19167, n19168,
    n19169, n19170, n19171, n19172, n19173, n19174,
    n19175, n19176, n19177, n19178, n19179, n19180,
    n19181, n19182, n19183, n19184, n19185, n19186,
    n19187, n19188, n19189, n19190, n19191, n19192,
    n19193, n19194, n19195, n19196, n19197, n19198,
    n19199, n19200, n19201, n19202, n19203, n19204,
    n19205, n19206, n19207, n19208, n19209, n19210,
    n19211, n19212, n19213, n19214, n19215, n19216,
    n19217, n19218, n19219, n19220, n19221, n19222,
    n19223, n19224, n19225, n19226, n19227, n19228,
    n19229, n19230, n19231, n19232, n19233, n19234,
    n19235, n19236, n19237, n19238, n19239, n19240,
    n19241, n19242, n19243, n19244, n19245, n19246,
    n19247, n19248, n19249, n19250, n19251, n19252,
    n19253, n19254, n19255, n19257, n19258, n19259,
    n19260, n19261, n19262, n19263, n19264, n19265,
    n19266, n19267, n19268, n19269, n19270, n19271,
    n19272, n19273, n19274, n19275, n19276, n19277,
    n19278, n19279, n19280, n19281, n19282, n19283,
    n19284, n19285, n19286, n19287, n19288, n19289,
    n19290, n19291, n19292, n19293, n19294, n19295,
    n19296, n19297, n19298, n19299, n19300, n19301,
    n19302, n19303, n19304, n19305, n19306, n19307,
    n19308, n19309, n19310, n19311, n19312, n19313,
    n19314, n19315, n19316, n19317, n19318, n19319,
    n19320, n19321, n19322, n19323, n19324, n19325,
    n19326, n19327, n19328, n19329, n19330, n19331,
    n19332, n19333, n19334, n19335, n19336, n19337,
    n19338, n19339, n19340, n19341, n19342, n19343,
    n19344, n19345, n19346, n19347, n19348, n19349,
    n19350, n19351, n19352, n19353, n19354, n19355,
    n19356, n19357, n19358, n19359, n19360, n19361,
    n19362, n19363, n19364, n19365, n19366, n19367,
    n19368, n19369, n19370, n19371, n19372, n19373,
    n19374, n19375, n19376, n19377, n19378, n19379,
    n19380, n19381, n19382, n19383, n19384, n19385,
    n19386, n19387, n19388, n19389, n19390, n19391,
    n19392, n19393, n19394, n19395, n19396, n19397,
    n19398, n19399, n19400, n19401, n19402, n19403,
    n19404, n19405, n19406, n19407, n19408, n19409,
    n19410, n19411, n19412, n19413, n19414, n19415,
    n19416, n19417, n19418, n19419, n19420, n19421,
    n19422, n19423, n19424, n19425, n19426, n19427,
    n19428, n19429, n19430, n19431, n19432, n19433,
    n19434, n19435, n19436, n19437, n19438, n19439,
    n19440, n19441, n19442, n19443, n19444, n19445,
    n19446, n19447, n19448, n19449, n19450, n19451,
    n19452, n19453, n19454, n19455, n19456, n19457,
    n19458, n19459, n19460, n19461, n19462, n19463,
    n19464, n19465, n19466, n19467, n19468, n19469,
    n19470, n19471, n19472, n19473, n19474, n19475,
    n19476, n19477, n19478, n19479, n19480, n19481,
    n19482, n19483, n19484, n19485, n19486, n19487,
    n19488, n19489, n19490, n19491, n19492, n19493,
    n19494, n19495, n19496, n19497, n19498, n19499,
    n19500, n19501, n19502, n19503, n19504, n19505,
    n19506, n19507, n19508, n19509, n19510, n19511,
    n19512, n19513, n19514, n19515, n19516, n19517,
    n19518, n19519, n19520, n19521, n19522, n19523,
    n19524, n19525, n19526, n19527, n19528, n19529,
    n19530, n19531, n19532, n19533, n19534, n19535,
    n19536, n19537, n19538, n19539, n19540, n19541,
    n19542, n19543, n19544, n19545, n19546, n19547,
    n19548, n19549, n19550, n19551, n19552, n19553,
    n19554, n19555, n19556, n19557, n19558, n19559,
    n19560, n19561, n19562, n19563, n19564, n19565,
    n19566, n19567, n19568, n19569, n19570, n19571,
    n19572, n19573, n19574, n19575, n19576, n19577,
    n19578, n19579, n19580, n19581, n19582, n19583,
    n19584, n19585, n19586, n19587, n19588, n19589,
    n19590, n19591, n19592, n19593, n19594, n19595,
    n19596, n19597, n19598, n19599, n19600, n19601,
    n19602, n19603, n19604, n19605, n19606, n19607,
    n19608, n19609, n19610, n19611, n19612, n19613,
    n19614, n19615, n19616, n19617, n19618, n19619,
    n19620, n19621, n19622, n19623, n19624, n19625,
    n19626, n19627, n19628, n19629, n19630, n19631,
    n19632, n19633, n19634, n19635, n19636, n19637,
    n19638, n19639, n19640, n19641, n19642, n19643,
    n19644, n19645, n19646, n19647, n19648, n19649,
    n19650, n19651, n19652, n19653, n19654, n19655,
    n19656, n19657, n19658, n19659, n19660, n19661,
    n19662, n19663, n19664, n19665, n19666, n19667,
    n19668, n19669, n19670, n19671, n19672, n19673,
    n19674, n19675, n19676, n19677, n19678, n19679,
    n19680, n19681, n19682, n19683, n19684, n19685,
    n19686, n19687, n19688, n19689, n19690, n19691,
    n19692, n19693, n19694, n19695, n19696, n19697,
    n19698, n19699, n19700, n19701, n19702, n19703,
    n19704, n19705, n19706, n19707, n19708, n19709,
    n19710, n19711, n19712, n19713, n19714, n19715,
    n19716, n19717, n19718, n19719, n19720, n19721,
    n19722, n19723, n19724, n19725, n19726, n19727,
    n19728, n19729, n19730, n19731, n19732, n19733,
    n19734, n19735, n19736, n19737, n19738, n19739,
    n19740, n19741, n19742, n19743, n19744, n19745,
    n19746, n19747, n19748, n19749, n19750, n19751,
    n19752, n19753, n19754, n19755, n19756, n19757,
    n19758, n19759, n19760, n19761, n19762, n19763,
    n19764, n19765, n19766, n19767, n19768, n19769,
    n19770, n19771, n19772, n19773, n19774, n19775,
    n19776, n19777, n19778, n19779, n19780, n19781,
    n19782, n19783, n19784, n19785, n19786, n19787,
    n19788, n19789, n19790, n19791, n19792, n19793,
    n19794, n19795, n19796, n19797, n19798, n19799,
    n19800, n19801, n19802, n19803, n19804, n19805,
    n19806, n19807, n19808, n19809, n19810, n19811,
    n19812, n19813, n19814, n19815, n19816, n19817,
    n19818, n19819, n19820, n19821, n19822, n19823,
    n19824, n19825, n19826, n19827, n19828, n19829,
    n19830, n19831, n19832, n19833, n19834, n19835,
    n19836, n19837, n19838, n19839, n19840, n19841,
    n19842, n19843, n19844, n19845, n19846, n19848,
    n19849, n19850, n19851, n19852, n19853, n19854,
    n19855, n19856, n19857, n19858, n19859, n19860,
    n19861, n19862, n19863, n19864, n19865, n19866,
    n19867, n19868, n19869, n19870, n19871, n19872,
    n19873, n19874, n19875, n19876, n19877, n19878,
    n19879, n19880, n19881, n19882, n19883, n19884,
    n19885, n19886, n19887, n19888, n19889, n19890,
    n19891, n19892, n19893, n19894, n19895, n19896,
    n19897, n19898, n19899, n19900, n19901, n19902,
    n19903, n19904, n19905, n19906, n19907, n19908,
    n19909, n19910, n19911, n19912, n19913, n19914,
    n19915, n19916, n19917, n19918, n19919, n19920,
    n19921, n19922, n19923, n19924, n19925, n19926,
    n19927, n19928, n19929, n19930, n19931, n19932,
    n19933, n19934, n19935, n19936, n19937, n19938,
    n19939, n19940, n19941, n19942, n19943, n19944,
    n19945, n19946, n19947, n19948, n19949, n19950,
    n19951, n19952, n19953, n19954, n19955, n19956,
    n19957, n19958, n19959, n19960, n19961, n19962,
    n19963, n19964, n19965, n19966, n19967, n19968,
    n19969, n19970, n19971, n19972, n19973, n19974,
    n19975, n19976, n19977, n19978, n19979, n19980,
    n19981, n19982, n19983, n19984, n19985, n19986,
    n19987, n19988, n19989, n19990, n19991, n19992,
    n19993, n19994, n19995, n19996, n19997, n19998,
    n19999, n20000, n20001, n20002, n20003, n20004,
    n20005, n20006, n20007, n20008, n20009, n20010,
    n20011, n20012, n20013, n20014, n20015, n20016,
    n20017, n20018, n20019, n20020, n20021, n20022,
    n20023, n20024, n20025, n20026, n20027, n20028,
    n20029, n20030, n20031, n20032, n20033, n20034,
    n20035, n20036, n20037, n20038, n20039, n20040,
    n20041, n20042, n20043, n20044, n20045, n20046,
    n20047, n20048, n20049, n20050, n20051, n20052,
    n20053, n20054, n20055, n20056, n20057, n20058,
    n20059, n20060, n20061, n20062, n20063, n20064,
    n20065, n20066, n20067, n20068, n20069, n20070,
    n20071, n20072, n20073, n20074, n20075, n20076,
    n20077, n20078, n20079, n20080, n20081, n20082,
    n20083, n20084, n20085, n20086, n20087, n20088,
    n20089, n20090, n20091, n20092, n20093, n20094,
    n20095, n20096, n20097, n20098, n20099, n20100,
    n20101, n20102, n20103, n20104, n20105, n20106,
    n20107, n20108, n20109, n20110, n20111, n20112,
    n20113, n20114, n20115, n20116, n20117, n20118,
    n20119, n20120, n20121, n20122, n20123, n20124,
    n20125, n20126, n20127, n20128, n20129, n20130,
    n20131, n20132, n20133, n20134, n20135, n20136,
    n20137, n20138, n20139, n20140, n20141, n20142,
    n20143, n20144, n20145, n20146, n20147, n20148,
    n20149, n20150, n20151, n20152, n20153, n20154,
    n20155, n20156, n20157, n20158, n20159, n20160,
    n20161, n20162, n20163, n20164, n20165, n20166,
    n20167, n20168, n20169, n20170, n20171, n20172,
    n20173, n20174, n20175, n20176, n20177, n20178,
    n20179, n20180, n20181, n20182, n20183, n20184,
    n20185, n20186, n20187, n20188, n20189, n20190,
    n20191, n20192, n20193, n20194, n20195, n20196,
    n20197, n20198, n20199, n20200, n20201, n20202,
    n20203, n20204, n20205, n20206, n20207, n20208,
    n20209, n20210, n20211, n20212, n20213, n20214,
    n20215, n20216, n20217, n20218, n20219, n20220,
    n20221, n20222, n20223, n20224, n20225, n20226,
    n20227, n20228, n20229, n20230, n20231, n20232,
    n20233, n20234, n20235, n20236, n20237, n20238,
    n20239, n20240, n20241, n20242, n20243, n20244,
    n20245, n20246, n20247, n20248, n20249, n20250,
    n20251, n20252, n20253, n20254, n20255, n20256,
    n20257, n20258, n20259, n20260, n20261, n20262,
    n20263, n20264, n20265, n20266, n20267, n20268,
    n20269, n20270, n20271, n20272, n20273, n20274,
    n20275, n20276, n20277, n20278, n20279, n20280,
    n20281, n20282, n20283, n20284, n20285, n20286,
    n20287, n20288, n20289, n20290, n20291, n20292,
    n20293, n20294, n20295, n20296, n20297, n20298,
    n20299, n20300, n20301, n20302, n20303, n20304,
    n20305, n20306, n20307, n20308, n20309, n20310,
    n20311, n20312, n20313, n20314, n20315, n20316,
    n20317, n20318, n20319, n20320, n20321, n20322,
    n20323, n20324, n20325, n20326, n20327, n20328,
    n20329, n20330, n20331, n20332, n20333, n20334,
    n20335, n20336, n20337, n20338, n20339, n20340,
    n20341, n20342, n20343, n20344, n20345, n20346,
    n20347, n20348, n20349, n20350, n20351, n20352,
    n20353, n20354, n20355, n20356, n20357, n20358,
    n20359, n20360, n20361, n20362, n20363, n20364,
    n20365, n20366, n20367, n20368, n20369, n20370,
    n20371, n20372, n20373, n20374, n20375, n20376,
    n20377, n20378, n20379, n20380, n20381, n20382,
    n20383, n20384, n20385, n20386, n20387, n20388,
    n20389, n20390, n20391, n20392, n20393, n20394,
    n20395, n20396, n20397, n20398, n20399, n20400,
    n20401, n20402, n20403, n20404, n20405, n20406,
    n20407, n20408, n20409, n20410, n20411, n20412,
    n20413, n20414, n20415, n20416, n20417, n20418,
    n20419, n20420, n20421, n20422, n20423, n20424,
    n20425, n20426, n20427, n20428, n20429, n20430,
    n20431, n20432, n20433, n20434, n20435, n20436,
    n20437, n20439, n20440, n20441, n20442, n20443,
    n20444, n20445, n20446, n20447, n20448, n20449,
    n20450, n20451, n20452, n20453, n20454, n20455,
    n20456, n20457, n20458, n20459, n20460, n20461,
    n20462, n20463, n20464, n20465, n20466, n20467,
    n20468, n20469, n20470, n20471, n20472, n20473,
    n20474, n20475, n20476, n20477, n20478, n20479,
    n20480, n20481, n20482, n20483, n20484, n20485,
    n20486, n20487, n20488, n20489, n20490, n20491,
    n20492, n20493, n20494, n20495, n20496, n20497,
    n20498, n20499, n20500, n20501, n20502, n20503,
    n20504, n20505, n20506, n20507, n20508, n20509,
    n20510, n20511, n20512, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521,
    n20522, n20523, n20524, n20525, n20526, n20527,
    n20528, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539,
    n20540, n20541, n20542, n20543, n20544, n20545,
    n20546, n20547, n20548, n20549, n20550, n20551,
    n20552, n20553, n20554, n20555, n20556, n20557,
    n20558, n20559, n20560, n20561, n20562, n20563,
    n20564, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581,
    n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599,
    n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617,
    n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20631, n20632, n20633, n20634, n20635,
    n20636, n20637, n20638, n20639, n20640, n20641,
    n20642, n20643, n20644, n20645, n20646, n20647,
    n20648, n20649, n20650, n20651, n20652, n20653,
    n20654, n20655, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665,
    n20666, n20667, n20668, n20669, n20670, n20671,
    n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683,
    n20684, n20685, n20686, n20687, n20688, n20689,
    n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701,
    n20702, n20703, n20704, n20705, n20706, n20707,
    n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719,
    n20720, n20721, n20722, n20723, n20724, n20725,
    n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737,
    n20738, n20739, n20740, n20741, n20742, n20743,
    n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755,
    n20756, n20757, n20758, n20759, n20760, n20761,
    n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773,
    n20774, n20775, n20776, n20777, n20778, n20779,
    n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20789, n20790, n20791,
    n20792, n20793, n20794, n20795, n20796, n20797,
    n20798, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809,
    n20810, n20811, n20812, n20813, n20814, n20815,
    n20816, n20817, n20818, n20819, n20820, n20821,
    n20822, n20823, n20824, n20825, n20826, n20827,
    n20828, n20829, n20830, n20831, n20832, n20833,
    n20834, n20835, n20836, n20837, n20838, n20839,
    n20840, n20841, n20842, n20843, n20844, n20845,
    n20846, n20847, n20848, n20849, n20850, n20851,
    n20852, n20853, n20854, n20855, n20856, n20857,
    n20858, n20859, n20860, n20861, n20862, n20863,
    n20864, n20865, n20866, n20867, n20868, n20869,
    n20870, n20871, n20872, n20873, n20874, n20875,
    n20876, n20877, n20878, n20879, n20880, n20881,
    n20882, n20883, n20884, n20885, n20886, n20887,
    n20888, n20889, n20890, n20891, n20892, n20893,
    n20894, n20895, n20896, n20897, n20898, n20899,
    n20900, n20901, n20902, n20903, n20904, n20905,
    n20906, n20907, n20908, n20909, n20910, n20911,
    n20912, n20913, n20914, n20915, n20916, n20917,
    n20918, n20919, n20920, n20921, n20922, n20923,
    n20924, n20925, n20926, n20927, n20928, n20929,
    n20930, n20931, n20932, n20933, n20934, n20935,
    n20936, n20937, n20938, n20939, n20940, n20941,
    n20942, n20943, n20944, n20945, n20946, n20947,
    n20948, n20949, n20950, n20951, n20952, n20953,
    n20954, n20955, n20956, n20957, n20958, n20959,
    n20960, n20961, n20962, n20963, n20964, n20965,
    n20966, n20967, n20968, n20969, n20970, n20971,
    n20972, n20973, n20974, n20975, n20976, n20977,
    n20978, n20979, n20980, n20981, n20982, n20983,
    n20984, n20985, n20986, n20987, n20988, n20989,
    n20990, n20991, n20992, n20993, n20994, n20995,
    n20996, n20997, n20998, n20999, n21000, n21001,
    n21002, n21003, n21004, n21005, n21006, n21007,
    n21008, n21009, n21010, n21011, n21012, n21013,
    n21014, n21015, n21016, n21017, n21019, n21020,
    n21021, n21022, n21023, n21024, n21025, n21026,
    n21027, n21028, n21029, n21030, n21031, n21032,
    n21033, n21034, n21035, n21036, n21037, n21038,
    n21039, n21040, n21041, n21042, n21043, n21044,
    n21045, n21046, n21047, n21048, n21049, n21050,
    n21051, n21052, n21053, n21054, n21055, n21056,
    n21057, n21058, n21059, n21060, n21061, n21062,
    n21063, n21064, n21065, n21066, n21067, n21068,
    n21069, n21070, n21071, n21072, n21073, n21074,
    n21075, n21076, n21077, n21078, n21079, n21080,
    n21081, n21082, n21083, n21084, n21085, n21086,
    n21087, n21088, n21089, n21090, n21091, n21092,
    n21093, n21094, n21095, n21096, n21097, n21098,
    n21099, n21100, n21101, n21102, n21103, n21104,
    n21105, n21106, n21107, n21108, n21109, n21110,
    n21111, n21112, n21113, n21114, n21115, n21116,
    n21117, n21118, n21119, n21120, n21121, n21122,
    n21123, n21124, n21125, n21126, n21127, n21128,
    n21129, n21130, n21131, n21132, n21133, n21134,
    n21135, n21136, n21137, n21138, n21139, n21140,
    n21141, n21142, n21143, n21144, n21145, n21146,
    n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158,
    n21159, n21160, n21161, n21162, n21163, n21164,
    n21165, n21166, n21167, n21168, n21169, n21170,
    n21171, n21172, n21173, n21174, n21175, n21176,
    n21177, n21178, n21179, n21180, n21181, n21182,
    n21183, n21184, n21185, n21186, n21187, n21188,
    n21189, n21190, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200,
    n21201, n21202, n21203, n21204, n21205, n21206,
    n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218,
    n21219, n21220, n21221, n21222, n21223, n21224,
    n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236,
    n21237, n21238, n21239, n21240, n21241, n21242,
    n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254,
    n21255, n21256, n21257, n21258, n21259, n21260,
    n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21268, n21269, n21270, n21271, n21272,
    n21273, n21274, n21275, n21276, n21277, n21278,
    n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290,
    n21291, n21292, n21293, n21294, n21295, n21296,
    n21297, n21298, n21299, n21300, n21301, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308,
    n21309, n21310, n21311, n21312, n21313, n21314,
    n21315, n21316, n21317, n21318, n21319, n21320,
    n21321, n21322, n21323, n21324, n21325, n21326,
    n21327, n21328, n21329, n21330, n21331, n21332,
    n21333, n21334, n21335, n21336, n21337, n21338,
    n21339, n21340, n21341, n21342, n21343, n21344,
    n21345, n21346, n21347, n21348, n21349, n21350,
    n21351, n21352, n21353, n21354, n21355, n21356,
    n21357, n21358, n21359, n21360, n21361, n21362,
    n21363, n21364, n21365, n21366, n21367, n21368,
    n21369, n21370, n21371, n21372, n21373, n21374,
    n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386,
    n21387, n21388, n21389, n21390, n21391, n21392,
    n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410,
    n21411, n21412, n21413, n21414, n21415, n21416,
    n21417, n21418, n21419, n21420, n21421, n21422,
    n21423, n21424, n21425, n21426, n21427, n21428,
    n21429, n21430, n21431, n21432, n21433, n21434,
    n21435, n21436, n21437, n21438, n21439, n21440,
    n21441, n21442, n21443, n21444, n21445, n21446,
    n21447, n21448, n21449, n21450, n21451, n21452,
    n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21463, n21464,
    n21465, n21466, n21467, n21468, n21469, n21470,
    n21471, n21472, n21473, n21474, n21475, n21476,
    n21477, n21478, n21479, n21480, n21481, n21482,
    n21483, n21484, n21485, n21486, n21487, n21488,
    n21489, n21490, n21491, n21492, n21493, n21494,
    n21495, n21496, n21497, n21498, n21499, n21500,
    n21501, n21502, n21503, n21504, n21505, n21506,
    n21507, n21508, n21509, n21510, n21511, n21512,
    n21513, n21514, n21515, n21516, n21517, n21518,
    n21519, n21520, n21521, n21522, n21523, n21524,
    n21525, n21526, n21527, n21528, n21529, n21530,
    n21531, n21532, n21533, n21534, n21535, n21536,
    n21537, n21538, n21539, n21540, n21541, n21542,
    n21543, n21544, n21545, n21546, n21547, n21548,
    n21549, n21550, n21551, n21552, n21553, n21554,
    n21555, n21556, n21557, n21558, n21559, n21560,
    n21561, n21562, n21563, n21564, n21565, n21566,
    n21568, n21569, n21570, n21571, n21572, n21573,
    n21574, n21575, n21576, n21577, n21578, n21579,
    n21580, n21581, n21582, n21583, n21584, n21585,
    n21586, n21587, n21588, n21589, n21590, n21591,
    n21592, n21593, n21594, n21595, n21596, n21597,
    n21598, n21599, n21600, n21601, n21602, n21603,
    n21604, n21605, n21606, n21607, n21608, n21609,
    n21610, n21611, n21612, n21613, n21614, n21615,
    n21616, n21617, n21618, n21619, n21620, n21621,
    n21622, n21623, n21624, n21625, n21626, n21627,
    n21628, n21629, n21630, n21631, n21632, n21633,
    n21634, n21635, n21636, n21637, n21638, n21639,
    n21640, n21641, n21642, n21643, n21644, n21645,
    n21646, n21647, n21648, n21649, n21650, n21651,
    n21652, n21653, n21654, n21655, n21656, n21657,
    n21658, n21659, n21660, n21661, n21662, n21663,
    n21664, n21665, n21666, n21667, n21668, n21669,
    n21670, n21671, n21672, n21673, n21674, n21675,
    n21676, n21677, n21678, n21679, n21680, n21681,
    n21682, n21683, n21684, n21685, n21686, n21687,
    n21688, n21689, n21690, n21691, n21692, n21693,
    n21694, n21695, n21696, n21697, n21698, n21699,
    n21700, n21701, n21702, n21703, n21704, n21705,
    n21706, n21707, n21708, n21709, n21710, n21711,
    n21712, n21713, n21714, n21715, n21716, n21717,
    n21718, n21719, n21720, n21721, n21722, n21723,
    n21724, n21725, n21726, n21727, n21728, n21729,
    n21730, n21731, n21732, n21733, n21734, n21735,
    n21736, n21737, n21738, n21739, n21740, n21741,
    n21742, n21743, n21744, n21745, n21746, n21747,
    n21748, n21749, n21750, n21751, n21752, n21753,
    n21754, n21755, n21756, n21757, n21758, n21759,
    n21760, n21761, n21762, n21763, n21764, n21765,
    n21766, n21767, n21768, n21769, n21770, n21771,
    n21772, n21773, n21774, n21775, n21776, n21777,
    n21778, n21779, n21780, n21781, n21782, n21783,
    n21784, n21785, n21786, n21787, n21788, n21789,
    n21790, n21791, n21792, n21793, n21794, n21795,
    n21796, n21797, n21798, n21799, n21800, n21801,
    n21802, n21803, n21804, n21805, n21806, n21807,
    n21808, n21809, n21810, n21811, n21812, n21813,
    n21814, n21815, n21816, n21817, n21818, n21819,
    n21820, n21821, n21822, n21823, n21824, n21825,
    n21826, n21827, n21828, n21829, n21830, n21831,
    n21832, n21833, n21834, n21835, n21836, n21837,
    n21838, n21839, n21840, n21841, n21842, n21843,
    n21844, n21845, n21846, n21847, n21848, n21849,
    n21850, n21851, n21852, n21853, n21854, n21855,
    n21856, n21857, n21858, n21859, n21860, n21861,
    n21862, n21863, n21864, n21865, n21866, n21867,
    n21868, n21869, n21870, n21871, n21872, n21873,
    n21874, n21875, n21876, n21877, n21878, n21879,
    n21880, n21881, n21882, n21883, n21884, n21885,
    n21886, n21887, n21888, n21889, n21890, n21891,
    n21892, n21893, n21894, n21895, n21896, n21897,
    n21898, n21899, n21900, n21901, n21902, n21903,
    n21904, n21905, n21906, n21907, n21908, n21909,
    n21910, n21911, n21912, n21913, n21914, n21915,
    n21916, n21917, n21918, n21919, n21920, n21921,
    n21922, n21923, n21924, n21925, n21926, n21927,
    n21928, n21929, n21930, n21931, n21932, n21933,
    n21934, n21935, n21936, n21937, n21938, n21939,
    n21940, n21941, n21942, n21943, n21944, n21945,
    n21946, n21947, n21948, n21949, n21950, n21951,
    n21952, n21953, n21954, n21955, n21956, n21957,
    n21958, n21959, n21960, n21961, n21962, n21963,
    n21964, n21965, n21966, n21967, n21968, n21969,
    n21970, n21971, n21972, n21973, n21974, n21975,
    n21976, n21977, n21978, n21979, n21980, n21981,
    n21982, n21983, n21984, n21985, n21986, n21987,
    n21988, n21989, n21990, n21991, n21992, n21993,
    n21994, n21995, n21996, n21997, n21998, n21999,
    n22000, n22001, n22002, n22003, n22004, n22005,
    n22006, n22007, n22008, n22009, n22010, n22011,
    n22012, n22013, n22014, n22015, n22016, n22017,
    n22018, n22019, n22020, n22021, n22022, n22023,
    n22024, n22025, n22026, n22027, n22028, n22029,
    n22030, n22031, n22032, n22033, n22034, n22035,
    n22036, n22037, n22038, n22039, n22040, n22041,
    n22042, n22043, n22044, n22045, n22046, n22047,
    n22048, n22049, n22050, n22051, n22052, n22053,
    n22054, n22055, n22056, n22057, n22058, n22059,
    n22060, n22061, n22062, n22063, n22064, n22065,
    n22066, n22067, n22068, n22069, n22070, n22071,
    n22072, n22073, n22074, n22075, n22076, n22077,
    n22078, n22079, n22080, n22081, n22082, n22083,
    n22084, n22085, n22086, n22087, n22088, n22089,
    n22090, n22091, n22092, n22093, n22094, n22095,
    n22096, n22097, n22098, n22099, n22100, n22101,
    n22102, n22103, n22104, n22105, n22106, n22107,
    n22108, n22109, n22110, n22111, n22112, n22113,
    n22114, n22115, n22117, n22118, n22119, n22120,
    n22121, n22122, n22123, n22124, n22125, n22126,
    n22127, n22128, n22129, n22130, n22131, n22132,
    n22133, n22134, n22135, n22136, n22137, n22138,
    n22139, n22140, n22141, n22142, n22143, n22144,
    n22145, n22146, n22147, n22148, n22149, n22150,
    n22151, n22152, n22153, n22154, n22155, n22156,
    n22157, n22158, n22159, n22160, n22161, n22162,
    n22163, n22164, n22165, n22166, n22167, n22168,
    n22169, n22170, n22171, n22172, n22173, n22174,
    n22175, n22176, n22177, n22178, n22179, n22180,
    n22181, n22182, n22183, n22184, n22185, n22186,
    n22187, n22188, n22189, n22190, n22191, n22192,
    n22193, n22194, n22195, n22196, n22197, n22198,
    n22199, n22200, n22201, n22202, n22203, n22204,
    n22205, n22206, n22207, n22208, n22209, n22210,
    n22211, n22212, n22213, n22214, n22215, n22216,
    n22217, n22218, n22219, n22220, n22221, n22222,
    n22223, n22224, n22225, n22226, n22227, n22228,
    n22229, n22230, n22231, n22232, n22233, n22234,
    n22235, n22236, n22237, n22238, n22239, n22240,
    n22241, n22242, n22243, n22244, n22245, n22246,
    n22247, n22248, n22249, n22250, n22251, n22252,
    n22253, n22254, n22255, n22256, n22257, n22258,
    n22259, n22260, n22261, n22262, n22263, n22264,
    n22265, n22266, n22267, n22268, n22269, n22270,
    n22271, n22272, n22273, n22274, n22275, n22276,
    n22277, n22278, n22279, n22280, n22281, n22282,
    n22283, n22284, n22285, n22286, n22287, n22288,
    n22289, n22290, n22291, n22292, n22293, n22294,
    n22295, n22296, n22297, n22298, n22299, n22300,
    n22301, n22302, n22303, n22304, n22305, n22306,
    n22307, n22308, n22309, n22310, n22311, n22312,
    n22313, n22314, n22315, n22316, n22317, n22318,
    n22319, n22320, n22321, n22322, n22323, n22324,
    n22325, n22326, n22327, n22328, n22329, n22330,
    n22331, n22332, n22333, n22334, n22335, n22336,
    n22337, n22338, n22339, n22340, n22341, n22342,
    n22343, n22344, n22345, n22346, n22347, n22348,
    n22349, n22350, n22351, n22352, n22353, n22354,
    n22355, n22356, n22357, n22358, n22359, n22360,
    n22361, n22362, n22363, n22364, n22365, n22366,
    n22367, n22368, n22369, n22370, n22371, n22372,
    n22373, n22374, n22375, n22376, n22377, n22378,
    n22379, n22380, n22381, n22382, n22383, n22384,
    n22385, n22386, n22387, n22388, n22389, n22390,
    n22391, n22392, n22393, n22394, n22395, n22396,
    n22397, n22398, n22399, n22400, n22401, n22402,
    n22403, n22404, n22405, n22406, n22407, n22408,
    n22409, n22410, n22411, n22412, n22413, n22414,
    n22415, n22416, n22417, n22418, n22419, n22420,
    n22421, n22422, n22423, n22424, n22425, n22426,
    n22427, n22428, n22429, n22430, n22431, n22432,
    n22433, n22434, n22435, n22436, n22437, n22438,
    n22439, n22440, n22441, n22442, n22443, n22444,
    n22445, n22446, n22447, n22448, n22449, n22450,
    n22451, n22452, n22453, n22454, n22455, n22456,
    n22457, n22458, n22459, n22460, n22461, n22462,
    n22463, n22464, n22465, n22466, n22467, n22468,
    n22469, n22470, n22471, n22472, n22473, n22474,
    n22475, n22476, n22477, n22478, n22479, n22480,
    n22481, n22482, n22483, n22484, n22485, n22486,
    n22487, n22488, n22489, n22490, n22491, n22492,
    n22493, n22494, n22495, n22496, n22497, n22498,
    n22499, n22500, n22501, n22502, n22503, n22504,
    n22505, n22506, n22507, n22508, n22509, n22510,
    n22511, n22512, n22513, n22514, n22515, n22516,
    n22517, n22518, n22519, n22520, n22521, n22522,
    n22523, n22524, n22525, n22526, n22527, n22528,
    n22529, n22530, n22531, n22532, n22533, n22534,
    n22535, n22536, n22537, n22538, n22539, n22540,
    n22541, n22542, n22543, n22544, n22545, n22546,
    n22547, n22548, n22549, n22550, n22551, n22552,
    n22553, n22554, n22555, n22556, n22557, n22558,
    n22559, n22560, n22561, n22562, n22563, n22564,
    n22565, n22566, n22567, n22568, n22569, n22570,
    n22571, n22572, n22573, n22574, n22575, n22576,
    n22577, n22578, n22579, n22580, n22581, n22582,
    n22583, n22584, n22585, n22586, n22587, n22588,
    n22589, n22590, n22591, n22592, n22593, n22594,
    n22595, n22596, n22597, n22598, n22599, n22600,
    n22601, n22602, n22603, n22604, n22605, n22606,
    n22607, n22608, n22609, n22610, n22611, n22612,
    n22613, n22614, n22615, n22616, n22617, n22618,
    n22619, n22620, n22621, n22622, n22623, n22624,
    n22625, n22626, n22627, n22628, n22629, n22630,
    n22631, n22632, n22633, n22634, n22635, n22636,
    n22637, n22638, n22639, n22640, n22641, n22642,
    n22643, n22644, n22645, n22646, n22647, n22648,
    n22649, n22650, n22651, n22652, n22653, n22654,
    n22655, n22656, n22657, n22658, n22659, n22660,
    n22661, n22662, n22663, n22664, n22666, n22667,
    n22668, n22669, n22670, n22671, n22672, n22673,
    n22674, n22675, n22676, n22677, n22678, n22679,
    n22680, n22681, n22682, n22683, n22684, n22685,
    n22686, n22687, n22688, n22689, n22690, n22691,
    n22692, n22693, n22694, n22695, n22696, n22697,
    n22698, n22699, n22700, n22701, n22702, n22703,
    n22704, n22705, n22706, n22707, n22708, n22709,
    n22710, n22711, n22712, n22713, n22714, n22715,
    n22716, n22717, n22718, n22719, n22720, n22721,
    n22722, n22723, n22724, n22725, n22726, n22727,
    n22728, n22729, n22730, n22731, n22732, n22733,
    n22734, n22735, n22736, n22737, n22738, n22739,
    n22740, n22741, n22742, n22743, n22744, n22745,
    n22746, n22747, n22748, n22749, n22750, n22751,
    n22752, n22753, n22754, n22755, n22756, n22757,
    n22758, n22759, n22760, n22761, n22762, n22763,
    n22764, n22765, n22766, n22767, n22768, n22769,
    n22770, n22771, n22772, n22773, n22774, n22775,
    n22776, n22777, n22778, n22779, n22780, n22781,
    n22782, n22783, n22784, n22785, n22786, n22787,
    n22788, n22789, n22790, n22791, n22792, n22793,
    n22794, n22795, n22796, n22797, n22798, n22799,
    n22800, n22801, n22802, n22803, n22804, n22805,
    n22806, n22807, n22808, n22809, n22810, n22811,
    n22812, n22813, n22814, n22815, n22816, n22817,
    n22818, n22819, n22820, n22821, n22822, n22823,
    n22824, n22825, n22826, n22827, n22828, n22829,
    n22830, n22831, n22832, n22833, n22834, n22835,
    n22836, n22837, n22838, n22839, n22840, n22841,
    n22842, n22843, n22844, n22845, n22846, n22847,
    n22848, n22849, n22850, n22851, n22852, n22853,
    n22854, n22855, n22856, n22857, n22858, n22859,
    n22860, n22861, n22862, n22863, n22864, n22865,
    n22866, n22867, n22868, n22869, n22870, n22871,
    n22872, n22873, n22874, n22875, n22876, n22877,
    n22878, n22879, n22880, n22881, n22882, n22883,
    n22884, n22885, n22886, n22887, n22888, n22889,
    n22890, n22891, n22892, n22893, n22894, n22895,
    n22896, n22897, n22898, n22899, n22900, n22901,
    n22902, n22903, n22904, n22905, n22906, n22907,
    n22908, n22909, n22910, n22911, n22912, n22913,
    n22914, n22915, n22916, n22917, n22918, n22919,
    n22920, n22921, n22922, n22923, n22924, n22925,
    n22926, n22927, n22928, n22929, n22930, n22931,
    n22932, n22933, n22934, n22935, n22936, n22937,
    n22938, n22939, n22940, n22941, n22942, n22943,
    n22944, n22945, n22946, n22947, n22948, n22949,
    n22950, n22951, n22952, n22953, n22954, n22955,
    n22956, n22957, n22958, n22959, n22960, n22961,
    n22962, n22963, n22964, n22965, n22966, n22967,
    n22968, n22969, n22970, n22971, n22972, n22973,
    n22974, n22975, n22976, n22977, n22978, n22979,
    n22980, n22981, n22982, n22983, n22984, n22985,
    n22986, n22987, n22988, n22989, n22990, n22991,
    n22992, n22993, n22994, n22995, n22996, n22997,
    n22998, n22999, n23000, n23001, n23002, n23003,
    n23004, n23005, n23006, n23007, n23008, n23009,
    n23010, n23011, n23012, n23013, n23014, n23015,
    n23016, n23017, n23018, n23019, n23020, n23021,
    n23022, n23023, n23024, n23025, n23026, n23027,
    n23028, n23029, n23030, n23031, n23032, n23033,
    n23034, n23035, n23036, n23037, n23038, n23039,
    n23040, n23041, n23042, n23043, n23044, n23045,
    n23046, n23047, n23048, n23049, n23050, n23051,
    n23052, n23053, n23054, n23055, n23056, n23057,
    n23058, n23059, n23060, n23061, n23062, n23063,
    n23064, n23065, n23066, n23067, n23068, n23069,
    n23070, n23071, n23072, n23073, n23074, n23075,
    n23076, n23077, n23078, n23079, n23080, n23081,
    n23082, n23083, n23084, n23085, n23086, n23087,
    n23088, n23089, n23090, n23091, n23092, n23093,
    n23094, n23095, n23096, n23097, n23098, n23099,
    n23100, n23101, n23102, n23103, n23104, n23105,
    n23106, n23107, n23108, n23109, n23110, n23111,
    n23112, n23113, n23114, n23115, n23116, n23117,
    n23118, n23119, n23120, n23121, n23122, n23123,
    n23124, n23125, n23126, n23127, n23128, n23129,
    n23130, n23131, n23132, n23133, n23134, n23135,
    n23136, n23137, n23138, n23139, n23140, n23141,
    n23142, n23143, n23144, n23145, n23146, n23147,
    n23148, n23149, n23150, n23151, n23152, n23153,
    n23154, n23155, n23156, n23157, n23158, n23159,
    n23160, n23161, n23162, n23163, n23164, n23165,
    n23166, n23167, n23168, n23169, n23170, n23171,
    n23172, n23173, n23174, n23175, n23176, n23177,
    n23178, n23179, n23180, n23181, n23182, n23183,
    n23184, n23185, n23186, n23187, n23188, n23189,
    n23190, n23191, n23192, n23193, n23194, n23195,
    n23196, n23197, n23198, n23199, n23201, n23202,
    n23203, n23204, n23205, n23206, n23207, n23208,
    n23209, n23210, n23211, n23212, n23213, n23214,
    n23215, n23216, n23217, n23218, n23219, n23220,
    n23221, n23222, n23223, n23224, n23225, n23226,
    n23227, n23228, n23229, n23230, n23231, n23232,
    n23233, n23234, n23235, n23236, n23237, n23238,
    n23239, n23240, n23241, n23242, n23243, n23244,
    n23245, n23246, n23247, n23248, n23249, n23250,
    n23251, n23252, n23253, n23254, n23255, n23256,
    n23257, n23258, n23259, n23260, n23261, n23262,
    n23263, n23264, n23265, n23266, n23267, n23268,
    n23269, n23270, n23271, n23272, n23273, n23274,
    n23275, n23276, n23277, n23278, n23279, n23280,
    n23281, n23282, n23283, n23284, n23285, n23286,
    n23287, n23288, n23289, n23290, n23291, n23292,
    n23293, n23294, n23295, n23296, n23297, n23298,
    n23299, n23300, n23301, n23302, n23303, n23304,
    n23305, n23306, n23307, n23308, n23309, n23310,
    n23311, n23312, n23313, n23314, n23315, n23316,
    n23317, n23318, n23319, n23320, n23321, n23322,
    n23323, n23324, n23325, n23326, n23327, n23328,
    n23329, n23330, n23331, n23332, n23333, n23334,
    n23335, n23336, n23337, n23338, n23339, n23340,
    n23341, n23342, n23343, n23344, n23345, n23346,
    n23347, n23348, n23349, n23350, n23351, n23352,
    n23353, n23354, n23355, n23356, n23357, n23358,
    n23359, n23360, n23361, n23362, n23363, n23364,
    n23365, n23366, n23367, n23368, n23369, n23370,
    n23371, n23372, n23373, n23374, n23375, n23376,
    n23377, n23378, n23379, n23380, n23381, n23382,
    n23383, n23384, n23385, n23386, n23387, n23388,
    n23389, n23390, n23391, n23392, n23393, n23394,
    n23395, n23396, n23397, n23398, n23399, n23400,
    n23401, n23402, n23403, n23404, n23405, n23406,
    n23407, n23408, n23409, n23410, n23411, n23412,
    n23413, n23414, n23415, n23416, n23417, n23418,
    n23419, n23420, n23421, n23422, n23423, n23424,
    n23425, n23426, n23427, n23428, n23429, n23430,
    n23431, n23432, n23433, n23434, n23435, n23436,
    n23437, n23438, n23439, n23440, n23441, n23442,
    n23443, n23444, n23445, n23446, n23447, n23448,
    n23449, n23450, n23451, n23452, n23453, n23454,
    n23455, n23456, n23457, n23458, n23459, n23460,
    n23461, n23462, n23463, n23464, n23465, n23466,
    n23467, n23468, n23469, n23470, n23471, n23472,
    n23473, n23474, n23475, n23476, n23477, n23478,
    n23479, n23480, n23481, n23482, n23483, n23484,
    n23485, n23486, n23487, n23488, n23489, n23490,
    n23491, n23492, n23493, n23494, n23495, n23496,
    n23497, n23498, n23499, n23500, n23501, n23502,
    n23503, n23504, n23505, n23506, n23507, n23508,
    n23509, n23510, n23511, n23512, n23513, n23514,
    n23515, n23516, n23517, n23518, n23519, n23520,
    n23521, n23522, n23523, n23524, n23525, n23526,
    n23527, n23528, n23529, n23530, n23531, n23532,
    n23533, n23534, n23535, n23536, n23537, n23538,
    n23539, n23540, n23541, n23542, n23543, n23544,
    n23545, n23546, n23547, n23548, n23549, n23550,
    n23551, n23552, n23553, n23554, n23555, n23556,
    n23557, n23558, n23559, n23560, n23561, n23562,
    n23563, n23564, n23565, n23566, n23567, n23568,
    n23569, n23570, n23571, n23572, n23573, n23574,
    n23575, n23576, n23577, n23578, n23579, n23580,
    n23581, n23582, n23583, n23584, n23585, n23586,
    n23587, n23588, n23589, n23590, n23591, n23592,
    n23593, n23594, n23595, n23596, n23597, n23598,
    n23599, n23600, n23601, n23602, n23603, n23604,
    n23605, n23606, n23607, n23608, n23609, n23610,
    n23611, n23612, n23613, n23614, n23615, n23616,
    n23617, n23618, n23619, n23620, n23621, n23622,
    n23623, n23624, n23625, n23626, n23627, n23628,
    n23629, n23630, n23631, n23632, n23633, n23634,
    n23635, n23636, n23637, n23638, n23639, n23640,
    n23641, n23642, n23643, n23644, n23645, n23646,
    n23647, n23648, n23649, n23650, n23651, n23652,
    n23653, n23654, n23655, n23656, n23657, n23658,
    n23659, n23660, n23661, n23662, n23663, n23664,
    n23665, n23666, n23667, n23668, n23669, n23670,
    n23671, n23672, n23673, n23674, n23675, n23676,
    n23677, n23678, n23679, n23680, n23681, n23682,
    n23683, n23684, n23685, n23686, n23687, n23688,
    n23689, n23690, n23691, n23692, n23693, n23694,
    n23695, n23696, n23697, n23698, n23699, n23700,
    n23701, n23702, n23703, n23704, n23705, n23706,
    n23707, n23708, n23709, n23710, n23711, n23712,
    n23713, n23714, n23715, n23716, n23717, n23718,
    n23719, n23720, n23721, n23722, n23723, n23724,
    n23725, n23726, n23727, n23728, n23729, n23730,
    n23731, n23732, n23733, n23734, n23735, n23736,
    n23737, n23738, n23739, n23740, n23741, n23742,
    n23743, n23744, n23745, n23746, n23747, n23748,
    n23749, n23750, n23751, n23752, n23753, n23754,
    n23755, n23756, n23757, n23758, n23759, n23760,
    n23761, n23762, n23763, n23764, n23765, n23766,
    n23767, n23768, n23769, n23770, n23771, n23772,
    n23773, n23774, n23775, n23776, n23777, n23778,
    n23779, n23780, n23781, n23782, n23783, n23784,
    n23785, n23786, n23787, n23788, n23789, n23790,
    n23791, n23792, n23793, n23794, n23795, n23796,
    n23797, n23798, n23799, n23800, n23801, n23802,
    n23803, n23804, n23805, n23806, n23807, n23808,
    n23809, n23810, n23812, n23813, n23814, n23815,
    n23816, n23817, n23818, n23819, n23820, n23821,
    n23822, n23823, n23824, n23825, n23826, n23827,
    n23828, n23829, n23830, n23831, n23832, n23833,
    n23834, n23835, n23836, n23837, n23838, n23839,
    n23840, n23841, n23842, n23843, n23844, n23845,
    n23846, n23847, n23848, n23849, n23850, n23851,
    n23852, n23853, n23854, n23855, n23856, n23857,
    n23858, n23859, n23860, n23861, n23862, n23863,
    n23864, n23865, n23866, n23867, n23868, n23869,
    n23870, n23871, n23872, n23873, n23874, n23875,
    n23876, n23877, n23878, n23879, n23880, n23881,
    n23882, n23883, n23884, n23885, n23886, n23887,
    n23888, n23889, n23890, n23891, n23892, n23893,
    n23894, n23895, n23896, n23897, n23898, n23899,
    n23900, n23901, n23902, n23903, n23904, n23905,
    n23906, n23907, n23908, n23909, n23910, n23911,
    n23912, n23913, n23914, n23915, n23916, n23917,
    n23918, n23919, n23920, n23921, n23922, n23923,
    n23924, n23925, n23926, n23927, n23928, n23929,
    n23930, n23931, n23932, n23933, n23934, n23935,
    n23936, n23937, n23938, n23939, n23940, n23941,
    n23942, n23943, n23944, n23945, n23946, n23947,
    n23948, n23949, n23950, n23951, n23952, n23953,
    n23954, n23955, n23956, n23957, n23958, n23959,
    n23960, n23961, n23962, n23963, n23964, n23965,
    n23966, n23967, n23968, n23969, n23970, n23971,
    n23972, n23973, n23974, n23975, n23976, n23977,
    n23978, n23979, n23980, n23981, n23982, n23983,
    n23984, n23985, n23986, n23987, n23988, n23989,
    n23990, n23991, n23992, n23993, n23994, n23995,
    n23996, n23997, n23998, n23999, n24000, n24001,
    n24002, n24003, n24004, n24005, n24006, n24007,
    n24008, n24009, n24010, n24011, n24012, n24013,
    n24014, n24015, n24016, n24017, n24018, n24019,
    n24020, n24021, n24022, n24023, n24024, n24025,
    n24026, n24027, n24028, n24029, n24030, n24031,
    n24032, n24033, n24034, n24035, n24036, n24037,
    n24038, n24039, n24040, n24041, n24042, n24043,
    n24044, n24045, n24046, n24047, n24048, n24049,
    n24050, n24051, n24052, n24053, n24054, n24055,
    n24056, n24057, n24058, n24059, n24060, n24061,
    n24062, n24063, n24064, n24065, n24066, n24067,
    n24068, n24069, n24070, n24071, n24072, n24073,
    n24074, n24075, n24076, n24077, n24078, n24079,
    n24080, n24081, n24082, n24083, n24084, n24085,
    n24086, n24087, n24088, n24089, n24090, n24091,
    n24092, n24093, n24094, n24095, n24096, n24097,
    n24098, n24099, n24100, n24101, n24102, n24103,
    n24104, n24105, n24106, n24107, n24108, n24109,
    n24110, n24111, n24112, n24113, n24114, n24115,
    n24116, n24117, n24118, n24119, n24120, n24121,
    n24122, n24123, n24124, n24125, n24126, n24127,
    n24128, n24129, n24130, n24131, n24132, n24133,
    n24134, n24135, n24136, n24137, n24138, n24139,
    n24140, n24141, n24142, n24143, n24144, n24145,
    n24146, n24147, n24148, n24149, n24150, n24151,
    n24152, n24153, n24154, n24155, n24156, n24157,
    n24158, n24159, n24160, n24161, n24162, n24163,
    n24164, n24165, n24166, n24167, n24168, n24169,
    n24170, n24171, n24172, n24173, n24174, n24175,
    n24176, n24177, n24178, n24179, n24180, n24181,
    n24182, n24183, n24184, n24185, n24186, n24187,
    n24188, n24189, n24190, n24191, n24192, n24193,
    n24194, n24195, n24196, n24197, n24198, n24199,
    n24200, n24201, n24202, n24203, n24204, n24205,
    n24206, n24207, n24208, n24209, n24210, n24211,
    n24212, n24213, n24214, n24215, n24216, n24217,
    n24218, n24219, n24220, n24221, n24222, n24223,
    n24224, n24225, n24226, n24227, n24228, n24229,
    n24230, n24231, n24232, n24233, n24234, n24235,
    n24236, n24237, n24238, n24239, n24240, n24241,
    n24242, n24243, n24244, n24245, n24246, n24247,
    n24248, n24249, n24250, n24251, n24252, n24253,
    n24254, n24255, n24256, n24257, n24258, n24259,
    n24260, n24261, n24262, n24263, n24264, n24265,
    n24266, n24267, n24268, n24269, n24270, n24271,
    n24272, n24273, n24274, n24275, n24276, n24277,
    n24278, n24279, n24280, n24281, n24282, n24283,
    n24284, n24285, n24286, n24287, n24288, n24289,
    n24290, n24291, n24292, n24293, n24294, n24295,
    n24296, n24297, n24298, n24299, n24300, n24301,
    n24302, n24303, n24304, n24305, n24306, n24307,
    n24308, n24309, n24310, n24311, n24312, n24313,
    n24314, n24315, n24316, n24317, n24318, n24319,
    n24320, n24321, n24322, n24323, n24324, n24325,
    n24326, n24327, n24328, n24329, n24330, n24331,
    n24332, n24333, n24334, n24335, n24336, n24337,
    n24338, n24339, n24340, n24341, n24342, n24343,
    n24344, n24345, n24346, n24347, n24348, n24349,
    n24350, n24351, n24352, n24353, n24354, n24355,
    n24356, n24357, n24358, n24359, n24360, n24361,
    n24362, n24363, n24364, n24365, n24366, n24367,
    n24368, n24369, n24370, n24371, n24372, n24373,
    n24374, n24375, n24376, n24377, n24378, n24379,
    n24380, n24381, n24382, n24383, n24384, n24385,
    n24386, n24387, n24388, n24389, n24390, n24391,
    n24392, n24393, n24394, n24395, n24396, n24397,
    n24398, n24399, n24400, n24401, n24402, n24403,
    n24404, n24405, n24406, n24407, n24408, n24409,
    n24410, n24411, n24412, n24413, n24414, n24415,
    n24416, n24417, n24418, n24419, n24420, n24421,
    n24422, n24423, n24424, n24425, n24426, n24427,
    n24428, n24429, n24430, n24431, n24432, n24433,
    n24434, n24435, n24436, n24437, n24438, n24439,
    n24440, n24441, n24442, n24443, n24444, n24445,
    n24446, n24447, n24448, n24449, n24450, n24451,
    n24452, n24453, n24454, n24455, n24456, n24457,
    n24458, n24459, n24460, n24461, n24462, n24463,
    n24464, n24465, n24466, n24467, n24468, n24469,
    n24470, n24471, n24472, n24473, n24474, n24475,
    n24476, n24477, n24478, n24479, n24480, n24481,
    n24482, n24483, n24484, n24485, n24486, n24487,
    n24488, n24489, n24490, n24491, n24492, n24493,
    n24494, n24495, n24496, n24497, n24498, n24499,
    n24500, n24501, n24502, n24503, n24504, n24505,
    n24506, n24507, n24508, n24509, n24510, n24511,
    n24512, n24513, n24514, n24515, n24516, n24517,
    n24518, n24519, n24520, n24521, n24522, n24523,
    n24524, n24525, n24526, n24527, n24528, n24529,
    n24530, n24531, n24532, n24533, n24534, n24535,
    n24536, n24537, n24538, n24539, n24540, n24541,
    n24542, n24543, n24544, n24545, n24546, n24547,
    n24548, n24549, n24550, n24551, n24552, n24553,
    n24554, n24555, n24556, n24557, n24558, n24559,
    n24560, n24561, n24562, n24563, n24564, n24565,
    n24566, n24567, n24568, n24569, n24570, n24571,
    n24572, n24573, n24574, n24575, n24576, n24577,
    n24578, n24579, n24580, n24581, n24582, n24583,
    n24584, n24585, n24586, n24587, n24588, n24589,
    n24590, n24591, n24592, n24593, n24594, n24595,
    n24596, n24597, n24598, n24599, n24600, n24601,
    n24602, n24603, n24604, n24605, n24606, n24607,
    n24608, n24609, n24610, n24611, n24612, n24613,
    n24614, n24615, n24616, n24617, n24618, n24619,
    n24620, n24621, n24622, n24623, n24624, n24625,
    n24626, n24627, n24628, n24629, n24630, n24631,
    n24632, n24633, n24634, n24635, n24636, n24637,
    n24638, n24639, n24640, n24641, n24642, n24643,
    n24644, n24645, n24646, n24647, n24648, n24649,
    n24650, n24651, n24652, n24653, n24654, n24655,
    n24656, n24657, n24658, n24659, n24660, n24661,
    n24662, n24663, n24664, n24665, n24666, n24667,
    n24668, n24669, n24670, n24671, n24672, n24673,
    n24674, n24675, n24676, n24677, n24678, n24679,
    n24680, n24681, n24682, n24683, n24684, n24685,
    n24686, n24687, n24688, n24689, n24690, n24691,
    n24692, n24693, n24694, n24695, n24696, n24697,
    n24698, n24699, n24700, n24701, n24702, n24703,
    n24704, n24705, n24706, n24707, n24708, n24709,
    n24710, n24711, n24712, n24713, n24714, n24715,
    n24716, n24717, n24718, n24719, n24720, n24721,
    n24722, n24723, n24724, n24725, n24726, n24727,
    n24728, n24729, n24730, n24731, n24732, n24733,
    n24734, n24735, n24736, n24737, n24738, n24739,
    n24740, n24741, n24742, n24743, n24744, n24745,
    n24746, n24747, n24748, n24749, n24750, n24751,
    n24752, n24753, n24754, n24755, n24756, n24757,
    n24758, n24759, n24760, n24761, n24762, n24763,
    n24764, n24765, n24766, n24767, n24768, n24769,
    n24770, n24771, n24772, n24773, n24774, n24775,
    n24776, n24777, n24778, n24779, n24780, n24781,
    n24782, n24783, n24784, n24785, n24786, n24787,
    n24788, n24789, n24790, n24791, n24792, n24793,
    n24794, n24795, n24796, n24797, n24798, n24799,
    n24800, n24801, n24802, n24803, n24804, n24805,
    n24806, n24807, n24808, n24809, n24810, n24811,
    n24812, n24813, n24814, n24815, n24816, n24817,
    n24818, n24819, n24820, n24821, n24822, n24823,
    n24824, n24825, n24826, n24827, n24828, n24829,
    n24830, n24831, n24832, n24833, n24834, n24835,
    n24836, n24837, n24838, n24839, n24840, n24841,
    n24842, n24843, n24844, n24845, n24846, n24847,
    n24848, n24849, n24850, n24851, n24852, n24853,
    n24854, n24855, n24856, n24857, n24858, n24859,
    n24860, n24861, n24862, n24863, n24864, n24865,
    n24866, n24867, n24868, n24869, n24870, n24871,
    n24872, n24873, n24874, n24875, n24876, n24877,
    n24878, n24879, n24880, n24881, n24882, n24883,
    n24884, n24885, n24886, n24887, n24888, n24889,
    n24890, n24891, n24892, n24893, n24894, n24895,
    n24896, n24897, n24898, n24899, n24900, n24901,
    n24902, n24903, n24904, n24905, n24906, n24907,
    n24908, n24909, n24910, n24911, n24912, n24913,
    n24914, n24915, n24916, n24917, n24918, n24919,
    n24920, n24921, n24922, n24923, n24924, n24925,
    n24926, n24927, n24928, n24929, n24930, n24931,
    n24932, n24933, n24934, n24935, n24936, n24937,
    n24938, n24939, n24940, n24941, n24942, n24943,
    n24944, n24945, n24946, n24947, n24948, n24949,
    n24950, n24951, n24952, n24953, n24954, n24955,
    n24956, n24957, n24958, n24959, n24960, n24961,
    n24962, n24963, n24964, n24965, n24966, n24967,
    n24968, n24969, n24970, n24971, n24972, n24973,
    n24974, n24975, n24976, n24977, n24978, n24979,
    n24980, n24981, n24982, n24983, n24984, n24985,
    n24986, n24987, n24988, n24989, n24990, n24991,
    n24992, n24993, n24994, n24995, n24996, n24997,
    n24998, n24999, n25000, n25001, n25002, n25003,
    n25004, n25005, n25006, n25007, n25008, n25009,
    n25010, n25011, n25012, n25013, n25014, n25015,
    n25016, n25017, n25018, n25019, n25020, n25021,
    n25022, n25023, n25024, n25025, n25026, n25027,
    n25028, n25029, n25030, n25031, n25032, n25033,
    n25034, n25035, n25036, n25037, n25038, n25039,
    n25040, n25041, n25042, n25043, n25044, n25045,
    n25046, n25047, n25048, n25049, n25050, n25051,
    n25052, n25053, n25054, n25055, n25056, n25057,
    n25058, n25059, n25060, n25061, n25062, n25063,
    n25064, n25065, n25066, n25067, n25068, n25069,
    n25070, n25071, n25072, n25073, n25074, n25075,
    n25076, n25077, n25078, n25079, n25080, n25081,
    n25082, n25083, n25084, n25085, n25086, n25087,
    n25088, n25089, n25090, n25091, n25092, n25093,
    n25094, n25095, n25096, n25097, n25098, n25099,
    n25100, n25101, n25102, n25103, n25104, n25105,
    n25106, n25107, n25108, n25109, n25110, n25111,
    n25112, n25113, n25114, n25115, n25116, n25117,
    n25118, n25119, n25120, n25121, n25122, n25123,
    n25124, n25125, n25126, n25127, n25128, n25129,
    n25130, n25131, n25132, n25133, n25134, n25135,
    n25136, n25137, n25138, n25139, n25140, n25141,
    n25142, n25143, n25144, n25145, n25146, n25147,
    n25148, n25149, n25150, n25151, n25152, n25153,
    n25154, n25155, n25156, n25157, n25158, n25159,
    n25160, n25161, n25162, n25163, n25164, n25165,
    n25166, n25167, n25168, n25169, n25170, n25171,
    n25172, n25173, n25174, n25175, n25176, n25177,
    n25178, n25179, n25180, n25181, n25182, n25183,
    n25184, n25185, n25186, n25187, n25188, n25189,
    n25190, n25191, n25192, n25193, n25194, n25195,
    n25196, n25197, n25198, n25199, n25200, n25201,
    n25202, n25203, n25204, n25205, n25206, n25207,
    n25208, n25209, n25210, n25211, n25212, n25213,
    n25214, n25215, n25216, n25217, n25218, n25219,
    n25220, n25221, n25222, n25223, n25224, n25225,
    n25226, n25227, n25228, n25229, n25230, n25231,
    n25232, n25233, n25234, n25235, n25236, n25237,
    n25238, n25239, n25240, n25241, n25242, n25243,
    n25244, n25245, n25246, n25247, n25248, n25249,
    n25250, n25251, n25252, n25253, n25254, n25255,
    n25256, n25257, n25258, n25259, n25260, n25261,
    n25262, n25263, n25264, n25265, n25266, n25267,
    n25268, n25269, n25270, n25271, n25272, n25273,
    n25274, n25275, n25276, n25277, n25278, n25279,
    n25280, n25281, n25282, n25283, n25284, n25285,
    n25286, n25287, n25288, n25289, n25290, n25291,
    n25292, n25293, n25294, n25295, n25296, n25297,
    n25298, n25299, n25300, n25301, n25302, n25303,
    n25304, n25305, n25306, n25307, n25308, n25309,
    n25310, n25311, n25312, n25313, n25314, n25315,
    n25316, n25317, n25318, n25319, n25320, n25321,
    n25322, n25323, n25324, n25325, n25326, n25327,
    n25328, n25329, n25330, n25331, n25332, n25333,
    n25334, n25335, n25336, n25337, n25338, n25339,
    n25340, n25341, n25342, n25343, n25344, n25345,
    n25346, n25347, n25348, n25349, n25350, n25351,
    n25352, n25353, n25354, n25355, n25356, n25357,
    n25358, n25359, n25360, n25361, n25362, n25363,
    n25364, n25365, n25366, n25367, n25368, n25369,
    n25370, n25371, n25372, n25373, n25374, n25375,
    n25376, n25377, n25378, n25379, n25380, n25381,
    n25382, n25383, n25384, n25385, n25386, n25387,
    n25388, n25389, n25390, n25391, n25392, n25393,
    n25394, n25395, n25396, n25397, n25398, n25399,
    n25400, n25401, n25402, n25403, n25404, n25405,
    n25406, n25407, n25408, n25409, n25410, n25411,
    n25412, n25413, n25414, n25415, n25416, n25417,
    n25418, n25419, n25420, n25421, n25422, n25423,
    n25424, n25425, n25426, n25427, n25428, n25429,
    n25430, n25431, n25432, n25433, n25434, n25435,
    n25436, n25437, n25438, n25439, n25440, n25441,
    n25442, n25443, n25444, n25445, n25446, n25447,
    n25448, n25449, n25450, n25451, n25452, n25453,
    n25454, n25455, n25456, n25457, n25458, n25459,
    n25460, n25461, n25462, n25463, n25464, n25465,
    n25466, n25467, n25468, n25469, n25470, n25471,
    n25472, n25473, n25474, n25475, n25476, n25477,
    n25478, n25479, n25480, n25481, n25482, n25483,
    n25484, n25485, n25486, n25487, n25488, n25489,
    n25490, n25491, n25492, n25493, n25494, n25495,
    n25496, n25497, n25498, n25499, n25500, n25501,
    n25502, n25503, n25504, n25505, n25506, n25507,
    n25508, n25509, n25510, n25511, n25512, n25513,
    n25514, n25515, n25516, n25517, n25518, n25519,
    n25520, n25521, n25522, n25523, n25524, n25525,
    n25526, n25527, n25528, n25529, n25530, n25531,
    n25532, n25533, n25534, n25535, n25536, n25537,
    n25538, n25539, n25540, n25541, n25542, n25543,
    n25544, n25545, n25546, n25547, n25548, n25549,
    n25550, n25551, n25552, n25553, n25554, n25555,
    n25556, n25557, n25558, n25559, n25560, n25561,
    n25562, n25563, n25564, n25565, n25566, n25567,
    n25568, n25569, n25570, n25571, n25572, n25573,
    n25574, n25575, n25576, n25577, n25578, n25579,
    n25580, n25581, n25582, n25583, n25584, n25585,
    n25586, n25587, n25588, n25589, n25590, n25591,
    n25592, n25593, n25594, n25595, n25596, n25597,
    n25598, n25599, n25600, n25601, n25602, n25603,
    n25604, n25605, n25606, n25607, n25608, n25609,
    n25610, n25611, n25612, n25613, n25614, n25615,
    n25616, n25617, n25618, n25619, n25620, n25621,
    n25622, n25623, n25624, n25625, n25626, n25627,
    n25628, n25629, n25630, n25631, n25632, n25633,
    n25634, n25635, n25636, n25637, n25638, n25639,
    n25640, n25641, n25642, n25643, n25644, n25645,
    n25646, n25647, n25648, n25649, n25650, n25651,
    n25652, n25653, n25654, n25655, n25656, n25657,
    n25658, n25659, n25660, n25661, n25662, n25663,
    n25664, n25665, n25666, n25667, n25668, n25669,
    n25670, n25671, n25672, n25673, n25674, n25675,
    n25676, n25677, n25678, n25679, n25680, n25681,
    n25682, n25683, n25684, n25685, n25686, n25687,
    n25688, n25689, n25690, n25691, n25692, n25693,
    n25694, n25695, n25696, n25697, n25698, n25699,
    n25700, n25701, n25702, n25703, n25704, n25705,
    n25706, n25707, n25708, n25709, n25710, n25711,
    n25712, n25713, n25714, n25715, n25716, n25717,
    n25718, n25719, n25720, n25721, n25722, n25723,
    n25724, n25725, n25726, n25727, n25728, n25729,
    n25730, n25731, n25732, n25733, n25734, n25735,
    n25736, n25737, n25738, n25739, n25740, n25741,
    n25742, n25743, n25744, n25745, n25746, n25747,
    n25748, n25749, n25750, n25751, n25752, n25753,
    n25754, n25755, n25756, n25757, n25758, n25759,
    n25760, n25761, n25762, n25763, n25764, n25765,
    n25766, n25767, n25768, n25769, n25770, n25771,
    n25772, n25773, n25774, n25775, n25776, n25777,
    n25778, n25779, n25780, n25781, n25782, n25783,
    n25784, n25785, n25786, n25787, n25788, n25789,
    n25790, n25791, n25792, n25793, n25794, n25795,
    n25796, n25797, n25798, n25799, n25800, n25801,
    n25802, n25803, n25804, n25805, n25806, n25807,
    n25808, n25809, n25810, n25811, n25812, n25813,
    n25814, n25815, n25816, n25817, n25818, n25819,
    n25820, n25821, n25822, n25823, n25824, n25825,
    n25826, n25827, n25828, n25829, n25830, n25831,
    n25832, n25833, n25834, n25835, n25836, n25837,
    n25838, n25839, n25840, n25841, n25842, n25843,
    n25844, n25845, n25846, n25847, n25848, n25849,
    n25850, n25851, n25852, n25853, n25854, n25855,
    n25856, n25857, n25858, n25859, n25860, n25861,
    n25862, n25863, n25864, n25865, n25866, n25867,
    n25868, n25869, n25870, n25871, n25872, n25873,
    n25874, n25875, n25876, n25877, n25878, n25879,
    n25880, n25881, n25882, n25883, n25884, n25885,
    n25886, n25887, n25888, n25889, n25890, n25891,
    n25892, n25893, n25894, n25895, n25896, n25897,
    n25898, n25899, n25900, n25901, n25902, n25903,
    n25904, n25905, n25906, n25907, n25908, n25909,
    n25910, n25911, n25912, n25913, n25914, n25915,
    n25916, n25917, n25918, n25919, n25920, n25921,
    n25922, n25923, n25924, n25925, n25926, n25927,
    n25928, n25929, n25930, n25931, n25932, n25933,
    n25934, n25935, n25936, n25937, n25938, n25939,
    n25940, n25941, n25942, n25943, n25944, n25945,
    n25946, n25947, n25948, n25949, n25950, n25951,
    n25952, n25953, n25954, n25955, n25956, n25957,
    n25958, n25959, n25960, n25961, n25962, n25963,
    n25964, n25965, n25966, n25967, n25968, n25969,
    n25970, n25971, n25972, n25973, n25974, n25975,
    n25976, n25977, n25978, n25979, n25980, n25981,
    n25982, n25983, n25984, n25985, n25986, n25987,
    n25988, n25989, n25990, n25991, n25992, n25993,
    n25994, n25995, n25996, n25997, n25998, n25999,
    n26000, n26001, n26002, n26003, n26004, n26005,
    n26006, n26007, n26008, n26009, n26010, n26011,
    n26012, n26013, n26014, n26015, n26016, n26017,
    n26018, n26019, n26020, n26021, n26022, n26023,
    n26024, n26025, n26026, n26027, n26028, n26029,
    n26030, n26031, n26032, n26033, n26034, n26035,
    n26036, n26037, n26038, n26039, n26040, n26041,
    n26042, n26043, n26044, n26045, n26046, n26047,
    n26048, n26049, n26050, n26051, n26052, n26053,
    n26054, n26055, n26056, n26057, n26058, n26059,
    n26060, n26061, n26062, n26063, n26064, n26065,
    n26066, n26067, n26068, n26069, n26070, n26071,
    n26072, n26073, n26074, n26075, n26076, n26077,
    n26078, n26079, n26080, n26081, n26082, n26083,
    n26084, n26085, n26086, n26087, n26088, n26089,
    n26090, n26091, n26092, n26093, n26094, n26095,
    n26096, n26097, n26098, n26099, n26100, n26101,
    n26102, n26103, n26104, n26105, n26106, n26107,
    n26108, n26109, n26110, n26111, n26112, n26113,
    n26114, n26115, n26116, n26117, n26118, n26119,
    n26120, n26121, n26122, n26123, n26124, n26125,
    n26126, n26127, n26128, n26129, n26130, n26131,
    n26132, n26133, n26134, n26135, n26136, n26137,
    n26138, n26139, n26140, n26141, n26142, n26143,
    n26144, n26145, n26146, n26147, n26148, n26149,
    n26150, n26151, n26152, n26153, n26154, n26155,
    n26156, n26157, n26158, n26159, n26160, n26161,
    n26162, n26163, n26164, n26165, n26166, n26167,
    n26168, n26169, n26170, n26171, n26172, n26173,
    n26174, n26175, n26176, n26177, n26178, n26179,
    n26180, n26181, n26182, n26183, n26184, n26185,
    n26186, n26187, n26188, n26189, n26190, n26191,
    n26192, n26193, n26194, n26195, n26196, n26197,
    n26198, n26199, n26200, n26201, n26202, n26203,
    n26204, n26205, n26206, n26207, n26208, n26209,
    n26210, n26211, n26212, n26213, n26214, n26215,
    n26216, n26217, n26218, n26219, n26220, n26221,
    n26222, n26223, n26224, n26225, n26226, n26227,
    n26228, n26229, n26230, n26231, n26232, n26233,
    n26234, n26235, n26236, n26237, n26238, n26239,
    n26240, n26241, n26242, n26243, n26244, n26245,
    n26246, n26247, n26248, n26249, n26250, n26251,
    n26252, n26253, n26254, n26255, n26256, n26257,
    n26258, n26259, n26260, n26261, n26262, n26263,
    n26264, n26265, n26266, n26267, n26268, n26269,
    n26270, n26271, n26272, n26273, n26274, n26275,
    n26276, n26277, n26278, n26279, n26280, n26281,
    n26282, n26283, n26284, n26285, n26286, n26287,
    n26288, n26289, n26290, n26291, n26292, n26293,
    n26294, n26295, n26296, n26297, n26298, n26299,
    n26300, n26301, n26302, n26303, n26304, n26305,
    n26306, n26307, n26308, n26309, n26310, n26311,
    n26312, n26313, n26314, n26315, n26316, n26317,
    n26318, n26319, n26320, n26321, n26322, n26323,
    n26324, n26325, n26326, n26327, n26328, n26329,
    n26330, n26331, n26332, n26333, n26334, n26335,
    n26336, n26337, n26338, n26339, n26340, n26341,
    n26342, n26343, n26344, n26345, n26346, n26347,
    n26348, n26349, n26350, n26351, n26352, n26353,
    n26354, n26355, n26356, n26357, n26358, n26359,
    n26360, n26361, n26362, n26363, n26364, n26365,
    n26366, n26367, n26368, n26369, n26370, n26371,
    n26372, n26373, n26374, n26375, n26376, n26377,
    n26378, n26379, n26380, n26381, n26382, n26383,
    n26384, n26385, n26386, n26387, n26388, n26389,
    n26390, n26391, n26392, n26393, n26394, n26395,
    n26396, n26397, n26398, n26399, n26400, n26401,
    n26402, n26403, n26404, n26405, n26406, n26407,
    n26408, n26409, n26410, n26411, n26412, n26413,
    n26414, n26415, n26416, n26417, n26418, n26419,
    n26420, n26421, n26422, n26423, n26424, n26425,
    n26426, n26427, n26428, n26429, n26430, n26431,
    n26432, n26433, n26434, n26435, n26436, n26437,
    n26438, n26439, n26440, n26441, n26442, n26443,
    n26444, n26445, n26446, n26447, n26448, n26449,
    n26450, n26451, n26452, n26453, n26454, n26455,
    n26456, n26457, n26458, n26459, n26460, n26461,
    n26462, n26463, n26464, n26465, n26466, n26467,
    n26468, n26469, n26470, n26471, n26472, n26473,
    n26474, n26475, n26476, n26477, n26478, n26479,
    n26480, n26481, n26482, n26483, n26484, n26485,
    n26486, n26487, n26488, n26489, n26490, n26491,
    n26492, n26493, n26494, n26495, n26496, n26497,
    n26498, n26499, n26500, n26501, n26502, n26503,
    n26504, n26505, n26506, n26507, n26508, n26509,
    n26510, n26511, n26512, n26513, n26514, n26515,
    n26516, n26517, n26518, n26519, n26520, n26521,
    n26522, n26523, n26524, n26525, n26526, n26527,
    n26528, n26529, n26530, n26531, n26532, n26533,
    n26534, n26535, n26536, n26537, n26538, n26539,
    n26540, n26541, n26542, n26543, n26544, n26545,
    n26546, n26547, n26548, n26549, n26550, n26551,
    n26552, n26553, n26554, n26555, n26556, n26557,
    n26558, n26559, n26560, n26561, n26562, n26563,
    n26564, n26565, n26566, n26567, n26568, n26569,
    n26570, n26571, n26572, n26573, n26574, n26575,
    n26576, n26577, n26578, n26579, n26580, n26581,
    n26582, n26583, n26584, n26585, n26586, n26587,
    n26588, n26589, n26590, n26591, n26592, n26593,
    n26594, n26595, n26596, n26597, n26598, n26599,
    n26600, n26601, n26602, n26603, n26604, n26605,
    n26606, n26607, n26608, n26609, n26610, n26611,
    n26612, n26613, n26614, n26615, n26616, n26617,
    n26618, n26619, n26620, n26621, n26622, n26623,
    n26624, n26625, n26626, n26627, n26628, n26629,
    n26630, n26631, n26632, n26633, n26634, n26635,
    n26636, n26637, n26638, n26639, n26640, n26641,
    n26642, n26643, n26644, n26645, n26646, n26647,
    n26648, n26649, n26650, n26651, n26652, n26653,
    n26654, n26655, n26656, n26657, n26658, n26659,
    n26660, n26661, n26662, n26663, n26664, n26665,
    n26666, n26667, n26668, n26669, n26670, n26671,
    n26672, n26673, n26674, n26675, n26676, n26677,
    n26678, n26679, n26680, n26681, n26682, n26683,
    n26684, n26685, n26686, n26687, n26688, n26689,
    n26690, n26691, n26692, n26693, n26694, n26695,
    n26696, n26697, n26698, n26699, n26700, n26701,
    n26702, n26703, n26704, n26705, n26706, n26707,
    n26708, n26709, n26710, n26711, n26712, n26713,
    n26714, n26715, n26716, n26717, n26718, n26719,
    n26720, n26721, n26722, n26723, n26724, n26725,
    n26726, n26727, n26728, n26729, n26730, n26731,
    n26732, n26733, n26734, n26735, n26736, n26737,
    n26738, n26739, n26740, n26741, n26742, n26743,
    n26744, n26745, n26746, n26747, n26748, n26749,
    n26750, n26751, n26752, n26753, n26754, n26755,
    n26756, n26757, n26758, n26759, n26760, n26761,
    n26762, n26763, n26764, n26765, n26766, n26767,
    n26768, n26769, n26770, n26771, n26772, n26773,
    n26774, n26775, n26776, n26777, n26778, n26779,
    n26780, n26781, n26782, n26783, n26784, n26785,
    n26786, n26787, n26788, n26789, n26790, n26791,
    n26792, n26793, n26794, n26795, n26796, n26797,
    n26798, n26799, n26800, n26801, n26802, n26803,
    n26804, n26805, n26806, n26807, n26808, n26809,
    n26810, n26811, n26812, n26813, n26814, n26815,
    n26816, n26817, n26818, n26819, n26820, n26821,
    n26822, n26823, n26824, n26825, n26826, n26827,
    n26828, n26829, n26830, n26831, n26832, n26833,
    n26834, n26835, n26836, n26837, n26838, n26839,
    n26840, n26841, n26842, n26843, n26844, n26845,
    n26846, n26847, n26848, n26849, n26850, n26851,
    n26852, n26853, n26854, n26855, n26856, n26857,
    n26858, n26859, n26860, n26861, n26862, n26863,
    n26864, n26865, n26866, n26867, n26868, n26869,
    n26870, n26871, n26872, n26873, n26874, n26875,
    n26876, n26877, n26878, n26879, n26880, n26881,
    n26882, n26883, n26884, n26885, n26886, n26887,
    n26888, n26889, n26890, n26891, n26892, n26893,
    n26894, n26895, n26896, n26897, n26898, n26899,
    n26900, n26901, n26902, n26903, n26904, n26905,
    n26906, n26907, n26908, n26909, n26910, n26911,
    n26912, n26913, n26914, n26915, n26916, n26917,
    n26918, n26919, n26920, n26921, n26922, n26923,
    n26924, n26925, n26926, n26927, n26928, n26929,
    n26930, n26931, n26932, n26933, n26934, n26935,
    n26936, n26937, n26938, n26939, n26940, n26941,
    n26942, n26943, n26944, n26945, n26946, n26947,
    n26948, n26949, n26950, n26951, n26952, n26953,
    n26954, n26955, n26956, n26957, n26958, n26959,
    n26960, n26961, n26962, n26963, n26964, n26965,
    n26966, n26967, n26968, n26969, n26970, n26971,
    n26972, n26973, n26974, n26975, n26976, n26977,
    n26978, n26979, n26980, n26981, n26982, n26983,
    n26984, n26985, n26986, n26987, n26988, n26989,
    n26990, n26991, n26992, n26993, n26994, n26995,
    n26996, n26997, n26998, n26999, n27000, n27001,
    n27002, n27003, n27004, n27005, n27006, n27007,
    n27008, n27009, n27010, n27011, n27012, n27013,
    n27014, n27015, n27016, n27017, n27018, n27019,
    n27020, n27021, n27022, n27023, n27024, n27025,
    n27026, n27027, n27028, n27029, n27030, n27031,
    n27032, n27033, n27034, n27035, n27036, n27037,
    n27038, n27039, n27040, n27041, n27042, n27043,
    n27044, n27045, n27046, n27047, n27048, n27049,
    n27050, n27051, n27052, n27053, n27054, n27055,
    n27056, n27057, n27058, n27059, n27060, n27061,
    n27062, n27063, n27064, n27065, n27066, n27067,
    n27068, n27069, n27070, n27071, n27072, n27073,
    n27074, n27075, n27076, n27077, n27078, n27079,
    n27080, n27081, n27082, n27083, n27084, n27085,
    n27086, n27087, n27088, n27089, n27090, n27091,
    n27092, n27093, n27094, n27095, n27096, n27097,
    n27098, n27099, n27100, n27101, n27102, n27103,
    n27104, n27105, n27106, n27107, n27108, n27109,
    n27110, n27111, n27112, n27113, n27114, n27115,
    n27116, n27117, n27118, n27119, n27120, n27121,
    n27122, n27123, n27124, n27125, n27126, n27127,
    n27128, n27129, n27130, n27131, n27132, n27133,
    n27134, n27135, n27136, n27137, n27138, n27139,
    n27140, n27141, n27142, n27143, n27144, n27145,
    n27146, n27147, n27148, n27149, n27150, n27151,
    n27152, n27153, n27154, n27155, n27156, n27157,
    n27158, n27159, n27160, n27161, n27162, n27163,
    n27164, n27165, n27166, n27167, n27168, n27169,
    n27170, n27171, n27172, n27173, n27174, n27175,
    n27176, n27177, n27178, n27179, n27180, n27181,
    n27182, n27183, n27184, n27185, n27186, n27187,
    n27188, n27189, n27190, n27191, n27192, n27193,
    n27194, n27195, n27196, n27197, n27198, n27199,
    n27200, n27201, n27202, n27203, n27204, n27205,
    n27206, n27207, n27208, n27209, n27210, n27211,
    n27212, n27213, n27214, n27215, n27216, n27217,
    n27218, n27219, n27220, n27221, n27222, n27223,
    n27224, n27225, n27226, n27227, n27228, n27229,
    n27230, n27231, n27232, n27233, n27234, n27235,
    n27236, n27237, n27238, n27239, n27240, n27241,
    n27242, n27243, n27244, n27245, n27246, n27247,
    n27248, n27249, n27250, n27251, n27252, n27253,
    n27254, n27255, n27256, n27257, n27258, n27259,
    n27260, n27261, n27262, n27263, n27264, n27265,
    n27266, n27267, n27268, n27269, n27270, n27271,
    n27272, n27273, n27274, n27275, n27276, n27277,
    n27278, n27279, n27280, n27281, n27282, n27283,
    n27284, n27285, n27286, n27287, n27288, n27289,
    n27290, n27291, n27292, n27293, n27294, n27295,
    n27296, n27297, n27298, n27299, n27300, n27301,
    n27302, n27303, n27304, n27305, n27306, n27307,
    n27308, n27309, n27310, n27311, n27312, n27313,
    n27314, n27315, n27316, n27317, n27318, n27319,
    n27320, n27321, n27322, n27323, n27324, n27325,
    n27326, n27327, n27328, n27329, n27330, n27331,
    n27332, n27333, n27334, n27335, n27336, n27337,
    n27338, n27339, n27340, n27341, n27342, n27343,
    n27344, n27345, n27346, n27347, n27348, n27349,
    n27350, n27351, n27352, n27353, n27354, n27355,
    n27356, n27357, n27358, n27359, n27360, n27361,
    n27362, n27363, n27364, n27365, n27366, n27367,
    n27368, n27369, n27370, n27371, n27372, n27373,
    n27374, n27375, n27376, n27377, n27378, n27379,
    n27380, n27381, n27382, n27383, n27384, n27385,
    n27386, n27387, n27388, n27389, n27390, n27391,
    n27392, n27393, n27394, n27395, n27396, n27397,
    n27398, n27399, n27400, n27401, n27402, n27403,
    n27404, n27405, n27406, n27407, n27408, n27409,
    n27410, n27411, n27412, n27413, n27414, n27415,
    n27416, n27417, n27418, n27419, n27420, n27421,
    n27422, n27423, n27424, n27425, n27426, n27427,
    n27428, n27429, n27430, n27431, n27432, n27433,
    n27434, n27435, n27436, n27437, n27438, n27439,
    n27440, n27441, n27442, n27443, n27444, n27445,
    n27446, n27447, n27448, n27449, n27450, n27451,
    n27452, n27453, n27454, n27455, n27456, n27457,
    n27458, n27459, n27460, n27461, n27462, n27463,
    n27464, n27465, n27466, n27467, n27468, n27469,
    n27470, n27471, n27472, n27473, n27474, n27475,
    n27476, n27477, n27478, n27479, n27480, n27481,
    n27482, n27483, n27484, n27485, n27486, n27487,
    n27488, n27489, n27490, n27491, n27492, n27493,
    n27494, n27495, n27496, n27497, n27498, n27499,
    n27500, n27501, n27502, n27503, n27504, n27505,
    n27506, n27507, n27508, n27509, n27510, n27511,
    n27512, n27513, n27514, n27515, n27516, n27517,
    n27518, n27519, n27520, n27521, n27522, n27523,
    n27524, n27525, n27526, n27527, n27528, n27529,
    n27530, n27531, n27532, n27533, n27534, n27535,
    n27536, n27537, n27538, n27539, n27540, n27541,
    n27542, n27543, n27544, n27545, n27546, n27547,
    n27548, n27549, n27550, n27551, n27552, n27553,
    n27554, n27555, n27556, n27557, n27558, n27559,
    n27560, n27561, n27562, n27563, n27564, n27565,
    n27566, n27567, n27568, n27569, n27570, n27571,
    n27572, n27573, n27574, n27575, n27576, n27577,
    n27578, n27579, n27580, n27581, n27582, n27583,
    n27584, n27585, n27586, n27587, n27588, n27589,
    n27590, n27591, n27592, n27593, n27594, n27595,
    n27596, n27597, n27598, n27599, n27600, n27601,
    n27602, n27603, n27604, n27605, n27606, n27607,
    n27608, n27609, n27610, n27611, n27612, n27613,
    n27614, n27615, n27616, n27617, n27618, n27619,
    n27620, n27621, n27622, n27623, n27624, n27625,
    n27626, n27627, n27628, n27629, n27630, n27631,
    n27632, n27633, n27634, n27635, n27636, n27637,
    n27638, n27639, n27640, n27641, n27642, n27643,
    n27644, n27645, n27646, n27647, n27648, n27649,
    n27650, n27651, n27652, n27653, n27654, n27655,
    n27656, n27657, n27658, n27659, n27660, n27661,
    n27662, n27663, n27664, n27665, n27666, n27667,
    n27668, n27669, n27670, n27671, n27672, n27673,
    n27674, n27675, n27676, n27677, n27678, n27679,
    n27680, n27681, n27682, n27683, n27684, n27685,
    n27686, n27687, n27688, n27689, n27690, n27691,
    n27692, n27693, n27694, n27695, n27696, n27697,
    n27698, n27699, n27700, n27701, n27702, n27703,
    n27704, n27705, n27706, n27707, n27708, n27709,
    n27710, n27711, n27712, n27713, n27714, n27715,
    n27716, n27717, n27718, n27719, n27720, n27721,
    n27722, n27723, n27724, n27725, n27726, n27727,
    n27728, n27729, n27730, n27731, n27732, n27733,
    n27734, n27735, n27736, n27737, n27738, n27739,
    n27740, n27741, n27742, n27743, n27744, n27745,
    n27746, n27747, n27748, n27749, n27750, n27751,
    n27752, n27753, n27754, n27755, n27756, n27757,
    n27758, n27759, n27760, n27761, n27762, n27763,
    n27764, n27765, n27766, n27767, n27768, n27769,
    n27770, n27771, n27772, n27773, n27774, n27775,
    n27776, n27777, n27778, n27779, n27780, n27781,
    n27782, n27783, n27784, n27785, n27786, n27787,
    n27788, n27789, n27790, n27791, n27792, n27793,
    n27794, n27795, n27796, n27797, n27798, n27799,
    n27800, n27801, n27802, n27803, n27804, n27805,
    n27806, n27807, n27808, n27809, n27810, n27811,
    n27812, n27813, n27814, n27815, n27816, n27817,
    n27818, n27819, n27820, n27821, n27822, n27823,
    n27824, n27825, n27826, n27827, n27828, n27829,
    n27830, n27831, n27832, n27833, n27834, n27835,
    n27836, n27837, n27838, n27839, n27840, n27841,
    n27842, n27843, n27844, n27845, n27846, n27847,
    n27848, n27849, n27850, n27851, n27852, n27853,
    n27854, n27855, n27856, n27857, n27858, n27859,
    n27860, n27861, n27862, n27863, n27864, n27865,
    n27866, n27867, n27868, n27869, n27870, n27871,
    n27872, n27873, n27874, n27875, n27876, n27877,
    n27878, n27879, n27880, n27881, n27882, n27883,
    n27884, n27885, n27886, n27887, n27888, n27889,
    n27890, n27891, n27892, n27893, n27894, n27895,
    n27896, n27897, n27898, n27899, n27900, n27901,
    n27902, n27903, n27904, n27905, n27906, n27907,
    n27908, n27909, n27910, n27911, n27912, n27913,
    n27914, n27915, n27916, n27917, n27918, n27919,
    n27920, n27921, n27922, n27923, n27924, n27925,
    n27926, n27927, n27928, n27929, n27930, n27931,
    n27932, n27933, n27934, n27935, n27936, n27937,
    n27938, n27939, n27940, n27941, n27942, n27943,
    n27944, n27945, n27946, n27947, n27948, n27949,
    n27950, n27951, n27952, n27953, n27954, n27955,
    n27956, n27957, n27958, n27959, n27960, n27961,
    n27962, n27963, n27964, n27965, n27966, n27967,
    n27968, n27969, n27970, n27971, n27972, n27973,
    n27974, n27975, n27976, n27977, n27978, n27979,
    n27980, n27981, n27982, n27983, n27984, n27985,
    n27986, n27987, n27988, n27989, n27990, n27991,
    n27992, n27993, n27994, n27995, n27996, n27997,
    n27998, n27999, n28000, n28001, n28002, n28003,
    n28004, n28005, n28006, n28007, n28008, n28009,
    n28010, n28011, n28012, n28013, n28014, n28015,
    n28016, n28017, n28018, n28019, n28020, n28021,
    n28022, n28023, n28024, n28025, n28026, n28027,
    n28028, n28029, n28030, n28031, n28032, n28033,
    n28034, n28035, n28036, n28037, n28038, n28039,
    n28040, n28041, n28042, n28043, n28044, n28045,
    n28046, n28047, n28048, n28049, n28050, n28051,
    n28052, n28053, n28054, n28055, n28056, n28057,
    n28058, n28059, n28060, n28061, n28062, n28063,
    n28064, n28065, n28066, n28067, n28068, n28069,
    n28070, n28071, n28072, n28073, n28074, n28075,
    n28076, n28077, n28078, n28079, n28080, n28081,
    n28082, n28083, n28084, n28085, n28086, n28087,
    n28088, n28089, n28090, n28091, n28092, n28093,
    n28094, n28095, n28096, n28097, n28098, n28099,
    n28100, n28101, n28102, n28103, n28104, n28105,
    n28106, n28107, n28108, n28109, n28110, n28111,
    n28112, n28113, n28114, n28115, n28116, n28117,
    n28118, n28119, n28120, n28121, n28122, n28123,
    n28124, n28125, n28126, n28127, n28128, n28129,
    n28130, n28131, n28132, n28133, n28134, n28135,
    n28136, n28137, n28138, n28139, n28140, n28141,
    n28142, n28143, n28144, n28145, n28146, n28147,
    n28148, n28149, n28150, n28151, n28152, n28153,
    n28154, n28155, n28156, n28157, n28158, n28159,
    n28160, n28161, n28162, n28163, n28164, n28165,
    n28166, n28167, n28168, n28169, n28170, n28171,
    n28172, n28173, n28174, n28175, n28176, n28177,
    n28178, n28179, n28180, n28181, n28182, n28183,
    n28184, n28185, n28186, n28187, n28188, n28189,
    n28190, n28191, n28192, n28193, n28194, n28195,
    n28196, n28197, n28198, n28199, n28200, n28201,
    n28202, n28203, n28204, n28205, n28206, n28207,
    n28208, n28209, n28210, n28211, n28212, n28213,
    n28214, n28215, n28216, n28217, n28218, n28219,
    n28220, n28221, n28222, n28223, n28224, n28225,
    n28226, n28227, n28228, n28229, n28230, n28231,
    n28232, n28233, n28234, n28235, n28236, n28237,
    n28238, n28239, n28240, n28241, n28242, n28243,
    n28244, n28245, n28246, n28247, n28248, n28249,
    n28250, n28251, n28252, n28253, n28254, n28255,
    n28256, n28257, n28258, n28259, n28260, n28261,
    n28262, n28263, n28264, n28265, n28266, n28267,
    n28268, n28269, n28270, n28271, n28272, n28273,
    n28274, n28275, n28276, n28277, n28278, n28279,
    n28280, n28282, n28283, n28284, n28285, n28286,
    n28287, n28288, n28289, n28290, n28291, n28292,
    n28293, n28294, n28295, n28296, n28297, n28298,
    n28299, n28300, n28301, n28302, n28303, n28304,
    n28305, n28306, n28307, n28308, n28309, n28310,
    n28311, n28312, n28313, n28314, n28315, n28316,
    n28317, n28318, n28319, n28320, n28321, n28322,
    n28323, n28324, n28325, n28326, n28327, n28328,
    n28329, n28330, n28331, n28332, n28333, n28334,
    n28335, n28336, n28337, n28338, n28339, n28340,
    n28341, n28342, n28343, n28344, n28345, n28346,
    n28347, n28348, n28349, n28350, n28351, n28352,
    n28353, n28354, n28355, n28356, n28357, n28358,
    n28359, n28360, n28361, n28362, n28363, n28364,
    n28365, n28366, n28367, n28368, n28369, n28370,
    n28371, n28372, n28373, n28374, n28375, n28376,
    n28377, n28378, n28379, n28380, n28381, n28382,
    n28383, n28384, n28385, n28386, n28387, n28388,
    n28389, n28390, n28391, n28392, n28393, n28394,
    n28395, n28396, n28397, n28398, n28399, n28400,
    n28401, n28402, n28403, n28404, n28405, n28406,
    n28407, n28408, n28409, n28410, n28411, n28412,
    n28413, n28414, n28415, n28416, n28417, n28418,
    n28419, n28420, n28421, n28422, n28423, n28424,
    n28425, n28426, n28427, n28428, n28429, n28430,
    n28431, n28432, n28433, n28434, n28435, n28436,
    n28437, n28438, n28439, n28440, n28441, n28442,
    n28443, n28444, n28445, n28446, n28447, n28448,
    n28449, n28450, n28451, n28452, n28453, n28454,
    n28455, n28456, n28457, n28458, n28459, n28460,
    n28461, n28462, n28463, n28464, n28465, n28466,
    n28467, n28468, n28469, n28470, n28471, n28472,
    n28473, n28474, n28475, n28476, n28477, n28478,
    n28479, n28480, n28481, n28482, n28483, n28484,
    n28485, n28486, n28487, n28488, n28489, n28490,
    n28491, n28492, n28493, n28494, n28495, n28496,
    n28497, n28498, n28499, n28500, n28501, n28502,
    n28503, n28504, n28505, n28506, n28507, n28508,
    n28509, n28510, n28511, n28512, n28513, n28514,
    n28515, n28516, n28517, n28518, n28519, n28520,
    n28521, n28522, n28523, n28524, n28525, n28526,
    n28527, n28528, n28529, n28530, n28531, n28532,
    n28533, n28534, n28535, n28536, n28537, n28538,
    n28539, n28540, n28541, n28542, n28543, n28544,
    n28545, n28546, n28547, n28548, n28549, n28550,
    n28551, n28552, n28553, n28554, n28555, n28556,
    n28557, n28558, n28559, n28560, n28561, n28562,
    n28563, n28564, n28565, n28566, n28567, n28568,
    n28569, n28570, n28571, n28572, n28573, n28574,
    n28575, n28576, n28577, n28578, n28579, n28580,
    n28581, n28582, n28583, n28584, n28585, n28586,
    n28587, n28588, n28589, n28590, n28591, n28592,
    n28593, n28594, n28595, n28596, n28597, n28598,
    n28600, n28601, n28603, n28604, n28605, n28606,
    n28607, n28608, n28609, n28610, n28611, n28612,
    n28613, n28614, n28615, n28616, n28617, n28618,
    n28619, n28620, n28621, n28622, n28623, n28624,
    n28625, n28626, n28627, n28628, n28629, n28630,
    n28631, n28632, n28633, n28634, n28635, n28636,
    n28637, n28638, n28639, n28640, n28641, n28642,
    n28643, n28644, n28645, n28646, n28647, n28648,
    n28649, n28650, n28651, n28652, n28653, n28654,
    n28655, n28656, n28657, n28658, n28659, n28660,
    n28661, n28662, n28663, n28664, n28665, n28666,
    n28667, n28668, n28669, n28670, n28671, n28672,
    n28673, n28674, n28675, n28676, n28677, n28678,
    n28679, n28680, n28681, n28682, n28683, n28684,
    n28685, n28686, n28687, n28688, n28689, n28690,
    n28691, n28692, n28693, n28694, n28695, n28696,
    n28697, n28698, n28699, n28700, n28701, n28702,
    n28703, n28704, n28705, n28706, n28707, n28708,
    n28709, n28710, n28711, n28712, n28713, n28714,
    n28715, n28716, n28717, n28718, n28719, n28720,
    n28721, n28722, n28723, n28724, n28725, n28726,
    n28727, n28728, n28729, n28730, n28731, n28732,
    n28733, n28734, n28735, n28736, n28737, n28738,
    n28739, n28740, n28741, n28742, n28743, n28744,
    n28745, n28746, n28747, n28748, n28749, n28750,
    n28751, n28752, n28753, n28754, n28755, n28756,
    n28757, n28758, n28759, n28760, n28761, n28762,
    n28763, n28764, n28765, n28766, n28767, n28768,
    n28769, n28770, n28771, n28772, n28773, n28774,
    n28775, n28776, n28777, n28778, n28779, n28780,
    n28781, n28782, n28783, n28784, n28785, n28786,
    n28787, n28788, n28789, n28790, n28791, n28792,
    n28793, n28794, n28795, n28796, n28797, n28798,
    n28799, n28800, n28801, n28802, n28803, n28804,
    n28805, n28806, n28807, n28808, n28809, n28810,
    n28811, n28812, n28813, n28814, n28815, n28816,
    n28817, n28818, n28819, n28820, n28821, n28822,
    n28823, n28824, n28825, n28826, n28827, n28828,
    n28829, n28830, n28831, n28832, n28833, n28834,
    n28835, n28836, n28837, n28838, n28839, n28840,
    n28841, n28842, n28843, n28844, n28845, n28846,
    n28847, n28848, n28849, n28850, n28851, n28852,
    n28853, n28854, n28855, n28856, n28857, n28858,
    n28859, n28860, n28861, n28862, n28863, n28864,
    n28865, n28866, n28867, n28868, n28869, n28870,
    n28871, n28872, n28873, n28874, n28875, n28876,
    n28877, n28878, n28879, n28880, n28881, n28882,
    n28883, n28884, n28885, n28886, n28887, n28888,
    n28889, n28890, n28891, n28892, n28893, n28894,
    n28895, n28896, n28897, n28898, n28899, n28900,
    n28901, n28902, n28903, n28904, n28905, n28906,
    n28907, n28908, n28909, n28910, n28911, n28912,
    n28913, n28914, n28915, n28916, n28917, n28918,
    n28919, n28920, n28921, n28922, n28923, n28924,
    n28925, n28926, n28927, n28928, n28929, n28930,
    n28931, n28932, n28933, n28934, n28935, n28936,
    n28937, n28938, n28939, n28940, n28941, n28942,
    n28943, n28944, n28945, n28946, n28947, n28948,
    n28949, n28950, n28951, n28952, n28953, n28954,
    n28955, n28956, n28957, n28958, n28959, n28960,
    n28961, n28962, n28963, n28964, n28965, n28966,
    n28967, n28968, n28969, n28970, n28971, n28972,
    n28973, n28974, n28975, n28976, n28977, n28978,
    n28979, n28980, n28981, n28982, n28983, n28984,
    n28985, n28986, n28987, n28988, n28989, n28990,
    n28991, n28992, n28993, n28994, n28995, n28996,
    n28997, n28998, n28999, n29000, n29001, n29002,
    n29003, n29004, n29005, n29006, n29007, n29008,
    n29009, n29010, n29011, n29012, n29013, n29014,
    n29015, n29016, n29017, n29018, n29019, n29020,
    n29021, n29022, n29023, n29024, n29025, n29026,
    n29027, n29028, n29029, n29030, n29031, n29032,
    n29033, n29034, n29035, n29036, n29037, n29038,
    n29039, n29040, n29041, n29042, n29043, n29044,
    n29045, n29046, n29047, n29048, n29049, n29050,
    n29051, n29052, n29053, n29054, n29055, n29056,
    n29057, n29058, n29059, n29060, n29061, n29062,
    n29063, n29064, n29065, n29066, n29067, n29068,
    n29069, n29070, n29071, n29072, n29073, n29074,
    n29075, n29076, n29077, n29078, n29079, n29080,
    n29081, n29082, n29083, n29084, n29085, n29086,
    n29087, n29088, n29089, n29090, n29091, n29092,
    n29093, n29094, n29095, n29096, n29097, n29098,
    n29099, n29100, n29101, n29102, n29103, n29104,
    n29105, n29106, n29107, n29108, n29109, n29110,
    n29111, n29112, n29113, n29114, n29115, n29116,
    n29117, n29118, n29119, n29120, n29121, n29122,
    n29123, n29124, n29125, n29126, n29127, n29128,
    n29129, n29130, n29131, n29132, n29133, n29134,
    n29135, n29136, n29137, n29138, n29139, n29140,
    n29141, n29142, n29143, n29144, n29145, n29146,
    n29147, n29148, n29149, n29150, n29151, n29152,
    n29153, n29154, n29155, n29156, n29157, n29158,
    n29159, n29160, n29161, n29162, n29163, n29164,
    n29165, n29166, n29167, n29168, n29169, n29170,
    n29171, n29172, n29173, n29174, n29175, n29176,
    n29177, n29178, n29179, n29180, n29181, n29182,
    n29183, n29184, n29185, n29186, n29187, n29188,
    n29189, n29190, n29191, n29192, n29193, n29194,
    n29195, n29196, n29197, n29198, n29199, n29200,
    n29201, n29202, n29203, n29204, n29205, n29206,
    n29207, n29208, n29209, n29210, n29211, n29212,
    n29213, n29214, n29215, n29216, n29217, n29218,
    n29219, n29220, n29221, n29222, n29223, n29224,
    n29225, n29226, n29227, n29228, n29229, n29230,
    n29231, n29232, n29233, n29234, n29235, n29236,
    n29237, n29238, n29239, n29240, n29241, n29242,
    n29243, n29244, n29245, n29246, n29247, n29248,
    n29249, n29250, n29251, n29252, n29253, n29254,
    n29255, n29256, n29257, n29258, n29259, n29260,
    n29261, n29262, n29263, n29264, n29265, n29266,
    n29267, n29268, n29269, n29270, n29271, n29272,
    n29273, n29274, n29275, n29276, n29277, n29278,
    n29279, n29280, n29281, n29282, n29283, n29284,
    n29285, n29286, n29287, n29288, n29289, n29290,
    n29291, n29292, n29293, n29294, n29295, n29296,
    n29297, n29298, n29299, n29300, n29301, n29302,
    n29303, n29304, n29305, n29306, n29307, n29308,
    n29309, n29310, n29311, n29312, n29313, n29314,
    n29315, n29316, n29317, n29318, n29319, n29320,
    n29321, n29322, n29323, n29324, n29325, n29326,
    n29327, n29328, n29329, n29330, n29331, n29332,
    n29333, n29334, n29335, n29336, n29337, n29338,
    n29339, n29340, n29341, n29342, n29343, n29344,
    n29345, n29346, n29347, n29348, n29349, n29350,
    n29351, n29352, n29353, n29354, n29355, n29356,
    n29357, n29358, n29359, n29360, n29361, n29362,
    n29363, n29364, n29365, n29366, n29367, n29368,
    n29369, n29370, n29371, n29372, n29373, n29374,
    n29375, n29376, n29377, n29378, n29379, n29380,
    n29381, n29382, n29383, n29384, n29385, n29386,
    n29387, n29388, n29389, n29390, n29391, n29392,
    n29393, n29394, n29395, n29396, n29397, n29398,
    n29399, n29400, n29401, n29402, n29403, n29404,
    n29405, n29406, n29407, n29408, n29409, n29410,
    n29411, n29412, n29413, n29414, n29415, n29416,
    n29417, n29418, n29419, n29420, n29421, n29422,
    n29423, n29424, n29425, n29426, n29427, n29428,
    n29429, n29430, n29431, n29432, n29433, n29434,
    n29435, n29436, n29437, n29438, n29439, n29440,
    n29441, n29442, n29443, n29444, n29445, n29446,
    n29447, n29448, n29449, n29450, n29451, n29452,
    n29453, n29454, n29455, n29456, n29457, n29458,
    n29459, n29460, n29461, n29462, n29463, n29464,
    n29465, n29466, n29467, n29468, n29469, n29470,
    n29471, n29472, n29473, n29474, n29475, n29476,
    n29477, n29478, n29479, n29480, n29481, n29482,
    n29483, n29484, n29485, n29486, n29487, n29488,
    n29489, n29490, n29491, n29492, n29493, n29494,
    n29495, n29496, n29497, n29498, n29499, n29500,
    n29501, n29502, n29503, n29504, n29505, n29506,
    n29507, n29508, n29509, n29510, n29511, n29512,
    n29513, n29514, n29515, n29516, n29517, n29518,
    n29519, n29520, n29521, n29522, n29523, n29524,
    n29525, n29526, n29527, n29528, n29529, n29530,
    n29531, n29532, n29533, n29534, n29535, n29536,
    n29537, n29538, n29539, n29540, n29541, n29542,
    n29543, n29544, n29545, n29546, n29547, n29548,
    n29549, n29550, n29551, n29552, n29553, n29554,
    n29555, n29556, n29557, n29558, n29559, n29560,
    n29561, n29562, n29563, n29564, n29565, n29566,
    n29567, n29568, n29569, n29570, n29571, n29572,
    n29573, n29574, n29575, n29576, n29577, n29578,
    n29579, n29580, n29581, n29582, n29583, n29584,
    n29585, n29586, n29587, n29588, n29589, n29590,
    n29591, n29592, n29593, n29594, n29595, n29596,
    n29597, n29598, n29599, n29600, n29601, n29602,
    n29603, n29604, n29605, n29606, n29607, n29608,
    n29609, n29610, n29611, n29612, n29613, n29614,
    n29615, n29616, n29617, n29618, n29619, n29620,
    n29621, n29622, n29623, n29624, n29625, n29626,
    n29627, n29628, n29629, n29630, n29631, n29632,
    n29633, n29634, n29635, n29636, n29637, n29638,
    n29639, n29640, n29641, n29642, n29643, n29644,
    n29645, n29646, n29647, n29648, n29649, n29650,
    n29651, n29652, n29653, n29654, n29655, n29656,
    n29657, n29658, n29659, n29660, n29661, n29662,
    n29663, n29664, n29665, n29666, n29667, n29668,
    n29669, n29670, n29671, n29672, n29673, n29674,
    n29675, n29676, n29677, n29678, n29679, n29680,
    n29681, n29682, n29683, n29684, n29685, n29686,
    n29687, n29688, n29689, n29690, n29691, n29692,
    n29693, n29694, n29695, n29696, n29697, n29698,
    n29699, n29700, n29701, n29702, n29703, n29704,
    n29705, n29706, n29707, n29708, n29709, n29710,
    n29711, n29712, n29713, n29714, n29715, n29716,
    n29717, n29718, n29719, n29720, n29721, n29722,
    n29723, n29724, n29725, n29726, n29727, n29728,
    n29729, n29730, n29731, n29732, n29733, n29734,
    n29735, n29736, n29737, n29738, n29739, n29740,
    n29741, n29742, n29743, n29744, n29745, n29746,
    n29747, n29748, n29749, n29750, n29751, n29752,
    n29753, n29754, n29755, n29756, n29757, n29758,
    n29759, n29760, n29761, n29762, n29763, n29764,
    n29765, n29766, n29767, n29768, n29769, n29770,
    n29771, n29772, n29773, n29774, n29775, n29776,
    n29777, n29778, n29779, n29780, n29781, n29782,
    n29783, n29784, n29785, n29786, n29787, n29788,
    n29789, n29790, n29791, n29792, n29793, n29794,
    n29795, n29796, n29797, n29798, n29799, n29800,
    n29801, n29802, n29803, n29804, n29805, n29806,
    n29807, n29808, n29809, n29810, n29811, n29812,
    n29813, n29814, n29815, n29816, n29817, n29818,
    n29819, n29820, n29821, n29822, n29823, n29824,
    n29825, n29826, n29827, n29828, n29829, n29830,
    n29831, n29832, n29833, n29834, n29835, n29836,
    n29837, n29838, n29839, n29840, n29841, n29842,
    n29843, n29844, n29845, n29846, n29847, n29848,
    n29849, n29850, n29851, n29852, n29853, n29854,
    n29855, n29856, n29857, n29858, n29859, n29860,
    n29861, n29862, n29863, n29864, n29865, n29866,
    n29867, n29868, n29869, n29870, n29871, n29872,
    n29873, n29874, n29875, n29876, n29877, n29878,
    n29879, n29880, n29881, n29882, n29883, n29884,
    n29885, n29886, n29887, n29888, n29889, n29890,
    n29891, n29892, n29893, n29894, n29895, n29896,
    n29897, n29898, n29899, n29900, n29901, n29902,
    n29903, n29904, n29905, n29906, n29907, n29908,
    n29909, n29910, n29911, n29912, n29913, n29914,
    n29915, n29916, n29917, n29918, n29919, n29920,
    n29921, n29922, n29923, n29924, n29925, n29926,
    n29927, n29928, n29929, n29930, n29931, n29932,
    n29933, n29934, n29935, n29936, n29937, n29938,
    n29939, n29940, n29941, n29942, n29944, n29945,
    n29946, n29947, n29948, n29949, n29950, n29951,
    n29952, n29953, n29954, n29955, n29956, n29957,
    n29958, n29959, n29960, n29961, n29962, n29963,
    n29964, n29965, n29966, n29967, n29968, n29969,
    n29970, n29971, n29972, n29973, n29974, n29975,
    n29976, n29977, n29978, n29979, n29980, n29981,
    n29982, n29983, n29984, n29985, n29986, n29987,
    n29988, n29989, n29990, n29991, n29992, n29993,
    n29994, n29995, n29996, n29997, n29998, n29999,
    n30000, n30001, n30002, n30003, n30004, n30005,
    n30006, n30007, n30008, n30009, n30010, n30011,
    n30012, n30013, n30014, n30015, n30016, n30017,
    n30018, n30019, n30020, n30021, n30022, n30023,
    n30024, n30025, n30026, n30027, n30028, n30029,
    n30030, n30031, n30032, n30033, n30034, n30035,
    n30036, n30037, n30038, n30039, n30040, n30041,
    n30042, n30043, n30044, n30045, n30046, n30047,
    n30048, n30049, n30050, n30051, n30052, n30053,
    n30054, n30055, n30056, n30057, n30058, n30059,
    n30060, n30061, n30062, n30063, n30064, n30065,
    n30066, n30067, n30068, n30069, n30070, n30071,
    n30072, n30073, n30074, n30075, n30076, n30077,
    n30078, n30079, n30080, n30081, n30082, n30083,
    n30084, n30085, n30086, n30087, n30088, n30089,
    n30090, n30091, n30092, n30093, n30094, n30095,
    n30096, n30097, n30098, n30099, n30100, n30101,
    n30102, n30103, n30104, n30105, n30106, n30107,
    n30108, n30109, n30110, n30111, n30112, n30113,
    n30114, n30115, n30116, n30117, n30118, n30119,
    n30120, n30121, n30122, n30123, n30124, n30125,
    n30126, n30127, n30128, n30129, n30130, n30131,
    n30132, n30133, n30134, n30135, n30136, n30137,
    n30138, n30139, n30140, n30141, n30142, n30143,
    n30144, n30145, n30146, n30147, n30148, n30149,
    n30150, n30151, n30152, n30153, n30154, n30155,
    n30156, n30157, n30158, n30159, n30160, n30161,
    n30162, n30163, n30164, n30165, n30166, n30167,
    n30168, n30169, n30170, n30171, n30172, n30173,
    n30174, n30175, n30176, n30177, n30178, n30179,
    n30180, n30181, n30182, n30183, n30184, n30185,
    n30186, n30187, n30188, n30189, n30190, n30191,
    n30192, n30193, n30194, n30195, n30196, n30197,
    n30198, n30199, n30200, n30201, n30202, n30203,
    n30204, n30205, n30206, n30207, n30208, n30209,
    n30210, n30211, n30212, n30213, n30214, n30215,
    n30216, n30217, n30218, n30219, n30220, n30221,
    n30222, n30223, n30224, n30225, n30226, n30227,
    n30228, n30229, n30230, n30231, n30232, n30233,
    n30234, n30235, n30236, n30237, n30238, n30239,
    n30240, n30241, n30242, n30243, n30244, n30245,
    n30246, n30247, n30248, n30249, n30250, n30251,
    n30252, n30253, n30254, n30255, n30256, n30257,
    n30258, n30259, n30260, n30261, n30262, n30263,
    n30264, n30265, n30266, n30267, n30268, n30269,
    n30270, n30271, n30272, n30273, n30274, n30275,
    n30276, n30277, n30278, n30279, n30280, n30281,
    n30282, n30283, n30284, n30285, n30286, n30287,
    n30288, n30289, n30290, n30291, n30292, n30293,
    n30294, n30295, n30296, n30297, n30298, n30299,
    n30300, n30301, n30302, n30303, n30304, n30305,
    n30306, n30307, n30308, n30309, n30310, n30311,
    n30312, n30313, n30314, n30315, n30316, n30317,
    n30318, n30319, n30320, n30321, n30322, n30323,
    n30324, n30325, n30326, n30327, n30328, n30329,
    n30330, n30331, n30332, n30333, n30334, n30335,
    n30336, n30337, n30338, n30339, n30340, n30341,
    n30342, n30343, n30344, n30345, n30346, n30347,
    n30348, n30349, n30350, n30351, n30352, n30353,
    n30354, n30355, n30356, n30357, n30358, n30359,
    n30360, n30361, n30362, n30363, n30364, n30365,
    n30366, n30367, n30368, n30369, n30370, n30371,
    n30372, n30373, n30374, n30375, n30376, n30377,
    n30378, n30379, n30380, n30381, n30382, n30383,
    n30384, n30385, n30386, n30387, n30388, n30389,
    n30390, n30391, n30392, n30393, n30394, n30395,
    n30396, n30397, n30398, n30399, n30400, n30401,
    n30402, n30403, n30404, n30405, n30406, n30407,
    n30408, n30409, n30410, n30411, n30412, n30413,
    n30414, n30415, n30416, n30417, n30418, n30419,
    n30420, n30421, n30422, n30423, n30424, n30425,
    n30426, n30427, n30428, n30429, n30430, n30431,
    n30432, n30433, n30434, n30435, n30436, n30437,
    n30438, n30439, n30440, n30441, n30442, n30443,
    n30444, n30445, n30446, n30447, n30448, n30449,
    n30450, n30451, n30452, n30453, n30454, n30455,
    n30456, n30457, n30458, n30459, n30460, n30461,
    n30462, n30463, n30464, n30465, n30466, n30467,
    n30468, n30469, n30470, n30471, n30472, n30473,
    n30474, n30475, n30476, n30477, n30478, n30479,
    n30480, n30481, n30482, n30483, n30484, n30485,
    n30486, n30487, n30488, n30489, n30490, n30491,
    n30492, n30493, n30494, n30495, n30496, n30497,
    n30498, n30499, n30500, n30501, n30502, n30503,
    n30504, n30505, n30506, n30507, n30508, n30509,
    n30510, n30511, n30512, n30513, n30514, n30515,
    n30516, n30517, n30518, n30519, n30520, n30521,
    n30522, n30523, n30524, n30525, n30526, n30527,
    n30528, n30529, n30530, n30531, n30532, n30533,
    n30534, n30535, n30536, n30537, n30538, n30539,
    n30540, n30541, n30542, n30543, n30544, n30545,
    n30546, n30547, n30548, n30549, n30550, n30551,
    n30552, n30553, n30554, n30555, n30556, n30557,
    n30558, n30559, n30560, n30561, n30562, n30563,
    n30564, n30565, n30566, n30567, n30568, n30569,
    n30570, n30571, n30572, n30573, n30574, n30575,
    n30576, n30577, n30578, n30579, n30580, n30581,
    n30582, n30583, n30584, n30585, n30586, n30587,
    n30588, n30589, n30590, n30591, n30592, n30593,
    n30594, n30595, n30596, n30597, n30598, n30599,
    n30600, n30601, n30602, n30603, n30604, n30605,
    n30606, n30607, n30608, n30609, n30610, n30611,
    n30612, n30613, n30614, n30615, n30616, n30617,
    n30618, n30619, n30620, n30621, n30622, n30623,
    n30624, n30625, n30626, n30627, n30628, n30629,
    n30630, n30631, n30632, n30633, n30634, n30635,
    n30636, n30637, n30638, n30639, n30640, n30641,
    n30642, n30643, n30644, n30645, n30646, n30647,
    n30648, n30649, n30650, n30651, n30652, n30653,
    n30654, n30655, n30656, n30657, n30658, n30659,
    n30660, n30661, n30662, n30663, n30664, n30665,
    n30666, n30667, n30668, n30669, n30670, n30671,
    n30672, n30673, n30674, n30675, n30676, n30677,
    n30678, n30679, n30680, n30681, n30682, n30683,
    n30684, n30685, n30686, n30687, n30688, n30689,
    n30690, n30691, n30692, n30693, n30694, n30695,
    n30696, n30697, n30698, n30699, n30700, n30701,
    n30702, n30703, n30704, n30705, n30706, n30707,
    n30708, n30709, n30710, n30711, n30712, n30713,
    n30714, n30715, n30716, n30717, n30718, n30719,
    n30720, n30721, n30722, n30723, n30724, n30725,
    n30726, n30727, n30728, n30729, n30730, n30731,
    n30732, n30733, n30734, n30735, n30736, n30737,
    n30738, n30739, n30740, n30741, n30742, n30743,
    n30744, n30745, n30746, n30747, n30748, n30749,
    n30750, n30751, n30752, n30753, n30754, n30755,
    n30756, n30757, n30758, n30759, n30760, n30761,
    n30762, n30763, n30764, n30765, n30766, n30767,
    n30768, n30769, n30770, n30771, n30772, n30773,
    n30774, n30775, n30776, n30777, n30778, n30779,
    n30780, n30781, n30782, n30783, n30784, n30785,
    n30786, n30787, n30788, n30789, n30790, n30791,
    n30792, n30793, n30794, n30795, n30796, n30797,
    n30798, n30799, n30800, n30801, n30802, n30803,
    n30804, n30805, n30806, n30807, n30808, n30809,
    n30810, n30811, n30812, n30813, n30814, n30815,
    n30816, n30817, n30818, n30819, n30820, n30821,
    n30822, n30823, n30824, n30825, n30826, n30827,
    n30828, n30829, n30830, n30831, n30832, n30833,
    n30834, n30835, n30836, n30837, n30838, n30839,
    n30840, n30841, n30842, n30843, n30844, n30845,
    n30846, n30847, n30848, n30849, n30850, n30851,
    n30852, n30853, n30854, n30855, n30856, n30857,
    n30858, n30859, n30860, n30861, n30862, n30863,
    n30864, n30865, n30866, n30867, n30868, n30869,
    n30870, n30871, n30872, n30873, n30874, n30875,
    n30876, n30877, n30878, n30879, n30880, n30881,
    n30882, n30883, n30884, n30885, n30886, n30887,
    n30888, n30889, n30890, n30891, n30892, n30893,
    n30894, n30895, n30896, n30897, n30898, n30899,
    n30900, n30901, n30902, n30903, n30904, n30905,
    n30906, n30907, n30908, n30909, n30910, n30911,
    n30912, n30913, n30914, n30915, n30916, n30917,
    n30918, n30919, n30920, n30921, n30922, n30923,
    n30924, n30925, n30926, n30927, n30928, n30929,
    n30930, n30931, n30932, n30933, n30934, n30935,
    n30936, n30937, n30938, n30939, n30940, n30941,
    n30942, n30943, n30944, n30945, n30946, n30947,
    n30948, n30949, n30950, n30951, n30952, n30953,
    n30954, n30955, n30956, n30957, n30958, n30959,
    n30960, n30961, n30962, n30963, n30964, n30965,
    n30966, n30967, n30968, n30969, n30970, n30971,
    n30972, n30973, n30974, n30975, n30976, n30977,
    n30978, n30979, n30980, n30981, n30982, n30983,
    n30984, n30985, n30986, n30987, n30988, n30989,
    n30990, n30991, n30992, n30993, n30994, n30995,
    n30996, n30997, n30998, n30999, n31000, n31001,
    n31002, n31003, n31004, n31005, n31006, n31007,
    n31008, n31009, n31010, n31011, n31012, n31013,
    n31014, n31015, n31016, n31017, n31018, n31019,
    n31020, n31021, n31022, n31023, n31024, n31025,
    n31026, n31027, n31028, n31029, n31030, n31031,
    n31032, n31033, n31034, n31035, n31036, n31037,
    n31038, n31039, n31040, n31041, n31042, n31043,
    n31044, n31045, n31046, n31047, n31048, n31049,
    n31050, n31051, n31052, n31053, n31054, n31055,
    n31056, n31057, n31058, n31059, n31060, n31061,
    n31062, n31063, n31064, n31065, n31066, n31067,
    n31068, n31069, n31070, n31071, n31072, n31073,
    n31074, n31075, n31076, n31077, n31078, n31079,
    n31080, n31081, n31082, n31083, n31084, n31085,
    n31086, n31087, n31088, n31089, n31090, n31091,
    n31092, n31093, n31094, n31095, n31096, n31097,
    n31098, n31099, n31100, n31101, n31102, n31103,
    n31104, n31105, n31106, n31107, n31108, n31109,
    n31110, n31111, n31112, n31113, n31114, n31115,
    n31116, n31117, n31118, n31119, n31120, n31121,
    n31122, n31123, n31124, n31125, n31126, n31127,
    n31128, n31129, n31130, n31131, n31132, n31133,
    n31134, n31135, n31136, n31137, n31138, n31139,
    n31140, n31141, n31142, n31143, n31144, n31145,
    n31146, n31147, n31148, n31149, n31150, n31151,
    n31152, n31153, n31154, n31155, n31156, n31157,
    n31158, n31159, n31160, n31161, n31162, n31163,
    n31164, n31165, n31166, n31167, n31168, n31169,
    n31170, n31171, n31172, n31173, n31174, n31175,
    n31176, n31177, n31178, n31179, n31180, n31181,
    n31182, n31183, n31184, n31185, n31186, n31187,
    n31188, n31189, n31190, n31191, n31192, n31193,
    n31194, n31195, n31196, n31197, n31198, n31199,
    n31200, n31201, n31202, n31203, n31204, n31205,
    n31206, n31207, n31208, n31209, n31210, n31211,
    n31212, n31213, n31214, n31215, n31216, n31217,
    n31218, n31219, n31220, n31221, n31222, n31223,
    n31224, n31225, n31226, n31227, n31228, n31229,
    n31230, n31231, n31232, n31233, n31234, n31235,
    n31236, n31237, n31238, n31239, n31240, n31241,
    n31242, n31243, n31244, n31245, n31246, n31247,
    n31248, n31249, n31250, n31251, n31252, n31253,
    n31254, n31255, n31256, n31257, n31258, n31259,
    n31260, n31261, n31262, n31263, n31264, n31265,
    n31266, n31267, n31268, n31269, n31270, n31271,
    n31272, n31273, n31274, n31275, n31276, n31277,
    n31278, n31279, n31280, n31281, n31282, n31283,
    n31284, n31285, n31286, n31287, n31288, n31289,
    n31290, n31291, n31292, n31293, n31294, n31295,
    n31296, n31297, n31298, n31299, n31300, n31301,
    n31302, n31303, n31304, n31305, n31306, n31307,
    n31308, n31309, n31310, n31311, n31312, n31313,
    n31314, n31315, n31316, n31317, n31318, n31319,
    n31320, n31321, n31322, n31323, n31324, n31325,
    n31326, n31327, n31328, n31329, n31330, n31331,
    n31332, n31333, n31334, n31335, n31336, n31337,
    n31338, n31339, n31340, n31341, n31342, n31343,
    n31344, n31345, n31346, n31347, n31348, n31349,
    n31350, n31351, n31352, n31353, n31354, n31355,
    n31356, n31357, n31358, n31359, n31360, n31361,
    n31362, n31363, n31364, n31365, n31366, n31367,
    n31368, n31369, n31370, n31371, n31372, n31373,
    n31374, n31375, n31376, n31377, n31378, n31379,
    n31380, n31381, n31382, n31383, n31384, n31385,
    n31386, n31387, n31389, n31390, n31391, n31392,
    n31393, n31394, n31395, n31396, n31397, n31398,
    n31399, n31400, n31401, n31402, n31403, n31404,
    n31405, n31406, n31407, n31408, n31409, n31410,
    n31411, n31412, n31413, n31414, n31415, n31416,
    n31417, n31418, n31419, n31420, n31421, n31422,
    n31423, n31424, n31425, n31426, n31427, n31428,
    n31429, n31430, n31431, n31432, n31433, n31434,
    n31435, n31436, n31437, n31438, n31439, n31440,
    n31441, n31442, n31443, n31444, n31445, n31446,
    n31447, n31448, n31449, n31450, n31451, n31452,
    n31453, n31454, n31455, n31456, n31457, n31458,
    n31459, n31460, n31461, n31462, n31463, n31464,
    n31465, n31466, n31467, n31468, n31469, n31470,
    n31471, n31472, n31473, n31474, n31475, n31476,
    n31477, n31478, n31479, n31480, n31481, n31482,
    n31483, n31484, n31485, n31486, n31487, n31488,
    n31489, n31490, n31491, n31492, n31493, n31494,
    n31495, n31496, n31497, n31498, n31499, n31500,
    n31501, n31502, n31503, n31504, n31505, n31506,
    n31507, n31508, n31509, n31510, n31511, n31512,
    n31513, n31514, n31515, n31516, n31517, n31518,
    n31519, n31520, n31521, n31522, n31523, n31524,
    n31525, n31526, n31527, n31528, n31529, n31530,
    n31531, n31532, n31533, n31534, n31535, n31536,
    n31537, n31538, n31539, n31540, n31541, n31542,
    n31543, n31544, n31545, n31546, n31547, n31548,
    n31549, n31550, n31551, n31552, n31553, n31554,
    n31555, n31556, n31557, n31558, n31559, n31560,
    n31561, n31562, n31563, n31564, n31565, n31566,
    n31567, n31568, n31569, n31570, n31571, n31572,
    n31573, n31574, n31575, n31576, n31577, n31578,
    n31580, n31581, n31582, n31583, n31584, n31585,
    n31586, n31587, n31588, n31589, n31590, n31591,
    n31592, n31593, n31594, n31595, n31596, n31597,
    n31598, n31599, n31600, n31601, n31602, n31603,
    n31604, n31605, n31606, n31607, n31608, n31609,
    n31610, n31611, n31612, n31613, n31614, n31615,
    n31616, n31617, n31618, n31619, n31620, n31621,
    n31622, n31623, n31624, n31625, n31626, n31627,
    n31628, n31629, n31630, n31631, n31632, n31633,
    n31634, n31635, n31636, n31637, n31638, n31639,
    n31640, n31641, n31642, n31643, n31644, n31645,
    n31646, n31647, n31648, n31649, n31650, n31651,
    n31652, n31653, n31654, n31655, n31656, n31657,
    n31658, n31659, n31660, n31661, n31662, n31663,
    n31664, n31665, n31666, n31667, n31668, n31669,
    n31670, n31671, n31672, n31673, n31674, n31675,
    n31676, n31677, n31678, n31679, n31680, n31681,
    n31682, n31683, n31684, n31685, n31686, n31687,
    n31688, n31689, n31690, n31691, n31692, n31693,
    n31694, n31695, n31696, n31697, n31698, n31699,
    n31700, n31701, n31702, n31703, n31704, n31705,
    n31706, n31707, n31708, n31709, n31710, n31711,
    n31712, n31713, n31714, n31715, n31716, n31717,
    n31718, n31719, n31720, n31721, n31722, n31723,
    n31724, n31725, n31726, n31727, n31728, n31729,
    n31730, n31731, n31732, n31733, n31735, n31736,
    n31737, n31738, n31739, n31740, n31741, n31742,
    n31743, n31744, n31745, n31746, n31747, n31748,
    n31749, n31750, n31751, n31752, n31753, n31754,
    n31755, n31756, n31757, n31758, n31759, n31760,
    n31761, n31762, n31763, n31764, n31765, n31766,
    n31767, n31768, n31769, n31770, n31771, n31772,
    n31773, n31774, n31775, n31776, n31777, n31778,
    n31779, n31780, n31781, n31782, n31783, n31784,
    n31785, n31786, n31787, n31788, n31789, n31790,
    n31791, n31792, n31793, n31794, n31795, n31796,
    n31797, n31798, n31799, n31800, n31801, n31802,
    n31803, n31804, n31805, n31806, n31807, n31808,
    n31809, n31810, n31811, n31812, n31813, n31814,
    n31815, n31816, n31817, n31818, n31819, n31820,
    n31821, n31822, n31823, n31824, n31825, n31826,
    n31827, n31828, n31829, n31830, n31831, n31832,
    n31833, n31834, n31835, n31836, n31837, n31838,
    n31839, n31840, n31841, n31842, n31843, n31844,
    n31845, n31846, n31847, n31848, n31849, n31850,
    n31851, n31852, n31853, n31854, n31855, n31856,
    n31857, n31858, n31859, n31860, n31861, n31862,
    n31864, n31865, n31866, n31867, n31868, n31869,
    n31870, n31871, n31872, n31873, n31874, n31875,
    n31876, n31877, n31878, n31879, n31880, n31881,
    n31882, n31883, n31884, n31885, n31886, n31887,
    n31888, n31889, n31890, n31891, n31892, n31893,
    n31894, n31895, n31896, n31897, n31898, n31899,
    n31900, n31901, n31902, n31903, n31904, n31905,
    n31906, n31907, n31908, n31909, n31910, n31911,
    n31912, n31913, n31914, n31915, n31916, n31917,
    n31918, n31919, n31920, n31921, n31922, n31923,
    n31924, n31925, n31926, n31927, n31928, n31929,
    n31930, n31931, n31932, n31933, n31934, n31935,
    n31936, n31937, n31938, n31939, n31940, n31941,
    n31942, n31943, n31944, n31945, n31946, n31947,
    n31948, n31949, n31950, n31951, n31952, n31953,
    n31954, n31955, n31956, n31957, n31958, n31959,
    n31960, n31961, n31962, n31963, n31964, n31965,
    n31966, n31967, n31968, n31969, n31970, n31971,
    n31972, n31973, n31974, n31975, n31976, n31977,
    n31978, n31979, n31980, n31981, n31982, n31983,
    n31984, n31985, n31986, n31987, n31988, n31989,
    n31991, n31992, n31993, n31994, n31995, n31996,
    n31997, n31998, n31999, n32000, n32001, n32002,
    n32003, n32004, n32005, n32006, n32007, n32008,
    n32009, n32010, n32011, n32012, n32013, n32014,
    n32015, n32016, n32017, n32018, n32019, n32020,
    n32021, n32022, n32023, n32024, n32025, n32026,
    n32027, n32028, n32029, n32030, n32031, n32032,
    n32033, n32034, n32035, n32036, n32037, n32038,
    n32039, n32040, n32041, n32042, n32043, n32044,
    n32045, n32046, n32047, n32048, n32049, n32050,
    n32051, n32052, n32053, n32054, n32055, n32056,
    n32057, n32058, n32059, n32060, n32061, n32062,
    n32063, n32064, n32065, n32066, n32067, n32068,
    n32069, n32070, n32071, n32072, n32073, n32074,
    n32075, n32076, n32077, n32078, n32079, n32080,
    n32081, n32082, n32083, n32084, n32085, n32087,
    n32088, n32089, n32090, n32091, n32092, n32093,
    n32094, n32095, n32096, n32097, n32098, n32099,
    n32100, n32101, n32102, n32103, n32104, n32105,
    n32106, n32107, n32108, n32109, n32110, n32111,
    n32112, n32113, n32114, n32115, n32116, n32117,
    n32118, n32119, n32120, n32121, n32122, n32123,
    n32124, n32125, n32126, n32127, n32128, n32129,
    n32130, n32131, n32132, n32133, n32134, n32135,
    n32136, n32137, n32138, n32139, n32140, n32141,
    n32142, n32143, n32144, n32145, n32146, n32147,
    n32148, n32149, n32150, n32151, n32152, n32153,
    n32154, n32155, n32156, n32157, n32158, n32159,
    n32160, n32161, n32162, n32163, n32164, n32165,
    n32166, n32167, n32168, n32169, n32170, n32171,
    n32172, n32173, n32174, n32175, n32176, n32177,
    n32178, n32179, n32180, n32181, n32183, n32184,
    n32185, n32186, n32187, n32188, n32189, n32190,
    n32191, n32192, n32193, n32194, n32195, n32196,
    n32197, n32198, n32199, n32200, n32201, n32202,
    n32203, n32204, n32205, n32206, n32207, n32208,
    n32209, n32210, n32211, n32212, n32213, n32214,
    n32215, n32216, n32217, n32218, n32219, n32220,
    n32221, n32222, n32223, n32224, n32225, n32226,
    n32227, n32228, n32229, n32230, n32231, n32232,
    n32233, n32234, n32235, n32236, n32237, n32238,
    n32239, n32240, n32241, n32242, n32243, n32244,
    n32245, n32246, n32247, n32248, n32249, n32250,
    n32251, n32252, n32253, n32254, n32255, n32256,
    n32257, n32258, n32259, n32260, n32261, n32262,
    n32263, n32264, n32265, n32266, n32267, n32268,
    n32269, n32270, n32271, n32272, n32273, n32274,
    n32275, n32276, n32277, n32279, n32280, n32281,
    n32282, n32283, n32284, n32285, n32286, n32287,
    n32288, n32289, n32290, n32291, n32292, n32293,
    n32294, n32295, n32296, n32297, n32298, n32299,
    n32300, n32301, n32302, n32303, n32304, n32305,
    n32306, n32307, n32308, n32309, n32310, n32311,
    n32312, n32313, n32314, n32315, n32316, n32317,
    n32318, n32319, n32320, n32321, n32322, n32323,
    n32324, n32325, n32326, n32327, n32328, n32329,
    n32330, n32331, n32332, n32333, n32334, n32335,
    n32336, n32337, n32338, n32339, n32340, n32341,
    n32342, n32343, n32344, n32345, n32346, n32347,
    n32348, n32349, n32350, n32351, n32352, n32353,
    n32354, n32355, n32356, n32357, n32358, n32359,
    n32360, n32361, n32362, n32363, n32364, n32365,
    n32366, n32367, n32368, n32369, n32370, n32371,
    n32372, n32373, n32375, n32376, n32377, n32378,
    n32379, n32380, n32381, n32382, n32383, n32384,
    n32385, n32386, n32387, n32388, n32389, n32390,
    n32391, n32392, n32393, n32394, n32395, n32396,
    n32397, n32398, n32399, n32400, n32401, n32402,
    n32403, n32404, n32405, n32406, n32407, n32408,
    n32409, n32410, n32411, n32412, n32413, n32414,
    n32415, n32416, n32417, n32418, n32419, n32420,
    n32421, n32422, n32423, n32424, n32425, n32426,
    n32427, n32428, n32429, n32430, n32431, n32432,
    n32433, n32434, n32435, n32436, n32437, n32438,
    n32439, n32440, n32441, n32442, n32443, n32444,
    n32445, n32446, n32447, n32448, n32449, n32450,
    n32451, n32452, n32453, n32454, n32455, n32456,
    n32457, n32458, n32459, n32460, n32461, n32462,
    n32463, n32464, n32465, n32466, n32467, n32469,
    n32470, n32471, n32472, n32473, n32474, n32475,
    n32476, n32477, n32478, n32479, n32480, n32481,
    n32482, n32483, n32484, n32485, n32486, n32487,
    n32488, n32489, n32490, n32491, n32492, n32493,
    n32494, n32495, n32496, n32497, n32498, n32499,
    n32500, n32501, n32502, n32503, n32504, n32505,
    n32506, n32507, n32508, n32509, n32510, n32511,
    n32512, n32513, n32514, n32515, n32516, n32517,
    n32518, n32519, n32520, n32521, n32522, n32523,
    n32524, n32525, n32526, n32527, n32528, n32529,
    n32530, n32531, n32532, n32533, n32534, n32535,
    n32536, n32537, n32538, n32539, n32540, n32541,
    n32543, n32544, n32545, n32546, n32547, n32548,
    n32549, n32550, n32551, n32552, n32553, n32554,
    n32555, n32556, n32557, n32558, n32559, n32560,
    n32561, n32562, n32563, n32564, n32565, n32566,
    n32567, n32568, n32569, n32570, n32571, n32572,
    n32573, n32574, n32575, n32576, n32577, n32578,
    n32579, n32580, n32581, n32582, n32583, n32584,
    n32585, n32586, n32587, n32588, n32589, n32590,
    n32591, n32592, n32593, n32594, n32595, n32596,
    n32597, n32598, n32599, n32600, n32601, n32602,
    n32603, n32604, n32605, n32606, n32607, n32608,
    n32609, n32610, n32611, n32612, n32613, n32614,
    n32615, n32616, n32617, n32618, n32619, n32620,
    n32621, n32622, n32623, n32624, n32625, n32626,
    n32627, n32628, n32629, n32630, n32631, n32632,
    n32633, n32634, n32635, n32636, n32637, n32638,
    n32639, n32640, n32641, n32642, n32643, n32644,
    n32645, n32646, n32648, n32649, n32650, n32651,
    n32652, n32653, n32654, n32655, n32656, n32657,
    n32658, n32659, n32660, n32661, n32662, n32663,
    n32664, n32665, n32666, n32667, n32668, n32669,
    n32670, n32671, n32672, n32673, n32674, n32675,
    n32676, n32677, n32678, n32679, n32680, n32681,
    n32682, n32683, n32684, n32685, n32686, n32687,
    n32688, n32689, n32690, n32691, n32692, n32693,
    n32694, n32695, n32696, n32697, n32698, n32699,
    n32700, n32701, n32702, n32703, n32704, n32705,
    n32706, n32707, n32708, n32709, n32710, n32712,
    n32713, n32714, n32715, n32716, n32717, n32718,
    n32719, n32720, n32721, n32722, n32723, n32724,
    n32725, n32726, n32727, n32728, n32729, n32730,
    n32731, n32732, n32733, n32734, n32735, n32736,
    n32737, n32738, n32739, n32740, n32741, n32742,
    n32743, n32744, n32745, n32746, n32747, n32748,
    n32749, n32750, n32751, n32752, n32753, n32754,
    n32755, n32756, n32757, n32758, n32759, n32760,
    n32761, n32762, n32763, n32764, n32765, n32766,
    n32767, n32768, n32769, n32770, n32771, n32772,
    n32773, n32774, n32775, n32776, n32777, n32778,
    n32779, n32780, n32781, n32782, n32783, n32784,
    n32785, n32786, n32787, n32788, n32789, n32790,
    n32791, n32792, n32793, n32794, n32795, n32796,
    n32797, n32798, n32799, n32800, n32801, n32802,
    n32803, n32804, n32805, n32806, n32807, n32808,
    n32809, n32810, n32811, n32812, n32813, n32814,
    n32815, n32816, n32817, n32818, n32819, n32820,
    n32821, n32822, n32823, n32824, n32825, n32826,
    n32827, n32828, n32829, n32830, n32831, n32832,
    n32833, n32834, n32835, n32836, n32837, n32838,
    n32839, n32840, n32841, n32842, n32843, n32844,
    n32845, n32846, n32847, n32848, n32849, n32850,
    n32851, n32852, n32853, n32854, n32855, n32856,
    n32857, n32858, n32859, n32860, n32861, n32862,
    n32863, n32864, n32865, n32866, n32867, n32868,
    n32869, n32870, n32871, n32872, n32873, n32874,
    n32875, n32876, n32877, n32878, n32879, n32880,
    n32881, n32882, n32883, n32884, n32885, n32886,
    n32887, n32888, n32889, n32890, n32891, n32892,
    n32893, n32894, n32895, n32896, n32897, n32898,
    n32899, n32900, n32901, n32902, n32903, n32904,
    n32905, n32906, n32907, n32908, n32909, n32910,
    n32911, n32912, n32913, n32914, n32915, n32916,
    n32917, n32918, n32919, n32920, n32921, n32922,
    n32923, n32924, n32925, n32926, n32927, n32928,
    n32929, n32930, n32931, n32932, n32933, n32934,
    n32935, n32936, n32937, n32938, n32939, n32940,
    n32941, n32942, n32943, n32944, n32945, n32946,
    n32947, n32948, n32949, n32950, n32951, n32952,
    n32953, n32954, n32955, n32956, n32957, n32958,
    n32959, n32960, n32961, n32962, n32963, n32964,
    n32965, n32966, n32967, n32968, n32969, n32970,
    n32971, n32972, n32973, n32974, n32975, n32976,
    n32977, n32978, n32979, n32980, n32981, n32982,
    n32983, n32984, n32985, n32986, n32987, n32988,
    n32989, n32990, n32991, n32992, n32993, n32994,
    n32995, n32996, n32997, n32998, n32999, n33000,
    n33001, n33002, n33003, n33004, n33005, n33006,
    n33007, n33008, n33009, n33010, n33011, n33012,
    n33013, n33014, n33015, n33016, n33017, n33018,
    n33019, n33020, n33021, n33022, n33023, n33024,
    n33025, n33026, n33027, n33028, n33029, n33030,
    n33031, n33032, n33033, n33034, n33035, n33036,
    n33037, n33038, n33039, n33040, n33041, n33042,
    n33043, n33044, n33045, n33046, n33047, n33048,
    n33049, n33050, n33051, n33052, n33053, n33054,
    n33055, n33056, n33057, n33058, n33059, n33060,
    n33061, n33062, n33063, n33064, n33065, n33066,
    n33067, n33068, n33069, n33070, n33071, n33072,
    n33073, n33074, n33075, n33076, n33077, n33078,
    n33079, n33080, n33081, n33082, n33083, n33084,
    n33085, n33086, n33087, n33088, n33089, n33090,
    n33091, n33092, n33093, n33094, n33095, n33096,
    n33097, n33098, n33099, n33100, n33101, n33102,
    n33103, n33104, n33105, n33106, n33107, n33108,
    n33109, n33110, n33111, n33112, n33113, n33114,
    n33115, n33116, n33117, n33118, n33119, n33120,
    n33121, n33122, n33123, n33124, n33125, n33126,
    n33127, n33128, n33129, n33130, n33131, n33132,
    n33133, n33134, n33135, n33136, n33137, n33138,
    n33139, n33140, n33141, n33142, n33143, n33144,
    n33145, n33146, n33147, n33148, n33149, n33150,
    n33151, n33152, n33153, n33154, n33155, n33156,
    n33157, n33158, n33159, n33160, n33161, n33162,
    n33163, n33164, n33165, n33166, n33167, n33168,
    n33169, n33170, n33171, n33172, n33173, n33174,
    n33175, n33176, n33177, n33178, n33179, n33180,
    n33181, n33182, n33183, n33184, n33185, n33186,
    n33187, n33188, n33189, n33190, n33191, n33192,
    n33193, n33194, n33195, n33196, n33197, n33198,
    n33199, n33200, n33201, n33202, n33203, n33204,
    n33205, n33206, n33207, n33208, n33209, n33210,
    n33211, n33212, n33213, n33214, n33215, n33216,
    n33217, n33218, n33219, n33220, n33221, n33222,
    n33223, n33224, n33225, n33226, n33227, n33228,
    n33229, n33231, n33232, n33233, n33234, n33235,
    n33236, n33237, n33238, n33239, n33240, n33241,
    n33242, n33243, n33244, n33245, n33246, n33247,
    n33248, n33249, n33250, n33251, n33252, n33253,
    n33254, n33255, n33256, n33257, n33258, n33259,
    n33260, n33261, n33262, n33263, n33264, n33265,
    n33266, n33267, n33268, n33269, n33270, n33271,
    n33272, n33273, n33274, n33275, n33276, n33277,
    n33278, n33279, n33280, n33281, n33282, n33283,
    n33284, n33285, n33286, n33287, n33288, n33289,
    n33290, n33291, n33292, n33293, n33294, n33295,
    n33296, n33297, n33298, n33299, n33300, n33301,
    n33302, n33303, n33304, n33305, n33306, n33307,
    n33308, n33309, n33310, n33311, n33312, n33313,
    n33314, n33315, n33316, n33317, n33318, n33319,
    n33320, n33321, n33322, n33323, n33324, n33325,
    n33326, n33327, n33328, n33329, n33330, n33331,
    n33332, n33333, n33334, n33335, n33336, n33337,
    n33338, n33339, n33340, n33341, n33342, n33343,
    n33344, n33345, n33346, n33347, n33348, n33349,
    n33350, n33351, n33352, n33353, n33354, n33355,
    n33356, n33357, n33358, n33359, n33360, n33361,
    n33362, n33363, n33364, n33365, n33366, n33367,
    n33368, n33369, n33370, n33371, n33372, n33373,
    n33374, n33375, n33376, n33377, n33378, n33379,
    n33380, n33381, n33382, n33383, n33384, n33385,
    n33386, n33387, n33389, n33390, n33391, n33392,
    n33393, n33394, n33395, n33396, n33397, n33398,
    n33399, n33400, n33401, n33402, n33403, n33404,
    n33405, n33406, n33407, n33408, n33409, n33410,
    n33411, n33412, n33413, n33414, n33415, n33416,
    n33417, n33418, n33419, n33420, n33421, n33422,
    n33423, n33424, n33425, n33426, n33427, n33428,
    n33429, n33430, n33431, n33432, n33433, n33434,
    n33435, n33436, n33437, n33438, n33439, n33440,
    n33441, n33442, n33443, n33444, n33445, n33446,
    n33447, n33448, n33449, n33450, n33451, n33452,
    n33453, n33454, n33455, n33456, n33457, n33458,
    n33459, n33460, n33462, n33463, n33464, n33465,
    n33466, n33467, n33468, n33469, n33470, n33471,
    n33472, n33473, n33474, n33475, n33476, n33477,
    n33478, n33479, n33480, n33481, n33482, n33483,
    n33484, n33485, n33486, n33487, n33488, n33489,
    n33490, n33491, n33492, n33493, n33494, n33495,
    n33496, n33497, n33498, n33499, n33500, n33501,
    n33502, n33503, n33504, n33505, n33506, n33507,
    n33508, n33509, n33510, n33511, n33512, n33513,
    n33514, n33515, n33516, n33517, n33518, n33519,
    n33520, n33521, n33522, n33523, n33524, n33525,
    n33526, n33527, n33528, n33529, n33530, n33531,
    n33532, n33533, n33534, n33535, n33536, n33537,
    n33538, n33539, n33540, n33541, n33542, n33543,
    n33544, n33545, n33546, n33547, n33548, n33549,
    n33550, n33551, n33553, n33554, n33555, n33556,
    n33557, n33558, n33559, n33560, n33561, n33562,
    n33563, n33564, n33565, n33566, n33567, n33568,
    n33569, n33570, n33571, n33572, n33573, n33574,
    n33575, n33576, n33577, n33578, n33579, n33580,
    n33581, n33582, n33583, n33584, n33585, n33586,
    n33587, n33588, n33589, n33590, n33591, n33592,
    n33593, n33594, n33595, n33596, n33597, n33598,
    n33599, n33600, n33601, n33602, n33603, n33604,
    n33605, n33606, n33607, n33608, n33609, n33610,
    n33611, n33612, n33613, n33614, n33615, n33616,
    n33617, n33618, n33619, n33620, n33621, n33622,
    n33623, n33624, n33625, n33626, n33627, n33628,
    n33629, n33630, n33631, n33632, n33633, n33634,
    n33635, n33636, n33637, n33638, n33639, n33640,
    n33641, n33642, n33643, n33644, n33645, n33646,
    n33647, n33648, n33649, n33650, n33651, n33652,
    n33653, n33654, n33655, n33656, n33657, n33658,
    n33659, n33660, n33661, n33662, n33663, n33664,
    n33665, n33666, n33667, n33668, n33669, n33670,
    n33671, n33672, n33673, n33674, n33675, n33676,
    n33677, n33678, n33679, n33680, n33681, n33682,
    n33683, n33684, n33685, n33686, n33687, n33688,
    n33689, n33690, n33691, n33692, n33693, n33694,
    n33695, n33696, n33697, n33698, n33699, n33700,
    n33701, n33702, n33703, n33704, n33705, n33706,
    n33707, n33708, n33709, n33710, n33711, n33712,
    n33713, n33714, n33715, n33716, n33717, n33718,
    n33719, n33720, n33721, n33722, n33723, n33724,
    n33725, n33726, n33727, n33728, n33729, n33730,
    n33731, n33732, n33733, n33734, n33735, n33736,
    n33737, n33738, n33739, n33740, n33741, n33742,
    n33743, n33744, n33745, n33746, n33747, n33748,
    n33749, n33750, n33751, n33752, n33753, n33754,
    n33755, n33756, n33757, n33758, n33759, n33760,
    n33761, n33762, n33763, n33764, n33765, n33766,
    n33767, n33768, n33769, n33770, n33771, n33772,
    n33773, n33774, n33775, n33776, n33777, n33778,
    n33779, n33780, n33781, n33782, n33783, n33784,
    n33785, n33786, n33787, n33788, n33789, n33790,
    n33791, n33792, n33793, n33794, n33795, n33796,
    n33797, n33798, n33799, n33800, n33801, n33802,
    n33803, n33804, n33805, n33806, n33807, n33808,
    n33809, n33810, n33811, n33813, n33814, n33815,
    n33816, n33817, n33818, n33819, n33820, n33821,
    n33822, n33823, n33824, n33825, n33826, n33827,
    n33828, n33829, n33830, n33831, n33832, n33833,
    n33834, n33835, n33836, n33837, n33838, n33839,
    n33840, n33841, n33842, n33843, n33844, n33845,
    n33846, n33847, n33848, n33849, n33850, n33851,
    n33852, n33853, n33854, n33855, n33856, n33857,
    n33859, n33860, n33861, n33862, n33863, n33864,
    n33865, n33866, n33867, n33868, n33869, n33870,
    n33871, n33872, n33873, n33874, n33875, n33876,
    n33877, n33878, n33879, n33880, n33881, n33882,
    n33883, n33884, n33885, n33886, n33887, n33888,
    n33889, n33890, n33892, n33893, n33894, n33895,
    n33896, n33897, n33898, n33899, n33900, n33901,
    n33902, n33903, n33904, n33905, n33906, n33907,
    n33908, n33909, n33910, n33911, n33912, n33913,
    n33914, n33915, n33916, n33917, n33918, n33919,
    n33920, n33921, n33922, n33923, n33924, n33925,
    n33926, n33927, n33928, n33929, n33930, n33931,
    n33932, n33933, n33934, n33935, n33936, n33937,
    n33938, n33939, n33940, n33941, n33942, n33943,
    n33944, n33945, n33946, n33947, n33948, n33949,
    n33950, n33951, n33952, n33953, n33954, n33955,
    n33956, n33957, n33958, n33959, n33960, n33961,
    n33962, n33963, n33964, n33965, n33966, n33967,
    n33968, n33969, n33970, n33971, n33972, n33973,
    n33974, n33976, n33977, n33978, n33979, n33980,
    n33981, n33982, n33983, n33984, n33985, n33986,
    n33987, n33988, n33989, n33990, n33991, n33992,
    n33993, n33994, n33995, n33996, n33997, n33998,
    n33999, n34000, n34001, n34002, n34003, n34004,
    n34005, n34006, n34007, n34008, n34009, n34010,
    n34011, n34012, n34013, n34014, n34015, n34016,
    n34017, n34018, n34019, n34020, n34021, n34022,
    n34023, n34024, n34025, n34026, n34027, n34028,
    n34029, n34030, n34031, n34032, n34033, n34034,
    n34035, n34036, n34037, n34038, n34039, n34040,
    n34041, n34042, n34043, n34044, n34045, n34046,
    n34047, n34049, n34050, n34051, n34052, n34053,
    n34054, n34055, n34056, n34057, n34058, n34059,
    n34060, n34061, n34062, n34063, n34064, n34065,
    n34066, n34067, n34068, n34069, n34070, n34071,
    n34072, n34073, n34074, n34075, n34076, n34077,
    n34078, n34079, n34080, n34081, n34082, n34083,
    n34084, n34085, n34086, n34087, n34088, n34089,
    n34090, n34091, n34092, n34093, n34094, n34095,
    n34096, n34097, n34098, n34099, n34100, n34101,
    n34102, n34103, n34104, n34105, n34106, n34107,
    n34108, n34109, n34110, n34111, n34112, n34113,
    n34114, n34115, n34116, n34117, n34118, n34119,
    n34120, n34122, n34123, n34124, n34125, n34126,
    n34127, n34128, n34129, n34130, n34131, n34132,
    n34133, n34134, n34135, n34136, n34137, n34138,
    n34139, n34140, n34141, n34142, n34143, n34144,
    n34145, n34146, n34147, n34148, n34149, n34150,
    n34151, n34152, n34153, n34154, n34155, n34156,
    n34157, n34158, n34159, n34160, n34161, n34162,
    n34163, n34164, n34165, n34166, n34167, n34168,
    n34169, n34170, n34171, n34172, n34173, n34174,
    n34175, n34176, n34177, n34178, n34179, n34180,
    n34181, n34182, n34183, n34184, n34185, n34186,
    n34187, n34188, n34189, n34190, n34191, n34192,
    n34193, n34194, n34195, n34196, n34197, n34198,
    n34199, n34200, n34201, n34202, n34203, n34205,
    n34206, n34207, n34208, n34209, n34210, n34211,
    n34212, n34213, n34214, n34215, n34216, n34217,
    n34218, n34219, n34220, n34221, n34222, n34223,
    n34224, n34225, n34226, n34227, n34228, n34229,
    n34230, n34231, n34232, n34233, n34234, n34235,
    n34236, n34237, n34238, n34239, n34240, n34241,
    n34242, n34243, n34244, n34245, n34246, n34247,
    n34248, n34249, n34250, n34251, n34252, n34253,
    n34254, n34255, n34256, n34257, n34258, n34259,
    n34260, n34261, n34262, n34263, n34264, n34265,
    n34266, n34267, n34268, n34269, n34270, n34271,
    n34272, n34273, n34274, n34275, n34276, n34277,
    n34278, n34279, n34280, n34281, n34282, n34283,
    n34284, n34285, n34286, n34287, n34288, n34289,
    n34290, n34291, n34292, n34293, n34294, n34295,
    n34296, n34297, n34298, n34299, n34300, n34301,
    n34302, n34303, n34304, n34305, n34306, n34307,
    n34308, n34309, n34310, n34311, n34312, n34313,
    n34314, n34315, n34316, n34317, n34318, n34319,
    n34320, n34321, n34322, n34323, n34324, n34325,
    n34326, n34327, n34328, n34329, n34330, n34331,
    n34332, n34333, n34334, n34335, n34336, n34337,
    n34338, n34339, n34340, n34341, n34342, n34343,
    n34344, n34345, n34346, n34347, n34348, n34349,
    n34350, n34351, n34352, n34353, n34354, n34355,
    n34356, n34357, n34358, n34359, n34360, n34361,
    n34362, n34363, n34364, n34365, n34366, n34367,
    n34368, n34369, n34370, n34371, n34372, n34373,
    n34374, n34375, n34376, n34377, n34378, n34379,
    n34380, n34381, n34382, n34384, n34385, n34386,
    n34387, n34388, n34389, n34390, n34391, n34392,
    n34393, n34394, n34395, n34396, n34397, n34398,
    n34399, n34400, n34401, n34402, n34403, n34404,
    n34405, n34406, n34407, n34408, n34409, n34410,
    n34411, n34412, n34413, n34414, n34415, n34416,
    n34417, n34418, n34419, n34420, n34421, n34422,
    n34423, n34424, n34425, n34426, n34427, n34428,
    n34429, n34430, n34431, n34432, n34433, n34434,
    n34435, n34436, n34437, n34438, n34439, n34440,
    n34441, n34442, n34443, n34444, n34445, n34446,
    n34447, n34448, n34449, n34450, n34451, n34452,
    n34453, n34454, n34455, n34456, n34457, n34458,
    n34459, n34460, n34461, n34462, n34463, n34464,
    n34465, n34467, n34468, n34469, n34470, n34471,
    n34472, n34473, n34474, n34475, n34476, n34477,
    n34478, n34479, n34480, n34481, n34482, n34483,
    n34484, n34485, n34486, n34487, n34488, n34489,
    n34490, n34491, n34492, n34493, n34494, n34495,
    n34496, n34497, n34498, n34499, n34500, n34501,
    n34502, n34503, n34504, n34505, n34506, n34507,
    n34508, n34509, n34510, n34512, n34513, n34514,
    n34515, n34516, n34517, n34518, n34519, n34520,
    n34521, n34522, n34523, n34524, n34525, n34526,
    n34527, n34528, n34529, n34530, n34531, n34532,
    n34533, n34534, n34535, n34536, n34537, n34538,
    n34539, n34540, n34541, n34542, n34543, n34544,
    n34545, n34546, n34547, n34548, n34549, n34550,
    n34551, n34552, n34553, n34554, n34555, n34557,
    n34558, n34559, n34560, n34561, n34562, n34563,
    n34564, n34565, n34566, n34567, n34568, n34569,
    n34570, n34571, n34572, n34573, n34574, n34575,
    n34576, n34577, n34578, n34579, n34580, n34581,
    n34582, n34583, n34584, n34585, n34586, n34587,
    n34588, n34589, n34590, n34591, n34592, n34593,
    n34594, n34595, n34596, n34597, n34598, n34599,
    n34600, n34601, n34602, n34603, n34604, n34605,
    n34606, n34607, n34608, n34609, n34610, n34611,
    n34612, n34613, n34614, n34615, n34616, n34617,
    n34618, n34619, n34620, n34621, n34622, n34623,
    n34624, n34625, n34626, n34627, n34628, n34629,
    n34630, n34631, n34632, n34633, n34634, n34635,
    n34636, n34637, n34638, n34639, n34640, n34641,
    n34642, n34643, n34644, n34645, n34646, n34647,
    n34648, n34649, n34650, n34651, n34652, n34653,
    n34654, n34655, n34656, n34657, n34658, n34659,
    n34660, n34661, n34662, n34663, n34664, n34665,
    n34666, n34667, n34668, n34669, n34670, n34671,
    n34672, n34673, n34674, n34675, n34676, n34677,
    n34678, n34679, n34680, n34681, n34682, n34683,
    n34684, n34685, n34686, n34687, n34688, n34689,
    n34690, n34691, n34692, n34693, n34694, n34695,
    n34696, n34697, n34698, n34699, n34700, n34701,
    n34702, n34703, n34704, n34705, n34706, n34708,
    n34709, n34710, n34711, n34712, n34713, n34714,
    n34715, n34716, n34717, n34718, n34719, n34720,
    n34721, n34722, n34723, n34724, n34725, n34726,
    n34727, n34728, n34729, n34730, n34731, n34732,
    n34733, n34734, n34735, n34736, n34737, n34738,
    n34739, n34740, n34741, n34742, n34743, n34744,
    n34745, n34746, n34747, n34748, n34749, n34750,
    n34751, n34752, n34753, n34754, n34755, n34756,
    n34757, n34758, n34759, n34760, n34761, n34762,
    n34763, n34764, n34765, n34766, n34767, n34768,
    n34769, n34770, n34771, n34772, n34773, n34774,
    n34775, n34776, n34777, n34778, n34779, n34780,
    n34781, n34782, n34783, n34784, n34785, n34786,
    n34787, n34788, n34789, n34790, n34791, n34792,
    n34793, n34794, n34795, n34796, n34797, n34798,
    n34799, n34800, n34801, n34802, n34803, n34804,
    n34805, n34806, n34807, n34808, n34809, n34810,
    n34811, n34812, n34813, n34814, n34815, n34816,
    n34817, n34818, n34819, n34820, n34821, n34822,
    n34823, n34824, n34825, n34826, n34827, n34828,
    n34829, n34830, n34831, n34832, n34833, n34834,
    n34835, n34836, n34837, n34838, n34839, n34840,
    n34841, n34842, n34843, n34844, n34845, n34846,
    n34847, n34848, n34849, n34850, n34851, n34852,
    n34853, n34854, n34855, n34856, n34857, n34858,
    n34859, n34860, n34861, n34862, n34863, n34864,
    n34865, n34866, n34867, n34868, n34869, n34870,
    n34871, n34872, n34873, n34874, n34875, n34876,
    n34877, n34878, n34879, n34880, n34881, n34882,
    n34883, n34884, n34885, n34886, n34887, n34888,
    n34889, n34890, n34891, n34892, n34893, n34894,
    n34895, n34896, n34897, n34898, n34899, n34900,
    n34901, n34902, n34903, n34904, n34905, n34906,
    n34907, n34908, n34909, n34910, n34911, n34912,
    n34913, n34914, n34915, n34916, n34917, n34918,
    n34919, n34920, n34921, n34922, n34923, n34924,
    n34925, n34926, n34927, n34928, n34929, n34930,
    n34931, n34932, n34933, n34934, n34935, n34936,
    n34937, n34938, n34939, n34940, n34941, n34942,
    n34943, n34944, n34945, n34946, n34947, n34948,
    n34949, n34950, n34951, n34952, n34953, n34954,
    n34955, n34956, n34957, n34958, n34959, n34960,
    n34961, n34962, n34963, n34964, n34965, n34966,
    n34967, n34968, n34969, n34970, n34971, n34972,
    n34973, n34974, n34975, n34976, n34977, n34978,
    n34979, n34980, n34981, n34982, n34983, n34984,
    n34985, n34986, n34987, n34988, n34989, n34990,
    n34991, n34992, n34993, n34994, n34995, n34996,
    n34997, n34998, n34999, n35000, n35001, n35002,
    n35003, n35004, n35005, n35006, n35007, n35008,
    n35009, n35010, n35011, n35012, n35013, n35014,
    n35015, n35016, n35017, n35018, n35019, n35020,
    n35021, n35022, n35023, n35024, n35025, n35026,
    n35027, n35028, n35029, n35030, n35031, n35032,
    n35033, n35034, n35035, n35036, n35037, n35038,
    n35039, n35040, n35041, n35042, n35043, n35044,
    n35045, n35046, n35047, n35048, n35049, n35050,
    n35051, n35052, n35053, n35054, n35055, n35056,
    n35057, n35058, n35059, n35060, n35061, n35062,
    n35063, n35064, n35065, n35066, n35067, n35068,
    n35069, n35070, n35071, n35072, n35073, n35074,
    n35075, n35076, n35077, n35078, n35079, n35080,
    n35081, n35082, n35083, n35084, n35085, n35086,
    n35087, n35088, n35089, n35090, n35091, n35092,
    n35093, n35094, n35095, n35096, n35097, n35098,
    n35099, n35100, n35101, n35102, n35103, n35104,
    n35105, n35106, n35107, n35108, n35109, n35110,
    n35111, n35112, n35113, n35114, n35115, n35116,
    n35117, n35118, n35119, n35120, n35121, n35122,
    n35123, n35124, n35125, n35126, n35127, n35128,
    n35129, n35130, n35131, n35132, n35133, n35134,
    n35135, n35136, n35137, n35138, n35139, n35140,
    n35141, n35142, n35143, n35144, n35145, n35146,
    n35147, n35148, n35149, n35150, n35151, n35152,
    n35153, n35154, n35155, n35156, n35157, n35158,
    n35159, n35160, n35161, n35162, n35163, n35164,
    n35165, n35166, n35167, n35168, n35169, n35170,
    n35171, n35172, n35173, n35174, n35175, n35176,
    n35177, n35178, n35179, n35180, n35181, n35182,
    n35183, n35184, n35185, n35186, n35187, n35188,
    n35189, n35190, n35191, n35192, n35193, n35194,
    n35195, n35196, n35197, n35198, n35199, n35200,
    n35201, n35202, n35203, n35204, n35205, n35206,
    n35207, n35208, n35209, n35210, n35211, n35212,
    n35213, n35214, n35215, n35216, n35217, n35218,
    n35219, n35220, n35221, n35222, n35223, n35224,
    n35225, n35226, n35227, n35228, n35229, n35230,
    n35231, n35232, n35233, n35234, n35235, n35236,
    n35237, n35238, n35239, n35240, n35241, n35242,
    n35243, n35244, n35245, n35246, n35247, n35248,
    n35249, n35250, n35251, n35252, n35253, n35254,
    n35255, n35256, n35257, n35258, n35259, n35260,
    n35261, n35262, n35263, n35264, n35265, n35266,
    n35267, n35268, n35269, n35270, n35271, n35273,
    n35274, n35275, n35276, n35277, n35278, n35279,
    n35280, n35281, n35282, n35283, n35284, n35285,
    n35287, n35288, n35289, n35290, n35291, n35292,
    n35293, n35294, n35295, n35296, n35297, n35298,
    n35299, n35300, n35301, n35302, n35303, n35304,
    n35305, n35306, n35307, n35308, n35309, n35310,
    n35311, n35312, n35313, n35314, n35315, n35316,
    n35317, n35318, n35319, n35320, n35321, n35322,
    n35323, n35324, n35325, n35326, n35327, n35328,
    n35329, n35330, n35331, n35332, n35333, n35334,
    n35335, n35336, n35337, n35338, n35339, n35340,
    n35341, n35342, n35343, n35344, n35345, n35346,
    n35347, n35348, n35349, n35350, n35351, n35352,
    n35353, n35354, n35355, n35356, n35357, n35358,
    n35359, n35360, n35361, n35362, n35363, n35364,
    n35365, n35366, n35367, n35368, n35369, n35370,
    n35371, n35372, n35373, n35374, n35375, n35376,
    n35377, n35378, n35379, n35380, n35381, n35382,
    n35383, n35384, n35385, n35386, n35387, n35388,
    n35389, n35390, n35391, n35392, n35393, n35394,
    n35395, n35396, n35397, n35398, n35399, n35400,
    n35401, n35402, n35403, n35404, n35405, n35406,
    n35407, n35408, n35409, n35410, n35411, n35412,
    n35413, n35414, n35415, n35416, n35417, n35418,
    n35419, n35420, n35421, n35422, n35423, n35424,
    n35425, n35426, n35427, n35428, n35429, n35430,
    n35431, n35432, n35433, n35434, n35435, n35436,
    n35437, n35438, n35439, n35440, n35441, n35442,
    n35443, n35444, n35445, n35446, n35447, n35448,
    n35449, n35450, n35451, n35452, n35453, n35454,
    n35455, n35456, n35457, n35458, n35459, n35460,
    n35461, n35462, n35463, n35464, n35465, n35466,
    n35467, n35468, n35469, n35470, n35471, n35472,
    n35473, n35474, n35475, n35476, n35477, n35478,
    n35479, n35480, n35481, n35482, n35483, n35484,
    n35485, n35486, n35487, n35488, n35489, n35490,
    n35491, n35492, n35493, n35494, n35495, n35496,
    n35497, n35498, n35499, n35500, n35501, n35502,
    n35503, n35504, n35505, n35506, n35507, n35508,
    n35509, n35510, n35511, n35512, n35513, n35514,
    n35515, n35516, n35517, n35518, n35519, n35520,
    n35521, n35522, n35523, n35524, n35525, n35526,
    n35527, n35528, n35529, n35530, n35531, n35532,
    n35533, n35534, n35535, n35536, n35537, n35538,
    n35539, n35540, n35541, n35542, n35543, n35544,
    n35545, n35546, n35547, n35548, n35549, n35550,
    n35551, n35552, n35553, n35554, n35555, n35556,
    n35557, n35558, n35559, n35560, n35561, n35562,
    n35563, n35564, n35565, n35566, n35567, n35568,
    n35569, n35570, n35572, n35573, n35574, n35575,
    n35576, n35577, n35578, n35579, n35580, n35581,
    n35582, n35583, n35584, n35585, n35586, n35587,
    n35588, n35589, n35590, n35591, n35592, n35593,
    n35594, n35595, n35596, n35597, n35598, n35599,
    n35600, n35601, n35602, n35604, n35605, n35606,
    n35607, n35608, n35609, n35610, n35611, n35612,
    n35613, n35614, n35615, n35616, n35617, n35618,
    n35619, n35620, n35621, n35622, n35623, n35624,
    n35625, n35626, n35627, n35628, n35629, n35630,
    n35631, n35632, n35633, n35634, n35635, n35636,
    n35637, n35638, n35639, n35640, n35641, n35643,
    n35644, n35645, n35646, n35647, n35648, n35649,
    n35650, n35651, n35652, n35653, n35654, n35655,
    n35657, n35658, n35659, n35660, n35661, n35662,
    n35663, n35664, n35665, n35666, n35667, n35668,
    n35669, n35670, n35671, n35672, n35673, n35674,
    n35675, n35676, n35677, n35678, n35679, n35680,
    n35681, n35682, n35683, n35684, n35685, n35686,
    n35687, n35688, n35689, n35690, n35691, n35692,
    n35693, n35694, n35695, n35696, n35697, n35698,
    n35699, n35700, n35701, n35702, n35703, n35704,
    n35705, n35706, n35707, n35708, n35709, n35710,
    n35711, n35712, n35713, n35714, n35715, n35716,
    n35717, n35718, n35719, n35720, n35721, n35722,
    n35723, n35724, n35725, n35726, n35727, n35728,
    n35729, n35730, n35731, n35732, n35733, n35734,
    n35735, n35736, n35737, n35738, n35739, n35740,
    n35741, n35742, n35743, n35744, n35745, n35746,
    n35747, n35748, n35749, n35750, n35751, n35752,
    n35753, n35754, n35755, n35756, n35757, n35758,
    n35759, n35760, n35761, n35762, n35763, n35764,
    n35765, n35766, n35767, n35768, n35769, n35770,
    n35771, n35772, n35773, n35774, n35775, n35776,
    n35777, n35778, n35779, n35780, n35781, n35782,
    n35783, n35784, n35785, n35786, n35787, n35788,
    n35789, n35790, n35791, n35792, n35793, n35794,
    n35795, n35796, n35797, n35798, n35799, n35800,
    n35801, n35802, n35803, n35804, n35805, n35806,
    n35807, n35808, n35809, n35810, n35811, n35812,
    n35813, n35814, n35815, n35816, n35817, n35818,
    n35819, n35820, n35821, n35822, n35823, n35824,
    n35825, n35826, n35827, n35828, n35829, n35830,
    n35831, n35832, n35833, n35834, n35835, n35836,
    n35837, n35838, n35839, n35840, n35841, n35842,
    n35843, n35844, n35845, n35846, n35847, n35848,
    n35849, n35850, n35851, n35852, n35853, n35854,
    n35855, n35856, n35857, n35858, n35859, n35860,
    n35861, n35862, n35863, n35864, n35865, n35866,
    n35867, n35868, n35869, n35870, n35871, n35872,
    n35873, n35874, n35875, n35876, n35877, n35878,
    n35879, n35880, n35881, n35882, n35883, n35884,
    n35885, n35886, n35887, n35888, n35889, n35890,
    n35891, n35892, n35893, n35894, n35895, n35896,
    n35897, n35898, n35899, n35900, n35901, n35902,
    n35903, n35904, n35905, n35906, n35907, n35908,
    n35909, n35910, n35911, n35912, n35913, n35914,
    n35915, n35916, n35917, n35918, n35919, n35920,
    n35921, n35922, n35923, n35924, n35925, n35926,
    n35927, n35928, n35929, n35930, n35931, n35932,
    n35933, n35934, n35935, n35936, n35937, n35938,
    n35939, n35940, n35941, n35942, n35943, n35944,
    n35945, n35947, n35948, n35949, n35950, n35951,
    n35952, n35953, n35954, n35955, n35956, n35957,
    n35958, n35959, n35960, n35961, n35962, n35963,
    n35964, n35965, n35966, n35967, n35968, n35969,
    n35970, n35971, n35972, n35973, n35974, n35975,
    n35976, n35977, n35978, n35979, n35980, n35981,
    n35982, n35983, n35984, n35985, n35986, n35987,
    n35988, n35989, n35990, n35991, n35992, n35993,
    n35994, n35995, n35996, n35997, n35998, n35999,
    n36000, n36001, n36002, n36003, n36004, n36005,
    n36006, n36007, n36008, n36009, n36010, n36011,
    n36012, n36013, n36014, n36015, n36016, n36017,
    n36018, n36019, n36020, n36021, n36022, n36023,
    n36024, n36025, n36026, n36027, n36028, n36029,
    n36030, n36031, n36032, n36033, n36034, n36035,
    n36036, n36037, n36038, n36039, n36040, n36041,
    n36042, n36043, n36044, n36045, n36046, n36047,
    n36048, n36049, n36050, n36051, n36052, n36053,
    n36054, n36055, n36056, n36057, n36058, n36059,
    n36060, n36061, n36062, n36063, n36064, n36065,
    n36066, n36067, n36068, n36069, n36070, n36071,
    n36072, n36073, n36074, n36075, n36076, n36077,
    n36078, n36079, n36080, n36081, n36082, n36083,
    n36085, n36086, n36087, n36088, n36089, n36090,
    n36091, n36092, n36093, n36094, n36095, n36096,
    n36097, n36098, n36099, n36100, n36101, n36102,
    n36103, n36104, n36105, n36106, n36107, n36108,
    n36109, n36110, n36111, n36112, n36113, n36114,
    n36115, n36116, n36117, n36118, n36119, n36120,
    n36121, n36122, n36123, n36124, n36125, n36126,
    n36127, n36128, n36129, n36130, n36131, n36132,
    n36133, n36134, n36135, n36136, n36137, n36138,
    n36139, n36140, n36141, n36142, n36143, n36144,
    n36145, n36146, n36147, n36148, n36149, n36150,
    n36151, n36152, n36153, n36154, n36155, n36156,
    n36157, n36158, n36159, n36160, n36161, n36162,
    n36163, n36164, n36165, n36166, n36167, n36168,
    n36169, n36170, n36171, n36172, n36173, n36174,
    n36175, n36176, n36177, n36178, n36179, n36180,
    n36181, n36182, n36183, n36185, n36186, n36187,
    n36188, n36189, n36190, n36191, n36192, n36193,
    n36194, n36195, n36196, n36197, n36198, n36199,
    n36200, n36201, n36202, n36203, n36204, n36205,
    n36206, n36207, n36208, n36209, n36210, n36211,
    n36212, n36213, n36214, n36215, n36216, n36217,
    n36218, n36219, n36220, n36221, n36222, n36223,
    n36224, n36225, n36226, n36227, n36228, n36229,
    n36230, n36231, n36232, n36233, n36234, n36235,
    n36236, n36237, n36238, n36239, n36240, n36241,
    n36242, n36243, n36244, n36245, n36246, n36247,
    n36248, n36249, n36250, n36251, n36252, n36253,
    n36254, n36255, n36256, n36257, n36258, n36259,
    n36260, n36261, n36262, n36263, n36264, n36266,
    n36267, n36268, n36269, n36270, n36271, n36272,
    n36273, n36274, n36275, n36276, n36277, n36278,
    n36279, n36280, n36281, n36282, n36283, n36284,
    n36285, n36286, n36287, n36288, n36289, n36290,
    n36291, n36293, n36294, n36295, n36296, n36297,
    n36298, n36299, n36300, n36301, n36302, n36303,
    n36304, n36306, n36307, n36308, n36309, n36310,
    n36311, n36312, n36313, n36314, n36315, n36316,
    n36317, n36318, n36319, n36320, n36321, n36322,
    n36323, n36324, n36325, n36326, n36327, n36328,
    n36329, n36330, n36331, n36332, n36333, n36334,
    n36335, n36336, n36337, n36338, n36339, n36340,
    n36341, n36342, n36343, n36344, n36345, n36346,
    n36347, n36348, n36349, n36350, n36351, n36352,
    n36353, n36354, n36355, n36356, n36357, n36358,
    n36359, n36360, n36361, n36362, n36363, n36364,
    n36365, n36366, n36367, n36368, n36369, n36370,
    n36371, n36372, n36373, n36374, n36375, n36376,
    n36377, n36378, n36379, n36380, n36381, n36382,
    n36383, n36384, n36385, n36386, n36387, n36388,
    n36389, n36390, n36391, n36392, n36393, n36394,
    n36395, n36396, n36397, n36398, n36399, n36400,
    n36401, n36402, n36403, n36404, n36405, n36406,
    n36407, n36408, n36409, n36410, n36411, n36412,
    n36413, n36414, n36415, n36416, n36417, n36418,
    n36419, n36420, n36421, n36422, n36423, n36424,
    n36425, n36426, n36427, n36428, n36429, n36430,
    n36431, n36432, n36433, n36434, n36435, n36436,
    n36437, n36438, n36439, n36440, n36441, n36442,
    n36443, n36444, n36445, n36446, n36447, n36448,
    n36449, n36450, n36451, n36452, n36453, n36454,
    n36455, n36456, n36457, n36458, n36459, n36460,
    n36461, n36462, n36463, n36464, n36465, n36466,
    n36467, n36468, n36469, n36470, n36471, n36472,
    n36473, n36474, n36475, n36476, n36477, n36478,
    n36479, n36480, n36481, n36482, n36483, n36484,
    n36485, n36486, n36487, n36488, n36489, n36490,
    n36491, n36492, n36493, n36494, n36495, n36496,
    n36497, n36498, n36499, n36500, n36501, n36502,
    n36503, n36504, n36505, n36506, n36507, n36508,
    n36509, n36510, n36511, n36512, n36513, n36514,
    n36515, n36516, n36517, n36518, n36519, n36520,
    n36521, n36522, n36523, n36524, n36525, n36526,
    n36527, n36528, n36529, n36530, n36531, n36532,
    n36533, n36534, n36535, n36536, n36537, n36538,
    n36539, n36540, n36541, n36542, n36543, n36544,
    n36545, n36546, n36547, n36548, n36549, n36550,
    n36551, n36552, n36553, n36554, n36555, n36556,
    n36557, n36558, n36559, n36560, n36561, n36562,
    n36563, n36564, n36565, n36566, n36567, n36568,
    n36569, n36570, n36571, n36572, n36573, n36574,
    n36575, n36576, n36577, n36578, n36579, n36580,
    n36581, n36582, n36583, n36584, n36585, n36586,
    n36587, n36588, n36589, n36590, n36591, n36592,
    n36593, n36594, n36595, n36596, n36597, n36598,
    n36599, n36600, n36601, n36602, n36603, n36604,
    n36605, n36606, n36607, n36608, n36609, n36610,
    n36611, n36612, n36613, n36614, n36615, n36616,
    n36617, n36618, n36619, n36620, n36621, n36622,
    n36623, n36624, n36625, n36626, n36627, n36628,
    n36629, n36630, n36631, n36632, n36633, n36634,
    n36635, n36636, n36637, n36638, n36639, n36640,
    n36641, n36642, n36643, n36644, n36645, n36646,
    n36647, n36648, n36649, n36650, n36651, n36652,
    n36653, n36654, n36655, n36656, n36657, n36658,
    n36659, n36660, n36661, n36662, n36663, n36664,
    n36665, n36666, n36667, n36668, n36669, n36670,
    n36671, n36672, n36673, n36674, n36675, n36676,
    n36677, n36678, n36679, n36680, n36681, n36682,
    n36683, n36684, n36685, n36686, n36687, n36688,
    n36689, n36690, n36691, n36692, n36693, n36694,
    n36695, n36696, n36697, n36698, n36699, n36700,
    n36701, n36702, n36703, n36704, n36705, n36706,
    n36707, n36708, n36709, n36710, n36711, n36712,
    n36713, n36714, n36715, n36716, n36717, n36718,
    n36719, n36720, n36721, n36722, n36723, n36724,
    n36725, n36726, n36727, n36728, n36729, n36730,
    n36731, n36732, n36733, n36734, n36735, n36736,
    n36737, n36738, n36739, n36740, n36741, n36742,
    n36743, n36744, n36745, n36746, n36747, n36748,
    n36749, n36750, n36751, n36752, n36753, n36754,
    n36755, n36756, n36757, n36758, n36759, n36760,
    n36761, n36762, n36763, n36764, n36765, n36766,
    n36767, n36768, n36769, n36770, n36771, n36772,
    n36773, n36774, n36775, n36776, n36777, n36778,
    n36779, n36780, n36781, n36782, n36783, n36784,
    n36785, n36786, n36787, n36788, n36789, n36790,
    n36791, n36792, n36793, n36794, n36795, n36796,
    n36797, n36798, n36799, n36800, n36801, n36802,
    n36803, n36804, n36805, n36806, n36807, n36808,
    n36809, n36810, n36811, n36812, n36813, n36814,
    n36815, n36816, n36817, n36818, n36819, n36820,
    n36821, n36822, n36823, n36824, n36825, n36826,
    n36827, n36828, n36829, n36830, n36831, n36832,
    n36833, n36834, n36835, n36836, n36837, n36838,
    n36839, n36840, n36841, n36842, n36843, n36844,
    n36845, n36846, n36847, n36848, n36849, n36850,
    n36851, n36852, n36853, n36854, n36855, n36856,
    n36857, n36858, n36859, n36860, n36861, n36862,
    n36863, n36864, n36865, n36866, n36867, n36868,
    n36869, n36870, n36871, n36872, n36873, n36874,
    n36875, n36876, n36877, n36878, n36879, n36880,
    n36881, n36882, n36883, n36884, n36885, n36886,
    n36887, n36888, n36889, n36890, n36891, n36892,
    n36893, n36894, n36895, n36896, n36897, n36898,
    n36899, n36900, n36901, n36902, n36903, n36904,
    n36905, n36906, n36907, n36908, n36909, n36910,
    n36911, n36912, n36913, n36914, n36915, n36916,
    n36917, n36918, n36919, n36920, n36921, n36922,
    n36923, n36924, n36925, n36926, n36927, n36928,
    n36929, n36930, n36931, n36932, n36933, n36934,
    n36935, n36936, n36937, n36938, n36939, n36940,
    n36941, n36942, n36943, n36944, n36945, n36946,
    n36947, n36948, n36949, n36950, n36951, n36952,
    n36953, n36954, n36955, n36956, n36957, n36958,
    n36959, n36960, n36961, n36962, n36963, n36964,
    n36965, n36966, n36967, n36968, n36969, n36970,
    n36971, n36972, n36973, n36974, n36975, n36976,
    n36977, n36978, n36979, n36980, n36981, n36982,
    n36983, n36984, n36985, n36986, n36987, n36988,
    n36989, n36990, n36991, n36992, n36993, n36994,
    n36995, n36996, n36997, n36998, n36999, n37000,
    n37001, n37002, n37003, n37004, n37005, n37006,
    n37007, n37008, n37009, n37010, n37011, n37012,
    n37013, n37014, n37015, n37016, n37017, n37018,
    n37019, n37020, n37021, n37022, n37023, n37024,
    n37025, n37026, n37027, n37028, n37029, n37030,
    n37031, n37032, n37033, n37034, n37035, n37036,
    n37037, n37038, n37039, n37040, n37041, n37042,
    n37043, n37044, n37045, n37046, n37047, n37049,
    n37050, n37051, n37052, n37053, n37054, n37055,
    n37057, n37058, n37059, n37060, n37061, n37062,
    n37063, n37064, n37065, n37066, n37067, n37068,
    n37070, n37071, n37072, n37073, n37074, n37075,
    n37076, n37077, n37078, n37079, n37080, n37081,
    n37082, n37083, n37084, n37085, n37086, n37087,
    n37088, n37089, n37090, n37091, n37092, n37093,
    n37094, n37095, n37096, n37097, n37098, n37099,
    n37100, n37101, n37102, n37103, n37104, n37105,
    n37106, n37107, n37108, n37109, n37110, n37111,
    n37112, n37113, n37114, n37115, n37116, n37117,
    n37118, n37119, n37120, n37121, n37122, n37123,
    n37124, n37125, n37126, n37127, n37128, n37129,
    n37130, n37131, n37132, n37133, n37134, n37135,
    n37136, n37137, n37138, n37139, n37140, n37141,
    n37142, n37143, n37144, n37145, n37146, n37147,
    n37148, n37149, n37150, n37151, n37152, n37153,
    n37154, n37155, n37156, n37157, n37158, n37159,
    n37160, n37161, n37162, n37163, n37164, n37165,
    n37166, n37167, n37168, n37169, n37170, n37171,
    n37172, n37173, n37174, n37175, n37176, n37177,
    n37178, n37179, n37180, n37181, n37182, n37183,
    n37184, n37185, n37186, n37187, n37188, n37189,
    n37190, n37191, n37192, n37193, n37194, n37195,
    n37196, n37197, n37198, n37199, n37200, n37201,
    n37202, n37203, n37204, n37205, n37206, n37207,
    n37208, n37209, n37210, n37211, n37212, n37213,
    n37214, n37215, n37216, n37217, n37218, n37219,
    n37220, n37221, n37222, n37223, n37224, n37225,
    n37226, n37227, n37228, n37229, n37230, n37231,
    n37232, n37233, n37234, n37235, n37236, n37237,
    n37238, n37239, n37240, n37241, n37242, n37243,
    n37244, n37245, n37246, n37247, n37248, n37249,
    n37250, n37251, n37252, n37253, n37255, n37256,
    n37257, n37259, n37260, n37261, n37262, n37263,
    n37264, n37265, n37266, n37267, n37268, n37269,
    n37270, n37271, n37272, n37273, n37274, n37275,
    n37276, n37277, n37278, n37279, n37280, n37281,
    n37282, n37283, n37284, n37285, n37286, n37287,
    n37288, n37289, n37290, n37291, n37292, n37293,
    n37294, n37295, n37296, n37297, n37298, n37299,
    n37300, n37301, n37302, n37304, n37305, n37306,
    n37307, n37308, n37309, n37310, n37311, n37312,
    n37313, n37314, n37315, n37316, n37317, n37318,
    n37319, n37320, n37321, n37322, n37323, n37324,
    n37325, n37326, n37327, n37328, n37329, n37330,
    n37331, n37332, n37333, n37334, n37335, n37336,
    n37337, n37338, n37339, n37340, n37341, n37342,
    n37343, n37344, n37345, n37346, n37347, n37348,
    n37349, n37350, n37351, n37352, n37353, n37354,
    n37355, n37356, n37357, n37358, n37359, n37360,
    n37361, n37362, n37363, n37364, n37365, n37366,
    n37368, n37369, n37370, n37371, n37372, n37373,
    n37374, n37375, n37376, n37377, n37378, n37379,
    n37380, n37381, n37382, n37383, n37384, n37385,
    n37386, n37387, n37388, n37389, n37390, n37391,
    n37392, n37393, n37394, n37395, n37396, n37397,
    n37398, n37399, n37400, n37401, n37402, n37403,
    n37404, n37405, n37406, n37407, n37408, n37409,
    n37410, n37411, n37412, n37413, n37414, n37415,
    n37416, n37417, n37418, n37419, n37420, n37421,
    n37422, n37423, n37424, n37425, n37426, n37427,
    n37428, n37429, n37430, n37431, n37432, n37433,
    n37434, n37435, n37436, n37437, n37438, n37439,
    n37440, n37441, n37442, n37444, n37445, n37446,
    n37447, n37448, n37449, n37450, n37451, n37452,
    n37453, n37454, n37455, n37456, n37457, n37458,
    n37459, n37460, n37461, n37462, n37463, n37464,
    n37465, n37466, n37467, n37468, n37469, n37470,
    n37471, n37472, n37473, n37474, n37475, n37476,
    n37477, n37478, n37479, n37480, n37481, n37482,
    n37483, n37484, n37485, n37486, n37487, n37488,
    n37489, n37490, n37491, n37492, n37493, n37494,
    n37495, n37496, n37497, n37498, n37499, n37500,
    n37501, n37502, n37503, n37504, n37505, n37506,
    n37507, n37508, n37509, n37510, n37511, n37512,
    n37513, n37514, n37515, n37516, n37517, n37518,
    n37519, n37520, n37521, n37522, n37523, n37524,
    n37525, n37526, n37527, n37528, n37529, n37530,
    n37531, n37532, n37533, n37534, n37535, n37536,
    n37537, n37538, n37539, n37540, n37541, n37542,
    n37543, n37544, n37546, n37547, n37548, n37549,
    n37550, n37551, n37552, n37553, n37554, n37555,
    n37556, n37557, n37558, n37559, n37560, n37561,
    n37562, n37563, n37564, n37565, n37566, n37567,
    n37568, n37569, n37570, n37571, n37572, n37573,
    n37574, n37575, n37576, n37577, n37578, n37579,
    n37580, n37581, n37582, n37583, n37584, n37585,
    n37586, n37587, n37588, n37589, n37590, n37591,
    n37592, n37593, n37594, n37595, n37596, n37597,
    n37598, n37599, n37600, n37601, n37602, n37603,
    n37604, n37605, n37606, n37607, n37608, n37609,
    n37610, n37611, n37612, n37613, n37614, n37615,
    n37616, n37617, n37618, n37619, n37620, n37621,
    n37622, n37623, n37624, n37625, n37626, n37627,
    n37628, n37629, n37630, n37631, n37632, n37633,
    n37634, n37635, n37636, n37637, n37638, n37639,
    n37640, n37641, n37642, n37643, n37644, n37645,
    n37646, n37647, n37648, n37649, n37650, n37651,
    n37652, n37653, n37654, n37655, n37656, n37657,
    n37658, n37659, n37660, n37661, n37662, n37663,
    n37664, n37665, n37666, n37667, n37668, n37669,
    n37670, n37671, n37672, n37673, n37674, n37675,
    n37676, n37677, n37678, n37679, n37680, n37681,
    n37682, n37683, n37684, n37685, n37686, n37687,
    n37688, n37689, n37690, n37691, n37692, n37693,
    n37694, n37695, n37696, n37697, n37698, n37699,
    n37700, n37701, n37702, n37703, n37704, n37705,
    n37706, n37707, n37708, n37709, n37710, n37711,
    n37712, n37713, n37714, n37715, n37716, n37717,
    n37718, n37719, n37720, n37721, n37722, n37723,
    n37724, n37725, n37726, n37727, n37728, n37729,
    n37730, n37731, n37732, n37733, n37734, n37735,
    n37736, n37737, n37738, n37739, n37740, n37741,
    n37742, n37743, n37744, n37745, n37746, n37747,
    n37748, n37749, n37750, n37751, n37752, n37753,
    n37754, n37755, n37756, n37757, n37758, n37759,
    n37760, n37761, n37762, n37763, n37764, n37765,
    n37766, n37767, n37768, n37769, n37770, n37771,
    n37772, n37773, n37774, n37775, n37776, n37777,
    n37778, n37779, n37780, n37781, n37782, n37783,
    n37784, n37785, n37786, n37787, n37788, n37789,
    n37790, n37791, n37792, n37793, n37794, n37795,
    n37796, n37797, n37798, n37799, n37800, n37801,
    n37802, n37803, n37804, n37805, n37806, n37807,
    n37808, n37809, n37810, n37811, n37812, n37813,
    n37814, n37815, n37816, n37817, n37818, n37819,
    n37820, n37821, n37822, n37823, n37824, n37825,
    n37826, n37827, n37828, n37829, n37830, n37831,
    n37832, n37833, n37834, n37835, n37836, n37837,
    n37838, n37839, n37840, n37841, n37842, n37843,
    n37844, n37845, n37846, n37847, n37848, n37849,
    n37850, n37851, n37852, n37853, n37854, n37855,
    n37856, n37857, n37858, n37859, n37860, n37861,
    n37862, n37863, n37864, n37865, n37866, n37867,
    n37868, n37869, n37870, n37871, n37872, n37873,
    n37874, n37875, n37876, n37877, n37878, n37879,
    n37880, n37881, n37882, n37883, n37884, n37885,
    n37886, n37887, n37888, n37889, n37890, n37891,
    n37892, n37893, n37894, n37895, n37896, n37897,
    n37898, n37899, n37900, n37901, n37902, n37903,
    n37904, n37905, n37906, n37907, n37908, n37909,
    n37910, n37911, n37912, n37913, n37914, n37915,
    n37916, n37917, n37918, n37919, n37920, n37921,
    n37922, n37923, n37924, n37925, n37926, n37927,
    n37928, n37929, n37930, n37931, n37932, n37933,
    n37934, n37935, n37936, n37937, n37938, n37939,
    n37940, n37941, n37942, n37943, n37944, n37945,
    n37946, n37947, n37948, n37949, n37950, n37951,
    n37952, n37953, n37954, n37955, n37956, n37957,
    n37958, n37959, n37960, n37961, n37962, n37963,
    n37964, n37965, n37966, n37967, n37968, n37969,
    n37970, n37971, n37972, n37973, n37974, n37975,
    n37976, n37977, n37978, n37979, n37980, n37981,
    n37982, n37983, n37984, n37985, n37986, n37987,
    n37988, n37989, n37990, n37991, n37992, n37993,
    n37994, n37995, n37996, n37997, n37998, n37999,
    n38000, n38001, n38002, n38003, n38004, n38005,
    n38006, n38007, n38008, n38009, n38010, n38011,
    n38012, n38013, n38014, n38015, n38016, n38017,
    n38018, n38019, n38020, n38021, n38022, n38023,
    n38024, n38025, n38026, n38027, n38028, n38029,
    n38030, n38031, n38032, n38033, n38034, n38035,
    n38036, n38037, n38038, n38039, n38040, n38041,
    n38042, n38043, n38044, n38045, n38046, n38047,
    n38049, n38050, n38051, n38052, n38053, n38054,
    n38055, n38056, n38057, n38058, n38059, n38060,
    n38061, n38062, n38063, n38064, n38065, n38066,
    n38067, n38068, n38069, n38070, n38071, n38072,
    n38073, n38074, n38075, n38076, n38077, n38078,
    n38079, n38080, n38081, n38082, n38083, n38084,
    n38085, n38086, n38087, n38088, n38089, n38090,
    n38091, n38092, n38093, n38094, n38095, n38096,
    n38097, n38098, n38099, n38101, n38102, n38103,
    n38104, n38105, n38106, n38107, n38108, n38109,
    n38110, n38111, n38112, n38113, n38114, n38115,
    n38116, n38117, n38118, n38119, n38120, n38121,
    n38122, n38123, n38124, n38125, n38126, n38127,
    n38128, n38129, n38130, n38131, n38132, n38133,
    n38134, n38135, n38136, n38137, n38138, n38139,
    n38140, n38141, n38142, n38143, n38144, n38145,
    n38146, n38147, n38149, n38150, n38151, n38152,
    n38153, n38154, n38155, n38156, n38157, n38158,
    n38159, n38160, n38161, n38162, n38163, n38164,
    n38165, n38166, n38167, n38168, n38169, n38170,
    n38171, n38172, n38173, n38174, n38175, n38176,
    n38177, n38178, n38179, n38180, n38181, n38182,
    n38183, n38184, n38185, n38186, n38187, n38188,
    n38189, n38190, n38191, n38192, n38193, n38194,
    n38195, n38196, n38197, n38198, n38199, n38200,
    n38201, n38202, n38203, n38204, n38205, n38207,
    n38208, n38209, n38210, n38211, n38212, n38213,
    n38214, n38215, n38216, n38217, n38218, n38219,
    n38220, n38221, n38222, n38223, n38224, n38225,
    n38226, n38227, n38228, n38229, n38230, n38231,
    n38232, n38233, n38234, n38235, n38236, n38237,
    n38238, n38239, n38240, n38241, n38242, n38243,
    n38244, n38245, n38246, n38247, n38248, n38249,
    n38250, n38251, n38252, n38253, n38254, n38255,
    n38256, n38257, n38258, n38259, n38260, n38261,
    n38262, n38263, n38264, n38265, n38266, n38267,
    n38268, n38269, n38270, n38271, n38272, n38273,
    n38274, n38275, n38276, n38277, n38278, n38279,
    n38280, n38281, n38282, n38283, n38284, n38285,
    n38286, n38287, n38288, n38289, n38290, n38291,
    n38292, n38293, n38294, n38295, n38296, n38297,
    n38298, n38299, n38300, n38301, n38302, n38303,
    n38304, n38305, n38306, n38307, n38308, n38309,
    n38310, n38311, n38312, n38313, n38314, n38315,
    n38316, n38317, n38318, n38319, n38320, n38321,
    n38322, n38323, n38324, n38325, n38326, n38327,
    n38328, n38329, n38330, n38331, n38332, n38333,
    n38334, n38335, n38336, n38337, n38338, n38339,
    n38340, n38341, n38342, n38343, n38344, n38345,
    n38346, n38347, n38348, n38349, n38350, n38351,
    n38352, n38353, n38354, n38355, n38356, n38357,
    n38358, n38359, n38360, n38361, n38362, n38363,
    n38364, n38365, n38366, n38367, n38368, n38369,
    n38370, n38371, n38372, n38373, n38374, n38375,
    n38376, n38377, n38378, n38379, n38380, n38381,
    n38382, n38383, n38384, n38385, n38386, n38387,
    n38388, n38389, n38390, n38391, n38392, n38393,
    n38394, n38395, n38396, n38397, n38398, n38399,
    n38400, n38401, n38402, n38403, n38404, n38405,
    n38406, n38407, n38408, n38409, n38410, n38411,
    n38412, n38413, n38414, n38415, n38416, n38417,
    n38418, n38419, n38420, n38421, n38422, n38423,
    n38424, n38425, n38426, n38427, n38428, n38429,
    n38430, n38431, n38432, n38433, n38434, n38435,
    n38436, n38437, n38438, n38439, n38440, n38441,
    n38442, n38443, n38444, n38445, n38446, n38447,
    n38448, n38449, n38450, n38451, n38452, n38453,
    n38454, n38455, n38456, n38457, n38458, n38459,
    n38460, n38461, n38462, n38463, n38464, n38465,
    n38466, n38467, n38468, n38469, n38470, n38471,
    n38472, n38473, n38474, n38475, n38476, n38477,
    n38478, n38479, n38480, n38481, n38482, n38483,
    n38484, n38485, n38486, n38487, n38488, n38489,
    n38490, n38491, n38492, n38493, n38494, n38495,
    n38496, n38497, n38498, n38499, n38500, n38501,
    n38502, n38503, n38504, n38505, n38506, n38507,
    n38508, n38509, n38510, n38511, n38512, n38513,
    n38514, n38515, n38516, n38517, n38518, n38519,
    n38520, n38521, n38522, n38523, n38524, n38525,
    n38526, n38527, n38528, n38529, n38530, n38531,
    n38532, n38533, n38534, n38535, n38536, n38537,
    n38538, n38539, n38540, n38541, n38542, n38543,
    n38544, n38545, n38546, n38547, n38548, n38549,
    n38550, n38551, n38552, n38553, n38554, n38555,
    n38556, n38557, n38558, n38559, n38560, n38561,
    n38562, n38563, n38564, n38565, n38566, n38567,
    n38568, n38569, n38570, n38571, n38572, n38573,
    n38574, n38575, n38576, n38577, n38578, n38579,
    n38580, n38581, n38582, n38583, n38584, n38585,
    n38586, n38587, n38588, n38589, n38590, n38591,
    n38592, n38593, n38594, n38595, n38596, n38597,
    n38598, n38599, n38600, n38601, n38602, n38603,
    n38604, n38605, n38606, n38607, n38608, n38609,
    n38610, n38611, n38612, n38613, n38614, n38615,
    n38616, n38617, n38618, n38619, n38620, n38621,
    n38622, n38623, n38624, n38625, n38626, n38627,
    n38628, n38629, n38630, n38631, n38632, n38633,
    n38634, n38635, n38636, n38637, n38638, n38639,
    n38640, n38641, n38642, n38643, n38644, n38645,
    n38646, n38647, n38648, n38649, n38650, n38651,
    n38652, n38653, n38654, n38655, n38656, n38657,
    n38658, n38659, n38660, n38661, n38662, n38663,
    n38664, n38665, n38666, n38667, n38668, n38669,
    n38670, n38671, n38672, n38673, n38674, n38675,
    n38676, n38677, n38678, n38679, n38680, n38681,
    n38682, n38683, n38684, n38685, n38686, n38687,
    n38688, n38689, n38690, n38691, n38692, n38693,
    n38694, n38695, n38696, n38697, n38698, n38699,
    n38700, n38701, n38702, n38703, n38704, n38705,
    n38706, n38707, n38708, n38709, n38710, n38711,
    n38712, n38713, n38714, n38715, n38716, n38717,
    n38718, n38719, n38720, n38721, n38722, n38723,
    n38724, n38725, n38726, n38727, n38728, n38729,
    n38730, n38731, n38732, n38733, n38734, n38735,
    n38736, n38737, n38738, n38739, n38740, n38741,
    n38742, n38743, n38744, n38745, n38746, n38747,
    n38748, n38749, n38750, n38751, n38752, n38753,
    n38754, n38755, n38756, n38757, n38758, n38759,
    n38760, n38761, n38762, n38763, n38764, n38765,
    n38766, n38767, n38768, n38769, n38770, n38771,
    n38772, n38773, n38774, n38775, n38776, n38777,
    n38778, n38779, n38780, n38781, n38782, n38783,
    n38784, n38785, n38786, n38787, n38788, n38789,
    n38790, n38791, n38792, n38793, n38794, n38795,
    n38796, n38797, n38798, n38799, n38800, n38801,
    n38802, n38803, n38804, n38805, n38806, n38807,
    n38808, n38809, n38810, n38811, n38812, n38813,
    n38814, n38815, n38816, n38817, n38818, n38819,
    n38820, n38821, n38822, n38823, n38824, n38825,
    n38826, n38827, n38828, n38829, n38830, n38831,
    n38832, n38833, n38834, n38835, n38836, n38837,
    n38838, n38839, n38840, n38841, n38842, n38843,
    n38844, n38845, n38846, n38847, n38848, n38849,
    n38850, n38851, n38852, n38853, n38854, n38855,
    n38856, n38857, n38858, n38859, n38860, n38861,
    n38862, n38863, n38864, n38865, n38866, n38867,
    n38868, n38869, n38870, n38871, n38872, n38873,
    n38874, n38875, n38876, n38877, n38878, n38879,
    n38880, n38881, n38882, n38883, n38884, n38885,
    n38886, n38887, n38888, n38889, n38890, n38891,
    n38892, n38893, n38894, n38895, n38896, n38898,
    n38899, n38900, n38901, n38902, n38903, n38904,
    n38905, n38906, n38907, n38908, n38909, n38910,
    n38911, n38912, n38913, n38914, n38915, n38916,
    n38918, n38919, n38920, n38921, n38922, n38923,
    n38924, n38925, n38926, n38927, n38928, n38929,
    n38930, n38931, n38932, n38933, n38934, n38935,
    n38936, n38937, n38938, n38939, n38940, n38941,
    n38942, n38943, n38944, n38945, n38946, n38947,
    n38948, n38949, n38950, n38951, n38952, n38953,
    n38954, n38955, n38956, n38957, n38958, n38959,
    n38960, n38961, n38962, n38963, n38964, n38965,
    n38966, n38967, n38968, n38969, n38970, n38971,
    n38972, n38973, n38974, n38975, n38976, n38977,
    n38978, n38979, n38980, n38981, n38982, n38983,
    n38984, n38985, n38986, n38987, n38988, n38989,
    n38990, n38991, n38992, n38993, n38994, n38995,
    n38996, n38997, n38998, n38999, n39000, n39001,
    n39002, n39003, n39004, n39005, n39006, n39007,
    n39008, n39009, n39010, n39011, n39012, n39013,
    n39014, n39015, n39016, n39017, n39018, n39019,
    n39020, n39021, n39022, n39023, n39024, n39025,
    n39026, n39027, n39028, n39029, n39030, n39031,
    n39032, n39033, n39034, n39035, n39036, n39037,
    n39038, n39039, n39040, n39041, n39042, n39043,
    n39044, n39045, n39046, n39047, n39048, n39049,
    n39050, n39051, n39052, n39053, n39054, n39055,
    n39056, n39057, n39058, n39059, n39060, n39061,
    n39062, n39063, n39064, n39065, n39066, n39067,
    n39068, n39069, n39070, n39071, n39072, n39073,
    n39074, n39075, n39076, n39077, n39078, n39079,
    n39080, n39081, n39082, n39083, n39084, n39085,
    n39086, n39087, n39088, n39089, n39090, n39091,
    n39092, n39093, n39094, n39095, n39096, n39097,
    n39098, n39099, n39100, n39101, n39102, n39103,
    n39104, n39105, n39106, n39107, n39108, n39109,
    n39110, n39111, n39112, n39113, n39114, n39115,
    n39116, n39117, n39118, n39119, n39120, n39121,
    n39122, n39123, n39124, n39125, n39126, n39127,
    n39128, n39129, n39130, n39131, n39132, n39133,
    n39134, n39135, n39136, n39137, n39138, n39139,
    n39140, n39141, n39142, n39143, n39144, n39145,
    n39146, n39147, n39148, n39149, n39150, n39151,
    n39152, n39153, n39154, n39155, n39156, n39157,
    n39158, n39159, n39160, n39161, n39162, n39163,
    n39164, n39165, n39166, n39167, n39168, n39169,
    n39170, n39171, n39172, n39173, n39174, n39175,
    n39176, n39177, n39178, n39179, n39180, n39181,
    n39182, n39183, n39184, n39185, n39186, n39187,
    n39188, n39189, n39190, n39191, n39192, n39193,
    n39194, n39195, n39196, n39197, n39198, n39199,
    n39200, n39201, n39202, n39203, n39204, n39205,
    n39206, n39207, n39208, n39209, n39210, n39211,
    n39212, n39213, n39214, n39215, n39216, n39217,
    n39218, n39219, n39220, n39221, n39222, n39223,
    n39224, n39225, n39226, n39227, n39228, n39229,
    n39230, n39231, n39232, n39233, n39234, n39235,
    n39236, n39237, n39238, n39239, n39240, n39241,
    n39242, n39243, n39244, n39245, n39246, n39247,
    n39248, n39249, n39250, n39251, n39252, n39253,
    n39254, n39255, n39256, n39257, n39258, n39259,
    n39260, n39261, n39262, n39263, n39264, n39265,
    n39266, n39267, n39268, n39269, n39270, n39271,
    n39272, n39273, n39274, n39275, n39276, n39277,
    n39278, n39279, n39280, n39281, n39282, n39283,
    n39284, n39285, n39286, n39287, n39288, n39289,
    n39290, n39291, n39292, n39293, n39294, n39295,
    n39296, n39297, n39298, n39299, n39300, n39301,
    n39302, n39303, n39304, n39305, n39306, n39307,
    n39308, n39309, n39310, n39311, n39312, n39313,
    n39314, n39315, n39316, n39317, n39318, n39319,
    n39320, n39321, n39322, n39323, n39324, n39325,
    n39326, n39327, n39328, n39329, n39330, n39331,
    n39332, n39333, n39334, n39335, n39336, n39337,
    n39338, n39339, n39340, n39341, n39342, n39343,
    n39344, n39345, n39346, n39347, n39348, n39349,
    n39350, n39351, n39352, n39353, n39354, n39355,
    n39356, n39357, n39358, n39359, n39360, n39361,
    n39362, n39363, n39364, n39365, n39366, n39367,
    n39368, n39369, n39370, n39371, n39372, n39373,
    n39374, n39375, n39376, n39377, n39378, n39379,
    n39380, n39381, n39382, n39383, n39384, n39385,
    n39386, n39387, n39388, n39389, n39390, n39391,
    n39392, n39393, n39394, n39395, n39396, n39397,
    n39398, n39399, n39400, n39401, n39402, n39403,
    n39404, n39405, n39406, n39407, n39408, n39409,
    n39410, n39411, n39412, n39413, n39414, n39415,
    n39416, n39417, n39418, n39419, n39420, n39421,
    n39422, n39423, n39424, n39425, n39426, n39427,
    n39428, n39429, n39430, n39431, n39432, n39433,
    n39434, n39435, n39436, n39437, n39438, n39439,
    n39440, n39441, n39442, n39443, n39444, n39445,
    n39446, n39447, n39448, n39449, n39450, n39451,
    n39452, n39453, n39454, n39455, n39456, n39457,
    n39458, n39459, n39460, n39461, n39462, n39463,
    n39464, n39465, n39466, n39467, n39468, n39469,
    n39470, n39471, n39472, n39473, n39474, n39475,
    n39476, n39477, n39478, n39479, n39480, n39481,
    n39482, n39483, n39484, n39485, n39486, n39487,
    n39488, n39489, n39490, n39491, n39492, n39493,
    n39494, n39495, n39496, n39497, n39498, n39499,
    n39500, n39501, n39502, n39503, n39504, n39505,
    n39506, n39507, n39508, n39509, n39510, n39511,
    n39512, n39513, n39514, n39515, n39516, n39517,
    n39518, n39519, n39520, n39521, n39522, n39523,
    n39524, n39525, n39526, n39527, n39528, n39529,
    n39530, n39531, n39532, n39533, n39534, n39535,
    n39536, n39537, n39538, n39539, n39540, n39541,
    n39542, n39543, n39544, n39545, n39546, n39547,
    n39548, n39549, n39550, n39551, n39552, n39553,
    n39554, n39555, n39556, n39557, n39558, n39559,
    n39560, n39561, n39562, n39563, n39564, n39565,
    n39566, n39567, n39568, n39569, n39570, n39571,
    n39572, n39573, n39574, n39575, n39576, n39577,
    n39578, n39579, n39580, n39581, n39582, n39583,
    n39584, n39585, n39586, n39587, n39588, n39589,
    n39590, n39591, n39592, n39593, n39594, n39595,
    n39596, n39597, n39598, n39599, n39600, n39601,
    n39602, n39603, n39604, n39605, n39606, n39607,
    n39608, n39609, n39610, n39611, n39612, n39613,
    n39614, n39615, n39616, n39617, n39618, n39619,
    n39620, n39621, n39622, n39623, n39624, n39625,
    n39626, n39627, n39628, n39629, n39630, n39631,
    n39632, n39633, n39634, n39635, n39636, n39637,
    n39638, n39639, n39640, n39641, n39642, n39643,
    n39644, n39645, n39646, n39647, n39648, n39649,
    n39650, n39651, n39652, n39653, n39654, n39655,
    n39656, n39657, n39658, n39659, n39660, n39661,
    n39662, n39663, n39664, n39665, n39666, n39667,
    n39668, n39669, n39670, n39671, n39672, n39673,
    n39674, n39675, n39676, n39677, n39678, n39679,
    n39680, n39681, n39682, n39683, n39684, n39685,
    n39686, n39687, n39688, n39689, n39690, n39691,
    n39692, n39693, n39694, n39695, n39696, n39697,
    n39698, n39699, n39700, n39701, n39702, n39703,
    n39704, n39705, n39706, n39707, n39708, n39709,
    n39710, n39711, n39712, n39713, n39714, n39715,
    n39716, n39717, n39718, n39719, n39720, n39721,
    n39722, n39723, n39724, n39725, n39726, n39727,
    n39728, n39729, n39730, n39731, n39732, n39733,
    n39734, n39735, n39736, n39737, n39738, n39739,
    n39740, n39741, n39742, n39743, n39744, n39745,
    n39746, n39747, n39748, n39749, n39750, n39751,
    n39752, n39753, n39754, n39755, n39756, n39757,
    n39758, n39759, n39760, n39761, n39762, n39763,
    n39764, n39765, n39766, n39767, n39768, n39769,
    n39770, n39771, n39772, n39773, n39774, n39775,
    n39776, n39777, n39778, n39779, n39780, n39781,
    n39782, n39783, n39784, n39785, n39786, n39787,
    n39788, n39789, n39790, n39791, n39792, n39793,
    n39794, n39795, n39796, n39797, n39798, n39799,
    n39800, n39801, n39802, n39803, n39804, n39805,
    n39806, n39807, n39808, n39809, n39810, n39811,
    n39812, n39813, n39814, n39815, n39816, n39817,
    n39818, n39819, n39820, n39821, n39822, n39823,
    n39824, n39825, n39826, n39827, n39828, n39829,
    n39830, n39831, n39832, n39833, n39834, n39835,
    n39836, n39837, n39838, n39839, n39840, n39841,
    n39842, n39843, n39844, n39845, n39846, n39847,
    n39848, n39849, n39850, n39851, n39852, n39853,
    n39854, n39855, n39856, n39857, n39858, n39859,
    n39860, n39861, n39862, n39863, n39864, n39865,
    n39866, n39867, n39868, n39869, n39870, n39871,
    n39872, n39873, n39874, n39875, n39876, n39877,
    n39878, n39879, n39880, n39881, n39882, n39883,
    n39884, n39885, n39886, n39887, n39888, n39889,
    n39890, n39891, n39892, n39893, n39894, n39895,
    n39896, n39897, n39898, n39899, n39900, n39901,
    n39902, n39903, n39904, n39905, n39906, n39907,
    n39908, n39909, n39910, n39911, n39912, n39913,
    n39914, n39915, n39916, n39917, n39918, n39919,
    n39920, n39921, n39922, n39923, n39924, n39925,
    n39926, n39927, n39928, n39929, n39930, n39931,
    n39932, n39933, n39934, n39935, n39936, n39937,
    n39938, n39939, n39940, n39941, n39942, n39943,
    n39944, n39945, n39946, n39947, n39948, n39949,
    n39950, n39951, n39952, n39953, n39954, n39955,
    n39956, n39957, n39958, n39959, n39960, n39961,
    n39962, n39963, n39964, n39965, n39966, n39967,
    n39968, n39969, n39970, n39971, n39972, n39973,
    n39974, n39975, n39976, n39977, n39978, n39979,
    n39980, n39981, n39982, n39983, n39984, n39985,
    n39986, n39987, n39988, n39989, n39990, n39991,
    n39992, n39993, n39994, n39995, n39996, n39997,
    n39998, n39999, n40000, n40001, n40002, n40003,
    n40004, n40005, n40006, n40007, n40008, n40009,
    n40010, n40011, n40012, n40013, n40014, n40015,
    n40016, n40017, n40018, n40019, n40020, n40021,
    n40022, n40023, n40024, n40025, n40026, n40027,
    n40028, n40029, n40030, n40031, n40032, n40033,
    n40034, n40035, n40036, n40037, n40038, n40039,
    n40040, n40041, n40042, n40043, n40044, n40045,
    n40046, n40047, n40048, n40049, n40050, n40051,
    n40052, n40053, n40054, n40055, n40056, n40057,
    n40058, n40059, n40060, n40061, n40062, n40063,
    n40064, n40065, n40066, n40067, n40068, n40069,
    n40070, n40071, n40072, n40073, n40074, n40075,
    n40076, n40077, n40078, n40079, n40080, n40081,
    n40082, n40083, n40084, n40085, n40086, n40087,
    n40088, n40089, n40090, n40091, n40092, n40093,
    n40094, n40095, n40096, n40097, n40098, n40099,
    n40100, n40101, n40102, n40103, n40104, n40105,
    n40106, n40107, n40108, n40109, n40110, n40111,
    n40112, n40113, n40114, n40115, n40116, n40117,
    n40118, n40119, n40120, n40121, n40122, n40123,
    n40124, n40125, n40126, n40127, n40128, n40129,
    n40130, n40131, n40132, n40133, n40134, n40135,
    n40136, n40137, n40138, n40139, n40140, n40141,
    n40142, n40143, n40144, n40145, n40146, n40147,
    n40148, n40149, n40150, n40151, n40152, n40153,
    n40154, n40155, n40156, n40157, n40158, n40159,
    n40160, n40161, n40162, n40163, n40164, n40165,
    n40166, n40167, n40168, n40169, n40170, n40171,
    n40172, n40173, n40174, n40175, n40176, n40177,
    n40178, n40179, n40180, n40181, n40182, n40183,
    n40184, n40185, n40186, n40187, n40188, n40189,
    n40190, n40191, n40192, n40193, n40194, n40195,
    n40196, n40197, n40198, n40199, n40200, n40201,
    n40202, n40203, n40204, n40205, n40206, n40207,
    n40208, n40209, n40210, n40211, n40212, n40213,
    n40214, n40215, n40216, n40217, n40218, n40219,
    n40220, n40221, n40222, n40223, n40224, n40225,
    n40226, n40227, n40228, n40229, n40230, n40231,
    n40232, n40233, n40234, n40235, n40236, n40237,
    n40238, n40239, n40240, n40241, n40242, n40243,
    n40244, n40245, n40246, n40247, n40248, n40249,
    n40250, n40251, n40252, n40253, n40254, n40255,
    n40256, n40257, n40258, n40259, n40260, n40261,
    n40262, n40263, n40264, n40265, n40266, n40267,
    n40268, n40269, n40270, n40271, n40272, n40273,
    n40274, n40275, n40276, n40277, n40278, n40279,
    n40280, n40281, n40282, n40283, n40284, n40285,
    n40286, n40287, n40288, n40289, n40290, n40291,
    n40292, n40293, n40294, n40295, n40296, n40297,
    n40298, n40299, n40300, n40301, n40302, n40303,
    n40304, n40305, n40306, n40307, n40309, n40310,
    n40311, n40312, n40313, n40314, n40315, n40316,
    n40317, n40318, n40319, n40320, n40321, n40322,
    n40323, n40324, n40325, n40326, n40327, n40328,
    n40329, n40330, n40331, n40332, n40333, n40334,
    n40335, n40336, n40337, n40338, n40339, n40340,
    n40341, n40342, n40343, n40344, n40345, n40346,
    n40347, n40348, n40349, n40350, n40351, n40352,
    n40353, n40354, n40355, n40356, n40357, n40358,
    n40359, n40360, n40361, n40362, n40363, n40364,
    n40365, n40366, n40367, n40368, n40369, n40370,
    n40371, n40372, n40373, n40374, n40375, n40376,
    n40377, n40378, n40379, n40380, n40381, n40382,
    n40383, n40384, n40385, n40386, n40387, n40388,
    n40389, n40390, n40391, n40392, n40393, n40394,
    n40395, n40396, n40397, n40398, n40399, n40400,
    n40401, n40402, n40403, n40404, n40405, n40406,
    n40407, n40408, n40409, n40410, n40411, n40412,
    n40413, n40414, n40415, n40416, n40417, n40418,
    n40419, n40420, n40421, n40422, n40423, n40424,
    n40425, n40426, n40427, n40428, n40429, n40430,
    n40431, n40432, n40433, n40434, n40435, n40436,
    n40437, n40438, n40439, n40440, n40441, n40442,
    n40443, n40444, n40445, n40446, n40447, n40448,
    n40449, n40450, n40451, n40452, n40453, n40454,
    n40455, n40456, n40457, n40458, n40459, n40460,
    n40461, n40462, n40463, n40464, n40465, n40466,
    n40467, n40468, n40469, n40470, n40471, n40472,
    n40473, n40474, n40475, n40476, n40477, n40478,
    n40479, n40480, n40481, n40482, n40483, n40484,
    n40485, n40486, n40487, n40488, n40489, n40490,
    n40491, n40492, n40493, n40494, n40495, n40496,
    n40497, n40498, n40499, n40500, n40501, n40502,
    n40503, n40504, n40505, n40506, n40507, n40508,
    n40509, n40510, n40511, n40512, n40513, n40514,
    n40515, n40516, n40517, n40518, n40519, n40520,
    n40521, n40522, n40523, n40524, n40525, n40526,
    n40527, n40528, n40529, n40530, n40531, n40532,
    n40533, n40534, n40535, n40536, n40537, n40538,
    n40539, n40540, n40541, n40542, n40543, n40544,
    n40545, n40546, n40547, n40548, n40549, n40550,
    n40551, n40552, n40553, n40554, n40555, n40556,
    n40557, n40558, n40559, n40560, n40561, n40562,
    n40563, n40564, n40565, n40566, n40567, n40568,
    n40569, n40570, n40571, n40572, n40573, n40574,
    n40575, n40576, n40577, n40578, n40579, n40580,
    n40581, n40582, n40583, n40584, n40585, n40586,
    n40587, n40588, n40589, n40590, n40591, n40592,
    n40593, n40594, n40595, n40596, n40597, n40598,
    n40599, n40600, n40601, n40602, n40603, n40604,
    n40605, n40606, n40607, n40608, n40609, n40610,
    n40611, n40612, n40613, n40614, n40615, n40616,
    n40617, n40618, n40619, n40620, n40621, n40622,
    n40623, n40624, n40625, n40626, n40627, n40628,
    n40629, n40630, n40631, n40632, n40633, n40634,
    n40635, n40636, n40637, n40638, n40639, n40640,
    n40641, n40642, n40643, n40644, n40645, n40646,
    n40647, n40648, n40649, n40650, n40651, n40652,
    n40653, n40654, n40655, n40656, n40657, n40658,
    n40659, n40660, n40661, n40662, n40663, n40664,
    n40665, n40666, n40667, n40668, n40669, n40670,
    n40671, n40672, n40673, n40674, n40675, n40676,
    n40677, n40678, n40679, n40680, n40681, n40682,
    n40683, n40684, n40685, n40686, n40687, n40688,
    n40689, n40690, n40691, n40692, n40693, n40694,
    n40695, n40696, n40697, n40698, n40699, n40700,
    n40701, n40702, n40703, n40704, n40705, n40706,
    n40707, n40708, n40709, n40710, n40711, n40712,
    n40713, n40714, n40715, n40717, n40718, n40719,
    n40720, n40721, n40722, n40723, n40724, n40725,
    n40726, n40727, n40728, n40729, n40730, n40731,
    n40732, n40733, n40734, n40735, n40736, n40738,
    n40739, n40740, n40741, n40742, n40743, n40744,
    n40745, n40746, n40747, n40748, n40749, n40750,
    n40751, n40752, n40753, n40754, n40755, n40756,
    n40757, n40758, n40759, n40760, n40761, n40762,
    n40763, n40764, n40765, n40766, n40767, n40768,
    n40769, n40770, n40771, n40772, n40773, n40774,
    n40775, n40777, n40778, n40779, n40780, n40781,
    n40782, n40783, n40784, n40785, n40786, n40787,
    n40788, n40789, n40790, n40791, n40792, n40793,
    n40794, n40795, n40796, n40797, n40798, n40799,
    n40800, n40801, n40802, n40803, n40804, n40805,
    n40806, n40807, n40808, n40809, n40810, n40811,
    n40812, n40813, n40814, n40815, n40816, n40817,
    n40818, n40819, n40820, n40821, n40822, n40823,
    n40824, n40825, n40826, n40827, n40828, n40829,
    n40830, n40831, n40832, n40833, n40834, n40835,
    n40836, n40837, n40838, n40839, n40840, n40841,
    n40842, n40843, n40844, n40845, n40846, n40847,
    n40848, n40849, n40850, n40851, n40852, n40853,
    n40854, n40855, n40856, n40857, n40858, n40859,
    n40860, n40861, n40862, n40863, n40864, n40865,
    n40866, n40867, n40868, n40869, n40870, n40871,
    n40872, n40873, n40874, n40875, n40876, n40877,
    n40878, n40879, n40880, n40881, n40882, n40883,
    n40884, n40885, n40886, n40887, n40888, n40889,
    n40890, n40891, n40892, n40893, n40894, n40895,
    n40896, n40897, n40898, n40899, n40900, n40901,
    n40902, n40903, n40904, n40905, n40906, n40907,
    n40908, n40909, n40910, n40911, n40912, n40913,
    n40915, n40916, n40917, n40918, n40919, n40920,
    n40921, n40922, n40923, n40924, n40925, n40926,
    n40927, n40928, n40929, n40930, n40931, n40932,
    n40933, n40934, n40935, n40936, n40937, n40938,
    n40939, n40940, n40941, n40942, n40943, n40944,
    n40945, n40946, n40947, n40948, n40949, n40950,
    n40951, n40952, n40953, n40954, n40955, n40956,
    n40957, n40958, n40959, n40960, n40961, n40962,
    n40963, n40964, n40965, n40966, n40967, n40968,
    n40969, n40970, n40971, n40972, n40973, n40974,
    n40975, n40976, n40977, n40978, n40979, n40980,
    n40981, n40982, n40983, n40984, n40985, n40986,
    n40987, n40988, n40989, n40990, n40991, n40992,
    n40993, n40994, n40995, n40996, n40997, n40998,
    n40999, n41000, n41001, n41002, n41003, n41004,
    n41005, n41006, n41007, n41008, n41009, n41010,
    n41011, n41012, n41013, n41014, n41015, n41016,
    n41017, n41018, n41019, n41020, n41021, n41022,
    n41023, n41024, n41025, n41026, n41027, n41028,
    n41029, n41030, n41031, n41032, n41033, n41034,
    n41035, n41036, n41037, n41038, n41039, n41040,
    n41041, n41042, n41043, n41044, n41045, n41046,
    n41047, n41048, n41049, n41050, n41051, n41052,
    n41053, n41054, n41055, n41056, n41057, n41058,
    n41059, n41060, n41061, n41062, n41063, n41064,
    n41065, n41066, n41067, n41068, n41069, n41070,
    n41071, n41072, n41073, n41074, n41075, n41076,
    n41077, n41078, n41079, n41080, n41081, n41082,
    n41083, n41084, n41085, n41086, n41087, n41088,
    n41089, n41090, n41091, n41092, n41093, n41094,
    n41095, n41096, n41097, n41098, n41099, n41100,
    n41101, n41102, n41103, n41104, n41105, n41106,
    n41107, n41108, n41109, n41110, n41111, n41112,
    n41113, n41114, n41115, n41116, n41117, n41118,
    n41119, n41120, n41121, n41122, n41123, n41124,
    n41125, n41126, n41127, n41128, n41129, n41130,
    n41131, n41132, n41133, n41134, n41135, n41136,
    n41137, n41138, n41139, n41140, n41141, n41142,
    n41143, n41144, n41145, n41146, n41147, n41148,
    n41149, n41150, n41151, n41152, n41153, n41154,
    n41155, n41156, n41157, n41158, n41159, n41160,
    n41161, n41162, n41163, n41164, n41165, n41166,
    n41167, n41168, n41169, n41170, n41171, n41172,
    n41173, n41174, n41175, n41176, n41177, n41178,
    n41179, n41180, n41181, n41182, n41183, n41184,
    n41185, n41186, n41187, n41188, n41189, n41190,
    n41191, n41192, n41193, n41194, n41195, n41196,
    n41197, n41198, n41199, n41200, n41201, n41202,
    n41203, n41204, n41205, n41206, n41207, n41208,
    n41209, n41210, n41211, n41212, n41213, n41214,
    n41215, n41216, n41217, n41218, n41219, n41220,
    n41221, n41222, n41223, n41224, n41225, n41226,
    n41227, n41228, n41229, n41230, n41231, n41232,
    n41233, n41234, n41235, n41236, n41237, n41238,
    n41239, n41240, n41241, n41242, n41243, n41244,
    n41245, n41246, n41247, n41248, n41249, n41250,
    n41251, n41252, n41253, n41254, n41255, n41256,
    n41257, n41258, n41259, n41260, n41261, n41262,
    n41263, n41264, n41265, n41266, n41267, n41268,
    n41269, n41270, n41271, n41272, n41273, n41274,
    n41275, n41276, n41277, n41278, n41279, n41280,
    n41281, n41282, n41283, n41284, n41285, n41286,
    n41287, n41288, n41289, n41290, n41291, n41292,
    n41293, n41294, n41295, n41296, n41297, n41298,
    n41299, n41300, n41301, n41302, n41303, n41304,
    n41305, n41306, n41307, n41308, n41309, n41310,
    n41311, n41312, n41313, n41314, n41315, n41316,
    n41317, n41318, n41319, n41320, n41321, n41322,
    n41323, n41324, n41325, n41326, n41327, n41328,
    n41329, n41330, n41331, n41332, n41333, n41334,
    n41335, n41336, n41337, n41338, n41339, n41340,
    n41341, n41342, n41343, n41344, n41345, n41346,
    n41347, n41348, n41349, n41350, n41351, n41352,
    n41353, n41354, n41355, n41356, n41357, n41358,
    n41359, n41360, n41361, n41362, n41363, n41364,
    n41365, n41366, n41367, n41368, n41369, n41370,
    n41371, n41372, n41373, n41374, n41375, n41376,
    n41377, n41378, n41379, n41380, n41381, n41382,
    n41383, n41384, n41385, n41386, n41387, n41388,
    n41389, n41390, n41391, n41392, n41393, n41394,
    n41395, n41396, n41397, n41398, n41399, n41400,
    n41401, n41402, n41403, n41404, n41405, n41406,
    n41407, n41408, n41409, n41410, n41411, n41412,
    n41413, n41414, n41415, n41416, n41417, n41418,
    n41419, n41420, n41421, n41422, n41423, n41424,
    n41425, n41426, n41427, n41428, n41429, n41430,
    n41431, n41432, n41433, n41434, n41435, n41436,
    n41437, n41438, n41439, n41440, n41441, n41442,
    n41443, n41444, n41445, n41446, n41447, n41448,
    n41449, n41450, n41451, n41452, n41453, n41454,
    n41455, n41456, n41457, n41458, n41459, n41460,
    n41461, n41462, n41463, n41464, n41465, n41466,
    n41467, n41468, n41469, n41470, n41471, n41472,
    n41473, n41474, n41475, n41476, n41477, n41478,
    n41479, n41480, n41481, n41482, n41483, n41484,
    n41485, n41486, n41487, n41488, n41489, n41490,
    n41491, n41492, n41493, n41494, n41495, n41496,
    n41497, n41498, n41499, n41500, n41501, n41502,
    n41503, n41504, n41505, n41506, n41507, n41508,
    n41509, n41510, n41511, n41512, n41513, n41514,
    n41515, n41516, n41517, n41518, n41519, n41520,
    n41521, n41522, n41523, n41524, n41525, n41526,
    n41527, n41528, n41529, n41530, n41531, n41532,
    n41533, n41534, n41535, n41536, n41537, n41538,
    n41539, n41540, n41541, n41542, n41543, n41544,
    n41545, n41546, n41547, n41548, n41549, n41550,
    n41551, n41552, n41553, n41554, n41555, n41556,
    n41557, n41558, n41559, n41560, n41561, n41562,
    n41563, n41564, n41565, n41566, n41567, n41568,
    n41569, n41570, n41571, n41572, n41573, n41574,
    n41575, n41576, n41577, n41578, n41579, n41580,
    n41581, n41582, n41583, n41584, n41585, n41586,
    n41587, n41588, n41589, n41590, n41591, n41592,
    n41593, n41594, n41595, n41596, n41597, n41598,
    n41599, n41600, n41601, n41602, n41603, n41604,
    n41605, n41606, n41607, n41608, n41609, n41610,
    n41611, n41612, n41613, n41614, n41615, n41616,
    n41617, n41618, n41619, n41620, n41621, n41622,
    n41623, n41624, n41625, n41626, n41627, n41628,
    n41629, n41630, n41631, n41632, n41633, n41634,
    n41635, n41636, n41637, n41638, n41639, n41640,
    n41641, n41642, n41643, n41644, n41645, n41646,
    n41647, n41648, n41649, n41650, n41651, n41652,
    n41653, n41654, n41655, n41656, n41657, n41658,
    n41659, n41660, n41661, n41662, n41663, n41664,
    n41665, n41666, n41667, n41668, n41669, n41670,
    n41671, n41672, n41673, n41674, n41675, n41676,
    n41677, n41678, n41679, n41680, n41681, n41682,
    n41683, n41684, n41685, n41686, n41687, n41688,
    n41689, n41690, n41691, n41692, n41693, n41694,
    n41695, n41696, n41697, n41698, n41699, n41700,
    n41701, n41702, n41703, n41704, n41705, n41706,
    n41707, n41708, n41709, n41710, n41711, n41712,
    n41713, n41714, n41715, n41716, n41717, n41718,
    n41719, n41720, n41721, n41722, n41723, n41724,
    n41725, n41726, n41727, n41728, n41729, n41730,
    n41731, n41732, n41733, n41734, n41735, n41736,
    n41737, n41738, n41739, n41740, n41741, n41742,
    n41743, n41744, n41745, n41746, n41747, n41748,
    n41749, n41750, n41751, n41752, n41753, n41754,
    n41755, n41756, n41757, n41758, n41759, n41760,
    n41761, n41762, n41763, n41764, n41765, n41766,
    n41767, n41768, n41769, n41770, n41771, n41772,
    n41773, n41774, n41775, n41776, n41777, n41778,
    n41779, n41780, n41781, n41782, n41783, n41784,
    n41785, n41786, n41787, n41788, n41789, n41790,
    n41791, n41792, n41793, n41794, n41795, n41796,
    n41797, n41798, n41799, n41800, n41801, n41802,
    n41803, n41804, n41805, n41806, n41807, n41808,
    n41809, n41810, n41811, n41812, n41813, n41814,
    n41815, n41816, n41817, n41818, n41819, n41820,
    n41821, n41822, n41823, n41824, n41825, n41826,
    n41827, n41828, n41829, n41830, n41831, n41832,
    n41833, n41834, n41835, n41836, n41837, n41838,
    n41839, n41840, n41841, n41842, n41843, n41844,
    n41845, n41846, n41847, n41848, n41849, n41850,
    n41851, n41852, n41853, n41854, n41855, n41856,
    n41857, n41858, n41859, n41860, n41861, n41862,
    n41863, n41864, n41865, n41866, n41867, n41868,
    n41869, n41870, n41871, n41872, n41873, n41874,
    n41875, n41876, n41877, n41878, n41879, n41880,
    n41881, n41882, n41883, n41884, n41885, n41886,
    n41887, n41888, n41889, n41890, n41891, n41892,
    n41893, n41894, n41895, n41896, n41897, n41898,
    n41899, n41900, n41901, n41902, n41903, n41904,
    n41905, n41906, n41907, n41908, n41909, n41910,
    n41911, n41912, n41913, n41914, n41915, n41916,
    n41917, n41918, n41919, n41920, n41921, n41922,
    n41923, n41924, n41925, n41926, n41927, n41928,
    n41929, n41930, n41931, n41932, n41933, n41934,
    n41935, n41936, n41937, n41938, n41939, n41940,
    n41941, n41942, n41943, n41944, n41945, n41946,
    n41947, n41948, n41949, n41950, n41951, n41952,
    n41953, n41954, n41955, n41956, n41957, n41958,
    n41959, n41960, n41961, n41962, n41963, n41964,
    n41965, n41966, n41967, n41968, n41969, n41970,
    n41971, n41972, n41973, n41974, n41975, n41976,
    n41977, n41978, n41979, n41980, n41981, n41982,
    n41983, n41984, n41985, n41986, n41987, n41988,
    n41989, n41990, n41991, n41992, n41993, n41994,
    n41995, n41996, n41997, n41998, n41999, n42000,
    n42001, n42002, n42003, n42004, n42005, n42006,
    n42007, n42008, n42009, n42010, n42011, n42012,
    n42013, n42014, n42015, n42016, n42017, n42018,
    n42019, n42020, n42021, n42022, n42023, n42024,
    n42025, n42026, n42027, n42028, n42029, n42030,
    n42031, n42032, n42033, n42034, n42035, n42036,
    n42037, n42038, n42039, n42040, n42041, n42042,
    n42043, n42044, n42045, n42046, n42047, n42048,
    n42049, n42050, n42051, n42052, n42053, n42054,
    n42055, n42056, n42057, n42058, n42059, n42060,
    n42061, n42062, n42063, n42064, n42065, n42066,
    n42067, n42068, n42069, n42070, n42071, n42072,
    n42073, n42074, n42075, n42076, n42077, n42078,
    n42079, n42080, n42081, n42082, n42083, n42084,
    n42085, n42086, n42087, n42088, n42089, n42090,
    n42091, n42092, n42093, n42094, n42095, n42096,
    n42097, n42098, n42099, n42100, n42101, n42102,
    n42103, n42104, n42105, n42106, n42107, n42108,
    n42109, n42110, n42111, n42112, n42113, n42114,
    n42115, n42116, n42117, n42118, n42119, n42120,
    n42121, n42122, n42123, n42124, n42125, n42126,
    n42127, n42128, n42129, n42130, n42131, n42132,
    n42133, n42134, n42135, n42136, n42137, n42138,
    n42139, n42140, n42141, n42142, n42143, n42144,
    n42145, n42146, n42147, n42148, n42149, n42150,
    n42151, n42152, n42153, n42154, n42155, n42156,
    n42157, n42158, n42159, n42160, n42161, n42162,
    n42163, n42164, n42165, n42166, n42167, n42168,
    n42169, n42170, n42171, n42172, n42173, n42174,
    n42175, n42176, n42177, n42178, n42179, n42180,
    n42181, n42182, n42183, n42184, n42185, n42186,
    n42187, n42188, n42189, n42190, n42191, n42192,
    n42193, n42194, n42195, n42196, n42197, n42198,
    n42199, n42200, n42201, n42202, n42203, n42204,
    n42205, n42206, n42207, n42208, n42209, n42210,
    n42211, n42212, n42213, n42214, n42215, n42216,
    n42217, n42218, n42219, n42220, n42221, n42222,
    n42223, n42224, n42225, n42226, n42227, n42228,
    n42229, n42230, n42231, n42232, n42233, n42234,
    n42235, n42236, n42237, n42238, n42239, n42240,
    n42241, n42242, n42243, n42244, n42245, n42246,
    n42247, n42248, n42249, n42250, n42251, n42252,
    n42253, n42254, n42255, n42256, n42257, n42258,
    n42259, n42260, n42261, n42262, n42263, n42264,
    n42265, n42266, n42267, n42268, n42269, n42270,
    n42271, n42272, n42273, n42274, n42275, n42276,
    n42277, n42278, n42279, n42280, n42281, n42282,
    n42283, n42284, n42285, n42286, n42287, n42288,
    n42289, n42290, n42291, n42292, n42293, n42294,
    n42295, n42296, n42297, n42298, n42299, n42300,
    n42301, n42302, n42303, n42304, n42305, n42306,
    n42307, n42308, n42309, n42310, n42311, n42312,
    n42313, n42314, n42315, n42316, n42317, n42318,
    n42319, n42320, n42321, n42322, n42323, n42324,
    n42325, n42326, n42327, n42328, n42329, n42330,
    n42331, n42332, n42333, n42334, n42335, n42336,
    n42337, n42338, n42339, n42340, n42341, n42342,
    n42343, n42344, n42345, n42346, n42347, n42348,
    n42349, n42350, n42351, n42352, n42353, n42354,
    n42355, n42356, n42357, n42358, n42359, n42360,
    n42361, n42362, n42363, n42364, n42365, n42366,
    n42367, n42368, n42369, n42370, n42371, n42372,
    n42373, n42374, n42375, n42376, n42377, n42378,
    n42379, n42380, n42381, n42382, n42383, n42384,
    n42385, n42386, n42387, n42388, n42389, n42390,
    n42391, n42392, n42393, n42394, n42395, n42396,
    n42397, n42398, n42399, n42400, n42401, n42402,
    n42403, n42404, n42405, n42406, n42407, n42408,
    n42409, n42410, n42411, n42412, n42413, n42414,
    n42415, n42416, n42417, n42418, n42419, n42420,
    n42421, n42422, n42423, n42424, n42425, n42426,
    n42427, n42428, n42429, n42430, n42431, n42432,
    n42433, n42434, n42435, n42436, n42437, n42438,
    n42439, n42440, n42441, n42442, n42443, n42444,
    n42445, n42446, n42447, n42448, n42449, n42450,
    n42451, n42452, n42453, n42454, n42455, n42456,
    n42457, n42458, n42459, n42460, n42461, n42462,
    n42463, n42464, n42465, n42466, n42467, n42468,
    n42469, n42470, n42471, n42472, n42473, n42474,
    n42475, n42476, n42477, n42478, n42479, n42480,
    n42481, n42482, n42483, n42484, n42485, n42486,
    n42487, n42488, n42489, n42490, n42491, n42492,
    n42493, n42494, n42495, n42496, n42497, n42498,
    n42499, n42500, n42501, n42502, n42503, n42504,
    n42505, n42506, n42507, n42508, n42509, n42510,
    n42511, n42512, n42513, n42514, n42515, n42516,
    n42517, n42518, n42519, n42520, n42521, n42522,
    n42523, n42524, n42525, n42526, n42527, n42528,
    n42529, n42530, n42531, n42532, n42533, n42534,
    n42535, n42536, n42537, n42538, n42539, n42540,
    n42541, n42542, n42543, n42544, n42545, n42546,
    n42547, n42548, n42549, n42550, n42551, n42552,
    n42553, n42554, n42555, n42556, n42557, n42558,
    n42559, n42560, n42561, n42562, n42563, n42564,
    n42565, n42566, n42567, n42568, n42569, n42570,
    n42571, n42572, n42573, n42574, n42575, n42576,
    n42577, n42578, n42579, n42580, n42581, n42582,
    n42583, n42584, n42585, n42586, n42587, n42588,
    n42589, n42590, n42591, n42592, n42593, n42594,
    n42595, n42596, n42597, n42598, n42599, n42600,
    n42601, n42602, n42603, n42604, n42605, n42606,
    n42607, n42608, n42609, n42610, n42611, n42612,
    n42613, n42614, n42615, n42616, n42617, n42618,
    n42619, n42620, n42621, n42622, n42623, n42624,
    n42625, n42626, n42627, n42628, n42629, n42630,
    n42631, n42632, n42633, n42634, n42635, n42636,
    n42637, n42638, n42639, n42640, n42641, n42642,
    n42643, n42644, n42645, n42646, n42647, n42648,
    n42649, n42650, n42651, n42652, n42653, n42654,
    n42655, n42656, n42657, n42658, n42659, n42660,
    n42661, n42662, n42663, n42664, n42665, n42666,
    n42667, n42668, n42669, n42670, n42671, n42672,
    n42673, n42674, n42675, n42676, n42677, n42678,
    n42679, n42680, n42681, n42682, n42683, n42684,
    n42685, n42686, n42687, n42688, n42689, n42690,
    n42691, n42692, n42693, n42694, n42695, n42696,
    n42697, n42698, n42699, n42700, n42701, n42702,
    n42703, n42704, n42705, n42706, n42707, n42708,
    n42709, n42710, n42711, n42712, n42713, n42714,
    n42715, n42716, n42717, n42718, n42719, n42720,
    n42721, n42722, n42723, n42724, n42725, n42726,
    n42727, n42728, n42729, n42730, n42731, n42732,
    n42733, n42734, n42735, n42736, n42737, n42738,
    n42739, n42740, n42741, n42742, n42743, n42744,
    n42745, n42746, n42747, n42748, n42749, n42750,
    n42751, n42752, n42753, n42754, n42755, n42756,
    n42757, n42758, n42759, n42760, n42761, n42762,
    n42763, n42764, n42765, n42766, n42767, n42768,
    n42769, n42770, n42771, n42772, n42773, n42774,
    n42775, n42776, n42777, n42778, n42779, n42780,
    n42781, n42782, n42783, n42784, n42785, n42786,
    n42787, n42788, n42789, n42790, n42791, n42792,
    n42793, n42794, n42795, n42796, n42797, n42798,
    n42799, n42800, n42801, n42802, n42803, n42804,
    n42805, n42806, n42807, n42808, n42809, n42810,
    n42811, n42812, n42813, n42814, n42815, n42816,
    n42817, n42818, n42819, n42820, n42821, n42822,
    n42823, n42824, n42825, n42826, n42827, n42828,
    n42829, n42830, n42831, n42832, n42833, n42834,
    n42835, n42836, n42837, n42838, n42839, n42840,
    n42841, n42842, n42843, n42844, n42845, n42846,
    n42847, n42848, n42849, n42850, n42851, n42852,
    n42853, n42854, n42855, n42856, n42857, n42858,
    n42859, n42860, n42861, n42862, n42863, n42864,
    n42865, n42866, n42867, n42868, n42869, n42870,
    n42871, n42872, n42873, n42874, n42875, n42876,
    n42877, n42878, n42879, n42880, n42881, n42882,
    n42883, n42884, n42885, n42886, n42887, n42888,
    n42889, n42890, n42891, n42892, n42893, n42894,
    n42895, n42896, n42897, n42898, n42899, n42900,
    n42901, n42902, n42903, n42904, n42905, n42906,
    n42907, n42908, n42909, n42910, n42911, n42912,
    n42913, n42914, n42915, n42916, n42917, n42918,
    n42919, n42920, n42921, n42922, n42923, n42924,
    n42925, n42926, n42927, n42928, n42929, n42930,
    n42931, n42932, n42933, n42934, n42935, n42936,
    n42937, n42938, n42939, n42940, n42941, n42942,
    n42943, n42944, n42945, n42946, n42947, n42948,
    n42949, n42950, n42951, n42952, n42953, n42954,
    n42955, n42956, n42957, n42958, n42959, n42960,
    n42961, n42962, n42963, n42964, n42965, n42966,
    n42967, n42968, n42969, n42970, n42971, n42973,
    n42974, n42975, n42976, n42977, n42978, n42979,
    n42980, n42981, n42982, n42983, n42984, n42985,
    n42986, n42987, n42988, n42989, n42990, n42991,
    n42992, n42993, n42994, n42995, n42996, n42997,
    n42998, n42999, n43000, n43001, n43002, n43003,
    n43004, n43005, n43006, n43007, n43008, n43009,
    n43010, n43011, n43012, n43013, n43014, n43015,
    n43016, n43017, n43018, n43019, n43020, n43021,
    n43022, n43023, n43024, n43025, n43026, n43027,
    n43028, n43029, n43030, n43031, n43032, n43033,
    n43034, n43035, n43036, n43037, n43038, n43039,
    n43040, n43041, n43042, n43043, n43044, n43045,
    n43046, n43047, n43048, n43049, n43050, n43051,
    n43052, n43053, n43054, n43055, n43056, n43057,
    n43058, n43059, n43060, n43061, n43062, n43063,
    n43064, n43065, n43066, n43067, n43068, n43069,
    n43070, n43071, n43072, n43073, n43074, n43075,
    n43076, n43077, n43078, n43079, n43080, n43081,
    n43082, n43083, n43084, n43085, n43086, n43087,
    n43088, n43089, n43090, n43091, n43092, n43093,
    n43094, n43095, n43096, n43097, n43098, n43099,
    n43100, n43101, n43102, n43103, n43104, n43105,
    n43106, n43107, n43108, n43109, n43110, n43111,
    n43112, n43113, n43114, n43115, n43116, n43117,
    n43118, n43119, n43120, n43121, n43122, n43123,
    n43124, n43125, n43126, n43127, n43128, n43129,
    n43130, n43131, n43132, n43133, n43134, n43135,
    n43136, n43137, n43138, n43139, n43140, n43141,
    n43142, n43143, n43144, n43145, n43146, n43147,
    n43148, n43149, n43150, n43151, n43152, n43153,
    n43154, n43155, n43156, n43157, n43158, n43159,
    n43160, n43161, n43162, n43163, n43164, n43165,
    n43166, n43167, n43168, n43169, n43170, n43171,
    n43172, n43173, n43174, n43175, n43176, n43177,
    n43178, n43179, n43180, n43181, n43182, n43183,
    n43184, n43185, n43186, n43187, n43188, n43189,
    n43190, n43191, n43192, n43193, n43194, n43195,
    n43196, n43197, n43198, n43199, n43200, n43201,
    n43202, n43203, n43204, n43205, n43206, n43207,
    n43208, n43209, n43210, n43211, n43212, n43213,
    n43214, n43215, n43216, n43217, n43218, n43219,
    n43220, n43221, n43222, n43223, n43224, n43225,
    n43226, n43227, n43228, n43229, n43230, n43231,
    n43232, n43233, n43234, n43235, n43236, n43237,
    n43238, n43239, n43240, n43241, n43242, n43243,
    n43244, n43245, n43246, n43247, n43248, n43249,
    n43250, n43251, n43252, n43253, n43254, n43255,
    n43256, n43257, n43258, n43259, n43260, n43261,
    n43262, n43263, n43264, n43265, n43266, n43267,
    n43268, n43269, n43270, n43271, n43272, n43273,
    n43274, n43275, n43276, n43277, n43278, n43279,
    n43280, n43281, n43282, n43283, n43284, n43285,
    n43286, n43287, n43288, n43289, n43290, n43291,
    n43292, n43293, n43294, n43295, n43296, n43297,
    n43298, n43299, n43300, n43301, n43302, n43303,
    n43304, n43305, n43306, n43307, n43308, n43309,
    n43310, n43311, n43312, n43313, n43314, n43315,
    n43316, n43317, n43318, n43319, n43320, n43321,
    n43322, n43323, n43324, n43325, n43326, n43327,
    n43328, n43329, n43330, n43331, n43332, n43333,
    n43334, n43335, n43336, n43337, n43338, n43339,
    n43340, n43341, n43342, n43344, n43345, n43346,
    n43347, n43348, n43349, n43350, n43351, n43352,
    n43353, n43354, n43355, n43356, n43357, n43358,
    n43359, n43360, n43361, n43362, n43363, n43364,
    n43365, n43366, n43367, n43368, n43369, n43370,
    n43371, n43372, n43373, n43374, n43375, n43376,
    n43377, n43378, n43379, n43380, n43381, n43382,
    n43383, n43384, n43385, n43386, n43387, n43388,
    n43389, n43390, n43391, n43392, n43393, n43394,
    n43395, n43396, n43397, n43398, n43399, n43400,
    n43401, n43402, n43403, n43404, n43405, n43406,
    n43407, n43408, n43409, n43410, n43411, n43412,
    n43413, n43414, n43415, n43416, n43417, n43418,
    n43419, n43420, n43421, n43422, n43423, n43424,
    n43425, n43426, n43427, n43428, n43429, n43430,
    n43431, n43432, n43433, n43434, n43435, n43436,
    n43437, n43438, n43439, n43440, n43441, n43442,
    n43443, n43444, n43445, n43446, n43447, n43448,
    n43449, n43450, n43451, n43452, n43453, n43454,
    n43455, n43456, n43457, n43458, n43459, n43460,
    n43461, n43462, n43463, n43464, n43465, n43466,
    n43467, n43468, n43469, n43470, n43471, n43472,
    n43473, n43474, n43475, n43476, n43477, n43478,
    n43479, n43480, n43481, n43482, n43483, n43484,
    n43485, n43486, n43487, n43488, n43489, n43490,
    n43491, n43492, n43493, n43494, n43495, n43496,
    n43497, n43498, n43499, n43500, n43501, n43502,
    n43503, n43504, n43505, n43506, n43507, n43508,
    n43509, n43510, n43511, n43512, n43513, n43514,
    n43515, n43516, n43517, n43518, n43519, n43520,
    n43521, n43522, n43523, n43524, n43525, n43526,
    n43527, n43528, n43529, n43530, n43531, n43532,
    n43533, n43534, n43535, n43536, n43537, n43538,
    n43539, n43540, n43541, n43542, n43543, n43544,
    n43545, n43546, n43547, n43548, n43549, n43550,
    n43551, n43552, n43553, n43554, n43555, n43556,
    n43557, n43558, n43559, n43560, n43561, n43562,
    n43563, n43564, n43565, n43566, n43567, n43568,
    n43569, n43570, n43571, n43572, n43573, n43574,
    n43575, n43576, n43577, n43578, n43579, n43580,
    n43581, n43582, n43583, n43584, n43585, n43586,
    n43587, n43588, n43589, n43590, n43591, n43592,
    n43593, n43594, n43595, n43596, n43597, n43598,
    n43599, n43601, n43602, n43603, n43604, n43605,
    n43606, n43607, n43608, n43609, n43610, n43611,
    n43612, n43613, n43614, n43615, n43616, n43617,
    n43618, n43619, n43620, n43621, n43622, n43623,
    n43624, n43625, n43626, n43627, n43628, n43629,
    n43630, n43631, n43632, n43633, n43634, n43635,
    n43636, n43637, n43638, n43639, n43640, n43641,
    n43642, n43643, n43644, n43645, n43646, n43647,
    n43648, n43649, n43650, n43651, n43652, n43653,
    n43654, n43655, n43656, n43657, n43658, n43659,
    n43660, n43661, n43662, n43663, n43664, n43665,
    n43666, n43667, n43668, n43669, n43670, n43671,
    n43672, n43673, n43674, n43675, n43676, n43677,
    n43678, n43679, n43680, n43681, n43682, n43683,
    n43684, n43685, n43686, n43687, n43688, n43689,
    n43690, n43691, n43692, n43693, n43694, n43695,
    n43696, n43697, n43698, n43699, n43700, n43701,
    n43702, n43703, n43704, n43705, n43706, n43707,
    n43708, n43709, n43710, n43711, n43712, n43713,
    n43714, n43715, n43716, n43717, n43718, n43719,
    n43720, n43721, n43722, n43723, n43724, n43725,
    n43726, n43727, n43728, n43729, n43730, n43731,
    n43732, n43733, n43734, n43735, n43736, n43737,
    n43738, n43739, n43740, n43741, n43742, n43743,
    n43744, n43745, n43746, n43747, n43748, n43749,
    n43750, n43751, n43752, n43753, n43754, n43755,
    n43756, n43757, n43758, n43759, n43760, n43761,
    n43762, n43763, n43764, n43765, n43766, n43767,
    n43768, n43769, n43770, n43771, n43772, n43773,
    n43774, n43775, n43776, n43777, n43778, n43779,
    n43780, n43781, n43782, n43783, n43784, n43785,
    n43786, n43787, n43788, n43789, n43790, n43791,
    n43792, n43793, n43794, n43795, n43796, n43797,
    n43798, n43799, n43800, n43801, n43802, n43803,
    n43804, n43805, n43806, n43807, n43808, n43809,
    n43810, n43811, n43812, n43813, n43814, n43815,
    n43816, n43817, n43818, n43819, n43820, n43821,
    n43822, n43823, n43824, n43825, n43826, n43827,
    n43828, n43829, n43830, n43831, n43832, n43833,
    n43834, n43835, n43836, n43837, n43838, n43839,
    n43840, n43841, n43842, n43843, n43844, n43845,
    n43846, n43847, n43848, n43849, n43850, n43851,
    n43852, n43853, n43854, n43855, n43856, n43857,
    n43858, n43859, n43860, n43861, n43862, n43863,
    n43864, n43865, n43866, n43867, n43868, n43869,
    n43870, n43871, n43872, n43873, n43874, n43875,
    n43876, n43877, n43878, n43879, n43880, n43881,
    n43882, n43883, n43884, n43885, n43886, n43887,
    n43888, n43889, n43890, n43891, n43892, n43893,
    n43894, n43895, n43896, n43897, n43898, n43899,
    n43900, n43901, n43902, n43903, n43904, n43905,
    n43906, n43907, n43908, n43909, n43910, n43911,
    n43912, n43913, n43914, n43915, n43916, n43917,
    n43918, n43919, n43920, n43921, n43922, n43923,
    n43924, n43925, n43926, n43927, n43928, n43929,
    n43930, n43931, n43932, n43933, n43934, n43935,
    n43936, n43937, n43938, n43939, n43940, n43941,
    n43942, n43943, n43944, n43945, n43946, n43947,
    n43948, n43949, n43950, n43951, n43952, n43953,
    n43954, n43955, n43956, n43957, n43958, n43959,
    n43960, n43961, n43962, n43963, n43964, n43965,
    n43966, n43967, n43968, n43969, n43970, n43971,
    n43972, n43973, n43974, n43975, n43976, n43977,
    n43978, n43979, n43980, n43981, n43982, n43983,
    n43984, n43985, n43986, n43987, n43988, n43989,
    n43990, n43991, n43992, n43993, n43994, n43995,
    n43996, n43997, n43998, n43999, n44000, n44001,
    n44002, n44003, n44004, n44005, n44006, n44007,
    n44008, n44009, n44010, n44011, n44012, n44013,
    n44014, n44015, n44016, n44017, n44018, n44019,
    n44020, n44021, n44022, n44023, n44024, n44025,
    n44026, n44027, n44028, n44029, n44030, n44031,
    n44032, n44033, n44034, n44035, n44036, n44037,
    n44038, n44039, n44040, n44041, n44042, n44043,
    n44044, n44045, n44046, n44047, n44048, n44049,
    n44050, n44051, n44052, n44053, n44054, n44055,
    n44056, n44057, n44058, n44059, n44060, n44061,
    n44062, n44063, n44064, n44065, n44066, n44067,
    n44068, n44069, n44070, n44071, n44072, n44073,
    n44074, n44075, n44076, n44077, n44078, n44079,
    n44080, n44081, n44082, n44083, n44084, n44085,
    n44086, n44087, n44088, n44089, n44090, n44091,
    n44092, n44093, n44094, n44095, n44096, n44097,
    n44098, n44099, n44100, n44101, n44102, n44103,
    n44104, n44105, n44106, n44107, n44108, n44109,
    n44110, n44111, n44112, n44113, n44114, n44115,
    n44116, n44117, n44118, n44119, n44120, n44121,
    n44122, n44123, n44124, n44125, n44126, n44127,
    n44128, n44129, n44130, n44131, n44132, n44133,
    n44134, n44135, n44136, n44137, n44138, n44139,
    n44140, n44141, n44142, n44143, n44144, n44145,
    n44146, n44147, n44148, n44149, n44150, n44151,
    n44152, n44153, n44154, n44155, n44156, n44157,
    n44158, n44159, n44160, n44161, n44162, n44163,
    n44164, n44165, n44166, n44167, n44168, n44169,
    n44170, n44171, n44172, n44173, n44174, n44175,
    n44176, n44177, n44178, n44179, n44180, n44181,
    n44182, n44183, n44184, n44185, n44186, n44187,
    n44188, n44189, n44190, n44191, n44192, n44193,
    n44194, n44195, n44196, n44197, n44198, n44199,
    n44200, n44201, n44202, n44203, n44204, n44205,
    n44206, n44207, n44208, n44209, n44210, n44211,
    n44212, n44213, n44214, n44215, n44216, n44217,
    n44218, n44219, n44220, n44221, n44222, n44223,
    n44224, n44225, n44226, n44227, n44228, n44229,
    n44230, n44231, n44232, n44233, n44234, n44235,
    n44236, n44237, n44238, n44239, n44240, n44241,
    n44242, n44243, n44244, n44245, n44246, n44247,
    n44248, n44249, n44250, n44251, n44252, n44253,
    n44254, n44255, n44256, n44257, n44258, n44259,
    n44260, n44261, n44262, n44263, n44264, n44265,
    n44266, n44267, n44268, n44269, n44270, n44271,
    n44272, n44273, n44274, n44275, n44276, n44277,
    n44278, n44279, n44280, n44281, n44282, n44283,
    n44284, n44285, n44286, n44287, n44288, n44289,
    n44290, n44291, n44292, n44293, n44294, n44295,
    n44296, n44297, n44298, n44299, n44300, n44301,
    n44302, n44303, n44304, n44305, n44306, n44307,
    n44308, n44309, n44310, n44311, n44312, n44313,
    n44314, n44315, n44316, n44317, n44318, n44319,
    n44320, n44321, n44322, n44323, n44324, n44325,
    n44326, n44327, n44328, n44329, n44330, n44331,
    n44332, n44333, n44334, n44335, n44336, n44337,
    n44338, n44339, n44340, n44341, n44342, n44343,
    n44344, n44345, n44346, n44347, n44348, n44349,
    n44350, n44351, n44352, n44353, n44354, n44355,
    n44356, n44357, n44358, n44359, n44360, n44361,
    n44362, n44363, n44364, n44365, n44366, n44367,
    n44368, n44369, n44370, n44371, n44372, n44373,
    n44374, n44375, n44376, n44377, n44378, n44379,
    n44380, n44381, n44382, n44383, n44384, n44385,
    n44386, n44387, n44388, n44389, n44390, n44391,
    n44392, n44393, n44394, n44395, n44396, n44397,
    n44398, n44399, n44400, n44401, n44402, n44403,
    n44404, n44405, n44406, n44407, n44408, n44409,
    n44410, n44411, n44412, n44413, n44414, n44415,
    n44416, n44417, n44418, n44419, n44420, n44421,
    n44422, n44423, n44424, n44425, n44426, n44427,
    n44428, n44429, n44430, n44431, n44432, n44433,
    n44434, n44435, n44436, n44437, n44438, n44439,
    n44440, n44441, n44442, n44443, n44444, n44445,
    n44446, n44447, n44448, n44449, n44450, n44451,
    n44452, n44453, n44454, n44455, n44456, n44457,
    n44458, n44459, n44460, n44461, n44462, n44463,
    n44464, n44465, n44466, n44467, n44468, n44469,
    n44470, n44471, n44472, n44473, n44474, n44475,
    n44476, n44477, n44478, n44480, n44481, n44482,
    n44483, n44484, n44485, n44486, n44487, n44488,
    n44489, n44490, n44491, n44492, n44493, n44494,
    n44495, n44496, n44497, n44498, n44499, n44500,
    n44501, n44502, n44503, n44504, n44505, n44506,
    n44507, n44508, n44509, n44510, n44511, n44512,
    n44513, n44515, n44516, n44517, n44518, n44519,
    n44520, n44521, n44522, n44523, n44524, n44525,
    n44526, n44527, n44528, n44529, n44530, n44531,
    n44533, n44534, n44535, n44536, n44537, n44538,
    n44539, n44541, n44542, n44543, n44544, n44545,
    n44546, n44547, n44548, n44549, n44550, n44551,
    n44552, n44553, n44554, n44556, n44557, n44558,
    n44559, n44560, n44561, n44562, n44563, n44564,
    n44565, n44566, n44567, n44568, n44569, n44570,
    n44571, n44572, n44573, n44574, n44575, n44576,
    n44577, n44578, n44579, n44580, n44581, n44582,
    n44583, n44584, n44585, n44586, n44587, n44588,
    n44589, n44590, n44591, n44592, n44593, n44594,
    n44595, n44596, n44597, n44598, n44599, n44600,
    n44601, n44602, n44603, n44604, n44605, n44606,
    n44607, n44608, n44609, n44610, n44611, n44612,
    n44613, n44614, n44615, n44616, n44617, n44618,
    n44619, n44620, n44621, n44622, n44623, n44624,
    n44625, n44626, n44627, n44628, n44629, n44630,
    n44631, n44632, n44633, n44634, n44635, n44636,
    n44637, n44638, n44639, n44640, n44641, n44642,
    n44643, n44644, n44645, n44646, n44647, n44648,
    n44649, n44650, n44651, n44652, n44653, n44654,
    n44655, n44656, n44657, n44658, n44659, n44660,
    n44661, n44662, n44663, n44664, n44665, n44666,
    n44667, n44668, n44669, n44670, n44671, n44672,
    n44673, n44674, n44675, n44676, n44677, n44678,
    n44679, n44680, n44681, n44682, n44683, n44684,
    n44685, n44686, n44687, n44688, n44689, n44690,
    n44691, n44692, n44693, n44694, n44695, n44696,
    n44697, n44698, n44699, n44700, n44701, n44702,
    n44703, n44704, n44705, n44706, n44707, n44708,
    n44709, n44710, n44711, n44712, n44713, n44714,
    n44715, n44716, n44717, n44718, n44719, n44720,
    n44721, n44722, n44723, n44724, n44725, n44726,
    n44727, n44728, n44729, n44730, n44731, n44732,
    n44733, n44734, n44735, n44736, n44737, n44738,
    n44739, n44740, n44741, n44742, n44743, n44744,
    n44745, n44746, n44747, n44748, n44749, n44750,
    n44751, n44752, n44753, n44754, n44755, n44756,
    n44757, n44758, n44759, n44760, n44761, n44762,
    n44763, n44764, n44765, n44766, n44767, n44768,
    n44769, n44770, n44771, n44772, n44773, n44774,
    n44775, n44776, n44777, n44778, n44779, n44780,
    n44781, n44782, n44783, n44784, n44786, n44787,
    n44788, n44789, n44790, n44791, n44792, n44794,
    n44795, n44796, n44797, n44798, n44799, n44800,
    n44802, n44803, n44804, n44805, n44806, n44807,
    n44808, n44809, n44810, n44811, n44812, n44813,
    n44814, n44815, n44816, n44817, n44818, n44819,
    n44820, n44821, n44822, n44823, n44824, n44825,
    n44826, n44827, n44828, n44829, n44830, n44831,
    n44832, n44833, n44834, n44835, n44836, n44837,
    n44838, n44839, n44840, n44841, n44842, n44843,
    n44844, n44845, n44846, n44847, n44848, n44849,
    n44850, n44851, n44852, n44853, n44854, n44855,
    n44856, n44857, n44858, n44859, n44860, n44861,
    n44862, n44863, n44864, n44865, n44866, n44867,
    n44868, n44869, n44870, n44871, n44872, n44873,
    n44874, n44875, n44876, n44877, n44878, n44879,
    n44880, n44881, n44882, n44883, n44884, n44885,
    n44886, n44887, n44888, n44889, n44890, n44891,
    n44892, n44893, n44894, n44895, n44896, n44897,
    n44898, n44899, n44900, n44901, n44902, n44903,
    n44904, n44905, n44906, n44907, n44908, n44909,
    n44910, n44911, n44912, n44913, n44914, n44916,
    n44917, n44918, n44919, n44920, n44921, n44923,
    n44924, n44925, n44926, n44927, n44928, n44929,
    n44931, n44932, n44933, n44934, n44935, n44936,
    n44938, n44939, n44940, n44941, n44942, n44943,
    n44945, n44946, n44947, n44948, n44949, n44950,
    n44951, n44952, n44953, n44954, n44955, n44956,
    n44957, n44958, n44959, n44960, n44961, n44962,
    n44963, n44964, n44965, n44967, n44968, n44969,
    n44970, n44971, n44972, n44973, n44974, n44975,
    n44976, n44977, n44978, n44979, n44980, n44981,
    n44982, n44983, n44984, n44985, n44986, n44987,
    n44988, n44989, n44990, n44991, n44992, n44993,
    n44994, n44995, n44996, n44997, n44998, n44999,
    n45000, n45001, n45002, n45003, n45004, n45005,
    n45006, n45007, n45008, n45009, n45010, n45011,
    n45012, n45013, n45014, n45015, n45016, n45017,
    n45018, n45019, n45020, n45021, n45022, n45023,
    n45024, n45025, n45026, n45027, n45028, n45029,
    n45030, n45031, n45032, n45033, n45034, n45035,
    n45036, n45037, n45038, n45039, n45040, n45041,
    n45042, n45043, n45044, n45045, n45046, n45047,
    n45048, n45049, n45050, n45051, n45052, n45053,
    n45054, n45055, n45056, n45057, n45058, n45059,
    n45060, n45061, n45062, n45063, n45064, n45066,
    n45067, n45068, n45069, n45070, n45071, n45072,
    n45073, n45074, n45075, n45076, n45077, n45078,
    n45079, n45080, n45081, n45082, n45083, n45084,
    n45085, n45087, n45088, n45089, n45090, n45091,
    n45092, n45093, n45094, n45095, n45096, n45097,
    n45098, n45099, n45100, n45101, n45102, n45103,
    n45104, n45105, n45106, n45107, n45108, n45109,
    n45110, n45111, n45112, n45113, n45114, n45115,
    n45116, n45117, n45118, n45119, n45120, n45121,
    n45122, n45123, n45124, n45125, n45126, n45127,
    n45128, n45129, n45130, n45131, n45132, n45133,
    n45134, n45135, n45136, n45137, n45138, n45140,
    n45141, n45142, n45143, n45144, n45145, n45146,
    n45147, n45148, n45150, n45151, n45152, n45153,
    n45154, n45155, n45156, n45157, n45158, n45159,
    n45160, n45161, n45162, n45163, n45165, n45166,
    n45167, n45168, n45169, n45170, n45171, n45172,
    n45173, n45174, n45175, n45176, n45177, n45178,
    n45179, n45180, n45181, n45182, n45183, n45184,
    n45185, n45186, n45187, n45189, n45190, n45191,
    n45192, n45193, n45194, n45195, n45196, n45197,
    n45198, n45199, n45200, n45201, n45203, n45204,
    n45205, n45206, n45207, n45208, n45209, n45210,
    n45211, n45212, n45213, n45214, n45215, n45216,
    n45217, n45218, n45219, n45220, n45221, n45222,
    n45223, n45224, n45225, n45226, n45227, n45228,
    n45229, n45230, n45231, n45232, n45233, n45234,
    n45235, n45236, n45237, n45238, n45239, n45240,
    n45241, n45242, n45243, n45244, n45245, n45246,
    n45247, n45248, n45249, n45250, n45251, n45252,
    n45253, n45254, n45255, n45256, n45257, n45258,
    n45259, n45260, n45261, n45262, n45263, n45264,
    n45265, n45266, n45267, n45268, n45269, n45270,
    n45271, n45272, n45273, n45274, n45275, n45276,
    n45277, n45278, n45279, n45280, n45281, n45282,
    n45283, n45284, n45285, n45286, n45287, n45288,
    n45289, n45290, n45291, n45292, n45293, n45294,
    n45295, n45296, n45297, n45298, n45299, n45300,
    n45301, n45302, n45303, n45304, n45305, n45306,
    n45307, n45308, n45309, n45310, n45311, n45312,
    n45313, n45314, n45315, n45316, n45317, n45318,
    n45319, n45320, n45321, n45322, n45323, n45324,
    n45325, n45326, n45327, n45328, n45329, n45330,
    n45331, n45332, n45333, n45334, n45335, n45336,
    n45337, n45338, n45339, n45340, n45341, n45342,
    n45343, n45344, n45345, n45346, n45347, n45348,
    n45349, n45350, n45351, n45352, n45353, n45354,
    n45355, n45356, n45357, n45358, n45359, n45360,
    n45361, n45362, n45363, n45364, n45365, n45366,
    n45367, n45368, n45369, n45370, n45371, n45372,
    n45373, n45374, n45375, n45376, n45377, n45378,
    n45379, n45380, n45381, n45382, n45383, n45384,
    n45385, n45386, n45387, n45388, n45389, n45390,
    n45391, n45392, n45393, n45394, n45395, n45396,
    n45397, n45398, n45399, n45401, n45402, n45403,
    n45404, n45405, n45406, n45407, n45408, n45409,
    n45410, n45411, n45412, n45413, n45414, n45415,
    n45417, n45419, n45420, n45421, n45422, n45423,
    n45424, n45425, n45426, n45427, n45428, n45429,
    n45430, n45431, n45432, n45433, n45434, n45435,
    n45436, n45437, n45438, n45440, n45441, n45442,
    n45443, n45444, n45445, n45446, n45447, n45448,
    n45449, n45450, n45451, n45452, n45454, n45455,
    n45456, n45457, n45458, n45459, n45460, n45461,
    n45462, n45463, n45464, n45465, n45466, n45467,
    n45468, n45469, n45470, n45471, n45472, n45473,
    n45474, n45475, n45476, n45477, n45478, n45479,
    n45480, n45481, n45482, n45483, n45484, n45485,
    n45486, n45487, n45488, n45489, n45490, n45491,
    n45492, n45493, n45494, n45495, n45496, n45497,
    n45499, n45500, n45501, n45502, n45503, n45504,
    n45505, n45506, n45507, n45508, n45509, n45510,
    n45511, n45512, n45513, n45514, n45515, n45516,
    n45517, n45518, n45519, n45520, n45521, n45522,
    n45523, n45524, n45525, n45526, n45528, n45529,
    n45530, n45531, n45532, n45533, n45534, n45535,
    n45536, n45537, n45538, n45539, n45540, n45541,
    n45542, n45543, n45544, n45545, n45546, n45547,
    n45548, n45550, n45551, n45552, n45553, n45554,
    n45555, n45556, n45557, n45558, n45559, n45560,
    n45561, n45562, n45563, n45564, n45565, n45566,
    n45567, n45568, n45570, n45572, n45573, n45574,
    n45575, n45576, n45577, n45578, n45579, n45580,
    n45581, n45582, n45583, n45584, n45585, n45586,
    n45588, n45589, n45590, n45591, n45592, n45593,
    n45594, n45595, n45596, n45597, n45598, n45599,
    n45600, n45601, n45603, n45604, n45605, n45606,
    n45607, n45608, n45609, n45611, n45612, n45613,
    n45614, n45615, n45616, n45618, n45619, n45620,
    n45621, n45622, n45624, n45625, n45626, n45627,
    n45628, n45629, n45630, n45631, n45632, n45633,
    n45634, n45635, n45636, n45637, n45638, n45639,
    n45640, n45641, n45642, n45643, n45644, n45645,
    n45646, n45647, n45648, n45649, n45650, n45651,
    n45652, n45653, n45654, n45656, n45657, n45658,
    n45659, n45660, n45661, n45663, n45664, n45665,
    n45666, n45668, n45669, n45670, n45671, n45672,
    n45673, n45675, n45676, n45677, n45679, n45680,
    n45681, n45682, n45683, n45684, n45685, n45686,
    n45687, n45688, n45689, n45691, n45692, n45693,
    n45694, n45695, n45696, n45697, n45698, n45699,
    n45700, n45701, n45702, n45703, n45704, n45705,
    n45707, n45708, n45709, n45710, n45711, n45712,
    n45713, n45714, n45715, n45716, n45717, n45718,
    n45719, n45720, n45721, n45722, n45723, n45724,
    n45725, n45726, n45727, n45728, n45729, n45731,
    n45732, n45733, n45734, n45735, n45736, n45737,
    n45738, n45739, n45740, n45741, n45742, n45743,
    n45744, n45745, n45746, n45747, n45748, n45749,
    n45750, n45751, n45752, n45753, n45754, n45755,
    n45756, n45757, n45758, n45759, n45760, n45761,
    n45762, n45763, n45764, n45765, n45766, n45767,
    n45768, n45769, n45770, n45771, n45773, n45774,
    n45775, n45777, n45778, n45779, n45780, n45781,
    n45782, n45783, n45784, n45785, n45786, n45788,
    n45789, n45790, n45791, n45792, n45793, n45794,
    n45795, n45796, n45798, n45799, n45800, n45801,
    n45802, n45803, n45804, n45805, n45806, n45808,
    n45809, n45810, n45811, n45813, n45814, n45815,
    n45816, n45817, n45818, n45819, n45820, n45821,
    n45822, n45823, n45824, n45825, n45826, n45827,
    n45828, n45829, n45830, n45831, n45832, n45833,
    n45834, n45835, n45836, n45837, n45838, n45839,
    n45840, n45841, n45842, n45843, n45844, n45846,
    n45847, n45848, n45849, n45851, n45852, n45853,
    n45854, n45855, n45856, n45857, n45858, n45859,
    n45860, n45861, n45862, n45863, n45864, n45865,
    n45866, n45867, n45868, n45869, n45870, n45871,
    n45872, n45873, n45874, n45875, n45876, n45877,
    n45878, n45879, n45880, n45881, n45882, n45884,
    n45885, n45886, n45887, n45889, n45890, n45891,
    n45892, n45893, n45894, n45895, n45896, n45897,
    n45898, n45900, n45901, n45902, n45903, n45904,
    n45907, n45908, n45910, n45911, n45913, n45915,
    n45916, n45918, n45919, n45920, n45921, n45922,
    n45923, n45924, n45925, n45926, n45927, n45928,
    n45929, n45930, n45931, n45932, n45933, n45934,
    n45935, n45936, n45937, n45938, n45939, n45940,
    n45942, n45943, n45944, n45945, n45946, n45947,
    n45948, n45949, n45950, n45951, n45952, n45953,
    n45954, n45955, n45956, n45957, n45958, n45959,
    n45960, n45961, n45962, n45963, n45964, n45965,
    n45966, n45967, n45968, n45969, n45970, n45971,
    n45972, n45973, n45974, n45975, n45976, n45977,
    n45978, n45979, n45980, n45981, n45982, n45984,
    n45985, n45986, n45987, n45988, n45989, n45990,
    n45991, n45992, n45993, n45994, n45995, n45996,
    n45997, n45998, n45999, n46000, n46001, n46002,
    n46003, n46004, n46005, n46006, n46007, n46008,
    n46009, n46010, n46011, n46012, n46013, n46014,
    n46015, n46016, n46017, n46018, n46019, n46020,
    n46021, n46022, n46023, n46024, n46025, n46026,
    n46027, n46028, n46029, n46030, n46031, n46032,
    n46033, n46034, n46035, n46036, n46037, n46038,
    n46039, n46040, n46041, n46042, n46043, n46044,
    n46045, n46046, n46047, n46048, n46049, n46050,
    n46051, n46052, n46053, n46054, n46055, n46056,
    n46057, n46058, n46059, n46060, n46061, n46062,
    n46063, n46064, n46065, n46066, n46067, n46068,
    n46069, n46070, n46071, n46072, n46073, n46074,
    n46075, n46076, n46077, n46078, n46079, n46080,
    n46081, n46082, n46083, n46084, n46085, n46086,
    n46087, n46088, n46089, n46090, n46091, n46092,
    n46093, n46094, n46095, n46096, n46097, n46098,
    n46099, n46100, n46101, n46102, n46103, n46104,
    n46105, n46106, n46107, n46108, n46109, n46110,
    n46111, n46112, n46113, n46114, n46115, n46116,
    n46117, n46118, n46119, n46120, n46121, n46122,
    n46123, n46124, n46125, n46126, n46127, n46128,
    n46129, n46130, n46131, n46132, n46133, n46134,
    n46135, n46136, n46137, n46138, n46139, n46140,
    n46141, n46142, n46143, n46144, n46145, n46146,
    n46147, n46148, n46149, n46150, n46151, n46152,
    n46153, n46154, n46155, n46156, n46157, n46158,
    n46159, n46160, n46161, n46162, n46163, n46164,
    n46165, n46166, n46167, n46168, n46169, n46170,
    n46171, n46172, n46173, n46174, n46175, n46176,
    n46177, n46178, n46179, n46180, n46181, n46182,
    n46183, n46184, n46185, n46186, n46187, n46188,
    n46189, n46190, n46191, n46192, n46193, n46194,
    n46195, n46196, n46197, n46198, n46199, n46200,
    n46201, n46202, n46203, n46204, n46205, n46206,
    n46207, n46208, n46209, n46210, n46211, n46212,
    n46213, n46214, n46215, n46216, n46217, n46218,
    n46219, n46220, n46221, n46222, n46223, n46224,
    n46225, n46226, n46227, n46228, n46229, n46230,
    n46231, n46232, n46233, n46234, n46235, n46236,
    n46237, n46238, n46239, n46240, n46241, n46242,
    n46243, n46244, n46245, n46246, n46247, n46248,
    n46249, n46250, n46251, n46252, n46253, n46254,
    n46255, n46256, n46257, n46258, n46259, n46260,
    n46261, n46262, n46263, n46264, n46265, n46266,
    n46267, n46268, n46269, n46270, n46271, n46272,
    n46273, n46274, n46275, n46276, n46277, n46278,
    n46279, n46280, n46281, n46282, n46283, n46284,
    n46285, n46286, n46287, n46288, n46289, n46290,
    n46291, n46292, n46293, n46294, n46295, n46296,
    n46297, n46298, n46299, n46300, n46301, n46302,
    n46303, n46304, n46305, n46306, n46307, n46308,
    n46309, n46310, n46311, n46312, n46313, n46314,
    n46315, n46316, n46317, n46318, n46319, n46320,
    n46321, n46322, n46323, n46324, n46325, n46326,
    n46327, n46328, n46329, n46330, n46331, n46332,
    n46333, n46334, n46335, n46336, n46337, n46338,
    n46339, n46340, n46341, n46342, n46343, n46344,
    n46345, n46346, n46347, n46348, n46349, n46350,
    n46351, n46352, n46353, n46354, n46355, n46356,
    n46357, n46358, n46359, n46360, n46361, n46362,
    n46363, n46364, n46365, n46366, n46367, n46368,
    n46369, n46370, n46371, n46372, n46373, n46374,
    n46375, n46376, n46377, n46378, n46379, n46380,
    n46381, n46382, n46383, n46384, n46385, n46386,
    n46387, n46388, n46389, n46390, n46391, n46392,
    n46393, n46394, n46395, n46396, n46397, n46398,
    n46399, n46400, n46401, n46402, n46403, n46404,
    n46405, n46406, n46407, n46408, n46409, n46410,
    n46411, n46412, n46413, n46414, n46415, n46416,
    n46417, n46418, n46419, n46420, n46421, n46422,
    n46423, n46424, n46425, n46426, n46427, n46428,
    n46429, n46430, n46431, n46432, n46433, n46434,
    n46435, n46436, n46437, n46438, n46439, n46440,
    n46441, n46442, n46443, n46444, n46445, n46446,
    n46447, n46448, n46449, n46450, n46451, n46452,
    n46453, n46454, n46455, n46456, n46457, n46458,
    n46459, n46460, n46461, n46462, n46463, n46464,
    n46465, n46466, n46467, n46468, n46469, n46470,
    n46471, n46472, n46473, n46474, n46475, n46476,
    n46477, n46478, n46479, n46480, n46481, n46482,
    n46483, n46484, n46485, n46486, n46487, n46488,
    n46489, n46490, n46491, n46492, n46493, n46494,
    n46496, n46497, n46498, n46499, n46500, n46501,
    n46502, n46503, n46504, n46505, n46506, n46507,
    n46508, n46509, n46510, n46511, n46512, n46513,
    n46514, n46515, n46516, n46517, n46518, n46519,
    n46520, n46521, n46522, n46523, n46524, n46525,
    n46526, n46527, n46528, n46529, n46530, n46531,
    n46532, n46533, n46534, n46535, n46536, n46537,
    n46538, n46539, n46540, n46541, n46542, n46543,
    n46544, n46545, n46546, n46547, n46548, n46549,
    n46550, n46551, n46552, n46553, n46554, n46555,
    n46556, n46557, n46558, n46559, n46560, n46561,
    n46562, n46563, n46564, n46565, n46566, n46567,
    n46568, n46569, n46570, n46571, n46572, n46573,
    n46574, n46575, n46576, n46577, n46578, n46579,
    n46580, n46581, n46582, n46583, n46584, n46585,
    n46586, n46587, n46588, n46589, n46590, n46591,
    n46592, n46593, n46594, n46595, n46596, n46597,
    n46598, n46599, n46600, n46601, n46602, n46603,
    n46604, n46605, n46606, n46607, n46608, n46609,
    n46610, n46611, n46612, n46613, n46614, n46615,
    n46616, n46617, n46618, n46619, n46620, n46621,
    n46622, n46623, n46624, n46625, n46626, n46627,
    n46628, n46629, n46630, n46631, n46632, n46633,
    n46634, n46635, n46636, n46637, n46638, n46639,
    n46640, n46641, n46642, n46643, n46644, n46645,
    n46646, n46647, n46648, n46649, n46650, n46651,
    n46652, n46653, n46654, n46655, n46656, n46657,
    n46658, n46659, n46660, n46661, n46662, n46663,
    n46664, n46665, n46666, n46667, n46668, n46669,
    n46670, n46671, n46672, n46673, n46674, n46675,
    n46676, n46677, n46678, n46679, n46680, n46681,
    n46682, n46683, n46684, n46685, n46686, n46687,
    n46688, n46689, n46690, n46691, n46692, n46693,
    n46694, n46695, n46696, n46697, n46698, n46699,
    n46700, n46701, n46702, n46703, n46704, n46705,
    n46706, n46707, n46708, n46709, n46710, n46711,
    n46712, n46713, n46714, n46715, n46716, n46717,
    n46718, n46719, n46720, n46721, n46722, n46723,
    n46724, n46725, n46726, n46727, n46728, n46729,
    n46730, n46731, n46732, n46733, n46734, n46735,
    n46736, n46737, n46738, n46739, n46740, n46741,
    n46742, n46743, n46744, n46745, n46746, n46747,
    n46748, n46749, n46750, n46751, n46752, n46753,
    n46754, n46755, n46756, n46757, n46758, n46759,
    n46760, n46761, n46762, n46763, n46764, n46765,
    n46766, n46767, n46768, n46769, n46770, n46771,
    n46772, n46773, n46774, n46775, n46776, n46777,
    n46778, n46779, n46780, n46781, n46782, n46783,
    n46784, n46785, n46786, n46787, n46788, n46789,
    n46790, n46791, n46792, n46793, n46794, n46795,
    n46796, n46797, n46798, n46799, n46800, n46801,
    n46802, n46803, n46804, n46805, n46806, n46807,
    n46808, n46809, n46810, n46811, n46813, n46814,
    n46815, n46816, n46817, n46818, n46819, n46820,
    n46821, n46822, n46823, n46824, n46825, n46826,
    n46827, n46828, n46829, n46830, n46831, n46832,
    n46833, n46834, n46835, n46836, n46837, n46838,
    n46839, n46840, n46841, n46842, n46843, n46844,
    n46845, n46846, n46847, n46848, n46849, n46850,
    n46851, n46852, n46853, n46854, n46855, n46856,
    n46857, n46858, n46859, n46860, n46861, n46862,
    n46863, n46864, n46865, n46866, n46867, n46868,
    n46869, n46870, n46871, n46872, n46873, n46874,
    n46875, n46876, n46877, n46878, n46879, n46880,
    n46881, n46882, n46883, n46884, n46885, n46886,
    n46887, n46888, n46889, n46890, n46891, n46892,
    n46893, n46894, n46895, n46896, n46897, n46898,
    n46899, n46900, n46901, n46902, n46903, n46904,
    n46905, n46906, n46907, n46908, n46909, n46910,
    n46911, n46912, n46913, n46914, n46915, n46916,
    n46917, n46918, n46919, n46920, n46921, n46922,
    n46923, n46924, n46925, n46926, n46927, n46928,
    n46929, n46930, n46931, n46932, n46933, n46934,
    n46935, n46936, n46937, n46938, n46939, n46940,
    n46941, n46942, n46943, n46944, n46945, n46946,
    n46947, n46948, n46949, n46950, n46951, n46952,
    n46953, n46954, n46955, n46956, n46957, n46958,
    n46959, n46960, n46961, n46962, n46963, n46964,
    n46965, n46966, n46967, n46968, n46969, n46970,
    n46971, n46972, n46973, n46974, n46975, n46976,
    n46977, n46978, n46979, n46980, n46981, n46982,
    n46983, n46984, n46985, n46986, n46987, n46988,
    n46989, n46990, n46991, n46992, n46993, n46994,
    n46995, n46996, n46997, n46998, n46999, n47000,
    n47001, n47002, n47003, n47004, n47005, n47006,
    n47007, n47008, n47009, n47010, n47011, n47012,
    n47013, n47014, n47015, n47016, n47017, n47018,
    n47019, n47020, n47021, n47022, n47023, n47024,
    n47025, n47026, n47027, n47028, n47029, n47030,
    n47031, n47032, n47033, n47034, n47035, n47036,
    n47037, n47038, n47039, n47040, n47041, n47042,
    n47043, n47044, n47045, n47046, n47047, n47048,
    n47049, n47050, n47051, n47052, n47053, n47054,
    n47055, n47056, n47057, n47058, n47059, n47060,
    n47061, n47062, n47063, n47064, n47065, n47066,
    n47067, n47068, n47069, n47070, n47071, n47072,
    n47073, n47074, n47075, n47076, n47077, n47078,
    n47079, n47080, n47081, n47082, n47083, n47084,
    n47085, n47086, n47087, n47088, n47089, n47090,
    n47091, n47092, n47093, n47094, n47095, n47096,
    n47097, n47098, n47099, n47100, n47101, n47102,
    n47103, n47104, n47105, n47106, n47107, n47108,
    n47109, n47110, n47111, n47112, n47113, n47114,
    n47115, n47116, n47117, n47118, n47119, n47120,
    n47121, n47123, n47124, n47125, n47126, n47127,
    n47128, n47129, n47130, n47131, n47132, n47133,
    n47134, n47135, n47136, n47137, n47138, n47139,
    n47140, n47141, n47142, n47143, n47144, n47145,
    n47146, n47147, n47148, n47149, n47150, n47151,
    n47152, n47153, n47154, n47155, n47156, n47157,
    n47158, n47159, n47160, n47161, n47162, n47163,
    n47164, n47165, n47166, n47167, n47168, n47169,
    n47170, n47171, n47172, n47173, n47174, n47175,
    n47176, n47177, n47178, n47179, n47180, n47181,
    n47182, n47183, n47184, n47185, n47186, n47187,
    n47188, n47189, n47190, n47191, n47192, n47193,
    n47194, n47195, n47196, n47197, n47198, n47199,
    n47200, n47201, n47202, n47203, n47204, n47205,
    n47206, n47207, n47208, n47209, n47210, n47211,
    n47212, n47213, n47214, n47215, n47216, n47217,
    n47218, n47219, n47220, n47221, n47222, n47223,
    n47224, n47225, n47226, n47227, n47228, n47229,
    n47230, n47231, n47232, n47233, n47234, n47235,
    n47236, n47237, n47238, n47239, n47240, n47241,
    n47242, n47243, n47244, n47245, n47246, n47247,
    n47248, n47249, n47250, n47251, n47252, n47253,
    n47254, n47255, n47256, n47257, n47258, n47259,
    n47260, n47261, n47262, n47263, n47264, n47265,
    n47266, n47267, n47268, n47269, n47270, n47271,
    n47272, n47273, n47274, n47275, n47276, n47277,
    n47278, n47279, n47280, n47281, n47282, n47283,
    n47284, n47285, n47286, n47287, n47288, n47289,
    n47290, n47291, n47292, n47293, n47294, n47295,
    n47296, n47297, n47298, n47299, n47300, n47301,
    n47302, n47303, n47304, n47305, n47306, n47307,
    n47308, n47309, n47310, n47311, n47312, n47313,
    n47314, n47315, n47316, n47317, n47318, n47319,
    n47320, n47321, n47322, n47323, n47324, n47325,
    n47326, n47327, n47328, n47329, n47330, n47331,
    n47332, n47333, n47334, n47335, n47336, n47337,
    n47338, n47339, n47340, n47341, n47342, n47343,
    n47344, n47345, n47346, n47347, n47348, n47349,
    n47350, n47351, n47352, n47353, n47354, n47355,
    n47356, n47357, n47358, n47359, n47360, n47361,
    n47362, n47363, n47364, n47365, n47366, n47367,
    n47368, n47369, n47370, n47371, n47372, n47373,
    n47374, n47375, n47376, n47377, n47378, n47379,
    n47380, n47381, n47382, n47383, n47384, n47385,
    n47386, n47387, n47388, n47390, n47391, n47392,
    n47393, n47394, n47395, n47396, n47397, n47398,
    n47399, n47400, n47401, n47402, n47403, n47404,
    n47405, n47406, n47407, n47408, n47409, n47410,
    n47411, n47412, n47413, n47414, n47415, n47416,
    n47417, n47418, n47419, n47420, n47421, n47422,
    n47423, n47424, n47425, n47426, n47427, n47428,
    n47429, n47430, n47431, n47432, n47433, n47434,
    n47435, n47436, n47437, n47438, n47439, n47440,
    n47441, n47442, n47443, n47444, n47445, n47446,
    n47447, n47448, n47449, n47450, n47451, n47452,
    n47453, n47454, n47455, n47456, n47457, n47458,
    n47459, n47460, n47461, n47462, n47463, n47464,
    n47465, n47466, n47467, n47468, n47469, n47470,
    n47471, n47472, n47473, n47474, n47475, n47476,
    n47477, n47478, n47479, n47480, n47481, n47482,
    n47483, n47484, n47485, n47486, n47487, n47488,
    n47489, n47490, n47491, n47492, n47493, n47494,
    n47495, n47496, n47497, n47498, n47499, n47500,
    n47501, n47502, n47503, n47504, n47505, n47506,
    n47507, n47508, n47509, n47510, n47511, n47512,
    n47513, n47514, n47515, n47516, n47517, n47518,
    n47519, n47520, n47521, n47522, n47523, n47524,
    n47525, n47526, n47527, n47528, n47529, n47530,
    n47531, n47532, n47533, n47534, n47535, n47536,
    n47537, n47538, n47539, n47540, n47541, n47542,
    n47543, n47544, n47545, n47546, n47547, n47548,
    n47549, n47550, n47551, n47552, n47553, n47554,
    n47555, n47556, n47557, n47558, n47559, n47560,
    n47561, n47562, n47563, n47564, n47565, n47566,
    n47567, n47568, n47569, n47570, n47571, n47572,
    n47573, n47574, n47575, n47576, n47577, n47578,
    n47579, n47580, n47581, n47582, n47583, n47584,
    n47585, n47586, n47587, n47588, n47589, n47590,
    n47591, n47592, n47593, n47594, n47595, n47596,
    n47597, n47598, n47599, n47600, n47601, n47602,
    n47603, n47604, n47605, n47606, n47607, n47608,
    n47609, n47610, n47611, n47612, n47613, n47614,
    n47615, n47616, n47617, n47618, n47619, n47620,
    n47621, n47622, n47623, n47624, n47625, n47626,
    n47627, n47628, n47629, n47630, n47631, n47632,
    n47633, n47634, n47635, n47636, n47637, n47638,
    n47639, n47640, n47641, n47642, n47643, n47645,
    n47646, n47647, n47648, n47649, n47650, n47651,
    n47652, n47653, n47654, n47655, n47656, n47657,
    n47658, n47659, n47660, n47661, n47662, n47663,
    n47664, n47665, n47666, n47667, n47668, n47669,
    n47670, n47671, n47672, n47673, n47674, n47675,
    n47676, n47677, n47678, n47679, n47680, n47681,
    n47682, n47683, n47684, n47685, n47686, n47687,
    n47688, n47689, n47690, n47691, n47692, n47693,
    n47694, n47695, n47696, n47697, n47698, n47699,
    n47700, n47701, n47702, n47703, n47704, n47705,
    n47706, n47707, n47708, n47709, n47710, n47711,
    n47712, n47713, n47714, n47715, n47716, n47717,
    n47718, n47719, n47720, n47721, n47722, n47723,
    n47724, n47725, n47726, n47727, n47728, n47729,
    n47730, n47731, n47732, n47733, n47734, n47735,
    n47736, n47737, n47738, n47739, n47740, n47741,
    n47742, n47743, n47744, n47745, n47746, n47747,
    n47748, n47749, n47750, n47751, n47752, n47753,
    n47754, n47755, n47756, n47757, n47758, n47759,
    n47760, n47761, n47762, n47763, n47764, n47765,
    n47766, n47767, n47768, n47769, n47770, n47771,
    n47772, n47773, n47774, n47775, n47776, n47777,
    n47778, n47779, n47780, n47781, n47782, n47783,
    n47784, n47785, n47786, n47787, n47788, n47789,
    n47790, n47791, n47792, n47793, n47794, n47795,
    n47796, n47797, n47798, n47799, n47800, n47801,
    n47802, n47803, n47804, n47805, n47806, n47807,
    n47808, n47809, n47810, n47811, n47812, n47813,
    n47814, n47815, n47816, n47817, n47818, n47819,
    n47820, n47821, n47822, n47823, n47824, n47825,
    n47826, n47827, n47828, n47829, n47830, n47831,
    n47832, n47833, n47834, n47835, n47836, n47837,
    n47838, n47839, n47840, n47841, n47842, n47843,
    n47844, n47845, n47846, n47847, n47848, n47849,
    n47850, n47851, n47852, n47853, n47854, n47855,
    n47856, n47857, n47858, n47859, n47860, n47861,
    n47862, n47863, n47864, n47865, n47866, n47867,
    n47868, n47869, n47870, n47871, n47872, n47873,
    n47874, n47875, n47876, n47877, n47878, n47879,
    n47880, n47881, n47882, n47883, n47884, n47885,
    n47886, n47887, n47888, n47889, n47890, n47891,
    n47892, n47893, n47894, n47895, n47896, n47897,
    n47898, n47899, n47900, n47901, n47902, n47903,
    n47904, n47905, n47906, n47907, n47908, n47909,
    n47910, n47911, n47912, n47913, n47914, n47915,
    n47916, n47917, n47918, n47919, n47920, n47921,
    n47922, n47923, n47924, n47925, n47926, n47927,
    n47928, n47929, n47930, n47931, n47932, n47933,
    n47934, n47935, n47936, n47937, n47938, n47939,
    n47940, n47941, n47942, n47943, n47944, n47945,
    n47946, n47947, n47948, n47949, n47950, n47951,
    n47952, n47953, n47954, n47955, n47956, n47957,
    n47958, n47959, n47960, n47961, n47962, n47963,
    n47964, n47965, n47966, n47967, n47968, n47969,
    n47970, n47971, n47972, n47973, n47974, n47975,
    n47976, n47977, n47978, n47979, n47980, n47981,
    n47982, n47983, n47984, n47985, n47986, n47987,
    n47988, n47989, n47990, n47991, n47992, n47993,
    n47994, n47995, n47996, n47997, n47998, n47999,
    n48000, n48001, n48002, n48003, n48004, n48005,
    n48006, n48007, n48008, n48009, n48010, n48011,
    n48012, n48013, n48014, n48015, n48016, n48017,
    n48018, n48019, n48020, n48021, n48022, n48023,
    n48024, n48025, n48026, n48027, n48028, n48029,
    n48030, n48031, n48032, n48033, n48034, n48035,
    n48036, n48037, n48038, n48039, n48040, n48041,
    n48042, n48043, n48044, n48045, n48046, n48047,
    n48048, n48049, n48050, n48051, n48052, n48053,
    n48054, n48055, n48056, n48057, n48058, n48059,
    n48060, n48061, n48062, n48063, n48064, n48065,
    n48066, n48067, n48068, n48069, n48070, n48071,
    n48072, n48073, n48074, n48075, n48076, n48077,
    n48078, n48079, n48080, n48081, n48082, n48083,
    n48084, n48085, n48086, n48087, n48088, n48089,
    n48090, n48091, n48092, n48093, n48094, n48095,
    n48096, n48097, n48098, n48099, n48100, n48101,
    n48102, n48103, n48104, n48105, n48106, n48107,
    n48108, n48109, n48110, n48111, n48112, n48113,
    n48114, n48115, n48116, n48117, n48118, n48119,
    n48120, n48121, n48122, n48123, n48124, n48125,
    n48126, n48127, n48128, n48129, n48130, n48131,
    n48132, n48133, n48134, n48135, n48136, n48137,
    n48138, n48139, n48140, n48141, n48142, n48143,
    n48144, n48145, n48146, n48147, n48148, n48149,
    n48150, n48151, n48152, n48153, n48154, n48155,
    n48156, n48157, n48158, n48159, n48160, n48161,
    n48162, n48163, n48164, n48165, n48166, n48167,
    n48168, n48169, n48170, n48171, n48172, n48173,
    n48174, n48175, n48176, n48177, n48178, n48179,
    n48180, n48181, n48182, n48183, n48184, n48185,
    n48186, n48187, n48188, n48189, n48190, n48191,
    n48192, n48193, n48194, n48195, n48196, n48197,
    n48198, n48199, n48200, n48201, n48203, n48204,
    n48205, n48206, n48207, n48208, n48209, n48210,
    n48211, n48212, n48213, n48214, n48215, n48216,
    n48217, n48218, n48219, n48220, n48221, n48222,
    n48223, n48224, n48225, n48226, n48227, n48228,
    n48229, n48230, n48231, n48232, n48233, n48234,
    n48235, n48236, n48237, n48238, n48239, n48240,
    n48241, n48242, n48243, n48244, n48245, n48246,
    n48247, n48248, n48249, n48250, n48251, n48252,
    n48253, n48254, n48255, n48256, n48257, n48258,
    n48259, n48260, n48261, n48262, n48263, n48264,
    n48265, n48266, n48267, n48268, n48269, n48270,
    n48271, n48272, n48273, n48274, n48275, n48276,
    n48277, n48278, n48279, n48280, n48281, n48282,
    n48283, n48284, n48285, n48286, n48287, n48288,
    n48289, n48290, n48291, n48292, n48293, n48294,
    n48295, n48296, n48297, n48298, n48299, n48300,
    n48301, n48302, n48303, n48304, n48305, n48306,
    n48307, n48308, n48309, n48310, n48311, n48312,
    n48313, n48314, n48315, n48316, n48317, n48318,
    n48319, n48320, n48321, n48322, n48323, n48324,
    n48325, n48326, n48327, n48328, n48329, n48330,
    n48331, n48332, n48333, n48334, n48335, n48336,
    n48337, n48338, n48339, n48340, n48341, n48342,
    n48343, n48344, n48345, n48346, n48347, n48348,
    n48349, n48350, n48351, n48352, n48353, n48354,
    n48355, n48356, n48357, n48358, n48359, n48360,
    n48361, n48362, n48363, n48364, n48365, n48366,
    n48367, n48368, n48369, n48370, n48371, n48372,
    n48373, n48374, n48375, n48376, n48377, n48378,
    n48379, n48380, n48381, n48382, n48383, n48384,
    n48385, n48386, n48387, n48388, n48389, n48390,
    n48391, n48392, n48393, n48394, n48395, n48396,
    n48397, n48398, n48399, n48400, n48401, n48402,
    n48403, n48404, n48405, n48406, n48407, n48408,
    n48409, n48410, n48411, n48412, n48413, n48414,
    n48415, n48416, n48417, n48418, n48419, n48420,
    n48421, n48422, n48423, n48424, n48425, n48426,
    n48427, n48429, n48430, n48431, n48432, n48433,
    n48434, n48435, n48436, n48437, n48438, n48439,
    n48440, n48441, n48442, n48443, n48444, n48445,
    n48446, n48447, n48448, n48449, n48450, n48451,
    n48452, n48453, n48454, n48455, n48456, n48457,
    n48458, n48459, n48460, n48461, n48462, n48463,
    n48464, n48465, n48466, n48467, n48468, n48469,
    n48470, n48471, n48472, n48473, n48474, n48475,
    n48476, n48477, n48478, n48479, n48480, n48481,
    n48482, n48483, n48484, n48485, n48486, n48487,
    n48488, n48489, n48490, n48491, n48492, n48493,
    n48494, n48495, n48496, n48497, n48498, n48499,
    n48500, n48501, n48502, n48503, n48504, n48505,
    n48506, n48507, n48508, n48509, n48510, n48511,
    n48512, n48513, n48514, n48515, n48517, n48518,
    n48519, n48520, n48521, n48522, n48523, n48524,
    n48525, n48526, n48527, n48528, n48529, n48530,
    n48531, n48532, n48533, n48534, n48535, n48536,
    n48537, n48538, n48539, n48540, n48541, n48542,
    n48543, n48544, n48545, n48546, n48547, n48548,
    n48549, n48550, n48551, n48552, n48553, n48554,
    n48555, n48556, n48557, n48558, n48559, n48560,
    n48561, n48562, n48563, n48564, n48565, n48566,
    n48567, n48568, n48569, n48570, n48571, n48572,
    n48573, n48574, n48575, n48576, n48577, n48578,
    n48579, n48580, n48581, n48582, n48583, n48584,
    n48585, n48586, n48587, n48588, n48589, n48590,
    n48591, n48592, n48593, n48594, n48595, n48596,
    n48597, n48598, n48599, n48600, n48601, n48602,
    n48603, n48604, n48605, n48606, n48607, n48608,
    n48609, n48610, n48611, n48612, n48613, n48614,
    n48615, n48616, n48617, n48618, n48619, n48620,
    n48621, n48622, n48623, n48624, n48625, n48626,
    n48627, n48628, n48629, n48630, n48631, n48632,
    n48633, n48634, n48635, n48636, n48637, n48638,
    n48639, n48640, n48641, n48642, n48643, n48644,
    n48645, n48646, n48647, n48648, n48649, n48650,
    n48651, n48652, n48653, n48654, n48655, n48656,
    n48657, n48658, n48659, n48660, n48661, n48662,
    n48663, n48664, n48665, n48666, n48667, n48668,
    n48669, n48670, n48671, n48672, n48673, n48674,
    n48675, n48676, n48677, n48678, n48679, n48680,
    n48681, n48682, n48683, n48684, n48685, n48686,
    n48687, n48688, n48689, n48690, n48691, n48692,
    n48693, n48694, n48695, n48696, n48697, n48698,
    n48699, n48700, n48701, n48702, n48703, n48704,
    n48705, n48706, n48707, n48708, n48709, n48710,
    n48711, n48712, n48713, n48714, n48715, n48716,
    n48717, n48718, n48719, n48720, n48721, n48722,
    n48723, n48724, n48725, n48726, n48727, n48728,
    n48729, n48730, n48731, n48732, n48733, n48734,
    n48735, n48736, n48737, n48738, n48739, n48740,
    n48741, n48742, n48743, n48744, n48745, n48746,
    n48747, n48748, n48749, n48750, n48751, n48752,
    n48753, n48754, n48755, n48756, n48757, n48758,
    n48759, n48760, n48761, n48762, n48763, n48764,
    n48765, n48766, n48767, n48768, n48769, n48770,
    n48771, n48772, n48773, n48774, n48775, n48776,
    n48777, n48778, n48779, n48780, n48781, n48782,
    n48783, n48784, n48785, n48786, n48787, n48788,
    n48789, n48790, n48791, n48792, n48793, n48794,
    n48795, n48796, n48797, n48798, n48799, n48800,
    n48801, n48802, n48803, n48804, n48805, n48806,
    n48807, n48808, n48809, n48810, n48811, n48812,
    n48813, n48814, n48815, n48816, n48817, n48818,
    n48819, n48820, n48821, n48822, n48823, n48824,
    n48825, n48826, n48827, n48828, n48829, n48830,
    n48831, n48832, n48833, n48834, n48835, n48836,
    n48837, n48838, n48839, n48840, n48841, n48842,
    n48843, n48844, n48845, n48846, n48847, n48848,
    n48849, n48850, n48851, n48852, n48853, n48854,
    n48855, n48856, n48857, n48858, n48859, n48860,
    n48861, n48862, n48863, n48864, n48865, n48866,
    n48867, n48868, n48869, n48870, n48871, n48872,
    n48873, n48874, n48875, n48876, n48877, n48878,
    n48879, n48880, n48881, n48882, n48883, n48884,
    n48885, n48886, n48887, n48888, n48889, n48890,
    n48891, n48892, n48893, n48894, n48895, n48896,
    n48897, n48898, n48899, n48900, n48901, n48902,
    n48903, n48904, n48905, n48906, n48907, n48908,
    n48909, n48910, n48911, n48912, n48913, n48914,
    n48915, n48916, n48917, n48918, n48919, n48920,
    n48921, n48922, n48923, n48924, n48925, n48926,
    n48927, n48928, n48929, n48930, n48931, n48932,
    n48933, n48934, n48935, n48936, n48937, n48938,
    n48939, n48940, n48941, n48942, n48943, n48944,
    n48945, n48946, n48947, n48948, n48949, n48950,
    n48951, n48952, n48953, n48954, n48955, n48956,
    n48957, n48958, n48959, n48960, n48961, n48962,
    n48963, n48964, n48965, n48966, n48967, n48968,
    n48969, n48970, n48971, n48972, n48973, n48974,
    n48975, n48976, n48977, n48978, n48979, n48980,
    n48981, n48982, n48983, n48984, n48985, n48986,
    n48987, n48988, n48989, n48990, n48991, n48992,
    n48993, n48994, n48995, n48996, n48997, n48998,
    n48999, n49000, n49001, n49002, n49003, n49004,
    n49005, n49006, n49007, n49008, n49009, n49010,
    n49011, n49012, n49013, n49014, n49015, n49016,
    n49017, n49018, n49019, n49020, n49021, n49022,
    n49023, n49024, n49025, n49026, n49027, n49028,
    n49029, n49030, n49031, n49032, n49033, n49034,
    n49035, n49036, n49037, n49038, n49039, n49040,
    n49041, n49042, n49043, n49044, n49045, n49046,
    n49047, n49048, n49049, n49050, n49051, n49052,
    n49053, n49054, n49055, n49056, n49057, n49058,
    n49059, n49060, n49061, n49062, n49063, n49064,
    n49065, n49066, n49067, n49068, n49069, n49070,
    n49071, n49072, n49073, n49074, n49075, n49076,
    n49077, n49078, n49079, n49080, n49081, n49082,
    n49083, n49084, n49085, n49086, n49087, n49088,
    n49089, n49090, n49091, n49092, n49093, n49094,
    n49095, n49096, n49097, n49098, n49099, n49100,
    n49101, n49102, n49103, n49104, n49105, n49106,
    n49107, n49108, n49109, n49110, n49111, n49112,
    n49113, n49114, n49115, n49116, n49117, n49118,
    n49119, n49120, n49121, n49122, n49123, n49124,
    n49125, n49126, n49127, n49128, n49129, n49130,
    n49131, n49132, n49133, n49134, n49135, n49136,
    n49137, n49138, n49140, n49141, n49142, n49143,
    n49144, n49145, n49146, n49147, n49148, n49149,
    n49150, n49151, n49152, n49153, n49154, n49155,
    n49156, n49157, n49158, n49159, n49160, n49161,
    n49162, n49163, n49164, n49165, n49166, n49167,
    n49168, n49169, n49170, n49171, n49172, n49173,
    n49174, n49175, n49176, n49177, n49178, n49179,
    n49180, n49181, n49182, n49183, n49184, n49185,
    n49186, n49187, n49188, n49189, n49190, n49191,
    n49192, n49193, n49194, n49195, n49196, n49197,
    n49198, n49199, n49200, n49201, n49202, n49203,
    n49204, n49205, n49206, n49207, n49208, n49209,
    n49210, n49211, n49212, n49213, n49214, n49215,
    n49216, n49217, n49218, n49219, n49220, n49221,
    n49222, n49223, n49224, n49225, n49226, n49227,
    n49228, n49229, n49230, n49231, n49232, n49233,
    n49234, n49235, n49236, n49237, n49238, n49239,
    n49240, n49241, n49242, n49243, n49244, n49245,
    n49246, n49247, n49248, n49249, n49250, n49251,
    n49252, n49253, n49254, n49255, n49256, n49257,
    n49258, n49259, n49260, n49261, n49262, n49263,
    n49264, n49265, n49266, n49267, n49268, n49269,
    n49270, n49271, n49272, n49273, n49274, n49275,
    n49276, n49277, n49278, n49279, n49280, n49281,
    n49282, n49283, n49284, n49285, n49286, n49287,
    n49288, n49289, n49290, n49291, n49292, n49293,
    n49294, n49295, n49296, n49297, n49298, n49299,
    n49300, n49301, n49302, n49303, n49304, n49305,
    n49306, n49307, n49308, n49309, n49310, n49311,
    n49312, n49313, n49314, n49315, n49316, n49317,
    n49318, n49319, n49320, n49321, n49322, n49323,
    n49324, n49325, n49326, n49327, n49328, n49329,
    n49330, n49331, n49332, n49333, n49334, n49335,
    n49336, n49337, n49338, n49339, n49340, n49343,
    n49344, n49345, n49346, n49347, n49348, n49349,
    n49350, n49351, n49352, n49353, n49354, n49355,
    n49356, n49357, n49358, n49359, n49360, n49361,
    n49362, n49363, n49364, n49365, n49366, n49367,
    n49368, n49369, n49370, n49371, n49372, n49373,
    n49374, n49375, n49376, n49377, n49378, n49379,
    n49380, n49381, n49382, n49383, n49384, n49385,
    n49386, n49387, n49388, n49389, n49390, n49391,
    n49392, n49393, n49394, n49395, n49396, n49397,
    n49398, n49399, n49400, n49401, n49402, n49403,
    n49404, n49405, n49406, n49407, n49408, n49409,
    n49410, n49411, n49412, n49413, n49414, n49415,
    n49416, n49417, n49418, n49419, n49420, n49421,
    n49422, n49423, n49424, n49425, n49426, n49427,
    n49428, n49429, n49430, n49431, n49432, n49433,
    n49434, n49435, n49436, n49437, n49438, n49439,
    n49440, n49441, n49442, n49443, n49444, n49445,
    n49446, n49447, n49448, n49449, n49450, n49451,
    n49452, n49453, n49454, n49455, n49456, n49457,
    n49458, n49459, n49460, n49461, n49462, n49463,
    n49464, n49465, n49466, n49467, n49468, n49469,
    n49470, n49471, n49472, n49473, n49474, n49475,
    n49476, n49477, n49478, n49479, n49480, n49481,
    n49482, n49483, n49484, n49485, n49486, n49487,
    n49488, n49489, n49490, n49491, n49492, n49493,
    n49494, n49495, n49496, n49497, n49498, n49499,
    n49500, n49501, n49502, n49503, n49504, n49505,
    n49506, n49507, n49508, n49509, n49510, n49511,
    n49512, n49513, n49514, n49515, n49516, n49517,
    n49518, n49519, n49520, n49521, n49522, n49523,
    n49524, n49525, n49526, n49527, n49528, n49529,
    n49530, n49531, n49532, n49533, n49534, n49535,
    n49536, n49537, n49538, n49539, n49540, n49541,
    n49542, n49543, n49544, n49545, n49546, n49547,
    n49548, n49549, n49550, n49551, n49552, n49553,
    n49554, n49555, n49556, n49557, n49558, n49559,
    n49560, n49561, n49562, n49563, n49564, n49565,
    n49566, n49567, n49568, n49569, n49570, n49571,
    n49572, n49573, n49574, n49575, n49576, n49577,
    n49578, n49579, n49580, n49581, n49582, n49583,
    n49584, n49585, n49586, n49587, n49588, n49589,
    n49590, n49591, n49592, n49593, n49594, n49595,
    n49596, n49597, n49598, n49599, n49600, n49601,
    n49602, n49603, n49604, n49605, n49606, n49607,
    n49608, n49609, n49610, n49611, n49612, n49613,
    n49614, n49615, n49616, n49617, n49618, n49619,
    n49620, n49621, n49622, n49623, n49624, n49625,
    n49626, n49627, n49628, n49629, n49630, n49631,
    n49632, n49633, n49634, n49635, n49636, n49637,
    n49638, n49639, n49640, n49641, n49642, n49643,
    n49644, n49645, n49646, n49647, n49648, n49649,
    n49650, n49651, n49652, n49653, n49654, n49655,
    n49656, n49657, n49658, n49659, n49660, n49661,
    n49662, n49663, n49664, n49665, n49666, n49667,
    n49668, n49669, n49670, n49671, n49672, n49673,
    n49674, n49675, n49676, n49677, n49678, n49679,
    n49680, n49681, n49682, n49683, n49684, n49685,
    n49686, n49687, n49688, n49689, n49690, n49691,
    n49692, n49693, n49694, n49695, n49696, n49697,
    n49698, n49699, n49700, n49701, n49702, n49703,
    n49704, n49705, n49706, n49707, n49708, n49709,
    n49710, n49711, n49712, n49713, n49714, n49715,
    n49716, n49717, n49718, n49719, n49720, n49721,
    n49722, n49723, n49724, n49725, n49726, n49727,
    n49728, n49729, n49730, n49731, n49732, n49733,
    n49734, n49735, n49736, n49737, n49738, n49739,
    n49740, n49741, n49742, n49743, n49744, n49745,
    n49746, n49747, n49748, n49749, n49750, n49751,
    n49752, n49753, n49754, n49755, n49756, n49757,
    n49758, n49759, n49760, n49761, n49762, n49763,
    n49764, n49765, n49766, n49767, n49768, n49769,
    n49770, n49771, n49772, n49773, n49774, n49775,
    n49776, n49777, n49778, n49779, n49780, n49781,
    n49782, n49783, n49784, n49785, n49786, n49787,
    n49788, n49789, n49790, n49791, n49792, n49793,
    n49794, n49795, n49796, n49797, n49798, n49799,
    n49800, n49801, n49802, n49803, n49804, n49805,
    n49806, n49807, n49808, n49809, n49810, n49811,
    n49812, n49813, n49814, n49815, n49816, n49817,
    n49818, n49819, n49820, n49821, n49822, n49823,
    n49824, n49825, n49826, n49827, n49828, n49829,
    n49830, n49831, n49832, n49833, n49834, n49835,
    n49836, n49837, n49838, n49839, n49840, n49841,
    n49842, n49843, n49844, n49845, n49846, n49847,
    n49848, n49849, n49850, n49851, n49852, n49853,
    n49854, n49855, n49856, n49857, n49858, n49859,
    n49860, n49861, n49862, n49863, n49864, n49865,
    n49866, n49867, n49868, n49869, n49870, n49871,
    n49872, n49873, n49874, n49875, n49876, n49877,
    n49878, n49879, n49880, n49881, n49882, n49883,
    n49884, n49885, n49886, n49887, n49888, n49889,
    n49890, n49891, n49892, n49893, n49894, n49895,
    n49896, n49897, n49898, n49899, n49900, n49901,
    n49902, n49903, n49904, n49905, n49906, n49907,
    n49908, n49909, n49910, n49911, n49912, n49913,
    n49914, n49915, n49916, n49917, n49918, n49919,
    n49920, n49921, n49922, n49923, n49924, n49925,
    n49926, n49927, n49928, n49929, n49930, n49931,
    n49932, n49933, n49934, n49935, n49936, n49937,
    n49938, n49939, n49940, n49941, n49942, n49943,
    n49944, n49945, n49946, n49947, n49948, n49949,
    n49950, n49951, n49952, n49953, n49954, n49955,
    n49956, n49957, n49958, n49959, n49960, n49961,
    n49962, n49963, n49964, n49965, n49966, n49967,
    n49968, n49969, n49970, n49971, n49972, n49973,
    n49974, n49975, n49976, n49977, n49978, n49979,
    n49980, n49981, n49982, n49983, n49984, n49985,
    n49986, n49987, n49988, n49989, n49990, n49991,
    n49992, n49993, n49994, n49995, n49996, n49997,
    n49998, n49999, n50000, n50001, n50002, n50003,
    n50004, n50005, n50006, n50007, n50008, n50009,
    n50010, n50011, n50012, n50013, n50014, n50015,
    n50016, n50017, n50018, n50019, n50020, n50021,
    n50022, n50023, n50024, n50025, n50026, n50027,
    n50028, n50029, n50030, n50031, n50032, n50033,
    n50034, n50035, n50036, n50037, n50038, n50039,
    n50040, n50041, n50042, n50043, n50044, n50045,
    n50046, n50047, n50048, n50049, n50050, n50051,
    n50052, n50053, n50054, n50055, n50056, n50057,
    n50058, n50059, n50060, n50061, n50062, n50063,
    n50064, n50065, n50066, n50067, n50068, n50069,
    n50070, n50071, n50072, n50073, n50074, n50075,
    n50076, n50077, n50078, n50079, n50080, n50081,
    n50082, n50083, n50084, n50085, n50086, n50087,
    n50088, n50089, n50090, n50091, n50092, n50093,
    n50094, n50095, n50096, n50097, n50098, n50099,
    n50100, n50101, n50102, n50103, n50104, n50105,
    n50106, n50107, n50108, n50109, n50110, n50111,
    n50112, n50113, n50114, n50115, n50116, n50117,
    n50118, n50119, n50120, n50121, n50122, n50123,
    n50124, n50125, n50126, n50127, n50128, n50129,
    n50130, n50131, n50132, n50133, n50134, n50135,
    n50136, n50137, n50138, n50139, n50140, n50141,
    n50142, n50143, n50144, n50145, n50146, n50147,
    n50148, n50149, n50150, n50151, n50152, n50153,
    n50154, n50155, n50156, n50157, n50158, n50159,
    n50160, n50161, n50162, n50163, n50164, n50165,
    n50166, n50167, n50168, n50169, n50170, n50171,
    n50172, n50173, n50174, n50175, n50176, n50177,
    n50178, n50179, n50180, n50181, n50182, n50183,
    n50184, n50185, n50186, n50187, n50188, n50189,
    n50190, n50191, n50192, n50193, n50194, n50195,
    n50196, n50197, n50198, n50199, n50200, n50201,
    n50202, n50203, n50204, n50205, n50206, n50207,
    n50208, n50209, n50210, n50211, n50212, n50213,
    n50214, n50215, n50216, n50217, n50218, n50219,
    n50220, n50221, n50222, n50223, n50224, n50225,
    n50226, n50227, n50228, n50229, n50230, n50231,
    n50232, n50233, n50234, n50235, n50236, n50237,
    n50238, n50239, n50240, n50241, n50242, n50243,
    n50244, n50245, n50246, n50247, n50248, n50249,
    n50250, n50251, n50252, n50253, n50254, n50255,
    n50256, n50257, n50258, n50259, n50260, n50261,
    n50262, n50263, n50264, n50265, n50266, n50267,
    n50268, n50269, n50270, n50271, n50272, n50273,
    n50274, n50275, n50276, n50277, n50278, n50279,
    n50280, n50281, n50282, n50283, n50284, n50285,
    n50286, n50287, n50288, n50289, n50290, n50291,
    n50292, n50293, n50294, n50295, n50296, n50297,
    n50298, n50299, n50300, n50301, n50302, n50303,
    n50304, n50305, n50306, n50307, n50308, n50309,
    n50310, n50311, n50312, n50313, n50314, n50315,
    n50316, n50317, n50318, n50319, n50320, n50321,
    n50322, n50323, n50324, n50325, n50326, n50327,
    n50328, n50329, n50330, n50331, n50332, n50333,
    n50334, n50335, n50336, n50337, n50338, n50339,
    n50340, n50341, n50342, n50343, n50344, n50345,
    n50346, n50347, n50348, n50349, n50350, n50351,
    n50352, n50353, n50354, n50355, n50356, n50357,
    n50358, n50359, n50360, n50361, n50362, n50363,
    n50364, n50365, n50366, n50367, n50368, n50369,
    n50370, n50371, n50372, n50373, n50374, n50375,
    n50376, n50377, n50378, n50379, n50380, n50382,
    n50383, n50384, n50385, n50386, n50387, n50388,
    n50389, n50390, n50391, n50392, n50393, n50394,
    n50395, n50396, n50397, n50398, n50399, n50400,
    n50401, n50402, n50403, n50404, n50405, n50406,
    n50407, n50408, n50409, n50410, n50411, n50412,
    n50413, n50414, n50415, n50416, n50417, n50418,
    n50419, n50420, n50421, n50422, n50423, n50424,
    n50425, n50426, n50427, n50428, n50429, n50430,
    n50431, n50432, n50433, n50434, n50435, n50436,
    n50437, n50438, n50439, n50440, n50441, n50442,
    n50443, n50444, n50445, n50446, n50447, n50448,
    n50449, n50450, n50451, n50452, n50453, n50454,
    n50455, n50456, n50457, n50458, n50459, n50460,
    n50461, n50462, n50463, n50464, n50465, n50466,
    n50467, n50468, n50469, n50470, n50471, n50473,
    n50474, n50475, n50476, n50477, n50478, n50479,
    n50480, n50481, n50482, n50483, n50484, n50485,
    n50486, n50487, n50488, n50489, n50490, n50491,
    n50492, n50493, n50494, n50495, n50496, n50497,
    n50498, n50499, n50500, n50501, n50502, n50503,
    n50504, n50505, n50506, n50507, n50508, n50509,
    n50510, n50511, n50512, n50513, n50514, n50515,
    n50516, n50517, n50518, n50519, n50520, n50521,
    n50522, n50523, n50524, n50525, n50526, n50527,
    n50528, n50529, n50530, n50531, n50532, n50533,
    n50534, n50535, n50536, n50537, n50538, n50539,
    n50540, n50541, n50542, n50543, n50544, n50545,
    n50546, n50547, n50548, n50549, n50550, n50551,
    n50552, n50553, n50554, n50555, n50556, n50557,
    n50558, n50559, n50560, n50561, n50562, n50563,
    n50564, n50565, n50566, n50567, n50568, n50569,
    n50570, n50571, n50572, n50573, n50574, n50575,
    n50576, n50577, n50578, n50579, n50580, n50581,
    n50582, n50583, n50584, n50585, n50586, n50587,
    n50588, n50589, n50590, n50591, n50592, n50593,
    n50594, n50595, n50596, n50597, n50598, n50599,
    n50600, n50601, n50602, n50603, n50604, n50605,
    n50606, n50607, n50608, n50609, n50610, n50611,
    n50612, n50613, n50614, n50615, n50616, n50617,
    n50618, n50619, n50620, n50621, n50622, n50623,
    n50624, n50625, n50626, n50627, n50628, n50629,
    n50630, n50631, n50632, n50633, n50634, n50635,
    n50636, n50637, n50638, n50639, n50640, n50641,
    n50642, n50643, n50644, n50645, n50646, n50647,
    n50648, n50649, n50650, n50651, n50652, n50653,
    n50654, n50655, n50656, n50657, n50658, n50659,
    n50660, n50661, n50662, n50663, n50664, n50665,
    n50666, n50667, n50668, n50669, n50670, n50671,
    n50672, n50673, n50674, n50675, n50676, n50677,
    n50678, n50679, n50680, n50681, n50682, n50683,
    n50684, n50685, n50686, n50687, n50688, n50689,
    n50690, n50691, n50692, n50693, n50694, n50695,
    n50696, n50697, n50698, n50699, n50700, n50701,
    n50702, n50703, n50704, n50705, n50706, n50707,
    n50708, n50709, n50710, n50711, n50712, n50713,
    n50714, n50715, n50716, n50717, n50718, n50719,
    n50720, n50721, n50722, n50723, n50724, n50725,
    n50726, n50727, n50728, n50729, n50730, n50731,
    n50732, n50733, n50734, n50735, n50736, n50737,
    n50738, n50739, n50740, n50741, n50742, n50743,
    n50744, n50745, n50746, n50747, n50748, n50749,
    n50750, n50751, n50752, n50753, n50754, n50755,
    n50756, n50757, n50758, n50759, n50760, n50761,
    n50762, n50763, n50764, n50765, n50766, n50767,
    n50768, n50769, n50770, n50771, n50772, n50773,
    n50774, n50775, n50776, n50777, n50778, n50779,
    n50780, n50781, n50782, n50783, n50784, n50785,
    n50786, n50787, n50788, n50789, n50790, n50791,
    n50792, n50793, n50794, n50795, n50796, n50797,
    n50798, n50799, n50800, n50801, n50802, n50803,
    n50804, n50805, n50806, n50807, n50808, n50809,
    n50810, n50811, n50812, n50813, n50814, n50815,
    n50816, n50817, n50818, n50819, n50820, n50821,
    n50822, n50823, n50824, n50825, n50826, n50827,
    n50828, n50829, n50830, n50831, n50832, n50833,
    n50834, n50835, n50836, n50837, n50838, n50839,
    n50840, n50841, n50842, n50843, n50844, n50845,
    n50846, n50847, n50848, n50849, n50850, n50851,
    n50852, n50853, n50854, n50855, n50856, n50857,
    n50858, n50859, n50860, n50861, n50862, n50863,
    n50864, n50865, n50866, n50867, n50868, n50869,
    n50870, n50871, n50872, n50873, n50874, n50875,
    n50876, n50877, n50878, n50879, n50880, n50881,
    n50882, n50883, n50884, n50885, n50886, n50887,
    n50888, n50889, n50890, n50891, n50892, n50893,
    n50894, n50895, n50896, n50897, n50898, n50899,
    n50900, n50901, n50902, n50903, n50904, n50905,
    n50906, n50907, n50908, n50909, n50910, n50911,
    n50912, n50913, n50914, n50915, n50916, n50917,
    n50918, n50919, n50920, n50921, n50922, n50923,
    n50924, n50925, n50926, n50927, n50928, n50929,
    n50930, n50931, n50932, n50933, n50934, n50935,
    n50936, n50937, n50938, n50939, n50940, n50941,
    n50942, n50943, n50944, n50945, n50946, n50947,
    n50948, n50949, n50950, n50951, n50952, n50953,
    n50954, n50955, n50956, n50957, n50958, n50959,
    n50960, n50961, n50962, n50963, n50964, n50965,
    n50966, n50967, n50968, n50969, n50970, n50971,
    n50972, n50973, n50974, n50975, n50976, n50977,
    n50978, n50979, n50980, n50981, n50982, n50983,
    n50984, n50985, n50986, n50987, n50988, n50989,
    n50990, n50991, n50992, n50993, n50994, n50995,
    n50996, n50997, n50998, n50999, n51000, n51002,
    n51003, n51004, n51005, n51006, n51007, n51008,
    n51009, n51010, n51011, n51012, n51013, n51014,
    n51015, n51016, n51017, n51018, n51019, n51020,
    n51021, n51022, n51023, n51024, n51025, n51026,
    n51027, n51028, n51029, n51030, n51031, n51032,
    n51033, n51034, n51035, n51036, n51037, n51038,
    n51039, n51040, n51041, n51042, n51043, n51044,
    n51045, n51046, n51047, n51048, n51049, n51050,
    n51051, n51052, n51053, n51054, n51055, n51056,
    n51057, n51058, n51059, n51060, n51061, n51062,
    n51063, n51064, n51065, n51066, n51067, n51068,
    n51069, n51070, n51071, n51072, n51073, n51074,
    n51075, n51076, n51077, n51078, n51079, n51080,
    n51081, n51082, n51083, n51084, n51085, n51086,
    n51087, n51088, n51089, n51090, n51091, n51092,
    n51093, n51094, n51095, n51096, n51097, n51098,
    n51099, n51100, n51101, n51102, n51103, n51104,
    n51105, n51106, n51107, n51108, n51109, n51110,
    n51111, n51112, n51113, n51114, n51115, n51116,
    n51117, n51118, n51119, n51120, n51121, n51122,
    n51123, n51124, n51125, n51126, n51127, n51128,
    n51129, n51130, n51131, n51132, n51133, n51134,
    n51135, n51136, n51137, n51138, n51139, n51140,
    n51141, n51142, n51143, n51144, n51145, n51146,
    n51147, n51148, n51149, n51150, n51151, n51152,
    n51153, n51154, n51155, n51156, n51157, n51158,
    n51159, n51160, n51161, n51162, n51163, n51164,
    n51165, n51166, n51167, n51168, n51169, n51170,
    n51171, n51172, n51173, n51174, n51175, n51176,
    n51177, n51178, n51179, n51180, n51181, n51182,
    n51183, n51184, n51185, n51186, n51187, n51188,
    n51189, n51190, n51191, n51192, n51193, n51194,
    n51195, n51196, n51197, n51198, n51199, n51200,
    n51201, n51202, n51203, n51204, n51205, n51206,
    n51207, n51208, n51209, n51210, n51211, n51212,
    n51213, n51214, n51215, n51216, n51217, n51218,
    n51219, n51220, n51221, n51222, n51223, n51224,
    n51225, n51226, n51227, n51228, n51229, n51230,
    n51231, n51232, n51233, n51234, n51235, n51236,
    n51237, n51238, n51239, n51240, n51241, n51242,
    n51243, n51244, n51245, n51246, n51247, n51248,
    n51249, n51250, n51251, n51252, n51253, n51254,
    n51255, n51256, n51257, n51258, n51259, n51260,
    n51261, n51262, n51263, n51264, n51265, n51266,
    n51267, n51268, n51269, n51270, n51271, n51272,
    n51273, n51274, n51275, n51276, n51277, n51278,
    n51279, n51280, n51281, n51282, n51283, n51284,
    n51285, n51286, n51287, n51288, n51289, n51290,
    n51291, n51292, n51293, n51294, n51295, n51296,
    n51297, n51298, n51299, n51300, n51301, n51302,
    n51303, n51304, n51305, n51306, n51307, n51308,
    n51309, n51310, n51311, n51312, n51313, n51314,
    n51315, n51316, n51317, n51318, n51319, n51320,
    n51321, n51322, n51323, n51324, n51325, n51326,
    n51327, n51328, n51329, n51330, n51331, n51332,
    n51333, n51334, n51335, n51336, n51337, n51338,
    n51339, n51340, n51341, n51342, n51343, n51344,
    n51345, n51346, n51347, n51348, n51349, n51350,
    n51351, n51352, n51353, n51354, n51355, n51356,
    n51357, n51358, n51359, n51360, n51361, n51362,
    n51363, n51364, n51365, n51366, n51367, n51368,
    n51369, n51370, n51371, n51372, n51373, n51374,
    n51375, n51376, n51377, n51378, n51379, n51380,
    n51381, n51382, n51383, n51384, n51385, n51386,
    n51387, n51388, n51389, n51390, n51391, n51392,
    n51393, n51394, n51395, n51396, n51397, n51398,
    n51399, n51400, n51401, n51402, n51403, n51404,
    n51405, n51406, n51407, n51408, n51409, n51410,
    n51411, n51412, n51413, n51414, n51415, n51416,
    n51417, n51418, n51419, n51420, n51421, n51422,
    n51423, n51424, n51425, n51426, n51427, n51428,
    n51429, n51430, n51431, n51432, n51433, n51434,
    n51435, n51436, n51437, n51438, n51439, n51440,
    n51441, n51442, n51443, n51444, n51445, n51446,
    n51447, n51448, n51449, n51450, n51451, n51452,
    n51453, n51454, n51455, n51456, n51457, n51458,
    n51459, n51460, n51461, n51462, n51463, n51464,
    n51466, n51467, n51468, n51469, n51470, n51471,
    n51472, n51473, n51474, n51475, n51476, n51477,
    n51478, n51479, n51480, n51481, n51482, n51483,
    n51484, n51485, n51486, n51487, n51488, n51489,
    n51490, n51491, n51492, n51493, n51494, n51495,
    n51496, n51497, n51498, n51499, n51500, n51501,
    n51502, n51503, n51504, n51505, n51506, n51507,
    n51508, n51509, n51510, n51511, n51512, n51513,
    n51514, n51515, n51516, n51517, n51518, n51519,
    n51520, n51521, n51522, n51523, n51524, n51525,
    n51526, n51527, n51528, n51529, n51530, n51531,
    n51532, n51533, n51534, n51535, n51536, n51537,
    n51538, n51539, n51540, n51541, n51542, n51543,
    n51544, n51545, n51546, n51547, n51548, n51549,
    n51550, n51551, n51552, n51553, n51554, n51555,
    n51556, n51557, n51558, n51559, n51560, n51561,
    n51562, n51563, n51564, n51565, n51566, n51567,
    n51568, n51569, n51570, n51571, n51572, n51573,
    n51574, n51575, n51576, n51577, n51578, n51579,
    n51580, n51581, n51582, n51583, n51584, n51585,
    n51586, n51587, n51588, n51589, n51590, n51591,
    n51592, n51593, n51594, n51595, n51596, n51597,
    n51598, n51599, n51600, n51601, n51602, n51603,
    n51604, n51605, n51606, n51607, n51608, n51609,
    n51610, n51611, n51612, n51613, n51614, n51615,
    n51616, n51617, n51618, n51619, n51620, n51621,
    n51622, n51623, n51624, n51625, n51626, n51627,
    n51628, n51629, n51630, n51631, n51632, n51633,
    n51634, n51635, n51636, n51637, n51638, n51639,
    n51640, n51641, n51642, n51643, n51644, n51645,
    n51646, n51647, n51648, n51649, n51650, n51651,
    n51652, n51653, n51654, n51655, n51656, n51657,
    n51658, n51659, n51660, n51661, n51662, n51663,
    n51664, n51665, n51666, n51667, n51668, n51669,
    n51670, n51671, n51672, n51673, n51674, n51675,
    n51676, n51677, n51678, n51679, n51680, n51681,
    n51682, n51683, n51684, n51685, n51686, n51687,
    n51688, n51689, n51690, n51691, n51692, n51693,
    n51694, n51695, n51696, n51697, n51698, n51699,
    n51700, n51701, n51702, n51703, n51704, n51705,
    n51706, n51707, n51708, n51709, n51710, n51711,
    n51712, n51713, n51714, n51715, n51716, n51717,
    n51718, n51719, n51720, n51721, n51722, n51723,
    n51724, n51725, n51726, n51727, n51728, n51729,
    n51730, n51731, n51732, n51733, n51734, n51735,
    n51736, n51737, n51738, n51739, n51740, n51741,
    n51742, n51743, n51744, n51745, n51746, n51747,
    n51748, n51749, n51750, n51751, n51752, n51753,
    n51754, n51755, n51756, n51757, n51758, n51759,
    n51760, n51761, n51762, n51763, n51764, n51765,
    n51766, n51767, n51768, n51769, n51770, n51771,
    n51772, n51773, n51774, n51775, n51776, n51777,
    n51778, n51779, n51780, n51781, n51782, n51783,
    n51784, n51785, n51786, n51787, n51788, n51789,
    n51790, n51791, n51792, n51793, n51794, n51795,
    n51796, n51797, n51798, n51799, n51800, n51801,
    n51802, n51803, n51804, n51805, n51806, n51807,
    n51808, n51809, n51810, n51811, n51812, n51813,
    n51814, n51815, n51816, n51817, n51818, n51819,
    n51820, n51821, n51822, n51823, n51824, n51825,
    n51826, n51827, n51828, n51829, n51830, n51831,
    n51832, n51833, n51834, n51835, n51836, n51837,
    n51838, n51839, n51840, n51841, n51842, n51843,
    n51844, n51845, n51846, n51847, n51848, n51849,
    n51850, n51851, n51852, n51853, n51854, n51855,
    n51856, n51857, n51858, n51859, n51860, n51861,
    n51862, n51863, n51864, n51865, n51866, n51867,
    n51868, n51869, n51870, n51871, n51872, n51873,
    n51874, n51875, n51876, n51877, n51878, n51879,
    n51880, n51881, n51882, n51883, n51884, n51885,
    n51886, n51887, n51888, n51889, n51890, n51891,
    n51892, n51893, n51894, n51895, n51896, n51897,
    n51898, n51899, n51900, n51901, n51902, n51903,
    n51904, n51905, n51906, n51907, n51908, n51909,
    n51910, n51911, n51912, n51913, n51914, n51915,
    n51916, n51917, n51918, n51919, n51920, n51921,
    n51922, n51923, n51924, n51925, n51926, n51927,
    n51928, n51929, n51930, n51931, n51932, n51933,
    n51934, n51935, n51936, n51937, n51938, n51939,
    n51940, n51941, n51942, n51943, n51944, n51945,
    n51946, n51947, n51948, n51949, n51950, n51951,
    n51952, n51953, n51954, n51955, n51956, n51957,
    n51958, n51959, n51960, n51961, n51962, n51963,
    n51964, n51965, n51966, n51967, n51968, n51969,
    n51970, n51971, n51972, n51973, n51974, n51975,
    n51976, n51977, n51978, n51979, n51980, n51981,
    n51982, n51983, n51984, n51985, n51986, n51987,
    n51988, n51989, n51990, n51991, n51992, n51993,
    n51994, n51995, n51996, n51997, n51998, n51999,
    n52000, n52001, n52002, n52003, n52004, n52005,
    n52006, n52007, n52008, n52009, n52010, n52011,
    n52012, n52013, n52014, n52015, n52016, n52017,
    n52018, n52019, n52020, n52021, n52022, n52023,
    n52024, n52025, n52026, n52027, n52028, n52029,
    n52030, n52031, n52032, n52033, n52034, n52035,
    n52036, n52037, n52038, n52039, n52040, n52041,
    n52042, n52043, n52044, n52045, n52046, n52047,
    n52048, n52049, n52050, n52051, n52052, n52053,
    n52054, n52055, n52056, n52057, n52058, n52059,
    n52060, n52061, n52062, n52063, n52064, n52065,
    n52066, n52067, n52068, n52069, n52070, n52071,
    n52072, n52073, n52074, n52075, n52076, n52077,
    n52078, n52079, n52080, n52081, n52082, n52083,
    n52084, n52085, n52086, n52087, n52088, n52089,
    n52090, n52091, n52092, n52093, n52094, n52095,
    n52096, n52097, n52098, n52099, n52100, n52101,
    n52102, n52103, n52104, n52105, n52106, n52107,
    n52108, n52109, n52110, n52111, n52112, n52113,
    n52114, n52115, n52116, n52117, n52118, n52119,
    n52120, n52121, n52122, n52123, n52124, n52125,
    n52126, n52127, n52128, n52129, n52130, n52131,
    n52132, n52133, n52134, n52135, n52136, n52137,
    n52138, n52139, n52140, n52141, n52142, n52143,
    n52144, n52145, n52146, n52147, n52148, n52149,
    n52150, n52151, n52152, n52153, n52154, n52155,
    n52156, n52157, n52158, n52159, n52160, n52161,
    n52162, n52163, n52164, n52165, n52166, n52167,
    n52168, n52169, n52170, n52171, n52172, n52173,
    n52174, n52175, n52176, n52177, n52178, n52179,
    n52180, n52181, n52182, n52183, n52184, n52185,
    n52186, n52187, n52188, n52189, n52190, n52191,
    n52192, n52193, n52194, n52195, n52196, n52197,
    n52198, n52199, n52200, n52201, n52202, n52203,
    n52204, n52205, n52206, n52207, n52208, n52209,
    n52210, n52211, n52212, n52213, n52214, n52215,
    n52216, n52217, n52218, n52219, n52220, n52221,
    n52222, n52223, n52224, n52225, n52226, n52227,
    n52228, n52229, n52230, n52231, n52232, n52233,
    n52234, n52235, n52236, n52237, n52238, n52239,
    n52240, n52241, n52242, n52243, n52244, n52245,
    n52246, n52247, n52248, n52249, n52250, n52251,
    n52252, n52253, n52254, n52255, n52256, n52257,
    n52258, n52259, n52260, n52261, n52262, n52263,
    n52264, n52265, n52266, n52267, n52268, n52269,
    n52270, n52271, n52272, n52273, n52274, n52275,
    n52276, n52277, n52278, n52279, n52280, n52281,
    n52282, n52283, n52284, n52285, n52286, n52287,
    n52288, n52289, n52290, n52291, n52292, n52293,
    n52294, n52295, n52296, n52297, n52298, n52299,
    n52300, n52301, n52302, n52303, n52304, n52305,
    n52306, n52307, n52308, n52309, n52310, n52311,
    n52312, n52313, n52314, n52315, n52316, n52317,
    n52318, n52319, n52320, n52321, n52322, n52323,
    n52324, n52325, n52326, n52327, n52328, n52329,
    n52330, n52331, n52332, n52333, n52334, n52335,
    n52336, n52337, n52338, n52339, n52340, n52341,
    n52342, n52343, n52344, n52345, n52346, n52347,
    n52348, n52349, n52350, n52351, n52352, n52353,
    n52354, n52355, n52356, n52357, n52358, n52359,
    n52360, n52361, n52362, n52363, n52364, n52365,
    n52366, n52367, n52368, n52369, n52370, n52371,
    n52372, n52373, n52374, n52375, n52376, n52377,
    n52378, n52379, n52380, n52381, n52382, n52383,
    n52384, n52385, n52386, n52387, n52388, n52389,
    n52390, n52391, n52392, n52393, n52394, n52395,
    n52396, n52397, n52398, n52399, n52400, n52401,
    n52402, n52403, n52404, n52405, n52406, n52407,
    n52408, n52409, n52410, n52411, n52412, n52413,
    n52414, n52415, n52416, n52417, n52418, n52419,
    n52420, n52421, n52422, n52423, n52424, n52425,
    n52426, n52427, n52428, n52429, n52430, n52431,
    n52432, n52433, n52434, n52436, n52437, n52438,
    n52439, n52440, n52441, n52442, n52443, n52444,
    n52445, n52446, n52447, n52448, n52449, n52450,
    n52451, n52452, n52453, n52454, n52455, n52456,
    n52457, n52458, n52459, n52460, n52461, n52462,
    n52463, n52464, n52465, n52466, n52467, n52468,
    n52469, n52470, n52471, n52472, n52473, n52474,
    n52475, n52476, n52477, n52478, n52479, n52480,
    n52481, n52482, n52483, n52484, n52485, n52486,
    n52487, n52488, n52489, n52490, n52491, n52492,
    n52493, n52494, n52495, n52496, n52497, n52499,
    n52500, n52501, n52502, n52503, n52504, n52505,
    n52506, n52507, n52508, n52509, n52510, n52511,
    n52512, n52513, n52514, n52515, n52516, n52517,
    n52518, n52519, n52520, n52521, n52522, n52523,
    n52524, n52525, n52526, n52527, n52528, n52529,
    n52530, n52531, n52532, n52533, n52534, n52535,
    n52536, n52537, n52538, n52539, n52540, n52541,
    n52542, n52543, n52544, n52545, n52546, n52547,
    n52548, n52549, n52550, n52551, n52552, n52553,
    n52554, n52555, n52556, n52557, n52558, n52559,
    n52560, n52561, n52562, n52563, n52564, n52565,
    n52566, n52567, n52568, n52569, n52570, n52571,
    n52572, n52573, n52574, n52575, n52576, n52577,
    n52578, n52579, n52580, n52581, n52582, n52583,
    n52584, n52585, n52586, n52587, n52588, n52589,
    n52590, n52591, n52592, n52593, n52594, n52595,
    n52596, n52597, n52598, n52599, n52600, n52601,
    n52602, n52603, n52604, n52605, n52606, n52607,
    n52608, n52609, n52610, n52611, n52612, n52613,
    n52614, n52615, n52616, n52617, n52618, n52619,
    n52620, n52621, n52622, n52623, n52624, n52625,
    n52626, n52627, n52628, n52629, n52630, n52631,
    n52632, n52633, n52634, n52635, n52636, n52637,
    n52638, n52639, n52640, n52641, n52642, n52643,
    n52644, n52645, n52646, n52647, n52648, n52649,
    n52650, n52651, n52652, n52653, n52654, n52655,
    n52656, n52657, n52658, n52659, n52660, n52661,
    n52662, n52663, n52664, n52665, n52666, n52667,
    n52668, n52669, n52670, n52671, n52672, n52673,
    n52674, n52675, n52676, n52677, n52678, n52679,
    n52680, n52681, n52682, n52683, n52684, n52685,
    n52686, n52687, n52688, n52689, n52690, n52691,
    n52692, n52693, n52694, n52695, n52696, n52697,
    n52698, n52699, n52700, n52701, n52702, n52703,
    n52704, n52705, n52706, n52707, n52708, n52709,
    n52710, n52711, n52712, n52713, n52714, n52715,
    n52716, n52717, n52718, n52719, n52720, n52721,
    n52722, n52723, n52724, n52725, n52726, n52727,
    n52728, n52729, n52730, n52731, n52732, n52733,
    n52734, n52735, n52736, n52737, n52738, n52739,
    n52740, n52741, n52742, n52743, n52744, n52745,
    n52746, n52747, n52748, n52749, n52750, n52751,
    n52752, n52753, n52754, n52755, n52756, n52757,
    n52758, n52759, n52760, n52761, n52762, n52763,
    n52764, n52765, n52766, n52767, n52768, n52769,
    n52770, n52771, n52772, n52773, n52774, n52775,
    n52776, n52777, n52778, n52779, n52780, n52781,
    n52782, n52783, n52784, n52785, n52786, n52787,
    n52788, n52789, n52790, n52791, n52792, n52793,
    n52794, n52795, n52796, n52797, n52798, n52799,
    n52800, n52801, n52802, n52803, n52804, n52805,
    n52806, n52807, n52808, n52809, n52810, n52811,
    n52812, n52813, n52814, n52815, n52816, n52817,
    n52818, n52819, n52820, n52821, n52822, n52823,
    n52824, n52825, n52826, n52827, n52828, n52829,
    n52830, n52831, n52832, n52833, n52834, n52835,
    n52836, n52837, n52838, n52839, n52840, n52841,
    n52842, n52843, n52844, n52845, n52846, n52847,
    n52848, n52849, n52850, n52851, n52852, n52853,
    n52854, n52855, n52856, n52857, n52858, n52859,
    n52860, n52861, n52862, n52863, n52864, n52865,
    n52866, n52867, n52868, n52869, n52870, n52871,
    n52872, n52873, n52874, n52875, n52876, n52877,
    n52878, n52879, n52880, n52881, n52882, n52883,
    n52884, n52885, n52886, n52887, n52888, n52889,
    n52890, n52891, n52892, n52893, n52894, n52895,
    n52896, n52897, n52898, n52899, n52900, n52901,
    n52902, n52903, n52904, n52905, n52906, n52907,
    n52908, n52909, n52910, n52911, n52912, n52913,
    n52914, n52915, n52916, n52917, n52918, n52919,
    n52920, n52921, n52922, n52923, n52924, n52925,
    n52926, n52927, n52928, n52929, n52930, n52931,
    n52932, n52933, n52934, n52935, n52936, n52937,
    n52938, n52939, n52940, n52941, n52942, n52943,
    n52944, n52945, n52946, n52947, n52948, n52949,
    n52950, n52951, n52952, n52953, n52954, n52955,
    n52956, n52957, n52958, n52959, n52960, n52961,
    n52962, n52963, n52964, n52965, n52966, n52967,
    n52968, n52969, n52970, n52971, n52972, n52973,
    n52974, n52975, n52976, n52977, n52978, n52979,
    n52980, n52981, n52982, n52983, n52984, n52985,
    n52986, n52987, n52988, n52989, n52990, n52991,
    n52992, n52993, n52994, n52995, n52996, n52997,
    n52998, n52999, n53000, n53001, n53002, n53003,
    n53004, n53005, n53006, n53007, n53008, n53009,
    n53010, n53011, n53012, n53013, n53014, n53015,
    n53016, n53017, n53018, n53019, n53020, n53021,
    n53022, n53023, n53024, n53025, n53026, n53027,
    n53028, n53029, n53030, n53031, n53032, n53033,
    n53034, n53035, n53036, n53037, n53038, n53039,
    n53040, n53041, n53042, n53043, n53044, n53045,
    n53046, n53047, n53048, n53049, n53050, n53051,
    n53052, n53053, n53054, n53055, n53056, n53057,
    n53058, n53059, n53060, n53061, n53062, n53063,
    n53064, n53065, n53066, n53067, n53068, n53069,
    n53070, n53071, n53072, n53073, n53074, n53075,
    n53076, n53077, n53078, n53079, n53080, n53081,
    n53082, n53083, n53084, n53085, n53086, n53087,
    n53088, n53089, n53090, n53091, n53092, n53093,
    n53094, n53095, n53096, n53097, n53098, n53099,
    n53100, n53101, n53102, n53103, n53104, n53105,
    n53106, n53107, n53108, n53109, n53110, n53111,
    n53112, n53113, n53114, n53115, n53116, n53117,
    n53118, n53119, n53120, n53121, n53122, n53123,
    n53124, n53125, n53126, n53127, n53128, n53129,
    n53130, n53131, n53132, n53133, n53134, n53135,
    n53136, n53137, n53138, n53139, n53140, n53141,
    n53142, n53143, n53144, n53145, n53146, n53147,
    n53148, n53149, n53150, n53151, n53152, n53153,
    n53154, n53155, n53156, n53157, n53158, n53159,
    n53160, n53161, n53162, n53163, n53164, n53165,
    n53166, n53167, n53168, n53169, n53170, n53171,
    n53172, n53173, n53174, n53175, n53176, n53177,
    n53178, n53179, n53180, n53181, n53182, n53183,
    n53184, n53185, n53186, n53187, n53188, n53189,
    n53190, n53191, n53192, n53193, n53194, n53195,
    n53196, n53197, n53198, n53199, n53200, n53201,
    n53202, n53203, n53204, n53205, n53206, n53207,
    n53208, n53209, n53210, n53211, n53212, n53213,
    n53214, n53215, n53216, n53217, n53218, n53219,
    n53220, n53221, n53222, n53223, n53224, n53225,
    n53226, n53227, n53228, n53229, n53230, n53231,
    n53232, n53233, n53234, n53235, n53236, n53237,
    n53238, n53239, n53240, n53241, n53242, n53243,
    n53244, n53245, n53246, n53247, n53248, n53249,
    n53250, n53251, n53252, n53253, n53254, n53255,
    n53256, n53257, n53258, n53259, n53260, n53261,
    n53262, n53263, n53264, n53265, n53266, n53267,
    n53268, n53269, n53270, n53271, n53272, n53273,
    n53274, n53275, n53276, n53277, n53278, n53279,
    n53280, n53281, n53282, n53283, n53284, n53285,
    n53286, n53287, n53288, n53289, n53290, n53291,
    n53292, n53293, n53294, n53295, n53296, n53297,
    n53298, n53299, n53300, n53301, n53302, n53303,
    n53304, n53305, n53306, n53307, n53308, n53309,
    n53310, n53311, n53312, n53313, n53314, n53315,
    n53316, n53317, n53318, n53319, n53320, n53321,
    n53322, n53323, n53324, n53325, n53326, n53327,
    n53328, n53329, n53330, n53331, n53332, n53333,
    n53334, n53335, n53336, n53337, n53338, n53339,
    n53340, n53341, n53342, n53343, n53344, n53345,
    n53346, n53347, n53348, n53349, n53350, n53351,
    n53352, n53353, n53354, n53355, n53356, n53357,
    n53358, n53359, n53360, n53361, n53362, n53363,
    n53364, n53365, n53366, n53367, n53368, n53369,
    n53370, n53371, n53372, n53373, n53374, n53375,
    n53376, n53377, n53378, n53379, n53380, n53381,
    n53382, n53383, n53384, n53385, n53386, n53387,
    n53388, n53389, n53390, n53391, n53392, n53393,
    n53394, n53395, n53396, n53397, n53398, n53399,
    n53400, n53401, n53402, n53403, n53404, n53405,
    n53406, n53407, n53408, n53409, n53410, n53411,
    n53412, n53413, n53414, n53415, n53416, n53417,
    n53418, n53419, n53420, n53421, n53422, n53423,
    n53424, n53425, n53426, n53427, n53428, n53429,
    n53430, n53431, n53432, n53433, n53434, n53435,
    n53436, n53437, n53438, n53439, n53440, n53441,
    n53442, n53443, n53444, n53445, n53446, n53447,
    n53448, n53449, n53450, n53451, n53452, n53453,
    n53454, n53455, n53456, n53457, n53458, n53459,
    n53460, n53461, n53462, n53463, n53464, n53465,
    n53466, n53467, n53468, n53469, n53470, n53471,
    n53472, n53473, n53474, n53475, n53476, n53477,
    n53478, n53479, n53480, n53481, n53482, n53483,
    n53484, n53485, n53486, n53487, n53488, n53489,
    n53490, n53491, n53492, n53493, n53494, n53495,
    n53496, n53497, n53498, n53499, n53500, n53501,
    n53502, n53503, n53504, n53505, n53506, n53507,
    n53508, n53509, n53510, n53511, n53512, n53513,
    n53514, n53515, n53516, n53517, n53518, n53519,
    n53520, n53521, n53522, n53523, n53524, n53525,
    n53526, n53527, n53528, n53529, n53530, n53531,
    n53532, n53533, n53534, n53535, n53536, n53537,
    n53538, n53539, n53540, n53541, n53542, n53543,
    n53544, n53545, n53546, n53547, n53548, n53549,
    n53550, n53551, n53552, n53553, n53554, n53555,
    n53556, n53557, n53558, n53559, n53560, n53561,
    n53562, n53563, n53564, n53565, n53566, n53567,
    n53568, n53569, n53570, n53571, n53572, n53573,
    n53574, n53575, n53576, n53577, n53578, n53579,
    n53580, n53581, n53582, n53583, n53584, n53585,
    n53586, n53587, n53588, n53589, n53590, n53591,
    n53592, n53593, n53594, n53595, n53596, n53597,
    n53598, n53599, n53600, n53601, n53602, n53603,
    n53604, n53605, n53606, n53607, n53608, n53609,
    n53610, n53611, n53612, n53613, n53614, n53615,
    n53616, n53617, n53618, n53619, n53620, n53621,
    n53622, n53623, n53624, n53625, n53626, n53627,
    n53628, n53629, n53630, n53631, n53632, n53633,
    n53634, n53635, n53636, n53637, n53638, n53639,
    n53640, n53641, n53642, n53643, n53644, n53645,
    n53646, n53647, n53648, n53649, n53650, n53651,
    n53652, n53653, n53654, n53655, n53656, n53657,
    n53658, n53659, n53660, n53661, n53662, n53663,
    n53664, n53665, n53666, n53667, n53668, n53669,
    n53670, n53671, n53672, n53673, n53674, n53675,
    n53676, n53677, n53678, n53679, n53680, n53681,
    n53682, n53683, n53684, n53685, n53686, n53687,
    n53688, n53689, n53690, n53691, n53692, n53693,
    n53694, n53695, n53696, n53697, n53698, n53699,
    n53700, n53701, n53702, n53703, n53704, n53705,
    n53706, n53707, n53708, n53709, n53710, n53711,
    n53712, n53713, n53714, n53715, n53716, n53717,
    n53718, n53719, n53720, n53721, n53722, n53723,
    n53724, n53725, n53726, n53727, n53728, n53729,
    n53730, n53731, n53732, n53733, n53734, n53735,
    n53736, n53737, n53738, n53739, n53740, n53741,
    n53742, n53743, n53744, n53745, n53746, n53747,
    n53748, n53749, n53750, n53751, n53752, n53753,
    n53754, n53755, n53756, n53757, n53758, n53759,
    n53760, n53761, n53762, n53763, n53764, n53765,
    n53766, n53767, n53768, n53769, n53770, n53771,
    n53772, n53773, n53774, n53775, n53776, n53777,
    n53778, n53779, n53780, n53781, n53782, n53783,
    n53784, n53785, n53786, n53787, n53788, n53789,
    n53790, n53791, n53792, n53793, n53794, n53795,
    n53796, n53797, n53798, n53799, n53800, n53801,
    n53802, n53803, n53804, n53805, n53806, n53807,
    n53808, n53809, n53810, n53811, n53812, n53813,
    n53814, n53815, n53816, n53817, n53818, n53819,
    n53820, n53821, n53822, n53823, n53824, n53825,
    n53826, n53827, n53828, n53829, n53830, n53831,
    n53832, n53833, n53834, n53835, n53836, n53837,
    n53838, n53839, n53840, n53841, n53842, n53843,
    n53844, n53845, n53846, n53847, n53848, n53849,
    n53850, n53851, n53852, n53853, n53854, n53855,
    n53856, n53857, n53858, n53859, n53860, n53861,
    n53862, n53863, n53864, n53865, n53866, n53867,
    n53868, n53869, n53870, n53871, n53872, n53873,
    n53874, n53875, n53876, n53877, n53878, n53879,
    n53880, n53881, n53882, n53883, n53884, n53885,
    n53886, n53887, n53888, n53889, n53890, n53891,
    n53892, n53893, n53894, n53895, n53896, n53897,
    n53898, n53899, n53900, n53901, n53902, n53903,
    n53904, n53905, n53906, n53907, n53908, n53909,
    n53910, n53911, n53912, n53913, n53914, n53915,
    n53916, n53917, n53918, n53919, n53920, n53921,
    n53922, n53923, n53924, n53925, n53926, n53927,
    n53928, n53929, n53930, n53931, n53932, n53933,
    n53934, n53935, n53936, n53937, n53938, n53939,
    n53940, n53941, n53942, n53943, n53944, n53945,
    n53946, n53947, n53948, n53949, n53950, n53951,
    n53952, n53953, n53954, n53955, n53956, n53957,
    n53958, n53959, n53960, n53961, n53962, n53963,
    n53964, n53965, n53966, n53967, n53968, n53969,
    n53970, n53971, n53972, n53973, n53974, n53975,
    n53976, n53977, n53978, n53980, n53981, n53982,
    n53983, n53984, n53985, n53986, n53987, n53988,
    n53989, n53990, n53991, n53992, n53993, n53994,
    n53995, n53996, n53997, n53998, n53999, n54000,
    n54001, n54002, n54003, n54004, n54005, n54006,
    n54007, n54008, n54009, n54010, n54011, n54012,
    n54013, n54014, n54015, n54016, n54017, n54018,
    n54019, n54020, n54021, n54022, n54023, n54024,
    n54025, n54026, n54027, n54028, n54029, n54030,
    n54031, n54032, n54033, n54034, n54035, n54036,
    n54037, n54038, n54039, n54040, n54041, n54042,
    n54043, n54044, n54045, n54046, n54047, n54048,
    n54049, n54050, n54051, n54052, n54053, n54054,
    n54055, n54056, n54057, n54058, n54059, n54060,
    n54061, n54062, n54063, n54064, n54065, n54066,
    n54067, n54068, n54069, n54070, n54071, n54072,
    n54073, n54074, n54075, n54076, n54077, n54078,
    n54079, n54080, n54081, n54082, n54083, n54084,
    n54085, n54086, n54087, n54088, n54089, n54090,
    n54091, n54092, n54093, n54094, n54095, n54096,
    n54097, n54098, n54099, n54100, n54101, n54102,
    n54103, n54104, n54105, n54106, n54107, n54108,
    n54109, n54110, n54111, n54112, n54113, n54114,
    n54115, n54116, n54117, n54118, n54119, n54120,
    n54121, n54122, n54123, n54124, n54125, n54126,
    n54127, n54128, n54129, n54130, n54131, n54132,
    n54133, n54134, n54135, n54136, n54137, n54138,
    n54139, n54140, n54141, n54142, n54143, n54144,
    n54145, n54146, n54147, n54148, n54149, n54150,
    n54151, n54152, n54153, n54154, n54155, n54156,
    n54157, n54158, n54160, n54161, n54162, n54163,
    n54164, n54165, n54166, n54167, n54168, n54169,
    n54170, n54171, n54172, n54173, n54174, n54175,
    n54176, n54177, n54178, n54179, n54180, n54181,
    n54182, n54183, n54184, n54185, n54186, n54187,
    n54188, n54189, n54190, n54191, n54192, n54193,
    n54194, n54195, n54196, n54197, n54198, n54199,
    n54200, n54201, n54202, n54203, n54204, n54205,
    n54206, n54207, n54208, n54209, n54211, n54212,
    n54213, n54214, n54215, n54216, n54217, n54218,
    n54219, n54220, n54221, n54222, n54223, n54224,
    n54225, n54226, n54227, n54228, n54229, n54230,
    n54231, n54232, n54233, n54234, n54235, n54236,
    n54237, n54238, n54239, n54240, n54241, n54242,
    n54243, n54244, n54245, n54246, n54247, n54248,
    n54249, n54250, n54251, n54252, n54253, n54254,
    n54255, n54256, n54257, n54258, n54259, n54260,
    n54261, n54262, n54263, n54264, n54265, n54266,
    n54267, n54268, n54269, n54270, n54271, n54272,
    n54273, n54274, n54275, n54276, n54277, n54278,
    n54279, n54280, n54281, n54282, n54283, n54284,
    n54285, n54286, n54287, n54288, n54289, n54290,
    n54291, n54292, n54293, n54294, n54295, n54296,
    n54297, n54298, n54299, n54300, n54301, n54302,
    n54303, n54304, n54305, n54306, n54307, n54308,
    n54309, n54310, n54311, n54312, n54313, n54314,
    n54315, n54316, n54317, n54318, n54320, n54321,
    n54322, n54323, n54324, n54325, n54326, n54327,
    n54328, n54329, n54330, n54331, n54332, n54333,
    n54334, n54335, n54336, n54337, n54338, n54339,
    n54340, n54341, n54342, n54343, n54344, n54345,
    n54346, n54347, n54348, n54349, n54350, n54351,
    n54352, n54353, n54354, n54355, n54356, n54357,
    n54358, n54359, n54360, n54361, n54362, n54363,
    n54364, n54365, n54366, n54367, n54368, n54369,
    n54370, n54371, n54372, n54373, n54374, n54375,
    n54376, n54377, n54378, n54379, n54380, n54381,
    n54382, n54383, n54384, n54385, n54386, n54387,
    n54388, n54389, n54390, n54391, n54392, n54393,
    n54394, n54395, n54396, n54397, n54398, n54399,
    n54400, n54401, n54402, n54403, n54404, n54405,
    n54406, n54407, n54408, n54409, n54410, n54411,
    n54412, n54413, n54414, n54415, n54416, n54417,
    n54418, n54419, n54420, n54421, n54422, n54423,
    n54424, n54425, n54426, n54427, n54428, n54429,
    n54430, n54431, n54432, n54433, n54434, n54435,
    n54436, n54437, n54438, n54439, n54440, n54441,
    n54442, n54443, n54444, n54445, n54446, n54447,
    n54448, n54449, n54450, n54451, n54452, n54453,
    n54454, n54455, n54456, n54457, n54458, n54459,
    n54460, n54461, n54462, n54463, n54464, n54465,
    n54466, n54467, n54468, n54469, n54470, n54471,
    n54472, n54473, n54474, n54475, n54476, n54477,
    n54478, n54479, n54480, n54481, n54482, n54484,
    n54485, n54486, n54487, n54488, n54489, n54490,
    n54491, n54492, n54493, n54494, n54495, n54496,
    n54497, n54498, n54499, n54500, n54501, n54502,
    n54503, n54504, n54505, n54506, n54507, n54508,
    n54509, n54510, n54511, n54512, n54513, n54514,
    n54515, n54516, n54517, n54518, n54519, n54520,
    n54521, n54522, n54523, n54524, n54525, n54526,
    n54527, n54528, n54529, n54530, n54531, n54532,
    n54533, n54534, n54535, n54536, n54537, n54538,
    n54539, n54540, n54541, n54542, n54543, n54544,
    n54545, n54547, n54548, n54549, n54550, n54551,
    n54552, n54553, n54554, n54555, n54556, n54557,
    n54558, n54559, n54560, n54561, n54562, n54563,
    n54564, n54565, n54566, n54567, n54568, n54569,
    n54570, n54571, n54572, n54573, n54574, n54575,
    n54576, n54577, n54578, n54579, n54580, n54581,
    n54582, n54583, n54584, n54585, n54586, n54587,
    n54588, n54589, n54590, n54591, n54592, n54593,
    n54594, n54595, n54596, n54597, n54598, n54599,
    n54600, n54601, n54602, n54603, n54604, n54605,
    n54606, n54607, n54608, n54609, n54610, n54611,
    n54612, n54613, n54614, n54615, n54616, n54617,
    n54618, n54619, n54620, n54621, n54622, n54623,
    n54624, n54625, n54626, n54627, n54628, n54629,
    n54630, n54631, n54632, n54633, n54634, n54635,
    n54636, n54637, n54638, n54639, n54640, n54641,
    n54642, n54643, n54644, n54645, n54646, n54647,
    n54648, n54649, n54650, n54651, n54653, n54654,
    n54655, n54656, n54657, n54658, n54659, n54660,
    n54661, n54662, n54663, n54664, n54665, n54666,
    n54667, n54668, n54669, n54670, n54671, n54672,
    n54673, n54674, n54675, n54676, n54677, n54678,
    n54679, n54680, n54681, n54682, n54683, n54684,
    n54685, n54686, n54687, n54688, n54689, n54690,
    n54691, n54692, n54693, n54694, n54696, n54697,
    n54698, n54699, n54700, n54701, n54702, n54703,
    n54704, n54705, n54706, n54707, n54708, n54709,
    n54710, n54711, n54712, n54713, n54714, n54715,
    n54716, n54717, n54718, n54719, n54720, n54721,
    n54722, n54723, n54724, n54725, n54726, n54727,
    n54728, n54729, n54730, n54731, n54732, n54733,
    n54734, n54735, n54736, n54737, n54738, n54739,
    n54740, n54741, n54742, n54743, n54744, n54745,
    n54746, n54747, n54748, n54749, n54750, n54751,
    n54752, n54753, n54754, n54755, n54756, n54757,
    n54758, n54759, n54760, n54761, n54762, n54763,
    n54764, n54765, n54766, n54767, n54768, n54769,
    n54770, n54771, n54772, n54773, n54774, n54775,
    n54776, n54777, n54778, n54779, n54780, n54781,
    n54782, n54783, n54784, n54785, n54786, n54787,
    n54788, n54789, n54790, n54791, n54792, n54793,
    n54794, n54795, n54796, n54797, n54798, n54799,
    n54800, n54801, n54802, n54803, n54804, n54805,
    n54806, n54807, n54808, n54809, n54810, n54811,
    n54812, n54813, n54814, n54815, n54816, n54817,
    n54818, n54819, n54820, n54821, n54822, n54823,
    n54824, n54825, n54826, n54827, n54828, n54829,
    n54830, n54831, n54832, n54833, n54834, n54835,
    n54836, n54837, n54838, n54839, n54840, n54841,
    n54842, n54843, n54844, n54845, n54846, n54847,
    n54848, n54849, n54850, n54851, n54852, n54853,
    n54854, n54855, n54856, n54857, n54858, n54859,
    n54860, n54861, n54862, n54863, n54864, n54865,
    n54866, n54867, n54868, n54869, n54870, n54871,
    n54872, n54873, n54874, n54875, n54876, n54877,
    n54878, n54879, n54880, n54881, n54882, n54883,
    n54884, n54885, n54886, n54887, n54888, n54889,
    n54890, n54891, n54892, n54893, n54894, n54895,
    n54896, n54897, n54898, n54899, n54900, n54901,
    n54902, n54903, n54904, n54905, n54906, n54907,
    n54908, n54909, n54910, n54911, n54912, n54913,
    n54914, n54915, n54916, n54917, n54918, n54919,
    n54920, n54921, n54922, n54923, n54924, n54925,
    n54926, n54927, n54928, n54929, n54930, n54931,
    n54932, n54933, n54934, n54935, n54936, n54937,
    n54938, n54939, n54940, n54941, n54942, n54943,
    n54944, n54945, n54946, n54947, n54948, n54949,
    n54950, n54951, n54952, n54953, n54954, n54955,
    n54956, n54957, n54958, n54959, n54960, n54961,
    n54962, n54963, n54964, n54965, n54966, n54967,
    n54968, n54969, n54971, n54972, n54973, n54974,
    n54975, n54976, n54977, n54978, n54979, n54980,
    n54981, n54982, n54983, n54984, n54985, n54986,
    n54987, n54988, n54989, n54990, n54991, n54992,
    n54993, n54994, n54995, n54996, n54997, n54998,
    n54999, n55000, n55001, n55002, n55003, n55004,
    n55005, n55006, n55007, n55008, n55009, n55010,
    n55011, n55012, n55014, n55015, n55016, n55017,
    n55018, n55019, n55020, n55021, n55022, n55023,
    n55024, n55025, n55026, n55027, n55028, n55029,
    n55030, n55031, n55032, n55033, n55034, n55035,
    n55036, n55037, n55038, n55039, n55040, n55041,
    n55042, n55043, n55044, n55045, n55046, n55047,
    n55048, n55049, n55050, n55051, n55052, n55053,
    n55054, n55055, n55056, n55057, n55058, n55059,
    n55060, n55061, n55062, n55063, n55064, n55065,
    n55066, n55068, n55069, n55071, n55072, n55073,
    n55074, n55075, n55076, n55077, n55078, n55079,
    n55080, n55081, n55082, n55083, n55084, n55085,
    n55086, n55087, n55088, n55089, n55090, n55091,
    n55092, n55093, n55095, n55096, n55097, n55098,
    n55099, n55100, n55101, n55102, n55103, n55104,
    n55105, n55106, n55107, n55108, n55109, n55110,
    n55111, n55113, n55114, n55115, n55116, n55117,
    n55118, n55119, n55120, n55122, n55123, n55124,
    n55125, n55126, n55127, n55128, n55129, n55130,
    n55131, n55132, n55133, n55134, n55135, n55136,
    n55137, n55138, n55139, n55140, n55141, n55142,
    n55143, n55144, n55145, n55146, n55147, n55148,
    n55149, n55150, n55151, n55152, n55153, n55154,
    n55155, n55156, n55157, n55158, n55159, n55160,
    n55161, n55162, n55163, n55164, n55165, n55166,
    n55167, n55168, n55169, n55170, n55171, n55172,
    n55173, n55174, n55175, n55176, n55177, n55178,
    n55179, n55180, n55181, n55182, n55183, n55184,
    n55185, n55186, n55187, n55188, n55189, n55190,
    n55191, n55192, n55193, n55194, n55195, n55196,
    n55197, n55198, n55199, n55200, n55202, n55203,
    n55204, n55205, n55206, n55207, n55208, n55209,
    n55210, n55211, n55212, n55213, n55214, n55215,
    n55216, n55217, n55218, n55219, n55220, n55222,
    n55223, n55224, n55225, n55226, n55227, n55228,
    n55229, n55230, n55231, n55232, n55233, n55234,
    n55235, n55236, n55237, n55238, n55239, n55240,
    n55241, n55242, n55243, n55244, n55245, n55246,
    n55247, n55248, n55249, n55250, n55251, n55252,
    n55253, n55254, n55255, n55256, n55257, n55258,
    n55259, n55260, n55261, n55262, n55263, n55264,
    n55265, n55266, n55267, n55268, n55269, n55270,
    n55271, n55272, n55273, n55274, n55275, n55276,
    n55277, n55278, n55279, n55280, n55281, n55282,
    n55283, n55284, n55285, n55286, n55287, n55288,
    n55289, n55290, n55291, n55292, n55293, n55294,
    n55295, n55296, n55297, n55298, n55299, n55300,
    n55301, n55302, n55303, n55304, n55305, n55306,
    n55307, n55308, n55309, n55310, n55312, n55314,
    n55316, n55317, n55318, n55320, n55322, n55324,
    n55326, n55328, n55330, n55332, n55333, n55334,
    n55335, n55336, n55337, n55338, n55339, n55340,
    n55341, n55342, n55343, n55344, n55345, n55346,
    n55347, n55348, n55349, n55350, n55351, n55352,
    n55353, n55354, n55355, n55356, n55357, n55358,
    n55360, n55361, n55362, n55363, n55364, n55365,
    n55366, n55367, n55368, n55369, n55370, n55371,
    n55372, n55373, n55374, n55375, n55376, n55377,
    n55378, n55379, n55380, n55381, n55382, n55383,
    n55384, n55385, n55386, n55387, n55388, n55389,
    n55390, n55391, n55392, n55393, n55394, n55395,
    n55396, n55397, n55398, n55399, n55400, n55401,
    n55402, n55403, n55404, n55405, n55406, n55407,
    n55408, n55409, n55410, n55411, n55412, n55413,
    n55414, n55415, n55416, n55417, n55418, n55419,
    n55420, n55421, n55422, n55423, n55424, n55425,
    n55426, n55427, n55428, n55429, n55430, n55431,
    n55432, n55433, n55434, n55435, n55436, n55437,
    n55438, n55439, n55440, n55441, n55442, n55443,
    n55444, n55445, n55446, n55447, n55449, n55450,
    n55451, n55452, n55453, n55454, n55455, n55456,
    n55457, n55458, n55459, n55460, n55461, n55462,
    n55463, n55464, n55465, n55466, n55467, n55468,
    n55469, n55470, n55471, n55472, n55473, n55474,
    n55475, n55476, n55477, n55478, n55479, n55480,
    n55481, n55482, n55483, n55484, n55485, n55486,
    n55487, n55488, n55489, n55490, n55491, n55492,
    n55493, n55494, n55495, n55496, n55497, n55498,
    n55499, n55500, n55501, n55502, n55503, n55504,
    n55505, n55506, n55507, n55508, n55509, n55510,
    n55511, n55512, n55513, n55514, n55515, n55516,
    n55517, n55518, n55519, n55520, n55521, n55522,
    n55523, n55524, n55525, n55526, n55527, n55528,
    n55529, n55530, n55531, n55532, n55533, n55534,
    n55535, n55536, n55537, n55538, n55539, n55540,
    n55541, n55542, n55543, n55544, n55545, n55546,
    n55547, n55548, n55549, n55550, n55551, n55552,
    n55553, n55554, n55555, n55556, n55557, n55558,
    n55559, n55560, n55561, n55562, n55563, n55564,
    n55565, n55566, n55567, n55568, n55569, n55570,
    n55571, n55572, n55573, n55574, n55575, n55576,
    n55577, n55578, n55579, n55580, n55581, n55582,
    n55583, n55584, n55586, n55587, n55588, n55589,
    n55590, n55591, n55592, n55593, n55594, n55595,
    n55596, n55597, n55599, n55600, n55601, n55602,
    n55603, n55604, n55605, n55606, n55607, n55608,
    n55609, n55610, n55612, n55613, n55614, n55615,
    n55616, n55617, n55618, n55619, n55620, n55621,
    n55622, n55623, n55624, n55625, n55626, n55627,
    n55628, n55629, n55630, n55631, n55632, n55633,
    n55634, n55635, n55636, n55637, n55638, n55639,
    n55640, n55641, n55642, n55643, n55644, n55645,
    n55646, n55647, n55648, n55649, n55650, n55651,
    n55652, n55653, n55654, n55655, n55656, n55657,
    n55658, n55659, n55660, n55661, n55662, n55663,
    n55664, n55665, n55666, n55667, n55668, n55669,
    n55670, n55671, n55672, n55673, n55674, n55675,
    n55676, n55677, n55678, n55679, n55680, n55681,
    n55682, n55683, n55684, n55685, n55686, n55687,
    n55688, n55689, n55690, n55691, n55692, n55693,
    n55694, n55695, n55696, n55697, n55698, n55699,
    n55700, n55701, n55702, n55703, n55704, n55705,
    n55706, n55707, n55708, n55709, n55710, n55711,
    n55712, n55713, n55714, n55715, n55716, n55717,
    n55718, n55719, n55720, n55721, n55722, n55723,
    n55724, n55725, n55726, n55727, n55728, n55729,
    n55730, n55731, n55732, n55733, n55734, n55735,
    n55736, n55737, n55738, n55739, n55740, n55741,
    n55742, n55743, n55744, n55745, n55746, n55747,
    n55748, n55749, n55750, n55751, n55752, n55753,
    n55754, n55755, n55756, n55757, n55758, n55759,
    n55760, n55761, n55762, n55763, n55764, n55765,
    n55766, n55767, n55768, n55769, n55770, n55771,
    n55772, n55773, n55774, n55775, n55776, n55777,
    n55778, n55779, n55780, n55781, n55782, n55783,
    n55784, n55785, n55786, n55787, n55788, n55789,
    n55790, n55791, n55792, n55793, n55794, n55795,
    n55796, n55797, n55798, n55799, n55800, n55801,
    n55802, n55803, n55804, n55805, n55806, n55807,
    n55808, n55809, n55810, n55811, n55812, n55813,
    n55814, n55815, n55816, n55817, n55818, n55819,
    n55820, n55821, n55822, n55823, n55824, n55825,
    n55826, n55827, n55828, n55829, n55830, n55831,
    n55832, n55833, n55834, n55835, n55836, n55837,
    n55838, n55839, n55840, n55841, n55842, n55843,
    n55844, n55845, n55846, n55847, n55848, n55849,
    n55850, n55851, n55852, n55853, n55854, n55855,
    n55856, n55857, n55858, n55859, n55860, n55861,
    n55862, n55863, n55864, n55865, n55866, n55867,
    n55868, n55869, n55870, n55871, n55872, n55873,
    n55874, n55875, n55876, n55877, n55878, n55879,
    n55880, n55881, n55882, n55883, n55884, n55885,
    n55886, n55887, n55888, n55889, n55890, n55891,
    n55892, n55893, n55894, n55895, n55896, n55897,
    n55898, n55899, n55900, n55901, n55902, n55903,
    n55904, n55905, n55906, n55907, n55908, n55909,
    n55910, n55911, n55912, n55913, n55914, n55915,
    n55916, n55917, n55918, n55919, n55920, n55921,
    n55922, n55923, n55924, n55925, n55926, n55927,
    n55928, n55929, n55930, n55931, n55932, n55933,
    n55934, n55935, n55936, n55937, n55938, n55939,
    n55940, n55941, n55942, n55943, n55944, n55945,
    n55946, n55947, n55948, n55949, n55950, n55951,
    n55952, n55953, n55954, n55955, n55956, n55957,
    n55958, n55959, n55960, n55961, n55962, n55963,
    n55964, n55965, n55966, n55967, n55968, n55969,
    n55970, n55971, n55972, n55973, n55974, n55975,
    n55976, n55977, n55978, n55979, n55980, n55981,
    n55982, n55983, n55984, n55985, n55986, n55987,
    n55988, n55989, n55990, n55991, n55992, n55993,
    n55994, n55995, n55996, n55997, n55998, n55999,
    n56000, n56001, n56002, n56003, n56004, n56005,
    n56006, n56007, n56008, n56009, n56010, n56011,
    n56012, n56013, n56014, n56015, n56016, n56017,
    n56018, n56019, n56020, n56021, n56022, n56023,
    n56024, n56025, n56026, n56027, n56028, n56029,
    n56030, n56031, n56032, n56033, n56034, n56035,
    n56036, n56037, n56038, n56039, n56040, n56041,
    n56042, n56043, n56044, n56045, n56046, n56047,
    n56048, n56049, n56050, n56051, n56052, n56053,
    n56054, n56055, n56056, n56057, n56058, n56059,
    n56060, n56061, n56062, n56063, n56064, n56065,
    n56066, n56067, n56068, n56069, n56070, n56071,
    n56072, n56073, n56074, n56075, n56076, n56077,
    n56078, n56079, n56080, n56081, n56082, n56083,
    n56084, n56085, n56086, n56087, n56088, n56089,
    n56090, n56091, n56092, n56093, n56094, n56095,
    n56096, n56097, n56098, n56099, n56100, n56101,
    n56102, n56103, n56104, n56105, n56106, n56107,
    n56108, n56109, n56110, n56111, n56112, n56113,
    n56114, n56115, n56116, n56117, n56118, n56119,
    n56120, n56121, n56122, n56123, n56124, n56125,
    n56126, n56127, n56128, n56129, n56130, n56131,
    n56132, n56133, n56134, n56135, n56136, n56137,
    n56138, n56139, n56140, n56141, n56142, n56143,
    n56144, n56145, n56146, n56147, n56148, n56149,
    n56150, n56151, n56152, n56153, n56154, n56155,
    n56156, n56157, n56158, n56159, n56160, n56161,
    n56162, n56163, n56164, n56165, n56166, n56167,
    n56168, n56169, n56170, n56171, n56172, n56173,
    n56174, n56175, n56176, n56177, n56178, n56179,
    n56180, n56181, n56182, n56183, n56184, n56185,
    n56186, n56187, n56188, n56189, n56190, n56191,
    n56192, n56193, n56194, n56195, n56196, n56197,
    n56198, n56199, n56200, n56201, n56202, n56203,
    n56204, n56205, n56206, n56207, n56208, n56209,
    n56210, n56211, n56212, n56213, n56214, n56215,
    n56216, n56217, n56218, n56219, n56220, n56221,
    n56222, n56223, n56224, n56225, n56226, n56227,
    n56228, n56229, n56230, n56231, n56232, n56233,
    n56234, n56235, n56236, n56237, n56238, n56239,
    n56240, n56241, n56242, n56243, n56244, n56245,
    n56246, n56247, n56248, n56249, n56250, n56251,
    n56252, n56253, n56254, n56255, n56256, n56257,
    n56258, n56259, n56260, n56261, n56262, n56263,
    n56264, n56265, n56266, n56267, n56268, n56269,
    n56270, n56271, n56272, n56273, n56274, n56275,
    n56276, n56277, n56278, n56279, n56280, n56281,
    n56282, n56283, n56284, n56285, n56286, n56287,
    n56288, n56289, n56290, n56291, n56292, n56293,
    n56294, n56295, n56296, n56297, n56298, n56299,
    n56300, n56301, n56302, n56303, n56304, n56305,
    n56306, n56307, n56308, n56309, n56310, n56311,
    n56312, n56313, n56314, n56315, n56316, n56317,
    n56318, n56319, n56320, n56321, n56322, n56323,
    n56324, n56325, n56326, n56327, n56328, n56329,
    n56330, n56331, n56332, n56333, n56334, n56335,
    n56336, n56337, n56338, n56339, n56340, n56341,
    n56342, n56343, n56344, n56345, n56346, n56347,
    n56348, n56349, n56350, n56351, n56352, n56353,
    n56354, n56355, n56356, n56357, n56358, n56359,
    n56360, n56361, n56362, n56363, n56364, n56365,
    n56366, n56367, n56368, n56369, n56370, n56371,
    n56372, n56373, n56374, n56375, n56376, n56377,
    n56378, n56379, n56380, n56381, n56382, n56383,
    n56384, n56385, n56386, n56387, n56388, n56389,
    n56390, n56391, n56392, n56393, n56394, n56395,
    n56396, n56397, n56398, n56399, n56400, n56401,
    n56402, n56403, n56404, n56405, n56406, n56407,
    n56408, n56409, n56410, n56411, n56412, n56413,
    n56414, n56415, n56416, n56417, n56418, n56419,
    n56420, n56421, n56422, n56423, n56424, n56425,
    n56426, n56427, n56428, n56429, n56430, n56431,
    n56432, n56433, n56434, n56435, n56436, n56437,
    n56438, n56439, n56440, n56441, n56442, n56443,
    n56444, n56445, n56446, n56447, n56448, n56449,
    n56450, n56451, n56452, n56453, n56454, n56455,
    n56456, n56457, n56458, n56459, n56460, n56461,
    n56462, n56463, n56464, n56465, n56466, n56467,
    n56468, n56469, n56470, n56471, n56472, n56473,
    n56474, n56475, n56476, n56477, n56478, n56479,
    n56480, n56481, n56482, n56483, n56484, n56485,
    n56486, n56487, n56488, n56489, n56490, n56491,
    n56492, n56493, n56494, n56495, n56496, n56497,
    n56498, n56499, n56500, n56501, n56502, n56503,
    n56504, n56505, n56506, n56507, n56508, n56509,
    n56510, n56511, n56512, n56513, n56514, n56515,
    n56516, n56517, n56518, n56519, n56520, n56521,
    n56522, n56523, n56524, n56525, n56526, n56527,
    n56528, n56529, n56530, n56531, n56532, n56533,
    n56534, n56535, n56536, n56537, n56538, n56539,
    n56540, n56541, n56542, n56543, n56544, n56545,
    n56546, n56547, n56548, n56549, n56550, n56551,
    n56552, n56553, n56554, n56555, n56556, n56557,
    n56558, n56559, n56560, n56561, n56562, n56563,
    n56564, n56565, n56566, n56567, n56568, n56569,
    n56570, n56571, n56572, n56573, n56574, n56575,
    n56576, n56577, n56578, n56579, n56580, n56581,
    n56582, n56583, n56584, n56585, n56586, n56587,
    n56588, n56589, n56590, n56591, n56592, n56593,
    n56594, n56595, n56596, n56597, n56598, n56599,
    n56600, n56601, n56602, n56603, n56604, n56605,
    n56606, n56607, n56608, n56609, n56610, n56611,
    n56612, n56613, n56614, n56615, n56616, n56617,
    n56618, n56619, n56620, n56621, n56622, n56623,
    n56624, n56625, n56626, n56627, n56628, n56629,
    n56630, n56631, n56632, n56633, n56634, n56635,
    n56636, n56637, n56638, n56639, n56640, n56641,
    n56642, n56643, n56644, n56645, n56646, n56647,
    n56648, n56649, n56650, n56651, n56652, n56653,
    n56655, n56656, n56658, n56659, n56660, n56661,
    n56662, n56663, n56664, n56665, n56666, n56667,
    n56668, n56669, n56670, n56671, n56672, n56673,
    n56674, n56675, n56676, n56677, n56678, n56679,
    n56680, n56681, n56682, n56683, n56684, n56685,
    n56686, n56687, n56688, n56689, n56690, n56691,
    n56692, n56693, n56694, n56695, n56696, n56697,
    n56698, n56699, n56700, n56701, n56702, n56703,
    n56704, n56705, n56706, n56707, n56708, n56709,
    n56711, n56712, n56713, n56714, n56715, n56716,
    n56717, n56718, n56719, n56720, n56721, n56722,
    n56723, n56724, n56725, n56726, n56727, n56728,
    n56729, n56730, n56731, n56732, n56733, n56734,
    n56735, n56736, n56737, n56738, n56739, n56740,
    n56741, n56742, n56743, n56744, n56745, n56746,
    n56747, n56748, n56749, n56750, n56751, n56752,
    n56753, n56754, n56755, n56756, n56757, n56758,
    n56759, n56760, n56761, n56762, n56763, n56764,
    n56765, n56766, n56767, n56768, n56770, n56771,
    n56772, n56773, n56774, n56775, n56776, n56777,
    n56778, n56779, n56780, n56781, n56782, n56783,
    n56784, n56785, n56786, n56787, n56788, n56789,
    n56790, n56791, n56792, n56793, n56794, n56795,
    n56796, n56797, n56798, n56799, n56800, n56801,
    n56802, n56803, n56804, n56805, n56806, n56807,
    n56808, n56809, n56810, n56811, n56812, n56813,
    n56814, n56815, n56816, n56817, n56818, n56819,
    n56820, n56821, n56822, n56823, n56824, n56825,
    n56826, n56827, n56828, n56829, n56830, n56831,
    n56832, n56833, n56834, n56835, n56836, n56837,
    n56839, n56840, n56841, n56842, n56843, n56844,
    n56845, n56846, n56847, n56848, n56849, n56850,
    n56851, n56852, n56853, n56854, n56855, n56856,
    n56857, n56858, n56859, n56860, n56861, n56862,
    n56863, n56864, n56865, n56866, n56867, n56868,
    n56869, n56870, n56871, n56872, n56873, n56874,
    n56875, n56876, n56877, n56878, n56879, n56880,
    n56881, n56882, n56883, n56884, n56885, n56886,
    n56887, n56888, n56889, n56890, n56891, n56892,
    n56893, n56894, n56895, n56896, n56897, n56898,
    n56899, n56900, n56901, n56902, n56903, n56904,
    n56905, n56906, n56907, n56908, n56909, n56910,
    n56911, n56912, n56913, n56914, n56915, n56916,
    n56917, n56918, n56919, n56920, n56921, n56922,
    n56923, n56924, n56925, n56926, n56927, n56928,
    n56929, n56930, n56931, n56932, n56933, n56934,
    n56935, n56936, n56937, n56938, n56939, n56940,
    n56941, n56942, n56943, n56944, n56945, n56946,
    n56947, n56948, n56949, n56950, n56951, n56952,
    n56953, n56954, n56955, n56956, n56957, n56958,
    n56959, n56960, n56961, n56962, n56963, n56964,
    n56965, n56966, n56967, n56968, n56969, n56970,
    n56971, n56972, n56973, n56974, n56975, n56976,
    n56977, n56978, n56979, n56980, n56981, n56982,
    n56983, n56984, n56985, n56986, n56987, n56988,
    n56989, n56990, n56991, n56992, n56993, n56994,
    n56995, n56996, n56997, n56998, n56999, n57000,
    n57001, n57002, n57003, n57004, n57005, n57006,
    n57007, n57008, n57009, n57010, n57011, n57012,
    n57013, n57014, n57015, n57016, n57017, n57018,
    n57019, n57020, n57021, n57022, n57023, n57024,
    n57025, n57026, n57027, n57028, n57029, n57030,
    n57031, n57032, n57033, n57034, n57035, n57036,
    n57037, n57038, n57039, n57040, n57041, n57042,
    n57043, n57044, n57045, n57046, n57047, n57048,
    n57049, n57050, n57051, n57052, n57053, n57054,
    n57055, n57056, n57057, n57058, n57059, n57060,
    n57061, n57062, n57063, n57064, n57065, n57066,
    n57067, n57068, n57069, n57070, n57071, n57072,
    n57073, n57074, n57075, n57076, n57077, n57078,
    n57079, n57080, n57082, n57083, n57084, n57085,
    n57086, n57087, n57088, n57089, n57090, n57091,
    n57092, n57093, n57094, n57095, n57096, n57097,
    n57098, n57099, n57100, n57101, n57102, n57103,
    n57104, n57105, n57106, n57107, n57108, n57109,
    n57110, n57111, n57112, n57113, n57114, n57115,
    n57116, n57117, n57118, n57119, n57120, n57121,
    n57122, n57123, n57124, n57125, n57126, n57127,
    n57128, n57129, n57130, n57131, n57132, n57133,
    n57134, n57135, n57136, n57137, n57138, n57139,
    n57140, n57141, n57142, n57143, n57144, n57145,
    n57146, n57147, n57148, n57149, n57150, n57151,
    n57152, n57153, n57154, n57155, n57156, n57157,
    n57158, n57159, n57160, n57161, n57162, n57163,
    n57164, n57165, n57166, n57167, n57168, n57169,
    n57170, n57171, n57172, n57173, n57174, n57175,
    n57176, n57177, n57178, n57179, n57180, n57181,
    n57182, n57183, n57184, n57185, n57186, n57187,
    n57188, n57189, n57190, n57191, n57192, n57193,
    n57194, n57195, n57196, n57197, n57198, n57199,
    n57200, n57201, n57202, n57203, n57204, n57205,
    n57206, n57207, n57208, n57209, n57210, n57211,
    n57212, n57213, n57214, n57215, n57216, n57217,
    n57218, n57219, n57220, n57221, n57222, n57223,
    n57224, n57225, n57226, n57227, n57228, n57229,
    n57230, n57231, n57232, n57233, n57234, n57235,
    n57236, n57237, n57238, n57239, n57240, n57241,
    n57242, n57243, n57244, n57245, n57246, n57247,
    n57248, n57249, n57250, n57251, n57252, n57253,
    n57254, n57255, n57256, n57257, n57258, n57259,
    n57260, n57261, n57262, n57263, n57264, n57265,
    n57266, n57267, n57268, n57269, n57270, n57271,
    n57272, n57273, n57274, n57275, n57276, n57277,
    n57278, n57279, n57280, n57281, n57282, n57283,
    n57284, n57285, n57286, n57287, n57288, n57289,
    n57290, n57291, n57292, n57293, n57294, n57295,
    n57296, n57297, n57298, n57299, n57300, n57301,
    n57302, n57303, n57304, n57305, n57306, n57307,
    n57308, n57309, n57310, n57311, n57312, n57313,
    n57314, n57315, n57316, n57317, n57318, n57319,
    n57320, n57321, n57322, n57323, n57324, n57325,
    n57326, n57327, n57328, n57329, n57330, n57331,
    n57332, n57333, n57334, n57335, n57336, n57337,
    n57338, n57339, n57340, n57341, n57342, n57343,
    n57344, n57345, n57346, n57347, n57348, n57349,
    n57350, n57351, n57352, n57353, n57354, n57355,
    n57356, n57357, n57358, n57359, n57360, n57361,
    n57362, n57363, n57364, n57365, n57366, n57367,
    n57368, n57369, n57370, n57371, n57372, n57373,
    n57374, n57375, n57376, n57377, n57378, n57379,
    n57380, n57381, n57382, n57383, n57384, n57385,
    n57386, n57387, n57388, n57389, n57390, n57391,
    n57392, n57393, n57394, n57395, n57396, n57397,
    n57398, n57399, n57400, n57401, n57402, n57403,
    n57404, n57405, n57406, n57407, n57408, n57409,
    n57410, n57411, n57412, n57413, n57414, n57415,
    n57416, n57417, n57418, n57419, n57420, n57421,
    n57422, n57423, n57424, n57425, n57426, n57427,
    n57428, n57429, n57431, n57432, n57433, n57434,
    n57435, n57436, n57437, n57438, n57439, n57440,
    n57441, n57442, n57443, n57444, n57445, n57446,
    n57447, n57448, n57449, n57450, n57451, n57452,
    n57453, n57454, n57455, n57456, n57457, n57458,
    n57459, n57460, n57461, n57462, n57463, n57464,
    n57465, n57466, n57467, n57468, n57469, n57470,
    n57471, n57472, n57473, n57474, n57475, n57476,
    n57477, n57478, n57480, n57481, n57482, n57483,
    n57484, n57485, n57486, n57487, n57488, n57489,
    n57490, n57491, n57492, n57493, n57494, n57495,
    n57496, n57497, n57498, n57499, n57500, n57501,
    n57502, n57503, n57504, n57505, n57506, n57507,
    n57508, n57509, n57510, n57511, n57512, n57513,
    n57514, n57515, n57516, n57517, n57518, n57519,
    n57520, n57521, n57522, n57523, n57524, n57525,
    n57526, n57527, n57529, n57530, n57531, n57532,
    n57533, n57534, n57535, n57536, n57537, n57538,
    n57539, n57540, n57541, n57542, n57543, n57544,
    n57545, n57546, n57547, n57548, n57549, n57550,
    n57551, n57552, n57553, n57554, n57555, n57556,
    n57557, n57558, n57559, n57560, n57561, n57562,
    n57563, n57564, n57565, n57566, n57567, n57568,
    n57569, n57570, n57571, n57572, n57573, n57574,
    n57575, n57576, n57578, n57579, n57580, n57581,
    n57582, n57583, n57584, n57585, n57586, n57587,
    n57588, n57589, n57590, n57591, n57592, n57593,
    n57594, n57595, n57596, n57597, n57598, n57599,
    n57600, n57601, n57602, n57603, n57604, n57605,
    n57606, n57607, n57608, n57609, n57610, n57611,
    n57612, n57613, n57614, n57615, n57616, n57617,
    n57618, n57619, n57620, n57621, n57622, n57623,
    n57624, n57625, n57626, n57627, n57628, n57629,
    n57630, n57631, n57632, n57633, n57634, n57635,
    n57636, n57637, n57638, n57639, n57640, n57641,
    n57642, n57643, n57644, n57645, n57646, n57647,
    n57648, n57649, n57650, n57651, n57652, n57653,
    n57654, n57655, n57656, n57657, n57658, n57659,
    n57660, n57661, n57662, n57663, n57664, n57665,
    n57666, n57667, n57668, n57669, n57670, n57671,
    n57672, n57673, n57674, n57675, n57676, n57677,
    n57678, n57679, n57680, n57681, n57682, n57683,
    n57684, n57685, n57686, n57687, n57688, n57689,
    n57690, n57691, n57692, n57693, n57694, n57695,
    n57696, n57697, n57698, n57699, n57700, n57701,
    n57702, n57703, n57704, n57705, n57706, n57707,
    n57708, n57709, n57710, n57711, n57712, n57713,
    n57714, n57715, n57716, n57717, n57718, n57719,
    n57720, n57721, n57722, n57723, n57724, n57725,
    n57726, n57727, n57728, n57729, n57730, n57731,
    n57732, n57733, n57734, n57735, n57736, n57737,
    n57738, n57739, n57740, n57741, n57742, n57743,
    n57744, n57745, n57746, n57747, n57748, n57749,
    n57750, n57751, n57752, n57753, n57754, n57755,
    n57756, n57757, n57758, n57759, n57760, n57761,
    n57762, n57763, n57764, n57765, n57766, n57767,
    n57768, n57769, n57770, n57771, n57772, n57773,
    n57774, n57775, n57776, n57777, n57778, n57779,
    n57780, n57781, n57782, n57783, n57784, n57785,
    n57786, n57787, n57788, n57789, n57790, n57791,
    n57792, n57793, n57794, n57795, n57796, n57797,
    n57798, n57799, n57800, n57801, n57802, n57803,
    n57804, n57805, n57806, n57807, n57808, n57809,
    n57810, n57811, n57812, n57813, n57814, n57815,
    n57816, n57817, n57818, n57819, n57820, n57821,
    n57822, n57823, n57824, n57825, n57826, n57827,
    n57828, n57829, n57830, n57831, n57832, n57833,
    n57834, n57835, n57836, n57837, n57838, n57839,
    n57840, n57841, n57842, n57843, n57844, n57845,
    n57846, n57847, n57848, n57849, n57850, n57851,
    n57852, n57853, n57854, n57855, n57856, n57857,
    n57858, n57859, n57860, n57861, n57862, n57863,
    n57864, n57865, n57866, n57867, n57868, n57869,
    n57870, n57871, n57872, n57874, n57875, n57876,
    n57877, n57878, n57879, n57880, n57881, n57882,
    n57883, n57884, n57885, n57886, n57887, n57888,
    n57889, n57890, n57891, n57892, n57893, n57894,
    n57895, n57896, n57897, n57898, n57899, n57900,
    n57901, n57902, n57903, n57904, n57905, n57906,
    n57907, n57908, n57909, n57910, n57911, n57912,
    n57913, n57914, n57915, n57916, n57917, n57918,
    n57919, n57920, n57921, n57922, n57923, n57924,
    n57925, n57926, n57927, n57928, n57929, n57930,
    n57931, n57932, n57933, n57934, n57935, n57936,
    n57937, n57938, n57939, n57940, n57941, n57942,
    n57943, n57944, n57945, n57946, n57947, n57948,
    n57949, n57951, n57952, n57953, n57954, n57955,
    n57956, n57957, n57958, n57959, n57960, n57961,
    n57962, n57963, n57964, n57965, n57966, n57967,
    n57968, n57969, n57970, n57971, n57972, n57973,
    n57974, n57975, n57976, n57977, n57978, n57979,
    n57980, n57981, n57982, n57983, n57984, n57985,
    n57986, n57987, n57988, n57989, n57990, n57991,
    n57992, n57993, n57994, n57995, n57996, n57997,
    n57998, n57999, n58000, n58001, n58002, n58003,
    n58004, n58005, n58006, n58007, n58008, n58009,
    n58010, n58011, n58012, n58013, n58014, n58015,
    n58016, n58017, n58018, n58019, n58020, n58021,
    n58022, n58023, n58024, n58025, n58026, n58027,
    n58028, n58029, n58031, n58032, n58033, n58034,
    n58035, n58036, n58037, n58038, n58039, n58040,
    n58041, n58042, n58043, n58044, n58045, n58046,
    n58047, n58048, n58049, n58050, n58051, n58052,
    n58053, n58054, n58055, n58056, n58057, n58058,
    n58059, n58060, n58061, n58062, n58063, n58065,
    n58066, n58067, n58068, n58069, n58071, n58072,
    n58074, n58075, n58076, n58077, n58079, n58080,
    n58081, n58083, n58084, n58086, n58087, n58088,
    n58089, n58090, n58091, n58092, n58094, n58095,
    n58097, n58098, n58099, n58100, n58101, n58102,
    n58103, n58104, n58105, n58106, n58107, n58108,
    n58109, n58110, n58111, n58112, n58113, n58114,
    n58115, n58116, n58117, n58118, n58119, n58120,
    n58121, n58122, n58123, n58124, n58125, n58126,
    n58127, n58128, n58129, n58130, n58131, n58132,
    n58133, n58134, n58135, n58136, n58137, n58138,
    n58139, n58140, n58141, n58142, n58143, n58144,
    n58145, n58146, n58147, n58148, n58149, n58150,
    n58151, n58152, n58153, n58154, n58155, n58156,
    n58157, n58158, n58159, n58160, n58161, n58162,
    n58163, n58164, n58165, n58166, n58167, n58168,
    n58169, n58170, n58171, n58172, n58173, n58174,
    n58175, n58176, n58177, n58178, n58179, n58180,
    n58181, n58182, n58183, n58184, n58185, n58186,
    n58187, n58188, n58189, n58190, n58191, n58192,
    n58193, n58194, n58195, n58196, n58197, n58198,
    n58199, n58200, n58201, n58202, n58203, n58204,
    n58205, n58206, n58207, n58208, n58209, n58210,
    n58211, n58212, n58213, n58214, n58215, n58217,
    n58218, n58219, n58220, n58221, n58222, n58223,
    n58224, n58225, n58226, n58227, n58228, n58229,
    n58230, n58231, n58232, n58233, n58234, n58235,
    n58236, n58237, n58238, n58239, n58240, n58241,
    n58242, n58243, n58244, n58245, n58246, n58247,
    n58248, n58249, n58250, n58251, n58252, n58254,
    n58255, n58257, n58258, n58259, n58260, n58261,
    n58262, n58263, n58264, n58265, n58266, n58267,
    n58268, n58269, n58271, n58272, n58273, n58274,
    n58275, n58276, n58277, n58278, n58279, n58280,
    n58281, n58282, n58283, n58284, n58285, n58287,
    n58288, n58289, n58290, n58291, n58292, n58293,
    n58294, n58295, n58296, n58297, n58298, n58299,
    n58300, n58301, n58302, n58303, n58304, n58305,
    n58306, n58307, n58308, n58310, n58311, n58312,
    n58313, n58314, n58315, n58316, n58317, n58318,
    n58319, n58320, n58321, n58322, n58323, n58324,
    n58325, n58326, n58327, n58328, n58329, n58330,
    n58331, n58332, n58333, n58334, n58335, n58336,
    n58337, n58338, n58339, n58340, n58341, n58342,
    n58343, n58344, n58345, n58346, n58347, n58348,
    n58349, n58350, n58351, n58352, n58353, n58354,
    n58355, n58356, n58357, n58358, n58359, n58361,
    n58362, n58363, n58364, n58365, n58366, n58367,
    n58368, n58370, n58371, n58372, n58373, n58374,
    n58375, n58376, n58377, n58378, n58379, n58380,
    n58382, n58383, n58384, n58385, n58386, n58387,
    n58388, n58389, n58391, n58392, n58393, n58394,
    n58395, n58397, n58398, n58399, n58400, n58401,
    n58402, n58404, n58405, n58406, n58407, n58408,
    n58409, n58410, n58411, n58412, n58413, n58414,
    n58415, n58416, n58417, n58418, n58419, n58420,
    n58421, n58422, n58423, n58424, n58425, n58426,
    n58427, n58428, n58429, n58430, n58431, n58432,
    n58433, n58434, n58435, n58436, n58437, n58438,
    n58439, n58440, n58441, n58442, n58443, n58444,
    n58445, n58446, n58447, n58448, n58449, n58450,
    n58451, n58452, n58453, n58454, n58455, n58456,
    n58457, n58458, n58459, n58460, n58461, n58462,
    n58463, n58464, n58465, n58466, n58467, n58468,
    n58469, n58470, n58471, n58472, n58473, n58474,
    n58475, n58476, n58477, n58478, n58479, n58480,
    n58481, n58482, n58483, n58484, n58485, n58486,
    n58487, n58488, n58489, n58490, n58491, n58492,
    n58493, n58494, n58495, n58496, n58497, n58498,
    n58499, n58500, n58501, n58502, n58503, n58504,
    n58505, n58506, n58507, n58508, n58509, n58510,
    n58511, n58512, n58513, n58514, n58515, n58516,
    n58517, n58518, n58519, n58520, n58521, n58522,
    n58523, n58524, n58525, n58526, n58527, n58528,
    n58529, n58530, n58531, n58532, n58533, n58534,
    n58535, n58536, n58537, n58538, n58539, n58540,
    n58541, n58542, n58543, n58544, n58545, n58546,
    n58547, n58548, n58549, n58550, n58551, n58552,
    n58553, n58554, n58555, n58556, n58557, n58558,
    n58559, n58560, n58561, n58562, n58563, n58564,
    n58565, n58566, n58567, n58568, n58569, n58570,
    n58571, n58572, n58573, n58574, n58575, n58576,
    n58577, n58578, n58579, n58580, n58581, n58582,
    n58583, n58584, n58585, n58586, n58587, n58588,
    n58589, n58590, n58591, n58592, n58593, n58594,
    n58595, n58596, n58597, n58598, n58599, n58600,
    n58601, n58602, n58603, n58604, n58605, n58606,
    n58607, n58608, n58609, n58610, n58611, n58612,
    n58613, n58614, n58615, n58616, n58617, n58618,
    n58619, n58620, n58621, n58622, n58623, n58624,
    n58625, n58626, n58627, n58628, n58629, n58630,
    n58631, n58632, n58633, n58634, n58635, n58636,
    n58637, n58638, n58639, n58640, n58641, n58642,
    n58643, n58644, n58645, n58646, n58647, n58648,
    n58649, n58650, n58651, n58652, n58653, n58654,
    n58655, n58656, n58657, n58658, n58659, n58660,
    n58661, n58662, n58663, n58664, n58665, n58666,
    n58667, n58668, n58669, n58670, n58671, n58672,
    n58673, n58674, n58675, n58676, n58677, n58678,
    n58679, n58680, n58681, n58682, n58683, n58684,
    n58685, n58686, n58687, n58688, n58689, n58690,
    n58691, n58692, n58693, n58694, n58695, n58696,
    n58697, n58698, n58699, n58700, n58701, n58702,
    n58703, n58704, n58705, n58706, n58707, n58708,
    n58709, n58710, n58711, n58712, n58713, n58714,
    n58715, n58716, n58717, n58718, n58720, n58721,
    n58722, n58723, n58724, n58725, n58726, n58727,
    n58728, n58729, n58730, n58731, n58732, n58733,
    n58734, n58735, n58736, n58737, n58738, n58739,
    n58740, n58741, n58742, n58743, n58744, n58745,
    n58746, n58747, n58748, n58749, n58750, n58751,
    n58752, n58753, n58754, n58755, n58756, n58757,
    n58758, n58759, n58760, n58761, n58763, n58764,
    n58765, n58766, n58767, n58768, n58781, n58782,
    n58783, n58784, n58785, n58786, n58787, n58788,
    n58789, n58790, n58791, n58792, n58793, n58794,
    n58795, n58796, n58797, n58798, n58799, n58800,
    n58801, n58802, n58803, n58804, n58805, n58806,
    n58807, n58808, n58809, n58810, n58811, n58812,
    n58813, n58814, n58815, n58816, n58817, n58818,
    n58819, n58820, n58821, n58822, n58823, n58824,
    n58825, n58826, n58827, n58828, n58829, n58830,
    n58831, n58832, n58833, n58834, n58835, n58836,
    n58837, n58838, n58839, n58840, n58841, n58842,
    n58843, n58844, n58845, n58846, n58847, n58848,
    n58849, n58850, n58851, n58852, n58853, n58854,
    n58855, n58856, n58857, n58858, n58859, n58860,
    n58861, n58862, n58863, n58864, n58865, n58866,
    n58867, n58868, n58869, n58870, n58871, n58872,
    n58873, n58874, n58875, n58876, n58877, n58878,
    n58879, n58880, n58881, n58882, n58883, n58884,
    n58885, n58886, n58887, n58888, n58889, n58890,
    n58891, n58892, n58893, n58894, n58895, n58896,
    n58897, n58898, n58899, n58900, n58901, n58902,
    n58903, n58904, n58905, n58906, n58907, n58908,
    n58909, n58910, n58911, n58912, n58913, n58914,
    n58915, n58916, n58917, n58918, n58919, n58920,
    n58921, n58922, n58923, n58924, n58925, n58926,
    n58927, n58928, n58929, n58930, n58931, n58932,
    n58933, n58934, n58935, n58936, n58937, n58938,
    n58939, n58940, n58941, n58942, n58943, n58944,
    n58945, n58946, n58947, n58948, n58949, n58950,
    n58951, n58952, n58953, n58954, n58955, n58956,
    n58957, n58958, n58959, n58960, n58961, n58962,
    n58963, n58964, n58965, n58966, n58967, n58968,
    n58969, n58970, n58971, n58972, n58973, n58974,
    n58975, n58976, n58977, n58978, n58979, n58980,
    n58981, n58982, n58983, n58984, n58985, n58986,
    n58987, n58988, n58989, n58990, n58991, n58992,
    n58993, n58994, n58995, n58996, n58997, n58998,
    n58999, n59000, n59001, n59002, n59003, n59004,
    n59005, n59006, n59007, n59008, n59009, n59010,
    n59011, n59012, n59013, n59014, n59015, n59016,
    n59017, n59018, n59019, n59020, n59021, n59022,
    n59023, n59024, n59025, n59026, n59027, n59028,
    n59029, n59030, n59031, n59032, n59033, n59034,
    n59035, n59036, n59037, n59038, n59039, n59040,
    n59041, n59042, n59043, n59044, n59045, n59046,
    n59047, n59048, n59049, n59050, n59051, n59052,
    n59053, n59054, n59055, n59056, n59057, n59058,
    n59059, n59060, n59061, n59062, n59063, n59064,
    n59065, n59066, n59067, n59068, n59069, n59070,
    n59071, n59072, n59073, n59074, n59075, n59076,
    n59077, n59078, n59079, n59080, n59081, n59082,
    n59083, n59084, n59085, n59086, n59087, n59088,
    n59089, n59090, n59091, n59092, n59093, n59094,
    n59095, n59096, n59097, n59098, n59099, n59100,
    n59101, n59102, n59103, n59104, n59105, n59106,
    n59107, n59108, n59109, n59110, n59111, n59112,
    n59113, n59114, n59115, n59116, n59117, n59118,
    n59119, n59120, n59121, n59122, n59123, n59124,
    n59125, n59126, n59127, n59128, n59129, n59130,
    n59131, n59132, n59133, n59134, n59135, n59136,
    n59137, n59138, n59139, n59140, n59141, n59142,
    n59143, n59144, n59145, n59146, n59147, n59148,
    n59149, n59150, n59151, n59152, n59153, n59154,
    n59155, n59156, n59157, n59158, n59159, n59160,
    n59161, n59162, n59163, n59164, n59165, n59166,
    n59167, n59168, n59169, n59170, n59171, n59172,
    n59173, n59174, n59175, n59176, n59177, n59178,
    n59179, n59180, n59181, n59182, n59183, n59184,
    n59185, n59186, n59187, n59188, n59189, n59190,
    n59191, n59192, n59193, n59194, n59195, n59196,
    n59197, n59198, n59199, n59200, n59201, n59202,
    n59203, n59204, n59205, n59206, n59207, n59208,
    n59209, n59210, n59211, n59212, n59213, n59214,
    n59215, n59216, n59217, n59218, n59219, n59220,
    n59221, n59222, n59223, n59224, n59225, n59226,
    n59227, n59228, n59229, n59230, n59231, n59232,
    n59233, n59234, n59235, n59236, n59237, n59238,
    n59239, n59240, n59241, n59242, n59243, n59244,
    n59245, n59246, n59247, n59248, n59249, n59250,
    n59251, n59252, n59253, n59254, n59255, n59256,
    n59257, n59258, n59259, n59260, n59261, n59262,
    n59263, n59264, n59265, n59266, n59267, n59268,
    n59269, n59270, n59271, n59272, n59273, n59274,
    n59275, n59276, n59277, n59278, n59279, n59280,
    n59281, n59282, n59283, n59284, n59285, n59286,
    n59287, n59288, n59289, n59290, n59291, n59292,
    n59293, n59294, n59295, n59296, n59297, n59298,
    n59299, n59300, n59301, n59302, n59303, n59304,
    n59305, n59306, n59307, n59308, n59309, n59310,
    n59311, n59312, n59313, n59314, n59315, n59316,
    n59317, n59318, n59319, n59320, n59321, n59322,
    n59323, n59324, n59325, n59326, n59327, n59328,
    n59329, n59330, n59331, n59332, n59333, n59334,
    n59335, n59336, n59337, n59338, n59339, n59340,
    n59341, n59342, n59343, n59344, n59345, n59346,
    n59347, n59348, n59349, n59350, n59351, n59352,
    n59353, n59354, n59355, n59356, n59357, n59358,
    n59359, n59360, n59361, n59362, n59363, n59364,
    n59365, n59366, n59367, n59368, n59369, n59370,
    n59371, n59372, n59373, n59374, n59375, n59376,
    n59377, n59378, n59379, n59380, n59381, n59382,
    n59383, n59384, n59385, n59386, n59387, n59388,
    n59389, n59390, n59391, n59392, n59393, n59394,
    n59395, n59396, n59397, n59398, n59399, n59400,
    n59401, n59402, n59403, n59404, n59405, n59406,
    n59407, n59408, n59409, n59410, n59411, n59412,
    n59413, n59414, n59415, n59416, n59417, n59418,
    n59419, n59420, n59421, n59422, n59423, n59424,
    n59425, n59426, n59427, n59428, n59429, n59430,
    n59431, n59432, n59433, n59434, n59435, n59436,
    n59437, n59438, n59439, n59440, n59441, n59442,
    n59443, n59444, n59445, n59446, n59447, n59448,
    n59449, n59450, n59451, n59452, n59453, n59454,
    n59455, n59456, n59457, n59458, n59459, n59460,
    n59461, n59462, n59463, n59464, n59465, n59466,
    n59467, n59468, n59469, n59470, n59471, n59472,
    n59473, n59474, n59475, n59476, n59477, n59478,
    n59479, n59480, n59481, n59482, n59483, n59484,
    n59485, n59486, n59487, n59488, n59489, n59490,
    n59491, n59492, n59493, n59494, n59495, n59496,
    n59497, n59498, n59499, n59500, n59501, n59502,
    n59503, n59504, n59505, n59506, n59507, n59508,
    n59509, n59510, n59511, n59512, n59513, n59514,
    n59515, n59516, n59517, n59518, n59519, n59520,
    n59521, n59522, n59523, n59524, n59525, n59526,
    n59527, n59528, n59529, n59530, n59531, n59532,
    n59533, n59534, n59535, n59536, n59537, n59538,
    n59539, n59540, n59541, n59542, n59543, n59544,
    n59545, n59546, n59547, n59548, n59549, n59550,
    n59551, n59552, n59553, n59554, n59555, n59556,
    n59557, n59558, n59559, n59560, n59561, n59562,
    n59563, n59564, n59565, n59566, n59567, n59568,
    n59569, n59570, n59571, n59572, n59573, n59574,
    n59575, n59576, n59577, n59578, n59579, n59580,
    n59581, n59582, n59583, n59584, n59585, n59586,
    n59587, n59588, n59589, n59590, n59591, n59592,
    n59593, n59594, n59595, n59596, n59597, n59598,
    n59599, n59600, n59601, n59602, n59603, n59604,
    n59605, n59606, n59607, n59608, n59609, n59610,
    n59611, n59612, n59613, n59614, n59615, n59616,
    n59617, n59618, n59619, n59620, n59621, n59622,
    n59623, n59624, n59625, n59626, n59627, n59628,
    n59629, n59630, n59631, n59632, n59633, n59634,
    n59635, n59636, n59637, n59638, n59639, n59640,
    n59641, n59642, n59643, n59644, n59645, n59646,
    n59647, n59648, n59649, n59650, n59651, n59652,
    n59653, n59654, n59655, n59656, n59657, n59658,
    n59659, n59660, n59661, n59662, n59663, n59664,
    n59665, n59666, n59667, n59668, n59669, n59670,
    n59671, n59672, n59673, n59674, n59675, n59676,
    n59677, n59678, n59679, n59680, n59681, n59682,
    n59683, n59684, n59685, n59686, n59687, n59688,
    n59689, n59690, n59691, n59692, n59693, n59694,
    n59695, n59696, n59697, n59698, n59699, n59700,
    n59701, n59702, n59703, n59704, n59705, n59706,
    n59707, n59708, n59709, n59710, n59711, n59712,
    n59713, n59714, n59715, n59716, n59717, n59718,
    n59719, n59720, n59721, n59722, n59723, n59724,
    n59725, n59726, n59727, n59728, n59729, n59730,
    n59731, n59732, n59733, n59734, n59735, n59736,
    n59737, n59738, n59739, n59740, n59741, n59742,
    n59743, n59744, n59745, n59746, n59747, n59748,
    n59749, n59750, n59751, n59752, n59753, n59754,
    n59755, n59756, n59757, n59758, n59759, n59760,
    n59761, n59762, n59763, n59764, n59765, n59766,
    n59767, n59768, n59769, n59770, n59771, n59772,
    n59773, n59774, n59775, n59776, n59777, n59778,
    n59779, n59780, n59781, n59782, n59783, n59784,
    n59785, n59786, n59787, n59788, n59789, n59790,
    n59791, n59792, n59793, n59794, n59795, n59796,
    n59797, n59798, n59799, n59800, n59801, n59802,
    n59803, n59804, n59805, n59806, n59807, n59808,
    n59809, n59810, n59811, n59812, n59813, n59814,
    n59815, n59816, n59817, n59818, n59819, n59820,
    n59821, n59822, n59823, n59824, n59825, n59826,
    n59827, n59828, n59829, n59830, n59831, n59832,
    n59833, n59834, n59835, n59836, n59837, n59838,
    n59839, n59840, n59841, n59842, n59843, n59844,
    n59845, n59846, n59847, n59848, n59849, n59850,
    n59851, n59852, n59853, n59854, n59855, n59856,
    n59857, n59858, n59859, n59860, n59861, n59862,
    n59863, n59864, n59865, n59866, n59867, n59868,
    n59869, n59870, n59871, n59872, n59873, n59874,
    n59875, n59876, n59877, n59878, n59879, n59880,
    n59882, n59883, n59884, n59885, n59886, n59887,
    n59888, n59889, n59890, n59891, n59892, n59893,
    n59894, n59895, n59896, n59897, n59898, n59899,
    n59900, n59901, n59902, n59903, n59904, n59905,
    n59906, n59907, n59908, n59909, n59910, n59911,
    n59912, n59913, n59914, n59915, n59916, n59917,
    n59918, n59919, n59920, n59921, n59922, n59923,
    n59924, n59925, n59926, n59927, n59928, n59929,
    n59930, n59931, n59932, n59933, n59934, n59935,
    n59936, n59937, n59938, n59939, n59940, n59941,
    n59942, n59943, n59944, n59945, n59946, n59947,
    n59948, n59949, n59950, n59951, n59952, n59953,
    n59954, n59955, n59956, n59957, n59958, n59959,
    n59960, n59961, n59962, n59963, n59964, n59965,
    n59966, n59967, n59968, n59969, n59970, n59971,
    n59972, n59973, n59974, n59975, n59976, n59977,
    n59978, n59979, n59980, n59981, n59982, n59983,
    n59984, n59985, n59986, n59987, n59988, n59989,
    n59990, n59991, n59992, n59993, n59994, n59995,
    n59996, n59997, n59998, n59999, n60000, n60001,
    n60002, n60004, n60005, n60006, n60007, n60008,
    n60009, n60010, n60011, n60012, n60013, n60014,
    n60015, n60016, n60017, n60018, n60019, n60020,
    n60021, n60022, n60023, n60024, n60025, n60026,
    n60027, n60028, n60029, n60030, n60031, n60032,
    n60033, n60034, n60036, n60037, n60038, n60039,
    n60040, n60041, n60042, n60043, n60044, n60045,
    n60046, n60047, n60048, n60049, n60050, n60051,
    n60052, n60053, n60054, n60055, n60056, n60057,
    n60058, n60059, n60060, n60061, n60062, n60063,
    n60064, n60065, n60066, n60067, n60068, n60069,
    n60070, n60071, n60072, n60073, n60074, n60075,
    n60076, n60077, n60078, n60079, n60080, n60081,
    n60082, n60083, n60084, n60085, n60086, n60087,
    n60088, n60089, n60090, n60091, n60092, n60093,
    n60094, n60095, n60096, n60097, n60098, n60099,
    n60100, n60101, n60102, n60103, n60104, n60105,
    n60106, n60107, n60108, n60109, n60110, n60111,
    n60112, n60113, n60114, n60115, n60116, n60117,
    n60118, n60119, n60120, n60121, n60122, n60123,
    n60124, n60125, n60126, n60127, n60128, n60129,
    n60130, n60131, n60132, n60133, n60134, n60135,
    n60136, n60137, n60138, n60139, n60140, n60141,
    n60142, n60143, n60144, n60145, n60146, n60147,
    n60148, n60149, n60150, n60151, n60152, n60153,
    n60154, n60155, n60156, n60157, n60158, n60159,
    n60160, n60161, n60162, n60163, n60164, n60165,
    n60166, n60167, n60168, n60169, n60170, n60171,
    n60172, n60173, n60174, n60175, n60176, n60177,
    n60178, n60179, n60180, n60181, n60182, n60183,
    n60184, n60185, n60186, n60187, n60188, n60189,
    n60190, n60191, n60192, n60193, n60194, n60195,
    n60196, n60197, n60198, n60199, n60200, n60201,
    n60202, n60203, n60204, n60205, n60206, n60207,
    n60208, n60209, n60210, n60211, n60212, n60213,
    n60214, n60215, n60216, n60217, n60218, n60219,
    n60220, n60221, n60222, n60223, n60224, n60225,
    n60226, n60227, n60228, n60229, n60230, n60231,
    n60232, n60233, n60234, n60235, n60236, n60237,
    n60238, n60239, n60240, n60241, n60242, n60243,
    n60244, n60245, n60246, n60247, n60248, n60249,
    n60250, n60251, n60252, n60253, n60254, n60255,
    n60256, n60257, n60258, n60259, n60260, n60261,
    n60262, n60263, n60264, n60265, n60266, n60267,
    n60268, n60269, n60270, n60271, n60272, n60273,
    n60274, n60275, n60276, n60277, n60278, n60279,
    n60280, n60281, n60282, n60283, n60284, n60285,
    n60286, n60287, n60288, n60289, n60290, n60291,
    n60292, n60293, n60294, n60295, n60296, n60297,
    n60298, n60299, n60300, n60301, n60302, n60303,
    n60304, n60305, n60306, n60307, n60308, n60309,
    n60310, n60311, n60312, n60313, n60314, n60315,
    n60316, n60317, n60318, n60319, n60320, n60321,
    n60322, n60323, n60324, n60325, n60326, n60327,
    n60328, n60329, n60330, n60331, n60332, n60333,
    n60334, n60335, n60336, n60337, n60338, n60339,
    n60340, n60341, n60342, n60343, n60344, n60345,
    n60346, n60347, n60348, n60349, n60350, n60351,
    n60352, n60353, n60354, n60355, n60356, n60357,
    n60358, n60359, n60360, n60361, n60362, n60363,
    n60364, n60365, n60366, n60367, n60368, n60369,
    n60370, n60371, n60372, n60373, n60374, n60375,
    n60376, n60377, n60378, n60379, n60380, n60381,
    n60382, n60383, n60384, n60385, n60386, n60387,
    n60388, n60389, n60390, n60391, n60392, n60393,
    n60394, n60395, n60396, n60397, n60398, n60399,
    n60400, n60401, n60402, n60403, n60404, n60405,
    n60406, n60407, n60408, n60409, n60410, n60411,
    n60412, n60413, n60414, n60415, n60416, n60417,
    n60418, n60419, n60420, n60421, n60422, n60423,
    n60424, n60425, n60426, n60427, n60428, n60429,
    n60430, n60431, n60432, n60433, n60434, n60435,
    n60436, n60437, n60438, n60439, n60440, n60441,
    n60442, n60443, n60444, n60445, n60446, n60447,
    n60448, n60449, n60450, n60451, n60452, n60453,
    n60454, n60455, n60456, n60457, n60458, n60459,
    n60460, n60461, n60462, n60463, n60464, n60465,
    n60466, n60467, n60468, n60469, n60470, n60471,
    n60472, n60473, n60474, n60475, n60476, n60477,
    n60478, n60480, n60481, n60482, n60483, n60484,
    n60485, n60486, n60487, n60488, n60489, n60490,
    n60491, n60492, n60493, n60494, n60495, n60496,
    n60497, n60498, n60499, n60500, n60501, n60502,
    n60503, n60504, n60505, n60506, n60507, n60508,
    n60509, n60510, n60511, n60512, n60513, n60514,
    n60515, n60516, n60517, n60518, n60519, n60520,
    n60521, n60522, n60523, n60524, n60525, n60526,
    n60527, n60528, n60529, n60530, n60531, n60532,
    n60533, n60534, n60535, n60536, n60537, n60538,
    n60539, n60541, n60542, n60543, n60544, n60545,
    n60546, n60547, n60548, n60549, n60550, n60551,
    n60552, n60553, n60554, n60555, n60556, n60557,
    n60558, n60559, n60560, n60561, n60562, n60563,
    n60564, n60565, n60566, n60567, n60569, n60570,
    n60571, n60572, n60573, n60574, n60575, n60576,
    n60577, n60578, n60579, n60580, n60581, n60582,
    n60583, n60584, n60585, n60586, n60587, n60588,
    n60589, n60590, n60591, n60592, n60593, n60594,
    n60595, n60596, n60597, n60598, n60599, n60600,
    n60601, n60602, n60603, n60604, n60605, n60606,
    n60607, n60608, n60609, n60610, n60611, n60612,
    n60613, n60614, n60615, n60616, n60617, n60618,
    n60619, n60620, n60621, n60622, n60623, n60624,
    n60625, n60626, n60627, n60628, n60629, n60630,
    n60631, n60632, n60633, n60634, n60635, n60636,
    n60637, n60638, n60639, n60640, n60641, n60642,
    n60643, n60644, n60645, n60646, n60647, n60648,
    n60649, n60650, n60651, n60652, n60653, n60654,
    n60655, n60656, n60657, n60658, n60659, n60660,
    n60661, n60662, n60663, n60664, n60665, n60666,
    n60667, n60668, n60669, n60670, n60671, n60672,
    n60673, n60674, n60675, n60676, n60677, n60678,
    n60679, n60680, n60681, n60682, n60683, n60684,
    n60685, n60686, n60687, n60688, n60689, n60691,
    n60692, n60693, n60694, n60695, n60696, n60697,
    n60698, n60699, n60700, n60701, n60702, n60703,
    n60704, n60705, n60706, n60707, n60708, n60709,
    n60710, n60711, n60712, n60713, n60714, n60715,
    n60716, n60717, n60718, n60719, n60720, n60721,
    n60722, n60723, n60724, n60725, n60726, n60727,
    n60728, n60730, n60731, n60732, n60733, n60734,
    n60735, n60736, n60737, n60739, n60740, n60741,
    n60742, n60743, n60744, n60745, n60746, n60747,
    n60748, n60749, n60750, n60751, n60752, n60754,
    n60755, n60756, n60757, n60758, n60759, n60760,
    n60761, n60763, n60764, n60765, n60766, n60767,
    n60768, n60769, n60770, n60771, n60772, n60773,
    n60774, n60775, n60776, n60777, n60778, n60779,
    n60780, n60781, n60782, n60783, n60784, n60785,
    n60786, n60787, n60788, n60789, n60790, n60791,
    n60792, n60793, n60794, n60795, n60796, n60797,
    n60798, n60799, n60800, n60801, n60802, n60803,
    n60804, n60805, n60806, n60807, n60808, n60809,
    n60812, n60813, n60814, n60815, n60816, n60817,
    n60818, n60819, n60820, n60821, n60822, n60823,
    n60824, n60825, n60826, n60827, n60828, n60829,
    n60830, n60831, n60832, n60833, n60834, n60835,
    n60836, n60837, n60838, n60839, n60840, n60841,
    n60842, n60843, n60844, n60846, n60847, n60848,
    n60850, n60851, n60852, n60853, n60854, n60855,
    n60856, n60859, n60860, n60861, n60862, n60863,
    n60865, n60867, n60870, n60871, n60872, n60873,
    n60874, n60879, n60880, n60881, n60882, n60883,
    n60885, n60890, n60891, n60892, n60893, n60894,
    n60895, n60896, n60897, n60898, n60899, n60900,
    n60901, n60902, n60903, n60904, n60905, n60906,
    n60907, n60908, n60909, n60910, n60911, n60912,
    n60913, n60914, n60915, n60916, n60917, n60918,
    n60919, n60920, n60921, n60922, n60923, n60924,
    n60925, n60926, n60927, n60928, n60929, n60930,
    n60931, n60932, n60933, n60934, n60935, n60936,
    n60937, n60938, n60939, n60940, n60941, n60942,
    n60943, n60944, n60945, n60946, n60947, n60948,
    n60949, n60950, n60951, n60952, n60953, n60954,
    n60955, n60956, n60957, n60958, n60959, n60960,
    n60961, n60962, n60963, n60964, n60965, n60966,
    n60967, n60968, n60969, n60970, n60971, n60972,
    n60973, n60974, n60975, n60976, n60977, n60978,
    n60979, n60980, n60981, n60982, n60983, n60984,
    n60985, n60986, n60987, n60988, n60989, n60990,
    n60991, n60992, n60993, n60994, n60995, n60996,
    n60997, n60998, n60999, n61000, n61001, n61002,
    n61003, n61004, n61005, n61006, n61007, n61008,
    n61009, n61010, n61011, n61012, n61013, n61014,
    n61015, n61016, n61017, n61018, n61019, n61020,
    n61021, n61022, n61023, n61024, n61025, n61026,
    n61027, n61028, n61029, n61030, n61031, n61032,
    n61033, n61034, n61035, n61036, n61037, n61038,
    n61039, n61040, n61041, n61042, n61043, n61044,
    n61045, n61046, n61047, n61048, n61049, n61050,
    n61051, n61052, n61053, n61054, n61055, n61056,
    n61057, n61058, n61059, n61060, n61061, n61062,
    n61063, n61064, n61065, n61066, n61067, n61081,
    n61082, n61083, n61084, n61085, n61086, n61087,
    n61088, n61089, n61090, n61091, n61092, n61093,
    n61094, n61095, n61096, n61097, n61098, n61099,
    n61100, n61101, n61102, n61103, n61104, n61105,
    n61106, n61107, n61108, n61109, n61110, n61111,
    n61112, n61113, n61114, n61115, n61116, n61117,
    n61118, n61119, n61120, n61121, n61122, n61123,
    n61124, n61125, n61126, n61127, n61128, n61129,
    n61130, n61131, n61132, n61133, n61134, n61135,
    n61136, n61137, n61138, n61139, n61140, n61141,
    n61142, n61143, n61144, n61145, n61146, n61147,
    n61148, n61149, n61150, n61151, n61152, n61153,
    n61154, n61155, n61156, n61157, n61158, n61159,
    n61160, n61161, n61162, n61163, n61164, n61165,
    n61166, n61167, n61168, n61169, n61170, n61171,
    n61172, n61173, n61174, n61175, n61176, n61177,
    n61178, n61179, n61180, n61181, n61182, n61183,
    n61184, n61185, n61186, n61187, n61188, n61189,
    n61190, n61191, n61192, n61193, n61194, n61195,
    n61196, n61197, n61198, n61199, n61200, n61201,
    n61202, n61203, n61204, n61205, n61206, n61207,
    n61208, n61209, n61210, n61211, n61212, n61213,
    n61214, n61215, n61216, n61217, n61218, n61219,
    n61220, n61221, n61222, n61223, n61224, n61225,
    n61226, n61227, n61228, n61230, n61231, n61232,
    n61233, n61234, n61235, n61236, n61237, n61238,
    n61239, n61240, n61241, n61242, n61243, n61244,
    n61245, n61246, n61247, n61248, n61249, n61250,
    n61251, n61252, n61254, n61255, n61256, n61257,
    n61258, n61259, n61260, n61261, n61262, n61263,
    n61264, n61265, n61266, n61267, n61268, n61269,
    n61270, n61271, n61272, n61273, n61274, n61275,
    n61276, n61277, n61278, n61280, n61281, n61282,
    n61283, n61284, n61285, n61286, n61287, n61288,
    n61289, n61290, n61291, n61292, n61293, n61294,
    n61295, n61296, n61297, n61298, n61299, n61300,
    n61302, n61303, n61304, n61305, n61306, n61307,
    n61308, n61309, n61310, n61311, n61312, n61314,
    n61315, n61316, n61317, n61318, n61319, n61320,
    n61321, n61322, n61323, n61324, n61325, n61326,
    n61327, n61329, n61330, n61331, n61332, n61333,
    n61334, n61335, n61336, n61337, n61338, n61340,
    n61341, n61342, n61343, n61344, n61345, n61346,
    n61347, n61348, n61349, n61350, n61351, n61352,
    n61353, n61354, n61355, n61356, n61357, n61358,
    n61359, n61360, n61361, n61362, n61363, n61364,
    n61365, n61366, n61367, n61368, n61369, n61370,
    n61371, n61372, n61373, n61374, n61375, n61376,
    n61377, n61378, n61379, n61380, n61381, n61382,
    n61383, n61384, n61385, n61386, n61387, n61388,
    n61389, n61390, n61391, n61393, n61394, n61395,
    n61396, n61397, n61398, n61399, n61400, n61401,
    n61402, n61403, n61407, n61409, n61410, n61411,
    n61412, n61413, n61414, n61415, n61416, n61417,
    n61419, n61420, n61425, n61426, n61427, n61428,
    n61429, n61430, n61431, n61432, n61433, n61434,
    n61435, n61436, n61437, n61438, n61439, n61440,
    n61441, n61442, n61443, n61444, n61445, n61446,
    n61447, n61448, n61449, n61450, n61451, n61452,
    n61453, n61454, n61455, n61456, n61457, n61458,
    n61459, n61460, n61461, n61462, n61463, n61464,
    n61465, n61466, n61467, n61468, n61547, n61548,
    n61549, n61550, n61551, n61552, n61553, n61554,
    n61555, n61556, n61557, n61558, n61559, n61560,
    n61561, n61562, n61563, n61564, n61565, n61566,
    n61567, n61568, n61569, n61570, n61571, n61572,
    n61573, n61574, n61575, n61576, n61577, n61579,
    n61580, n61581, n61598, n61599, n61600, n61601,
    n61602, n61603, n61604, n61605, n61606, n61607,
    n61608, n61609, n61610, n61611, n61612, n61613,
    n61614, n61615, n61616, n61617, n61618, n61619,
    n61630, n61631, n61632, n61633, n61634, n61635,
    n61636, n61637, n61638, n61639, n61641, n61645,
    n61646, n61647, n61648, n61649, n61650, n61651,
    n61652, n61654, n61655, n61656, n61657, n61658,
    n61659, n61660, n61661, n61662, n61663, n61664,
    n61665, n61666, n61667, n61668, n61669, n61670,
    n61671, n61672, n61673, n61674, n61675, n61676,
    n61677, n61678, n61679, n61680, n61681, n61682,
    n61683, n61684, n61685, n61686, n61687, n61688,
    n61689, n61690, n61691, n61692, n61693, n61694,
    n61695, n61696, n61697;
  assign po166 = 1'b1;
  assign n2437 = pi351 & pi1199;
  assign n2438 = ~pi54 & ~pi92;
  assign n2439 = ~pi74 & n2438;
  assign n2440 = ~pi122 & pi829;
  assign n2441 = pi950 & pi1092;
  assign n2442 = ~pi824 & ~pi829;
  assign n2443 = n2441 & ~n2442;
  assign n2444 = ~pi35 & ~pi70;
  assign n2445 = ~pi58 & ~pi90;
  assign n2446 = ~pi63 & ~pi107;
  assign n2447 = ~pi83 & ~pi103;
  assign n2448 = ~pi61 & ~pi76;
  assign n2449 = ~pi85 & ~pi106;
  assign n2450 = n2448 & n2449;
  assign n2451 = ~pi48 & n2450;
  assign n2452 = ~pi89 & n2451;
  assign n2453 = ~pi49 & n2452;
  assign n2454 = ~pi104 & n2453;
  assign n2455 = ~pi45 & n2454;
  assign n2456 = ~pi68 & ~pi84;
  assign n2457 = ~pi82 & ~pi111;
  assign n2458 = ~pi36 & n2457;
  assign n2459 = n2456 & n2458;
  assign n2460 = ~pi66 & ~pi73;
  assign n2461 = n2459 & n2460;
  assign n2462 = n2455 & n2459;
  assign n2463 = n2460 & n2462;
  assign n2464 = n2455 & n2461;
  assign n2465 = ~pi67 & ~pi69;
  assign n2466 = ~pi67 & n58781;
  assign n2467 = ~pi69 & n2466;
  assign n2468 = n58781 & n2465;
  assign n2469 = n2447 & n58782;
  assign n2470 = ~pi88 & ~pi98;
  assign n2471 = ~pi50 & ~pi77;
  assign n2472 = ~pi77 & n2470;
  assign n2473 = ~pi50 & n2472;
  assign n2474 = n2470 & n2471;
  assign n2475 = ~pi64 & ~pi81;
  assign n2476 = ~pi65 & ~pi102;
  assign n2477 = n2475 & n2476;
  assign n2478 = ~pi65 & ~pi71;
  assign n2479 = ~pi102 & n2475;
  assign n2480 = n2478 & n2479;
  assign n2481 = ~pi71 & n2477;
  assign n2482 = ~pi102 & n58783;
  assign n2483 = n2475 & n2482;
  assign n2484 = n2478 & n2483;
  assign n2485 = n58783 & n58784;
  assign n2486 = n2469 & n2478;
  assign n2487 = n2483 & n2486;
  assign n2488 = n2469 & n58785;
  assign n2489 = ~pi53 & ~pi60;
  assign n2490 = ~pi109 & ~pi110;
  assign n2491 = ~pi46 & n2490;
  assign n2492 = ~pi47 & ~pi91;
  assign n2493 = ~pi97 & ~pi108;
  assign n2494 = n2492 & n2493;
  assign n2495 = ~pi46 & ~pi97;
  assign n2496 = ~pi46 & n2493;
  assign n2497 = ~pi108 & n2495;
  assign n2498 = n2490 & n58787;
  assign n2499 = n2492 & n2498;
  assign n2500 = n2491 & n2494;
  assign n2501 = ~pi86 & ~pi94;
  assign n2502 = n58788 & n2501;
  assign n2503 = ~pi86 & n2489;
  assign n2504 = ~pi94 & n2493;
  assign n2505 = ~pi94 & n2498;
  assign n2506 = n2491 & n2504;
  assign n2507 = n2489 & n2501;
  assign n2508 = ~pi46 & n2503;
  assign n2509 = n2504 & n2508;
  assign n2510 = n58787 & n2507;
  assign n2511 = n2490 & n58790;
  assign n2512 = n2503 & n58789;
  assign n2513 = n2492 & n58791;
  assign n2514 = n2489 & n2502;
  assign n2515 = ~pi60 & n58786;
  assign n2516 = ~pi53 & n2502;
  assign n2517 = n2515 & n2516;
  assign n2518 = n58786 & n58792;
  assign n2519 = n2446 & n2486;
  assign n2520 = ~pi64 & n2519;
  assign n2521 = ~pi81 & n2520;
  assign n2522 = n2482 & n2521;
  assign n2523 = n2446 & n58786;
  assign n2524 = n58792 & n58794;
  assign n2525 = n2446 & n58793;
  assign n2526 = n2445 & n58795;
  assign n2527 = ~pi841 & n2526;
  assign n2528 = pi93 & ~n2527;
  assign n2529 = n2444 & ~n2528;
  assign n2530 = ~pi58 & ~pi91;
  assign n2531 = ~pi47 & n2530;
  assign n2532 = n2490 & n2531;
  assign n2533 = ~pi47 & n2490;
  assign n2534 = ~pi47 & n58791;
  assign n2535 = n58790 & n2533;
  assign n2536 = n2530 & n58796;
  assign n2537 = ~pi58 & n58788;
  assign n2538 = n58787 & n2532;
  assign n2539 = ~pi109 & n58787;
  assign n2540 = ~pi47 & ~pi110;
  assign n2541 = ~pi110 & n2531;
  assign n2542 = n2530 & n2540;
  assign n2543 = n2539 & n58799;
  assign n2544 = n2498 & n2531;
  assign n2545 = n2507 & n58798;
  assign n2546 = n58790 & n2532;
  assign n2547 = n2483 & n58797;
  assign n2548 = n58790 & n58794;
  assign n2549 = n2533 & n2548;
  assign n2550 = n58794 & n58796;
  assign n2551 = n2530 & n58800;
  assign n2552 = n2532 & n2548;
  assign n2553 = n2519 & n2547;
  assign n2554 = ~pi841 & n58801;
  assign n2555 = pi90 & n2554;
  assign n2556 = ~pi93 & ~n2555;
  assign n2557 = n2529 & ~n2556;
  assign n2558 = ~pi51 & ~n2557;
  assign n2559 = ~pi102 & n2521;
  assign n2560 = ~pi88 & pi98;
  assign n2561 = n2471 & n2560;
  assign n2562 = ~pi50 & n2489;
  assign n2563 = ~pi77 & n2562;
  assign n2564 = n2471 & n2489;
  assign n2565 = n2501 & n58802;
  assign n2566 = n2560 & n2565;
  assign n2567 = n2507 & n2561;
  assign n2568 = ~pi94 & n2471;
  assign n2569 = n2471 & n2559;
  assign n2570 = ~pi94 & n2569;
  assign n2571 = n2559 & n2568;
  assign n2572 = n2503 & n2560;
  assign n2573 = n58804 & n2572;
  assign n2574 = n2507 & n2560;
  assign n2575 = n2569 & n2574;
  assign n2576 = n2559 & n58803;
  assign n2577 = ~pi90 & n58798;
  assign n2578 = n58805 & n2577;
  assign n2579 = ~pi90 & ~pi93;
  assign n2580 = ~pi35 & n2579;
  assign n2581 = ~pi70 & n2580;
  assign n2582 = ~pi97 & ~n58805;
  assign n2583 = n58798 & ~n2582;
  assign n2584 = n2581 & n2583;
  assign n2585 = n2529 & n2577;
  assign n2586 = n58805 & n2585;
  assign n2587 = n2529 & n2578;
  assign n2588 = n2558 & ~n58806;
  assign n2589 = ~pi93 & n2445;
  assign n2590 = ~pi93 & n2526;
  assign n2591 = n58795 & n2589;
  assign n2592 = ~pi35 & ~pi93;
  assign n2593 = n2526 & n2592;
  assign n2594 = ~pi70 & n2593;
  assign n2595 = n2444 & n58807;
  assign n2596 = pi51 & ~n58808;
  assign n2597 = ~pi40 & ~pi72;
  assign n2598 = ~pi32 & ~pi95;
  assign n2599 = n2597 & n2598;
  assign n2600 = ~pi72 & ~pi96;
  assign n2601 = ~pi40 & n2600;
  assign n2602 = n2598 & n2601;
  assign n2603 = ~pi96 & n2599;
  assign n2604 = ~pi96 & ~n2596;
  assign n2605 = n2599 & n2604;
  assign n2606 = ~n2596 & n58809;
  assign n2607 = ~n2588 & ~n2596;
  assign n2608 = n58809 & n2607;
  assign n2609 = ~n2588 & n58810;
  assign n2610 = n2443 & n58811;
  assign n2611 = ~n2440 & n2610;
  assign n2612 = ~pi96 & ~n2607;
  assign n2613 = n2440 & n2441;
  assign n2614 = ~pi51 & n2444;
  assign n2615 = ~pi841 & n58807;
  assign n2616 = n2614 & n2615;
  assign n2617 = pi96 & ~n2616;
  assign n2618 = n2597 & ~n2617;
  assign n2619 = n2598 & n2618;
  assign n2620 = ~pi32 & ~pi40;
  assign n2621 = ~pi95 & n2620;
  assign n2622 = ~n2617 & n2621;
  assign n2623 = ~pi72 & n2622;
  assign n2624 = n2599 & ~n2617;
  assign n2625 = ~pi72 & n2613;
  assign n2626 = n2622 & n2625;
  assign n2627 = n2613 & n58812;
  assign n2628 = ~n2612 & n2622;
  assign n2629 = n2625 & n2628;
  assign n2630 = ~n2612 & n58813;
  assign n2631 = ~n2611 & ~n58814;
  assign n2632 = ~pi1093 & ~n2631;
  assign n2633 = ~pi87 & ~n2632;
  assign n2634 = ~pi38 & ~pi39;
  assign n2635 = ~pi75 & ~pi100;
  assign n2636 = ~pi38 & ~pi100;
  assign n2637 = ~pi100 & n2634;
  assign n2638 = ~pi39 & n2636;
  assign n2639 = ~pi75 & n58815;
  assign n2640 = n2634 & n2635;
  assign n2641 = ~pi70 & ~pi96;
  assign n2642 = ~pi51 & ~pi72;
  assign n2643 = ~pi51 & ~pi70;
  assign n2644 = n2600 & n2643;
  assign n2645 = n2641 & n2642;
  assign n2646 = ~pi70 & n58809;
  assign n2647 = n2599 & n2641;
  assign n2648 = ~pi51 & n58818;
  assign n2649 = n2601 & n2643;
  assign n2650 = ~pi40 & n58817;
  assign n2651 = n2598 & n58820;
  assign n2652 = n2621 & n58817;
  assign n2653 = ~pi51 & ~pi96;
  assign n2654 = ~pi51 & n58809;
  assign n2655 = n2599 & n2653;
  assign n2656 = n58808 & n58821;
  assign n2657 = n2600 & n2614;
  assign n2658 = ~pi35 & n58817;
  assign n2659 = n2593 & n58817;
  assign n2660 = n58807 & n58823;
  assign n2661 = n2620 & n58824;
  assign n2662 = ~pi95 & n2661;
  assign n2663 = n2593 & n58819;
  assign po740 = ~pi1093 & n2443;
  assign n2665 = n58822 & po740;
  assign n2666 = pi87 & ~n2665;
  assign n2667 = n58816 & ~n2666;
  assign n2668 = ~n2633 & n2667;
  assign n2669 = ~pi567 & ~n2668;
  assign n2670 = n2439 & ~n2669;
  assign n2671 = ~pi39 & ~pi87;
  assign n2672 = n2636 & n2671;
  assign n2673 = ~pi144 & ~pi174;
  assign n2674 = ~pi189 & n2673;
  assign n2675 = ~pi299 & ~n2674;
  assign n2676 = ~pi152 & ~pi161;
  assign n2677 = ~pi166 & n2676;
  assign n2678 = pi299 & ~n2677;
  assign n2679 = ~n2675 & ~n2678;
  assign n2680 = ~pi332 & ~pi468;
  assign n2681 = pi232 & n2680;
  assign n2682 = n2679 & n2681;
  assign n2683 = n2672 & ~n2682;
  assign n2684 = pi252 & n2621;
  assign n2685 = pi252 & n58822;
  assign n2686 = n58824 & n2684;
  assign n2687 = ~pi24 & n2593;
  assign n2688 = n58819 & n2687;
  assign n2689 = ~pi24 & n58822;
  assign n2690 = pi252 & n58826;
  assign n2691 = ~pi24 & n58825;
  assign n2692 = ~pi833 & pi957;
  assign n2693 = ~pi41 & ~pi99;
  assign n2694 = ~pi101 & n2693;
  assign n2695 = ~pi113 & ~pi116;
  assign n2696 = ~pi52 & n2695;
  assign n2697 = ~pi42 & ~pi43;
  assign n2698 = ~pi114 & ~pi115;
  assign n2699 = ~pi114 & n2697;
  assign n2700 = ~pi115 & n2699;
  assign n2701 = n2697 & n2698;
  assign n2702 = ~pi52 & n2697;
  assign n2703 = n2695 & n2698;
  assign n2704 = n2702 & n2703;
  assign n2705 = n2696 & n58828;
  assign n2706 = n2694 & n58829;
  assign n2707 = ~pi44 & n2706;
  assign n2708 = ~n2692 & ~n2707;
  assign n2709 = pi1091 & n2708;
  assign n2710 = n2613 & n2709;
  assign n2711 = n58827 & n2710;
  assign n2712 = pi1093 & n2711;
  assign n2713 = n2683 & n2712;
  assign n2714 = pi75 & ~n2713;
  assign n2715 = pi1093 & n2613;
  assign n2716 = n2708 & n2715;
  assign n2717 = n58822 & n2716;
  assign n2718 = pi1091 & n2717;
  assign n2719 = pi228 & ~n2682;
  assign n2720 = n2634 & n2719;
  assign n2721 = pi228 & n2718;
  assign n2722 = n2634 & ~n2682;
  assign n2723 = n2721 & n2722;
  assign n2724 = n2718 & n2720;
  assign n2725 = pi100 & ~n58830;
  assign n2726 = pi1093 & ~n2692;
  assign n2727 = pi824 & n2441;
  assign n2728 = ~n2558 & n58810;
  assign n2729 = n2727 & n2728;
  assign n2730 = ~pi829 & n2729;
  assign n2731 = pi91 & n58800;
  assign n2732 = ~pi24 & n2731;
  assign n2733 = n2470 & n2559;
  assign n2734 = ~pi77 & n2733;
  assign n2735 = n2472 & n2559;
  assign n2736 = n2501 & n2562;
  assign n2737 = ~pi50 & n2507;
  assign n2738 = n2565 & n2733;
  assign n2739 = n58802 & n2733;
  assign n2740 = n2562 & n58831;
  assign n2741 = n2501 & n58834;
  assign n2742 = n58831 & n58832;
  assign n2743 = ~pi46 & pi97;
  assign n2744 = ~pi108 & n2743;
  assign n2745 = n2533 & n2744;
  assign n2746 = ~pi108 & n58833;
  assign n2747 = n2533 & n2743;
  assign n2748 = n2746 & n2747;
  assign n2749 = n58833 & n2745;
  assign n2750 = ~pi91 & n58835;
  assign n2751 = ~n2732 & ~n2750;
  assign n2752 = n2445 & n2529;
  assign n2753 = ~n2751 & n2752;
  assign n2754 = n2558 & ~n2753;
  assign n2755 = ~n2596 & ~n2754;
  assign n2756 = ~pi96 & ~n2755;
  assign n2757 = pi829 & n2441;
  assign n2758 = ~pi72 & pi950;
  assign n2759 = n2622 & n2758;
  assign n2760 = pi950 & n58812;
  assign n2761 = pi829 & pi1092;
  assign n2762 = n58836 & n2761;
  assign n2763 = n58812 & n2757;
  assign n2764 = ~n2756 & n58837;
  assign n2765 = ~n2730 & ~n2764;
  assign n2766 = ~pi122 & ~n2765;
  assign n2767 = pi122 & n2443;
  assign n2768 = n2728 & n2767;
  assign n2769 = ~n2766 & ~n2768;
  assign n2770 = n2726 & ~n2769;
  assign n2771 = pi1091 & ~n2770;
  assign n2772 = ~n2632 & n2771;
  assign n2773 = ~pi1091 & ~n2632;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = ~pi39 & ~n2774;
  assign n2776 = pi603 & ~pi642;
  assign n2777 = ~pi614 & ~pi616;
  assign n2778 = n2776 & n2777;
  assign n2779 = ~pi662 & pi680;
  assign n2780 = ~pi661 & n2779;
  assign n2781 = ~pi681 & n2780;
  assign n2782 = ~n2778 & ~n2781;
  assign n2783 = ~n2680 & ~n2782;
  assign n2784 = ~pi969 & ~pi971;
  assign n2785 = ~pi974 & ~pi977;
  assign n2786 = n2784 & n2785;
  assign n2787 = ~pi587 & ~pi602;
  assign n2788 = ~pi961 & ~pi967;
  assign n2789 = n2787 & n2788;
  assign n2790 = n2786 & n2789;
  assign n2791 = n2680 & ~n2790;
  assign n2792 = ~n2783 & ~n2791;
  assign n2793 = pi1091 & ~n2692;
  assign n2794 = pi1092 & pi1093;
  assign n2795 = pi829 & pi950;
  assign n2796 = n2794 & n2795;
  assign n2797 = pi1091 & pi1093;
  assign n2798 = ~n2692 & n2797;
  assign n2799 = n2757 & n2798;
  assign n2800 = n2793 & n2796;
  assign n2801 = ~pi287 & n58822;
  assign n2802 = pi835 & pi984;
  assign n2803 = ~pi252 & ~pi1001;
  assign n2804 = ~pi979 & ~n2803;
  assign n2805 = ~n2802 & n2804;
  assign n2806 = pi835 & n2805;
  assign n2807 = n2801 & n2806;
  assign n2808 = n2795 & n2807;
  assign n2809 = pi1092 & n2808;
  assign n2810 = n2757 & n2807;
  assign n2811 = ~n2692 & n2795;
  assign n2812 = ~n2692 & n2808;
  assign n2813 = n2807 & n2811;
  assign n2814 = n2794 & n58840;
  assign n2815 = n2726 & n58839;
  assign n2816 = pi1091 & n58841;
  assign n2817 = n2798 & n58839;
  assign n2818 = n58838 & n2807;
  assign n2819 = n2783 & n58842;
  assign n2820 = n2790 & ~n2819;
  assign n2821 = ~n2680 & ~n2778;
  assign n2822 = ~n2781 & n2821;
  assign n2823 = n58842 & ~n2822;
  assign n2824 = ~n2790 & ~n2823;
  assign n2825 = ~n2820 & ~n2824;
  assign n2826 = ~n2792 & n58842;
  assign n2827 = pi222 & ~pi224;
  assign n2828 = ~pi223 & ~pi299;
  assign n2829 = pi222 & ~pi223;
  assign n2830 = ~pi299 & n2829;
  assign n2831 = pi222 & n2828;
  assign n2832 = ~pi224 & n58844;
  assign n2833 = n2827 & n2828;
  assign n2834 = n58843 & n58845;
  assign n2835 = ~pi960 & ~pi963;
  assign n2836 = ~pi970 & ~pi972;
  assign n2837 = ~pi975 & ~pi978;
  assign n2838 = n2836 & n2837;
  assign n2839 = n2835 & n2838;
  assign n2840 = ~pi907 & ~pi947;
  assign n2841 = ~pi907 & n2839;
  assign n2842 = ~pi947 & n2841;
  assign n2843 = n2839 & n2840;
  assign n2844 = n2680 & ~n58846;
  assign n2845 = ~n2783 & ~n2844;
  assign n2846 = ~n2819 & n58846;
  assign n2847 = ~n2823 & ~n58846;
  assign n2848 = ~n2846 & ~n2847;
  assign n2849 = n58842 & ~n2845;
  assign n2850 = ~pi216 & pi221;
  assign n2851 = ~pi215 & pi299;
  assign n2852 = ~pi215 & pi221;
  assign n2853 = pi299 & n2852;
  assign n2854 = ~pi216 & n2853;
  assign n2855 = n2850 & n2851;
  assign n2856 = n58847 & n58848;
  assign n2857 = pi39 & ~n2856;
  assign n2858 = ~n2834 & n2857;
  assign n2859 = ~pi38 & ~n2858;
  assign n2860 = ~n2775 & n2859;
  assign n2861 = ~pi100 & ~n2860;
  assign n2862 = pi824 & pi1093;
  assign n2863 = pi1093 & n2727;
  assign n2864 = n2441 & n2862;
  assign n2865 = pi1093 & n2729;
  assign n2866 = n2728 & n58849;
  assign n2867 = n2859 & n58850;
  assign n2868 = ~n2771 & n2867;
  assign n2869 = n2861 & ~n2868;
  assign n2870 = ~n2725 & ~n2869;
  assign n2871 = ~pi87 & ~n2870;
  assign n2872 = pi824 & pi950;
  assign n2873 = pi950 & n58822;
  assign n2874 = pi824 & n2873;
  assign n2875 = n58822 & n2872;
  assign n2876 = pi1092 & n58851;
  assign n2877 = n58822 & n2727;
  assign n2878 = ~pi1091 & pi1093;
  assign n2879 = ~n58852 & n2878;
  assign n2880 = pi1093 & n2692;
  assign n2881 = n2443 & ~n2880;
  assign n2882 = n58822 & n2881;
  assign n2883 = ~n2878 & ~n2882;
  assign n2884 = n58815 & ~n2883;
  assign n2885 = ~n2879 & n2884;
  assign n2886 = pi87 & ~n2885;
  assign n2887 = ~n2871 & ~n2886;
  assign n2888 = ~pi75 & ~n2887;
  assign n2889 = ~n2714 & ~n2888;
  assign n2890 = pi567 & ~n2889;
  assign n2891 = n2670 & ~n2890;
  assign n2892 = ~pi452 & ~pi455;
  assign n2893 = pi452 & pi455;
  assign n2894 = pi452 & ~pi455;
  assign n2895 = ~pi452 & pi455;
  assign n2896 = ~n2894 & ~n2895;
  assign n2897 = ~n2892 & ~n2893;
  assign n2898 = n2891 & n58853;
  assign n2899 = ~pi87 & ~n2725;
  assign n2900 = ~n2861 & n2899;
  assign n2901 = ~pi1091 & ~n2665;
  assign n2902 = pi1091 & ~n2882;
  assign n2903 = pi87 & ~pi100;
  assign n2904 = pi87 & n58815;
  assign n2905 = n2634 & n2903;
  assign n2906 = ~n2902 & n58854;
  assign n2907 = ~n2901 & n2906;
  assign n2908 = ~pi75 & ~n2907;
  assign n2909 = ~n2900 & n2908;
  assign n2910 = ~n2714 & ~n2909;
  assign n2911 = pi567 & ~n2910;
  assign n2912 = n2670 & ~n2911;
  assign n2913 = ~pi592 & ~n2912;
  assign n2914 = pi592 & ~n2891;
  assign n2915 = ~n2913 & ~n2914;
  assign n2916 = ~n58853 & n2915;
  assign n2917 = pi455 & ~n2915;
  assign n2918 = ~pi455 & ~n2891;
  assign n2919 = ~n2917 & ~n2918;
  assign n2920 = ~pi452 & ~n2919;
  assign n2921 = ~pi455 & ~n2915;
  assign n2922 = pi455 & ~n2891;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = pi452 & ~n2923;
  assign n2925 = ~n2920 & ~n2924;
  assign n2926 = ~n58853 & ~n2915;
  assign n2927 = ~n2891 & n58853;
  assign n2928 = ~n2926 & ~n2927;
  assign n2929 = ~n2898 & ~n2916;
  assign n2930 = ~pi355 & n58855;
  assign n2931 = n58853 & n2915;
  assign n2932 = n2891 & ~n58853;
  assign n2933 = ~pi455 & n2915;
  assign n2934 = pi455 & n2891;
  assign n2935 = ~pi452 & ~n2934;
  assign n2936 = ~pi452 & ~n2923;
  assign n2937 = ~n2933 & n2935;
  assign n2938 = pi455 & n2915;
  assign n2939 = ~pi455 & n2891;
  assign n2940 = pi452 & ~n2939;
  assign n2941 = pi452 & ~n2919;
  assign n2942 = ~n2938 & n2940;
  assign n2943 = ~n58856 & ~n58857;
  assign n2944 = ~n2931 & ~n2932;
  assign n2945 = pi355 & n58858;
  assign n2946 = pi355 & ~n58858;
  assign n2947 = ~pi355 & ~n58855;
  assign n2948 = ~n2946 & ~n2947;
  assign n2949 = ~n2930 & ~n2945;
  assign n2950 = pi458 & ~n58859;
  assign n2951 = ~pi320 & ~pi460;
  assign n2952 = pi320 & pi460;
  assign n2953 = pi320 & ~pi460;
  assign n2954 = ~pi320 & pi460;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = ~n2951 & ~n2952;
  assign n2957 = pi342 & ~n58860;
  assign n2958 = ~pi342 & n58860;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = pi361 & ~pi441;
  assign n2961 = ~pi361 & pi441;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = n2959 & n2962;
  assign n2964 = ~n2959 & ~n2962;
  assign n2965 = ~n2963 & ~n2964;
  assign n2966 = pi355 & n58855;
  assign n2967 = ~pi355 & n58858;
  assign n2968 = ~pi355 & ~n58858;
  assign n2969 = pi355 & ~n58855;
  assign n2970 = ~n2968 & ~n2969;
  assign n2971 = ~n2966 & ~n2967;
  assign n2972 = ~pi458 & ~n58861;
  assign n2973 = ~n2965 & ~n2972;
  assign n2974 = ~n2950 & ~n2965;
  assign n2975 = ~n2972 & n2974;
  assign n2976 = ~n2950 & n2973;
  assign n2977 = pi458 & ~n58861;
  assign n2978 = ~pi458 & ~n58859;
  assign n2979 = n2965 & ~n2978;
  assign n2980 = n2965 & ~n2977;
  assign n2981 = ~n2978 & n2980;
  assign n2982 = ~n2977 & n2979;
  assign n2983 = pi1196 & ~n58863;
  assign n2984 = ~n58862 & n2983;
  assign n2985 = ~pi1196 & ~n2891;
  assign n2986 = ~pi1198 & ~n2985;
  assign n2987 = ~n2984 & n2986;
  assign n2988 = ~pi345 & ~pi346;
  assign n2989 = pi345 & pi346;
  assign n2990 = pi345 & ~pi346;
  assign n2991 = ~pi345 & pi346;
  assign n2992 = ~n2990 & ~n2991;
  assign n2993 = ~n2988 & ~n2989;
  assign n2994 = pi450 & ~n58864;
  assign n2995 = ~pi450 & n58864;
  assign n2996 = ~n2994 & ~n2995;
  assign n2997 = pi323 & ~pi358;
  assign n2998 = ~pi323 & pi358;
  assign n2999 = ~n2997 & ~n2998;
  assign n3000 = n2996 & n2999;
  assign n3001 = ~n2996 & ~n2999;
  assign n3002 = pi323 & ~n58864;
  assign n3003 = ~pi323 & n58864;
  assign n3004 = ~n3002 & ~n3003;
  assign n3005 = pi358 & ~pi450;
  assign n3006 = ~pi358 & pi450;
  assign n3007 = ~n3005 & ~n3006;
  assign n3008 = n3004 & ~n3007;
  assign n3009 = ~n3004 & n3007;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = pi358 & ~n3004;
  assign n3012 = ~pi358 & n3004;
  assign n3013 = ~n3011 & ~n3012;
  assign n3014 = pi450 & n3013;
  assign n3015 = ~pi450 & ~n3013;
  assign n3016 = ~n3014 & ~n3015;
  assign n3017 = ~n3000 & ~n3001;
  assign n3018 = pi327 & ~pi362;
  assign n3019 = ~pi327 & pi362;
  assign n3020 = ~pi327 & ~pi362;
  assign n3021 = pi327 & pi362;
  assign n3022 = ~n3020 & ~n3021;
  assign n3023 = ~n3018 & ~n3019;
  assign n3024 = pi343 & ~pi344;
  assign n3025 = ~pi343 & pi344;
  assign n3026 = ~n3024 & ~n3025;
  assign n3027 = ~n58866 & n3026;
  assign n3028 = n58866 & ~n3026;
  assign n3029 = pi343 & ~n58866;
  assign n3030 = ~pi343 & n58866;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = pi344 & n3031;
  assign n3033 = ~pi344 & ~n3031;
  assign n3034 = ~n3032 & ~n3033;
  assign n3035 = ~n3027 & ~n3028;
  assign n3036 = ~n58865 & n58867;
  assign n3037 = n58865 & ~n58867;
  assign n3038 = pi1197 & ~n3037;
  assign n3039 = ~n3036 & n3038;
  assign n3040 = ~pi350 & ~pi592;
  assign n3041 = ~n2891 & ~n3040;
  assign n3042 = pi315 & ~pi359;
  assign n3043 = ~pi315 & pi359;
  assign n3044 = ~n3042 & ~n3043;
  assign n3045 = ~pi321 & ~pi347;
  assign n3046 = pi321 & pi347;
  assign n3047 = pi321 & ~pi347;
  assign n3048 = ~pi321 & pi347;
  assign n3049 = ~n3047 & ~n3048;
  assign n3050 = ~n3045 & ~n3046;
  assign n3051 = pi348 & ~n58868;
  assign n3052 = ~pi348 & n58868;
  assign n3053 = ~n3051 & ~n3052;
  assign n3054 = ~pi316 & ~pi349;
  assign n3055 = pi316 & pi349;
  assign n3056 = pi316 & ~pi349;
  assign n3057 = ~pi316 & pi349;
  assign n3058 = ~n3056 & ~n3057;
  assign n3059 = ~n3054 & ~n3055;
  assign n3060 = pi322 & ~n58869;
  assign n3061 = ~pi322 & n58869;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = n3053 & ~n3062;
  assign n3064 = ~n3053 & n3062;
  assign n3065 = pi322 & ~pi348;
  assign n3066 = ~pi322 & pi348;
  assign n3067 = ~n3065 & ~n3066;
  assign n3068 = n58869 & n3067;
  assign n3069 = ~n58869 & ~n3067;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = n58868 & ~n3070;
  assign n3072 = ~n58868 & n3070;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = ~n3063 & ~n3064;
  assign n3075 = n3044 & ~n58870;
  assign n3076 = ~n3044 & n58870;
  assign n3077 = pi348 & n58869;
  assign n3078 = ~pi348 & ~n58869;
  assign n3079 = ~n3077 & ~n3078;
  assign n3080 = pi322 & n3044;
  assign n3081 = ~pi322 & ~n3044;
  assign n3082 = ~n3080 & ~n3081;
  assign n3083 = n3079 & ~n3082;
  assign n3084 = ~n3079 & n3082;
  assign n3085 = ~n3083 & ~n3084;
  assign n3086 = n58868 & n3085;
  assign n3087 = ~n58868 & ~n3085;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = n3044 & n58870;
  assign n3090 = ~n3044 & ~n58870;
  assign n3091 = ~n3089 & ~n3090;
  assign n3092 = ~n3075 & ~n3076;
  assign n3093 = ~n2912 & n3040;
  assign n3094 = n58871 & ~n3093;
  assign n3095 = ~n3041 & n3094;
  assign n3096 = pi355 & ~pi458;
  assign n3097 = ~pi355 & pi458;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = n2965 & n3098;
  assign n3100 = ~n2965 & ~n3098;
  assign n3101 = pi458 & n2965;
  assign n3102 = ~pi458 & ~n2965;
  assign n3103 = ~n3101 & ~n3102;
  assign n3104 = pi355 & ~n3103;
  assign n3105 = ~pi355 & n3103;
  assign n3106 = ~n3104 & ~n3105;
  assign n3107 = pi355 & ~n2965;
  assign n3108 = ~pi355 & n2965;
  assign n3109 = ~n3107 & ~n3108;
  assign n3110 = pi458 & n3109;
  assign n3111 = ~pi458 & ~n3109;
  assign n3112 = ~n3110 & ~n3111;
  assign n3113 = ~n3099 & ~n3100;
  assign n3114 = ~n58853 & n58872;
  assign n3115 = n58853 & ~n58872;
  assign n3116 = pi355 & n58853;
  assign n3117 = ~pi355 & ~n58853;
  assign n3118 = ~n3116 & ~n3117;
  assign n3119 = n3103 & n3118;
  assign n3120 = ~n3103 & ~n3118;
  assign n3121 = ~n3119 & ~n3120;
  assign n3122 = n58853 & n58872;
  assign n3123 = ~n58853 & ~n58872;
  assign n3124 = ~n3122 & ~n3123;
  assign n3125 = ~n3114 & ~n3115;
  assign n3126 = pi1196 & n58873;
  assign n3127 = pi350 & ~pi592;
  assign n3128 = ~n2891 & ~n3127;
  assign n3129 = ~n2912 & n3127;
  assign n3130 = ~n58871 & ~n3129;
  assign n3131 = ~n3128 & n3130;
  assign n3132 = ~n3126 & ~n3131;
  assign n3133 = ~n3095 & ~n3126;
  assign n3134 = ~n3131 & n3133;
  assign n3135 = ~n3095 & n3132;
  assign n3136 = ~n2915 & n3126;
  assign n3137 = pi1198 & ~n3136;
  assign n3138 = ~n58874 & n3137;
  assign n3139 = ~n3039 & ~n3138;
  assign n3140 = ~n2987 & n3139;
  assign n3141 = ~n2915 & n3039;
  assign n3142 = ~n2987 & ~n3138;
  assign n3143 = ~n3039 & ~n3142;
  assign n3144 = n2915 & n3039;
  assign n3145 = ~n3143 & ~n3144;
  assign n3146 = ~n3140 & ~n3141;
  assign n3147 = ~n2437 & n58875;
  assign n3148 = pi1199 & ~n2915;
  assign n3149 = pi351 & n3148;
  assign n3150 = ~n3147 & ~n3149;
  assign n3151 = ~pi461 & ~n3150;
  assign n3152 = ~pi351 & pi1199;
  assign n3153 = n58875 & ~n3152;
  assign n3154 = ~pi351 & n3148;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = pi461 & ~n3155;
  assign n3157 = ~n3151 & ~n3156;
  assign n3158 = ~pi357 & ~n3157;
  assign n3159 = ~pi461 & ~n3155;
  assign n3160 = pi461 & ~n3150;
  assign n3161 = ~n3159 & ~n3160;
  assign n3162 = pi357 & ~n3161;
  assign n3163 = ~n3158 & ~n3162;
  assign n3164 = pi356 & n3163;
  assign n3165 = ~pi360 & ~pi462;
  assign n3166 = pi360 & pi462;
  assign n3167 = pi360 & ~pi462;
  assign n3168 = ~pi360 & pi462;
  assign n3169 = ~n3167 & ~n3168;
  assign n3170 = ~n3165 & ~n3166;
  assign n3171 = pi352 & ~pi353;
  assign n3172 = ~pi352 & pi353;
  assign n3173 = ~n3171 & ~n3172;
  assign n3174 = ~n58876 & n3173;
  assign n3175 = n58876 & ~n3173;
  assign n3176 = n58876 & n3173;
  assign n3177 = ~n58876 & ~n3173;
  assign n3178 = ~n3176 & ~n3177;
  assign n3179 = ~n3174 & ~n3175;
  assign n3180 = pi354 & ~n58877;
  assign n3181 = ~pi354 & n58877;
  assign n3182 = pi354 & n58877;
  assign n3183 = ~pi354 & ~n58877;
  assign n3184 = ~n3182 & ~n3183;
  assign n3185 = ~n3180 & ~n3181;
  assign n3186 = ~pi357 & ~n3161;
  assign n3187 = pi357 & ~n3157;
  assign n3188 = ~n3186 & ~n3187;
  assign n3189 = ~pi356 & n3188;
  assign n3190 = n58878 & ~n3189;
  assign n3191 = ~pi356 & ~n3188;
  assign n3192 = pi356 & ~n3163;
  assign n3193 = ~n3191 & ~n3192;
  assign n3194 = n58878 & ~n3193;
  assign n3195 = ~n3164 & n3190;
  assign n3196 = pi356 & n3188;
  assign n3197 = ~pi356 & n3163;
  assign n3198 = ~n58878 & ~n3197;
  assign n3199 = ~pi356 & ~n3163;
  assign n3200 = pi356 & ~n3188;
  assign n3201 = ~n3199 & ~n3200;
  assign n3202 = ~n58878 & ~n3201;
  assign n3203 = ~n3196 & n3198;
  assign n3204 = ~pi591 & ~n58880;
  assign n3205 = ~pi591 & ~n58879;
  assign n3206 = ~n58880 & n3205;
  assign n3207 = ~n58879 & n3204;
  assign n3208 = pi591 & n2891;
  assign n3209 = pi590 & ~n3208;
  assign n3210 = ~n58881 & n3209;
  assign n3211 = ~pi285 & ~pi286;
  assign n3212 = ~pi289 & n3211;
  assign n3213 = ~pi288 & n3212;
  assign n3214 = pi333 & pi1197;
  assign n3215 = ~pi75 & ~pi592;
  assign n3216 = ~n2889 & ~n3215;
  assign n3217 = ~pi1196 & ~n2888;
  assign n3218 = ~pi319 & ~pi324;
  assign n3219 = pi319 & pi324;
  assign n3220 = pi319 & ~pi324;
  assign n3221 = ~pi319 & pi324;
  assign n3222 = ~n3220 & ~n3221;
  assign n3223 = ~n3218 & ~n3219;
  assign n3224 = pi456 & ~n58882;
  assign n3225 = ~pi456 & n58882;
  assign n3226 = ~n3224 & ~n3225;
  assign n3227 = pi412 & ~n3226;
  assign n3228 = ~pi412 & n3226;
  assign n3229 = ~n3227 & ~n3228;
  assign n3230 = ~pi397 & ~pi404;
  assign n3231 = pi397 & pi404;
  assign n3232 = pi397 & ~pi404;
  assign n3233 = ~pi397 & pi404;
  assign n3234 = ~n3232 & ~n3233;
  assign n3235 = ~n3230 & ~n3231;
  assign n3236 = ~pi390 & ~pi410;
  assign n3237 = pi390 & pi410;
  assign n3238 = pi390 & ~pi410;
  assign n3239 = ~pi390 & pi410;
  assign n3240 = ~n3238 & ~n3239;
  assign n3241 = ~n3236 & ~n3237;
  assign n3242 = pi411 & ~n58884;
  assign n3243 = ~pi411 & n58884;
  assign n3244 = ~n3242 & ~n3243;
  assign n3245 = ~n58883 & ~n3244;
  assign n3246 = n58883 & n3244;
  assign n3247 = pi411 & ~n58883;
  assign n3248 = ~pi411 & n58883;
  assign n3249 = ~n3247 & ~n3248;
  assign n3250 = ~n58884 & n3249;
  assign n3251 = n58884 & ~n3249;
  assign n3252 = ~n3250 & ~n3251;
  assign n3253 = n58884 & n3249;
  assign n3254 = ~n58884 & ~n3249;
  assign n3255 = ~n3253 & ~n3254;
  assign n3256 = ~n3245 & ~n3246;
  assign n3257 = n3229 & ~n58885;
  assign n3258 = ~n3229 & n58885;
  assign n3259 = pi412 & ~n58883;
  assign n3260 = ~pi412 & n58883;
  assign n3261 = pi397 & ~pi412;
  assign n3262 = ~pi397 & pi412;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = pi404 & n3263;
  assign n3265 = ~pi404 & ~n3263;
  assign n3266 = ~n3264 & ~n3265;
  assign n3267 = ~n3259 & ~n3260;
  assign n3268 = ~n58884 & ~n58886;
  assign n3269 = n58884 & n58886;
  assign n3270 = ~n3268 & ~n3269;
  assign n3271 = n3226 & n3270;
  assign n3272 = ~n3226 & ~n3270;
  assign n3273 = ~n3226 & n58886;
  assign n3274 = n3226 & ~n58886;
  assign n3275 = ~n3273 & ~n3274;
  assign n3276 = n58884 & n3275;
  assign n3277 = ~n58884 & ~n3275;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = ~n3271 & ~n3272;
  assign n3280 = pi411 & n58887;
  assign n3281 = ~pi411 & ~n58887;
  assign n3282 = ~n3280 & ~n3281;
  assign n3283 = ~n3257 & ~n3258;
  assign n3284 = n2868 & n58888;
  assign n3285 = n2861 & ~n3284;
  assign n3286 = n2899 & ~n3285;
  assign n3287 = n58852 & n58888;
  assign n3288 = n2878 & ~n3287;
  assign n3289 = pi87 & n2884;
  assign n3290 = ~n2883 & n58854;
  assign n3291 = ~n3288 & n58889;
  assign n3292 = n3215 & ~n3291;
  assign n3293 = ~n3286 & n3292;
  assign n3294 = pi1196 & ~n3293;
  assign n3295 = ~pi1199 & ~n3294;
  assign n3296 = pi1196 & n3215;
  assign n3297 = ~n3291 & n3296;
  assign n3298 = ~n3286 & n3297;
  assign n3299 = ~pi1196 & n2888;
  assign n3300 = ~n3298 & ~n3299;
  assign n3301 = ~pi1199 & ~n3300;
  assign n3302 = ~n3217 & n3295;
  assign n3303 = ~pi318 & ~pi409;
  assign n3304 = pi318 & pi409;
  assign n3305 = pi318 & ~pi409;
  assign n3306 = ~pi318 & pi409;
  assign n3307 = ~n3305 & ~n3306;
  assign n3308 = ~n3303 & ~n3304;
  assign n3309 = pi325 & ~n58891;
  assign n3310 = ~pi325 & n58891;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = pi326 & ~n3311;
  assign n3313 = ~pi326 & n3311;
  assign n3314 = ~n3312 & ~n3313;
  assign n3315 = pi403 & ~pi405;
  assign n3316 = ~pi403 & pi405;
  assign n3317 = ~pi403 & ~pi405;
  assign n3318 = pi403 & pi405;
  assign n3319 = ~n3317 & ~n3318;
  assign n3320 = ~n3315 & ~n3316;
  assign n3321 = pi406 & ~n58892;
  assign n3322 = ~pi406 & n58892;
  assign n3323 = ~n3321 & ~n3322;
  assign n3324 = ~pi401 & ~pi402;
  assign n3325 = pi401 & pi402;
  assign n3326 = pi401 & ~pi402;
  assign n3327 = ~pi401 & pi402;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = ~n3324 & ~n3325;
  assign n3330 = n3323 & n58893;
  assign n3331 = ~n3323 & ~n58893;
  assign n3332 = ~n3330 & ~n3331;
  assign n3333 = n3314 & n3332;
  assign n3334 = ~n3314 & ~n3332;
  assign n3335 = pi406 & n58893;
  assign n3336 = ~pi406 & ~n58893;
  assign n3337 = ~n3335 & ~n3336;
  assign n3338 = pi325 & ~pi326;
  assign n3339 = ~pi325 & pi326;
  assign n3340 = ~n3338 & ~n3339;
  assign n3341 = n58892 & n3340;
  assign n3342 = ~n58892 & ~n3340;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = n3337 & ~n3343;
  assign n3345 = ~n3337 & n3343;
  assign n3346 = ~n3344 & ~n3345;
  assign n3347 = n58891 & n3346;
  assign n3348 = ~n58891 & ~n3346;
  assign n3349 = ~n3347 & ~n3348;
  assign n3350 = pi326 & ~pi406;
  assign n3351 = ~pi326 & pi406;
  assign n3352 = ~n3350 & ~n3351;
  assign n3353 = n58893 & n3352;
  assign n3354 = ~n58893 & ~n3352;
  assign n3355 = ~n3353 & ~n3354;
  assign n3356 = n58892 & ~n3355;
  assign n3357 = ~n58892 & n3355;
  assign n3358 = ~n3356 & ~n3357;
  assign n3359 = n3311 & n3358;
  assign n3360 = ~n3311 & ~n3358;
  assign n3361 = ~n3359 & ~n3360;
  assign n3362 = ~n3333 & ~n3334;
  assign n3363 = pi1196 & ~n58888;
  assign n3364 = ~pi75 & n3363;
  assign n3365 = ~n58894 & ~n3364;
  assign n3366 = n2868 & n3365;
  assign n3367 = n2861 & ~n3366;
  assign n3368 = n2899 & ~n3367;
  assign n3369 = ~n58894 & ~n3363;
  assign n3370 = n58852 & n3369;
  assign n3371 = n2878 & ~n3370;
  assign n3372 = pi1196 & n3288;
  assign n3373 = n58852 & ~n58894;
  assign n3374 = n2878 & ~n3373;
  assign n3375 = n58889 & ~n3374;
  assign n3376 = ~n3372 & n3375;
  assign n3377 = n58889 & ~n3371;
  assign n3378 = pi1199 & n3215;
  assign n3379 = ~n3288 & n3375;
  assign n3380 = ~pi1196 & n3375;
  assign n3381 = n3378 & ~n3380;
  assign n3382 = ~n3379 & n3381;
  assign n3383 = ~n58895 & n3378;
  assign n3384 = ~n3368 & n58896;
  assign n3385 = ~n58890 & ~n3384;
  assign n3386 = ~n3216 & ~n3384;
  assign n3387 = ~n58890 & n3386;
  assign n3388 = ~n3216 & n3385;
  assign n3389 = pi567 & ~n58897;
  assign n3390 = pi328 & ~pi408;
  assign n3391 = ~pi328 & pi408;
  assign n3392 = ~n3390 & ~n3391;
  assign n3393 = ~pi329 & ~pi395;
  assign n3394 = pi329 & pi395;
  assign n3395 = pi329 & ~pi395;
  assign n3396 = ~pi329 & pi395;
  assign n3397 = ~n3395 & ~n3396;
  assign n3398 = ~n3393 & ~n3394;
  assign n3399 = pi396 & ~n58898;
  assign n3400 = ~pi396 & n58898;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = ~pi398 & ~pi399;
  assign n3403 = pi398 & pi399;
  assign n3404 = pi398 & ~pi399;
  assign n3405 = ~pi398 & pi399;
  assign n3406 = ~n3404 & ~n3405;
  assign n3407 = ~n3402 & ~n3403;
  assign n3408 = pi394 & ~pi400;
  assign n3409 = ~pi394 & pi400;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = ~n58899 & n3410;
  assign n3412 = n58899 & ~n3410;
  assign n3413 = ~n3411 & ~n3412;
  assign n3414 = n3401 & ~n3413;
  assign n3415 = ~n3401 & n3413;
  assign n3416 = ~n3414 & ~n3415;
  assign n3417 = n3392 & n3416;
  assign n3418 = ~n3392 & ~n3416;
  assign n3419 = ~pi394 & ~pi396;
  assign n3420 = pi394 & pi396;
  assign n3421 = ~n3419 & ~n3420;
  assign n3422 = n3392 & ~n3421;
  assign n3423 = ~n3392 & n3421;
  assign n3424 = ~n3422 & ~n3423;
  assign n3425 = pi395 & n58899;
  assign n3426 = ~pi395 & ~n58899;
  assign n3427 = ~n3425 & ~n3426;
  assign n3428 = pi329 & ~n3427;
  assign n3429 = ~pi329 & n3427;
  assign n3430 = ~n3428 & ~n3429;
  assign n3431 = pi400 & ~n3430;
  assign n3432 = ~pi400 & n3430;
  assign n3433 = ~n3431 & ~n3432;
  assign n3434 = n3424 & n3433;
  assign n3435 = ~n3424 & ~n3433;
  assign n3436 = ~n3434 & ~n3435;
  assign n3437 = pi400 & ~n58899;
  assign n3438 = ~pi400 & n58899;
  assign n3439 = ~n3437 & ~n3438;
  assign n3440 = pi394 & ~n3392;
  assign n3441 = ~pi394 & n3392;
  assign n3442 = ~n3440 & ~n3441;
  assign n3443 = n3439 & ~n3442;
  assign n3444 = ~n3439 & n3442;
  assign n3445 = ~n3443 & ~n3444;
  assign n3446 = n3401 & n3445;
  assign n3447 = ~n3401 & ~n3445;
  assign n3448 = ~n3446 & ~n3447;
  assign n3449 = ~n3417 & ~n3418;
  assign n3450 = pi1198 & ~n58900;
  assign n3451 = n2670 & ~n3450;
  assign n3452 = ~n3389 & n3451;
  assign n3453 = n2915 & n3450;
  assign n3454 = ~n3452 & ~n3453;
  assign n3455 = ~n3214 & n3454;
  assign n3456 = pi1197 & ~n2915;
  assign n3457 = pi333 & n3456;
  assign n3458 = ~pi1197 & n3454;
  assign n3459 = ~n3456 & ~n3458;
  assign n3460 = pi333 & ~n3459;
  assign n3461 = ~pi333 & n3454;
  assign n3462 = ~n3460 & ~n3461;
  assign n3463 = ~n3455 & ~n3457;
  assign n3464 = ~pi391 & ~n58901;
  assign n3465 = ~pi333 & pi1197;
  assign n3466 = n3454 & ~n3465;
  assign n3467 = ~pi333 & n3456;
  assign n3468 = pi333 & ~n3454;
  assign n3469 = ~pi333 & n3459;
  assign n3470 = ~n3468 & ~n3469;
  assign n3471 = ~pi333 & ~n3459;
  assign n3472 = pi333 & n3454;
  assign n3473 = ~n3471 & ~n3472;
  assign n3474 = ~n3466 & ~n3467;
  assign n3475 = pi391 & n58902;
  assign n3476 = ~n3464 & ~n3475;
  assign n3477 = ~pi392 & ~n3476;
  assign n3478 = pi391 & ~n58901;
  assign n3479 = ~pi391 & n58902;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = pi392 & ~n3480;
  assign n3482 = ~n3477 & ~n3481;
  assign n3483 = pi393 & ~n3482;
  assign n3484 = ~pi407 & ~pi463;
  assign n3485 = pi407 & pi463;
  assign n3486 = pi407 & ~pi463;
  assign n3487 = ~pi407 & pi463;
  assign n3488 = ~n3486 & ~n3487;
  assign n3489 = ~n3484 & ~n3485;
  assign n3490 = pi335 & ~pi413;
  assign n3491 = ~pi335 & pi413;
  assign n3492 = ~n3490 & ~n3491;
  assign n3493 = ~n58903 & n3492;
  assign n3494 = n58903 & ~n3492;
  assign n3495 = n58903 & n3492;
  assign n3496 = ~n58903 & ~n3492;
  assign n3497 = ~n3495 & ~n3496;
  assign n3498 = ~n3493 & ~n3494;
  assign n3499 = pi334 & n58904;
  assign n3500 = ~pi334 & ~n58904;
  assign n3501 = pi334 & ~n58904;
  assign n3502 = ~pi334 & n58904;
  assign n3503 = ~n3501 & ~n3502;
  assign n3504 = ~n3499 & ~n3500;
  assign n3505 = ~pi392 & ~n3480;
  assign n3506 = pi392 & ~n3476;
  assign n3507 = ~n3505 & ~n3506;
  assign n3508 = ~pi393 & ~n3507;
  assign n3509 = ~n58905 & ~n3508;
  assign n3510 = ~n3483 & n3509;
  assign n3511 = pi393 & ~n3507;
  assign n3512 = ~pi393 & ~n3482;
  assign n3513 = n58905 & ~n3512;
  assign n3514 = ~n3511 & n3513;
  assign n3515 = pi591 & ~n3514;
  assign n3516 = ~n3510 & n3515;
  assign n3517 = ~pi370 & ~pi371;
  assign n3518 = pi370 & pi371;
  assign n3519 = pi370 & ~pi371;
  assign n3520 = ~pi370 & pi371;
  assign n3521 = ~n3519 & ~n3520;
  assign n3522 = ~n3517 & ~n3518;
  assign n3523 = ~pi338 & ~pi388;
  assign n3524 = pi338 & pi388;
  assign n3525 = pi338 & ~pi388;
  assign n3526 = ~pi338 & pi388;
  assign n3527 = ~n3525 & ~n3526;
  assign n3528 = ~n3523 & ~n3524;
  assign n3529 = pi337 & ~n58907;
  assign n3530 = ~pi337 & n58907;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = pi339 & ~pi386;
  assign n3533 = ~pi339 & pi386;
  assign n3534 = ~n3532 & ~n3533;
  assign n3535 = pi363 & ~pi372;
  assign n3536 = ~pi363 & pi372;
  assign n3537 = ~pi363 & ~pi372;
  assign n3538 = pi363 & pi372;
  assign n3539 = ~n3537 & ~n3538;
  assign n3540 = ~n3535 & ~n3536;
  assign n3541 = ~pi380 & ~pi387;
  assign n3542 = pi380 & pi387;
  assign n3543 = pi380 & ~pi387;
  assign n3544 = ~pi380 & pi387;
  assign n3545 = ~n3543 & ~n3544;
  assign n3546 = ~n3541 & ~n3542;
  assign n3547 = ~n58908 & n58909;
  assign n3548 = n58908 & ~n58909;
  assign n3549 = ~n3547 & ~n3548;
  assign n3550 = n3534 & n3549;
  assign n3551 = ~n3534 & ~n3549;
  assign n3552 = ~n3550 & ~n3551;
  assign n3553 = n3531 & ~n3552;
  assign n3554 = ~n3531 & n3552;
  assign n3555 = pi1196 & ~n3554;
  assign n3556 = pi386 & ~n58908;
  assign n3557 = ~pi386 & n58908;
  assign n3558 = ~n3556 & ~n3557;
  assign n3559 = pi337 & ~pi339;
  assign n3560 = ~pi337 & pi339;
  assign n3561 = ~n3559 & ~n3560;
  assign n3562 = n58907 & n3561;
  assign n3563 = ~n58907 & ~n3561;
  assign n3564 = ~n3562 & ~n3563;
  assign n3565 = n3558 & ~n3564;
  assign n3566 = ~n3558 & n3564;
  assign n3567 = ~n3565 & ~n3566;
  assign n3568 = n58909 & n3567;
  assign n3569 = ~n58909 & ~n3567;
  assign n3570 = pi387 & n3561;
  assign n3571 = ~pi387 & ~n3561;
  assign n3572 = ~n3570 & ~n3571;
  assign n3573 = pi380 & ~n3572;
  assign n3574 = ~pi380 & n3572;
  assign n3575 = ~n3573 & ~n3574;
  assign n3576 = n58907 & ~n3575;
  assign n3577 = ~n58907 & n3575;
  assign n3578 = ~n3576 & ~n3577;
  assign n3579 = n3558 & n3578;
  assign n3580 = ~n3558 & ~n3578;
  assign n3581 = ~n3579 & ~n3580;
  assign n3582 = ~n3568 & ~n3569;
  assign n3583 = pi1196 & ~n58910;
  assign n3584 = ~n3553 & n3555;
  assign n3585 = pi368 & ~pi389;
  assign n3586 = ~pi368 & pi389;
  assign n3587 = ~pi368 & ~pi389;
  assign n3588 = pi368 & pi389;
  assign n3589 = ~n3587 & ~n3588;
  assign n3590 = ~n3585 & ~n3586;
  assign n3591 = ~pi365 & ~pi447;
  assign n3592 = pi365 & pi447;
  assign n3593 = pi365 & ~pi447;
  assign n3594 = ~pi365 & pi447;
  assign n3595 = ~n3593 & ~n3594;
  assign n3596 = ~n3591 & ~n3592;
  assign n3597 = pi367 & n58913;
  assign n3598 = ~pi367 & ~n58913;
  assign n3599 = pi367 & ~n58913;
  assign n3600 = ~pi367 & n58913;
  assign n3601 = ~n3599 & ~n3600;
  assign n3602 = ~n3597 & ~n3598;
  assign n3603 = ~pi336 & ~pi383;
  assign n3604 = pi336 & pi383;
  assign n3605 = pi336 & ~pi383;
  assign n3606 = ~pi336 & pi383;
  assign n3607 = ~n3605 & ~n3606;
  assign n3608 = ~n3603 & ~n3604;
  assign n3609 = pi364 & ~pi366;
  assign n3610 = ~pi364 & pi366;
  assign n3611 = ~n3609 & ~n3610;
  assign n3612 = ~n58915 & n3611;
  assign n3613 = n58915 & ~n3611;
  assign n3614 = n58915 & n3611;
  assign n3615 = ~n58915 & ~n3611;
  assign n3616 = ~n3614 & ~n3615;
  assign n3617 = ~n3612 & ~n3613;
  assign n3618 = ~n58914 & ~n58916;
  assign n3619 = n58914 & n58916;
  assign n3620 = n58913 & n58916;
  assign n3621 = ~n58913 & ~n58916;
  assign n3622 = ~n3620 & ~n3621;
  assign n3623 = pi367 & ~n3622;
  assign n3624 = ~pi367 & n3622;
  assign n3625 = ~n3623 & ~n3624;
  assign n3626 = ~n3618 & ~n3619;
  assign n3627 = ~n58912 & ~n58917;
  assign n3628 = n58912 & n58917;
  assign n3629 = pi1197 & ~n3628;
  assign n3630 = ~n58912 & n58914;
  assign n3631 = n58912 & ~n58914;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = n58916 & n3632;
  assign n3634 = ~n58916 & ~n3632;
  assign n3635 = n58912 & n3622;
  assign n3636 = ~n58912 & ~n3622;
  assign n3637 = ~n3635 & ~n3636;
  assign n3638 = pi367 & ~n3637;
  assign n3639 = ~pi367 & n3637;
  assign n3640 = ~n3638 & ~n3639;
  assign n3641 = ~n3633 & ~n3634;
  assign n3642 = pi1197 & n58918;
  assign n3643 = ~n3627 & n3629;
  assign n3644 = ~n58911 & ~n58919;
  assign n3645 = pi317 & ~pi385;
  assign n3646 = ~pi317 & pi385;
  assign n3647 = ~n3645 & ~n3646;
  assign n3648 = ~pi379 & ~pi382;
  assign n3649 = pi379 & pi382;
  assign n3650 = pi379 & ~pi382;
  assign n3651 = ~pi379 & pi382;
  assign n3652 = ~n3650 & ~n3651;
  assign n3653 = ~n3648 & ~n3649;
  assign n3654 = pi381 & ~n58920;
  assign n3655 = ~pi381 & n58920;
  assign n3656 = ~n3654 & ~n3655;
  assign n3657 = ~pi376 & ~pi439;
  assign n3658 = pi376 & pi439;
  assign n3659 = pi376 & ~pi439;
  assign n3660 = ~pi376 & pi439;
  assign n3661 = ~n3659 & ~n3660;
  assign n3662 = ~n3657 & ~n3658;
  assign n3663 = pi378 & ~n58921;
  assign n3664 = ~pi378 & n58921;
  assign n3665 = ~n3663 & ~n3664;
  assign n3666 = n3656 & ~n3665;
  assign n3667 = ~n3656 & n3665;
  assign n3668 = pi378 & ~pi381;
  assign n3669 = ~pi378 & pi381;
  assign n3670 = ~n3668 & ~n3669;
  assign n3671 = n58921 & n3670;
  assign n3672 = ~n58921 & ~n3670;
  assign n3673 = ~n3671 & ~n3672;
  assign n3674 = n58920 & ~n3673;
  assign n3675 = ~n58920 & n3673;
  assign n3676 = ~n3674 & ~n3675;
  assign n3677 = ~n3666 & ~n3667;
  assign n3678 = n3647 & ~n58922;
  assign n3679 = ~n3647 & n58922;
  assign n3680 = pi381 & n58921;
  assign n3681 = ~pi381 & ~n58921;
  assign n3682 = ~n3680 & ~n3681;
  assign n3683 = pi378 & n3647;
  assign n3684 = ~pi378 & ~n3647;
  assign n3685 = ~n3683 & ~n3684;
  assign n3686 = n3682 & ~n3685;
  assign n3687 = ~n3682 & n3685;
  assign n3688 = ~n3686 & ~n3687;
  assign n3689 = n58920 & n3688;
  assign n3690 = ~n58920 & ~n3688;
  assign n3691 = ~n3689 & ~n3690;
  assign n3692 = n3647 & n58922;
  assign n3693 = ~n3647 & ~n58922;
  assign n3694 = ~n3692 & ~n3693;
  assign n3695 = ~n3678 & ~n3679;
  assign n3696 = ~pi377 & ~n58923;
  assign n3697 = pi377 & n58923;
  assign n3698 = pi377 & ~n58923;
  assign n3699 = ~pi377 & n58923;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = ~n3696 & ~n3697;
  assign n3702 = pi1199 & ~n58924;
  assign n3703 = n3644 & ~n3702;
  assign n3704 = pi592 & ~n3703;
  assign n3705 = ~n2912 & n3704;
  assign n3706 = ~n2891 & ~n3704;
  assign n3707 = pi377 & pi592;
  assign n3708 = ~n2912 & n3707;
  assign n3709 = ~n58923 & ~n3708;
  assign n3710 = ~n2891 & ~n3707;
  assign n3711 = n3709 & ~n3710;
  assign n3712 = ~pi377 & pi592;
  assign n3713 = ~n2912 & n3712;
  assign n3714 = n58923 & ~n3713;
  assign n3715 = ~n2891 & ~n3712;
  assign n3716 = n3714 & ~n3715;
  assign n3717 = ~n3711 & ~n3716;
  assign n3718 = n3644 & ~n3717;
  assign n3719 = pi592 & ~n2912;
  assign n3720 = ~pi592 & ~n2891;
  assign n3721 = ~n3719 & ~n3720;
  assign n3722 = ~n3644 & n3721;
  assign n3723 = ~n3718 & ~n3722;
  assign n3724 = pi1199 & n3723;
  assign n3725 = n2891 & ~n58919;
  assign n3726 = n58919 & n3721;
  assign n3727 = ~n3725 & ~n3726;
  assign n3728 = n58910 & ~n3727;
  assign n3729 = ~pi1196 & ~n58919;
  assign n3730 = n3721 & ~n3729;
  assign n3731 = ~pi1196 & n3725;
  assign n3732 = ~n3730 & ~n3731;
  assign n3733 = ~n58910 & ~n3732;
  assign n3734 = ~pi1199 & ~n3733;
  assign n3735 = ~pi1199 & ~n3728;
  assign n3736 = ~n3733 & n3735;
  assign n3737 = ~n3728 & n3734;
  assign n3738 = ~n3724 & ~n58925;
  assign n3739 = ~n3705 & ~n3706;
  assign n3740 = ~pi374 & ~n58926;
  assign n3741 = ~pi1198 & ~n58926;
  assign n3742 = pi1198 & ~n3721;
  assign n3743 = ~pi1198 & n58925;
  assign n3744 = ~pi1198 & pi1199;
  assign n3745 = n3723 & n3744;
  assign n3746 = ~n3742 & ~n3745;
  assign n3747 = ~n3743 & n3746;
  assign n3748 = ~n3741 & ~n3742;
  assign n3749 = pi374 & ~n58927;
  assign n3750 = ~n3740 & ~n3749;
  assign n3751 = ~pi369 & ~n3750;
  assign n3752 = ~pi374 & ~n58927;
  assign n3753 = pi374 & ~n58926;
  assign n3754 = ~n3752 & ~n3753;
  assign n3755 = pi369 & ~n3754;
  assign n3756 = ~n3751 & ~n3755;
  assign n3757 = n58906 & n3756;
  assign n3758 = pi369 & ~pi374;
  assign n3759 = ~pi369 & pi374;
  assign n3760 = ~pi369 & ~pi374;
  assign n3761 = pi369 & pi374;
  assign n3762 = ~n3760 & ~n3761;
  assign n3763 = ~n3758 & ~n3759;
  assign n3764 = n58927 & ~n58928;
  assign n3765 = n58926 & n58928;
  assign n3766 = pi369 & ~n3750;
  assign n3767 = ~pi369 & ~n3754;
  assign n3768 = ~n3766 & ~n3767;
  assign n3769 = ~n3764 & ~n3765;
  assign n3770 = ~n58906 & n58929;
  assign n3771 = ~pi370 & ~n3756;
  assign n3772 = pi370 & ~n58929;
  assign n3773 = ~n3771 & ~n3772;
  assign n3774 = ~pi371 & ~n3773;
  assign n3775 = ~pi370 & ~n58929;
  assign n3776 = pi370 & ~n3756;
  assign n3777 = ~n3775 & ~n3776;
  assign n3778 = pi371 & ~n3777;
  assign n3779 = ~n3774 & ~n3778;
  assign n3780 = ~n3757 & ~n3770;
  assign n3781 = ~pi373 & ~n58930;
  assign n3782 = ~pi384 & ~pi442;
  assign n3783 = pi384 & pi442;
  assign n3784 = pi384 & ~pi442;
  assign n3785 = ~pi384 & pi442;
  assign n3786 = ~n3784 & ~n3785;
  assign n3787 = ~n3782 & ~n3783;
  assign n3788 = pi440 & ~n58931;
  assign n3789 = ~pi440 & n58931;
  assign n3790 = ~n3788 & ~n3789;
  assign n3791 = pi375 & ~n3790;
  assign n3792 = ~pi375 & n3790;
  assign n3793 = pi375 & n3790;
  assign n3794 = ~pi375 & ~n3790;
  assign n3795 = ~n3793 & ~n3794;
  assign n3796 = ~n3791 & ~n3792;
  assign n3797 = n58906 & ~n58929;
  assign n3798 = ~n58906 & ~n3756;
  assign n3799 = pi370 & n3756;
  assign n3800 = ~pi370 & n58929;
  assign n3801 = ~pi371 & ~n3800;
  assign n3802 = ~pi371 & ~n3777;
  assign n3803 = ~n3799 & n3801;
  assign n3804 = pi370 & n58929;
  assign n3805 = ~pi370 & n3756;
  assign n3806 = pi371 & ~n3805;
  assign n3807 = pi371 & ~n3773;
  assign n3808 = ~n3804 & n3806;
  assign n3809 = ~n58933 & ~n58934;
  assign n3810 = ~n3797 & ~n3798;
  assign n3811 = pi373 & ~n58935;
  assign n3812 = ~n58932 & ~n3811;
  assign n3813 = ~n3781 & n3812;
  assign n3814 = pi373 & ~n58930;
  assign n3815 = ~pi373 & ~n58935;
  assign n3816 = n58932 & ~n3815;
  assign n3817 = ~n3814 & n3816;
  assign n3818 = ~pi591 & ~n3817;
  assign n3819 = ~n3813 & n3818;
  assign n3820 = ~n3516 & ~n3819;
  assign n3821 = ~pi373 & n58930;
  assign n3822 = pi373 & n58935;
  assign n3823 = ~n3781 & ~n3811;
  assign n3824 = ~n3821 & ~n3822;
  assign n3825 = ~pi375 & n58936;
  assign n3826 = pi373 & n58930;
  assign n3827 = ~pi373 & n58935;
  assign n3828 = ~n3814 & ~n3815;
  assign n3829 = ~n3826 & ~n3827;
  assign n3830 = pi375 & n58937;
  assign n3831 = ~n3790 & ~n3830;
  assign n3832 = ~n3825 & n3831;
  assign n3833 = ~pi375 & n58937;
  assign n3834 = pi375 & n58936;
  assign n3835 = n3790 & ~n3834;
  assign n3836 = n3790 & ~n3833;
  assign n3837 = ~n3834 & n3836;
  assign n3838 = ~n3833 & n3835;
  assign n3839 = ~pi591 & ~n58938;
  assign n3840 = ~n3832 & n3839;
  assign n3841 = ~n3483 & ~n3508;
  assign n3842 = ~pi334 & n3841;
  assign n3843 = ~n3511 & ~n3512;
  assign n3844 = pi334 & n3843;
  assign n3845 = n58904 & ~n3844;
  assign n3846 = n58904 & ~n3842;
  assign n3847 = ~n3844 & n3846;
  assign n3848 = ~n3842 & n3845;
  assign n3849 = pi334 & n3841;
  assign n3850 = ~pi334 & n3843;
  assign n3851 = ~n58904 & ~n3850;
  assign n3852 = ~n3849 & n3851;
  assign n3853 = pi591 & ~n3852;
  assign n3854 = pi591 & ~n58939;
  assign n3855 = ~n3852 & n3854;
  assign n3856 = ~n58939 & n3853;
  assign n3857 = ~pi590 & ~n58940;
  assign n3858 = ~n3840 & n3857;
  assign n3859 = ~pi590 & ~n3820;
  assign n3860 = n3213 & ~n58941;
  assign n3861 = ~n3210 & n3860;
  assign n3862 = n58827 & n2716;
  assign n3863 = pi1091 & ~n3862;
  assign n3864 = n2683 & ~n3863;
  assign n3865 = ~pi122 & pi1093;
  assign n3866 = ~pi98 & n2727;
  assign n3867 = n3865 & n3866;
  assign n3868 = ~pi1091 & ~n3867;
  assign n3869 = n3864 & ~n3868;
  assign n3870 = n2727 & n3865;
  assign n3871 = ~pi1091 & n3870;
  assign n3872 = ~pi1091 & n3867;
  assign n3873 = ~pi98 & n3871;
  assign n3874 = ~n2683 & n58942;
  assign n3875 = pi75 & ~n3874;
  assign n3876 = ~n3869 & n3875;
  assign n3877 = ~pi39 & ~n2772;
  assign n3878 = ~pi122 & n3866;
  assign n3879 = pi122 & n2729;
  assign n3880 = ~n3878 & ~n3879;
  assign n3881 = pi1093 & ~n3880;
  assign n3882 = n2773 & ~n3881;
  assign n3883 = n3877 & ~n3882;
  assign n3884 = pi1091 & ~n58841;
  assign n3885 = ~n3868 & ~n3884;
  assign n3886 = ~n2822 & n3885;
  assign n3887 = n2822 & n58942;
  assign n3888 = ~n3886 & ~n3887;
  assign n3889 = ~n2790 & n3888;
  assign n3890 = ~pi223 & n2827;
  assign n3891 = ~n2783 & ~n58942;
  assign n3892 = n2783 & ~n3885;
  assign n3893 = n2783 & n3885;
  assign n3894 = ~n2783 & n58942;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = ~n3891 & ~n3892;
  assign n3897 = n2790 & n58943;
  assign n3898 = n3890 & ~n3897;
  assign n3899 = ~n3889 & n3898;
  assign n3900 = n3871 & ~n3890;
  assign n3901 = ~pi98 & n3900;
  assign n3902 = n58942 & ~n3890;
  assign n3903 = ~pi299 & ~n58944;
  assign n3904 = ~n3899 & n3903;
  assign n3905 = n58846 & n58943;
  assign n3906 = ~pi216 & n2852;
  assign n3907 = ~n58846 & n3888;
  assign n3908 = n3906 & ~n3907;
  assign n3909 = ~n3905 & n3906;
  assign n3910 = ~n3907 & n3909;
  assign n3911 = ~n3905 & n3908;
  assign n3912 = n3871 & ~n3906;
  assign n3913 = ~pi98 & n3912;
  assign n3914 = n58942 & ~n3906;
  assign n3915 = pi299 & ~n58946;
  assign n3916 = ~n58945 & n3915;
  assign n3917 = pi39 & ~n3916;
  assign n3918 = pi39 & ~n3904;
  assign n3919 = ~n3916 & n3918;
  assign n3920 = ~n3904 & n3917;
  assign n3921 = ~n3883 & ~n58947;
  assign n3922 = ~pi38 & ~n3921;
  assign n3923 = pi38 & n3871;
  assign n3924 = ~pi98 & n3923;
  assign n3925 = pi38 & n58942;
  assign n3926 = ~pi100 & ~n58948;
  assign n3927 = ~n3922 & n3926;
  assign n3928 = n2719 & ~n58942;
  assign n3929 = pi1091 & ~n2717;
  assign n3930 = ~n3868 & ~n3929;
  assign n3931 = n2719 & ~n3930;
  assign n3932 = ~n2718 & n3928;
  assign n3933 = ~n2719 & ~n58942;
  assign n3934 = n2634 & ~n3933;
  assign n3935 = ~n58949 & n3934;
  assign n3936 = ~n2634 & n58942;
  assign n3937 = pi100 & ~n3936;
  assign n3938 = ~n3935 & n3937;
  assign n3939 = ~pi87 & ~n3938;
  assign n3940 = ~n3927 & n3939;
  assign n3941 = pi122 & n58852;
  assign n3942 = ~n3878 & ~n3941;
  assign n3943 = pi1093 & ~n3942;
  assign n3944 = n2901 & ~n3943;
  assign n3945 = n58815 & ~n2902;
  assign n3946 = ~n3944 & n3945;
  assign n3947 = ~n58942 & ~n3946;
  assign n3948 = pi87 & ~n3947;
  assign n3949 = ~pi75 & ~n3948;
  assign n3950 = ~n3940 & n3949;
  assign n3951 = ~n3876 & ~n3950;
  assign n3952 = pi567 & ~n3951;
  assign n3953 = n2670 & ~n3952;
  assign n3954 = pi567 & n58942;
  assign n3955 = ~n2439 & n3954;
  assign n3956 = ~n3953 & ~n3955;
  assign n3957 = pi592 & n3956;
  assign n3958 = ~n2913 & ~n3957;
  assign n3959 = pi1198 & n3126;
  assign n3960 = ~n3039 & ~n3959;
  assign n3961 = ~n3958 & ~n3960;
  assign n3962 = ~n3040 & n3956;
  assign n3963 = n3094 & ~n3962;
  assign n3964 = pi1198 & ~n3126;
  assign n3965 = ~n3127 & n3956;
  assign n3966 = n3130 & ~n3965;
  assign n3967 = n3964 & ~n3966;
  assign n3968 = ~n3963 & n3967;
  assign n3969 = pi1196 & n58872;
  assign n3970 = n3958 & n3969;
  assign n3971 = ~n58872 & ~n3956;
  assign n3972 = n58853 & ~n3971;
  assign n3973 = ~n3970 & n3972;
  assign n3974 = pi1196 & ~n58872;
  assign n3975 = n3958 & n3974;
  assign n3976 = n58872 & ~n3956;
  assign n3977 = ~n58853 & ~n3976;
  assign n3978 = ~n3975 & n3977;
  assign n3979 = ~n3973 & ~n3978;
  assign n3980 = ~pi1196 & ~n3956;
  assign n3981 = ~pi1198 & ~n3980;
  assign n3982 = ~n3979 & n3981;
  assign n3983 = ~n3968 & ~n3982;
  assign n3984 = ~n3039 & ~n3983;
  assign n3985 = ~pi455 & ~n3958;
  assign n3986 = pi455 & n3956;
  assign n3987 = ~n3985 & ~n3986;
  assign n3988 = pi452 & ~n3987;
  assign n3989 = pi455 & ~n3958;
  assign n3990 = ~pi455 & n3956;
  assign n3991 = ~n3989 & ~n3990;
  assign n3992 = ~pi452 & ~n3991;
  assign n3993 = ~n58872 & ~n3992;
  assign n3994 = ~n3988 & n3993;
  assign n3995 = pi452 & ~n3991;
  assign n3996 = ~pi452 & ~n3987;
  assign n3997 = n58872 & ~n3996;
  assign n3998 = ~n3995 & n3997;
  assign n3999 = pi1196 & ~n3998;
  assign n4000 = pi1196 & ~n3994;
  assign n4001 = ~n3998 & n4000;
  assign n4002 = ~n3994 & n3999;
  assign n4003 = ~pi1196 & n3956;
  assign n4004 = ~pi1198 & ~n4003;
  assign n4005 = ~n58950 & n4004;
  assign n4006 = ~n3126 & ~n3963;
  assign n4007 = ~n3126 & ~n3966;
  assign n4008 = ~n3963 & n4007;
  assign n4009 = ~n3966 & n4006;
  assign n4010 = n3126 & ~n3958;
  assign n4011 = pi1198 & ~n4010;
  assign n4012 = ~n58951 & n4011;
  assign n4013 = ~n3039 & ~n4012;
  assign n4014 = ~n4005 & n4013;
  assign n4015 = n3039 & ~n3958;
  assign n4016 = ~n4014 & ~n4015;
  assign n4017 = ~n3961 & ~n3984;
  assign n4018 = ~n2437 & ~n58952;
  assign n4019 = pi1199 & ~n3958;
  assign n4020 = pi351 & n4019;
  assign n4021 = ~n4018 & ~n4020;
  assign n4022 = ~pi461 & ~n4021;
  assign n4023 = ~n3152 & ~n58952;
  assign n4024 = ~pi351 & n4019;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = pi461 & ~n4025;
  assign n4027 = ~n4022 & ~n4026;
  assign n4028 = ~pi357 & ~n4027;
  assign n4029 = ~pi461 & ~n4025;
  assign n4030 = pi461 & ~n4021;
  assign n4031 = ~n4029 & ~n4030;
  assign n4032 = pi357 & ~n4031;
  assign n4033 = ~n4028 & ~n4032;
  assign n4034 = pi356 & n4033;
  assign n4035 = ~pi357 & ~n4031;
  assign n4036 = pi357 & ~n4027;
  assign n4037 = ~n4035 & ~n4036;
  assign n4038 = ~pi356 & n4037;
  assign n4039 = n58878 & ~n4038;
  assign n4040 = ~pi356 & ~n4037;
  assign n4041 = pi356 & ~n4033;
  assign n4042 = ~n4040 & ~n4041;
  assign n4043 = n58878 & ~n4042;
  assign n4044 = ~n4034 & n4039;
  assign n4045 = pi356 & n4037;
  assign n4046 = ~pi356 & n4033;
  assign n4047 = ~n58878 & ~n4046;
  assign n4048 = ~pi356 & ~n4033;
  assign n4049 = pi356 & ~n4037;
  assign n4050 = ~n4048 & ~n4049;
  assign n4051 = ~n58878 & ~n4050;
  assign n4052 = ~n4045 & n4047;
  assign n4053 = ~pi591 & ~n58954;
  assign n4054 = ~pi591 & ~n58953;
  assign n4055 = ~n58954 & n4054;
  assign n4056 = ~n58953 & n4053;
  assign n4057 = pi591 & ~n3956;
  assign n4058 = pi590 & ~n4057;
  assign n4059 = ~n58955 & n4058;
  assign n4060 = ~pi592 & n3956;
  assign n4061 = ~n3719 & ~n4060;
  assign n4062 = ~n3644 & n4061;
  assign n4063 = n3644 & ~n3956;
  assign n4064 = ~pi1199 & ~n4063;
  assign n4065 = ~n4062 & n4064;
  assign n4066 = ~n3707 & n3956;
  assign n4067 = n3709 & ~n4066;
  assign n4068 = ~n3712 & n3956;
  assign n4069 = n3714 & ~n4068;
  assign n4070 = ~n4067 & ~n4069;
  assign n4071 = n3644 & ~n4070;
  assign n4072 = pi1199 & ~n4062;
  assign n4073 = ~n4071 & n4072;
  assign n4074 = pi1199 & ~n4070;
  assign n4075 = ~pi1199 & ~n3956;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = n3644 & ~n4076;
  assign n4078 = ~n4062 & ~n4077;
  assign n4079 = ~n4065 & ~n4073;
  assign n4080 = pi374 & ~n58956;
  assign n4081 = ~pi1198 & ~n58956;
  assign n4082 = pi1198 & n4061;
  assign n4083 = ~pi1198 & n58956;
  assign n4084 = pi1198 & ~n4061;
  assign n4085 = ~n4083 & ~n4084;
  assign n4086 = ~n4081 & ~n4082;
  assign n4087 = ~pi374 & n58957;
  assign n4088 = ~pi374 & ~n58957;
  assign n4089 = pi374 & n58956;
  assign n4090 = ~n4088 & ~n4089;
  assign n4091 = ~n4080 & ~n4087;
  assign n4092 = ~pi369 & n58958;
  assign n4093 = pi374 & n58957;
  assign n4094 = ~pi374 & ~n58956;
  assign n4095 = ~pi374 & n58956;
  assign n4096 = pi374 & ~n58957;
  assign n4097 = ~n4095 & ~n4096;
  assign n4098 = ~n4093 & ~n4094;
  assign n4099 = pi369 & n58959;
  assign n4100 = pi369 & ~n58959;
  assign n4101 = ~pi369 & ~n58958;
  assign n4102 = ~n4100 & ~n4101;
  assign n4103 = ~n4092 & ~n4099;
  assign n4104 = pi370 & n58960;
  assign n4105 = pi369 & n58958;
  assign n4106 = ~pi369 & n58959;
  assign n4107 = ~pi369 & ~n58959;
  assign n4108 = pi369 & ~n58958;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = ~n4105 & ~n4106;
  assign n4111 = ~pi370 & n58961;
  assign n4112 = ~pi370 & ~n58961;
  assign n4113 = pi370 & ~n58960;
  assign n4114 = ~n4112 & ~n4113;
  assign n4115 = ~n4104 & ~n4111;
  assign n4116 = pi371 & ~n58962;
  assign n4117 = pi373 & ~pi375;
  assign n4118 = ~pi373 & pi375;
  assign n4119 = ~n4117 & ~n4118;
  assign n4120 = n3790 & n4119;
  assign n4121 = ~n3790 & ~n4119;
  assign n4122 = pi373 & ~n58932;
  assign n4123 = ~pi373 & n58932;
  assign n4124 = ~n4122 & ~n4123;
  assign n4125 = pi373 & ~n3790;
  assign n4126 = ~pi373 & n3790;
  assign n4127 = ~n4125 & ~n4126;
  assign n4128 = pi375 & n4127;
  assign n4129 = ~pi375 & ~n4127;
  assign n4130 = ~n4128 & ~n4129;
  assign n4131 = ~n4120 & ~n4121;
  assign n4132 = pi370 & n58961;
  assign n4133 = ~pi370 & n58960;
  assign n4134 = ~pi370 & ~n58960;
  assign n4135 = pi370 & ~n58961;
  assign n4136 = ~n4134 & ~n4135;
  assign n4137 = ~n4132 & ~n4133;
  assign n4138 = ~pi371 & ~n58964;
  assign n4139 = ~n58963 & ~n4138;
  assign n4140 = ~n4116 & n4139;
  assign n4141 = pi371 & ~n58964;
  assign n4142 = ~pi371 & ~n58962;
  assign n4143 = n58963 & ~n4142;
  assign n4144 = ~n4141 & n4143;
  assign n4145 = ~n4140 & ~n4144;
  assign n4146 = pi371 & n58964;
  assign n4147 = ~pi371 & n58962;
  assign n4148 = n58963 & ~n4147;
  assign n4149 = ~n4141 & ~n4142;
  assign n4150 = n58963 & ~n4149;
  assign n4151 = ~n4146 & n4148;
  assign n4152 = pi371 & n58962;
  assign n4153 = ~pi371 & n58964;
  assign n4154 = ~n58963 & ~n4153;
  assign n4155 = ~n4116 & ~n4138;
  assign n4156 = ~n58963 & ~n4155;
  assign n4157 = ~n4152 & n4154;
  assign n4158 = ~pi591 & ~n58966;
  assign n4159 = ~n58965 & n4158;
  assign n4160 = ~pi591 & ~n58965;
  assign n4161 = ~n58966 & n4160;
  assign n4162 = ~pi591 & ~n4145;
  assign n4163 = n2773 & ~n58888;
  assign n4164 = n3883 & ~n4163;
  assign n4165 = n2729 & ~n58894;
  assign n4166 = pi122 & ~n4165;
  assign n4167 = ~n58894 & n3866;
  assign n4168 = ~pi122 & ~n4167;
  assign n4169 = pi1093 & ~n4168;
  assign n4170 = ~n58894 & n3881;
  assign n4171 = ~n4166 & n4169;
  assign n4172 = n2773 & ~n58968;
  assign n4173 = n4164 & ~n4172;
  assign n4174 = n58888 & n3867;
  assign n4175 = ~pi1091 & n4174;
  assign n4176 = n58888 & n58942;
  assign n4177 = n3865 & n4167;
  assign n4178 = ~n58894 & n3867;
  assign n4179 = ~pi1091 & n58970;
  assign n4180 = ~n58894 & n58942;
  assign n4181 = n58888 & n58971;
  assign n4182 = ~n58894 & n58969;
  assign n4183 = ~n58843 & ~n58972;
  assign n4184 = ~n2823 & ~n58972;
  assign n4185 = ~n2790 & n4184;
  assign n4186 = ~n2819 & ~n58972;
  assign n4187 = n2790 & n4186;
  assign n4188 = n3890 & ~n4187;
  assign n4189 = ~n4185 & n4188;
  assign n4190 = n3890 & ~n4185;
  assign n4191 = ~n4187 & n4190;
  assign n4192 = n3890 & ~n4183;
  assign n4193 = ~n3890 & n58972;
  assign n4194 = ~n3890 & n58969;
  assign n4195 = ~pi299 & ~n4194;
  assign n4196 = ~n3890 & n58971;
  assign n4197 = ~pi299 & ~n4196;
  assign n4198 = ~n4195 & ~n4197;
  assign n4199 = ~pi299 & ~n4193;
  assign n4200 = ~n58973 & ~n58974;
  assign n4201 = pi1093 & ~n2783;
  assign n4202 = n58846 & n4201;
  assign n4203 = n2822 & ~n58846;
  assign n4204 = n3906 & ~n4203;
  assign n4205 = ~n4202 & n4204;
  assign n4206 = n58847 & n3906;
  assign n4207 = n58842 & n4205;
  assign n4208 = pi299 & ~n58972;
  assign n4209 = ~n3906 & n58969;
  assign n4210 = pi299 & ~n4209;
  assign n4211 = ~n3906 & n58971;
  assign n4212 = pi299 & ~n4211;
  assign n4213 = ~n4210 & ~n4212;
  assign n4214 = n58846 & n4186;
  assign n4215 = ~n58846 & n4184;
  assign n4216 = n3906 & ~n4215;
  assign n4217 = n3906 & ~n4214;
  assign n4218 = ~n4215 & n4217;
  assign n4219 = ~n4214 & n4216;
  assign n4220 = ~n4213 & ~n58976;
  assign n4221 = ~n58975 & n4208;
  assign n4222 = pi39 & ~n58977;
  assign n4223 = pi39 & ~n4200;
  assign n4224 = ~n58977 & n4223;
  assign n4225 = ~n4200 & n4222;
  assign n4226 = ~n4173 & ~n58978;
  assign n4227 = ~pi38 & ~n4226;
  assign n4228 = pi38 & n58969;
  assign n4229 = ~pi100 & ~n4228;
  assign n4230 = pi38 & n58971;
  assign n4231 = ~pi100 & ~n4230;
  assign n4232 = ~n4229 & ~n4231;
  assign n4233 = ~n4227 & ~n4232;
  assign n4234 = ~n2717 & ~n58972;
  assign n4235 = ~pi1091 & ~n58972;
  assign n4236 = ~n2720 & ~n58972;
  assign n4237 = ~n4235 & ~n4236;
  assign n4238 = ~n4234 & n4237;
  assign n4239 = n2675 & n2718;
  assign n4240 = ~n2678 & n2680;
  assign n4241 = ~n2675 & ~n4240;
  assign n4242 = ~n4235 & n4241;
  assign n4243 = ~n3929 & n4242;
  assign n4244 = ~n4239 & ~n4243;
  assign n4245 = pi228 & ~n4244;
  assign n4246 = pi228 & n4241;
  assign n4247 = n58972 & ~n4246;
  assign n4248 = pi232 & ~n4247;
  assign n4249 = ~n4245 & n4248;
  assign n4250 = ~pi232 & ~n58972;
  assign n4251 = ~n2721 & n4250;
  assign n4252 = n2634 & ~n4251;
  assign n4253 = ~n4249 & n4252;
  assign n4254 = ~n2634 & n58972;
  assign n4255 = pi100 & ~n4254;
  assign n4256 = ~n4253 & n4255;
  assign n4257 = pi100 & ~n4238;
  assign n4258 = ~n4233 & ~n58979;
  assign n4259 = ~pi87 & ~n4258;
  assign n4260 = ~n58815 & n58969;
  assign n4261 = pi87 & ~n4260;
  assign n4262 = ~n58815 & n58971;
  assign n4263 = pi87 & ~n4262;
  assign n4264 = ~n4261 & ~n4263;
  assign n4265 = n2901 & ~n58888;
  assign n4266 = n2901 & n58894;
  assign n4267 = n3946 & ~n4266;
  assign n4268 = ~n4265 & n4267;
  assign n4269 = ~n4264 & ~n4268;
  assign n4270 = ~n4259 & ~n4269;
  assign n4271 = ~pi75 & ~n4270;
  assign n4272 = ~n2683 & n58969;
  assign n4273 = pi75 & ~n4272;
  assign n4274 = ~n2683 & n58971;
  assign n4275 = pi75 & ~n4274;
  assign n4276 = ~n4273 & ~n4275;
  assign n4277 = n3864 & ~n4235;
  assign n4278 = ~n4276 & ~n4277;
  assign n4279 = ~n4271 & ~n4278;
  assign n4280 = ~pi592 & pi1196;
  assign n4281 = pi567 & n58969;
  assign n4282 = ~n2439 & n4281;
  assign n4283 = n4167 & n4282;
  assign n4284 = n4280 & ~n4283;
  assign n4285 = ~n4279 & n4284;
  assign n4286 = pi567 & n58971;
  assign n4287 = ~n2439 & n4286;
  assign n4288 = ~pi592 & ~pi1196;
  assign n4289 = ~n4287 & n4288;
  assign n4290 = n4263 & ~n4267;
  assign n4291 = n2725 & ~n58971;
  assign n4292 = n3877 & ~n4172;
  assign n4293 = ~n2834 & ~n2856;
  assign n4294 = ~n58971 & n4293;
  assign n4295 = ~n2819 & ~n58971;
  assign n4296 = n2790 & n4295;
  assign n4297 = ~n2823 & ~n58971;
  assign n4298 = ~n2790 & n4297;
  assign n4299 = n3890 & ~n4298;
  assign n4300 = ~n4296 & n4299;
  assign n4301 = n4197 & ~n4300;
  assign n4302 = n58846 & n4295;
  assign n4303 = ~n58846 & n4297;
  assign n4304 = n3906 & ~n4303;
  assign n4305 = ~n4302 & n4304;
  assign n4306 = n4212 & ~n4305;
  assign n4307 = pi39 & ~n4306;
  assign n4308 = ~n4301 & n4307;
  assign n4309 = pi39 & ~n4301;
  assign n4310 = ~n4306 & n4309;
  assign n4311 = pi39 & ~n4294;
  assign n4312 = ~n4292 & ~n58980;
  assign n4313 = ~pi38 & ~n4312;
  assign n4314 = n4231 & ~n4313;
  assign n4315 = ~n4291 & ~n4314;
  assign n4316 = ~pi87 & ~n4315;
  assign n4317 = ~n4290 & ~n4316;
  assign n4318 = ~pi75 & ~n4317;
  assign n4319 = ~pi1091 & ~n58970;
  assign n4320 = n3864 & ~n4319;
  assign n4321 = n4275 & ~n4320;
  assign n4322 = ~n4318 & ~n4321;
  assign n4323 = n4289 & ~n4322;
  assign n4324 = ~n4285 & ~n4323;
  assign n4325 = pi567 & ~n4324;
  assign n4326 = ~n4284 & ~n4289;
  assign n4327 = ~n2670 & ~n4326;
  assign n4328 = pi1199 & ~n4327;
  assign n4329 = ~n4325 & n4328;
  assign n4330 = pi299 & ~n58969;
  assign n4331 = ~n2819 & ~n58969;
  assign n4332 = n58846 & n4331;
  assign n4333 = ~n2823 & ~n58969;
  assign n4334 = ~n58846 & n4333;
  assign n4335 = n3906 & ~n4334;
  assign n4336 = ~n4332 & n4335;
  assign n4337 = n4210 & ~n4336;
  assign n4338 = ~n58975 & n4330;
  assign n4339 = n2790 & n4201;
  assign n4340 = ~n2790 & n2822;
  assign n4341 = n3890 & ~n4340;
  assign n4342 = ~n4339 & n4341;
  assign n4343 = n58843 & n3890;
  assign n4344 = n58842 & n4342;
  assign n4345 = ~pi299 & ~n58969;
  assign n4346 = n2790 & n4331;
  assign n4347 = ~n2790 & n4333;
  assign n4348 = n3890 & ~n4347;
  assign n4349 = ~n4346 & n4348;
  assign n4350 = n4195 & ~n4349;
  assign n4351 = ~n58982 & n4345;
  assign n4352 = pi39 & ~n58983;
  assign n4353 = pi39 & ~n58981;
  assign n4354 = ~n58983 & n4353;
  assign n4355 = ~n58981 & n4352;
  assign n4356 = ~n4164 & ~n58984;
  assign n4357 = ~pi38 & ~n4356;
  assign n4358 = n4229 & ~n4357;
  assign n4359 = n2725 & ~n58969;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = ~pi87 & ~n4360;
  assign n4362 = n3946 & ~n4265;
  assign n4363 = n4261 & ~n4362;
  assign n4364 = ~n4361 & ~n4363;
  assign n4365 = ~pi75 & ~n4364;
  assign n4366 = ~pi1091 & ~n4174;
  assign n4367 = n3864 & ~n4366;
  assign n4368 = n4273 & ~n4367;
  assign n4369 = ~n4365 & ~n4368;
  assign n4370 = pi567 & ~n4369;
  assign n4371 = n2670 & ~n4370;
  assign n4372 = n4280 & ~n4282;
  assign n4373 = ~n4371 & n4372;
  assign n4374 = ~pi1199 & ~n4003;
  assign n4375 = ~n4373 & n4374;
  assign n4376 = ~n3450 & ~n4375;
  assign n4377 = ~n4329 & n4376;
  assign n4378 = n2913 & n3450;
  assign n4379 = ~n3957 & ~n4378;
  assign n4380 = ~n4377 & n4379;
  assign n4381 = ~n3214 & n4380;
  assign n4382 = n3214 & n3958;
  assign n4383 = ~pi333 & ~n4380;
  assign n4384 = ~pi1197 & ~n4380;
  assign n4385 = pi1197 & ~n3958;
  assign n4386 = ~n4384 & ~n4385;
  assign n4387 = pi333 & ~n4386;
  assign n4388 = ~n4383 & ~n4387;
  assign n4389 = ~n4381 & ~n4382;
  assign n4390 = pi391 & n58985;
  assign n4391 = n3465 & ~n3958;
  assign n4392 = ~n3465 & ~n4380;
  assign n4393 = ~pi333 & ~n4386;
  assign n4394 = pi333 & ~n4380;
  assign n4395 = ~n4393 & ~n4394;
  assign n4396 = ~n4391 & ~n4392;
  assign n4397 = ~pi391 & n58986;
  assign n4398 = ~pi391 & ~n58986;
  assign n4399 = pi391 & ~n58985;
  assign n4400 = ~n4398 & ~n4399;
  assign n4401 = ~n4390 & ~n4397;
  assign n4402 = pi392 & n58987;
  assign n4403 = pi393 & ~n58905;
  assign n4404 = ~pi393 & n58905;
  assign n4405 = pi393 & n58905;
  assign n4406 = ~pi393 & ~n58905;
  assign n4407 = ~n4405 & ~n4406;
  assign n4408 = ~n4403 & ~n4404;
  assign n4409 = ~pi391 & ~n58985;
  assign n4410 = pi391 & ~n58986;
  assign n4411 = ~n4409 & ~n4410;
  assign n4412 = ~pi392 & n4411;
  assign n4413 = n58988 & ~n4412;
  assign n4414 = ~pi392 & ~n4411;
  assign n4415 = pi392 & ~n58987;
  assign n4416 = ~n4414 & ~n4415;
  assign n4417 = n58988 & ~n4416;
  assign n4418 = ~n4402 & n4413;
  assign n4419 = ~pi392 & n58987;
  assign n4420 = pi392 & n4411;
  assign n4421 = ~n58988 & ~n4420;
  assign n4422 = ~pi392 & ~n58987;
  assign n4423 = pi392 & ~n4411;
  assign n4424 = ~n4422 & ~n4423;
  assign n4425 = ~n58988 & ~n4424;
  assign n4426 = ~n4419 & n4421;
  assign n4427 = pi591 & ~n58990;
  assign n4428 = pi591 & ~n58989;
  assign n4429 = ~n58990 & n4428;
  assign n4430 = ~n58989 & n4427;
  assign n4431 = ~pi590 & ~n58991;
  assign n4432 = ~n58967 & n4431;
  assign n4433 = ~n3213 & ~n4432;
  assign n4434 = ~n4059 & n4433;
  assign n4435 = ~pi588 & ~n4434;
  assign n4436 = ~n3861 & n4435;
  assign n4437 = ~pi56 & ~pi62;
  assign n4438 = ~pi57 & ~pi59;
  assign n4439 = n4437 & n4438;
  assign n4440 = ~pi55 & n4437;
  assign n4441 = ~pi59 & n4440;
  assign n4442 = ~pi57 & n4441;
  assign n4443 = ~pi55 & n4439;
  assign n4444 = pi426 & ~pi430;
  assign n4445 = ~pi426 & pi430;
  assign n4446 = ~n4444 & ~n4445;
  assign n4447 = ~pi433 & ~pi451;
  assign n4448 = pi433 & pi451;
  assign n4449 = pi433 & ~pi451;
  assign n4450 = ~pi433 & pi451;
  assign n4451 = ~n4449 & ~n4450;
  assign n4452 = ~n4447 & ~n4448;
  assign n4453 = pi449 & n58993;
  assign n4454 = ~pi449 & ~n58993;
  assign n4455 = ~n4453 & ~n4454;
  assign n4456 = pi445 & ~pi448;
  assign n4457 = ~pi445 & pi448;
  assign n4458 = ~pi445 & ~pi448;
  assign n4459 = pi445 & pi448;
  assign n4460 = ~n4458 & ~n4459;
  assign n4461 = ~n4456 & ~n4457;
  assign n4462 = n4455 & ~n58994;
  assign n4463 = ~n4455 & n58994;
  assign n4464 = pi448 & n4455;
  assign n4465 = ~pi448 & ~n4455;
  assign n4466 = pi448 & ~n4455;
  assign n4467 = ~pi448 & n4455;
  assign n4468 = ~n4466 & ~n4467;
  assign n4469 = ~n4464 & ~n4465;
  assign n4470 = pi445 & n58995;
  assign n4471 = ~pi445 & ~n58995;
  assign n4472 = ~n4470 & ~n4471;
  assign n4473 = ~n4462 & ~n4463;
  assign n4474 = n4446 & ~n58996;
  assign n4475 = ~n4446 & n58996;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = ~pi437 & ~pi453;
  assign n4478 = pi437 & pi453;
  assign n4479 = pi437 & ~pi453;
  assign n4480 = ~pi437 & pi453;
  assign n4481 = ~n4479 & ~n4480;
  assign n4482 = ~n4477 & ~n4478;
  assign n4483 = pi464 & ~n58997;
  assign n4484 = ~pi464 & n58997;
  assign n4485 = ~n4483 & ~n4484;
  assign n4486 = pi417 & ~pi418;
  assign n4487 = ~pi417 & pi418;
  assign n4488 = ~pi417 & ~pi418;
  assign n4489 = pi417 & pi418;
  assign n4490 = ~n4488 & ~n4489;
  assign n4491 = ~n4486 & ~n4487;
  assign n4492 = n4485 & ~n58998;
  assign n4493 = ~n4485 & n58998;
  assign n4494 = pi437 & n58998;
  assign n4495 = ~pi437 & ~n58998;
  assign n4496 = ~n4494 & ~n4495;
  assign n4497 = pi453 & ~pi464;
  assign n4498 = ~pi453 & pi464;
  assign n4499 = ~n4497 & ~n4498;
  assign n4500 = n4496 & n4499;
  assign n4501 = ~n4496 & ~n4499;
  assign n4502 = ~n4500 & ~n4501;
  assign n4503 = pi464 & ~n58998;
  assign n4504 = ~pi464 & n58998;
  assign n4505 = ~n4503 & ~n4504;
  assign n4506 = n58997 & n4505;
  assign n4507 = ~n58997 & ~n4505;
  assign n4508 = ~n4506 & ~n4507;
  assign n4509 = ~n4492 & ~n4493;
  assign n4510 = ~pi415 & ~pi431;
  assign n4511 = pi415 & pi431;
  assign n4512 = pi415 & ~pi431;
  assign n4513 = ~pi415 & pi431;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = ~n4510 & ~n4511;
  assign n4516 = pi416 & ~pi438;
  assign n4517 = ~pi416 & pi438;
  assign n4518 = ~n4516 & ~n4517;
  assign n4519 = ~n59000 & n4518;
  assign n4520 = n59000 & ~n4518;
  assign n4521 = n59000 & n4518;
  assign n4522 = ~n59000 & ~n4518;
  assign n4523 = ~n4521 & ~n4522;
  assign n4524 = ~n4519 & ~n4520;
  assign n4525 = ~n58999 & n59001;
  assign n4526 = n58999 & ~n59001;
  assign n4527 = pi1197 & ~n4526;
  assign n4528 = ~n4525 & n4527;
  assign n4529 = pi421 & ~pi454;
  assign n4530 = ~pi421 & pi454;
  assign n4531 = ~n4529 & ~n4530;
  assign n4532 = pi432 & ~pi459;
  assign n4533 = ~pi432 & pi459;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = n4531 & ~n4534;
  assign n4536 = ~n4531 & n4534;
  assign n4537 = ~n4535 & ~n4536;
  assign n4538 = ~pi423 & ~pi424;
  assign n4539 = pi423 & pi424;
  assign n4540 = pi423 & ~pi424;
  assign n4541 = ~pi423 & pi424;
  assign n4542 = ~n4540 & ~n4541;
  assign n4543 = ~n4538 & ~n4539;
  assign n4544 = pi419 & ~pi420;
  assign n4545 = ~pi419 & pi420;
  assign n4546 = ~pi419 & ~pi420;
  assign n4547 = pi419 & pi420;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = ~n4544 & ~n4545;
  assign n4550 = ~n59002 & n59003;
  assign n4551 = n59002 & ~n59003;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = n4537 & n4552;
  assign n4554 = ~n4537 & ~n4552;
  assign n4555 = pi432 & ~n59002;
  assign n4556 = ~pi432 & n59002;
  assign n4557 = ~n4555 & ~n4556;
  assign n4558 = pi459 & ~n59003;
  assign n4559 = ~pi459 & n59003;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = n4557 & ~n4560;
  assign n4562 = ~n4557 & n4560;
  assign n4563 = ~n4561 & ~n4562;
  assign n4564 = n4531 & n4563;
  assign n4565 = ~n4531 & ~n4563;
  assign n4566 = ~n4564 & ~n4565;
  assign n4567 = pi432 & ~n4531;
  assign n4568 = ~pi432 & n4531;
  assign n4569 = ~n4567 & ~n4568;
  assign n4570 = n59002 & ~n4569;
  assign n4571 = ~n59002 & n4569;
  assign n4572 = ~n4570 & ~n4571;
  assign n4573 = n4560 & n4572;
  assign n4574 = ~n4560 & ~n4572;
  assign n4575 = ~n4573 & ~n4574;
  assign n4576 = ~n4553 & ~n4554;
  assign n4577 = ~pi425 & n59004;
  assign n4578 = pi425 & ~n59004;
  assign n4579 = pi1198 & ~n4578;
  assign n4580 = ~n4577 & n4579;
  assign n4581 = ~n4528 & ~n4580;
  assign n4582 = n2915 & ~n4581;
  assign n4583 = pi429 & ~pi435;
  assign n4584 = ~pi429 & pi435;
  assign n4585 = ~pi429 & ~pi435;
  assign n4586 = pi429 & pi435;
  assign n4587 = ~n4585 & ~n4586;
  assign n4588 = ~n4583 & ~n4584;
  assign n4589 = ~pi434 & ~pi446;
  assign n4590 = pi434 & pi446;
  assign n4591 = pi434 & ~pi446;
  assign n4592 = ~pi434 & pi446;
  assign n4593 = ~n4591 & ~n4592;
  assign n4594 = ~n4589 & ~n4590;
  assign n4595 = pi414 & ~pi422;
  assign n4596 = ~pi414 & pi422;
  assign n4597 = ~n4595 & ~n4596;
  assign n4598 = ~n59006 & n4597;
  assign n4599 = n59006 & ~n4597;
  assign n4600 = n59006 & n4597;
  assign n4601 = ~n59006 & ~n4597;
  assign n4602 = ~n4600 & ~n4601;
  assign n4603 = ~n4598 & ~n4599;
  assign n4604 = n59005 & n59007;
  assign n4605 = ~n59005 & ~n59007;
  assign n4606 = pi429 & ~n59007;
  assign n4607 = ~pi429 & n59007;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = pi435 & n4608;
  assign n4610 = ~pi435 & ~n4608;
  assign n4611 = ~n4609 & ~n4610;
  assign n4612 = ~n4604 & ~n4605;
  assign n4613 = ~pi436 & ~pi444;
  assign n4614 = pi436 & pi444;
  assign n4615 = pi436 & ~pi444;
  assign n4616 = ~pi436 & pi444;
  assign n4617 = ~n4615 & ~n4616;
  assign n4618 = ~n4613 & ~n4614;
  assign n4619 = ~n59008 & n59009;
  assign n4620 = n59008 & ~n59009;
  assign n4621 = ~n59008 & ~n59009;
  assign n4622 = n59008 & n59009;
  assign n4623 = ~n4621 & ~n4622;
  assign n4624 = ~n4619 & ~n4620;
  assign n4625 = ~pi443 & ~n2891;
  assign n4626 = pi443 & ~pi592;
  assign n4627 = ~n2912 & n4626;
  assign n4628 = ~n4625 & ~n4627;
  assign n4629 = ~n59010 & ~n4628;
  assign n4630 = pi443 & ~n2891;
  assign n4631 = ~pi443 & ~pi592;
  assign n4632 = ~n2912 & n4631;
  assign n4633 = ~n4630 & ~n4632;
  assign n4634 = n59010 & ~n4633;
  assign n4635 = ~n2914 & ~n4634;
  assign n4636 = ~n4629 & n4635;
  assign n4637 = ~n2891 & ~n4631;
  assign n4638 = ~n4632 & ~n4637;
  assign n4639 = ~pi444 & ~n4638;
  assign n4640 = ~n2891 & ~n4626;
  assign n4641 = ~n4627 & ~n4640;
  assign n4642 = pi444 & ~n4641;
  assign n4643 = ~n4639 & ~n4642;
  assign n4644 = pi436 & ~n4643;
  assign n4645 = ~pi444 & ~n4641;
  assign n4646 = pi444 & ~n4638;
  assign n4647 = ~n4645 & ~n4646;
  assign n4648 = ~pi436 & ~n4647;
  assign n4649 = n59008 & ~n4648;
  assign n4650 = ~n4644 & n4649;
  assign n4651 = pi436 & ~n4647;
  assign n4652 = ~pi436 & ~n4643;
  assign n4653 = ~n59008 & ~n4652;
  assign n4654 = ~n4651 & n4653;
  assign n4655 = pi1196 & ~n4654;
  assign n4656 = ~n4650 & n4655;
  assign n4657 = pi1196 & ~n4650;
  assign n4658 = ~n4654 & n4657;
  assign n4659 = pi1196 & ~n4636;
  assign n4660 = ~n2985 & n4581;
  assign n4661 = ~n59011 & n4660;
  assign n4662 = ~n4582 & ~n4661;
  assign n4663 = n4476 & ~n4662;
  assign n4664 = pi427 & ~pi428;
  assign n4665 = ~pi427 & pi428;
  assign n4666 = ~pi427 & ~pi428;
  assign n4667 = pi427 & pi428;
  assign n4668 = ~n4666 & ~n4667;
  assign n4669 = ~n4664 & ~n4665;
  assign n4670 = ~n3148 & ~n4476;
  assign n4671 = n59012 & ~n4670;
  assign n4672 = ~n4663 & n4671;
  assign n4673 = ~n3148 & n4476;
  assign n4674 = ~n59012 & ~n4673;
  assign n4675 = pi1199 & ~n4674;
  assign n4676 = n4662 & ~n4675;
  assign n4677 = ~pi590 & ~pi591;
  assign n4678 = n4476 & n4674;
  assign n4679 = n4677 & ~n4678;
  assign n4680 = ~n4676 & n4679;
  assign n4681 = pi428 & ~n4662;
  assign n4682 = ~pi428 & n2915;
  assign n4683 = ~n4681 & ~n4682;
  assign n4684 = ~pi427 & ~n4683;
  assign n4685 = ~pi428 & ~n4662;
  assign n4686 = pi428 & n2915;
  assign n4687 = ~n4685 & ~n4686;
  assign n4688 = pi427 & ~n4687;
  assign n4689 = ~n4684 & ~n4688;
  assign n4690 = pi430 & ~n4689;
  assign n4691 = pi427 & ~n4683;
  assign n4692 = ~pi427 & ~n4687;
  assign n4693 = ~n4691 & ~n4692;
  assign n4694 = ~pi430 & ~n4693;
  assign n4695 = ~n4690 & ~n4694;
  assign n4696 = pi426 & ~n4695;
  assign n4697 = pi430 & ~n4693;
  assign n4698 = ~pi430 & ~n4689;
  assign n4699 = ~n4697 & ~n4698;
  assign n4700 = ~pi426 & ~n4699;
  assign n4701 = ~n4696 & ~n4700;
  assign n4702 = ~pi445 & n4701;
  assign n4703 = pi426 & ~n4699;
  assign n4704 = ~pi426 & ~n4695;
  assign n4705 = ~n4703 & ~n4704;
  assign n4706 = pi445 & n4705;
  assign n4707 = n58995 & ~n4706;
  assign n4708 = pi445 & ~n4705;
  assign n4709 = ~pi445 & ~n4701;
  assign n4710 = ~n4708 & ~n4709;
  assign n4711 = n58995 & ~n4710;
  assign n4712 = ~n4702 & n4707;
  assign n4713 = ~pi445 & n4705;
  assign n4714 = pi445 & n4701;
  assign n4715 = ~n58995 & ~n4714;
  assign n4716 = pi445 & ~n4701;
  assign n4717 = ~pi445 & ~n4705;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = ~n58995 & ~n4718;
  assign n4720 = ~n4713 & n4715;
  assign n4721 = pi1199 & ~n59014;
  assign n4722 = ~n59013 & n4721;
  assign n4723 = ~pi1199 & n4662;
  assign n4724 = n4677 & ~n4723;
  assign n4725 = ~n4722 & n4724;
  assign n4726 = ~n4672 & n4680;
  assign n4727 = n2891 & ~n4677;
  assign n4728 = n3213 & ~n4727;
  assign n4729 = ~n59015 & n4728;
  assign n4730 = n3958 & ~n59012;
  assign n4731 = ~n3958 & ~n4581;
  assign n4732 = n3956 & ~n4631;
  assign n4733 = n59010 & ~n4632;
  assign n4734 = ~n4732 & n4733;
  assign n4735 = n3956 & ~n4626;
  assign n4736 = ~n59010 & ~n4627;
  assign n4737 = ~n4735 & n4736;
  assign n4738 = ~n4734 & ~n4737;
  assign n4739 = pi1196 & ~n4738;
  assign n4740 = ~n3980 & n4581;
  assign n4741 = pi1196 & ~n4737;
  assign n4742 = pi1196 & ~n4734;
  assign n4743 = ~n4737 & n4742;
  assign n4744 = ~n4734 & n4741;
  assign n4745 = ~n4003 & ~n59016;
  assign n4746 = n4581 & ~n4745;
  assign n4747 = ~n4739 & n4740;
  assign n4748 = ~n4731 & ~n59017;
  assign n4749 = n59012 & n4748;
  assign n4750 = ~n4730 & ~n4749;
  assign n4751 = pi430 & ~n4750;
  assign n4752 = ~n59012 & n4748;
  assign n4753 = n3958 & n59012;
  assign n4754 = pi428 & n4748;
  assign n4755 = ~pi428 & n3958;
  assign n4756 = pi427 & ~n4755;
  assign n4757 = ~n4754 & n4756;
  assign n4758 = ~pi428 & n4748;
  assign n4759 = pi428 & n3958;
  assign n4760 = ~pi427 & ~n4759;
  assign n4761 = ~n4758 & n4760;
  assign n4762 = ~n4757 & ~n4761;
  assign n4763 = ~n4752 & ~n4753;
  assign n4764 = ~pi430 & n59018;
  assign n4765 = ~pi430 & ~n59018;
  assign n4766 = pi430 & n4750;
  assign n4767 = ~n4765 & ~n4766;
  assign n4768 = ~n4751 & ~n4764;
  assign n4769 = pi426 & n58996;
  assign n4770 = ~pi426 & ~n58996;
  assign n4771 = ~pi426 & n58996;
  assign n4772 = pi426 & ~n58996;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = ~n4769 & ~n4770;
  assign n4775 = n59019 & n59020;
  assign n4776 = ~pi430 & ~n4750;
  assign n4777 = pi430 & n59018;
  assign n4778 = pi430 & ~n59018;
  assign n4779 = ~pi430 & n4750;
  assign n4780 = ~n4778 & ~n4779;
  assign n4781 = ~n4776 & ~n4777;
  assign n4782 = ~n59020 & n59021;
  assign n4783 = pi426 & ~n59019;
  assign n4784 = ~pi426 & ~n59021;
  assign n4785 = ~n4783 & ~n4784;
  assign n4786 = ~pi445 & ~n4785;
  assign n4787 = ~pi426 & ~n59019;
  assign n4788 = pi426 & ~n59021;
  assign n4789 = ~n4787 & ~n4788;
  assign n4790 = pi445 & ~n4789;
  assign n4791 = ~n4786 & ~n4790;
  assign n4792 = ~pi448 & n4791;
  assign n4793 = ~pi445 & ~n4789;
  assign n4794 = pi445 & ~n4785;
  assign n4795 = ~n4793 & ~n4794;
  assign n4796 = pi448 & n4795;
  assign n4797 = ~n4455 & ~n4796;
  assign n4798 = ~n4792 & n4797;
  assign n4799 = pi448 & n4791;
  assign n4800 = ~pi448 & n4795;
  assign n4801 = n4455 & ~n4800;
  assign n4802 = ~n4799 & n4801;
  assign n4803 = ~n4798 & ~n4802;
  assign n4804 = ~n4775 & ~n4782;
  assign n4805 = ~n58996 & ~n4788;
  assign n4806 = ~n4787 & n4805;
  assign n4807 = n58996 & ~n4784;
  assign n4808 = ~n4783 & n4807;
  assign n4809 = pi1199 & ~n4808;
  assign n4810 = ~n4806 & n4809;
  assign n4811 = pi1199 & ~n59022;
  assign n4812 = ~pi1199 & ~n4748;
  assign n4813 = n4677 & ~n4812;
  assign n4814 = pi1199 & n59022;
  assign n4815 = ~pi1199 & n4748;
  assign n4816 = ~n4814 & ~n4815;
  assign n4817 = n4677 & ~n4816;
  assign n4818 = ~n59023 & n4813;
  assign n4819 = ~n3956 & ~n4677;
  assign n4820 = ~n3213 & ~n4819;
  assign n4821 = ~n59024 & n4820;
  assign n4822 = ~n4729 & ~n4821;
  assign n4823 = pi588 & ~n4822;
  assign n4824 = n58992 & ~n4823;
  assign n4825 = ~n4436 & n4824;
  assign n4826 = ~pi592 & n58873;
  assign n4827 = n3954 & ~n4826;
  assign n4828 = ~n2959 & n3954;
  assign n4829 = ~n4826 & n4828;
  assign n4830 = pi355 & ~pi361;
  assign n4831 = ~pi355 & pi361;
  assign n4832 = ~n4830 & ~n4831;
  assign n4833 = pi458 & ~n58853;
  assign n4834 = ~pi458 & n58853;
  assign n4835 = ~n4833 & ~n4834;
  assign n4836 = n4832 & n4835;
  assign n4837 = ~n4832 & ~n4835;
  assign n4838 = pi361 & ~pi458;
  assign n4839 = ~pi361 & pi458;
  assign n4840 = ~n4838 & ~n4839;
  assign n4841 = n3118 & n4840;
  assign n4842 = ~n3118 & ~n4840;
  assign n4843 = ~n4841 & ~n4842;
  assign n4844 = ~n4836 & ~n4837;
  assign n4845 = pi441 & ~n59025;
  assign n4846 = ~pi441 & n59025;
  assign n4847 = ~pi592 & ~n4846;
  assign n4848 = ~n4845 & n4847;
  assign n4849 = n2959 & n3954;
  assign n4850 = ~n4848 & n4849;
  assign n4851 = pi1196 & ~n4850;
  assign n4852 = ~n4829 & n4851;
  assign n4853 = pi1196 & ~n4827;
  assign n4854 = ~pi1198 & ~n59026;
  assign n4855 = pi350 & ~n58871;
  assign n4856 = ~pi350 & n58871;
  assign n4857 = ~n4855 & ~n4856;
  assign n4858 = ~pi592 & n3954;
  assign n4859 = n4857 & n4858;
  assign n4860 = ~n3126 & n4857;
  assign n4861 = pi1198 & n4858;
  assign n4862 = n4860 & n4861;
  assign n4863 = n3964 & n4859;
  assign n4864 = ~n4854 & ~n59027;
  assign n4865 = ~n3039 & ~n4864;
  assign n4866 = ~pi592 & ~n4865;
  assign n4867 = n3954 & ~n4866;
  assign n4868 = ~n2437 & ~n4867;
  assign n4869 = ~pi356 & ~pi357;
  assign n4870 = pi356 & pi357;
  assign n4871 = pi356 & ~pi357;
  assign n4872 = ~pi356 & pi357;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = ~n4869 & ~n4870;
  assign n4875 = pi461 & n58878;
  assign n4876 = ~pi461 & ~n58878;
  assign n4877 = ~n4875 & ~n4876;
  assign n4878 = ~n59028 & n4877;
  assign n4879 = n59028 & ~n4877;
  assign n4880 = ~n4878 & ~n4879;
  assign n4881 = pi592 & n3954;
  assign n4882 = pi1199 & ~n4881;
  assign n4883 = pi351 & n4882;
  assign n4884 = ~n4880 & ~n4883;
  assign n4885 = ~n4868 & n4884;
  assign n4886 = ~n3152 & ~n4867;
  assign n4887 = ~pi351 & n4882;
  assign n4888 = n4880 & ~n4887;
  assign n4889 = ~n4886 & n4888;
  assign n4890 = pi590 & ~n4889;
  assign n4891 = ~n4885 & n4890;
  assign n4892 = pi592 & ~n3644;
  assign n4893 = n3644 & n58924;
  assign n4894 = pi592 & ~n4893;
  assign n4895 = n3954 & ~n4894;
  assign n4896 = pi1199 & ~n4895;
  assign n4897 = ~n4892 & ~n4896;
  assign n4898 = n58906 & ~n58963;
  assign n4899 = ~n58906 & n58963;
  assign n4900 = pi371 & n58963;
  assign n4901 = ~pi371 & ~n58963;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = pi370 & ~n4902;
  assign n4904 = ~pi370 & n4902;
  assign n4905 = ~n4903 & ~n4904;
  assign n4906 = n58906 & n58963;
  assign n4907 = ~n58906 & ~n58963;
  assign n4908 = ~n4906 & ~n4907;
  assign n4909 = ~n4898 & ~n4899;
  assign n4910 = n58928 & n59029;
  assign n4911 = ~n58928 & ~n59029;
  assign n4912 = pi1198 & ~n4911;
  assign n4913 = ~n4910 & n4912;
  assign n4914 = n4881 & ~n4913;
  assign n4915 = n4897 & n4914;
  assign n4916 = ~pi590 & ~n4858;
  assign n4917 = ~n4915 & n4916;
  assign n4918 = ~n4891 & ~n4917;
  assign n4919 = ~n4868 & ~n4883;
  assign n4920 = pi461 & n4919;
  assign n4921 = n58878 & n59028;
  assign n4922 = ~n58878 & ~n59028;
  assign n4923 = ~n4921 & ~n4922;
  assign n4924 = ~n4886 & ~n4887;
  assign n4925 = ~pi461 & n4924;
  assign n4926 = ~n4923 & ~n4925;
  assign n4927 = ~n4920 & n4926;
  assign n4928 = pi461 & n4924;
  assign n4929 = ~pi461 & n4919;
  assign n4930 = n4923 & ~n4929;
  assign n4931 = ~n4928 & n4930;
  assign n4932 = pi590 & ~n4931;
  assign n4933 = ~pi461 & ~n4924;
  assign n4934 = pi461 & ~n4919;
  assign n4935 = ~n4933 & ~n4934;
  assign n4936 = ~pi357 & ~n4935;
  assign n4937 = ~pi461 & ~n4919;
  assign n4938 = pi461 & ~n4924;
  assign n4939 = ~n4937 & ~n4938;
  assign n4940 = pi357 & ~n4939;
  assign n4941 = ~n4936 & ~n4940;
  assign n4942 = pi356 & ~n4941;
  assign n4943 = ~pi357 & ~n4939;
  assign n4944 = pi357 & ~n4935;
  assign n4945 = ~n4943 & ~n4944;
  assign n4946 = ~pi356 & ~n4945;
  assign n4947 = ~n58878 & ~n4946;
  assign n4948 = ~n4942 & n4947;
  assign n4949 = pi356 & ~n4945;
  assign n4950 = ~pi356 & ~n4941;
  assign n4951 = n58878 & ~n4950;
  assign n4952 = ~n4949 & n4951;
  assign n4953 = ~n4948 & ~n4952;
  assign n4954 = pi590 & ~n4953;
  assign n4955 = ~n4927 & n4932;
  assign n4956 = n4881 & n4897;
  assign n4957 = ~pi370 & ~n58928;
  assign n4958 = pi370 & n58928;
  assign n4959 = ~n4957 & ~n4958;
  assign n4960 = ~pi371 & ~n4959;
  assign n4961 = pi371 & n4959;
  assign n4962 = ~n4960 & ~n4961;
  assign n4963 = ~pi373 & ~n4962;
  assign n4964 = pi373 & n4962;
  assign n4965 = ~n4963 & ~n4964;
  assign n4966 = pi375 & ~n4965;
  assign n4967 = ~pi375 & n4965;
  assign n4968 = ~n4966 & ~n4967;
  assign n4969 = ~n3790 & ~n4968;
  assign n4970 = n3790 & n4968;
  assign n4971 = ~n4969 & ~n4970;
  assign n4972 = n4956 & n4971;
  assign n4973 = ~pi1198 & n4956;
  assign n4974 = ~n4858 & ~n4973;
  assign n4975 = ~n4972 & n4974;
  assign n4976 = ~n4858 & ~n4915;
  assign n4977 = ~pi590 & ~n59031;
  assign n4978 = ~pi591 & ~n4977;
  assign n4979 = ~n59030 & n4978;
  assign n4980 = ~pi591 & ~n4918;
  assign n4981 = ~pi392 & ~n58988;
  assign n4982 = pi392 & n58988;
  assign n4983 = ~n4981 & ~n4982;
  assign n4984 = ~pi391 & n4983;
  assign n4985 = pi391 & ~n4983;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = pi333 & n4986;
  assign n4988 = ~pi333 & ~n4986;
  assign n4989 = pi1197 & ~n4988;
  assign n4990 = ~n4987 & n4989;
  assign n4991 = ~n3450 & ~n4990;
  assign n4992 = ~n4881 & ~n4991;
  assign n4993 = ~pi592 & ~n3363;
  assign n4994 = ~pi592 & n4286;
  assign n4995 = ~n3363 & n4994;
  assign n4996 = n4286 & n4993;
  assign n4997 = n4882 & ~n59033;
  assign n4998 = n4280 & n4281;
  assign n4999 = n3954 & ~n4280;
  assign n5000 = ~pi1199 & ~n4999;
  assign n5001 = ~n4998 & n5000;
  assign n5002 = ~n4997 & ~n5001;
  assign n5003 = n3214 & n58900;
  assign n5004 = ~n4986 & n5003;
  assign n5005 = ~n5002 & ~n5004;
  assign n5006 = ~pi590 & ~n5005;
  assign n5007 = pi1197 & ~n4881;
  assign n5008 = ~pi1197 & ~n5002;
  assign n5009 = ~n5007 & ~n5008;
  assign n5010 = ~pi333 & ~n5009;
  assign n5011 = pi1198 & ~n4881;
  assign n5012 = n5002 & ~n5011;
  assign n5013 = ~n58900 & ~n5012;
  assign n5014 = n5002 & ~n5013;
  assign n5015 = ~n5010 & n5014;
  assign n5016 = ~pi391 & ~n5015;
  assign n5017 = pi333 & ~n5009;
  assign n5018 = ~pi333 & ~n5002;
  assign n5019 = ~n5013 & ~n5018;
  assign n5020 = ~n5017 & n5019;
  assign n5021 = pi391 & ~n5020;
  assign n5022 = ~n5016 & ~n5021;
  assign n5023 = pi392 & ~n5022;
  assign n5024 = ~pi391 & ~n5020;
  assign n5025 = pi391 & ~n5015;
  assign n5026 = ~n5024 & ~n5025;
  assign n5027 = ~pi392 & ~n5026;
  assign n5028 = n58988 & ~n5027;
  assign n5029 = ~n5023 & n5028;
  assign n5030 = pi392 & ~n5026;
  assign n5031 = ~pi392 & ~n5022;
  assign n5032 = ~n58988 & ~n5031;
  assign n5033 = ~n5030 & n5032;
  assign n5034 = ~n5030 & ~n5031;
  assign n5035 = pi393 & ~n5034;
  assign n5036 = ~n5023 & ~n5027;
  assign n5037 = ~pi393 & ~n5036;
  assign n5038 = n58905 & ~n5037;
  assign n5039 = ~n5035 & n5038;
  assign n5040 = pi393 & ~n5036;
  assign n5041 = ~pi393 & ~n5034;
  assign n5042 = ~n58905 & ~n5041;
  assign n5043 = ~n5040 & n5042;
  assign n5044 = ~n5039 & ~n5043;
  assign n5045 = ~n5029 & ~n5033;
  assign n5046 = ~pi590 & ~n59034;
  assign n5047 = ~n4992 & n5006;
  assign n5048 = pi590 & n3954;
  assign n5049 = pi591 & ~n5048;
  assign n5050 = ~n59035 & n5049;
  assign n5051 = ~n59032 & ~n5050;
  assign n5052 = ~pi588 & ~n5051;
  assign n5053 = ~n3213 & ~n58992;
  assign n5054 = ~pi436 & ~pi443;
  assign n5055 = pi436 & pi443;
  assign n5056 = pi436 & ~pi443;
  assign n5057 = ~pi436 & pi443;
  assign n5058 = ~n5056 & ~n5057;
  assign n5059 = ~n5054 & ~n5055;
  assign n5060 = ~pi444 & n59036;
  assign n5061 = pi444 & ~n59036;
  assign n5062 = ~n5060 & ~n5061;
  assign n5063 = n59008 & ~n5062;
  assign n5064 = ~n59008 & n5062;
  assign n5065 = n4280 & ~n5064;
  assign n5066 = n4280 & ~n5063;
  assign n5067 = ~n5064 & n5066;
  assign n5068 = ~n5063 & n5065;
  assign n5069 = n4581 & ~n59037;
  assign n5070 = n4446 & n4455;
  assign n5071 = ~n4446 & ~n4455;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = ~n58994 & ~n59012;
  assign n5074 = n58994 & n59012;
  assign n5075 = pi445 & n59012;
  assign n5076 = ~pi445 & ~n59012;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = pi448 & ~n5077;
  assign n5079 = ~pi448 & n5077;
  assign n5080 = ~n5078 & ~n5079;
  assign n5081 = ~n5073 & ~n5074;
  assign n5082 = ~n5072 & n59038;
  assign n5083 = n5072 & ~n59038;
  assign n5084 = pi1199 & ~n5083;
  assign n5085 = ~n5082 & n5084;
  assign n5086 = n4677 & n4858;
  assign n5087 = ~n5085 & n5086;
  assign n5088 = n5069 & n5087;
  assign n5089 = ~pi592 & n4677;
  assign n5090 = n3954 & ~n5089;
  assign n5091 = pi588 & ~n5090;
  assign n5092 = n4858 & n5069;
  assign n5093 = n4446 & n59038;
  assign n5094 = ~n4446 & ~n59038;
  assign n5095 = pi430 & n59012;
  assign n5096 = ~pi430 & ~n59012;
  assign n5097 = ~n5095 & ~n5096;
  assign n5098 = ~pi426 & ~n5097;
  assign n5099 = pi426 & n5097;
  assign n5100 = ~n5098 & ~n5099;
  assign n5101 = ~pi445 & ~n5100;
  assign n5102 = pi445 & n5100;
  assign n5103 = ~n5101 & ~n5102;
  assign n5104 = ~pi448 & ~n5103;
  assign n5105 = pi448 & n5103;
  assign n5106 = ~n5104 & ~n5105;
  assign n5107 = ~n5093 & ~n5094;
  assign n5108 = n5092 & ~n59039;
  assign n5109 = ~n4881 & ~n5108;
  assign n5110 = n4455 & ~n5109;
  assign n5111 = n5092 & n59039;
  assign n5112 = ~n4881 & ~n5111;
  assign n5113 = ~n4455 & ~n5112;
  assign n5114 = pi1199 & ~n5113;
  assign n5115 = pi1199 & ~n5110;
  assign n5116 = ~n5113 & n5115;
  assign n5117 = ~n5110 & n5114;
  assign n5118 = ~pi1199 & ~n4881;
  assign n5119 = ~n5092 & n5118;
  assign n5120 = n4677 & ~n5119;
  assign n5121 = ~n59040 & n5120;
  assign n5122 = n3954 & ~n4677;
  assign n5123 = pi588 & ~n5122;
  assign n5124 = ~n5121 & n5123;
  assign n5125 = ~n5088 & n5091;
  assign n5126 = n5053 & ~n59041;
  assign n5127 = ~n5052 & n5126;
  assign n5128 = ~pi217 & ~n5127;
  assign n5129 = ~n4825 & n5128;
  assign n5130 = ~n2891 & n3213;
  assign n5131 = ~n3213 & n3956;
  assign n5132 = n58992 & ~n5131;
  assign n5133 = ~n5130 & n5132;
  assign n5134 = n3954 & n5053;
  assign n5135 = pi217 & ~n5134;
  assign n5136 = ~n5133 & n5135;
  assign n5137 = ~pi1161 & ~pi1162;
  assign n5138 = ~pi1163 & n5137;
  assign n5139 = ~n5136 & n5138;
  assign n5140 = ~n5129 & n5139;
  assign n5141 = pi1161 & ~pi1163;
  assign n5142 = n2794 & n5141;
  assign n5143 = ~pi31 & pi1162;
  assign n5144 = n5142 & n5143;
  assign n5145 = ~n5140 & ~n5144;
  assign n5146 = pi98 & pi1092;
  assign n5147 = pi1093 & n5146;
  assign n5148 = ~pi567 & n2794;
  assign n5149 = ~n5147 & ~n5148;
  assign n5150 = ~pi592 & ~n5149;
  assign n5151 = ~pi88 & n2503;
  assign n5152 = n2539 & n5151;
  assign n5153 = n58799 & n5152;
  assign n5154 = n58798 & n5151;
  assign n5155 = n58804 & n59042;
  assign n5156 = n2581 & n5155;
  assign n5157 = n58821 & n2872;
  assign n5158 = n5156 & n5157;
  assign n5159 = ~pi98 & ~n5158;
  assign n5160 = pi1092 & ~n5159;
  assign n5161 = pi1091 & n5147;
  assign n5162 = n58815 & ~n5161;
  assign n5163 = pi87 & n5162;
  assign n5164 = n58854 & ~n5161;
  assign n5165 = ~n5160 & n59043;
  assign n5166 = n58854 & ~n5160;
  assign n5167 = pi51 & n5156;
  assign n5168 = pi90 & pi93;
  assign n5169 = ~pi841 & ~n2579;
  assign n5170 = ~n5168 & n5169;
  assign n5171 = n2614 & n5170;
  assign n5172 = n5155 & n5171;
  assign n5173 = ~n5167 & ~n5172;
  assign n5174 = n58809 & n2872;
  assign n5175 = ~n5173 & n5174;
  assign n5176 = ~pi98 & ~n5175;
  assign n5177 = pi1092 & ~n5176;
  assign n5178 = ~pi87 & n5162;
  assign n5179 = n2672 & ~n5161;
  assign n5180 = ~n5177 & n59045;
  assign n5181 = n2672 & ~n5177;
  assign n5182 = ~n59044 & ~n59046;
  assign n5183 = pi122 & ~n5182;
  assign n5184 = ~n3871 & ~n5147;
  assign n5185 = ~pi122 & n5184;
  assign n5186 = n2878 & ~n5185;
  assign n5187 = n58815 & ~n5186;
  assign n5188 = ~n5183 & ~n5187;
  assign n5189 = ~pi75 & ~n5161;
  assign n5190 = n5162 & ~n5186;
  assign n5191 = ~n5183 & ~n5190;
  assign n5192 = ~pi75 & ~n5191;
  assign n5193 = ~n5188 & n5189;
  assign n5194 = ~n58816 & n5184;
  assign n5195 = pi567 & n2439;
  assign n5196 = ~n5194 & n5195;
  assign n5197 = ~n59047 & n5196;
  assign n5198 = ~n2439 & ~n5184;
  assign n5199 = ~n5148 & ~n5198;
  assign n5200 = ~n5197 & n5199;
  assign n5201 = pi592 & ~n5200;
  assign n5202 = ~n5150 & ~n5201;
  assign n5203 = ~pi367 & ~n5202;
  assign n5204 = pi367 & ~n5149;
  assign n5205 = ~n5203 & ~n5204;
  assign n5206 = n58912 & ~n5205;
  assign n5207 = pi367 & ~n5202;
  assign n5208 = ~pi367 & ~n5149;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = ~n58912 & ~n5209;
  assign n5211 = ~n5206 & ~n5210;
  assign n5212 = ~n58913 & ~n5211;
  assign n5213 = n58912 & ~n5209;
  assign n5214 = ~n58912 & ~n5205;
  assign n5215 = ~n58912 & n5205;
  assign n5216 = n58912 & n5209;
  assign n5217 = ~n5215 & ~n5216;
  assign n5218 = ~n5213 & ~n5214;
  assign n5219 = n58913 & n59048;
  assign n5220 = n58916 & ~n5219;
  assign n5221 = n58916 & ~n5212;
  assign n5222 = ~n5219 & n5221;
  assign n5223 = ~n5212 & n5220;
  assign n5224 = ~n58913 & n59048;
  assign n5225 = n58913 & ~n5211;
  assign n5226 = ~n58916 & ~n5225;
  assign n5227 = ~n58916 & ~n5224;
  assign n5228 = ~n5225 & n5227;
  assign n5229 = ~n5224 & n5226;
  assign n5230 = pi1197 & ~n59050;
  assign n5231 = pi1197 & ~n59049;
  assign n5232 = ~n59050 & n5231;
  assign n5233 = ~n59049 & n5230;
  assign n5234 = ~pi1197 & ~n5149;
  assign n5235 = ~n58911 & ~n5234;
  assign n5236 = ~n59051 & n5235;
  assign n5237 = n58911 & n5202;
  assign n5238 = ~pi1199 & ~n5237;
  assign n5239 = ~n5236 & n5238;
  assign n5240 = ~n4893 & n5202;
  assign n5241 = n4893 & n5149;
  assign n5242 = pi1199 & ~n5241;
  assign n5243 = ~n5240 & ~n5241;
  assign n5244 = pi1199 & n5243;
  assign n5245 = ~n5240 & n5242;
  assign n5246 = ~n5239 & ~n59052;
  assign n5247 = ~pi374 & ~n5246;
  assign n5248 = ~pi1198 & n5239;
  assign n5249 = pi1198 & ~n5202;
  assign n5250 = n3744 & n5243;
  assign n5251 = ~n5249 & ~n5250;
  assign n5252 = ~pi1198 & ~n5246;
  assign n5253 = ~n5249 & ~n5252;
  assign n5254 = ~n5248 & n5251;
  assign n5255 = pi374 & ~n59053;
  assign n5256 = ~n5247 & ~n5255;
  assign n5257 = pi369 & ~n5256;
  assign n5258 = ~pi374 & ~n59053;
  assign n5259 = pi374 & ~n5246;
  assign n5260 = ~n5258 & ~n5259;
  assign n5261 = ~pi369 & ~n5260;
  assign n5262 = n59029 & ~n5261;
  assign n5263 = n59029 & ~n5257;
  assign n5264 = ~n5261 & n5263;
  assign n5265 = ~n5257 & n5262;
  assign n5266 = ~pi369 & ~n5256;
  assign n5267 = pi369 & ~n5260;
  assign n5268 = ~n59029 & ~n5267;
  assign n5269 = ~n59029 & ~n5266;
  assign n5270 = ~n5267 & n5269;
  assign n5271 = ~n5266 & n5268;
  assign n5272 = ~pi591 & ~n59055;
  assign n5273 = ~pi591 & ~n59054;
  assign n5274 = ~n59055 & n5273;
  assign n5275 = ~n59054 & n5272;
  assign n5276 = pi592 & ~n5149;
  assign n5277 = ~pi592 & ~n5200;
  assign n5278 = ~n5276 & ~n5277;
  assign n5279 = n3450 & ~n5278;
  assign n5280 = ~n58883 & n3244;
  assign n5281 = n58883 & ~n3244;
  assign n5282 = n2727 & ~n5281;
  assign n5283 = n2727 & n58885;
  assign n5284 = ~n5280 & n5282;
  assign n5285 = ~n5146 & ~n59057;
  assign n5286 = ~pi412 & ~n5285;
  assign n5287 = n2727 & ~n58885;
  assign n5288 = ~n5146 & ~n5287;
  assign n5289 = pi412 & ~n5288;
  assign n5290 = ~n3226 & ~n5289;
  assign n5291 = ~n5286 & n5290;
  assign n5292 = ~pi412 & ~n5288;
  assign n5293 = pi412 & ~n5285;
  assign n5294 = n3226 & ~n5293;
  assign n5295 = n3226 & ~n5292;
  assign n5296 = ~n5293 & n5295;
  assign n5297 = ~n5292 & n5294;
  assign n5298 = ~pi122 & ~n59058;
  assign n5299 = ~n5291 & n5298;
  assign n5300 = ~n5146 & ~n5299;
  assign n5301 = n2878 & ~n5300;
  assign n5302 = ~n5161 & ~n5301;
  assign n5303 = pi567 & ~n5302;
  assign n5304 = ~pi122 & n2727;
  assign n5305 = ~n5146 & ~n5304;
  assign n5306 = ~n2878 & ~n5161;
  assign n5307 = n2727 & n58894;
  assign n5308 = ~pi122 & ~n5146;
  assign n5309 = ~n5307 & n5308;
  assign n5310 = ~n5306 & ~n5309;
  assign n5311 = ~n5305 & n5310;
  assign n5312 = pi567 & n5311;
  assign n5313 = ~n5148 & ~n5312;
  assign n5314 = ~n5303 & n5313;
  assign n5315 = n2439 & ~n5148;
  assign n5316 = ~n5314 & ~n5315;
  assign n5317 = n58815 & ~n5310;
  assign n5318 = ~n5301 & n5317;
  assign n5319 = n58894 & n5177;
  assign n5320 = ~n58894 & n5146;
  assign n5321 = ~n5319 & ~n5320;
  assign n5322 = n59045 & n5321;
  assign n5323 = n58888 & ~n5146;
  assign n5324 = ~n58888 & ~n5177;
  assign n5325 = pi411 & n5177;
  assign n5326 = ~pi411 & n5146;
  assign n5327 = n58887 & ~n5326;
  assign n5328 = ~n5325 & n5327;
  assign n5329 = ~pi411 & n5177;
  assign n5330 = ~n58887 & ~n5146;
  assign n5331 = ~n3281 & ~n5330;
  assign n5332 = ~n5329 & ~n5331;
  assign n5333 = ~n5328 & ~n5332;
  assign n5334 = n58888 & n5146;
  assign n5335 = ~n58888 & n5177;
  assign n5336 = ~n5334 & ~n5335;
  assign n5337 = ~n5323 & ~n5324;
  assign n5338 = pi411 & n58888;
  assign n5339 = ~n58887 & ~n5329;
  assign n5340 = ~n5328 & ~n5339;
  assign n5341 = n59059 & ~n5338;
  assign n5342 = n5322 & ~n59060;
  assign n5343 = ~n58888 & ~n5160;
  assign n5344 = pi411 & n5160;
  assign n5345 = n5327 & ~n5344;
  assign n5346 = ~pi411 & n5160;
  assign n5347 = ~n5331 & ~n5346;
  assign n5348 = ~n5345 & ~n5347;
  assign n5349 = ~n5323 & ~n5343;
  assign n5350 = n58894 & n5160;
  assign n5351 = n59043 & ~n5350;
  assign n5352 = n58854 & ~n59061;
  assign n5353 = ~n5350 & n5352;
  assign n5354 = ~n59061 & n5351;
  assign n5355 = ~n5342 & ~n59062;
  assign n5356 = ~pi122 & n5307;
  assign n5357 = ~n5299 & ~n5356;
  assign n5358 = ~n5355 & n5357;
  assign n5359 = ~n5318 & ~n5358;
  assign n5360 = ~pi75 & ~n5359;
  assign n5361 = ~n58816 & ~n5311;
  assign n5362 = ~n5301 & n5361;
  assign n5363 = n5195 & ~n5362;
  assign n5364 = ~n5360 & n5363;
  assign n5365 = ~n5316 & ~n5364;
  assign n5366 = n4280 & ~n5365;
  assign n5367 = ~n5313 & ~n5315;
  assign n5368 = ~n5320 & ~n5350;
  assign n5369 = n59043 & n5368;
  assign n5370 = ~n5322 & ~n5369;
  assign n5371 = pi122 & ~n5370;
  assign n5372 = ~n5317 & ~n5371;
  assign n5373 = ~pi75 & ~n5372;
  assign n5374 = n5195 & ~n5361;
  assign n5375 = ~n5373 & n5374;
  assign n5376 = ~n5367 & ~n5375;
  assign n5377 = n4288 & ~n5376;
  assign n5378 = pi1199 & ~n5377;
  assign n5379 = ~n5366 & n5378;
  assign n5380 = ~pi1196 & ~n5149;
  assign n5381 = ~pi1199 & ~n5380;
  assign n5382 = ~n5148 & ~n5303;
  assign n5383 = ~n5315 & ~n5382;
  assign n5384 = n59045 & ~n59059;
  assign n5385 = ~n5352 & ~n5384;
  assign n5386 = ~n5299 & ~n5385;
  assign n5387 = ~pi122 & ~n5299;
  assign n5388 = n2878 & ~n5387;
  assign n5389 = n5162 & ~n5388;
  assign n5390 = ~n5386 & ~n5389;
  assign n5391 = ~pi75 & ~n5390;
  assign n5392 = ~n58816 & n5302;
  assign n5393 = n5195 & ~n5392;
  assign n5394 = pi122 & n59059;
  assign n5395 = ~n5299 & ~n5394;
  assign n5396 = n2878 & ~n5395;
  assign n5397 = n59045 & ~n5396;
  assign n5398 = ~n58815 & n5302;
  assign n5399 = pi122 & n59061;
  assign n5400 = ~n5299 & ~n5399;
  assign n5401 = n2878 & ~n5400;
  assign n5402 = n59043 & ~n5401;
  assign n5403 = ~n5398 & ~n5402;
  assign n5404 = ~n5397 & n5403;
  assign n5405 = ~pi75 & ~n5404;
  assign n5406 = pi75 & n5302;
  assign n5407 = n5195 & ~n5406;
  assign n5408 = ~n5405 & n5407;
  assign n5409 = ~n5391 & n5393;
  assign n5410 = ~n5383 & ~n59063;
  assign n5411 = n4280 & ~n5410;
  assign n5412 = n5381 & ~n5411;
  assign n5413 = ~n5379 & ~n5412;
  assign n5414 = ~n5380 & ~n5411;
  assign n5415 = ~pi1199 & ~n5414;
  assign n5416 = ~n5366 & ~n5377;
  assign n5417 = pi1199 & ~n5416;
  assign n5418 = ~n5276 & ~n5417;
  assign n5419 = ~n5415 & n5418;
  assign n5420 = ~n5276 & ~n5413;
  assign n5421 = ~n3450 & ~n59064;
  assign n5422 = ~n5279 & ~n5421;
  assign n5423 = pi333 & n5422;
  assign n5424 = ~pi1197 & ~n3450;
  assign n5425 = ~n5278 & ~n5424;
  assign n5426 = ~n59064 & n5424;
  assign n5427 = n5278 & ~n5424;
  assign n5428 = n59064 & n5424;
  assign n5429 = ~n5427 & ~n5428;
  assign n5430 = ~n5425 & ~n5426;
  assign n5431 = ~pi333 & ~n59065;
  assign n5432 = n58988 & ~n5431;
  assign n5433 = ~n5423 & n5432;
  assign n5434 = ~pi391 & ~pi392;
  assign n5435 = pi391 & pi392;
  assign n5436 = ~n5434 & ~n5435;
  assign n5437 = pi333 & n59065;
  assign n5438 = ~pi333 & ~n5422;
  assign n5439 = pi333 & ~n59065;
  assign n5440 = ~pi333 & n5422;
  assign n5441 = ~n5439 & ~n5440;
  assign n5442 = ~n5437 & ~n5438;
  assign n5443 = ~n58988 & n59066;
  assign n5444 = n5436 & ~n5443;
  assign n5445 = ~n5433 & n5444;
  assign n5446 = ~n58988 & ~n5431;
  assign n5447 = ~n5423 & n5446;
  assign n5448 = n58988 & n59066;
  assign n5449 = ~n5436 & ~n5448;
  assign n5450 = ~n5447 & n5449;
  assign n5451 = pi591 & ~n5450;
  assign n5452 = pi391 & ~n59066;
  assign n5453 = pi333 & ~n5422;
  assign n5454 = ~pi333 & n59065;
  assign n5455 = ~n5453 & ~n5454;
  assign n5456 = ~pi391 & n5455;
  assign n5457 = ~n5452 & ~n5456;
  assign n5458 = pi392 & ~n5457;
  assign n5459 = pi391 & ~n5455;
  assign n5460 = ~pi391 & n59066;
  assign n5461 = ~n5459 & ~n5460;
  assign n5462 = ~pi392 & n5461;
  assign n5463 = ~n5458 & ~n5462;
  assign n5464 = ~pi393 & n5463;
  assign n5465 = pi392 & ~n5461;
  assign n5466 = ~pi392 & n5457;
  assign n5467 = ~pi392 & ~n5457;
  assign n5468 = pi392 & n5461;
  assign n5469 = ~n5467 & ~n5468;
  assign n5470 = ~n5465 & ~n5466;
  assign n5471 = pi393 & n59067;
  assign n5472 = n58905 & ~n5471;
  assign n5473 = pi393 & ~n59067;
  assign n5474 = ~pi393 & ~n5463;
  assign n5475 = ~n5473 & ~n5474;
  assign n5476 = n58905 & ~n5475;
  assign n5477 = ~n5464 & n5472;
  assign n5478 = pi393 & n5463;
  assign n5479 = ~pi393 & n59067;
  assign n5480 = ~n58905 & ~n5479;
  assign n5481 = pi393 & ~n5463;
  assign n5482 = ~pi393 & ~n59067;
  assign n5483 = ~n5481 & ~n5482;
  assign n5484 = ~n58905 & ~n5483;
  assign n5485 = ~n5478 & n5480;
  assign n5486 = pi591 & ~n59069;
  assign n5487 = ~n59068 & n5486;
  assign n5488 = pi591 & ~n59068;
  assign n5489 = ~n59069 & n5488;
  assign n5490 = ~n5445 & n5451;
  assign n5491 = ~pi590 & ~n59070;
  assign n5492 = ~n59056 & n5491;
  assign n5493 = pi591 & ~n5149;
  assign n5494 = pi590 & ~n5493;
  assign n5495 = n4860 & n5149;
  assign n5496 = ~n4860 & n5278;
  assign n5497 = ~n5495 & ~n5496;
  assign n5498 = pi1198 & ~n5497;
  assign n5499 = ~pi1198 & ~n5380;
  assign n5500 = n58853 & n5149;
  assign n5501 = ~n58853 & n5278;
  assign n5502 = ~n5500 & ~n5501;
  assign n5503 = ~pi355 & ~n5502;
  assign n5504 = pi455 & ~n5149;
  assign n5505 = ~pi455 & ~n5278;
  assign n5506 = ~n5504 & ~n5505;
  assign n5507 = ~pi452 & ~n5506;
  assign n5508 = ~pi455 & ~n5149;
  assign n5509 = pi455 & ~n5278;
  assign n5510 = ~n5508 & ~n5509;
  assign n5511 = pi452 & ~n5510;
  assign n5512 = ~n5507 & ~n5511;
  assign n5513 = pi355 & n5512;
  assign n5514 = ~n5503 & ~n5513;
  assign n5515 = ~pi458 & n5514;
  assign n5516 = pi355 & ~n5502;
  assign n5517 = ~pi355 & n5512;
  assign n5518 = ~n5516 & ~n5517;
  assign n5519 = pi458 & n5518;
  assign n5520 = n2965 & ~n5519;
  assign n5521 = n2965 & ~n5515;
  assign n5522 = ~n5519 & n5521;
  assign n5523 = ~n5515 & n5520;
  assign n5524 = ~pi458 & n5518;
  assign n5525 = pi458 & n5514;
  assign n5526 = ~n2965 & ~n5525;
  assign n5527 = ~n2965 & ~n5524;
  assign n5528 = ~n5525 & n5527;
  assign n5529 = ~n5524 & n5526;
  assign n5530 = pi1196 & ~n59072;
  assign n5531 = pi1196 & ~n59071;
  assign n5532 = ~n59072 & n5531;
  assign n5533 = ~n59071 & n5530;
  assign n5534 = n5499 & ~n59073;
  assign n5535 = ~n5498 & ~n5534;
  assign n5536 = ~n3039 & ~n5535;
  assign n5537 = n3039 & n5278;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = ~n3152 & n5538;
  assign n5540 = pi1199 & ~n5278;
  assign n5541 = ~pi351 & n5540;
  assign n5542 = n4880 & ~n5541;
  assign n5543 = ~n5539 & n5542;
  assign n5544 = ~n2437 & n5538;
  assign n5545 = pi351 & n5540;
  assign n5546 = ~n4880 & ~n5545;
  assign n5547 = ~n5544 & n5546;
  assign n5548 = ~pi591 & ~n5547;
  assign n5549 = ~n5544 & ~n5545;
  assign n5550 = ~pi461 & ~n5549;
  assign n5551 = ~n5539 & ~n5541;
  assign n5552 = pi461 & ~n5551;
  assign n5553 = ~n5550 & ~n5552;
  assign n5554 = pi357 & n5553;
  assign n5555 = ~pi461 & ~n5551;
  assign n5556 = pi461 & ~n5549;
  assign n5557 = ~n5555 & ~n5556;
  assign n5558 = ~pi357 & n5557;
  assign n5559 = ~pi356 & ~n5558;
  assign n5560 = ~pi357 & ~n5557;
  assign n5561 = pi357 & ~n5553;
  assign n5562 = ~n5560 & ~n5561;
  assign n5563 = ~pi356 & ~n5562;
  assign n5564 = ~n5554 & n5559;
  assign n5565 = pi357 & n5557;
  assign n5566 = ~pi357 & n5553;
  assign n5567 = pi356 & ~n5566;
  assign n5568 = ~pi357 & ~n5553;
  assign n5569 = pi357 & ~n5557;
  assign n5570 = ~n5568 & ~n5569;
  assign n5571 = pi356 & ~n5570;
  assign n5572 = ~n5565 & n5567;
  assign n5573 = ~n59074 & ~n59075;
  assign n5574 = ~pi354 & ~n5573;
  assign n5575 = n59028 & n5553;
  assign n5576 = ~n59028 & n5557;
  assign n5577 = ~pi356 & ~n5570;
  assign n5578 = pi356 & ~n5562;
  assign n5579 = ~n5577 & ~n5578;
  assign n5580 = ~n5575 & ~n5576;
  assign n5581 = pi354 & ~n59076;
  assign n5582 = n58877 & ~n5581;
  assign n5583 = n58877 & ~n5574;
  assign n5584 = ~n5581 & n5583;
  assign n5585 = ~n5574 & n5582;
  assign n5586 = pi354 & ~n5573;
  assign n5587 = ~pi354 & ~n59076;
  assign n5588 = ~n58877 & ~n5587;
  assign n5589 = ~n5586 & n5588;
  assign n5590 = ~pi591 & ~n5589;
  assign n5591 = ~n59077 & n5590;
  assign n5592 = ~n5543 & n5548;
  assign n5593 = n5494 & ~n59078;
  assign n5594 = ~pi588 & ~n5593;
  assign n5595 = ~pi588 & ~n5492;
  assign n5596 = ~n5593 & n5595;
  assign n5597 = ~n5492 & n5594;
  assign n5598 = ~n4677 & n5149;
  assign n5599 = pi588 & ~n5598;
  assign n5600 = ~n4581 & n5278;
  assign n5601 = n4581 & ~n5380;
  assign n5602 = pi443 & ~n5149;
  assign n5603 = ~pi443 & ~n5278;
  assign n5604 = ~n5602 & ~n5603;
  assign n5605 = n59009 & n5604;
  assign n5606 = ~pi443 & ~n5149;
  assign n5607 = pi443 & ~n5278;
  assign n5608 = ~n5606 & ~n5607;
  assign n5609 = ~n59009 & n5608;
  assign n5610 = ~n59008 & ~n5609;
  assign n5611 = ~n5605 & n5610;
  assign n5612 = n59009 & n5608;
  assign n5613 = ~n59009 & n5604;
  assign n5614 = n59008 & ~n5613;
  assign n5615 = ~n5612 & n5614;
  assign n5616 = ~n5611 & ~n5615;
  assign n5617 = ~n5612 & ~n5613;
  assign n5618 = ~pi435 & ~n5617;
  assign n5619 = ~pi444 & n5604;
  assign n5620 = pi444 & n5608;
  assign n5621 = ~pi436 & ~n5620;
  assign n5622 = ~pi436 & ~n5619;
  assign n5623 = ~n5620 & n5622;
  assign n5624 = ~n5619 & n5621;
  assign n5625 = ~pi444 & n5608;
  assign n5626 = pi444 & n5604;
  assign n5627 = pi436 & ~n5626;
  assign n5628 = pi436 & ~n5625;
  assign n5629 = ~n5626 & n5628;
  assign n5630 = ~n5625 & n5627;
  assign n5631 = ~n59080 & ~n59081;
  assign n5632 = pi435 & n5631;
  assign n5633 = ~n5618 & ~n5632;
  assign n5634 = ~pi429 & n5633;
  assign n5635 = pi435 & ~n5617;
  assign n5636 = ~pi435 & n5631;
  assign n5637 = ~n5635 & ~n5636;
  assign n5638 = pi429 & n5637;
  assign n5639 = ~n59007 & ~n5638;
  assign n5640 = ~n59007 & ~n5634;
  assign n5641 = ~n5638 & n5640;
  assign n5642 = ~n5634 & n5639;
  assign n5643 = ~pi429 & n5637;
  assign n5644 = pi429 & n5633;
  assign n5645 = n59007 & ~n5644;
  assign n5646 = n59007 & ~n5643;
  assign n5647 = ~n5644 & n5646;
  assign n5648 = ~n5643 & n5645;
  assign n5649 = pi1196 & ~n59083;
  assign n5650 = ~n59082 & n5649;
  assign n5651 = pi1196 & ~n59082;
  assign n5652 = ~n59083 & n5651;
  assign n5653 = pi1196 & ~n5616;
  assign n5654 = n5601 & ~n59084;
  assign n5655 = ~n5600 & ~n5654;
  assign n5656 = pi428 & ~n5655;
  assign n5657 = ~pi428 & n5278;
  assign n5658 = ~n5656 & ~n5657;
  assign n5659 = pi427 & ~n5658;
  assign n5660 = pi428 & ~n5278;
  assign n5661 = ~pi428 & n5655;
  assign n5662 = ~pi428 & ~n5655;
  assign n5663 = pi428 & n5278;
  assign n5664 = ~n5662 & ~n5663;
  assign n5665 = ~n5660 & ~n5661;
  assign n5666 = ~pi427 & ~n59085;
  assign n5667 = ~n5659 & ~n5666;
  assign n5668 = ~pi430 & n5667;
  assign n5669 = ~pi427 & ~n5658;
  assign n5670 = pi427 & ~n59085;
  assign n5671 = ~n5669 & ~n5670;
  assign n5672 = pi430 & n5671;
  assign n5673 = n59020 & ~n5672;
  assign n5674 = ~n5668 & n5673;
  assign n5675 = ~pi430 & n5671;
  assign n5676 = pi430 & n5667;
  assign n5677 = ~n59020 & ~n5676;
  assign n5678 = ~n5675 & n5677;
  assign n5679 = pi1199 & ~n5678;
  assign n5680 = pi430 & ~n5667;
  assign n5681 = ~pi430 & ~n5671;
  assign n5682 = ~n5680 & ~n5681;
  assign n5683 = pi426 & ~n5682;
  assign n5684 = pi430 & ~n5671;
  assign n5685 = ~pi430 & ~n5667;
  assign n5686 = ~n5684 & ~n5685;
  assign n5687 = ~pi426 & ~n5686;
  assign n5688 = ~n5683 & ~n5687;
  assign n5689 = pi445 & ~n5688;
  assign n5690 = pi426 & ~n5686;
  assign n5691 = ~pi426 & ~n5682;
  assign n5692 = ~n5690 & ~n5691;
  assign n5693 = ~pi445 & ~n5692;
  assign n5694 = ~n5689 & ~n5693;
  assign n5695 = pi448 & n5694;
  assign n5696 = pi445 & ~n5692;
  assign n5697 = ~pi445 & ~n5688;
  assign n5698 = ~n5696 & ~n5697;
  assign n5699 = ~pi448 & n5698;
  assign n5700 = n4455 & ~n5699;
  assign n5701 = ~n5695 & n5700;
  assign n5702 = pi448 & n5698;
  assign n5703 = ~pi448 & n5694;
  assign n5704 = ~n4455 & ~n5703;
  assign n5705 = ~n4455 & ~n5702;
  assign n5706 = ~n5703 & n5705;
  assign n5707 = ~n5702 & n5704;
  assign n5708 = pi1199 & ~n59086;
  assign n5709 = ~n5701 & n5708;
  assign n5710 = pi1199 & ~n5701;
  assign n5711 = ~n59086 & n5710;
  assign n5712 = ~n5674 & n5679;
  assign n5713 = ~pi1199 & n5655;
  assign n5714 = n4677 & ~n5713;
  assign n5715 = ~n59087 & n5714;
  assign n5716 = n5599 & ~n5715;
  assign n5717 = ~n3213 & ~n5716;
  assign n5718 = ~n3213 & ~n59079;
  assign n5719 = ~n5716 & n5718;
  assign n5720 = ~n59079 & n5717;
  assign n5721 = ~n2439 & n5149;
  assign n5722 = pi75 & n5147;
  assign n5723 = n2672 & ~n5306;
  assign n5724 = n5177 & n5723;
  assign n5725 = n58854 & ~n5306;
  assign n5726 = n5160 & n5725;
  assign n5727 = ~n58815 & n5147;
  assign n5728 = ~n5726 & ~n5727;
  assign n5729 = ~n5724 & n5728;
  assign n5730 = ~pi75 & ~n5729;
  assign n5731 = ~n5722 & ~n5730;
  assign n5732 = pi567 & ~n5731;
  assign n5733 = n5315 & ~n5732;
  assign n5734 = ~n5721 & ~n5733;
  assign n5735 = ~pi592 & n5734;
  assign n5736 = ~n5276 & ~n5735;
  assign n5737 = ~n4581 & n5736;
  assign n5738 = pi443 & ~n5736;
  assign n5739 = ~n5606 & ~n5738;
  assign n5740 = n59009 & n5739;
  assign n5741 = ~pi443 & ~n5736;
  assign n5742 = ~n5602 & ~n5741;
  assign n5743 = ~n59009 & n5742;
  assign n5744 = ~n5740 & ~n5743;
  assign n5745 = n59007 & ~n5744;
  assign n5746 = n59009 & n5742;
  assign n5747 = ~n59009 & n5739;
  assign n5748 = ~pi444 & n5742;
  assign n5749 = pi444 & n5739;
  assign n5750 = ~pi436 & ~n5749;
  assign n5751 = ~pi436 & ~n5748;
  assign n5752 = ~n5749 & n5751;
  assign n5753 = ~n5748 & n5750;
  assign n5754 = ~pi444 & n5739;
  assign n5755 = pi444 & n5742;
  assign n5756 = pi436 & ~n5755;
  assign n5757 = pi436 & ~n5754;
  assign n5758 = ~n5755 & n5757;
  assign n5759 = ~n5754 & n5756;
  assign n5760 = ~n59089 & ~n59090;
  assign n5761 = ~n5746 & ~n5747;
  assign n5762 = ~n59007 & n59091;
  assign n5763 = n59005 & ~n5762;
  assign n5764 = ~n5745 & n5763;
  assign n5765 = ~n59007 & ~n5744;
  assign n5766 = n59007 & n59091;
  assign n5767 = ~n59005 & ~n5766;
  assign n5768 = ~n5765 & n5767;
  assign n5769 = ~n5764 & ~n5768;
  assign n5770 = ~pi435 & ~n5744;
  assign n5771 = pi435 & n59091;
  assign n5772 = ~n5770 & ~n5771;
  assign n5773 = ~pi429 & n5772;
  assign n5774 = pi435 & ~n5744;
  assign n5775 = ~pi435 & n59091;
  assign n5776 = ~n5774 & ~n5775;
  assign n5777 = pi429 & n5776;
  assign n5778 = ~n59007 & ~n5777;
  assign n5779 = ~n59007 & ~n5773;
  assign n5780 = ~n5777 & n5779;
  assign n5781 = ~n5773 & n5778;
  assign n5782 = ~pi429 & n5776;
  assign n5783 = pi429 & n5772;
  assign n5784 = n59007 & ~n5783;
  assign n5785 = n59007 & ~n5782;
  assign n5786 = ~n5783 & n5785;
  assign n5787 = ~n5782 & n5784;
  assign n5788 = pi1196 & ~n59093;
  assign n5789 = ~n59092 & n5788;
  assign n5790 = pi1196 & ~n59092;
  assign n5791 = ~n59093 & n5790;
  assign n5792 = pi1196 & ~n5769;
  assign n5793 = n5601 & ~n59094;
  assign n5794 = ~n5737 & ~n5793;
  assign n5795 = pi428 & ~n5794;
  assign n5796 = ~pi428 & n5736;
  assign n5797 = ~n5795 & ~n5796;
  assign n5798 = pi427 & ~n5797;
  assign n5799 = pi428 & ~n5736;
  assign n5800 = ~pi428 & n5794;
  assign n5801 = ~pi428 & ~n5794;
  assign n5802 = pi428 & n5736;
  assign n5803 = ~n5801 & ~n5802;
  assign n5804 = ~n5799 & ~n5800;
  assign n5805 = ~pi427 & ~n59095;
  assign n5806 = ~n5798 & ~n5805;
  assign n5807 = pi430 & n5806;
  assign n5808 = ~pi427 & ~n5797;
  assign n5809 = pi427 & ~n59095;
  assign n5810 = ~n5808 & ~n5809;
  assign n5811 = ~pi430 & n5810;
  assign n5812 = ~n59020 & ~n5811;
  assign n5813 = ~n5807 & n5812;
  assign n5814 = ~pi430 & n5806;
  assign n5815 = pi430 & n5810;
  assign n5816 = n59020 & ~n5815;
  assign n5817 = ~n5814 & n5816;
  assign n5818 = pi1199 & ~n5817;
  assign n5819 = pi430 & ~n5810;
  assign n5820 = ~pi430 & ~n5806;
  assign n5821 = ~n5819 & ~n5820;
  assign n5822 = pi426 & ~n5821;
  assign n5823 = pi430 & ~n5806;
  assign n5824 = ~pi430 & ~n5810;
  assign n5825 = ~n5823 & ~n5824;
  assign n5826 = ~pi426 & ~n5825;
  assign n5827 = ~n5822 & ~n5826;
  assign n5828 = pi445 & ~n5827;
  assign n5829 = pi426 & ~n5825;
  assign n5830 = ~pi426 & ~n5821;
  assign n5831 = ~n5829 & ~n5830;
  assign n5832 = ~pi445 & ~n5831;
  assign n5833 = ~n5828 & ~n5832;
  assign n5834 = pi448 & n5833;
  assign n5835 = pi445 & ~n5831;
  assign n5836 = ~pi445 & ~n5827;
  assign n5837 = ~n5835 & ~n5836;
  assign n5838 = ~pi448 & n5837;
  assign n5839 = ~n4455 & ~n5838;
  assign n5840 = ~n4455 & ~n5834;
  assign n5841 = ~n5838 & n5840;
  assign n5842 = ~n5834 & n5839;
  assign n5843 = pi448 & n5837;
  assign n5844 = ~pi448 & n5833;
  assign n5845 = n4455 & ~n5844;
  assign n5846 = n4455 & ~n5843;
  assign n5847 = ~n5844 & n5846;
  assign n5848 = ~n5843 & n5845;
  assign n5849 = pi1199 & ~n59097;
  assign n5850 = ~n59096 & n5849;
  assign n5851 = ~n5813 & n5818;
  assign n5852 = ~pi1199 & n5794;
  assign n5853 = n4677 & ~n5852;
  assign n5854 = ~n59098 & n5853;
  assign n5855 = n5599 & ~n5854;
  assign n5856 = ~n4860 & n5736;
  assign n5857 = ~n5495 & ~n5856;
  assign n5858 = pi1198 & ~n5857;
  assign n5859 = ~n58853 & n5736;
  assign n5860 = ~n5500 & ~n5859;
  assign n5861 = pi355 & ~n5860;
  assign n5862 = ~pi455 & ~n5736;
  assign n5863 = ~n5504 & ~n5862;
  assign n5864 = ~pi452 & ~n5863;
  assign n5865 = pi455 & ~n5736;
  assign n5866 = ~n5508 & ~n5865;
  assign n5867 = pi452 & ~n5866;
  assign n5868 = ~n5864 & ~n5867;
  assign n5869 = ~pi355 & n5868;
  assign n5870 = ~n5861 & ~n5869;
  assign n5871 = ~pi458 & n5870;
  assign n5872 = ~pi355 & ~n5860;
  assign n5873 = pi355 & n5868;
  assign n5874 = ~n5872 & ~n5873;
  assign n5875 = pi458 & n5874;
  assign n5876 = ~n2965 & ~n5875;
  assign n5877 = ~n2965 & ~n5871;
  assign n5878 = ~n5875 & n5877;
  assign n5879 = ~n5871 & n5876;
  assign n5880 = pi458 & n5870;
  assign n5881 = ~pi458 & n5874;
  assign n5882 = n2965 & ~n5881;
  assign n5883 = ~n5880 & n5882;
  assign n5884 = pi1196 & ~n5883;
  assign n5885 = pi1196 & ~n59099;
  assign n5886 = ~n5883 & n5885;
  assign n5887 = ~n59099 & n5884;
  assign n5888 = n5499 & ~n59100;
  assign n5889 = ~n5858 & ~n5888;
  assign n5890 = ~n3039 & ~n5889;
  assign n5891 = n3039 & n5736;
  assign n5892 = ~n5890 & ~n5891;
  assign n5893 = ~n2437 & n5892;
  assign n5894 = pi1199 & ~n5736;
  assign n5895 = pi351 & n5894;
  assign n5896 = ~n4880 & ~n5895;
  assign n5897 = ~n5893 & n5896;
  assign n5898 = ~n3152 & n5892;
  assign n5899 = ~pi351 & n5894;
  assign n5900 = n4880 & ~n5899;
  assign n5901 = ~n5898 & n5900;
  assign n5902 = ~pi591 & ~n5901;
  assign n5903 = ~n5893 & ~n5895;
  assign n5904 = ~pi461 & ~n5903;
  assign n5905 = ~n5898 & ~n5899;
  assign n5906 = pi461 & ~n5905;
  assign n5907 = ~n5904 & ~n5906;
  assign n5908 = pi357 & n5907;
  assign n5909 = ~pi461 & ~n5905;
  assign n5910 = pi461 & ~n5903;
  assign n5911 = ~n5909 & ~n5910;
  assign n5912 = ~pi357 & n5911;
  assign n5913 = ~pi356 & ~n5912;
  assign n5914 = ~pi357 & ~n5911;
  assign n5915 = pi357 & ~n5907;
  assign n5916 = ~n5914 & ~n5915;
  assign n5917 = ~pi356 & ~n5916;
  assign n5918 = ~n5908 & n5913;
  assign n5919 = pi357 & n5911;
  assign n5920 = ~pi357 & n5907;
  assign n5921 = pi356 & ~n5920;
  assign n5922 = ~pi357 & ~n5907;
  assign n5923 = pi357 & ~n5911;
  assign n5924 = ~n5922 & ~n5923;
  assign n5925 = pi356 & ~n5924;
  assign n5926 = ~n5919 & n5921;
  assign n5927 = ~n59101 & ~n59102;
  assign n5928 = ~pi354 & ~n5927;
  assign n5929 = n59028 & n5907;
  assign n5930 = ~n59028 & n5911;
  assign n5931 = ~pi356 & ~n5924;
  assign n5932 = pi356 & ~n5916;
  assign n5933 = ~n5931 & ~n5932;
  assign n5934 = ~n5929 & ~n5930;
  assign n5935 = pi354 & ~n59103;
  assign n5936 = n58877 & ~n5935;
  assign n5937 = n58877 & ~n5928;
  assign n5938 = ~n5935 & n5937;
  assign n5939 = ~n5928 & n5936;
  assign n5940 = pi354 & ~n5927;
  assign n5941 = ~pi354 & ~n59103;
  assign n5942 = ~n58877 & ~n5941;
  assign n5943 = ~n5940 & n5942;
  assign n5944 = ~pi591 & ~n5943;
  assign n5945 = ~n59104 & n5944;
  assign n5946 = ~n5897 & n5902;
  assign n5947 = n5494 & ~n59105;
  assign n5948 = n3450 & ~n5736;
  assign n5949 = ~n5276 & ~n5380;
  assign n5950 = ~pi1199 & n5949;
  assign n5951 = ~n5276 & n5381;
  assign n5952 = n4280 & ~n5721;
  assign n5953 = n59059 & n5723;
  assign n5954 = n59061 & n5725;
  assign n5955 = ~n5727 & ~n5954;
  assign n5956 = ~n5953 & n5955;
  assign n5957 = ~pi75 & ~n5956;
  assign n5958 = ~n5722 & ~n5957;
  assign n5959 = pi567 & ~n5958;
  assign n5960 = n5315 & ~n5959;
  assign n5961 = n5952 & ~n5960;
  assign n5962 = n59106 & ~n5961;
  assign n5963 = ~n5321 & n5724;
  assign n5964 = n58894 & n5726;
  assign n5965 = ~n5963 & ~n5964;
  assign n5966 = n5956 & n5965;
  assign n5967 = n5952 & ~n5966;
  assign n5968 = ~n5368 & n5726;
  assign n5969 = ~n5727 & ~n5968;
  assign n5970 = ~n5963 & n5969;
  assign n5971 = n4288 & ~n5721;
  assign n5972 = ~n5970 & n5971;
  assign n5973 = ~n5967 & ~n5972;
  assign n5974 = ~pi75 & pi567;
  assign n5975 = ~n5973 & n5974;
  assign n5976 = n3215 & n5315;
  assign n5977 = ~n5149 & ~n5976;
  assign n5978 = pi1199 & ~n5977;
  assign n5979 = ~n5975 & n5978;
  assign n5980 = ~n3450 & ~n5979;
  assign n5981 = ~n5962 & n5980;
  assign n5982 = ~n5948 & ~n5981;
  assign n5983 = pi333 & ~pi391;
  assign n5984 = ~pi333 & pi391;
  assign n5985 = ~n5983 & ~n5984;
  assign n5986 = n5982 & n5985;
  assign n5987 = ~n5424 & ~n5736;
  assign n5988 = ~pi1197 & n5981;
  assign n5989 = ~n5987 & ~n5988;
  assign n5990 = ~n5985 & n5989;
  assign n5991 = pi333 & ~n5989;
  assign n5992 = ~pi333 & ~n5982;
  assign n5993 = ~n5991 & ~n5992;
  assign n5994 = ~pi391 & ~n5993;
  assign n5995 = ~pi333 & ~n5989;
  assign n5996 = pi333 & ~n5982;
  assign n5997 = ~n5995 & ~n5996;
  assign n5998 = pi391 & ~n5997;
  assign n5999 = ~n5994 & ~n5998;
  assign n6000 = ~n5986 & ~n5990;
  assign n6001 = pi392 & n59107;
  assign n6002 = ~n5982 & ~n5985;
  assign n6003 = n5985 & ~n5989;
  assign n6004 = ~pi391 & ~n5997;
  assign n6005 = pi391 & ~n5993;
  assign n6006 = ~n6004 & ~n6005;
  assign n6007 = ~n6002 & ~n6003;
  assign n6008 = ~pi392 & n59108;
  assign n6009 = ~n58988 & ~n6008;
  assign n6010 = ~n6001 & n6009;
  assign n6011 = pi392 & n59108;
  assign n6012 = ~pi392 & n59107;
  assign n6013 = n58988 & ~n6012;
  assign n6014 = ~n6011 & n6013;
  assign n6015 = ~n6010 & ~n6014;
  assign n6016 = ~pi392 & ~n59108;
  assign n6017 = pi392 & ~n59107;
  assign n6018 = ~n6016 & ~n6017;
  assign n6019 = pi393 & ~n6018;
  assign n6020 = ~pi392 & ~n59107;
  assign n6021 = pi392 & ~n59108;
  assign n6022 = ~n6020 & ~n6021;
  assign n6023 = ~pi393 & ~n6022;
  assign n6024 = n58905 & ~n6023;
  assign n6025 = ~n6019 & n6024;
  assign n6026 = ~pi393 & ~n6018;
  assign n6027 = pi393 & ~n6022;
  assign n6028 = ~n58905 & ~n6027;
  assign n6029 = ~n58905 & ~n6026;
  assign n6030 = ~n6027 & n6029;
  assign n6031 = ~n6026 & n6028;
  assign n6032 = pi591 & ~n59109;
  assign n6033 = ~n6025 & n6032;
  assign n6034 = pi591 & ~n6025;
  assign n6035 = ~n59109 & n6034;
  assign n6036 = pi591 & ~n6015;
  assign n6037 = n3703 & ~n5149;
  assign n6038 = pi592 & n5734;
  assign n6039 = ~n5150 & ~n6038;
  assign n6040 = ~n3703 & ~n6039;
  assign n6041 = n58918 & n6039;
  assign n6042 = ~n58918 & n5149;
  assign n6043 = pi1197 & ~n6042;
  assign n6044 = ~n6041 & n6043;
  assign n6045 = n5235 & ~n6044;
  assign n6046 = n58911 & n6039;
  assign n6047 = ~pi1199 & ~n6046;
  assign n6048 = ~n6045 & n6047;
  assign n6049 = ~n4893 & n6039;
  assign n6050 = n5242 & ~n6049;
  assign n6051 = ~n6048 & ~n6050;
  assign n6052 = ~n6037 & ~n6040;
  assign n6053 = n59029 & n59111;
  assign n6054 = pi1198 & ~n6039;
  assign n6055 = ~n59029 & ~n6054;
  assign n6056 = n58928 & ~n6055;
  assign n6057 = ~n6053 & n6056;
  assign n6058 = n59029 & ~n6054;
  assign n6059 = ~n58928 & ~n6058;
  assign n6060 = n59029 & n6059;
  assign n6061 = n59111 & ~n6060;
  assign n6062 = pi1198 & ~n6059;
  assign n6063 = ~n6061 & ~n6062;
  assign n6064 = ~n6057 & ~n6063;
  assign n6065 = ~pi1198 & ~n59111;
  assign n6066 = ~n6054 & ~n6065;
  assign n6067 = ~pi374 & ~n6066;
  assign n6068 = pi374 & ~n59111;
  assign n6069 = ~n6067 & ~n6068;
  assign n6070 = ~pi369 & ~n6069;
  assign n6071 = ~pi374 & ~n59111;
  assign n6072 = pi374 & ~n6066;
  assign n6073 = ~n6071 & ~n6072;
  assign n6074 = pi369 & ~n6073;
  assign n6075 = n59029 & ~n6074;
  assign n6076 = ~n6070 & n6075;
  assign n6077 = pi369 & ~n6069;
  assign n6078 = ~pi369 & ~n6073;
  assign n6079 = ~n59029 & ~n6078;
  assign n6080 = ~n6077 & n6079;
  assign n6081 = ~pi591 & ~n6080;
  assign n6082 = ~n6076 & n6081;
  assign n6083 = ~pi591 & ~n6076;
  assign n6084 = ~n6080 & n6083;
  assign n6085 = ~pi591 & ~n6064;
  assign n6086 = ~pi590 & ~n59112;
  assign n6087 = ~n59110 & n6086;
  assign n6088 = ~pi588 & ~n6087;
  assign n6089 = ~n5947 & n6088;
  assign n6090 = n3213 & ~n6089;
  assign n6091 = ~n5855 & n6090;
  assign n6092 = ~pi80 & n58992;
  assign n6093 = ~n6091 & n6092;
  assign n6094 = ~n59088 & n6092;
  assign n6095 = ~n6091 & n6094;
  assign n6096 = ~n59088 & n6093;
  assign n6097 = ~n4858 & n5149;
  assign n6098 = ~n4881 & n5149;
  assign n6099 = n4865 & n6098;
  assign n6100 = ~n2437 & n6099;
  assign n6101 = ~n6097 & ~n6100;
  assign n6102 = pi461 & ~n6101;
  assign n6103 = ~n3152 & n6099;
  assign n6104 = ~n6097 & ~n6103;
  assign n6105 = ~pi461 & ~n6104;
  assign n6106 = ~n6102 & ~n6105;
  assign n6107 = n59028 & n6106;
  assign n6108 = pi461 & ~n6104;
  assign n6109 = ~pi461 & ~n6101;
  assign n6110 = ~n6108 & ~n6109;
  assign n6111 = ~n59028 & n6110;
  assign n6112 = pi357 & ~n6106;
  assign n6113 = ~pi357 & ~n6110;
  assign n6114 = ~n6112 & ~n6113;
  assign n6115 = pi356 & ~n6114;
  assign n6116 = pi357 & ~n6110;
  assign n6117 = ~pi357 & ~n6106;
  assign n6118 = ~n6116 & ~n6117;
  assign n6119 = ~pi356 & ~n6118;
  assign n6120 = ~n6115 & ~n6119;
  assign n6121 = ~n6107 & ~n6111;
  assign n6122 = pi354 & n59114;
  assign n6123 = ~n59028 & ~n6106;
  assign n6124 = n59028 & ~n6110;
  assign n6125 = pi357 & n6110;
  assign n6126 = ~pi357 & n6106;
  assign n6127 = pi356 & ~n6126;
  assign n6128 = pi356 & ~n6118;
  assign n6129 = ~n6125 & n6127;
  assign n6130 = pi357 & n6106;
  assign n6131 = ~pi357 & n6110;
  assign n6132 = ~pi356 & ~n6131;
  assign n6133 = ~pi356 & ~n6114;
  assign n6134 = ~n6130 & n6132;
  assign n6135 = ~n59115 & ~n59116;
  assign n6136 = ~n6123 & ~n6124;
  assign n6137 = ~pi354 & n59117;
  assign n6138 = ~n58877 & ~n6137;
  assign n6139 = ~n58877 & ~n6122;
  assign n6140 = ~n6137 & n6139;
  assign n6141 = ~n6122 & n6138;
  assign n6142 = ~pi354 & n59114;
  assign n6143 = pi354 & n59117;
  assign n6144 = n58877 & ~n6143;
  assign n6145 = n58877 & ~n6142;
  assign n6146 = ~n6143 & n6145;
  assign n6147 = ~n6142 & n6144;
  assign n6148 = ~pi591 & ~n59119;
  assign n6149 = ~pi591 & ~n59118;
  assign n6150 = ~n59119 & n6149;
  assign n6151 = ~n59118 & n6148;
  assign n6152 = n5494 & ~n59120;
  assign n6153 = ~pi1196 & n5313;
  assign n6154 = ~pi592 & ~n6153;
  assign n6155 = ~n5314 & n6154;
  assign n6156 = pi1199 & ~n5276;
  assign n6157 = ~n6155 & n6156;
  assign n6158 = n4280 & ~n5382;
  assign n6159 = n59106 & ~n6158;
  assign n6160 = n4991 & ~n6159;
  assign n6161 = ~n6157 & n6160;
  assign n6162 = ~n4991 & ~n6097;
  assign n6163 = pi591 & ~n6162;
  assign n6164 = ~n6161 & n6163;
  assign n6165 = n3954 & ~n4897;
  assign n6166 = ~pi1198 & ~n6165;
  assign n6167 = ~n4915 & ~n5011;
  assign n6168 = ~n5011 & ~n6166;
  assign n6169 = ~n4915 & n6168;
  assign n6170 = ~n6166 & n6167;
  assign n6171 = ~pi591 & n5149;
  assign n6172 = ~n59121 & n6171;
  assign n6173 = ~n6164 & ~n6172;
  assign n6174 = ~n5424 & ~n6097;
  assign n6175 = n5949 & ~n6158;
  assign n6176 = ~pi1199 & ~n6175;
  assign n6177 = n4280 & ~n5314;
  assign n6178 = n4288 & ~n5313;
  assign n6179 = ~n5276 & ~n6178;
  assign n6180 = ~n6177 & n6179;
  assign n6181 = pi1199 & ~n6180;
  assign n6182 = ~n6176 & ~n6181;
  assign n6183 = n5424 & ~n6182;
  assign n6184 = ~n6174 & ~n6183;
  assign n6185 = ~pi333 & ~n6184;
  assign n6186 = n3450 & ~n6097;
  assign n6187 = ~n3450 & ~n6182;
  assign n6188 = ~n6186 & ~n6187;
  assign n6189 = pi333 & ~n6188;
  assign n6190 = ~n6185 & ~n6189;
  assign n6191 = ~pi391 & ~n6190;
  assign n6192 = pi333 & ~n6184;
  assign n6193 = ~pi333 & ~n6188;
  assign n6194 = ~n6192 & ~n6193;
  assign n6195 = pi391 & ~n6194;
  assign n6196 = ~n4983 & ~n6195;
  assign n6197 = ~n6191 & n6196;
  assign n6198 = ~pi391 & ~n6194;
  assign n6199 = pi391 & ~n6190;
  assign n6200 = n4983 & ~n6199;
  assign n6201 = ~n6198 & n6200;
  assign n6202 = pi591 & ~n6201;
  assign n6203 = pi591 & ~n6197;
  assign n6204 = ~n6201 & n6203;
  assign n6205 = ~n6197 & n6202;
  assign n6206 = n5149 & ~n59121;
  assign n6207 = ~pi591 & ~n6206;
  assign n6208 = ~pi590 & ~n6207;
  assign n6209 = ~n59122 & n6208;
  assign n6210 = ~pi590 & ~n6173;
  assign n6211 = ~pi588 & ~n59123;
  assign n6212 = ~pi588 & ~n6152;
  assign n6213 = ~n59123 & n6212;
  assign n6214 = ~n6152 & n6211;
  assign n6215 = ~n59012 & ~n6097;
  assign n6216 = pi592 & ~n4581;
  assign n6217 = n3954 & ~n5069;
  assign n6218 = ~n6216 & n6217;
  assign n6219 = n5149 & ~n6218;
  assign n6220 = n59012 & ~n6219;
  assign n6221 = pi428 & ~n6219;
  assign n6222 = ~pi428 & ~n6097;
  assign n6223 = ~n6221 & ~n6222;
  assign n6224 = ~pi427 & ~n6223;
  assign n6225 = ~pi428 & ~n6219;
  assign n6226 = pi428 & ~n6097;
  assign n6227 = ~n6225 & ~n6226;
  assign n6228 = pi427 & ~n6227;
  assign n6229 = ~n6224 & ~n6228;
  assign n6230 = ~n6215 & ~n6220;
  assign n6231 = ~pi430 & n59125;
  assign n6232 = ~n59012 & n6219;
  assign n6233 = n59012 & n6097;
  assign n6234 = ~pi428 & n6219;
  assign n6235 = pi428 & n6097;
  assign n6236 = ~pi427 & ~n6235;
  assign n6237 = ~pi427 & ~n6227;
  assign n6238 = ~n6234 & n6236;
  assign n6239 = pi428 & n6219;
  assign n6240 = ~pi428 & n6097;
  assign n6241 = pi427 & ~n6240;
  assign n6242 = pi427 & ~n6223;
  assign n6243 = ~n6239 & n6241;
  assign n6244 = ~n59126 & ~n59127;
  assign n6245 = ~n6232 & ~n6233;
  assign n6246 = pi430 & n59128;
  assign n6247 = pi430 & ~n59128;
  assign n6248 = ~pi430 & ~n59125;
  assign n6249 = ~n6247 & ~n6248;
  assign n6250 = ~n6231 & ~n6246;
  assign n6251 = pi426 & n59129;
  assign n6252 = ~pi430 & ~n59128;
  assign n6253 = pi430 & ~n59125;
  assign n6254 = ~pi426 & ~n6253;
  assign n6255 = ~n6252 & n6254;
  assign n6256 = ~n58996 & ~n6255;
  assign n6257 = ~n6251 & n6256;
  assign n6258 = n4446 & n59125;
  assign n6259 = ~n4446 & n59128;
  assign n6260 = n58996 & ~n6259;
  assign n6261 = ~n6258 & n6260;
  assign n6262 = ~n6257 & ~n6261;
  assign n6263 = ~n6252 & ~n6253;
  assign n6264 = ~pi426 & ~n6263;
  assign n6265 = pi426 & ~n59129;
  assign n6266 = ~n6264 & ~n6265;
  assign n6267 = ~pi445 & ~n6266;
  assign n6268 = ~pi426 & ~n59129;
  assign n6269 = pi426 & ~n6263;
  assign n6270 = ~n6268 & ~n6269;
  assign n6271 = pi445 & ~n6270;
  assign n6272 = ~n6267 & ~n6271;
  assign n6273 = pi448 & ~n6272;
  assign n6274 = ~pi445 & ~n6270;
  assign n6275 = pi445 & ~n6266;
  assign n6276 = ~n6274 & ~n6275;
  assign n6277 = ~pi448 & ~n6276;
  assign n6278 = ~n4455 & ~n6277;
  assign n6279 = ~n6273 & n6278;
  assign n6280 = pi448 & ~n6276;
  assign n6281 = ~pi448 & ~n6272;
  assign n6282 = n4455 & ~n6281;
  assign n6283 = n4455 & ~n6280;
  assign n6284 = ~n6281 & n6283;
  assign n6285 = ~n6280 & n6282;
  assign n6286 = pi1199 & ~n59130;
  assign n6287 = ~n6279 & n6286;
  assign n6288 = pi1199 & ~n6262;
  assign n6289 = ~pi1199 & ~n6219;
  assign n6290 = n4677 & ~n6289;
  assign n6291 = ~n59131 & n6290;
  assign n6292 = n5599 & ~n6291;
  assign n6293 = ~n3213 & ~n6292;
  assign n6294 = ~n59124 & n6293;
  assign n6295 = n3213 & n5149;
  assign n6296 = ~pi80 & ~n58992;
  assign n6297 = ~n6295 & n6296;
  assign n6298 = ~n6294 & n6297;
  assign n6299 = ~pi217 & ~n6298;
  assign n6300 = ~n59113 & n6299;
  assign n6301 = ~pi80 & ~n5149;
  assign n6302 = pi217 & ~n6301;
  assign n6303 = n5138 & ~n6302;
  assign po238 = ~n6300 & n6303;
  assign n6305 = ~pi87 & ~pi100;
  assign n6306 = ~pi54 & ~pi74;
  assign n6307 = ~pi75 & ~pi92;
  assign n6308 = n6306 & n6307;
  assign n6309 = ~pi75 & ~pi87;
  assign n6310 = ~pi92 & n6309;
  assign n6311 = n6306 & n6310;
  assign n6312 = ~pi100 & n6311;
  assign n6313 = n6305 & n6308;
  assign n6314 = pi140 & ~n59132;
  assign n6315 = pi40 & ~n58824;
  assign n6316 = n2598 & ~n6315;
  assign n6317 = n2471 & n5151;
  assign n6318 = ~pi66 & ~pi84;
  assign n6319 = n2475 & n6318;
  assign n6320 = ~pi36 & ~pi67;
  assign n6321 = ~pi103 & n6320;
  assign n6322 = n6319 & n6321;
  assign n6323 = ~pi68 & ~pi73;
  assign n6324 = ~pi69 & ~pi83;
  assign n6325 = n2478 & n6324;
  assign n6326 = n6323 & n6325;
  assign n6327 = n6322 & n6326;
  assign n6328 = pi45 & n2446;
  assign n6329 = pi45 & n2457;
  assign n6330 = n2446 & n6329;
  assign n6331 = n2457 & n6328;
  assign n6332 = n6327 & n59133;
  assign n6333 = n2454 & n6332;
  assign n6334 = ~pi102 & ~n6333;
  assign n6335 = pi102 & ~n2521;
  assign n6336 = ~pi98 & ~n6335;
  assign n6337 = ~n6334 & n6336;
  assign n6338 = n6317 & n6337;
  assign n6339 = ~pi94 & n58798;
  assign n6340 = n58789 & n2531;
  assign n6341 = ~pi96 & n2581;
  assign n6342 = n2580 & n2641;
  assign n6343 = ~pi35 & ~pi51;
  assign n6344 = ~pi96 & n2614;
  assign n6345 = n2641 & n6343;
  assign n6346 = ~pi72 & ~pi93;
  assign n6347 = n59136 & n6346;
  assign n6348 = ~pi93 & n58823;
  assign n6349 = n2592 & n58817;
  assign n6350 = ~pi90 & n59137;
  assign n6351 = n2579 & n58823;
  assign n6352 = n2642 & n59135;
  assign n6353 = n59134 & n59138;
  assign n6354 = n6338 & n6353;
  assign n6355 = ~pi40 & ~n6354;
  assign n6356 = n6316 & ~n6355;
  assign n6357 = ~pi252 & ~n6356;
  assign n6358 = pi47 & n58794;
  assign n6359 = n58791 & n6358;
  assign n6360 = pi47 & ~n6359;
  assign n6361 = ~pi91 & ~n6360;
  assign n6362 = n2530 & ~n6360;
  assign n6363 = n2579 & n6362;
  assign n6364 = n2589 & n6361;
  assign n6365 = ~pi97 & n58833;
  assign n6366 = ~pi46 & pi108;
  assign n6367 = pi108 & n2491;
  assign n6368 = n2490 & n6366;
  assign n6369 = n6365 & n59140;
  assign n6370 = pi314 & n6369;
  assign n6371 = n58789 & n6338;
  assign n6372 = ~pi47 & ~n6371;
  assign n6373 = ~n6370 & n6372;
  assign n6374 = n59139 & ~n6373;
  assign n6375 = ~pi35 & ~n6374;
  assign n6376 = pi35 & ~n2615;
  assign n6377 = n58817 & ~n6376;
  assign n6378 = ~pi40 & n6377;
  assign n6379 = ~n6375 & n6378;
  assign n6380 = pi40 & n58824;
  assign n6381 = pi252 & ~n6380;
  assign n6382 = ~n6379 & n6381;
  assign n6383 = ~n6357 & ~n6382;
  assign n6384 = n2598 & n6383;
  assign n6385 = pi1092 & ~n2872;
  assign n6386 = pi1092 & n6384;
  assign n6387 = ~n2872 & n6386;
  assign n6388 = n6384 & n6385;
  assign n6389 = ~pi98 & n2559;
  assign n6390 = pi88 & ~n6389;
  assign n6391 = n2471 & ~n6390;
  assign n6392 = ~pi88 & ~n6337;
  assign n6393 = n6391 & ~n6392;
  assign n6394 = n58791 & n6393;
  assign n6395 = ~pi47 & ~n6394;
  assign n6396 = ~pi47 & ~n6370;
  assign n6397 = ~n6394 & n6396;
  assign n6398 = ~n6370 & n6395;
  assign n6399 = n59139 & ~n59142;
  assign n6400 = ~pi35 & ~n6399;
  assign n6401 = pi252 & n6377;
  assign n6402 = ~n6400 & n6401;
  assign n6403 = n58797 & n59138;
  assign n6404 = ~pi252 & n6403;
  assign n6405 = n6393 & n6404;
  assign n6406 = ~pi40 & ~n6405;
  assign n6407 = ~n6402 & n6406;
  assign n6408 = n2727 & n6316;
  assign n6409 = ~n6407 & n6408;
  assign n6410 = ~n59141 & ~n6409;
  assign n6411 = pi1093 & ~n6410;
  assign n6412 = ~n2692 & ~n6411;
  assign n6413 = pi1092 & n2797;
  assign n6414 = pi1091 & n2794;
  assign po1106 = n2692 & n59143;
  assign n6416 = n2692 & n2797;
  assign n6417 = n6386 & n6416;
  assign n6418 = n6384 & po1106;
  assign n6419 = ~n2793 & ~n59144;
  assign n6420 = ~n6412 & ~n6419;
  assign n6421 = ~pi1091 & n6411;
  assign n6422 = ~n6420 & ~n6421;
  assign n6423 = ~pi198 & n6422;
  assign n6424 = ~n6315 & ~n6407;
  assign n6425 = ~pi32 & ~n6424;
  assign n6426 = n2601 & n2616;
  assign n6427 = pi32 & ~n6426;
  assign n6428 = ~pi95 & n2441;
  assign n6429 = ~n6427 & n6428;
  assign n6430 = pi824 & n6429;
  assign n6431 = ~n6425 & n6429;
  assign n6432 = pi824 & n6431;
  assign n6433 = ~n6425 & n6430;
  assign n6434 = ~n59141 & ~n59145;
  assign n6435 = n2878 & ~n6434;
  assign n6436 = ~pi32 & ~n6383;
  assign n6437 = ~pi824 & n6429;
  assign n6438 = ~n6436 & n6437;
  assign n6439 = n6429 & ~n6436;
  assign n6440 = ~pi824 & pi829;
  assign n6441 = n6439 & n6440;
  assign n6442 = pi829 & n6438;
  assign n6443 = n6434 & ~n59146;
  assign n6444 = pi1093 & ~n6443;
  assign n6445 = ~n2692 & ~n6444;
  assign n6446 = ~n6419 & ~n6445;
  assign n6447 = ~n6435 & ~n6446;
  assign n6448 = pi198 & n6447;
  assign n6449 = ~n6423 & ~n6448;
  assign n6450 = ~pi299 & n6449;
  assign n6451 = ~pi210 & n6422;
  assign n6452 = pi210 & n6447;
  assign n6453 = ~n6451 & ~n6452;
  assign n6454 = pi299 & n6453;
  assign n6455 = pi299 & ~n6453;
  assign n6456 = ~pi299 & ~n6449;
  assign n6457 = ~n6455 & ~n6456;
  assign n6458 = ~n6450 & ~n6454;
  assign n6459 = ~pi39 & ~n59147;
  assign n6460 = n2801 & ~n2805;
  assign n6461 = ~pi120 & ~n6460;
  assign n6462 = pi120 & ~n58822;
  assign n6463 = ~n6461 & ~n6462;
  assign n6464 = n2794 & n6463;
  assign n6465 = ~n2680 & n6464;
  assign n6466 = n2794 & n6460;
  assign n6467 = ~pi120 & ~n6466;
  assign n6468 = n58822 & n2794;
  assign n6469 = ~pi287 & n2805;
  assign n6470 = pi835 & pi950;
  assign n6471 = n6469 & n6470;
  assign n6472 = ~n2442 & ~n2692;
  assign n6473 = n6471 & n6472;
  assign n6474 = n6468 & ~n6473;
  assign n6475 = pi120 & ~n6474;
  assign n6476 = pi1091 & ~n6475;
  assign n6477 = ~n6467 & n6476;
  assign n6478 = pi120 & ~n6468;
  assign n6479 = ~pi1091 & ~n6478;
  assign n6480 = pi120 & pi824;
  assign n6481 = n6471 & n6480;
  assign n6482 = n6479 & ~n6481;
  assign n6483 = ~n6467 & n6482;
  assign n6484 = ~n6477 & ~n6483;
  assign n6485 = n2680 & ~n6484;
  assign n6486 = ~n6465 & ~n6485;
  assign n6487 = ~n2776 & ~n6464;
  assign n6488 = n2680 & ~n6464;
  assign n6489 = ~n2680 & n6484;
  assign n6490 = ~n6488 & ~n6489;
  assign n6491 = n2776 & ~n6490;
  assign n6492 = ~n6487 & ~n6491;
  assign n6493 = ~pi614 & ~n6492;
  assign n6494 = ~pi616 & n6493;
  assign n6495 = n2777 & ~n6492;
  assign n6496 = ~n6486 & ~n59148;
  assign n6497 = pi681 & ~n6496;
  assign n6498 = pi616 & ~n6464;
  assign n6499 = pi614 & ~n6464;
  assign n6500 = ~n6493 & ~n6499;
  assign n6501 = ~pi616 & ~n6500;
  assign n6502 = ~n6498 & ~n6501;
  assign n6503 = ~n2779 & ~n6502;
  assign n6504 = n2779 & n6484;
  assign n6505 = ~n2680 & ~n6504;
  assign n6506 = ~n6503 & n6505;
  assign n6507 = ~n6485 & ~n6506;
  assign n6508 = ~pi661 & ~n6507;
  assign n6509 = pi661 & n6496;
  assign n6510 = ~pi681 & ~n6509;
  assign n6511 = ~n6508 & n6510;
  assign n6512 = ~n6497 & ~n6511;
  assign n6513 = ~n2790 & n6512;
  assign n6514 = n2781 & n6490;
  assign n6515 = ~n2781 & n6502;
  assign n6516 = pi681 & ~n6502;
  assign n6517 = ~pi661 & ~pi681;
  assign n6518 = ~pi662 & n6517;
  assign n6519 = ~pi616 & ~n6518;
  assign n6520 = n6500 & n6519;
  assign n6521 = ~pi680 & n6501;
  assign n6522 = pi680 & ~n6490;
  assign n6523 = ~pi616 & n6518;
  assign n6524 = ~n6522 & n6523;
  assign n6525 = ~n6521 & n6524;
  assign n6526 = ~n6520 & ~n6525;
  assign n6527 = ~pi680 & ~n6464;
  assign n6528 = pi616 & n6518;
  assign n6529 = ~n6527 & n6528;
  assign n6530 = ~n6522 & n6529;
  assign n6531 = pi616 & n6464;
  assign n6532 = ~n6518 & n6531;
  assign n6533 = ~n6530 & ~n6532;
  assign n6534 = ~pi681 & n6533;
  assign n6535 = n6526 & n6534;
  assign n6536 = ~n6516 & ~n6535;
  assign n6537 = ~n6514 & ~n6515;
  assign n6538 = n2790 & n59149;
  assign n6539 = n2790 & ~n59149;
  assign n6540 = ~n2790 & ~n6512;
  assign n6541 = ~n6539 & ~n6540;
  assign n6542 = ~n6513 & ~n6538;
  assign n6543 = pi223 & ~n59150;
  assign n6544 = ~pi222 & ~pi224;
  assign n6545 = n2692 & n6466;
  assign n6546 = ~pi824 & ~n6460;
  assign n6547 = ~pi824 & n2441;
  assign n6548 = ~pi984 & ~n2441;
  assign n6549 = pi835 & ~n6548;
  assign n6550 = n2804 & ~n6549;
  assign n6551 = n2801 & ~n6550;
  assign n6552 = pi1092 & n6551;
  assign n6553 = ~n6547 & ~n6552;
  assign n6554 = ~n6546 & ~n6553;
  assign n6555 = ~pi829 & ~n6554;
  assign n6556 = pi829 & ~n6552;
  assign n6557 = n2726 & ~n6556;
  assign n6558 = ~n6555 & n6557;
  assign n6559 = ~n6545 & ~n6558;
  assign n6560 = pi1091 & ~n6559;
  assign n6561 = ~pi120 & ~n6560;
  assign n6562 = ~n6478 & ~n6561;
  assign n6563 = pi1093 & n6554;
  assign n6564 = ~pi120 & ~n6563;
  assign n6565 = n6479 & ~n6564;
  assign n6566 = ~n6562 & ~n6565;
  assign n6567 = n2680 & ~n6566;
  assign n6568 = ~n6465 & ~n6567;
  assign n6569 = ~n2778 & n6568;
  assign n6570 = n2778 & n6566;
  assign n6571 = n2778 & ~n6566;
  assign n6572 = ~n2778 & ~n6568;
  assign n6573 = ~n6571 & ~n6572;
  assign n6574 = ~n6569 & ~n6570;
  assign n6575 = ~n2781 & n59151;
  assign n6576 = n2781 & n6566;
  assign n6577 = ~n2780 & ~n59151;
  assign n6578 = n2780 & ~n6566;
  assign n6579 = ~pi681 & ~n6578;
  assign n6580 = ~n6577 & n6579;
  assign n6581 = pi681 & n59151;
  assign n6582 = ~n6580 & ~n6581;
  assign n6583 = ~n6575 & ~n6576;
  assign n6584 = ~n2790 & n59152;
  assign n6585 = ~pi603 & ~n6464;
  assign n6586 = ~n2680 & n6566;
  assign n6587 = ~n6488 & ~n6586;
  assign n6588 = pi603 & ~n6587;
  assign n6589 = ~n6585 & ~n6588;
  assign n6590 = ~pi642 & ~n6589;
  assign n6591 = ~n6487 & ~n6590;
  assign n6592 = ~pi614 & ~n6591;
  assign n6593 = ~n6499 & ~n6592;
  assign n6594 = ~pi616 & ~n6593;
  assign n6595 = ~n6498 & ~n6594;
  assign n6596 = pi681 & ~n6595;
  assign n6597 = ~pi616 & ~n6591;
  assign n6598 = ~pi614 & ~n2781;
  assign n6599 = ~n6498 & n6598;
  assign n6600 = ~n6498 & ~n6597;
  assign n6601 = n6598 & n6600;
  assign n6602 = ~n6597 & n6599;
  assign n6603 = ~pi614 & n2781;
  assign n6604 = n6587 & n6603;
  assign n6605 = ~n59153 & ~n6604;
  assign n6606 = pi680 & ~n6587;
  assign n6607 = pi614 & n6518;
  assign n6608 = ~n6527 & n6607;
  assign n6609 = ~n6606 & n6608;
  assign n6610 = pi614 & n6464;
  assign n6611 = ~n6518 & n6610;
  assign n6612 = ~n6609 & ~n6611;
  assign n6613 = ~pi681 & n6612;
  assign n6614 = n6605 & n6613;
  assign n6615 = ~n6596 & ~n6614;
  assign n6616 = n2790 & n6615;
  assign n6617 = n2790 & ~n6615;
  assign n6618 = ~n2790 & ~n59152;
  assign n6619 = ~n6617 & ~n6618;
  assign n6620 = ~n6584 & ~n6616;
  assign n6621 = ~n6544 & n59154;
  assign n6622 = n6463 & n6544;
  assign n6623 = n6468 & n6622;
  assign n6624 = n6464 & n6544;
  assign n6625 = ~pi223 & ~n59155;
  assign n6626 = ~n6621 & n6625;
  assign n6627 = ~n6543 & ~n6626;
  assign n6628 = ~pi299 & ~n6627;
  assign n6629 = ~pi216 & ~pi221;
  assign n6630 = n2839 & ~n6615;
  assign n6631 = ~n2839 & ~n59152;
  assign n6632 = n2840 & ~n6631;
  assign n6633 = ~n6630 & n6632;
  assign n6634 = ~n6629 & n6633;
  assign n6635 = ~n2840 & n59152;
  assign n6636 = ~n6629 & n6635;
  assign n6637 = n6464 & n6629;
  assign n6638 = ~pi215 & ~n6637;
  assign n6639 = ~n6464 & n6629;
  assign n6640 = ~n6629 & ~n6635;
  assign n6641 = ~n6639 & ~n6640;
  assign n6642 = ~pi215 & ~n6641;
  assign n6643 = ~n6636 & n6638;
  assign n6644 = ~n6634 & n59156;
  assign n6645 = ~n2840 & n6512;
  assign n6646 = ~n2839 & ~n6512;
  assign n6647 = n2839 & ~n59149;
  assign n6648 = n2840 & ~n6647;
  assign n6649 = ~n6646 & n6648;
  assign n6650 = ~n6645 & ~n6649;
  assign n6651 = pi215 & n6650;
  assign n6652 = ~n6644 & ~n6651;
  assign n6653 = pi299 & ~n6652;
  assign n6654 = ~n6628 & ~n6653;
  assign n6655 = pi39 & ~n6654;
  assign n6656 = ~n6459 & ~n6655;
  assign n6657 = pi761 & n6656;
  assign n6658 = pi621 & n6420;
  assign n6659 = ~pi198 & ~n6658;
  assign n6660 = pi621 & n6446;
  assign n6661 = pi198 & ~n6660;
  assign n6662 = ~n6659 & ~n6661;
  assign n6663 = pi621 & ~n6421;
  assign n6664 = ~n6422 & ~n6663;
  assign n6665 = ~pi198 & n6664;
  assign n6666 = pi621 & ~n6435;
  assign n6667 = ~n6447 & ~n6666;
  assign n6668 = pi198 & n6667;
  assign n6669 = ~n6665 & ~n6668;
  assign n6670 = ~pi603 & ~n6669;
  assign n6671 = ~n6662 & ~n6670;
  assign n6672 = ~pi299 & ~n6671;
  assign n6673 = ~pi210 & ~n6658;
  assign n6674 = pi210 & ~n6660;
  assign n6675 = ~n6673 & ~n6674;
  assign n6676 = pi603 & ~n6675;
  assign n6677 = n6453 & ~n6676;
  assign n6678 = pi299 & n6677;
  assign n6679 = pi299 & ~n6677;
  assign n6680 = ~pi299 & n6671;
  assign n6681 = ~n6679 & ~n6680;
  assign n6682 = ~n6672 & ~n6678;
  assign n6683 = ~pi39 & n59157;
  assign n6684 = pi621 & pi1091;
  assign n6685 = n6562 & n6684;
  assign n6686 = pi621 & ~n6565;
  assign n6687 = ~n6566 & ~n6686;
  assign n6688 = ~pi603 & n6687;
  assign n6689 = ~n6685 & ~n6688;
  assign n6690 = n59152 & ~n6689;
  assign n6691 = ~n58846 & n6690;
  assign n6692 = n6464 & n6684;
  assign n6693 = n2680 & ~n6692;
  assign n6694 = ~n2680 & ~n6685;
  assign n6695 = ~n6693 & ~n6694;
  assign n6696 = pi603 & ~n6695;
  assign n6697 = n6587 & ~n6696;
  assign n6698 = n2781 & ~n6697;
  assign n6699 = ~pi614 & ~pi642;
  assign n6700 = ~pi616 & n6699;
  assign n6701 = pi603 & ~n6684;
  assign n6702 = n6464 & ~n6701;
  assign n6703 = ~n6700 & n6702;
  assign n6704 = ~n6585 & n6700;
  assign n6705 = ~n6696 & n6704;
  assign n6706 = ~n6703 & ~n6705;
  assign n6707 = ~n2781 & n6706;
  assign n6708 = ~n6698 & ~n6707;
  assign n6709 = n58846 & n6708;
  assign n6710 = ~n6691 & ~n6709;
  assign n6711 = n58846 & ~n6708;
  assign n6712 = ~n58846 & ~n6690;
  assign n6713 = ~n6629 & ~n6712;
  assign n6714 = ~n6711 & n6713;
  assign n6715 = ~n6629 & ~n6711;
  assign n6716 = ~n6712 & n6715;
  assign n6717 = ~n6629 & ~n6710;
  assign n6718 = n6629 & n6702;
  assign n6719 = ~pi215 & ~n6718;
  assign n6720 = ~n59158 & n6719;
  assign n6721 = pi621 & n6477;
  assign n6722 = ~n2680 & ~n6721;
  assign n6723 = ~n6693 & ~n6722;
  assign n6724 = pi603 & ~n6723;
  assign n6725 = n6514 & ~n6724;
  assign n6726 = n6704 & ~n6724;
  assign n6727 = ~n6703 & ~n6726;
  assign n6728 = ~n2781 & ~n6727;
  assign n6729 = ~n6725 & ~n6728;
  assign n6730 = n58846 & ~n6729;
  assign n6731 = n2794 & ~n6701;
  assign n6732 = ~n6486 & n6731;
  assign n6733 = n2778 & ~n6477;
  assign n6734 = n6732 & ~n6733;
  assign n6735 = ~n2781 & ~n6734;
  assign n6736 = ~n6484 & n6731;
  assign n6737 = pi680 & ~n6736;
  assign n6738 = n6518 & n6737;
  assign n6739 = n2781 & ~n6736;
  assign n6740 = ~n6735 & ~n59159;
  assign n6741 = ~n58846 & n6740;
  assign n6742 = pi215 & ~n6741;
  assign n6743 = ~n6730 & n6742;
  assign n6744 = ~n59158 & ~n6718;
  assign n6745 = ~pi215 & ~n6744;
  assign n6746 = n58846 & n6729;
  assign n6747 = ~n58846 & ~n6740;
  assign n6748 = pi215 & ~n6747;
  assign n6749 = ~n6746 & n6748;
  assign n6750 = ~n6745 & ~n6749;
  assign n6751 = ~n6720 & ~n6743;
  assign n6752 = pi299 & n59160;
  assign n6753 = n2790 & n6708;
  assign n6754 = ~n2790 & n6690;
  assign n6755 = ~n6753 & ~n6754;
  assign n6756 = n2790 & ~n6708;
  assign n6757 = ~n2790 & ~n6690;
  assign n6758 = ~n6544 & ~n6757;
  assign n6759 = ~n6756 & n6758;
  assign n6760 = ~n6544 & ~n6756;
  assign n6761 = ~n6757 & n6760;
  assign n6762 = ~n6544 & ~n6755;
  assign n6763 = n6544 & n6702;
  assign n6764 = ~pi223 & ~n6763;
  assign n6765 = ~n59161 & n6764;
  assign n6766 = n2790 & ~n6729;
  assign n6767 = ~n2790 & n6740;
  assign n6768 = pi223 & ~n6767;
  assign n6769 = ~n6766 & n6768;
  assign n6770 = ~n59161 & ~n6763;
  assign n6771 = ~pi223 & ~n6770;
  assign n6772 = n2790 & n6729;
  assign n6773 = ~n2790 & ~n6740;
  assign n6774 = pi223 & ~n6773;
  assign n6775 = ~n6772 & n6774;
  assign n6776 = ~n6771 & ~n6775;
  assign n6777 = ~n6765 & ~n6769;
  assign n6778 = ~pi299 & n59162;
  assign n6779 = pi299 & ~n59160;
  assign n6780 = ~pi299 & ~n59162;
  assign n6781 = ~n6779 & ~n6780;
  assign n6782 = ~n6752 & ~n6778;
  assign n6783 = pi39 & ~n59163;
  assign n6784 = ~pi39 & ~n59157;
  assign n6785 = pi39 & n59163;
  assign n6786 = ~n6784 & ~n6785;
  assign n6787 = ~n6683 & ~n6783;
  assign n6788 = ~pi761 & n59164;
  assign n6789 = ~pi140 & ~n6788;
  assign n6790 = ~n6657 & n6789;
  assign n6791 = pi603 & ~n6669;
  assign n6792 = ~pi299 & ~n6791;
  assign n6793 = ~pi210 & ~n6664;
  assign n6794 = pi210 & ~n6667;
  assign n6795 = ~n6793 & ~n6794;
  assign n6796 = pi603 & n6795;
  assign n6797 = pi299 & ~n6796;
  assign n6798 = ~n6792 & ~n6797;
  assign n6799 = ~pi39 & ~n6798;
  assign n6800 = n6587 & n6701;
  assign n6801 = n2781 & ~n6800;
  assign n6802 = n6700 & ~n6800;
  assign n6803 = n6464 & n6701;
  assign n6804 = ~n6700 & ~n6803;
  assign n6805 = ~n6700 & n6803;
  assign n6806 = n6700 & n6800;
  assign n6807 = ~n6805 & ~n6806;
  assign n6808 = ~n6802 & ~n6804;
  assign n6809 = ~n2781 & n59165;
  assign n6810 = n2781 & n6800;
  assign n6811 = ~n2781 & ~n59165;
  assign n6812 = ~n6810 & ~n6811;
  assign n6813 = ~n6801 & ~n6809;
  assign n6814 = n58846 & n59166;
  assign n6815 = n59152 & n6701;
  assign n6816 = ~n58846 & ~n6815;
  assign n6817 = ~n6629 & ~n6816;
  assign n6818 = ~n6629 & ~n6814;
  assign n6819 = ~n6816 & n6818;
  assign n6820 = ~n6814 & n6817;
  assign n6821 = n6463 & n6629;
  assign n6822 = n2794 & n6701;
  assign n6823 = n6629 & n6803;
  assign n6824 = n6821 & n6822;
  assign n6825 = ~pi215 & ~n59168;
  assign n6826 = ~n59167 & n6825;
  assign n6827 = ~n6489 & n6803;
  assign n6828 = ~n6486 & n6803;
  assign n6829 = n6489 & n6700;
  assign n6830 = n6828 & ~n6829;
  assign n6831 = ~n2781 & n6830;
  assign n6832 = ~n6827 & ~n6831;
  assign n6833 = ~n58846 & n6486;
  assign n6834 = ~n6832 & ~n6833;
  assign n6835 = pi215 & ~n6834;
  assign n6836 = pi299 & ~n6835;
  assign n6837 = ~n6826 & n6836;
  assign n6838 = n59155 & n6701;
  assign n6839 = n6622 & n6822;
  assign n6840 = ~pi223 & ~n59169;
  assign n6841 = n2790 & n59166;
  assign n6842 = ~n2790 & ~n6815;
  assign n6843 = ~n6544 & ~n6842;
  assign n6844 = ~n6544 & ~n6841;
  assign n6845 = ~n6842 & n6844;
  assign n6846 = ~n6841 & n6843;
  assign n6847 = n6840 & ~n59170;
  assign n6848 = ~n2790 & n6486;
  assign n6849 = ~n6832 & ~n6848;
  assign n6850 = pi223 & ~n6849;
  assign n6851 = ~pi299 & ~n6850;
  assign n6852 = ~n6847 & n6851;
  assign n6853 = ~n6837 & ~n6852;
  assign n6854 = pi39 & n6853;
  assign n6855 = ~n6799 & ~n6854;
  assign n6856 = pi140 & ~pi761;
  assign n6857 = n6855 & n6856;
  assign n6858 = ~n6790 & ~n6857;
  assign n6859 = ~pi38 & ~n6858;
  assign n6860 = ~pi39 & ~pi95;
  assign n6861 = n2661 & n6860;
  assign n6862 = ~pi39 & n58822;
  assign n6863 = n2794 & n59171;
  assign n6864 = ~pi140 & ~n6863;
  assign n6865 = n6822 & n59171;
  assign n6866 = ~pi761 & n6865;
  assign n6867 = ~n6864 & ~n6866;
  assign n6868 = pi38 & ~n6867;
  assign n6869 = ~n6859 & ~n6868;
  assign n6870 = pi738 & ~n6869;
  assign n6871 = pi680 & ~n6518;
  assign n6872 = pi665 & pi1091;
  assign n6873 = ~n6701 & ~n6872;
  assign n6874 = n6464 & ~n6873;
  assign n6875 = pi616 & ~n6874;
  assign n6876 = pi614 & ~n6874;
  assign n6877 = pi642 & ~n6874;
  assign n6878 = n6589 & ~n6873;
  assign n6879 = ~pi642 & ~n6878;
  assign n6880 = ~n6877 & ~n6879;
  assign n6881 = ~pi614 & ~n6880;
  assign n6882 = ~n6876 & ~n6881;
  assign n6883 = ~pi616 & ~n6882;
  assign n6884 = ~n6875 & ~n6883;
  assign n6885 = n6871 & ~n6884;
  assign n6886 = ~pi680 & ~n6595;
  assign n6887 = n6464 & n6872;
  assign n6888 = n2680 & ~n6887;
  assign n6889 = n6562 & n6872;
  assign n6890 = ~n2680 & ~n6889;
  assign n6891 = ~n6888 & ~n6890;
  assign n6892 = ~pi603 & ~n6891;
  assign n6893 = pi603 & ~pi665;
  assign n6894 = n6684 & n6893;
  assign n6895 = ~n6588 & ~n6894;
  assign n6896 = ~n6892 & n6895;
  assign n6897 = n2781 & ~n6896;
  assign n6898 = ~n6886 & ~n6897;
  assign n6899 = ~n6885 & n6898;
  assign n6900 = n2790 & n6899;
  assign n6901 = ~n59151 & ~n6873;
  assign n6902 = n6871 & ~n6901;
  assign n6903 = ~pi680 & n59151;
  assign n6904 = pi603 & n6687;
  assign n6905 = pi603 & ~pi621;
  assign n6906 = n6889 & ~n6905;
  assign n6907 = n2781 & ~n6906;
  assign n6908 = ~n6904 & n6907;
  assign n6909 = ~n6903 & ~n6908;
  assign n6910 = ~n6902 & n6909;
  assign n6911 = ~n2790 & n6910;
  assign n6912 = ~n6544 & ~n6911;
  assign n6913 = ~n6900 & n6912;
  assign n6914 = pi680 & n6873;
  assign n6915 = n6464 & ~n6914;
  assign n6916 = n6544 & ~n6915;
  assign n6917 = ~pi223 & ~n6916;
  assign n6918 = ~n6913 & n6917;
  assign n6919 = pi665 & n6477;
  assign n6920 = ~n6484 & n6803;
  assign n6921 = ~n6919 & ~n6920;
  assign n6922 = n6465 & n6872;
  assign n6923 = ~pi603 & n6922;
  assign n6924 = n6921 & ~n6923;
  assign n6925 = ~n2680 & ~n6919;
  assign n6926 = ~n6888 & ~n6925;
  assign n6927 = ~pi642 & ~n6926;
  assign n6928 = ~n6827 & n6927;
  assign n6929 = n6924 & n6928;
  assign n6930 = ~n6877 & ~n6929;
  assign n6931 = ~pi614 & ~n6930;
  assign n6932 = ~n6876 & ~n6931;
  assign n6933 = ~pi616 & ~n6932;
  assign n6934 = ~n6875 & ~n6933;
  assign n6935 = n6871 & ~n6934;
  assign n6936 = ~pi680 & ~n6502;
  assign n6937 = n2781 & ~n6926;
  assign n6938 = ~n6827 & n6937;
  assign n6939 = ~n6936 & ~n6938;
  assign n6940 = ~n6935 & n6939;
  assign n6941 = n2790 & ~n6940;
  assign n6942 = ~pi680 & ~n6496;
  assign n6943 = ~n6919 & ~n6922;
  assign n6944 = ~n6828 & n6943;
  assign n6945 = ~n6700 & n6944;
  assign n6946 = n6700 & n6924;
  assign n6947 = ~n6945 & ~n6946;
  assign n6948 = n6871 & ~n6947;
  assign n6949 = n2781 & n6921;
  assign n6950 = ~n6948 & ~n6949;
  assign n6951 = ~n6942 & ~n6949;
  assign n6952 = ~n6948 & n6951;
  assign n6953 = ~n6942 & n6950;
  assign n6954 = ~n2790 & ~n59172;
  assign n6955 = pi223 & ~n6954;
  assign n6956 = ~n6941 & n6955;
  assign n6957 = ~n6900 & ~n6911;
  assign n6958 = ~n6544 & ~n6957;
  assign n6959 = n6544 & n6915;
  assign n6960 = ~pi223 & ~n6959;
  assign n6961 = ~n6958 & n6960;
  assign n6962 = n2790 & n6940;
  assign n6963 = ~n2790 & n59172;
  assign n6964 = pi223 & ~n6963;
  assign n6965 = ~n6962 & n6964;
  assign n6966 = ~n6961 & ~n6965;
  assign n6967 = ~n6918 & ~n6956;
  assign n6968 = ~pi299 & ~n59173;
  assign n6969 = n58846 & n6899;
  assign n6970 = ~n58846 & n6910;
  assign n6971 = ~n6629 & ~n6970;
  assign n6972 = ~n58846 & ~n6910;
  assign n6973 = n58846 & ~n6899;
  assign n6974 = ~n6972 & ~n6973;
  assign n6975 = ~n6969 & ~n6970;
  assign n6976 = ~n6629 & ~n59174;
  assign n6977 = ~n6969 & n6971;
  assign n6978 = n6629 & ~n6915;
  assign n6979 = ~pi215 & ~n6978;
  assign n6980 = ~n59175 & n6979;
  assign n6981 = n58846 & ~n6940;
  assign n6982 = ~n58846 & ~n59172;
  assign n6983 = pi215 & ~n6982;
  assign n6984 = ~n6981 & n6983;
  assign n6985 = ~n6629 & n59174;
  assign n6986 = n6629 & n6915;
  assign n6987 = ~pi215 & ~n6986;
  assign n6988 = ~n6985 & n6987;
  assign n6989 = n58846 & n6940;
  assign n6990 = ~n58846 & n59172;
  assign n6991 = pi215 & ~n6990;
  assign n6992 = ~n6989 & n6991;
  assign n6993 = ~n6988 & ~n6992;
  assign n6994 = ~n6980 & ~n6984;
  assign n6995 = pi299 & ~n59176;
  assign n6996 = ~pi299 & n59173;
  assign n6997 = pi299 & n59176;
  assign n6998 = ~n6996 & ~n6997;
  assign n6999 = ~n6968 & ~n6995;
  assign n7000 = ~pi140 & n59177;
  assign n7001 = pi665 & ~n6565;
  assign n7002 = ~pi665 & n6562;
  assign n7003 = ~n6565 & ~n7002;
  assign n7004 = ~n6566 & ~n7001;
  assign n7005 = ~pi603 & n6568;
  assign n7006 = n2680 & n6685;
  assign n7007 = n6465 & n6684;
  assign n7008 = pi603 & ~n7007;
  assign n7009 = n2680 & n6562;
  assign n7010 = ~n6465 & ~n7009;
  assign n7011 = pi603 & n7010;
  assign n7012 = ~n6701 & ~n7011;
  assign n7013 = ~n7006 & n7008;
  assign n7014 = ~n7005 & n59179;
  assign n7015 = ~n59178 & n7014;
  assign n7016 = pi616 & ~n7015;
  assign n7017 = ~n6699 & n7015;
  assign n7018 = n6684 & n7002;
  assign n7019 = ~pi665 & n6685;
  assign n7020 = pi603 & ~n59180;
  assign n7021 = ~n6568 & ~n59178;
  assign n7022 = ~pi603 & ~n7021;
  assign n7023 = ~n7020 & ~n7022;
  assign n7024 = n6699 & n7023;
  assign n7025 = ~pi616 & ~n7024;
  assign n7026 = ~n7015 & n7025;
  assign n7027 = ~n7017 & n7025;
  assign n7028 = ~n7016 & ~n59181;
  assign n7029 = ~n6518 & ~n7028;
  assign n7030 = n2781 & ~n59178;
  assign n7031 = ~n7020 & n7030;
  assign n7032 = ~n6871 & ~n7031;
  assign n7033 = ~n7029 & ~n7032;
  assign n7034 = ~n58846 & ~n7033;
  assign n7035 = n6464 & ~n6872;
  assign n7036 = ~n6701 & n7035;
  assign n7037 = n6702 & ~n6872;
  assign n7038 = pi616 & ~n59182;
  assign n7039 = n6871 & ~n7038;
  assign n7040 = pi603 & pi665;
  assign n7041 = ~pi603 & ~n7035;
  assign n7042 = ~n7040 & ~n7041;
  assign n7043 = ~n6696 & n7042;
  assign n7044 = n6699 & n7043;
  assign n7045 = ~n6699 & n59182;
  assign n7046 = ~pi616 & ~n7045;
  assign n7047 = ~n7044 & n7046;
  assign n7048 = n7039 & ~n7047;
  assign n7049 = n6587 & n6897;
  assign n7050 = ~n7048 & ~n7049;
  assign n7051 = n58846 & n7050;
  assign n7052 = ~n6629 & ~n7051;
  assign n7053 = ~n7034 & n7052;
  assign n7054 = pi680 & ~n6872;
  assign n7055 = n2794 & n7054;
  assign n7056 = ~n6701 & n7055;
  assign n7057 = n6637 & n6914;
  assign n7058 = n6821 & n7056;
  assign n7059 = ~pi215 & ~n59183;
  assign n7060 = ~n7053 & n7059;
  assign n7061 = n6732 & n7042;
  assign n7062 = ~n6724 & n7042;
  assign n7063 = ~pi642 & ~n7062;
  assign n7064 = n2777 & n7063;
  assign n7065 = ~pi614 & n7063;
  assign n7066 = n7061 & ~n7065;
  assign n7067 = pi614 & ~pi616;
  assign n7068 = ~n7061 & n7067;
  assign n7069 = n7061 & ~n7063;
  assign n7070 = n2777 & ~n7069;
  assign n7071 = ~n7068 & ~n7070;
  assign n7072 = ~pi616 & ~n7066;
  assign n7073 = pi616 & ~n7061;
  assign n7074 = n59184 & ~n7073;
  assign n7075 = n7061 & ~n7064;
  assign n7076 = ~n6518 & ~n59185;
  assign n7077 = ~n6484 & n6914;
  assign n7078 = ~n6871 & ~n7077;
  assign n7079 = ~n7076 & ~n7078;
  assign n7080 = ~n58846 & n7079;
  assign n7081 = ~n6727 & ~n6872;
  assign n7082 = ~pi616 & ~n7081;
  assign n7083 = n7039 & ~n7082;
  assign n7084 = n6725 & n7042;
  assign n7085 = n6514 & n7062;
  assign n7086 = ~n7083 & ~n59186;
  assign n7087 = n58846 & ~n7086;
  assign n7088 = pi215 & ~n7087;
  assign n7089 = ~n7080 & n7088;
  assign n7090 = ~n7060 & ~n7089;
  assign n7091 = pi299 & ~n7090;
  assign n7092 = ~n2790 & n7033;
  assign n7093 = n2790 & ~n7050;
  assign n7094 = ~n6544 & ~n7093;
  assign n7095 = ~n7092 & n7094;
  assign n7096 = ~n6701 & ~n7054;
  assign n7097 = ~n6822 & ~n7056;
  assign n7098 = n6464 & ~n7097;
  assign n7099 = n6464 & ~n7096;
  assign n7100 = n6544 & ~n59187;
  assign n7101 = ~pi223 & ~n7100;
  assign n7102 = ~n59169 & n7101;
  assign n7103 = n6840 & ~n7100;
  assign n7104 = ~n7095 & n59188;
  assign n7105 = ~n2790 & ~n7079;
  assign n7106 = n2790 & n7086;
  assign n7107 = pi223 & ~n7106;
  assign n7108 = ~n7105 & n7107;
  assign n7109 = ~pi299 & ~n7108;
  assign n7110 = ~n7104 & n7109;
  assign n7111 = ~n7091 & ~n7110;
  assign n7112 = pi140 & n7111;
  assign n7113 = pi761 & ~n7112;
  assign n7114 = ~n7000 & n7113;
  assign n7115 = ~n6904 & ~n7023;
  assign n7116 = n6700 & ~n7115;
  assign n7117 = ~n6568 & n6701;
  assign n7118 = ~n7021 & ~n7117;
  assign n7119 = ~n6700 & ~n7118;
  assign n7120 = n6871 & ~n7119;
  assign n7121 = ~n6700 & n7118;
  assign n7122 = n6700 & ~n7023;
  assign n7123 = ~n6904 & n7122;
  assign n7124 = ~n7121 & ~n7123;
  assign n7125 = n6871 & ~n7124;
  assign n7126 = ~n7116 & n7120;
  assign n7127 = ~n6871 & ~n7030;
  assign n7128 = ~n6815 & n7127;
  assign n7129 = ~n59189 & ~n7128;
  assign n7130 = ~n58846 & ~n7129;
  assign n7131 = n6872 & ~n6905;
  assign n7132 = n6464 & ~n7131;
  assign n7133 = ~n6700 & n7132;
  assign n7134 = n6871 & ~n7133;
  assign n7135 = ~n6800 & ~n7043;
  assign n7136 = n6700 & ~n7135;
  assign n7137 = n7134 & ~n7136;
  assign n7138 = ~pi680 & n59165;
  assign n7139 = n6587 & ~n59178;
  assign n7140 = n2781 & ~n7139;
  assign n7141 = ~n6800 & n7140;
  assign n7142 = n6801 & ~n7139;
  assign n7143 = ~n7138 & ~n59190;
  assign n7144 = ~n7137 & n7143;
  assign n7145 = n58846 & ~n7144;
  assign n7146 = ~n6629 & ~n7145;
  assign n7147 = ~n58846 & n7129;
  assign n7148 = n58846 & n7144;
  assign n7149 = ~n7147 & ~n7148;
  assign n7150 = ~n6629 & ~n7149;
  assign n7151 = ~n7130 & n7146;
  assign n7152 = n6637 & ~n7096;
  assign n7153 = n6629 & n59187;
  assign n7154 = ~pi215 & ~n59192;
  assign n7155 = ~n59191 & n7154;
  assign n7156 = ~n2778 & n7035;
  assign n7157 = ~n6489 & n7035;
  assign n7158 = ~n7156 & ~n7157;
  assign n7159 = ~n6827 & n7158;
  assign n7160 = n6700 & ~n7159;
  assign n7161 = n7134 & ~n7160;
  assign n7162 = n6518 & ~n7157;
  assign n7163 = pi680 & ~n7162;
  assign n7164 = n6832 & ~n7163;
  assign n7165 = ~n7161 & ~n7164;
  assign n7166 = n58846 & n7165;
  assign n7167 = ~n6831 & ~n6920;
  assign n7168 = ~n7158 & n7163;
  assign n7169 = ~n6486 & n7035;
  assign n7170 = n7168 & n7169;
  assign n7171 = n7167 & ~n7170;
  assign n7172 = ~n58846 & ~n7171;
  assign n7173 = pi215 & ~n7172;
  assign n7174 = ~n7166 & n7173;
  assign n7175 = ~n7155 & ~n7174;
  assign n7176 = pi299 & ~n7175;
  assign n7177 = ~n2790 & n7129;
  assign n7178 = n2790 & n7144;
  assign n7179 = ~n6544 & ~n7178;
  assign n7180 = ~n7177 & n7179;
  assign n7181 = n7101 & ~n7180;
  assign n7182 = n2790 & ~n7165;
  assign n7183 = ~n2790 & n7171;
  assign n7184 = pi223 & ~n7183;
  assign n7185 = ~n7182 & n7184;
  assign n7186 = ~pi299 & ~n7185;
  assign n7187 = ~n7181 & n7186;
  assign n7188 = ~n7176 & ~n7187;
  assign n7189 = pi140 & n7188;
  assign n7190 = ~pi680 & n6706;
  assign n7191 = n6705 & n6872;
  assign n7192 = n6887 & ~n6905;
  assign n7193 = ~n6700 & n7192;
  assign n7194 = n6871 & ~n7193;
  assign n7195 = ~n7191 & n7194;
  assign n7196 = n6891 & n7131;
  assign n7197 = n2781 & ~n7196;
  assign n7198 = ~n7195 & ~n7197;
  assign n7199 = ~n7190 & ~n7197;
  assign n7200 = ~n7195 & n7199;
  assign n7201 = ~n7190 & n7198;
  assign n7202 = n2790 & ~n59193;
  assign n7203 = ~n59151 & ~n6701;
  assign n7204 = ~pi680 & ~n7203;
  assign n7205 = ~n2821 & n6889;
  assign n7206 = ~n2778 & n6887;
  assign n7207 = ~n2778 & n6922;
  assign n7208 = ~n2680 & n7206;
  assign n7209 = ~n7205 & ~n59194;
  assign n7210 = n7131 & ~n7209;
  assign n7211 = n6871 & ~n7210;
  assign n7212 = ~n6907 & ~n7211;
  assign n7213 = ~n7204 & n7212;
  assign n7214 = ~n2790 & ~n7213;
  assign n7215 = ~n6544 & ~n7214;
  assign n7216 = ~n2790 & n7213;
  assign n7217 = n2790 & n59193;
  assign n7218 = ~n7216 & ~n7217;
  assign n7219 = ~n7202 & ~n7214;
  assign n7220 = ~n6544 & ~n59195;
  assign n7221 = ~n7202 & n7215;
  assign n7222 = n6468 & n7096;
  assign n7223 = ~n6461 & n7222;
  assign n7224 = n6544 & n7223;
  assign n7225 = ~pi223 & ~n7224;
  assign n7226 = ~n59196 & n7225;
  assign n7227 = n6728 & ~n7054;
  assign n7228 = n2781 & ~n6905;
  assign n7229 = n6926 & n7228;
  assign n7230 = ~n7227 & ~n7229;
  assign n7231 = n2790 & ~n7230;
  assign n7232 = ~n6727 & ~n6943;
  assign n7233 = n6871 & ~n7232;
  assign n7234 = ~pi680 & ~n6734;
  assign n7235 = pi680 & ~n6919;
  assign n7236 = ~n6905 & ~n7235;
  assign n7237 = n2781 & ~n7236;
  assign n7238 = ~n7234 & ~n7237;
  assign n7239 = ~n7233 & n7238;
  assign n7240 = ~n2790 & n7239;
  assign n7241 = pi223 & ~n7240;
  assign n7242 = pi223 & ~n7231;
  assign n7243 = ~n7240 & n7242;
  assign n7244 = ~n7231 & n7241;
  assign n7245 = ~n6544 & n59195;
  assign n7246 = n6544 & ~n7223;
  assign n7247 = ~pi223 & ~n7246;
  assign n7248 = ~n7245 & n7247;
  assign n7249 = ~n2790 & ~n7239;
  assign n7250 = n2790 & n7230;
  assign n7251 = pi223 & ~n7250;
  assign n7252 = ~n7249 & n7251;
  assign n7253 = ~n7248 & ~n7252;
  assign n7254 = ~n7226 & ~n59197;
  assign n7255 = ~pi299 & ~n59198;
  assign n7256 = n58846 & ~n59193;
  assign n7257 = ~n58846 & ~n7213;
  assign n7258 = ~n6629 & ~n7257;
  assign n7259 = ~n58846 & n7213;
  assign n7260 = n58846 & n59193;
  assign n7261 = ~n7259 & ~n7260;
  assign n7262 = ~n7256 & ~n7257;
  assign n7263 = ~n6629 & ~n59199;
  assign n7264 = ~n7256 & n7258;
  assign n7265 = n6629 & n7223;
  assign n7266 = ~pi215 & ~n7265;
  assign n7267 = ~n59200 & n7266;
  assign n7268 = n58846 & ~n7230;
  assign n7269 = ~n58846 & n7239;
  assign n7270 = pi215 & ~n7269;
  assign n7271 = pi215 & ~n7268;
  assign n7272 = ~n7269 & n7271;
  assign n7273 = ~n7268 & n7270;
  assign n7274 = ~n6629 & n59199;
  assign n7275 = n6629 & ~n7223;
  assign n7276 = ~pi215 & ~n7275;
  assign n7277 = ~n7274 & n7276;
  assign n7278 = ~n58846 & ~n7239;
  assign n7279 = n58846 & n7230;
  assign n7280 = pi215 & ~n7279;
  assign n7281 = ~n7278 & n7280;
  assign n7282 = ~n7277 & ~n7281;
  assign n7283 = ~n7267 & ~n59201;
  assign n7284 = pi299 & ~n59202;
  assign n7285 = ~pi299 & n59198;
  assign n7286 = pi299 & n59202;
  assign n7287 = ~n7285 & ~n7286;
  assign n7288 = ~n7255 & ~n7284;
  assign n7289 = ~pi140 & ~n59203;
  assign n7290 = ~pi761 & ~n7289;
  assign n7291 = ~n7189 & n7290;
  assign n7292 = ~n7114 & ~n7291;
  assign n7293 = pi39 & ~n7292;
  assign n7294 = pi665 & n6446;
  assign n7295 = pi198 & ~n7294;
  assign n7296 = pi665 & n6420;
  assign n7297 = ~pi198 & ~n7296;
  assign n7298 = ~n7295 & ~n7297;
  assign n7299 = pi680 & ~n7298;
  assign n7300 = n6449 & ~n7299;
  assign n7301 = ~pi299 & ~n7300;
  assign n7302 = ~pi210 & ~n7296;
  assign n7303 = pi210 & ~n7294;
  assign n7304 = ~n7302 & ~n7303;
  assign n7305 = pi680 & ~n7304;
  assign n7306 = n6453 & ~n7305;
  assign n7307 = pi299 & ~n7306;
  assign n7308 = ~n7301 & ~n7307;
  assign n7309 = pi680 & n6798;
  assign n7310 = ~n7308 & ~n7309;
  assign n7311 = ~pi140 & ~n7310;
  assign n7312 = pi665 & ~n6421;
  assign n7313 = ~n6422 & ~n7312;
  assign n7314 = ~pi198 & ~n7313;
  assign n7315 = pi665 & ~n6435;
  assign n7316 = ~n6447 & ~n7315;
  assign n7317 = pi198 & ~n7316;
  assign n7318 = ~n7314 & ~n7317;
  assign n7319 = ~pi603 & ~n7318;
  assign n7320 = pi603 & ~n6662;
  assign n7321 = ~n7040 & ~n7320;
  assign n7322 = ~n7319 & n7321;
  assign n7323 = pi680 & n7322;
  assign n7324 = ~pi299 & ~n7323;
  assign n7325 = pi210 & ~n7316;
  assign n7326 = ~pi210 & ~n7313;
  assign n7327 = ~n7325 & ~n7326;
  assign n7328 = ~pi603 & ~n7327;
  assign n7329 = ~n6676 & ~n7040;
  assign n7330 = ~n7328 & n7329;
  assign n7331 = pi680 & n7330;
  assign n7332 = pi299 & ~n7331;
  assign n7333 = ~n7324 & ~n7332;
  assign n7334 = pi140 & ~n7333;
  assign n7335 = pi761 & ~n7334;
  assign n7336 = pi761 & ~n7311;
  assign n7337 = ~n7334 & n7336;
  assign n7338 = ~n7311 & n7335;
  assign n7339 = n59157 & n7308;
  assign n7340 = ~pi140 & n7339;
  assign n7341 = pi680 & n7318;
  assign n7342 = ~pi299 & ~n7341;
  assign n7343 = pi680 & n7327;
  assign n7344 = pi299 & ~n7343;
  assign n7345 = ~n7342 & ~n7344;
  assign n7346 = pi140 & ~n7345;
  assign n7347 = ~n6798 & ~n7345;
  assign n7348 = pi140 & n7347;
  assign n7349 = ~n6798 & n7346;
  assign n7350 = ~pi761 & ~n59205;
  assign n7351 = ~n7340 & n7350;
  assign n7352 = ~pi39 & ~n7351;
  assign n7353 = ~n7340 & ~n59205;
  assign n7354 = ~pi761 & ~n7353;
  assign n7355 = pi140 & n7333;
  assign n7356 = ~pi140 & n7310;
  assign n7357 = pi761 & ~n7356;
  assign n7358 = ~n7355 & n7357;
  assign n7359 = ~n7354 & ~n7358;
  assign n7360 = ~pi39 & ~n7359;
  assign n7361 = ~n59204 & n7352;
  assign n7362 = ~pi38 & ~n59206;
  assign n7363 = ~n7293 & n7362;
  assign n7364 = pi761 & n6701;
  assign n7365 = n6863 & ~n7096;
  assign n7366 = n6468 & ~n7096;
  assign n7367 = ~pi39 & n7366;
  assign n7368 = n59171 & ~n7097;
  assign n7369 = ~n7364 & n59207;
  assign n7370 = ~n6864 & ~n7369;
  assign n7371 = ~pi761 & n7366;
  assign n7372 = ~pi140 & ~n6468;
  assign n7373 = n6468 & n6914;
  assign n7374 = n58822 & n7056;
  assign n7375 = pi761 & n59208;
  assign n7376 = ~pi39 & ~n7375;
  assign n7377 = ~n7372 & n7376;
  assign n7378 = ~pi140 & ~n7222;
  assign n7379 = pi140 & ~n7097;
  assign n7380 = n58822 & n7379;
  assign n7381 = ~pi761 & ~n7380;
  assign n7382 = ~n7378 & n7381;
  assign n7383 = pi761 & ~n7372;
  assign n7384 = ~n59208 & n7383;
  assign n7385 = ~n7382 & ~n7384;
  assign n7386 = ~pi39 & ~n7385;
  assign n7387 = ~n7371 & n7377;
  assign n7388 = pi39 & pi140;
  assign n7389 = pi38 & ~n7388;
  assign n7390 = ~n59209 & n7389;
  assign n7391 = pi38 & ~n7370;
  assign n7392 = ~n7363 & ~n59210;
  assign n7393 = ~pi738 & ~n7392;
  assign n7394 = n59132 & ~n7393;
  assign n7395 = n59132 & ~n6870;
  assign n7396 = ~n7393 & n7395;
  assign n7397 = ~n6870 & n7394;
  assign n7398 = ~n6314 & ~n59211;
  assign n7399 = ~pi778 & ~n7398;
  assign n7400 = pi625 & n7398;
  assign n7401 = n59132 & n6869;
  assign n7402 = ~n6314 & ~n7401;
  assign n7403 = ~pi625 & n7402;
  assign n7404 = pi1153 & ~n7403;
  assign n7405 = ~n7400 & n7404;
  assign n7406 = ~pi140 & n7308;
  assign n7407 = ~n7346 & ~n7406;
  assign n7408 = ~pi140 & ~n7308;
  assign n7409 = pi140 & n7345;
  assign n7410 = ~pi39 & ~n7409;
  assign n7411 = ~n7408 & n7410;
  assign n7412 = ~pi39 & ~n7408;
  assign n7413 = ~n7409 & n7412;
  assign n7414 = ~pi39 & ~n7407;
  assign n7415 = n2778 & n6891;
  assign n7416 = pi680 & ~n7206;
  assign n7417 = ~n7415 & n7416;
  assign n7418 = ~n6886 & ~n7417;
  assign n7419 = ~n6518 & n7418;
  assign n7420 = pi680 & ~n6891;
  assign n7421 = n6518 & ~n7420;
  assign n7422 = ~n6886 & n7421;
  assign n7423 = ~n7419 & ~n7422;
  assign n7424 = n58846 & n7423;
  assign n7425 = ~n6518 & ~n7209;
  assign n7426 = n6518 & n6889;
  assign n7427 = pi680 & ~n7426;
  assign n7428 = ~n7425 & n7427;
  assign n7429 = ~n6903 & ~n7428;
  assign n7430 = ~n58846 & ~n7429;
  assign n7431 = ~n6629 & ~n7430;
  assign n7432 = ~n7424 & n7431;
  assign n7433 = n2794 & ~n7054;
  assign n7434 = n6637 & ~n7054;
  assign n7435 = n6821 & n7433;
  assign n7436 = ~pi215 & ~n59213;
  assign n7437 = ~n7432 & n7436;
  assign n7438 = ~n6926 & n7416;
  assign n7439 = ~n6937 & ~n7438;
  assign n7440 = ~n6936 & ~n7438;
  assign n7441 = ~n6937 & n7440;
  assign n7442 = ~n6936 & n7439;
  assign n7443 = n58846 & n59214;
  assign n7444 = ~n59194 & n7235;
  assign n7445 = ~n6942 & ~n7444;
  assign n7446 = n7439 & n7445;
  assign n7447 = ~n58846 & n7446;
  assign n7448 = pi215 & ~n7447;
  assign n7449 = pi215 & ~n7443;
  assign n7450 = ~n7447 & n7449;
  assign n7451 = ~n7443 & n7448;
  assign n7452 = ~n7432 & ~n59213;
  assign n7453 = ~pi215 & ~n7452;
  assign n7454 = n58846 & ~n59214;
  assign n7455 = ~n58846 & ~n7446;
  assign n7456 = pi215 & ~n7455;
  assign n7457 = ~n7454 & n7456;
  assign n7458 = ~n7453 & ~n7457;
  assign n7459 = ~n7437 & ~n59215;
  assign n7460 = pi299 & ~n59216;
  assign n7461 = n2790 & n7423;
  assign n7462 = ~n2790 & ~n7429;
  assign n7463 = ~n6544 & ~n7462;
  assign n7464 = ~n7461 & n7463;
  assign n7465 = n59155 & ~n7054;
  assign n7466 = n6622 & n7433;
  assign n7467 = ~pi223 & ~n59217;
  assign n7468 = ~n7464 & n7467;
  assign n7469 = n2790 & n59214;
  assign n7470 = ~n2790 & n7446;
  assign n7471 = pi223 & ~n7470;
  assign n7472 = pi223 & ~n7469;
  assign n7473 = ~n7470 & n7472;
  assign n7474 = ~n7469 & n7471;
  assign n7475 = ~n7464 & ~n59217;
  assign n7476 = ~pi223 & ~n7475;
  assign n7477 = n2790 & ~n59214;
  assign n7478 = ~n2790 & ~n7446;
  assign n7479 = pi223 & ~n7478;
  assign n7480 = ~n7477 & n7479;
  assign n7481 = ~n7476 & ~n7480;
  assign n7482 = ~n7468 & ~n59218;
  assign n7483 = ~pi299 & ~n59219;
  assign n7484 = ~pi299 & n59219;
  assign n7485 = pi299 & n59216;
  assign n7486 = ~n7484 & ~n7485;
  assign n7487 = ~n7460 & ~n7483;
  assign n7488 = ~pi140 & ~n59220;
  assign n7489 = n59155 & n7054;
  assign n7490 = ~n59151 & n7054;
  assign n7491 = ~n6518 & n7490;
  assign n7492 = ~n7030 & ~n7491;
  assign n7493 = ~n2790 & n7492;
  assign n7494 = n2778 & n7139;
  assign n7495 = ~n7156 & ~n7494;
  assign n7496 = ~n6518 & n7495;
  assign n7497 = n6518 & ~n7139;
  assign n7498 = pi680 & ~n7497;
  assign n7499 = ~n7496 & n7498;
  assign n7500 = n2790 & ~n7499;
  assign n7501 = ~n6544 & ~n7500;
  assign n7502 = ~n6544 & ~n7493;
  assign n7503 = ~n7500 & n7502;
  assign n7504 = ~n7493 & n7501;
  assign n7505 = ~n7489 & ~n59221;
  assign n7506 = ~pi223 & ~n7505;
  assign n7507 = pi680 & ~n7158;
  assign n7508 = ~n6848 & n7507;
  assign n7509 = pi223 & ~n7162;
  assign n7510 = n7508 & n7509;
  assign n7511 = ~n7506 & ~n7510;
  assign n7512 = ~pi299 & ~n7511;
  assign n7513 = ~n58846 & ~n7492;
  assign n7514 = n58846 & n7499;
  assign n7515 = ~n6629 & ~n7514;
  assign n7516 = ~n7513 & n7515;
  assign n7517 = pi680 & n7035;
  assign n7518 = n6464 & n7054;
  assign n7519 = n6629 & ~n59222;
  assign n7520 = ~pi215 & ~n7519;
  assign n7521 = n58846 & ~n7499;
  assign n7522 = ~n58846 & n7492;
  assign n7523 = ~n6629 & ~n7522;
  assign n7524 = ~n7521 & n7523;
  assign n7525 = n6629 & n59222;
  assign n7526 = n6637 & n7054;
  assign n7527 = ~n7524 & ~n59223;
  assign n7528 = ~pi215 & ~n7527;
  assign n7529 = ~n7516 & n7520;
  assign n7530 = pi215 & ~n6833;
  assign n7531 = ~n6833 & n7507;
  assign n7532 = pi215 & ~n7162;
  assign n7533 = n7531 & n7532;
  assign n7534 = n7168 & n7530;
  assign n7535 = ~n59224 & ~n59225;
  assign n7536 = pi299 & ~n7535;
  assign n7537 = ~n7512 & ~n7536;
  assign n7538 = pi140 & ~n7537;
  assign n7539 = pi39 & ~n7538;
  assign n7540 = pi39 & n59220;
  assign n7541 = ~n7388 & ~n7540;
  assign n7542 = ~n7538 & ~n7541;
  assign n7543 = ~n7488 & n7539;
  assign n7544 = ~n59212 & ~n59226;
  assign n7545 = ~pi38 & ~n7544;
  assign n7546 = n59171 & n7055;
  assign n7547 = pi38 & ~n7546;
  assign n7548 = ~n6864 & n7547;
  assign n7549 = ~pi738 & ~n7548;
  assign n7550 = ~n7545 & n7549;
  assign n7551 = ~pi38 & ~n6656;
  assign n7552 = pi38 & ~n6863;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = ~pi140 & pi738;
  assign n7555 = ~n7553 & n7554;
  assign n7556 = n59132 & ~n7555;
  assign n7557 = ~n7550 & n7556;
  assign n7558 = ~n6314 & ~n7557;
  assign n7559 = ~pi625 & n7558;
  assign n7560 = n59132 & n7553;
  assign n7561 = ~pi140 & ~n7560;
  assign n7562 = pi625 & n7561;
  assign n7563 = ~pi1153 & ~n7562;
  assign n7564 = ~n7559 & n7563;
  assign n7565 = pi608 & ~n7564;
  assign n7566 = ~n7405 & n7565;
  assign n7567 = ~pi625 & n7398;
  assign n7568 = pi625 & n7402;
  assign n7569 = ~pi1153 & ~n7568;
  assign n7570 = ~n7567 & n7569;
  assign n7571 = pi625 & n7558;
  assign n7572 = ~pi625 & n7561;
  assign n7573 = pi1153 & ~n7572;
  assign n7574 = ~n7571 & n7573;
  assign n7575 = ~pi608 & ~n7574;
  assign n7576 = ~n7570 & n7575;
  assign n7577 = pi778 & ~n7576;
  assign n7578 = pi778 & ~n7566;
  assign n7579 = ~n7576 & n7578;
  assign n7580 = ~n7566 & n7577;
  assign n7581 = ~n7566 & ~n7576;
  assign n7582 = pi778 & ~n7581;
  assign n7583 = ~pi778 & n7398;
  assign n7584 = ~n7582 & ~n7583;
  assign n7585 = ~n7399 & ~n59227;
  assign n7586 = ~pi609 & ~n59228;
  assign n7587 = ~pi778 & ~n7558;
  assign n7588 = ~n7564 & ~n7574;
  assign n7589 = pi778 & ~n7588;
  assign n7590 = ~n7587 & ~n7589;
  assign n7591 = pi609 & n7590;
  assign n7592 = ~pi1155 & ~n7591;
  assign n7593 = ~n7586 & n7592;
  assign n7594 = pi608 & ~pi1153;
  assign n7595 = ~pi608 & pi1153;
  assign n7596 = ~n7594 & ~n7595;
  assign n7597 = pi778 & ~n7596;
  assign n7598 = pi609 & ~n7597;
  assign n7599 = ~n7561 & ~n7598;
  assign n7600 = ~n7402 & ~n7597;
  assign n7601 = pi609 & n7600;
  assign n7602 = ~n7599 & ~n7601;
  assign n7603 = pi1155 & ~n7602;
  assign n7604 = ~pi660 & ~n7603;
  assign n7605 = ~n7593 & n7604;
  assign n7606 = pi609 & ~n59228;
  assign n7607 = ~pi609 & n7590;
  assign n7608 = pi1155 & ~n7607;
  assign n7609 = ~n7606 & n7608;
  assign n7610 = ~pi609 & ~n7597;
  assign n7611 = ~n7561 & ~n7610;
  assign n7612 = ~pi609 & n7600;
  assign n7613 = ~n7611 & ~n7612;
  assign n7614 = ~pi1155 & ~n7613;
  assign n7615 = pi660 & ~n7614;
  assign n7616 = ~n7609 & n7615;
  assign n7617 = ~n7605 & ~n7616;
  assign n7618 = pi785 & ~n7617;
  assign n7619 = ~pi785 & ~n59228;
  assign n7620 = ~n7618 & ~n7619;
  assign n7621 = ~pi618 & ~n7620;
  assign n7622 = pi660 & ~pi1155;
  assign n7623 = ~pi660 & pi1155;
  assign n7624 = ~n7622 & ~n7623;
  assign n7625 = ~pi660 & ~pi1155;
  assign n7626 = pi660 & pi1155;
  assign n7627 = pi785 & ~n7626;
  assign n7628 = ~n7625 & n7627;
  assign n7629 = pi785 & ~n7625;
  assign n7630 = ~n7626 & n7629;
  assign n7631 = pi785 & ~n7624;
  assign n7632 = n7590 & ~n59229;
  assign n7633 = n7561 & n59229;
  assign n7634 = ~n7561 & n59229;
  assign n7635 = ~n7590 & ~n59229;
  assign n7636 = ~n7634 & ~n7635;
  assign n7637 = ~n7632 & ~n7633;
  assign n7638 = pi618 & n59230;
  assign n7639 = ~pi1154 & ~n7638;
  assign n7640 = ~n7621 & n7639;
  assign n7641 = ~n7561 & n7597;
  assign n7642 = ~n7600 & ~n7641;
  assign n7643 = ~pi785 & ~n7642;
  assign n7644 = ~n7603 & ~n7614;
  assign n7645 = pi785 & ~n7644;
  assign n7646 = ~n7643 & ~n7645;
  assign n7647 = pi618 & n7646;
  assign n7648 = ~pi618 & n7561;
  assign n7649 = pi1154 & ~n7648;
  assign n7650 = ~n7647 & n7649;
  assign n7651 = ~pi627 & ~n7650;
  assign n7652 = ~n7640 & n7651;
  assign n7653 = pi618 & ~n7620;
  assign n7654 = ~pi618 & n59230;
  assign n7655 = pi1154 & ~n7654;
  assign n7656 = ~n7653 & n7655;
  assign n7657 = ~pi618 & n7646;
  assign n7658 = pi618 & n7561;
  assign n7659 = ~pi1154 & ~n7658;
  assign n7660 = ~n7657 & n7659;
  assign n7661 = pi627 & ~n7660;
  assign n7662 = ~n7656 & n7661;
  assign n7663 = ~n7652 & ~n7662;
  assign n7664 = pi781 & ~n7663;
  assign n7665 = ~pi781 & ~n7620;
  assign n7666 = ~n7664 & ~n7665;
  assign n7667 = ~pi619 & ~n7666;
  assign n7668 = pi627 & ~pi1154;
  assign n7669 = ~pi627 & pi1154;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = ~pi627 & ~pi1154;
  assign n7672 = pi627 & pi1154;
  assign n7673 = pi781 & ~n7672;
  assign n7674 = ~n7671 & n7673;
  assign n7675 = pi781 & ~n7671;
  assign n7676 = ~n7672 & n7675;
  assign n7677 = pi781 & ~n7670;
  assign n7678 = ~n59230 & ~n59231;
  assign n7679 = ~n7561 & n59231;
  assign n7680 = n59230 & ~n59231;
  assign n7681 = n7561 & n59231;
  assign n7682 = ~n7680 & ~n7681;
  assign n7683 = ~n7678 & ~n7679;
  assign n7684 = pi619 & ~n59232;
  assign n7685 = ~pi1159 & ~n7684;
  assign n7686 = ~n7667 & n7685;
  assign n7687 = ~pi781 & ~n7646;
  assign n7688 = ~n7650 & ~n7660;
  assign n7689 = pi781 & ~n7688;
  assign n7690 = ~n7687 & ~n7689;
  assign n7691 = pi619 & n7690;
  assign n7692 = ~pi619 & n7561;
  assign n7693 = pi1159 & ~n7692;
  assign n7694 = ~n7691 & n7693;
  assign n7695 = ~pi648 & ~n7694;
  assign n7696 = ~n7686 & n7695;
  assign n7697 = pi619 & ~n7666;
  assign n7698 = ~pi619 & ~n59232;
  assign n7699 = pi1159 & ~n7698;
  assign n7700 = ~n7697 & n7699;
  assign n7701 = ~pi619 & n7690;
  assign n7702 = pi619 & n7561;
  assign n7703 = ~pi1159 & ~n7702;
  assign n7704 = ~n7701 & n7703;
  assign n7705 = pi648 & ~n7704;
  assign n7706 = ~n7700 & n7705;
  assign n7707 = ~n7696 & ~n7706;
  assign n7708 = pi789 & ~n7707;
  assign n7709 = ~pi789 & ~n7666;
  assign n7710 = ~n7708 & ~n7709;
  assign n7711 = ~pi788 & n7710;
  assign n7712 = ~pi626 & n7710;
  assign n7713 = ~pi648 & pi1159;
  assign n7714 = pi648 & ~pi1159;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = pi789 & ~n7715;
  assign n7717 = ~n59232 & ~n7716;
  assign n7718 = n7561 & n7716;
  assign n7719 = ~n7561 & n7716;
  assign n7720 = n59232 & ~n7716;
  assign n7721 = ~n7719 & ~n7720;
  assign n7722 = ~n7717 & ~n7718;
  assign n7723 = pi626 & ~n59233;
  assign n7724 = ~pi641 & ~n7723;
  assign n7725 = ~n7712 & n7724;
  assign n7726 = ~pi641 & ~pi1158;
  assign n7727 = ~pi789 & ~n7690;
  assign n7728 = ~n7694 & ~n7704;
  assign n7729 = pi789 & ~n7728;
  assign n7730 = ~n7727 & ~n7729;
  assign n7731 = ~pi626 & n7730;
  assign n7732 = pi626 & n7561;
  assign n7733 = ~pi1158 & ~n7732;
  assign n7734 = ~n7731 & n7733;
  assign n7735 = ~n7726 & ~n7734;
  assign n7736 = ~n7725 & ~n7735;
  assign n7737 = pi626 & n7710;
  assign n7738 = ~pi626 & ~n59233;
  assign n7739 = pi641 & ~n7738;
  assign n7740 = ~n7737 & n7739;
  assign n7741 = pi641 & pi1158;
  assign n7742 = pi626 & n7730;
  assign n7743 = ~pi626 & n7561;
  assign n7744 = pi1158 & ~n7743;
  assign n7745 = ~n7742 & n7744;
  assign n7746 = ~n7741 & ~n7745;
  assign n7747 = ~n7740 & ~n7746;
  assign n7748 = ~n7736 & ~n7747;
  assign n7749 = pi788 & ~n7748;
  assign n7750 = ~n7711 & ~n7749;
  assign n7751 = ~pi628 & n7750;
  assign n7752 = ~n7734 & ~n7745;
  assign n7753 = pi788 & ~n7752;
  assign n7754 = ~pi788 & ~n7730;
  assign n7755 = ~n7753 & ~n7754;
  assign n7756 = pi628 & n7755;
  assign n7757 = ~pi1156 & ~n7756;
  assign n7758 = ~n7751 & n7757;
  assign n7759 = ~pi641 & pi1158;
  assign n7760 = pi641 & ~pi1158;
  assign n7761 = ~n7759 & ~n7760;
  assign n7762 = pi788 & ~n7761;
  assign n7763 = ~n59233 & ~n7762;
  assign n7764 = ~n7561 & n7762;
  assign n7765 = n59233 & ~n7762;
  assign n7766 = n7561 & n7762;
  assign n7767 = ~n7765 & ~n7766;
  assign n7768 = ~n7763 & ~n7764;
  assign n7769 = pi628 & ~n59234;
  assign n7770 = ~pi628 & n7561;
  assign n7771 = pi1156 & ~n7770;
  assign n7772 = ~n7769 & n7771;
  assign n7773 = ~pi629 & ~n7772;
  assign n7774 = ~n7758 & n7773;
  assign n7775 = pi628 & n7750;
  assign n7776 = ~pi628 & n7755;
  assign n7777 = pi1156 & ~n7776;
  assign n7778 = ~n7775 & n7777;
  assign n7779 = ~pi628 & ~n59234;
  assign n7780 = pi628 & n7561;
  assign n7781 = ~pi1156 & ~n7780;
  assign n7782 = ~n7779 & n7781;
  assign n7783 = pi629 & ~n7782;
  assign n7784 = ~n7778 & n7783;
  assign n7785 = ~n7774 & ~n7784;
  assign n7786 = pi792 & ~n7785;
  assign n7787 = ~pi792 & n7750;
  assign n7788 = ~n7786 & ~n7787;
  assign n7789 = ~pi647 & ~n7788;
  assign n7790 = ~pi629 & pi1156;
  assign n7791 = pi629 & ~pi1156;
  assign n7792 = ~n7790 & ~n7791;
  assign n7793 = pi792 & ~n7792;
  assign n7794 = n7755 & ~n7793;
  assign n7795 = n7561 & n7793;
  assign n7796 = ~n7794 & ~n7795;
  assign n7797 = pi647 & ~n7796;
  assign n7798 = ~pi1157 & ~n7797;
  assign n7799 = ~n7789 & n7798;
  assign n7800 = ~pi792 & n59234;
  assign n7801 = ~n7772 & ~n7782;
  assign n7802 = pi792 & ~n7801;
  assign n7803 = ~n7800 & ~n7802;
  assign n7804 = pi647 & n7803;
  assign n7805 = ~pi647 & n7561;
  assign n7806 = pi1157 & ~n7805;
  assign n7807 = ~n7804 & n7806;
  assign n7808 = ~pi630 & ~n7807;
  assign n7809 = ~n7799 & n7808;
  assign n7810 = pi647 & ~n7788;
  assign n7811 = ~pi647 & ~n7796;
  assign n7812 = pi1157 & ~n7811;
  assign n7813 = ~n7810 & n7812;
  assign n7814 = ~pi647 & n7803;
  assign n7815 = pi647 & n7561;
  assign n7816 = ~pi1157 & ~n7815;
  assign n7817 = ~n7814 & n7816;
  assign n7818 = pi630 & ~n7817;
  assign n7819 = ~n7813 & n7818;
  assign n7820 = ~n7809 & ~n7819;
  assign n7821 = pi787 & ~n7820;
  assign n7822 = ~pi787 & ~n7788;
  assign n7823 = ~n7821 & ~n7822;
  assign n7824 = pi644 & ~n7823;
  assign n7825 = ~pi787 & ~n7803;
  assign n7826 = ~n7807 & ~n7817;
  assign n7827 = pi787 & ~n7826;
  assign n7828 = ~n7825 & ~n7827;
  assign n7829 = ~pi644 & n7828;
  assign n7830 = pi715 & ~n7829;
  assign n7831 = ~n7824 & n7830;
  assign n7832 = ~pi630 & pi1157;
  assign n7833 = pi630 & ~pi1157;
  assign n7834 = ~n7832 & ~n7833;
  assign n7835 = pi787 & ~n7834;
  assign n7836 = ~n7796 & ~n7835;
  assign n7837 = n7561 & n7835;
  assign n7838 = ~n7561 & n7835;
  assign n7839 = n7796 & ~n7835;
  assign n7840 = ~n7838 & ~n7839;
  assign n7841 = ~n7836 & ~n7837;
  assign n7842 = pi644 & n59235;
  assign n7843 = ~pi644 & n7561;
  assign n7844 = ~pi715 & ~n7843;
  assign n7845 = ~n7842 & n7844;
  assign n7846 = pi1160 & ~n7845;
  assign n7847 = ~n7831 & n7846;
  assign n7848 = ~pi644 & ~n7823;
  assign n7849 = pi644 & n7828;
  assign n7850 = ~pi715 & ~n7849;
  assign n7851 = ~n7848 & n7850;
  assign n7852 = ~pi644 & n59235;
  assign n7853 = pi644 & n7561;
  assign n7854 = pi715 & ~n7853;
  assign n7855 = ~n7852 & n7854;
  assign n7856 = ~pi1160 & ~n7855;
  assign n7857 = ~n7851 & n7856;
  assign n7858 = pi790 & ~n7857;
  assign n7859 = pi790 & ~n7847;
  assign n7860 = ~n7857 & n7859;
  assign n7861 = ~n7847 & n7858;
  assign n7862 = ~pi790 & n7823;
  assign n7863 = n58992 & ~n7862;
  assign n7864 = ~n59236 & n7863;
  assign n7865 = ~pi140 & ~n58992;
  assign n7866 = ~pi832 & ~n7865;
  assign n7867 = ~n7864 & n7866;
  assign n7868 = pi630 & ~pi647;
  assign n7869 = pi1157 & n7868;
  assign n7870 = ~pi630 & pi647;
  assign n7871 = ~pi1157 & n7870;
  assign n7872 = ~n7869 & ~n7871;
  assign n7873 = ~pi140 & ~n2794;
  assign n7874 = n7793 & ~n7873;
  assign n7875 = n2794 & n7597;
  assign n7876 = ~pi761 & n6822;
  assign n7877 = ~n7873 & ~n7876;
  assign n7878 = ~n7875 & ~n7877;
  assign n7879 = ~pi785 & ~n7878;
  assign n7880 = n2794 & ~n7598;
  assign n7881 = ~n7877 & ~n7880;
  assign n7882 = pi1155 & ~n7881;
  assign n7883 = pi609 & n2794;
  assign n7884 = n7878 & ~n7883;
  assign n7885 = ~pi1155 & ~n7884;
  assign n7886 = ~n7882 & ~n7885;
  assign n7887 = pi785 & ~n7886;
  assign n7888 = ~n7879 & ~n7887;
  assign n7889 = ~pi781 & ~n7888;
  assign n7890 = ~pi618 & n2794;
  assign n7891 = n7888 & ~n7890;
  assign n7892 = pi1154 & ~n7891;
  assign n7893 = pi618 & n2794;
  assign n7894 = n7888 & ~n7893;
  assign n7895 = ~pi1154 & ~n7894;
  assign n7896 = ~n7892 & ~n7895;
  assign n7897 = pi781 & ~n7896;
  assign n7898 = ~n7889 & ~n7897;
  assign n7899 = ~pi789 & ~n7898;
  assign n7900 = pi619 & n7898;
  assign n7901 = ~pi619 & n7873;
  assign n7902 = pi1159 & ~n7901;
  assign n7903 = ~n7900 & n7902;
  assign n7904 = ~pi619 & n7898;
  assign n7905 = pi619 & n7873;
  assign n7906 = ~pi1159 & ~n7905;
  assign n7907 = ~n7904 & n7906;
  assign n7908 = ~n7903 & ~n7907;
  assign n7909 = pi789 & ~n7908;
  assign n7910 = ~n7899 & ~n7909;
  assign n7911 = ~pi626 & pi1158;
  assign n7912 = pi626 & ~pi1158;
  assign n7913 = ~n7911 & ~n7912;
  assign n7914 = n7910 & n7913;
  assign n7915 = n7873 & ~n7913;
  assign n7916 = pi626 & n7910;
  assign n7917 = ~pi626 & n7873;
  assign n7918 = pi1158 & ~n7917;
  assign n7919 = ~n7916 & n7918;
  assign n7920 = ~pi626 & n7910;
  assign n7921 = pi626 & n7873;
  assign n7922 = ~pi1158 & ~n7921;
  assign n7923 = ~n7920 & n7922;
  assign n7924 = ~n7919 & ~n7923;
  assign n7925 = ~n7914 & ~n7915;
  assign n7926 = pi788 & n59237;
  assign n7927 = ~pi788 & n7910;
  assign n7928 = ~pi788 & ~n7910;
  assign n7929 = pi788 & ~n59237;
  assign n7930 = ~n7928 & ~n7929;
  assign n7931 = ~n7926 & ~n7927;
  assign n7932 = ~n7793 & ~n59238;
  assign n7933 = ~n7793 & n59238;
  assign n7934 = n7793 & n7873;
  assign n7935 = ~n7933 & ~n7934;
  assign n7936 = ~n7874 & ~n7932;
  assign n7937 = ~n7872 & n59239;
  assign n7938 = ~pi738 & n7055;
  assign n7939 = ~n7873 & ~n7938;
  assign n7940 = ~pi778 & n7939;
  assign n7941 = ~pi625 & n7938;
  assign n7942 = ~n7939 & ~n7941;
  assign n7943 = pi1153 & ~n7942;
  assign n7944 = ~pi1153 & ~n7873;
  assign n7945 = ~n7941 & n7944;
  assign n7946 = ~n7943 & ~n7945;
  assign n7947 = pi778 & ~n7946;
  assign n7948 = ~n7940 & ~n7947;
  assign n7949 = n2794 & n59229;
  assign n7950 = n7948 & ~n7949;
  assign n7951 = n2794 & n59231;
  assign n7952 = n7950 & ~n7951;
  assign n7953 = n2794 & n7716;
  assign n7954 = n7952 & ~n7953;
  assign n7955 = n2794 & n7762;
  assign n7956 = n7954 & ~n7955;
  assign n7957 = ~pi628 & pi1156;
  assign n7958 = pi628 & ~pi1156;
  assign n7959 = ~n7957 & ~n7958;
  assign n7960 = ~pi628 & ~pi1156;
  assign n7961 = pi628 & pi1156;
  assign n7962 = pi792 & ~n7961;
  assign n7963 = ~n7960 & n7962;
  assign n7964 = pi792 & ~n7960;
  assign n7965 = ~n7961 & n7964;
  assign n7966 = pi792 & ~n7959;
  assign n7967 = n2794 & n59240;
  assign n7968 = n7956 & ~n7967;
  assign n7969 = ~pi647 & n7968;
  assign n7970 = pi647 & n7873;
  assign n7971 = ~pi1157 & ~n7970;
  assign n7972 = ~n7969 & n7971;
  assign n7973 = pi630 & n7972;
  assign n7974 = ~pi647 & ~n7873;
  assign n7975 = pi647 & ~n7968;
  assign n7976 = ~n7974 & ~n7975;
  assign n7977 = n7832 & ~n7976;
  assign n7978 = ~n7973 & ~n7977;
  assign n7979 = ~n7937 & n7978;
  assign n7980 = pi787 & ~n7979;
  assign n7981 = ~pi626 & pi641;
  assign n7982 = pi626 & ~pi641;
  assign n7983 = ~n7981 & ~n7982;
  assign n7984 = ~n7913 & ~n7983;
  assign n7985 = n7954 & n7984;
  assign n7986 = ~n7761 & n59237;
  assign n7987 = ~n7985 & ~n7986;
  assign n7988 = pi788 & ~n7987;
  assign n7989 = ~n6701 & ~n7939;
  assign n7990 = pi625 & n7989;
  assign n7991 = n7877 & ~n7989;
  assign n7992 = ~n7990 & ~n7991;
  assign n7993 = n7944 & ~n7992;
  assign n7994 = ~pi608 & ~n7943;
  assign n7995 = ~n7993 & n7994;
  assign n7996 = pi1153 & n7877;
  assign n7997 = ~n7990 & n7996;
  assign n7998 = pi608 & ~n7945;
  assign n7999 = ~n7997 & n7998;
  assign n8000 = ~n7995 & ~n7999;
  assign n8001 = pi778 & ~n8000;
  assign n8002 = ~pi778 & ~n7991;
  assign n8003 = ~n8001 & ~n8002;
  assign n8004 = ~pi609 & ~n8003;
  assign n8005 = pi609 & n7948;
  assign n8006 = ~pi1155 & ~n8005;
  assign n8007 = ~n8004 & n8006;
  assign n8008 = ~pi660 & ~n7882;
  assign n8009 = ~n8007 & n8008;
  assign n8010 = pi609 & ~n8003;
  assign n8011 = ~pi609 & n7948;
  assign n8012 = pi1155 & ~n8011;
  assign n8013 = ~n8010 & n8012;
  assign n8014 = pi660 & ~n7885;
  assign n8015 = ~n8013 & n8014;
  assign n8016 = ~n8009 & ~n8015;
  assign n8017 = pi785 & ~n8016;
  assign n8018 = ~pi785 & ~n8003;
  assign n8019 = ~n8017 & ~n8018;
  assign n8020 = ~pi618 & ~n8019;
  assign n8021 = pi618 & n7950;
  assign n8022 = ~pi1154 & ~n8021;
  assign n8023 = ~n8020 & n8022;
  assign n8024 = ~pi627 & ~n7892;
  assign n8025 = ~n8023 & n8024;
  assign n8026 = pi618 & ~n8019;
  assign n8027 = ~pi618 & n7950;
  assign n8028 = pi1154 & ~n8027;
  assign n8029 = ~n8026 & n8028;
  assign n8030 = pi627 & ~n7895;
  assign n8031 = ~n8029 & n8030;
  assign n8032 = ~n8025 & ~n8031;
  assign n8033 = pi781 & ~n8032;
  assign n8034 = ~pi781 & ~n8019;
  assign n8035 = ~n8033 & ~n8034;
  assign n8036 = ~pi619 & ~n8035;
  assign n8037 = pi619 & n7952;
  assign n8038 = ~pi1159 & ~n8037;
  assign n8039 = ~n8036 & n8038;
  assign n8040 = ~pi648 & ~n7903;
  assign n8041 = ~n8039 & n8040;
  assign n8042 = pi619 & ~n8035;
  assign n8043 = ~pi619 & n7952;
  assign n8044 = pi1159 & ~n8043;
  assign n8045 = ~n8042 & n8044;
  assign n8046 = pi648 & ~n7907;
  assign n8047 = ~n8045 & n8046;
  assign n8048 = pi789 & ~n8047;
  assign n8049 = pi789 & ~n8041;
  assign n8050 = ~n8047 & n8049;
  assign n8051 = ~n8041 & n8048;
  assign n8052 = ~pi789 & n8035;
  assign n8053 = n7913 & n7983;
  assign n8054 = pi788 & ~n7913;
  assign n8055 = ~n7762 & ~n8054;
  assign n8056 = pi788 & ~n8053;
  assign n8057 = ~n8052 & n59242;
  assign n8058 = ~n59241 & n8057;
  assign n8059 = ~n7988 & ~n8058;
  assign n8060 = pi628 & n8059;
  assign n8061 = ~pi628 & ~n59238;
  assign n8062 = pi1156 & ~n8061;
  assign n8063 = ~n8060 & n8062;
  assign n8064 = pi628 & n2794;
  assign n8065 = ~pi1156 & ~n8064;
  assign n8066 = n7956 & n8065;
  assign n8067 = pi629 & ~n8066;
  assign n8068 = ~n8063 & n8067;
  assign n8069 = ~pi628 & n8059;
  assign n8070 = pi628 & ~n59238;
  assign n8071 = ~pi1156 & ~n8070;
  assign n8072 = ~n8069 & n8071;
  assign n8073 = ~pi628 & n2794;
  assign n8074 = pi1156 & ~n8073;
  assign n8075 = n7956 & n8074;
  assign n8076 = ~pi629 & ~n8075;
  assign n8077 = ~n8072 & n8076;
  assign n8078 = pi792 & ~n8077;
  assign n8079 = ~pi628 & ~n8059;
  assign n8080 = pi628 & n59238;
  assign n8081 = ~pi1156 & ~n8080;
  assign n8082 = ~n8079 & n8081;
  assign n8083 = n7956 & ~n8073;
  assign n8084 = pi1156 & ~n8083;
  assign n8085 = ~pi629 & ~n8084;
  assign n8086 = ~n8082 & n8085;
  assign n8087 = pi628 & ~n8059;
  assign n8088 = ~pi628 & n59238;
  assign n8089 = pi1156 & ~n8088;
  assign n8090 = ~n8087 & n8089;
  assign n8091 = n7956 & ~n8064;
  assign n8092 = ~pi1156 & ~n8091;
  assign n8093 = pi629 & ~n8092;
  assign n8094 = ~n8090 & n8093;
  assign n8095 = ~n8086 & ~n8094;
  assign n8096 = pi792 & ~n8095;
  assign n8097 = ~n8068 & n8078;
  assign n8098 = ~pi792 & ~n8059;
  assign n8099 = ~pi630 & ~pi647;
  assign n8100 = ~pi1157 & n8099;
  assign n8101 = pi630 & pi647;
  assign n8102 = pi1157 & n8101;
  assign n8103 = ~pi647 & pi1157;
  assign n8104 = pi647 & ~pi1157;
  assign n8105 = ~n8103 & ~n8104;
  assign n8106 = n7834 & n8105;
  assign n8107 = ~n8100 & ~n8102;
  assign n8108 = pi787 & ~n59244;
  assign n8109 = ~n8098 & ~n8108;
  assign n8110 = ~n59243 & n8109;
  assign n8111 = ~n59243 & ~n8098;
  assign n8112 = ~pi647 & ~n8111;
  assign n8113 = pi647 & ~n59239;
  assign n8114 = ~pi1157 & ~n8113;
  assign n8115 = ~n8112 & n8114;
  assign n8116 = pi647 & n7968;
  assign n8117 = ~pi647 & n7873;
  assign n8118 = pi1157 & ~n8117;
  assign n8119 = pi1157 & ~n7976;
  assign n8120 = ~n8116 & n8118;
  assign n8121 = ~pi630 & ~n59245;
  assign n8122 = ~n8115 & n8121;
  assign n8123 = pi647 & ~n8111;
  assign n8124 = ~pi647 & ~n59239;
  assign n8125 = pi1157 & ~n8124;
  assign n8126 = ~n8123 & n8125;
  assign n8127 = pi630 & ~n7972;
  assign n8128 = ~n8126 & n8127;
  assign n8129 = ~n8122 & ~n8128;
  assign n8130 = pi787 & ~n8129;
  assign n8131 = ~pi787 & ~n8111;
  assign n8132 = ~n8130 & ~n8131;
  assign n8133 = ~n7980 & ~n8110;
  assign n8134 = pi644 & ~n59246;
  assign n8135 = ~pi787 & ~n7968;
  assign n8136 = ~n7972 & ~n59245;
  assign n8137 = pi787 & ~n8136;
  assign n8138 = ~n8135 & ~n8137;
  assign n8139 = ~pi644 & n8138;
  assign n8140 = pi715 & ~n8139;
  assign n8141 = ~n8134 & n8140;
  assign n8142 = n7835 & ~n7873;
  assign n8143 = ~n7835 & n59239;
  assign n8144 = ~n8142 & ~n8143;
  assign n8145 = pi644 & n8144;
  assign n8146 = ~pi644 & n7873;
  assign n8147 = ~pi715 & ~n8146;
  assign n8148 = ~n8145 & n8147;
  assign n8149 = pi1160 & ~n8148;
  assign n8150 = ~n8141 & n8149;
  assign n8151 = ~pi644 & ~n59246;
  assign n8152 = pi644 & n8138;
  assign n8153 = ~pi715 & ~n8152;
  assign n8154 = ~n8151 & n8153;
  assign n8155 = ~pi644 & n8144;
  assign n8156 = pi644 & n7873;
  assign n8157 = pi715 & ~n8156;
  assign n8158 = ~n8155 & n8157;
  assign n8159 = ~pi1160 & ~n8158;
  assign n8160 = ~n8154 & n8159;
  assign n8161 = ~n8150 & ~n8160;
  assign n8162 = pi790 & ~n8161;
  assign n8163 = ~pi790 & ~n59246;
  assign n8164 = pi832 & ~n8163;
  assign n8165 = ~n8162 & n8164;
  assign po297 = ~n7867 & ~n8165;
  assign n8167 = pi141 & ~n59132;
  assign n8168 = ~pi141 & ~n6863;
  assign n8169 = pi749 & n6865;
  assign n8170 = ~n8168 & ~n8169;
  assign n8171 = pi38 & ~n8170;
  assign n8172 = ~pi749 & n6654;
  assign n8173 = pi141 & n6853;
  assign n8174 = ~n8172 & ~n8173;
  assign n8175 = pi39 & ~n8174;
  assign n8176 = ~pi141 & n59164;
  assign n8177 = pi141 & n6799;
  assign n8178 = pi749 & ~n8177;
  assign n8179 = ~n8176 & n8178;
  assign n8180 = ~pi39 & n59147;
  assign n8181 = ~pi141 & ~pi749;
  assign n8182 = ~n8180 & n8181;
  assign n8183 = ~n8179 & ~n8182;
  assign n8184 = ~pi38 & ~n8183;
  assign n8185 = ~n8175 & n8184;
  assign n8186 = ~n8171 & ~n8185;
  assign n8187 = ~pi706 & ~n8186;
  assign n8188 = ~pi141 & n59177;
  assign n8189 = pi141 & n7111;
  assign n8190 = ~pi749 & ~n8189;
  assign n8191 = ~n8188 & n8190;
  assign n8192 = pi141 & n7188;
  assign n8193 = ~pi141 & ~n59203;
  assign n8194 = pi749 & ~n8193;
  assign n8195 = ~n8192 & n8194;
  assign n8196 = pi39 & ~n8195;
  assign n8197 = ~n8191 & n8196;
  assign n8198 = ~pi141 & n7310;
  assign n8199 = pi141 & n7333;
  assign n8200 = ~pi749 & ~n8199;
  assign n8201 = ~pi749 & ~n8198;
  assign n8202 = ~n8199 & n8201;
  assign n8203 = ~n8198 & n8200;
  assign n8204 = ~pi141 & ~n7339;
  assign n8205 = pi141 & ~n7347;
  assign n8206 = pi749 & ~n8205;
  assign n8207 = ~n8204 & n8206;
  assign n8208 = ~pi39 & ~n8207;
  assign n8209 = ~n59247 & n8208;
  assign n8210 = ~pi38 & ~n8209;
  assign n8211 = ~pi39 & ~n7310;
  assign n8212 = pi39 & ~n59177;
  assign n8213 = ~n8211 & ~n8212;
  assign n8214 = ~pi141 & n8213;
  assign n8215 = pi39 & ~n7111;
  assign n8216 = ~pi39 & ~n7333;
  assign n8217 = ~n8215 & ~n8216;
  assign n8218 = pi141 & n8217;
  assign n8219 = ~pi749 & ~n8218;
  assign n8220 = ~n8214 & n8219;
  assign n8221 = pi39 & ~n8193;
  assign n8222 = ~n8192 & n8221;
  assign n8223 = ~pi39 & ~n8205;
  assign n8224 = ~n8204 & n8223;
  assign n8225 = ~n8222 & ~n8224;
  assign n8226 = pi749 & ~n8225;
  assign n8227 = ~n8220 & ~n8226;
  assign n8228 = ~pi38 & ~n8227;
  assign n8229 = ~n8197 & n8210;
  assign n8230 = ~n6701 & n7546;
  assign n8231 = n59171 & n7056;
  assign n8232 = ~pi39 & n59208;
  assign n8233 = pi38 & ~n59249;
  assign n8234 = n8170 & n8233;
  assign n8235 = pi706 & ~n8234;
  assign n8236 = ~n59248 & n8235;
  assign n8237 = n59132 & ~n8236;
  assign n8238 = n59132 & ~n8187;
  assign n8239 = ~n8236 & n8238;
  assign n8240 = ~n8187 & n8237;
  assign n8241 = ~n8167 & ~n59250;
  assign n8242 = ~pi625 & n8241;
  assign n8243 = n59132 & n8186;
  assign n8244 = ~n8167 & ~n8243;
  assign n8245 = pi625 & n8244;
  assign n8246 = ~pi1153 & ~n8245;
  assign n8247 = ~n8242 & n8246;
  assign n8248 = ~pi39 & n7308;
  assign n8249 = ~n7540 & ~n8248;
  assign n8250 = ~pi141 & n8249;
  assign n8251 = ~pi39 & n7345;
  assign n8252 = pi39 & ~n7537;
  assign n8253 = ~pi39 & ~n7345;
  assign n8254 = pi39 & n7537;
  assign n8255 = ~n8253 & ~n8254;
  assign n8256 = ~n8251 & ~n8252;
  assign n8257 = pi141 & n59251;
  assign n8258 = ~pi38 & ~n8257;
  assign n8259 = ~n8250 & n8258;
  assign n8260 = n7547 & ~n8168;
  assign n8261 = pi706 & ~n8260;
  assign n8262 = ~n8259 & n8261;
  assign n8263 = ~pi141 & ~pi706;
  assign n8264 = ~n7553 & n8263;
  assign n8265 = n59132 & ~n8264;
  assign n8266 = ~n8262 & n8265;
  assign n8267 = ~n8167 & ~n8266;
  assign n8268 = pi625 & n8267;
  assign n8269 = ~pi141 & ~n7560;
  assign n8270 = ~pi625 & n8269;
  assign n8271 = pi1153 & ~n8270;
  assign n8272 = ~n8268 & n8271;
  assign n8273 = ~pi608 & ~n8272;
  assign n8274 = ~n8247 & n8273;
  assign n8275 = pi625 & n8241;
  assign n8276 = ~pi625 & n8244;
  assign n8277 = pi1153 & ~n8276;
  assign n8278 = ~n8275 & n8277;
  assign n8279 = ~pi625 & n8267;
  assign n8280 = pi625 & n8269;
  assign n8281 = ~pi1153 & ~n8280;
  assign n8282 = ~n8279 & n8281;
  assign n8283 = pi608 & ~n8282;
  assign n8284 = ~n8278 & n8283;
  assign n8285 = ~n8274 & ~n8284;
  assign n8286 = pi778 & ~n8285;
  assign n8287 = ~pi778 & n8241;
  assign n8288 = ~pi778 & ~n8241;
  assign n8289 = pi778 & ~n8284;
  assign n8290 = ~n8274 & n8289;
  assign n8291 = ~n8288 & ~n8290;
  assign n8292 = ~n8286 & ~n8287;
  assign n8293 = ~pi609 & n59252;
  assign n8294 = ~pi778 & ~n8267;
  assign n8295 = ~n8272 & ~n8282;
  assign n8296 = pi778 & ~n8295;
  assign n8297 = ~n8294 & ~n8296;
  assign n8298 = pi609 & n8297;
  assign n8299 = ~pi1155 & ~n8298;
  assign n8300 = ~n8293 & n8299;
  assign n8301 = ~n7598 & ~n8269;
  assign n8302 = ~n7597 & ~n8244;
  assign n8303 = pi609 & n8302;
  assign n8304 = ~n8301 & ~n8303;
  assign n8305 = pi1155 & ~n8304;
  assign n8306 = ~pi660 & ~n8305;
  assign n8307 = ~n8300 & n8306;
  assign n8308 = pi609 & n59252;
  assign n8309 = ~pi609 & n8297;
  assign n8310 = pi1155 & ~n8309;
  assign n8311 = ~n8308 & n8310;
  assign n8312 = ~n7610 & ~n8269;
  assign n8313 = ~pi609 & n8302;
  assign n8314 = ~n8312 & ~n8313;
  assign n8315 = ~pi1155 & ~n8314;
  assign n8316 = pi660 & ~n8315;
  assign n8317 = ~n8311 & n8316;
  assign n8318 = ~n8307 & ~n8317;
  assign n8319 = pi785 & ~n8318;
  assign n8320 = ~pi785 & n59252;
  assign n8321 = ~n8319 & ~n8320;
  assign n8322 = ~pi618 & ~n8321;
  assign n8323 = ~n59229 & n8297;
  assign n8324 = n59229 & n8269;
  assign n8325 = n59229 & ~n8269;
  assign n8326 = ~n59229 & ~n8297;
  assign n8327 = ~n8325 & ~n8326;
  assign n8328 = ~n8323 & ~n8324;
  assign n8329 = pi618 & n59253;
  assign n8330 = ~pi1154 & ~n8329;
  assign n8331 = ~n8322 & n8330;
  assign n8332 = n7597 & ~n8269;
  assign n8333 = ~n8302 & ~n8332;
  assign n8334 = ~pi785 & ~n8333;
  assign n8335 = ~n8305 & ~n8315;
  assign n8336 = pi785 & ~n8335;
  assign n8337 = ~n8334 & ~n8336;
  assign n8338 = pi618 & n8337;
  assign n8339 = ~pi618 & n8269;
  assign n8340 = pi1154 & ~n8339;
  assign n8341 = ~n8338 & n8340;
  assign n8342 = ~pi627 & ~n8341;
  assign n8343 = ~n8331 & n8342;
  assign n8344 = pi618 & ~n8321;
  assign n8345 = ~pi618 & n59253;
  assign n8346 = pi1154 & ~n8345;
  assign n8347 = ~n8344 & n8346;
  assign n8348 = ~pi618 & n8337;
  assign n8349 = pi618 & n8269;
  assign n8350 = ~pi1154 & ~n8349;
  assign n8351 = ~n8348 & n8350;
  assign n8352 = pi627 & ~n8351;
  assign n8353 = ~n8347 & n8352;
  assign n8354 = ~n8343 & ~n8353;
  assign n8355 = pi781 & ~n8354;
  assign n8356 = ~pi781 & ~n8321;
  assign n8357 = ~n8355 & ~n8356;
  assign n8358 = ~pi619 & ~n8357;
  assign n8359 = n59231 & ~n8269;
  assign n8360 = ~n59231 & ~n59253;
  assign n8361 = ~n59231 & n59253;
  assign n8362 = n59231 & n8269;
  assign n8363 = ~n8361 & ~n8362;
  assign n8364 = ~n8359 & ~n8360;
  assign n8365 = pi619 & ~n59254;
  assign n8366 = ~pi1159 & ~n8365;
  assign n8367 = ~n8358 & n8366;
  assign n8368 = ~pi781 & ~n8337;
  assign n8369 = ~n8341 & ~n8351;
  assign n8370 = pi781 & ~n8369;
  assign n8371 = ~n8368 & ~n8370;
  assign n8372 = pi619 & n8371;
  assign n8373 = ~pi619 & n8269;
  assign n8374 = pi1159 & ~n8373;
  assign n8375 = ~n8372 & n8374;
  assign n8376 = ~pi648 & ~n8375;
  assign n8377 = ~n8367 & n8376;
  assign n8378 = pi619 & ~n8357;
  assign n8379 = ~pi619 & ~n59254;
  assign n8380 = pi1159 & ~n8379;
  assign n8381 = ~n8378 & n8380;
  assign n8382 = ~pi619 & n8371;
  assign n8383 = pi619 & n8269;
  assign n8384 = ~pi1159 & ~n8383;
  assign n8385 = ~n8382 & n8384;
  assign n8386 = pi648 & ~n8385;
  assign n8387 = ~n8381 & n8386;
  assign n8388 = ~n8377 & ~n8387;
  assign n8389 = pi789 & ~n8388;
  assign n8390 = ~pi789 & ~n8357;
  assign n8391 = ~n8389 & ~n8390;
  assign n8392 = ~pi788 & n8391;
  assign n8393 = ~pi626 & n8391;
  assign n8394 = ~n7716 & ~n59254;
  assign n8395 = n7716 & n8269;
  assign n8396 = n7716 & ~n8269;
  assign n8397 = ~n7716 & n59254;
  assign n8398 = ~n8396 & ~n8397;
  assign n8399 = ~n8394 & ~n8395;
  assign n8400 = pi626 & ~n59255;
  assign n8401 = ~pi641 & ~n8400;
  assign n8402 = ~n8393 & n8401;
  assign n8403 = ~pi789 & ~n8371;
  assign n8404 = ~n8375 & ~n8385;
  assign n8405 = pi789 & ~n8404;
  assign n8406 = ~n8403 & ~n8405;
  assign n8407 = ~pi626 & n8406;
  assign n8408 = pi626 & n8269;
  assign n8409 = ~pi1158 & ~n8408;
  assign n8410 = ~n8407 & n8409;
  assign n8411 = ~n7726 & ~n8410;
  assign n8412 = ~n8402 & ~n8411;
  assign n8413 = pi626 & n8391;
  assign n8414 = ~pi626 & ~n59255;
  assign n8415 = pi641 & ~n8414;
  assign n8416 = ~n8413 & n8415;
  assign n8417 = pi626 & n8406;
  assign n8418 = ~pi626 & n8269;
  assign n8419 = pi1158 & ~n8418;
  assign n8420 = ~n8417 & n8419;
  assign n8421 = ~n7741 & ~n8420;
  assign n8422 = ~n8416 & ~n8421;
  assign n8423 = ~n8412 & ~n8422;
  assign n8424 = pi788 & ~n8423;
  assign n8425 = ~n8392 & ~n8424;
  assign n8426 = ~pi628 & n8425;
  assign n8427 = ~n8410 & ~n8420;
  assign n8428 = pi788 & ~n8427;
  assign n8429 = ~pi788 & ~n8406;
  assign n8430 = ~n8428 & ~n8429;
  assign n8431 = pi628 & n8430;
  assign n8432 = ~pi1156 & ~n8431;
  assign n8433 = ~n8426 & n8432;
  assign n8434 = n7762 & ~n8269;
  assign n8435 = ~n7762 & ~n59255;
  assign n8436 = ~n7762 & n59255;
  assign n8437 = n7762 & n8269;
  assign n8438 = ~n8436 & ~n8437;
  assign n8439 = ~n8434 & ~n8435;
  assign n8440 = pi628 & ~n59256;
  assign n8441 = ~pi628 & n8269;
  assign n8442 = pi1156 & ~n8441;
  assign n8443 = ~n8440 & n8442;
  assign n8444 = ~pi629 & ~n8443;
  assign n8445 = ~n8433 & n8444;
  assign n8446 = pi628 & n8425;
  assign n8447 = ~pi628 & n8430;
  assign n8448 = pi1156 & ~n8447;
  assign n8449 = ~n8446 & n8448;
  assign n8450 = ~pi628 & ~n59256;
  assign n8451 = pi628 & n8269;
  assign n8452 = ~pi1156 & ~n8451;
  assign n8453 = ~n8450 & n8452;
  assign n8454 = pi629 & ~n8453;
  assign n8455 = ~n8449 & n8454;
  assign n8456 = ~n8445 & ~n8455;
  assign n8457 = pi792 & ~n8456;
  assign n8458 = ~pi792 & n8425;
  assign n8459 = ~n8457 & ~n8458;
  assign n8460 = ~pi647 & ~n8459;
  assign n8461 = ~n7793 & n8430;
  assign n8462 = n7793 & n8269;
  assign n8463 = ~n8461 & ~n8462;
  assign n8464 = pi647 & ~n8463;
  assign n8465 = ~pi1157 & ~n8464;
  assign n8466 = ~n8460 & n8465;
  assign n8467 = ~pi792 & n59256;
  assign n8468 = ~n8443 & ~n8453;
  assign n8469 = pi792 & ~n8468;
  assign n8470 = ~n8467 & ~n8469;
  assign n8471 = pi647 & n8470;
  assign n8472 = ~pi647 & n8269;
  assign n8473 = pi1157 & ~n8472;
  assign n8474 = ~n8471 & n8473;
  assign n8475 = ~pi630 & ~n8474;
  assign n8476 = ~n8466 & n8475;
  assign n8477 = pi647 & ~n8459;
  assign n8478 = ~pi647 & ~n8463;
  assign n8479 = pi1157 & ~n8478;
  assign n8480 = ~n8477 & n8479;
  assign n8481 = ~pi647 & n8470;
  assign n8482 = pi647 & n8269;
  assign n8483 = ~pi1157 & ~n8482;
  assign n8484 = ~n8481 & n8483;
  assign n8485 = pi630 & ~n8484;
  assign n8486 = ~n8480 & n8485;
  assign n8487 = ~n8476 & ~n8486;
  assign n8488 = pi787 & ~n8487;
  assign n8489 = ~pi787 & ~n8459;
  assign n8490 = ~n8488 & ~n8489;
  assign n8491 = pi644 & ~n8490;
  assign n8492 = ~pi787 & ~n8470;
  assign n8493 = ~n8474 & ~n8484;
  assign n8494 = pi787 & ~n8493;
  assign n8495 = ~n8492 & ~n8494;
  assign n8496 = ~pi644 & n8495;
  assign n8497 = pi715 & ~n8496;
  assign n8498 = ~n8491 & n8497;
  assign n8499 = ~n7835 & ~n8463;
  assign n8500 = n7835 & n8269;
  assign n8501 = n7835 & ~n8269;
  assign n8502 = ~n7835 & n8463;
  assign n8503 = ~n8501 & ~n8502;
  assign n8504 = ~n8499 & ~n8500;
  assign n8505 = pi644 & n59257;
  assign n8506 = ~pi644 & n8269;
  assign n8507 = ~pi715 & ~n8506;
  assign n8508 = ~n8505 & n8507;
  assign n8509 = pi1160 & ~n8508;
  assign n8510 = ~n8498 & n8509;
  assign n8511 = ~pi644 & ~n8490;
  assign n8512 = pi644 & n8495;
  assign n8513 = ~pi715 & ~n8512;
  assign n8514 = ~n8511 & n8513;
  assign n8515 = ~pi644 & n59257;
  assign n8516 = pi644 & n8269;
  assign n8517 = pi715 & ~n8516;
  assign n8518 = ~n8515 & n8517;
  assign n8519 = ~pi1160 & ~n8518;
  assign n8520 = ~n8514 & n8519;
  assign n8521 = pi790 & ~n8520;
  assign n8522 = pi790 & ~n8510;
  assign n8523 = ~n8520 & n8522;
  assign n8524 = ~n8510 & n8521;
  assign n8525 = ~pi790 & n8490;
  assign n8526 = n58992 & ~n8525;
  assign n8527 = ~n59258 & n8526;
  assign n8528 = ~pi141 & ~n58992;
  assign n8529 = ~pi832 & ~n8528;
  assign n8530 = ~n8527 & n8529;
  assign n8531 = ~pi141 & ~n2794;
  assign n8532 = n7793 & ~n8531;
  assign n8533 = pi749 & n6822;
  assign n8534 = ~n8531 & ~n8533;
  assign n8535 = ~n7875 & ~n8534;
  assign n8536 = ~pi785 & ~n8535;
  assign n8537 = ~n7880 & ~n8534;
  assign n8538 = pi1155 & ~n8537;
  assign n8539 = ~n7883 & n8535;
  assign n8540 = ~pi1155 & ~n8539;
  assign n8541 = ~n8538 & ~n8540;
  assign n8542 = pi785 & ~n8541;
  assign n8543 = ~n8536 & ~n8542;
  assign n8544 = ~pi781 & ~n8543;
  assign n8545 = ~n7890 & n8543;
  assign n8546 = pi1154 & ~n8545;
  assign n8547 = ~n7893 & n8543;
  assign n8548 = ~pi1154 & ~n8547;
  assign n8549 = ~n8546 & ~n8548;
  assign n8550 = pi781 & ~n8549;
  assign n8551 = ~n8544 & ~n8550;
  assign n8552 = ~pi789 & ~n8551;
  assign n8553 = pi619 & n8551;
  assign n8554 = ~pi619 & n8531;
  assign n8555 = pi1159 & ~n8554;
  assign n8556 = ~n8553 & n8555;
  assign n8557 = ~pi619 & n8551;
  assign n8558 = pi619 & n8531;
  assign n8559 = ~pi1159 & ~n8558;
  assign n8560 = ~n8557 & n8559;
  assign n8561 = ~n8556 & ~n8560;
  assign n8562 = pi789 & ~n8561;
  assign n8563 = ~n8552 & ~n8562;
  assign n8564 = n7913 & n8563;
  assign n8565 = ~n7913 & n8531;
  assign n8566 = pi626 & n8563;
  assign n8567 = ~pi626 & n8531;
  assign n8568 = pi1158 & ~n8567;
  assign n8569 = ~n8566 & n8568;
  assign n8570 = ~pi626 & n8563;
  assign n8571 = pi626 & n8531;
  assign n8572 = ~pi1158 & ~n8571;
  assign n8573 = ~n8570 & n8572;
  assign n8574 = ~n8569 & ~n8573;
  assign n8575 = ~n8564 & ~n8565;
  assign n8576 = pi788 & n59259;
  assign n8577 = ~pi788 & n8563;
  assign n8578 = ~pi788 & ~n8563;
  assign n8579 = pi788 & ~n59259;
  assign n8580 = ~n8578 & ~n8579;
  assign n8581 = ~n8576 & ~n8577;
  assign n8582 = ~n7793 & ~n59260;
  assign n8583 = ~n7793 & n59260;
  assign n8584 = n7793 & n8531;
  assign n8585 = ~n8583 & ~n8584;
  assign n8586 = ~n8532 & ~n8582;
  assign n8587 = ~n7872 & n59261;
  assign n8588 = pi706 & n7055;
  assign n8589 = ~n8531 & ~n8588;
  assign n8590 = ~pi778 & n8589;
  assign n8591 = ~pi625 & n8588;
  assign n8592 = ~n8589 & ~n8591;
  assign n8593 = pi1153 & ~n8592;
  assign n8594 = ~pi1153 & ~n8531;
  assign n8595 = ~n8591 & n8594;
  assign n8596 = ~n8593 & ~n8595;
  assign n8597 = pi778 & ~n8596;
  assign n8598 = ~n8590 & ~n8597;
  assign n8599 = ~n7949 & n8598;
  assign n8600 = ~n7951 & n8599;
  assign n8601 = ~n7953 & n8600;
  assign n8602 = ~n7955 & n8601;
  assign n8603 = ~n7967 & n8602;
  assign n8604 = ~pi647 & n8603;
  assign n8605 = pi647 & n8531;
  assign n8606 = ~pi1157 & ~n8605;
  assign n8607 = ~n8604 & n8606;
  assign n8608 = pi630 & n8607;
  assign n8609 = ~pi647 & ~n8531;
  assign n8610 = pi647 & ~n8603;
  assign n8611 = ~n8609 & ~n8610;
  assign n8612 = n7832 & ~n8611;
  assign n8613 = ~n8608 & ~n8612;
  assign n8614 = ~n8587 & n8613;
  assign n8615 = pi787 & ~n8614;
  assign n8616 = n7984 & n8601;
  assign n8617 = ~n7761 & n59259;
  assign n8618 = ~n8616 & ~n8617;
  assign n8619 = pi788 & ~n8618;
  assign n8620 = ~n6701 & ~n8589;
  assign n8621 = pi625 & n8620;
  assign n8622 = n8534 & ~n8620;
  assign n8623 = ~n8621 & ~n8622;
  assign n8624 = n8594 & ~n8623;
  assign n8625 = ~pi608 & ~n8593;
  assign n8626 = ~n8624 & n8625;
  assign n8627 = pi1153 & n8534;
  assign n8628 = ~n8621 & n8627;
  assign n8629 = pi608 & ~n8595;
  assign n8630 = ~n8628 & n8629;
  assign n8631 = ~n8626 & ~n8630;
  assign n8632 = pi778 & ~n8631;
  assign n8633 = ~pi778 & ~n8622;
  assign n8634 = ~n8632 & ~n8633;
  assign n8635 = ~pi609 & ~n8634;
  assign n8636 = pi609 & n8598;
  assign n8637 = ~pi1155 & ~n8636;
  assign n8638 = ~n8635 & n8637;
  assign n8639 = ~pi660 & ~n8538;
  assign n8640 = ~n8638 & n8639;
  assign n8641 = pi609 & ~n8634;
  assign n8642 = ~pi609 & n8598;
  assign n8643 = pi1155 & ~n8642;
  assign n8644 = ~n8641 & n8643;
  assign n8645 = pi660 & ~n8540;
  assign n8646 = ~n8644 & n8645;
  assign n8647 = ~n8640 & ~n8646;
  assign n8648 = pi785 & ~n8647;
  assign n8649 = ~pi785 & ~n8634;
  assign n8650 = ~n8648 & ~n8649;
  assign n8651 = ~pi618 & ~n8650;
  assign n8652 = pi618 & n8599;
  assign n8653 = ~pi1154 & ~n8652;
  assign n8654 = ~n8651 & n8653;
  assign n8655 = ~pi627 & ~n8546;
  assign n8656 = ~n8654 & n8655;
  assign n8657 = pi618 & ~n8650;
  assign n8658 = ~pi618 & n8599;
  assign n8659 = pi1154 & ~n8658;
  assign n8660 = ~n8657 & n8659;
  assign n8661 = pi627 & ~n8548;
  assign n8662 = ~n8660 & n8661;
  assign n8663 = ~n8656 & ~n8662;
  assign n8664 = pi781 & ~n8663;
  assign n8665 = ~pi781 & ~n8650;
  assign n8666 = ~n8664 & ~n8665;
  assign n8667 = ~pi619 & ~n8666;
  assign n8668 = pi619 & n8600;
  assign n8669 = ~pi1159 & ~n8668;
  assign n8670 = ~n8667 & n8669;
  assign n8671 = ~pi648 & ~n8556;
  assign n8672 = ~n8670 & n8671;
  assign n8673 = pi619 & ~n8666;
  assign n8674 = ~pi619 & n8600;
  assign n8675 = pi1159 & ~n8674;
  assign n8676 = ~n8673 & n8675;
  assign n8677 = pi648 & ~n8560;
  assign n8678 = ~n8676 & n8677;
  assign n8679 = pi789 & ~n8678;
  assign n8680 = pi789 & ~n8672;
  assign n8681 = ~n8678 & n8680;
  assign n8682 = ~n8672 & n8679;
  assign n8683 = ~pi789 & n8666;
  assign n8684 = n59242 & ~n8683;
  assign n8685 = ~n59262 & n8684;
  assign n8686 = ~n8619 & ~n8685;
  assign n8687 = ~pi628 & n8686;
  assign n8688 = pi628 & ~n59260;
  assign n8689 = ~pi1156 & ~n8688;
  assign n8690 = ~n8687 & n8689;
  assign n8691 = n8074 & n8602;
  assign n8692 = ~pi629 & ~n8691;
  assign n8693 = ~n8690 & n8692;
  assign n8694 = pi628 & n8686;
  assign n8695 = ~pi628 & ~n59260;
  assign n8696 = pi1156 & ~n8695;
  assign n8697 = ~n8694 & n8696;
  assign n8698 = n8065 & n8602;
  assign n8699 = pi629 & ~n8698;
  assign n8700 = ~n8697 & n8699;
  assign n8701 = pi792 & ~n8700;
  assign n8702 = ~pi628 & ~n8686;
  assign n8703 = pi628 & n59260;
  assign n8704 = ~pi1156 & ~n8703;
  assign n8705 = ~n8702 & n8704;
  assign n8706 = ~n8073 & n8602;
  assign n8707 = pi1156 & ~n8706;
  assign n8708 = ~pi629 & ~n8707;
  assign n8709 = ~n8705 & n8708;
  assign n8710 = pi628 & ~n8686;
  assign n8711 = ~pi628 & n59260;
  assign n8712 = pi1156 & ~n8711;
  assign n8713 = ~n8710 & n8712;
  assign n8714 = ~n8064 & n8602;
  assign n8715 = ~pi1156 & ~n8714;
  assign n8716 = pi629 & ~n8715;
  assign n8717 = ~n8713 & n8716;
  assign n8718 = ~n8709 & ~n8717;
  assign n8719 = pi792 & ~n8718;
  assign n8720 = ~n8693 & n8701;
  assign n8721 = ~pi792 & ~n8686;
  assign n8722 = ~n8108 & ~n8721;
  assign n8723 = ~n59263 & n8722;
  assign n8724 = ~n59263 & ~n8721;
  assign n8725 = ~pi647 & ~n8724;
  assign n8726 = pi647 & ~n59261;
  assign n8727 = ~pi1157 & ~n8726;
  assign n8728 = ~n8725 & n8727;
  assign n8729 = pi647 & n8603;
  assign n8730 = ~pi647 & n8531;
  assign n8731 = pi1157 & ~n8730;
  assign n8732 = pi1157 & ~n8611;
  assign n8733 = ~n8729 & n8731;
  assign n8734 = ~pi630 & ~n59264;
  assign n8735 = ~n8728 & n8734;
  assign n8736 = pi647 & ~n8724;
  assign n8737 = ~pi647 & ~n59261;
  assign n8738 = pi1157 & ~n8737;
  assign n8739 = ~n8736 & n8738;
  assign n8740 = pi630 & ~n8607;
  assign n8741 = ~n8739 & n8740;
  assign n8742 = ~n8735 & ~n8741;
  assign n8743 = pi787 & ~n8742;
  assign n8744 = ~pi787 & ~n8724;
  assign n8745 = ~n8743 & ~n8744;
  assign n8746 = ~n8615 & ~n8723;
  assign n8747 = pi644 & ~n59265;
  assign n8748 = ~pi787 & ~n8603;
  assign n8749 = ~n8607 & ~n59264;
  assign n8750 = pi787 & ~n8749;
  assign n8751 = ~n8748 & ~n8750;
  assign n8752 = ~pi644 & n8751;
  assign n8753 = pi715 & ~n8752;
  assign n8754 = ~n8747 & n8753;
  assign n8755 = n7835 & ~n8531;
  assign n8756 = ~n7835 & n59261;
  assign n8757 = ~n8755 & ~n8756;
  assign n8758 = pi644 & n8757;
  assign n8759 = ~pi644 & n8531;
  assign n8760 = ~pi715 & ~n8759;
  assign n8761 = ~n8758 & n8760;
  assign n8762 = pi1160 & ~n8761;
  assign n8763 = ~n8754 & n8762;
  assign n8764 = ~pi644 & ~n59265;
  assign n8765 = pi644 & n8751;
  assign n8766 = ~pi715 & ~n8765;
  assign n8767 = ~n8764 & n8766;
  assign n8768 = ~pi644 & n8757;
  assign n8769 = pi644 & n8531;
  assign n8770 = pi715 & ~n8769;
  assign n8771 = ~n8768 & n8770;
  assign n8772 = ~pi1160 & ~n8771;
  assign n8773 = ~n8767 & n8772;
  assign n8774 = ~n8763 & ~n8773;
  assign n8775 = pi790 & ~n8774;
  assign n8776 = ~pi790 & ~n59265;
  assign n8777 = pi832 & ~n8776;
  assign n8778 = ~n8775 & n8777;
  assign po298 = ~n8530 & ~n8778;
  assign n8780 = pi142 & ~n59132;
  assign n8781 = pi142 & ~n59193;
  assign n8782 = ~pi142 & n7144;
  assign n8783 = pi743 & ~n8782;
  assign n8784 = ~n8781 & n8783;
  assign n8785 = pi142 & ~n6899;
  assign n8786 = ~pi142 & ~n7050;
  assign n8787 = ~pi743 & ~n8786;
  assign n8788 = ~n8785 & n8787;
  assign n8789 = pi142 & n6899;
  assign n8790 = ~pi142 & n7050;
  assign n8791 = ~pi743 & ~n8790;
  assign n8792 = ~n8789 & n8791;
  assign n8793 = pi142 & n59193;
  assign n8794 = ~pi142 & ~n7144;
  assign n8795 = pi743 & ~n8794;
  assign n8796 = pi743 & ~n8793;
  assign n8797 = ~n8794 & n8796;
  assign n8798 = ~n8793 & n8795;
  assign n8799 = ~n8792 & ~n59266;
  assign n8800 = ~n8784 & ~n8788;
  assign n8801 = pi735 & n59267;
  assign n8802 = pi142 & n6708;
  assign n8803 = ~pi142 & n59166;
  assign n8804 = pi743 & ~n8803;
  assign n8805 = ~n8802 & n8804;
  assign n8806 = pi142 & ~n6615;
  assign n8807 = ~pi743 & n8806;
  assign n8808 = ~n8802 & ~n8803;
  assign n8809 = pi743 & ~n8808;
  assign n8810 = ~pi743 & ~n8806;
  assign n8811 = ~n8809 & ~n8810;
  assign n8812 = ~n8805 & ~n8807;
  assign n8813 = ~pi735 & ~n59268;
  assign n8814 = pi735 & ~n59267;
  assign n8815 = ~pi735 & n59268;
  assign n8816 = ~n8814 & ~n8815;
  assign n8817 = ~n8801 & ~n8813;
  assign n8818 = n2790 & ~n59269;
  assign n8819 = ~pi142 & n7129;
  assign n8820 = pi142 & ~n7213;
  assign n8821 = pi743 & ~n8820;
  assign n8822 = ~n8819 & n8821;
  assign n8823 = ~pi142 & n7033;
  assign n8824 = pi142 & ~n6910;
  assign n8825 = ~pi743 & ~n8824;
  assign n8826 = ~n8823 & n8825;
  assign n8827 = ~pi142 & ~n7129;
  assign n8828 = pi142 & n7213;
  assign n8829 = pi743 & ~n8828;
  assign n8830 = ~n8827 & n8829;
  assign n8831 = ~pi142 & ~n7033;
  assign n8832 = pi142 & n6910;
  assign n8833 = ~pi743 & ~n8832;
  assign n8834 = ~n8831 & n8833;
  assign n8835 = ~n8830 & ~n8834;
  assign n8836 = ~n8822 & ~n8826;
  assign n8837 = pi735 & n59270;
  assign n8838 = pi142 & ~n59152;
  assign n8839 = ~pi743 & ~n8838;
  assign n8840 = pi142 & ~n6690;
  assign n8841 = pi743 & ~n6815;
  assign n8842 = ~n8840 & n8841;
  assign n8843 = ~n8839 & ~n8842;
  assign n8844 = ~pi735 & ~n8843;
  assign n8845 = pi735 & ~n59270;
  assign n8846 = ~pi735 & n8843;
  assign n8847 = ~n8845 & ~n8846;
  assign n8848 = ~n8837 & ~n8844;
  assign n8849 = ~n2790 & ~n59271;
  assign n8850 = ~n6544 & ~n8849;
  assign n8851 = ~n8818 & n8850;
  assign n8852 = pi142 & ~n6464;
  assign n8853 = pi743 & n6822;
  assign n8854 = pi743 & n6803;
  assign n8855 = n6463 & n8853;
  assign n8856 = ~n8852 & ~n59272;
  assign n8857 = ~pi735 & n8856;
  assign n8858 = pi142 & ~n6468;
  assign n8859 = n58822 & n8853;
  assign n8860 = ~n8858 & ~n8859;
  assign n8861 = ~n59208 & n8860;
  assign n8862 = ~n6461 & ~n8861;
  assign n8863 = pi735 & ~n8862;
  assign n8864 = ~n8852 & n8863;
  assign n8865 = ~n8857 & ~n8864;
  assign n8866 = n6544 & ~n8865;
  assign n8867 = ~pi223 & ~n8866;
  assign n8868 = ~n8851 & n8867;
  assign n8869 = pi142 & ~n7239;
  assign n8870 = ~pi142 & ~n7171;
  assign n8871 = pi743 & ~n8870;
  assign n8872 = ~n8869 & n8871;
  assign n8873 = pi142 & ~n59172;
  assign n8874 = ~pi142 & n7079;
  assign n8875 = ~pi743 & ~n8874;
  assign n8876 = ~n8873 & n8875;
  assign n8877 = pi142 & n7239;
  assign n8878 = ~pi142 & n7171;
  assign n8879 = pi743 & ~n8878;
  assign n8880 = ~n8877 & n8879;
  assign n8881 = ~pi142 & ~n7079;
  assign n8882 = pi142 & n59172;
  assign n8883 = ~pi743 & ~n8882;
  assign n8884 = ~n8881 & n8883;
  assign n8885 = ~n8880 & ~n8884;
  assign n8886 = ~n8872 & ~n8876;
  assign n8887 = pi735 & n59273;
  assign n8888 = pi142 & ~n6512;
  assign n8889 = ~pi743 & ~n8888;
  assign n8890 = pi142 & ~n6740;
  assign n8891 = pi743 & n7167;
  assign n8892 = ~n8890 & n8891;
  assign n8893 = ~n8889 & ~n8892;
  assign n8894 = ~pi735 & ~n8893;
  assign n8895 = pi735 & ~n59273;
  assign n8896 = ~pi735 & n8893;
  assign n8897 = ~n8895 & ~n8896;
  assign n8898 = ~n8887 & ~n8894;
  assign n8899 = ~n2790 & n59274;
  assign n8900 = pi142 & n7230;
  assign n8901 = ~pi142 & n7165;
  assign n8902 = pi743 & ~n8901;
  assign n8903 = ~n8900 & n8902;
  assign n8904 = pi142 & ~n6940;
  assign n8905 = ~pi142 & ~n7086;
  assign n8906 = ~pi743 & ~n8905;
  assign n8907 = ~n8904 & n8906;
  assign n8908 = ~pi142 & ~n7165;
  assign n8909 = pi142 & ~n7230;
  assign n8910 = pi743 & ~n8909;
  assign n8911 = pi743 & ~n8908;
  assign n8912 = ~n8909 & n8911;
  assign n8913 = ~n8908 & n8910;
  assign n8914 = pi142 & n6940;
  assign n8915 = ~pi142 & n7086;
  assign n8916 = ~pi743 & ~n8915;
  assign n8917 = ~n8914 & n8916;
  assign n8918 = ~n59275 & ~n8917;
  assign n8919 = ~n8903 & ~n8907;
  assign n8920 = pi735 & n59276;
  assign n8921 = pi142 & n6729;
  assign n8922 = n6832 & ~n8921;
  assign n8923 = pi743 & ~n8922;
  assign n8924 = pi142 & ~n59149;
  assign n8925 = ~pi743 & n8924;
  assign n8926 = ~pi743 & ~n8924;
  assign n8927 = pi743 & n6832;
  assign n8928 = ~n8921 & n8927;
  assign n8929 = ~n8926 & ~n8928;
  assign n8930 = ~n8923 & ~n8925;
  assign n8931 = ~pi735 & ~n59277;
  assign n8932 = pi735 & ~n59276;
  assign n8933 = ~pi735 & n59277;
  assign n8934 = ~n8932 & ~n8933;
  assign n8935 = ~n8920 & ~n8931;
  assign n8936 = n2790 & n59278;
  assign n8937 = pi223 & ~n8936;
  assign n8938 = ~n8899 & n8937;
  assign n8939 = ~n8868 & ~n8938;
  assign n8940 = ~pi299 & ~n8939;
  assign n8941 = ~n58846 & n59274;
  assign n8942 = n58846 & n59278;
  assign n8943 = pi215 & ~n8942;
  assign n8944 = ~n8941 & n8943;
  assign n8945 = n58846 & ~n59269;
  assign n8946 = ~n58846 & ~n59271;
  assign n8947 = ~n6629 & ~n8946;
  assign n8948 = ~n8945 & n8947;
  assign n8949 = n6629 & ~n8865;
  assign n8950 = ~pi215 & ~n8949;
  assign n8951 = ~n8948 & n8950;
  assign n8952 = ~n8944 & ~n8951;
  assign n8953 = pi299 & ~n8952;
  assign n8954 = pi39 & ~n8953;
  assign n8955 = pi39 & ~n8940;
  assign n8956 = ~n8953 & n8955;
  assign n8957 = ~n8940 & n8954;
  assign n8958 = pi142 & n6677;
  assign n8959 = ~n7305 & n8958;
  assign n8960 = ~pi142 & ~n6796;
  assign n8961 = ~n7343 & n8960;
  assign n8962 = pi299 & ~n8961;
  assign n8963 = ~n8959 & n8962;
  assign n8964 = pi142 & ~n6671;
  assign n8965 = n7300 & n8964;
  assign n8966 = ~pi142 & ~n6791;
  assign n8967 = ~n7341 & n8966;
  assign n8968 = ~pi299 & ~n8967;
  assign n8969 = ~n8965 & n8968;
  assign n8970 = pi743 & ~n8969;
  assign n8971 = ~n8963 & n8970;
  assign n8972 = ~pi142 & n7331;
  assign n8973 = pi142 & ~n7306;
  assign n8974 = ~n6796 & n8973;
  assign n8975 = pi299 & ~n8974;
  assign n8976 = ~n8972 & n8975;
  assign n8977 = ~pi142 & n7323;
  assign n8978 = pi142 & ~n7300;
  assign n8979 = ~n6791 & n8978;
  assign n8980 = ~pi299 & ~n8979;
  assign n8981 = ~n8977 & n8980;
  assign n8982 = ~n8976 & ~n8981;
  assign n8983 = ~pi743 & ~n8982;
  assign n8984 = pi735 & ~n8983;
  assign n8985 = ~n8965 & ~n8967;
  assign n8986 = pi743 & ~n8985;
  assign n8987 = ~pi743 & ~n8979;
  assign n8988 = ~n8977 & n8987;
  assign n8989 = ~pi299 & ~n8988;
  assign n8990 = ~n8986 & n8989;
  assign n8991 = ~n8959 & ~n8961;
  assign n8992 = pi743 & ~n8991;
  assign n8993 = ~pi743 & ~n8974;
  assign n8994 = ~n8972 & n8993;
  assign n8995 = pi299 & ~n8994;
  assign n8996 = pi299 & ~n8992;
  assign n8997 = ~n8994 & n8996;
  assign n8998 = ~n8992 & n8995;
  assign n8999 = ~n8990 & ~n59280;
  assign n9000 = pi735 & ~n8999;
  assign n9001 = ~n8971 & n8984;
  assign n9002 = pi142 & ~n6453;
  assign n9003 = ~pi743 & ~n9002;
  assign n9004 = pi743 & ~n8960;
  assign n9005 = ~n9002 & ~n9004;
  assign n9006 = ~n8960 & ~n9003;
  assign n9007 = ~n8958 & ~n59282;
  assign n9008 = pi299 & ~n9007;
  assign n9009 = pi743 & ~n8966;
  assign n9010 = ~n8964 & n9009;
  assign n9011 = pi142 & ~pi743;
  assign n9012 = ~n6449 & n9011;
  assign n9013 = ~pi299 & ~n9012;
  assign n9014 = ~n9010 & n9013;
  assign n9015 = ~n9008 & ~n9014;
  assign n9016 = ~pi735 & n9015;
  assign n9017 = ~pi39 & ~n9016;
  assign n9018 = ~n59281 & n9017;
  assign n9019 = ~n59279 & ~n9018;
  assign n9020 = ~pi38 & ~n9019;
  assign n9021 = pi39 & pi142;
  assign n9022 = pi38 & ~n9021;
  assign n9023 = pi735 & n7056;
  assign n9024 = pi735 & n7055;
  assign n9025 = n58822 & n9024;
  assign n9026 = ~n6701 & n9025;
  assign n9027 = pi735 & n59208;
  assign n9028 = n58822 & n9023;
  assign n9029 = n8860 & ~n59283;
  assign n9030 = ~pi39 & ~n9029;
  assign n9031 = n9022 & ~n9030;
  assign n9032 = n59132 & ~n9031;
  assign n9033 = ~n9020 & n9032;
  assign n9034 = ~n8780 & ~n9033;
  assign n9035 = pi625 & n9034;
  assign n9036 = n2790 & n59268;
  assign n9037 = ~n2790 & n8843;
  assign n9038 = ~n6544 & ~n9037;
  assign n9039 = ~n9036 & n9038;
  assign n9040 = n6544 & n8856;
  assign n9041 = ~pi223 & ~n9040;
  assign n9042 = ~n9039 & n9041;
  assign n9043 = ~n2790 & ~n8893;
  assign n9044 = n2790 & ~n59277;
  assign n9045 = pi223 & ~n9044;
  assign n9046 = ~n9043 & n9045;
  assign n9047 = ~pi299 & ~n9046;
  assign n9048 = ~n2790 & n8893;
  assign n9049 = n2790 & n59277;
  assign n9050 = pi223 & ~n9049;
  assign n9051 = ~n9048 & n9050;
  assign n9052 = ~n9036 & ~n9037;
  assign n9053 = ~n6544 & ~n9052;
  assign n9054 = n6544 & ~n8856;
  assign n9055 = ~pi223 & ~n9054;
  assign n9056 = ~n9053 & n9055;
  assign n9057 = ~n9051 & ~n9056;
  assign n9058 = ~pi299 & ~n9057;
  assign n9059 = ~n9042 & n9047;
  assign n9060 = n58846 & n59268;
  assign n9061 = ~n58846 & n8843;
  assign n9062 = ~n6629 & ~n9061;
  assign n9063 = ~n9060 & n9062;
  assign n9064 = n6629 & n8856;
  assign n9065 = ~pi215 & ~n9064;
  assign n9066 = ~n9063 & n9065;
  assign n9067 = ~n58846 & ~n8893;
  assign n9068 = n58846 & ~n59277;
  assign n9069 = pi215 & ~n9068;
  assign n9070 = ~n9067 & n9069;
  assign n9071 = pi299 & ~n9070;
  assign n9072 = n58846 & ~n59268;
  assign n9073 = ~n58846 & ~n8843;
  assign n9074 = ~n6629 & ~n9073;
  assign n9075 = ~n9060 & ~n9061;
  assign n9076 = ~n6629 & ~n9075;
  assign n9077 = ~n9072 & n9074;
  assign n9078 = n6629 & ~n8856;
  assign n9079 = ~pi215 & ~n9078;
  assign n9080 = ~n59285 & n9079;
  assign n9081 = ~n58846 & n8893;
  assign n9082 = n58846 & n59277;
  assign n9083 = pi215 & ~n9082;
  assign n9084 = ~n9081 & n9083;
  assign n9085 = ~n9080 & ~n9084;
  assign n9086 = pi299 & ~n9085;
  assign n9087 = ~n9066 & n9071;
  assign n9088 = pi39 & ~n59286;
  assign n9089 = pi39 & ~n59284;
  assign n9090 = ~n59286 & n9089;
  assign n9091 = ~n59284 & n9088;
  assign n9092 = ~pi39 & n9015;
  assign n9093 = ~pi38 & ~n9092;
  assign n9094 = ~n59287 & n9093;
  assign n9095 = ~pi39 & ~n8860;
  assign n9096 = n9022 & ~n9095;
  assign n9097 = n59132 & ~n9096;
  assign n9098 = ~n9094 & n9097;
  assign n9099 = ~n8780 & ~n9098;
  assign n9100 = ~pi625 & n9099;
  assign n9101 = pi1153 & ~n9100;
  assign n9102 = ~n9035 & n9101;
  assign n9103 = pi142 & ~n7423;
  assign n9104 = ~pi142 & ~n7499;
  assign n9105 = ~n9103 & ~n9104;
  assign n9106 = pi735 & ~n9105;
  assign n9107 = ~pi735 & ~n8806;
  assign n9108 = ~n9106 & ~n9107;
  assign n9109 = n2790 & n9108;
  assign n9110 = ~pi142 & n7492;
  assign n9111 = pi142 & n7429;
  assign n9112 = ~n9110 & ~n9111;
  assign n9113 = pi735 & ~n9112;
  assign n9114 = ~pi735 & ~n8838;
  assign n9115 = ~n9113 & ~n9114;
  assign n9116 = ~n2790 & n9115;
  assign n9117 = ~n6544 & ~n9116;
  assign n9118 = ~n9109 & n9117;
  assign n9119 = pi735 & n7054;
  assign n9120 = n6464 & n9119;
  assign n9121 = n6463 & n9024;
  assign n9122 = ~n8852 & ~n59288;
  assign n9123 = n6544 & n9122;
  assign n9124 = ~pi223 & ~n9123;
  assign n9125 = ~n9118 & n9124;
  assign n9126 = ~pi735 & ~n8888;
  assign n9127 = pi142 & ~n7446;
  assign n9128 = ~pi142 & n7168;
  assign n9129 = n7169 & n9128;
  assign n9130 = pi735 & ~n9129;
  assign n9131 = ~n9127 & n9130;
  assign n9132 = ~n9126 & ~n9131;
  assign n9133 = ~n2790 & ~n9132;
  assign n9134 = ~pi735 & ~n8924;
  assign n9135 = pi142 & ~n59214;
  assign n9136 = pi735 & ~n9128;
  assign n9137 = ~n9135 & n9136;
  assign n9138 = ~n9134 & ~n9137;
  assign n9139 = n2790 & ~n9138;
  assign n9140 = pi223 & ~n9139;
  assign n9141 = ~n9133 & n9140;
  assign n9142 = ~pi299 & ~n9141;
  assign n9143 = ~n9125 & n9142;
  assign n9144 = n58846 & n9108;
  assign n9145 = ~n58846 & n9115;
  assign n9146 = ~n6629 & ~n9145;
  assign n9147 = ~n9144 & n9146;
  assign n9148 = n6629 & n9122;
  assign n9149 = ~pi215 & ~n9148;
  assign n9150 = ~n9147 & n9149;
  assign n9151 = ~n58846 & ~n9132;
  assign n9152 = n58846 & ~n9138;
  assign n9153 = pi215 & ~n9152;
  assign n9154 = ~n9151 & n9153;
  assign n9155 = pi299 & ~n9154;
  assign n9156 = ~n9150 & n9155;
  assign n9157 = pi39 & ~n9156;
  assign n9158 = ~n9143 & n9157;
  assign n9159 = ~pi142 & ~n7345;
  assign n9160 = pi142 & n7308;
  assign n9161 = pi735 & ~n9160;
  assign n9162 = pi735 & ~n9159;
  assign n9163 = ~n9160 & n9162;
  assign n9164 = ~n9159 & n9161;
  assign n9165 = pi142 & ~pi735;
  assign n9166 = ~n59147 & n9165;
  assign n9167 = ~n59289 & ~n9166;
  assign n9168 = ~pi39 & ~n9167;
  assign n9169 = ~pi38 & ~n9168;
  assign n9170 = ~n9143 & ~n9156;
  assign n9171 = pi39 & ~n9170;
  assign n9172 = ~pi39 & ~n9166;
  assign n9173 = ~n59289 & n9172;
  assign n9174 = ~n9171 & ~n9173;
  assign n9175 = ~pi38 & ~n9174;
  assign n9176 = ~n9158 & n9169;
  assign n9177 = ~n8858 & ~n9025;
  assign n9178 = ~pi39 & ~n9177;
  assign n9179 = n9022 & ~n9178;
  assign n9180 = n59132 & ~n9179;
  assign n9181 = ~n59290 & n9180;
  assign n9182 = ~n8780 & ~n9181;
  assign n9183 = ~pi625 & n9182;
  assign n9184 = n59132 & ~n7552;
  assign n9185 = pi142 & ~n9184;
  assign n9186 = ~pi38 & ~pi87;
  assign n9187 = ~pi100 & n9186;
  assign n9188 = ~pi38 & n6305;
  assign n9189 = n6307 & n59291;
  assign n9190 = ~pi38 & n59132;
  assign n9191 = n6306 & n9189;
  assign n9192 = ~n58846 & ~n8888;
  assign n9193 = n58846 & ~n8924;
  assign n9194 = pi39 & pi215;
  assign n9195 = pi299 & n9194;
  assign n9196 = ~n9193 & n9195;
  assign n9197 = ~n9192 & n9196;
  assign n9198 = ~n58846 & n59152;
  assign n9199 = n58846 & n6615;
  assign n9200 = ~n6633 & ~n6635;
  assign n9201 = ~n9198 & ~n9199;
  assign n9202 = ~n6629 & ~n59293;
  assign n9203 = n2851 & ~n6637;
  assign n9204 = ~n9202 & n9203;
  assign n9205 = pi39 & ~n9204;
  assign n9206 = ~n6628 & n9205;
  assign n9207 = pi142 & ~n8180;
  assign n9208 = ~n9206 & n9207;
  assign n9209 = pi39 & ~n6628;
  assign n9210 = n9207 & ~n9209;
  assign n9211 = pi215 & ~n9193;
  assign n9212 = ~n9192 & n9211;
  assign n9213 = n58846 & n8806;
  assign n9214 = ~n58846 & n8838;
  assign n9215 = ~n6629 & ~n9214;
  assign n9216 = ~n58846 & ~n8838;
  assign n9217 = n58846 & ~n8806;
  assign n9218 = ~n9216 & ~n9217;
  assign n9219 = ~n6629 & ~n9218;
  assign n9220 = ~n9213 & n9215;
  assign n9221 = n6629 & ~n8852;
  assign n9222 = ~pi215 & ~n9221;
  assign n9223 = ~n59294 & n9222;
  assign n9224 = ~n9212 & ~n9223;
  assign n9225 = pi39 & pi299;
  assign n9226 = ~n9224 & n9225;
  assign n9227 = ~n9210 & ~n9226;
  assign n9228 = ~n9197 & ~n9208;
  assign n9229 = n59292 & ~n59295;
  assign n9230 = ~n9185 & ~n9229;
  assign n9231 = pi625 & n9230;
  assign n9232 = ~pi1153 & ~n9231;
  assign n9233 = ~n9183 & n9232;
  assign n9234 = pi608 & ~n9233;
  assign n9235 = ~n9102 & n9234;
  assign n9236 = ~pi625 & n9034;
  assign n9237 = pi625 & n9099;
  assign n9238 = ~pi1153 & ~n9237;
  assign n9239 = ~n9236 & n9238;
  assign n9240 = pi625 & n9182;
  assign n9241 = ~pi625 & n9230;
  assign n9242 = pi1153 & ~n9241;
  assign n9243 = ~n9240 & n9242;
  assign n9244 = ~pi608 & ~n9243;
  assign n9245 = ~n9239 & n9244;
  assign n9246 = ~n9235 & ~n9245;
  assign n9247 = pi778 & ~n9246;
  assign n9248 = ~pi778 & n9034;
  assign n9249 = ~n9247 & ~n9248;
  assign n9250 = ~pi609 & ~n9249;
  assign n9251 = ~pi778 & ~n9182;
  assign n9252 = ~n9233 & ~n9243;
  assign n9253 = pi778 & ~n9252;
  assign n9254 = ~n9251 & ~n9253;
  assign n9255 = pi609 & n9254;
  assign n9256 = ~pi1155 & ~n9255;
  assign n9257 = ~n9250 & n9256;
  assign n9258 = ~n7598 & ~n9230;
  assign n9259 = ~n7597 & ~n9099;
  assign n9260 = pi609 & n9259;
  assign n9261 = ~n9258 & ~n9260;
  assign n9262 = pi1155 & ~n9261;
  assign n9263 = ~pi660 & ~n9262;
  assign n9264 = ~n9257 & n9263;
  assign n9265 = pi609 & ~n9249;
  assign n9266 = ~pi609 & n9254;
  assign n9267 = pi1155 & ~n9266;
  assign n9268 = ~n9265 & n9267;
  assign n9269 = ~n7610 & ~n9230;
  assign n9270 = ~pi609 & n9259;
  assign n9271 = ~n9269 & ~n9270;
  assign n9272 = ~pi1155 & ~n9271;
  assign n9273 = pi660 & ~n9272;
  assign n9274 = ~n9268 & n9273;
  assign n9275 = ~n9264 & ~n9274;
  assign n9276 = pi785 & ~n9275;
  assign n9277 = ~pi785 & ~n9249;
  assign n9278 = ~n9276 & ~n9277;
  assign n9279 = ~pi618 & ~n9278;
  assign n9280 = ~n59229 & ~n9254;
  assign n9281 = n59229 & ~n9230;
  assign n9282 = ~n59229 & n9254;
  assign n9283 = n59229 & n9230;
  assign n9284 = ~n9282 & ~n9283;
  assign n9285 = ~n9280 & ~n9281;
  assign n9286 = pi618 & ~n59296;
  assign n9287 = ~pi1154 & ~n9286;
  assign n9288 = ~n9279 & n9287;
  assign n9289 = n7597 & ~n9230;
  assign n9290 = ~n9259 & ~n9289;
  assign n9291 = ~pi785 & ~n9290;
  assign n9292 = ~n9262 & ~n9272;
  assign n9293 = pi785 & ~n9292;
  assign n9294 = ~n9291 & ~n9293;
  assign n9295 = pi618 & n9294;
  assign n9296 = ~pi618 & n9230;
  assign n9297 = pi1154 & ~n9296;
  assign n9298 = ~n9295 & n9297;
  assign n9299 = ~pi627 & ~n9298;
  assign n9300 = ~n9288 & n9299;
  assign n9301 = pi618 & ~n9278;
  assign n9302 = ~pi618 & ~n59296;
  assign n9303 = pi1154 & ~n9302;
  assign n9304 = ~n9301 & n9303;
  assign n9305 = ~pi618 & n9294;
  assign n9306 = pi618 & n9230;
  assign n9307 = ~pi1154 & ~n9306;
  assign n9308 = ~n9305 & n9307;
  assign n9309 = pi627 & ~n9308;
  assign n9310 = ~n9304 & n9309;
  assign n9311 = ~n9300 & ~n9310;
  assign n9312 = pi781 & ~n9311;
  assign n9313 = ~pi781 & ~n9278;
  assign n9314 = ~n9312 & ~n9313;
  assign n9315 = ~pi619 & ~n9314;
  assign n9316 = ~n59231 & ~n59296;
  assign n9317 = n59231 & n9230;
  assign n9318 = n59231 & ~n9230;
  assign n9319 = ~n59231 & n59296;
  assign n9320 = ~n9318 & ~n9319;
  assign n9321 = ~n9316 & ~n9317;
  assign n9322 = pi619 & n59297;
  assign n9323 = ~pi1159 & ~n9322;
  assign n9324 = ~n9315 & n9323;
  assign n9325 = ~pi781 & ~n9294;
  assign n9326 = ~n9298 & ~n9308;
  assign n9327 = pi781 & ~n9326;
  assign n9328 = ~n9325 & ~n9327;
  assign n9329 = pi619 & n9328;
  assign n9330 = ~pi619 & n9230;
  assign n9331 = pi1159 & ~n9330;
  assign n9332 = ~n9329 & n9331;
  assign n9333 = ~pi648 & ~n9332;
  assign n9334 = ~n9324 & n9333;
  assign n9335 = pi619 & ~n9314;
  assign n9336 = ~pi619 & n59297;
  assign n9337 = pi1159 & ~n9336;
  assign n9338 = ~n9335 & n9337;
  assign n9339 = ~pi619 & n9328;
  assign n9340 = pi619 & n9230;
  assign n9341 = ~pi1159 & ~n9340;
  assign n9342 = ~n9339 & n9341;
  assign n9343 = pi648 & ~n9342;
  assign n9344 = ~n9338 & n9343;
  assign n9345 = ~n9334 & ~n9344;
  assign n9346 = pi789 & ~n9345;
  assign n9347 = ~pi789 & ~n9314;
  assign n9348 = ~n9346 & ~n9347;
  assign n9349 = ~pi788 & n9348;
  assign n9350 = ~pi626 & n9348;
  assign n9351 = n7716 & ~n9230;
  assign n9352 = ~n7716 & ~n59297;
  assign n9353 = ~n7716 & n59297;
  assign n9354 = n7716 & n9230;
  assign n9355 = ~n9353 & ~n9354;
  assign n9356 = ~n9351 & ~n9352;
  assign n9357 = pi626 & n59298;
  assign n9358 = ~pi641 & ~n9357;
  assign n9359 = ~n9350 & n9358;
  assign n9360 = ~pi789 & ~n9328;
  assign n9361 = ~n9332 & ~n9342;
  assign n9362 = pi789 & ~n9361;
  assign n9363 = ~n9360 & ~n9362;
  assign n9364 = ~pi626 & n9363;
  assign n9365 = pi626 & n9230;
  assign n9366 = ~pi1158 & ~n9365;
  assign n9367 = ~n9364 & n9366;
  assign n9368 = ~n7726 & ~n9367;
  assign n9369 = ~n9359 & ~n9368;
  assign n9370 = pi626 & n9348;
  assign n9371 = ~pi626 & n59298;
  assign n9372 = pi641 & ~n9371;
  assign n9373 = ~n9370 & n9372;
  assign n9374 = pi626 & n9363;
  assign n9375 = ~pi626 & n9230;
  assign n9376 = pi1158 & ~n9375;
  assign n9377 = ~n9374 & n9376;
  assign n9378 = ~n7741 & ~n9377;
  assign n9379 = ~n9373 & ~n9378;
  assign n9380 = ~n9369 & ~n9379;
  assign n9381 = pi788 & ~n9380;
  assign n9382 = ~n9349 & ~n9381;
  assign n9383 = ~pi628 & n9382;
  assign n9384 = ~n9367 & ~n9377;
  assign n9385 = pi788 & ~n9384;
  assign n9386 = ~pi788 & ~n9363;
  assign n9387 = ~n9385 & ~n9386;
  assign n9388 = pi628 & n9387;
  assign n9389 = ~pi1156 & ~n9388;
  assign n9390 = ~n9383 & n9389;
  assign n9391 = ~n7762 & n59298;
  assign n9392 = n7762 & ~n9230;
  assign n9393 = ~n7762 & ~n59298;
  assign n9394 = n7762 & n9230;
  assign n9395 = ~n9393 & ~n9394;
  assign n9396 = ~n9391 & ~n9392;
  assign n9397 = pi628 & ~n59299;
  assign n9398 = ~pi628 & n9230;
  assign n9399 = pi1156 & ~n9398;
  assign n9400 = ~n9397 & n9399;
  assign n9401 = ~pi629 & ~n9400;
  assign n9402 = ~n9390 & n9401;
  assign n9403 = pi628 & n9382;
  assign n9404 = ~pi628 & n9387;
  assign n9405 = pi1156 & ~n9404;
  assign n9406 = ~n9403 & n9405;
  assign n9407 = ~pi628 & ~n59299;
  assign n9408 = pi628 & n9230;
  assign n9409 = ~pi1156 & ~n9408;
  assign n9410 = ~n9407 & n9409;
  assign n9411 = pi629 & ~n9410;
  assign n9412 = ~n9406 & n9411;
  assign n9413 = ~n9402 & ~n9412;
  assign n9414 = pi792 & ~n9413;
  assign n9415 = ~pi792 & n9382;
  assign n9416 = ~n9414 & ~n9415;
  assign n9417 = ~pi647 & ~n9416;
  assign n9418 = ~n7793 & ~n9387;
  assign n9419 = n7793 & ~n9230;
  assign n9420 = ~n7793 & n9387;
  assign n9421 = n7793 & n9230;
  assign n9422 = ~n9420 & ~n9421;
  assign n9423 = ~n9418 & ~n9419;
  assign n9424 = pi647 & ~n59300;
  assign n9425 = ~pi1157 & ~n9424;
  assign n9426 = ~n9417 & n9425;
  assign n9427 = ~pi792 & n59299;
  assign n9428 = ~n9400 & ~n9410;
  assign n9429 = pi792 & ~n9428;
  assign n9430 = ~n9427 & ~n9429;
  assign n9431 = pi647 & n9430;
  assign n9432 = ~pi647 & n9230;
  assign n9433 = pi1157 & ~n9432;
  assign n9434 = ~n9431 & n9433;
  assign n9435 = ~pi630 & ~n9434;
  assign n9436 = ~n9426 & n9435;
  assign n9437 = pi647 & ~n9416;
  assign n9438 = ~pi647 & ~n59300;
  assign n9439 = pi1157 & ~n9438;
  assign n9440 = ~n9437 & n9439;
  assign n9441 = ~pi647 & n9430;
  assign n9442 = pi647 & n9230;
  assign n9443 = ~pi1157 & ~n9442;
  assign n9444 = ~n9441 & n9443;
  assign n9445 = pi630 & ~n9444;
  assign n9446 = ~n9440 & n9445;
  assign n9447 = ~n9436 & ~n9446;
  assign n9448 = pi787 & ~n9447;
  assign n9449 = ~pi787 & ~n9416;
  assign n9450 = ~n9448 & ~n9449;
  assign n9451 = pi644 & ~n9450;
  assign n9452 = ~pi787 & ~n9430;
  assign n9453 = ~n9434 & ~n9444;
  assign n9454 = pi787 & ~n9453;
  assign n9455 = ~n9452 & ~n9454;
  assign n9456 = ~pi644 & n9455;
  assign n9457 = pi715 & ~n9456;
  assign n9458 = ~n9451 & n9457;
  assign n9459 = ~n7835 & ~n59300;
  assign n9460 = n7835 & n9230;
  assign n9461 = n7835 & ~n9230;
  assign n9462 = ~n7835 & n59300;
  assign n9463 = ~n9461 & ~n9462;
  assign n9464 = ~n9459 & ~n9460;
  assign n9465 = pi644 & n59301;
  assign n9466 = ~pi644 & n9230;
  assign n9467 = ~pi715 & ~n9466;
  assign n9468 = ~n9465 & n9467;
  assign n9469 = pi1160 & ~n9468;
  assign n9470 = ~n9458 & n9469;
  assign n9471 = ~pi644 & ~n9450;
  assign n9472 = pi644 & n9455;
  assign n9473 = ~pi715 & ~n9472;
  assign n9474 = ~n9471 & n9473;
  assign n9475 = ~pi644 & n59301;
  assign n9476 = pi644 & n9230;
  assign n9477 = pi715 & ~n9476;
  assign n9478 = ~n9475 & n9477;
  assign n9479 = ~pi1160 & ~n9478;
  assign n9480 = ~n9474 & n9479;
  assign n9481 = pi790 & ~n9480;
  assign n9482 = pi790 & ~n9470;
  assign n9483 = ~n9480 & n9482;
  assign n9484 = ~n9470 & n9481;
  assign n9485 = ~pi790 & n9450;
  assign n9486 = n4441 & ~n9485;
  assign n9487 = ~n59302 & n9486;
  assign n9488 = ~pi142 & ~n4441;
  assign n9489 = ~pi57 & ~n9488;
  assign n9490 = ~n9487 & n9489;
  assign n9491 = pi57 & pi142;
  assign n9492 = ~pi832 & ~n9491;
  assign n9493 = ~n9490 & n9492;
  assign n9494 = ~n7597 & n8853;
  assign n9495 = pi609 & n9494;
  assign n9496 = pi142 & ~n2794;
  assign n9497 = pi1155 & ~n9496;
  assign n9498 = ~n9495 & n9497;
  assign n9499 = ~pi609 & n9494;
  assign n9500 = ~pi1155 & ~n9496;
  assign n9501 = ~n9499 & n9500;
  assign n9502 = ~n9498 & ~n9501;
  assign n9503 = pi785 & ~n9502;
  assign n9504 = ~pi785 & ~n9496;
  assign n9505 = ~n9494 & n9504;
  assign n9506 = ~n9503 & ~n9505;
  assign n9507 = ~pi781 & ~n9506;
  assign n9508 = pi618 & n9506;
  assign n9509 = ~pi618 & n9496;
  assign n9510 = pi1154 & ~n9509;
  assign n9511 = ~n9508 & n9510;
  assign n9512 = ~pi618 & n9506;
  assign n9513 = pi618 & n9496;
  assign n9514 = ~pi1154 & ~n9513;
  assign n9515 = ~n9512 & n9514;
  assign n9516 = ~n9511 & ~n9515;
  assign n9517 = pi781 & ~n9516;
  assign n9518 = ~n9507 & ~n9517;
  assign n9519 = ~pi789 & ~n9518;
  assign n9520 = pi619 & n9518;
  assign n9521 = ~pi619 & n9496;
  assign n9522 = pi1159 & ~n9521;
  assign n9523 = ~n9520 & n9522;
  assign n9524 = ~pi619 & n9518;
  assign n9525 = pi619 & n9496;
  assign n9526 = ~pi1159 & ~n9525;
  assign n9527 = ~n9524 & n9526;
  assign n9528 = ~n9523 & ~n9527;
  assign n9529 = pi789 & ~n9528;
  assign n9530 = ~n9519 & ~n9529;
  assign n9531 = n7913 & n9530;
  assign n9532 = ~n7913 & n9496;
  assign n9533 = pi626 & n9530;
  assign n9534 = ~pi626 & n9496;
  assign n9535 = pi1158 & ~n9534;
  assign n9536 = ~n9533 & n9535;
  assign n9537 = ~pi626 & n9530;
  assign n9538 = pi626 & n9496;
  assign n9539 = ~pi1158 & ~n9538;
  assign n9540 = ~n9537 & n9539;
  assign n9541 = ~n9536 & ~n9540;
  assign n9542 = ~n9531 & ~n9532;
  assign n9543 = ~n7761 & n59303;
  assign n9544 = pi625 & pi1153;
  assign n9545 = ~pi625 & ~pi1153;
  assign n9546 = pi778 & ~n9545;
  assign n9547 = ~pi625 & pi1153;
  assign n9548 = pi625 & ~pi1153;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = pi778 & ~n9549;
  assign n9551 = ~n9544 & n9546;
  assign n9552 = n9024 & ~n59304;
  assign n9553 = ~n9496 & ~n9552;
  assign n9554 = ~n59229 & ~n59231;
  assign n9555 = ~n59229 & ~n9553;
  assign n9556 = ~n59231 & n9555;
  assign n9557 = ~n9553 & n9554;
  assign n9558 = ~n9496 & ~n59305;
  assign n9559 = n7716 & ~n9496;
  assign n9560 = n7984 & ~n9559;
  assign n9561 = ~n9558 & n9560;
  assign n9562 = ~n9543 & ~n9561;
  assign n9563 = pi788 & ~n9562;
  assign n9564 = pi625 & n9023;
  assign n9565 = ~n8853 & ~n9496;
  assign n9566 = ~n9023 & n9565;
  assign n9567 = ~n9564 & ~n9566;
  assign n9568 = ~pi1153 & ~n9567;
  assign n9569 = pi625 & n9024;
  assign n9570 = pi1153 & ~n9496;
  assign n9571 = ~n9569 & n9570;
  assign n9572 = ~pi608 & ~n9571;
  assign n9573 = ~n9568 & n9572;
  assign n9574 = ~n8853 & ~n9564;
  assign n9575 = pi1153 & ~n9574;
  assign n9576 = n9024 & n9545;
  assign n9577 = ~n9496 & ~n9576;
  assign n9578 = ~n9575 & n9577;
  assign n9579 = pi608 & ~n9578;
  assign n9580 = ~n9573 & ~n9579;
  assign n9581 = pi778 & ~n9580;
  assign n9582 = ~pi778 & ~n9566;
  assign n9583 = ~n9581 & ~n9582;
  assign n9584 = ~pi609 & ~n9583;
  assign n9585 = pi609 & ~n9553;
  assign n9586 = ~pi1155 & ~n9585;
  assign n9587 = ~n9584 & n9586;
  assign n9588 = ~pi660 & ~n9498;
  assign n9589 = ~n9587 & n9588;
  assign n9590 = pi609 & ~n9583;
  assign n9591 = ~pi609 & ~n9553;
  assign n9592 = pi1155 & ~n9591;
  assign n9593 = ~n9590 & n9592;
  assign n9594 = pi660 & ~n9501;
  assign n9595 = ~n9593 & n9594;
  assign n9596 = ~n9589 & ~n9595;
  assign n9597 = pi785 & ~n9596;
  assign n9598 = ~pi785 & ~n9583;
  assign n9599 = ~n9597 & ~n9598;
  assign n9600 = ~pi618 & ~n9599;
  assign n9601 = n59229 & ~n9496;
  assign n9602 = ~n9496 & ~n9555;
  assign n9603 = ~n59229 & n9552;
  assign n9604 = ~n9496 & ~n9603;
  assign n9605 = ~n9553 & ~n9601;
  assign n9606 = pi618 & ~n59306;
  assign n9607 = ~pi1154 & ~n9606;
  assign n9608 = ~n9600 & n9607;
  assign n9609 = ~pi627 & ~n9511;
  assign n9610 = ~n9608 & n9609;
  assign n9611 = pi618 & ~n9599;
  assign n9612 = ~pi618 & ~n59306;
  assign n9613 = pi1154 & ~n9612;
  assign n9614 = ~n9611 & n9613;
  assign n9615 = pi627 & ~n9515;
  assign n9616 = ~n9614 & n9615;
  assign n9617 = ~n9610 & ~n9616;
  assign n9618 = pi781 & ~n9617;
  assign n9619 = ~pi781 & ~n9599;
  assign n9620 = ~n9618 & ~n9619;
  assign n9621 = ~pi619 & ~n9620;
  assign n9622 = pi619 & ~n9558;
  assign n9623 = ~pi1159 & ~n9622;
  assign n9624 = ~n9621 & n9623;
  assign n9625 = ~pi648 & ~n9523;
  assign n9626 = ~n9624 & n9625;
  assign n9627 = pi619 & ~n9620;
  assign n9628 = ~pi619 & ~n9558;
  assign n9629 = pi1159 & ~n9628;
  assign n9630 = ~n9627 & n9629;
  assign n9631 = pi648 & ~n9527;
  assign n9632 = ~n9630 & n9631;
  assign n9633 = pi789 & ~n9632;
  assign n9634 = pi789 & ~n9626;
  assign n9635 = ~n9632 & n9634;
  assign n9636 = ~n9626 & n9633;
  assign n9637 = ~pi789 & n9620;
  assign n9638 = n59242 & ~n9637;
  assign n9639 = ~n59307 & n9638;
  assign n9640 = ~n9563 & ~n9639;
  assign n9641 = ~pi628 & ~n9640;
  assign n9642 = pi788 & n59303;
  assign n9643 = ~pi788 & n9530;
  assign n9644 = ~pi788 & ~n9530;
  assign n9645 = pi788 & ~n59303;
  assign n9646 = ~n9644 & ~n9645;
  assign n9647 = ~n9642 & ~n9643;
  assign n9648 = pi628 & n59308;
  assign n9649 = ~pi1156 & ~n9648;
  assign n9650 = ~n9641 & n9649;
  assign n9651 = ~n7716 & ~n7762;
  assign n9652 = n9554 & n9651;
  assign n9653 = n59305 & n9651;
  assign n9654 = ~n9553 & n9652;
  assign n9655 = pi628 & n59309;
  assign n9656 = pi1156 & ~n9496;
  assign n9657 = ~n9655 & n9656;
  assign n9658 = ~pi629 & ~n9657;
  assign n9659 = ~n9650 & n9658;
  assign n9660 = pi628 & ~n9640;
  assign n9661 = ~pi628 & n59308;
  assign n9662 = pi1156 & ~n9661;
  assign n9663 = ~n9660 & n9662;
  assign n9664 = ~pi628 & n59309;
  assign n9665 = ~pi1156 & ~n9496;
  assign n9666 = ~n9664 & n9665;
  assign n9667 = pi629 & ~n9666;
  assign n9668 = ~n9663 & n9667;
  assign n9669 = ~pi628 & n9640;
  assign n9670 = pi628 & ~n59308;
  assign n9671 = ~pi1156 & ~n9670;
  assign n9672 = ~n9669 & n9671;
  assign n9673 = ~n9496 & ~n9655;
  assign n9674 = pi1156 & ~n9673;
  assign n9675 = ~pi629 & ~n9674;
  assign n9676 = ~n9672 & n9675;
  assign n9677 = pi628 & n9640;
  assign n9678 = ~pi628 & ~n59308;
  assign n9679 = pi1156 & ~n9678;
  assign n9680 = ~n9677 & n9679;
  assign n9681 = ~n9496 & ~n9664;
  assign n9682 = ~pi1156 & ~n9681;
  assign n9683 = pi629 & ~n9682;
  assign n9684 = ~n9680 & n9683;
  assign n9685 = ~n9676 & ~n9684;
  assign n9686 = ~n9659 & ~n9668;
  assign n9687 = pi792 & n59310;
  assign n9688 = ~pi792 & ~n9640;
  assign n9689 = pi792 & ~n59310;
  assign n9690 = ~pi792 & n9640;
  assign n9691 = ~n9689 & ~n9690;
  assign n9692 = ~n9687 & ~n9688;
  assign n9693 = ~pi647 & ~n59311;
  assign n9694 = n7793 & ~n9496;
  assign n9695 = ~n7793 & ~n59308;
  assign n9696 = ~n7793 & n59308;
  assign n9697 = n7793 & n9496;
  assign n9698 = ~n9696 & ~n9697;
  assign n9699 = ~n9694 & ~n9695;
  assign n9700 = pi647 & n59312;
  assign n9701 = ~pi1157 & ~n9700;
  assign n9702 = ~n9693 & n9701;
  assign n9703 = ~n59240 & n59309;
  assign n9704 = pi647 & n9703;
  assign n9705 = ~n9496 & ~n9704;
  assign n9706 = pi1157 & ~n9705;
  assign n9707 = ~pi630 & ~n9706;
  assign n9708 = ~n9702 & n9707;
  assign n9709 = pi647 & ~n59311;
  assign n9710 = ~pi647 & n59312;
  assign n9711 = pi1157 & ~n9710;
  assign n9712 = ~n9709 & n9711;
  assign n9713 = ~pi647 & n9703;
  assign n9714 = ~n9496 & ~n9713;
  assign n9715 = ~pi1157 & ~n9714;
  assign n9716 = pi630 & ~n9715;
  assign n9717 = ~n9712 & n9716;
  assign n9718 = ~pi647 & n59311;
  assign n9719 = pi647 & ~n59312;
  assign n9720 = ~pi1157 & ~n9719;
  assign n9721 = ~n9718 & n9720;
  assign n9722 = pi1157 & ~n9496;
  assign n9723 = ~n9704 & n9722;
  assign n9724 = ~pi630 & ~n9723;
  assign n9725 = ~n9721 & n9724;
  assign n9726 = pi647 & n59311;
  assign n9727 = ~pi647 & ~n59312;
  assign n9728 = pi1157 & ~n9727;
  assign n9729 = ~n9726 & n9728;
  assign n9730 = ~pi1157 & ~n9496;
  assign n9731 = ~n9713 & n9730;
  assign n9732 = pi630 & ~n9731;
  assign n9733 = ~n9729 & n9732;
  assign n9734 = ~n9725 & ~n9733;
  assign n9735 = ~n9708 & ~n9717;
  assign n9736 = pi787 & n59313;
  assign n9737 = ~pi787 & ~n59311;
  assign n9738 = pi787 & ~n59313;
  assign n9739 = ~pi787 & n59311;
  assign n9740 = ~n9738 & ~n9739;
  assign n9741 = ~n9736 & ~n9737;
  assign n9742 = pi644 & ~n59314;
  assign n9743 = pi787 & ~n8105;
  assign n9744 = n9703 & ~n9743;
  assign n9745 = ~n9496 & ~n9744;
  assign n9746 = ~pi644 & ~n9745;
  assign n9747 = pi715 & ~n9746;
  assign n9748 = ~n9742 & n9747;
  assign n9749 = ~n7835 & ~n59312;
  assign n9750 = n7835 & n9496;
  assign n9751 = n7835 & ~n9496;
  assign n9752 = ~n7835 & n59312;
  assign n9753 = ~n9751 & ~n9752;
  assign n9754 = ~n9749 & ~n9750;
  assign n9755 = pi644 & n59315;
  assign n9756 = ~pi644 & n9496;
  assign n9757 = ~pi715 & ~n9756;
  assign n9758 = ~n9755 & n9757;
  assign n9759 = pi1160 & ~n9758;
  assign n9760 = ~n9748 & n9759;
  assign n9761 = ~pi644 & ~n59314;
  assign n9762 = pi644 & ~n9745;
  assign n9763 = ~pi715 & ~n9762;
  assign n9764 = ~n9761 & n9763;
  assign n9765 = ~pi644 & n59315;
  assign n9766 = pi644 & n9496;
  assign n9767 = pi715 & ~n9766;
  assign n9768 = ~n9765 & n9767;
  assign n9769 = ~pi1160 & ~n9768;
  assign n9770 = ~n9764 & n9769;
  assign n9771 = ~n9760 & ~n9770;
  assign n9772 = pi790 & ~n9771;
  assign n9773 = ~pi790 & ~n59314;
  assign n9774 = pi832 & ~n9773;
  assign n9775 = ~n9772 & n9774;
  assign po299 = ~n9493 & ~n9775;
  assign n9777 = pi143 & ~n59132;
  assign n9778 = ~pi143 & ~n7553;
  assign n9779 = pi774 & ~n9778;
  assign n9780 = pi38 & n6865;
  assign n9781 = ~pi38 & n6855;
  assign n9782 = pi143 & ~n9781;
  assign n9783 = ~pi38 & ~n59164;
  assign n9784 = ~n6701 & n6863;
  assign n9785 = n6731 & n59171;
  assign n9786 = pi38 & ~n59316;
  assign n9787 = ~n9783 & ~n9786;
  assign n9788 = ~pi143 & ~pi774;
  assign n9789 = n9787 & n9788;
  assign n9790 = ~n9782 & ~n9789;
  assign n9791 = ~n9780 & ~n9790;
  assign n9792 = ~n9779 & ~n9791;
  assign n9793 = ~pi687 & n9792;
  assign n9794 = n6863 & ~n6914;
  assign n9795 = pi38 & n9794;
  assign n9796 = ~pi38 & ~n8213;
  assign n9797 = ~n9795 & ~n9796;
  assign n9798 = ~pi143 & n9797;
  assign n9799 = ~pi38 & n8217;
  assign n9800 = pi143 & n9799;
  assign n9801 = pi38 & n59249;
  assign n9802 = pi774 & ~n9801;
  assign n9803 = ~n9800 & n9802;
  assign n9804 = ~n9798 & n9803;
  assign n9805 = pi39 & ~n7188;
  assign n9806 = ~n6798 & n8253;
  assign n9807 = n6799 & ~n7345;
  assign n9808 = ~n9805 & ~n59317;
  assign n9809 = ~pi38 & ~n9808;
  assign n9810 = pi38 & ~n59207;
  assign n9811 = ~n9809 & ~n9810;
  assign n9812 = pi143 & n9811;
  assign n9813 = ~pi39 & ~n7339;
  assign n9814 = ~pi38 & n9813;
  assign n9815 = pi39 & ~n59203;
  assign n9816 = n6863 & ~n7054;
  assign n9817 = n59171 & n7433;
  assign n9818 = ~pi39 & n7222;
  assign n9819 = ~n6701 & n59318;
  assign n9820 = pi38 & ~n59319;
  assign n9821 = ~n9815 & ~n9820;
  assign n9822 = ~n9814 & ~n9820;
  assign n9823 = ~n9815 & n9822;
  assign n9824 = ~n9814 & n9821;
  assign n9825 = ~pi143 & ~n59320;
  assign n9826 = ~pi774 & ~n9825;
  assign n9827 = ~n9812 & n9826;
  assign n9828 = pi687 & ~n9827;
  assign n9829 = ~n9804 & n9828;
  assign n9830 = n59132 & ~n9829;
  assign n9831 = ~n9793 & n9830;
  assign n9832 = ~n9777 & ~n9831;
  assign n9833 = pi625 & n9832;
  assign n9834 = n59132 & ~n9792;
  assign n9835 = ~n9777 & ~n9834;
  assign n9836 = ~pi625 & n9835;
  assign n9837 = pi1153 & ~n9836;
  assign n9838 = ~n9833 & n9837;
  assign n9839 = ~pi143 & n8249;
  assign n9840 = pi143 & n59251;
  assign n9841 = ~pi38 & ~n9840;
  assign n9842 = ~n9839 & n9841;
  assign n9843 = ~pi143 & ~n6863;
  assign n9844 = n7547 & ~n9843;
  assign n9845 = pi687 & ~n9844;
  assign n9846 = ~n9842 & n9845;
  assign n9847 = ~pi687 & n9778;
  assign n9848 = n59132 & ~n9847;
  assign n9849 = ~n9846 & n9848;
  assign n9850 = ~n9777 & ~n9849;
  assign n9851 = ~pi625 & n9850;
  assign n9852 = ~pi143 & ~n7560;
  assign n9853 = pi625 & n9852;
  assign n9854 = ~pi1153 & ~n9853;
  assign n9855 = ~n9851 & n9854;
  assign n9856 = pi608 & ~n9855;
  assign n9857 = ~n9838 & n9856;
  assign n9858 = ~pi625 & n9832;
  assign n9859 = pi625 & n9835;
  assign n9860 = ~pi1153 & ~n9859;
  assign n9861 = ~n9858 & n9860;
  assign n9862 = pi625 & n9850;
  assign n9863 = ~pi625 & n9852;
  assign n9864 = pi1153 & ~n9863;
  assign n9865 = ~n9862 & n9864;
  assign n9866 = ~pi608 & ~n9865;
  assign n9867 = ~n9861 & n9866;
  assign n9868 = ~n9857 & ~n9867;
  assign n9869 = pi778 & ~n9868;
  assign n9870 = ~pi778 & n9832;
  assign n9871 = ~pi778 & ~n9832;
  assign n9872 = pi778 & ~n9867;
  assign n9873 = ~n9857 & n9872;
  assign n9874 = ~n9871 & ~n9873;
  assign n9875 = ~n9869 & ~n9870;
  assign n9876 = ~pi609 & n59321;
  assign n9877 = ~pi778 & ~n9850;
  assign n9878 = ~n9855 & ~n9865;
  assign n9879 = pi778 & ~n9878;
  assign n9880 = ~n9877 & ~n9879;
  assign n9881 = pi609 & n9880;
  assign n9882 = ~pi1155 & ~n9881;
  assign n9883 = ~n9876 & n9882;
  assign n9884 = ~n7598 & ~n9852;
  assign n9885 = ~n7597 & ~n9835;
  assign n9886 = pi609 & n9885;
  assign n9887 = ~n9884 & ~n9886;
  assign n9888 = pi1155 & ~n9887;
  assign n9889 = ~pi660 & ~n9888;
  assign n9890 = ~n9883 & n9889;
  assign n9891 = pi609 & n59321;
  assign n9892 = ~pi609 & n9880;
  assign n9893 = pi1155 & ~n9892;
  assign n9894 = ~n9891 & n9893;
  assign n9895 = ~n7610 & ~n9852;
  assign n9896 = ~pi609 & n9885;
  assign n9897 = ~n9895 & ~n9896;
  assign n9898 = ~pi1155 & ~n9897;
  assign n9899 = pi660 & ~n9898;
  assign n9900 = ~n9894 & n9899;
  assign n9901 = ~n9890 & ~n9900;
  assign n9902 = pi785 & ~n9901;
  assign n9903 = ~pi785 & n59321;
  assign n9904 = ~n9902 & ~n9903;
  assign n9905 = ~pi618 & ~n9904;
  assign n9906 = ~n59229 & n9880;
  assign n9907 = n59229 & n9852;
  assign n9908 = n59229 & ~n9852;
  assign n9909 = ~n59229 & ~n9880;
  assign n9910 = ~n9908 & ~n9909;
  assign n9911 = ~n9906 & ~n9907;
  assign n9912 = pi618 & n59322;
  assign n9913 = ~pi1154 & ~n9912;
  assign n9914 = ~n9905 & n9913;
  assign n9915 = n7597 & ~n9852;
  assign n9916 = ~n9885 & ~n9915;
  assign n9917 = ~pi785 & ~n9916;
  assign n9918 = ~n9888 & ~n9898;
  assign n9919 = pi785 & ~n9918;
  assign n9920 = ~n9917 & ~n9919;
  assign n9921 = pi618 & n9920;
  assign n9922 = ~pi618 & n9852;
  assign n9923 = pi1154 & ~n9922;
  assign n9924 = ~n9921 & n9923;
  assign n9925 = ~pi627 & ~n9924;
  assign n9926 = ~n9914 & n9925;
  assign n9927 = pi618 & ~n9904;
  assign n9928 = ~pi618 & n59322;
  assign n9929 = pi1154 & ~n9928;
  assign n9930 = ~n9927 & n9929;
  assign n9931 = ~pi618 & n9920;
  assign n9932 = pi618 & n9852;
  assign n9933 = ~pi1154 & ~n9932;
  assign n9934 = ~n9931 & n9933;
  assign n9935 = pi627 & ~n9934;
  assign n9936 = ~n9930 & n9935;
  assign n9937 = ~n9926 & ~n9936;
  assign n9938 = pi781 & ~n9937;
  assign n9939 = ~pi781 & ~n9904;
  assign n9940 = ~n9938 & ~n9939;
  assign n9941 = ~pi619 & ~n9940;
  assign n9942 = n59231 & ~n9852;
  assign n9943 = ~n59231 & ~n59322;
  assign n9944 = ~n59231 & n59322;
  assign n9945 = n59231 & n9852;
  assign n9946 = ~n9944 & ~n9945;
  assign n9947 = ~n9942 & ~n9943;
  assign n9948 = pi619 & ~n59323;
  assign n9949 = ~pi1159 & ~n9948;
  assign n9950 = ~n9941 & n9949;
  assign n9951 = ~pi781 & ~n9920;
  assign n9952 = ~n9924 & ~n9934;
  assign n9953 = pi781 & ~n9952;
  assign n9954 = ~n9951 & ~n9953;
  assign n9955 = pi619 & n9954;
  assign n9956 = ~pi619 & n9852;
  assign n9957 = pi1159 & ~n9956;
  assign n9958 = ~n9955 & n9957;
  assign n9959 = ~pi648 & ~n9958;
  assign n9960 = ~n9950 & n9959;
  assign n9961 = pi619 & ~n9940;
  assign n9962 = ~pi619 & ~n59323;
  assign n9963 = pi1159 & ~n9962;
  assign n9964 = ~n9961 & n9963;
  assign n9965 = ~pi619 & n9954;
  assign n9966 = pi619 & n9852;
  assign n9967 = ~pi1159 & ~n9966;
  assign n9968 = ~n9965 & n9967;
  assign n9969 = pi648 & ~n9968;
  assign n9970 = ~n9964 & n9969;
  assign n9971 = ~n9960 & ~n9970;
  assign n9972 = pi789 & ~n9971;
  assign n9973 = ~pi789 & ~n9940;
  assign n9974 = ~n9972 & ~n9973;
  assign n9975 = ~pi788 & n9974;
  assign n9976 = ~pi626 & n9974;
  assign n9977 = ~n7716 & ~n59323;
  assign n9978 = n7716 & n9852;
  assign n9979 = n7716 & ~n9852;
  assign n9980 = ~n7716 & n59323;
  assign n9981 = ~n9979 & ~n9980;
  assign n9982 = ~n9977 & ~n9978;
  assign n9983 = pi626 & ~n59324;
  assign n9984 = ~pi641 & ~n9983;
  assign n9985 = ~n9976 & n9984;
  assign n9986 = ~pi789 & ~n9954;
  assign n9987 = ~n9958 & ~n9968;
  assign n9988 = pi789 & ~n9987;
  assign n9989 = ~n9986 & ~n9988;
  assign n9990 = ~pi626 & n9989;
  assign n9991 = pi626 & n9852;
  assign n9992 = ~pi1158 & ~n9991;
  assign n9993 = ~n9990 & n9992;
  assign n9994 = ~n7726 & ~n9993;
  assign n9995 = ~n9985 & ~n9994;
  assign n9996 = pi626 & n9974;
  assign n9997 = ~pi626 & ~n59324;
  assign n9998 = pi641 & ~n9997;
  assign n9999 = ~n9996 & n9998;
  assign n10000 = pi626 & n9989;
  assign n10001 = ~pi626 & n9852;
  assign n10002 = pi1158 & ~n10001;
  assign n10003 = ~n10000 & n10002;
  assign n10004 = ~n7741 & ~n10003;
  assign n10005 = ~n9999 & ~n10004;
  assign n10006 = ~n9995 & ~n10005;
  assign n10007 = pi788 & ~n10006;
  assign n10008 = ~n9975 & ~n10007;
  assign n10009 = ~pi628 & n10008;
  assign n10010 = ~n9993 & ~n10003;
  assign n10011 = pi788 & ~n10010;
  assign n10012 = ~pi788 & ~n9989;
  assign n10013 = ~n10011 & ~n10012;
  assign n10014 = pi628 & n10013;
  assign n10015 = ~pi1156 & ~n10014;
  assign n10016 = ~n10009 & n10015;
  assign n10017 = n7762 & ~n9852;
  assign n10018 = ~n7762 & ~n59324;
  assign n10019 = ~n7762 & n59324;
  assign n10020 = n7762 & n9852;
  assign n10021 = ~n10019 & ~n10020;
  assign n10022 = ~n10017 & ~n10018;
  assign n10023 = pi628 & ~n59325;
  assign n10024 = ~pi628 & n9852;
  assign n10025 = pi1156 & ~n10024;
  assign n10026 = ~n10023 & n10025;
  assign n10027 = ~pi629 & ~n10026;
  assign n10028 = ~n10016 & n10027;
  assign n10029 = pi628 & n10008;
  assign n10030 = ~pi628 & n10013;
  assign n10031 = pi1156 & ~n10030;
  assign n10032 = ~n10029 & n10031;
  assign n10033 = ~pi628 & ~n59325;
  assign n10034 = pi628 & n9852;
  assign n10035 = ~pi1156 & ~n10034;
  assign n10036 = ~n10033 & n10035;
  assign n10037 = pi629 & ~n10036;
  assign n10038 = ~n10032 & n10037;
  assign n10039 = ~n10028 & ~n10038;
  assign n10040 = pi792 & ~n10039;
  assign n10041 = ~pi792 & n10008;
  assign n10042 = ~n10040 & ~n10041;
  assign n10043 = ~pi647 & ~n10042;
  assign n10044 = ~n7793 & n10013;
  assign n10045 = n7793 & n9852;
  assign n10046 = ~n10044 & ~n10045;
  assign n10047 = pi647 & ~n10046;
  assign n10048 = ~pi1157 & ~n10047;
  assign n10049 = ~n10043 & n10048;
  assign n10050 = ~pi792 & n59325;
  assign n10051 = ~n10026 & ~n10036;
  assign n10052 = pi792 & ~n10051;
  assign n10053 = ~n10050 & ~n10052;
  assign n10054 = pi647 & n10053;
  assign n10055 = ~pi647 & n9852;
  assign n10056 = pi1157 & ~n10055;
  assign n10057 = ~n10054 & n10056;
  assign n10058 = ~pi630 & ~n10057;
  assign n10059 = ~n10049 & n10058;
  assign n10060 = pi647 & ~n10042;
  assign n10061 = ~pi647 & ~n10046;
  assign n10062 = pi1157 & ~n10061;
  assign n10063 = ~n10060 & n10062;
  assign n10064 = ~pi647 & n10053;
  assign n10065 = pi647 & n9852;
  assign n10066 = ~pi1157 & ~n10065;
  assign n10067 = ~n10064 & n10066;
  assign n10068 = pi630 & ~n10067;
  assign n10069 = ~n10063 & n10068;
  assign n10070 = ~n10059 & ~n10069;
  assign n10071 = pi787 & ~n10070;
  assign n10072 = ~pi787 & ~n10042;
  assign n10073 = ~n10071 & ~n10072;
  assign n10074 = pi644 & ~n10073;
  assign n10075 = ~pi787 & ~n10053;
  assign n10076 = ~n10057 & ~n10067;
  assign n10077 = pi787 & ~n10076;
  assign n10078 = ~n10075 & ~n10077;
  assign n10079 = ~pi644 & n10078;
  assign n10080 = pi715 & ~n10079;
  assign n10081 = ~n10074 & n10080;
  assign n10082 = ~n7835 & ~n10046;
  assign n10083 = n7835 & n9852;
  assign n10084 = n7835 & ~n9852;
  assign n10085 = ~n7835 & n10046;
  assign n10086 = ~n10084 & ~n10085;
  assign n10087 = ~n10082 & ~n10083;
  assign n10088 = pi644 & n59326;
  assign n10089 = ~pi644 & n9852;
  assign n10090 = ~pi715 & ~n10089;
  assign n10091 = ~n10088 & n10090;
  assign n10092 = pi1160 & ~n10091;
  assign n10093 = ~n10081 & n10092;
  assign n10094 = ~pi644 & ~n10073;
  assign n10095 = pi644 & n10078;
  assign n10096 = ~pi715 & ~n10095;
  assign n10097 = ~n10094 & n10096;
  assign n10098 = ~pi644 & n59326;
  assign n10099 = pi644 & n9852;
  assign n10100 = pi715 & ~n10099;
  assign n10101 = ~n10098 & n10100;
  assign n10102 = ~pi1160 & ~n10101;
  assign n10103 = ~n10097 & n10102;
  assign n10104 = pi790 & ~n10103;
  assign n10105 = pi790 & ~n10093;
  assign n10106 = ~n10103 & n10105;
  assign n10107 = ~n10093 & n10104;
  assign n10108 = ~pi790 & n10073;
  assign n10109 = n58992 & ~n10108;
  assign n10110 = ~n59327 & n10109;
  assign n10111 = ~pi143 & ~n58992;
  assign n10112 = ~pi832 & ~n10111;
  assign n10113 = ~n10110 & n10112;
  assign n10114 = ~pi143 & ~n2794;
  assign n10115 = n7793 & ~n10114;
  assign n10116 = ~pi774 & n6822;
  assign n10117 = ~n10114 & ~n10116;
  assign n10118 = ~n7875 & ~n10117;
  assign n10119 = ~pi785 & ~n10118;
  assign n10120 = ~n7880 & ~n10117;
  assign n10121 = pi1155 & ~n10120;
  assign n10122 = ~n7883 & n10118;
  assign n10123 = ~pi1155 & ~n10122;
  assign n10124 = ~n10121 & ~n10123;
  assign n10125 = pi785 & ~n10124;
  assign n10126 = ~n10119 & ~n10125;
  assign n10127 = ~pi781 & ~n10126;
  assign n10128 = ~n7890 & n10126;
  assign n10129 = pi1154 & ~n10128;
  assign n10130 = ~n7893 & n10126;
  assign n10131 = ~pi1154 & ~n10130;
  assign n10132 = ~n10129 & ~n10131;
  assign n10133 = pi781 & ~n10132;
  assign n10134 = ~n10127 & ~n10133;
  assign n10135 = ~pi789 & ~n10134;
  assign n10136 = pi619 & n10134;
  assign n10137 = ~pi619 & n10114;
  assign n10138 = pi1159 & ~n10137;
  assign n10139 = ~n10136 & n10138;
  assign n10140 = ~pi619 & n10134;
  assign n10141 = pi619 & n10114;
  assign n10142 = ~pi1159 & ~n10141;
  assign n10143 = ~n10140 & n10142;
  assign n10144 = ~n10139 & ~n10143;
  assign n10145 = pi789 & ~n10144;
  assign n10146 = ~n10135 & ~n10145;
  assign n10147 = n7913 & n10146;
  assign n10148 = ~n7913 & n10114;
  assign n10149 = pi626 & n10146;
  assign n10150 = ~pi626 & n10114;
  assign n10151 = pi1158 & ~n10150;
  assign n10152 = ~n10149 & n10151;
  assign n10153 = ~pi626 & n10146;
  assign n10154 = pi626 & n10114;
  assign n10155 = ~pi1158 & ~n10154;
  assign n10156 = ~n10153 & n10155;
  assign n10157 = ~n10152 & ~n10156;
  assign n10158 = ~n10147 & ~n10148;
  assign n10159 = pi788 & n59328;
  assign n10160 = ~pi788 & n10146;
  assign n10161 = ~pi788 & ~n10146;
  assign n10162 = pi788 & ~n59328;
  assign n10163 = ~n10161 & ~n10162;
  assign n10164 = ~n10159 & ~n10160;
  assign n10165 = ~n7793 & ~n59329;
  assign n10166 = ~n7793 & n59329;
  assign n10167 = n7793 & n10114;
  assign n10168 = ~n10166 & ~n10167;
  assign n10169 = ~n10115 & ~n10165;
  assign n10170 = ~n7872 & n59330;
  assign n10171 = pi687 & n7055;
  assign n10172 = ~n10114 & ~n10171;
  assign n10173 = ~pi778 & n10172;
  assign n10174 = ~pi625 & n10171;
  assign n10175 = ~n10172 & ~n10174;
  assign n10176 = pi1153 & ~n10175;
  assign n10177 = ~pi1153 & ~n10114;
  assign n10178 = ~n10174 & n10177;
  assign n10179 = ~n10176 & ~n10178;
  assign n10180 = pi778 & ~n10179;
  assign n10181 = ~n10173 & ~n10180;
  assign n10182 = ~n7949 & n10181;
  assign n10183 = ~n7951 & n10182;
  assign n10184 = ~n7953 & n10183;
  assign n10185 = ~n7955 & n10184;
  assign n10186 = ~n7967 & n10185;
  assign n10187 = ~pi647 & n10186;
  assign n10188 = pi647 & n10114;
  assign n10189 = ~pi1157 & ~n10188;
  assign n10190 = ~n10187 & n10189;
  assign n10191 = pi630 & n10190;
  assign n10192 = ~pi647 & ~n10114;
  assign n10193 = pi647 & ~n10186;
  assign n10194 = ~n10192 & ~n10193;
  assign n10195 = n7832 & ~n10194;
  assign n10196 = ~n10191 & ~n10195;
  assign n10197 = ~n10170 & n10196;
  assign n10198 = pi787 & ~n10197;
  assign n10199 = n7984 & n10184;
  assign n10200 = ~n7761 & n59328;
  assign n10201 = ~n10199 & ~n10200;
  assign n10202 = pi788 & ~n10201;
  assign n10203 = ~n6701 & ~n10172;
  assign n10204 = pi625 & n10203;
  assign n10205 = n10117 & ~n10203;
  assign n10206 = ~n10204 & ~n10205;
  assign n10207 = n10177 & ~n10206;
  assign n10208 = ~pi608 & ~n10176;
  assign n10209 = ~n10207 & n10208;
  assign n10210 = pi1153 & n10117;
  assign n10211 = ~n10204 & n10210;
  assign n10212 = pi608 & ~n10178;
  assign n10213 = ~n10211 & n10212;
  assign n10214 = ~n10209 & ~n10213;
  assign n10215 = pi778 & ~n10214;
  assign n10216 = ~pi778 & ~n10205;
  assign n10217 = ~n10215 & ~n10216;
  assign n10218 = ~pi609 & ~n10217;
  assign n10219 = pi609 & n10181;
  assign n10220 = ~pi1155 & ~n10219;
  assign n10221 = ~n10218 & n10220;
  assign n10222 = ~pi660 & ~n10121;
  assign n10223 = ~n10221 & n10222;
  assign n10224 = pi609 & ~n10217;
  assign n10225 = ~pi609 & n10181;
  assign n10226 = pi1155 & ~n10225;
  assign n10227 = ~n10224 & n10226;
  assign n10228 = pi660 & ~n10123;
  assign n10229 = ~n10227 & n10228;
  assign n10230 = ~n10223 & ~n10229;
  assign n10231 = pi785 & ~n10230;
  assign n10232 = ~pi785 & ~n10217;
  assign n10233 = ~n10231 & ~n10232;
  assign n10234 = ~pi618 & ~n10233;
  assign n10235 = pi618 & n10182;
  assign n10236 = ~pi1154 & ~n10235;
  assign n10237 = ~n10234 & n10236;
  assign n10238 = ~pi627 & ~n10129;
  assign n10239 = ~n10237 & n10238;
  assign n10240 = pi618 & ~n10233;
  assign n10241 = ~pi618 & n10182;
  assign n10242 = pi1154 & ~n10241;
  assign n10243 = ~n10240 & n10242;
  assign n10244 = pi627 & ~n10131;
  assign n10245 = ~n10243 & n10244;
  assign n10246 = ~n10239 & ~n10245;
  assign n10247 = pi781 & ~n10246;
  assign n10248 = ~pi781 & ~n10233;
  assign n10249 = ~n10247 & ~n10248;
  assign n10250 = ~pi619 & ~n10249;
  assign n10251 = pi619 & n10183;
  assign n10252 = ~pi1159 & ~n10251;
  assign n10253 = ~n10250 & n10252;
  assign n10254 = ~pi648 & ~n10139;
  assign n10255 = ~n10253 & n10254;
  assign n10256 = pi619 & ~n10249;
  assign n10257 = ~pi619 & n10183;
  assign n10258 = pi1159 & ~n10257;
  assign n10259 = ~n10256 & n10258;
  assign n10260 = pi648 & ~n10143;
  assign n10261 = ~n10259 & n10260;
  assign n10262 = pi789 & ~n10261;
  assign n10263 = pi789 & ~n10255;
  assign n10264 = ~n10261 & n10263;
  assign n10265 = ~n10255 & n10262;
  assign n10266 = ~pi789 & n10249;
  assign n10267 = n59242 & ~n10266;
  assign n10268 = ~n59331 & n10267;
  assign n10269 = ~n10202 & ~n10268;
  assign n10270 = ~pi628 & n10269;
  assign n10271 = pi628 & ~n59329;
  assign n10272 = ~pi1156 & ~n10271;
  assign n10273 = ~n10270 & n10272;
  assign n10274 = n8074 & n10185;
  assign n10275 = ~pi629 & ~n10274;
  assign n10276 = ~n10273 & n10275;
  assign n10277 = pi628 & n10269;
  assign n10278 = ~pi628 & ~n59329;
  assign n10279 = pi1156 & ~n10278;
  assign n10280 = ~n10277 & n10279;
  assign n10281 = n8065 & n10185;
  assign n10282 = pi629 & ~n10281;
  assign n10283 = ~n10280 & n10282;
  assign n10284 = pi792 & ~n10283;
  assign n10285 = ~pi628 & ~n10269;
  assign n10286 = pi628 & n59329;
  assign n10287 = ~pi1156 & ~n10286;
  assign n10288 = ~n10285 & n10287;
  assign n10289 = ~n8073 & n10185;
  assign n10290 = pi1156 & ~n10289;
  assign n10291 = ~pi629 & ~n10290;
  assign n10292 = ~n10288 & n10291;
  assign n10293 = pi628 & ~n10269;
  assign n10294 = ~pi628 & n59329;
  assign n10295 = pi1156 & ~n10294;
  assign n10296 = ~n10293 & n10295;
  assign n10297 = ~n8064 & n10185;
  assign n10298 = ~pi1156 & ~n10297;
  assign n10299 = pi629 & ~n10298;
  assign n10300 = ~n10296 & n10299;
  assign n10301 = ~n10292 & ~n10300;
  assign n10302 = pi792 & ~n10301;
  assign n10303 = ~n10276 & n10284;
  assign n10304 = ~pi792 & ~n10269;
  assign n10305 = ~n8108 & ~n10304;
  assign n10306 = ~n59332 & n10305;
  assign n10307 = ~n59332 & ~n10304;
  assign n10308 = ~pi647 & ~n10307;
  assign n10309 = pi647 & ~n59330;
  assign n10310 = ~pi1157 & ~n10309;
  assign n10311 = ~n10308 & n10310;
  assign n10312 = pi647 & n10186;
  assign n10313 = ~pi647 & n10114;
  assign n10314 = pi1157 & ~n10313;
  assign n10315 = pi1157 & ~n10194;
  assign n10316 = ~n10312 & n10314;
  assign n10317 = ~pi630 & ~n59333;
  assign n10318 = ~n10311 & n10317;
  assign n10319 = pi647 & ~n10307;
  assign n10320 = ~pi647 & ~n59330;
  assign n10321 = pi1157 & ~n10320;
  assign n10322 = ~n10319 & n10321;
  assign n10323 = pi630 & ~n10190;
  assign n10324 = ~n10322 & n10323;
  assign n10325 = ~n10318 & ~n10324;
  assign n10326 = pi787 & ~n10325;
  assign n10327 = ~pi787 & ~n10307;
  assign n10328 = ~n10326 & ~n10327;
  assign n10329 = ~n10198 & ~n10306;
  assign n10330 = pi644 & ~n59334;
  assign n10331 = ~pi787 & ~n10186;
  assign n10332 = ~n10190 & ~n59333;
  assign n10333 = pi787 & ~n10332;
  assign n10334 = ~n10331 & ~n10333;
  assign n10335 = ~pi644 & n10334;
  assign n10336 = pi715 & ~n10335;
  assign n10337 = ~n10330 & n10336;
  assign n10338 = n7835 & ~n10114;
  assign n10339 = ~n7835 & n59330;
  assign n10340 = ~n10338 & ~n10339;
  assign n10341 = pi644 & n10340;
  assign n10342 = ~pi644 & n10114;
  assign n10343 = ~pi715 & ~n10342;
  assign n10344 = ~n10341 & n10343;
  assign n10345 = pi1160 & ~n10344;
  assign n10346 = ~n10337 & n10345;
  assign n10347 = ~pi644 & ~n59334;
  assign n10348 = pi644 & n10334;
  assign n10349 = ~pi715 & ~n10348;
  assign n10350 = ~n10347 & n10349;
  assign n10351 = ~pi644 & n10340;
  assign n10352 = pi644 & n10114;
  assign n10353 = pi715 & ~n10352;
  assign n10354 = ~n10351 & n10353;
  assign n10355 = ~pi1160 & ~n10354;
  assign n10356 = ~n10350 & n10355;
  assign n10357 = ~n10346 & ~n10356;
  assign n10358 = pi790 & ~n10357;
  assign n10359 = ~pi790 & ~n59334;
  assign n10360 = pi832 & ~n10359;
  assign n10361 = ~n10358 & n10360;
  assign po300 = ~n10113 & ~n10361;
  assign n10363 = pi144 & ~n59132;
  assign n10364 = ~pi758 & ~n6654;
  assign n10365 = pi758 & n59163;
  assign n10366 = ~n10364 & ~n10365;
  assign n10367 = pi39 & ~n10366;
  assign n10368 = pi758 & n59157;
  assign n10369 = ~pi758 & n59147;
  assign n10370 = ~pi39 & ~n10369;
  assign n10371 = ~n10368 & n10370;
  assign n10372 = ~n10367 & ~n10371;
  assign n10373 = pi144 & ~n10372;
  assign n10374 = ~pi144 & pi758;
  assign n10375 = n6855 & n10374;
  assign n10376 = ~n10373 & ~n10375;
  assign n10377 = ~pi38 & ~n10376;
  assign n10378 = pi758 & n6701;
  assign n10379 = n6863 & ~n10378;
  assign n10380 = ~pi144 & ~n6863;
  assign n10381 = pi38 & ~n10380;
  assign n10382 = ~n10379 & n10381;
  assign n10383 = ~n10377 & ~n10382;
  assign n10384 = ~pi736 & n10383;
  assign n10385 = pi144 & ~n59177;
  assign n10386 = ~pi144 & ~n7111;
  assign n10387 = ~pi758 & ~n10386;
  assign n10388 = ~n10385 & n10387;
  assign n10389 = ~pi144 & ~n7188;
  assign n10390 = pi144 & n59203;
  assign n10391 = pi758 & ~n10390;
  assign n10392 = ~n10389 & n10391;
  assign n10393 = pi39 & ~n10392;
  assign n10394 = ~n10388 & n10393;
  assign n10395 = ~pi144 & ~n7333;
  assign n10396 = pi144 & ~n7310;
  assign n10397 = ~pi758 & ~n10396;
  assign n10398 = ~pi758 & ~n10395;
  assign n10399 = ~n10396 & n10398;
  assign n10400 = ~n10395 & n10397;
  assign n10401 = pi144 & n7339;
  assign n10402 = ~pi144 & n7347;
  assign n10403 = pi758 & ~n10402;
  assign n10404 = ~n10401 & n10403;
  assign n10405 = ~pi39 & ~n10404;
  assign n10406 = pi144 & ~n7339;
  assign n10407 = ~pi144 & ~n7347;
  assign n10408 = pi758 & ~n10407;
  assign n10409 = ~n10406 & n10408;
  assign n10410 = pi144 & n7310;
  assign n10411 = ~pi144 & n7333;
  assign n10412 = ~pi758 & ~n10411;
  assign n10413 = ~n10410 & n10412;
  assign n10414 = ~n10409 & ~n10413;
  assign n10415 = ~pi39 & ~n10414;
  assign n10416 = ~n59335 & n10405;
  assign n10417 = ~pi38 & ~n59336;
  assign n10418 = ~n10394 & n10417;
  assign n10419 = pi736 & ~n9801;
  assign n10420 = ~n10382 & n10419;
  assign n10421 = ~n10418 & n10420;
  assign n10422 = n59132 & ~n10421;
  assign n10423 = ~n10384 & n10422;
  assign n10424 = ~n10363 & ~n10423;
  assign n10425 = ~pi625 & n10424;
  assign n10426 = n59132 & ~n10383;
  assign n10427 = ~n10363 & ~n10426;
  assign n10428 = pi625 & n10427;
  assign n10429 = ~pi1153 & ~n10428;
  assign n10430 = ~n10425 & n10429;
  assign n10431 = pi736 & n59132;
  assign n10432 = pi38 & ~n59318;
  assign n10433 = ~n10380 & n10432;
  assign n10434 = pi144 & ~n8249;
  assign n10435 = ~pi144 & ~n59251;
  assign n10436 = ~pi38 & ~n10435;
  assign n10437 = ~n10434 & n10436;
  assign n10438 = ~n10433 & ~n10437;
  assign n10439 = n10431 & ~n10438;
  assign n10440 = pi144 & ~n7560;
  assign n10441 = ~n10431 & n10440;
  assign n10442 = ~n10431 & ~n10440;
  assign n10443 = n10431 & ~n10433;
  assign n10444 = ~n10437 & n10443;
  assign n10445 = ~n10442 & ~n10444;
  assign n10446 = ~n10439 & ~n10441;
  assign n10447 = pi625 & ~n59337;
  assign n10448 = ~pi625 & ~n10440;
  assign n10449 = pi1153 & ~n10448;
  assign n10450 = ~n10447 & n10449;
  assign n10451 = ~pi608 & ~n10450;
  assign n10452 = ~n10430 & n10451;
  assign n10453 = pi625 & n10424;
  assign n10454 = ~pi625 & n10427;
  assign n10455 = pi1153 & ~n10454;
  assign n10456 = ~n10453 & n10455;
  assign n10457 = ~pi625 & ~n59337;
  assign n10458 = pi625 & ~n10440;
  assign n10459 = ~pi1153 & ~n10458;
  assign n10460 = ~n10457 & n10459;
  assign n10461 = pi608 & ~n10460;
  assign n10462 = ~n10456 & n10461;
  assign n10463 = ~n10452 & ~n10462;
  assign n10464 = pi778 & ~n10463;
  assign n10465 = ~pi778 & n10424;
  assign n10466 = ~n10464 & ~n10465;
  assign n10467 = ~pi609 & ~n10466;
  assign n10468 = ~pi778 & n59337;
  assign n10469 = ~n10450 & ~n10460;
  assign n10470 = pi778 & ~n10469;
  assign n10471 = ~n10468 & ~n10470;
  assign n10472 = pi609 & n10471;
  assign n10473 = ~pi1155 & ~n10472;
  assign n10474 = ~n10467 & n10473;
  assign n10475 = n7597 & ~n10440;
  assign n10476 = ~n7597 & n10427;
  assign n10477 = ~n7597 & ~n10427;
  assign n10478 = n7597 & n10440;
  assign n10479 = ~n10477 & ~n10478;
  assign n10480 = ~n10475 & ~n10476;
  assign n10481 = pi609 & n59338;
  assign n10482 = ~pi609 & ~n10440;
  assign n10483 = pi1155 & ~n10482;
  assign n10484 = ~n10481 & n10483;
  assign n10485 = ~pi660 & ~n10484;
  assign n10486 = ~n10474 & n10485;
  assign n10487 = pi609 & ~n10466;
  assign n10488 = ~pi609 & n10471;
  assign n10489 = pi1155 & ~n10488;
  assign n10490 = ~n10487 & n10489;
  assign n10491 = ~pi609 & n59338;
  assign n10492 = pi609 & ~n10440;
  assign n10493 = ~pi1155 & ~n10492;
  assign n10494 = ~n10491 & n10493;
  assign n10495 = pi660 & ~n10494;
  assign n10496 = ~n10490 & n10495;
  assign n10497 = ~n10486 & ~n10496;
  assign n10498 = pi785 & ~n10497;
  assign n10499 = ~pi785 & ~n10466;
  assign n10500 = ~n10498 & ~n10499;
  assign n10501 = ~pi618 & ~n10500;
  assign n10502 = ~n59229 & ~n10471;
  assign n10503 = n59229 & n10440;
  assign n10504 = n59229 & ~n10440;
  assign n10505 = ~n59229 & n10471;
  assign n10506 = ~n10504 & ~n10505;
  assign n10507 = ~n10502 & ~n10503;
  assign n10508 = pi618 & ~n59339;
  assign n10509 = ~pi1154 & ~n10508;
  assign n10510 = ~n10501 & n10509;
  assign n10511 = ~pi785 & ~n59338;
  assign n10512 = ~n10484 & ~n10494;
  assign n10513 = pi785 & ~n10512;
  assign n10514 = ~n10511 & ~n10513;
  assign n10515 = pi618 & n10514;
  assign n10516 = ~pi618 & ~n10440;
  assign n10517 = pi1154 & ~n10516;
  assign n10518 = ~n10515 & n10517;
  assign n10519 = ~pi627 & ~n10518;
  assign n10520 = ~n10510 & n10519;
  assign n10521 = pi618 & ~n10500;
  assign n10522 = ~pi618 & ~n59339;
  assign n10523 = pi1154 & ~n10522;
  assign n10524 = ~n10521 & n10523;
  assign n10525 = ~pi618 & n10514;
  assign n10526 = pi618 & ~n10440;
  assign n10527 = ~pi1154 & ~n10526;
  assign n10528 = ~n10525 & n10527;
  assign n10529 = pi627 & ~n10528;
  assign n10530 = ~n10524 & n10529;
  assign n10531 = ~n10520 & ~n10530;
  assign n10532 = pi781 & ~n10531;
  assign n10533 = ~pi781 & ~n10500;
  assign n10534 = ~n10532 & ~n10533;
  assign n10535 = ~pi619 & ~n10534;
  assign n10536 = n59231 & ~n10440;
  assign n10537 = ~n59231 & ~n59339;
  assign n10538 = ~n59231 & n59339;
  assign n10539 = n59231 & n10440;
  assign n10540 = ~n10538 & ~n10539;
  assign n10541 = ~n10536 & ~n10537;
  assign n10542 = pi619 & n59340;
  assign n10543 = ~pi1159 & ~n10542;
  assign n10544 = ~n10535 & n10543;
  assign n10545 = ~pi781 & ~n10514;
  assign n10546 = ~n10518 & ~n10528;
  assign n10547 = pi781 & ~n10546;
  assign n10548 = ~n10545 & ~n10547;
  assign n10549 = pi619 & n10548;
  assign n10550 = ~pi619 & ~n10440;
  assign n10551 = pi1159 & ~n10550;
  assign n10552 = ~n10549 & n10551;
  assign n10553 = ~pi648 & ~n10552;
  assign n10554 = ~n10544 & n10553;
  assign n10555 = pi619 & ~n10534;
  assign n10556 = ~pi619 & n59340;
  assign n10557 = pi1159 & ~n10556;
  assign n10558 = ~n10555 & n10557;
  assign n10559 = ~pi619 & n10548;
  assign n10560 = pi619 & ~n10440;
  assign n10561 = ~pi1159 & ~n10560;
  assign n10562 = ~n10559 & n10561;
  assign n10563 = pi648 & ~n10562;
  assign n10564 = ~n10558 & n10563;
  assign n10565 = ~n10554 & ~n10564;
  assign n10566 = pi789 & ~n10565;
  assign n10567 = ~pi789 & ~n10534;
  assign n10568 = ~n10566 & ~n10567;
  assign n10569 = ~pi788 & n10568;
  assign n10570 = ~pi626 & n10568;
  assign n10571 = ~n7716 & ~n59340;
  assign n10572 = n7716 & n10440;
  assign n10573 = n7716 & ~n10440;
  assign n10574 = ~n7716 & n59340;
  assign n10575 = ~n10573 & ~n10574;
  assign n10576 = ~n10571 & ~n10572;
  assign n10577 = pi626 & n59341;
  assign n10578 = ~pi641 & ~n10577;
  assign n10579 = ~n10570 & n10578;
  assign n10580 = ~pi789 & ~n10548;
  assign n10581 = ~n10552 & ~n10562;
  assign n10582 = pi789 & ~n10581;
  assign n10583 = ~n10580 & ~n10582;
  assign n10584 = ~pi626 & n10583;
  assign n10585 = pi626 & ~n10440;
  assign n10586 = ~pi1158 & ~n10585;
  assign n10587 = ~n10584 & n10586;
  assign n10588 = ~n7726 & ~n10587;
  assign n10589 = ~n10579 & ~n10588;
  assign n10590 = pi626 & n10568;
  assign n10591 = ~pi626 & n59341;
  assign n10592 = pi641 & ~n10591;
  assign n10593 = ~n10590 & n10592;
  assign n10594 = pi626 & n10583;
  assign n10595 = ~pi626 & ~n10440;
  assign n10596 = pi1158 & ~n10595;
  assign n10597 = ~n10594 & n10596;
  assign n10598 = ~n7741 & ~n10597;
  assign n10599 = ~n10593 & ~n10598;
  assign n10600 = ~n10589 & ~n10599;
  assign n10601 = pi788 & ~n10600;
  assign n10602 = ~n10569 & ~n10601;
  assign n10603 = ~pi628 & n10602;
  assign n10604 = ~n10587 & ~n10597;
  assign n10605 = pi788 & ~n10604;
  assign n10606 = ~pi788 & ~n10583;
  assign n10607 = ~n10605 & ~n10606;
  assign n10608 = pi628 & n10607;
  assign n10609 = ~pi1156 & ~n10608;
  assign n10610 = ~n10603 & n10609;
  assign n10611 = n7762 & ~n10440;
  assign n10612 = ~n7762 & ~n59341;
  assign n10613 = ~n7762 & n59341;
  assign n10614 = n7762 & n10440;
  assign n10615 = ~n10613 & ~n10614;
  assign n10616 = ~n10611 & ~n10612;
  assign n10617 = pi628 & n59342;
  assign n10618 = ~pi628 & ~n10440;
  assign n10619 = pi1156 & ~n10618;
  assign n10620 = ~n10617 & n10619;
  assign n10621 = ~pi629 & ~n10620;
  assign n10622 = ~n10610 & n10621;
  assign n10623 = pi628 & n10602;
  assign n10624 = ~pi628 & n10607;
  assign n10625 = pi1156 & ~n10624;
  assign n10626 = ~n10623 & n10625;
  assign n10627 = ~pi628 & n59342;
  assign n10628 = pi628 & ~n10440;
  assign n10629 = ~pi1156 & ~n10628;
  assign n10630 = ~n10627 & n10629;
  assign n10631 = pi629 & ~n10630;
  assign n10632 = ~n10626 & n10631;
  assign n10633 = ~n10622 & ~n10632;
  assign n10634 = pi792 & ~n10633;
  assign n10635 = ~pi792 & n10602;
  assign n10636 = ~n10634 & ~n10635;
  assign n10637 = ~pi647 & ~n10636;
  assign n10638 = ~n7793 & ~n10607;
  assign n10639 = n7793 & n10440;
  assign n10640 = ~n10638 & ~n10639;
  assign n10641 = pi647 & n10640;
  assign n10642 = ~pi1157 & ~n10641;
  assign n10643 = ~n10637 & n10642;
  assign n10644 = ~pi792 & ~n59342;
  assign n10645 = ~n10620 & ~n10630;
  assign n10646 = pi792 & ~n10645;
  assign n10647 = ~n10644 & ~n10646;
  assign n10648 = pi647 & n10647;
  assign n10649 = ~pi647 & ~n10440;
  assign n10650 = pi1157 & ~n10649;
  assign n10651 = ~n10648 & n10650;
  assign n10652 = ~pi630 & ~n10651;
  assign n10653 = ~n10643 & n10652;
  assign n10654 = pi647 & ~n10636;
  assign n10655 = ~pi647 & n10640;
  assign n10656 = pi1157 & ~n10655;
  assign n10657 = ~n10654 & n10656;
  assign n10658 = ~pi647 & n10647;
  assign n10659 = pi647 & ~n10440;
  assign n10660 = ~pi1157 & ~n10659;
  assign n10661 = ~n10658 & n10660;
  assign n10662 = pi630 & ~n10661;
  assign n10663 = ~n10657 & n10662;
  assign n10664 = ~n10653 & ~n10663;
  assign n10665 = pi787 & ~n10664;
  assign n10666 = ~pi787 & ~n10636;
  assign n10667 = ~n10665 & ~n10666;
  assign n10668 = pi644 & ~n10667;
  assign n10669 = ~pi787 & ~n10647;
  assign n10670 = ~n10651 & ~n10661;
  assign n10671 = pi787 & ~n10670;
  assign n10672 = ~n10669 & ~n10671;
  assign n10673 = ~pi644 & n10672;
  assign n10674 = pi715 & ~n10673;
  assign n10675 = ~n10668 & n10674;
  assign n10676 = ~n7835 & ~n10640;
  assign n10677 = n7835 & n10440;
  assign n10678 = n7835 & ~n10440;
  assign n10679 = ~n7835 & n10640;
  assign n10680 = ~n10678 & ~n10679;
  assign n10681 = ~n10676 & ~n10677;
  assign n10682 = pi644 & ~n59343;
  assign n10683 = ~pi644 & ~n10440;
  assign n10684 = ~pi715 & ~n10683;
  assign n10685 = ~n10682 & n10684;
  assign n10686 = pi1160 & ~n10685;
  assign n10687 = ~n10675 & n10686;
  assign n10688 = ~pi644 & ~n10667;
  assign n10689 = pi644 & n10672;
  assign n10690 = ~pi715 & ~n10689;
  assign n10691 = ~n10688 & n10690;
  assign n10692 = ~pi644 & ~n59343;
  assign n10693 = pi644 & ~n10440;
  assign n10694 = pi715 & ~n10693;
  assign n10695 = ~n10692 & n10694;
  assign n10696 = ~pi1160 & ~n10695;
  assign n10697 = ~n10691 & n10696;
  assign n10698 = pi790 & ~n10697;
  assign n10699 = pi790 & ~n10687;
  assign n10700 = ~n10697 & n10699;
  assign n10701 = ~n10687 & n10698;
  assign n10702 = ~pi790 & n10667;
  assign n10703 = n4441 & ~n10702;
  assign n10704 = ~n59344 & n10703;
  assign n10705 = ~pi144 & ~n4441;
  assign n10706 = ~pi57 & ~n10705;
  assign n10707 = ~n10704 & n10706;
  assign n10708 = pi57 & pi144;
  assign n10709 = ~pi832 & ~n10708;
  assign n10710 = ~n10707 & n10709;
  assign n10711 = pi144 & ~n2794;
  assign n10712 = pi736 & n7055;
  assign n10713 = ~n10711 & ~n10712;
  assign n10714 = ~pi778 & n10713;
  assign n10715 = pi625 & n10712;
  assign n10716 = ~n10713 & ~n10715;
  assign n10717 = ~pi1153 & ~n10716;
  assign n10718 = pi1153 & ~n10711;
  assign n10719 = ~n10715 & n10718;
  assign n10720 = ~n10717 & ~n10719;
  assign n10721 = pi778 & ~n10720;
  assign n10722 = ~n10714 & ~n10721;
  assign n10723 = ~n59229 & n10722;
  assign n10724 = ~n59231 & n10723;
  assign n10725 = ~n7716 & n10724;
  assign n10726 = ~n7762 & n10725;
  assign n10727 = n9652 & n10722;
  assign n10728 = ~pi628 & n59345;
  assign n10729 = pi629 & ~n10728;
  assign n10730 = ~pi609 & ~pi1155;
  assign n10731 = pi609 & pi1155;
  assign n10732 = pi785 & ~n10731;
  assign n10733 = pi785 & ~n10730;
  assign n10734 = ~n10731 & n10733;
  assign n10735 = ~n10730 & n10732;
  assign n10736 = pi758 & n6822;
  assign n10737 = ~n59346 & n10736;
  assign n10738 = ~pi619 & pi1159;
  assign n10739 = pi619 & ~pi1159;
  assign n10740 = ~n10738 & ~n10739;
  assign n10741 = pi789 & ~n10740;
  assign n10742 = ~pi618 & ~pi1154;
  assign n10743 = pi618 & pi1154;
  assign n10744 = pi781 & ~n10743;
  assign n10745 = pi781 & ~n10742;
  assign n10746 = ~n10743 & n10745;
  assign n10747 = ~n10742 & n10744;
  assign n10748 = ~n7597 & ~n59347;
  assign n10749 = ~n7597 & ~n10741;
  assign n10750 = ~n59347 & n10749;
  assign n10751 = ~n10741 & n10748;
  assign n10752 = n10737 & n59348;
  assign n10753 = ~n8054 & n10752;
  assign n10754 = pi628 & ~n10753;
  assign n10755 = ~n10729 & ~n10754;
  assign n10756 = ~pi1156 & ~n10755;
  assign n10757 = pi628 & n59345;
  assign n10758 = ~pi628 & ~n10753;
  assign n10759 = pi629 & ~n10758;
  assign n10760 = pi1156 & ~n10759;
  assign n10761 = ~n10757 & n10760;
  assign n10762 = ~n10756 & ~n10761;
  assign n10763 = ~n10711 & ~n10762;
  assign n10764 = pi792 & n10763;
  assign n10765 = ~n10711 & ~n10724;
  assign n10766 = n7716 & ~n10711;
  assign n10767 = ~n10765 & ~n10766;
  assign n10768 = ~n10711 & ~n10725;
  assign n10769 = n7912 & n59349;
  assign n10770 = pi626 & n10752;
  assign n10771 = ~n10711 & ~n10770;
  assign n10772 = pi1158 & ~n10771;
  assign n10773 = ~pi641 & ~n10772;
  assign n10774 = ~n10769 & n10773;
  assign n10775 = n7911 & n59349;
  assign n10776 = ~pi626 & n10752;
  assign n10777 = ~n10711 & ~n10776;
  assign n10778 = ~pi1158 & ~n10777;
  assign n10779 = pi641 & ~n10778;
  assign n10780 = ~n10775 & n10779;
  assign n10781 = pi788 & ~n10780;
  assign n10782 = ~n10774 & n10781;
  assign n10783 = pi736 & n7056;
  assign n10784 = ~n6701 & n10712;
  assign n10785 = ~n10711 & ~n10736;
  assign n10786 = ~n59350 & n10785;
  assign n10787 = pi625 & n59350;
  assign n10788 = ~n6701 & n10715;
  assign n10789 = ~n10786 & ~n59351;
  assign n10790 = ~pi1153 & ~n10789;
  assign n10791 = ~pi608 & ~n10719;
  assign n10792 = ~n10790 & n10791;
  assign n10793 = pi1153 & n10785;
  assign n10794 = n10718 & ~n10736;
  assign n10795 = ~n59351 & n59352;
  assign n10796 = pi608 & ~n10717;
  assign n10797 = ~n10795 & n10796;
  assign n10798 = ~n10792 & ~n10797;
  assign n10799 = pi778 & ~n10798;
  assign n10800 = ~pi778 & ~n10786;
  assign n10801 = ~n10799 & ~n10800;
  assign n10802 = ~pi609 & ~n10801;
  assign n10803 = pi609 & n10722;
  assign n10804 = ~pi1155 & ~n10803;
  assign n10805 = ~n10802 & n10804;
  assign n10806 = n7598 & n10736;
  assign n10807 = pi1155 & ~n10711;
  assign n10808 = ~n10806 & n10807;
  assign n10809 = ~pi660 & ~n10808;
  assign n10810 = ~n10805 & n10809;
  assign n10811 = pi609 & ~n10801;
  assign n10812 = ~pi609 & n10722;
  assign n10813 = pi1155 & ~n10812;
  assign n10814 = ~n10811 & n10813;
  assign n10815 = n7610 & n10736;
  assign n10816 = ~pi1155 & ~n10711;
  assign n10817 = ~n10815 & n10816;
  assign n10818 = pi660 & ~n10817;
  assign n10819 = ~n10814 & n10818;
  assign n10820 = ~n10810 & ~n10819;
  assign n10821 = pi785 & ~n10820;
  assign n10822 = ~pi785 & ~n10801;
  assign n10823 = ~pi618 & n7671;
  assign n10824 = pi627 & n10743;
  assign n10825 = pi781 & ~n10824;
  assign n10826 = ~n10823 & n10825;
  assign n10827 = ~n10822 & ~n10826;
  assign n10828 = ~n10821 & n10827;
  assign n10829 = pi618 & n7671;
  assign n10830 = ~pi618 & pi627;
  assign n10831 = pi1154 & n10830;
  assign n10832 = ~n10829 & ~n10831;
  assign n10833 = ~n10723 & ~n10832;
  assign n10834 = ~n7670 & ~n10737;
  assign n10835 = pi618 & ~n7597;
  assign n10836 = n7669 & ~n10835;
  assign n10837 = ~pi618 & ~n7597;
  assign n10838 = n7668 & ~n10837;
  assign n10839 = ~n10836 & ~n10838;
  assign n10840 = ~n10834 & n10839;
  assign n10841 = ~n10833 & n10840;
  assign n10842 = pi781 & ~n10711;
  assign n10843 = ~n10841 & n10842;
  assign n10844 = ~n10821 & ~n10822;
  assign n10845 = ~pi618 & ~n10844;
  assign n10846 = ~n10711 & ~n10723;
  assign n10847 = pi618 & ~n10846;
  assign n10848 = ~pi1154 & ~n10847;
  assign n10849 = ~n10845 & n10848;
  assign n10850 = n10737 & n10835;
  assign n10851 = pi1154 & ~n10711;
  assign n10852 = ~n10850 & n10851;
  assign n10853 = ~pi627 & ~n10852;
  assign n10854 = ~n10849 & n10853;
  assign n10855 = pi618 & ~n10844;
  assign n10856 = ~pi618 & ~n10846;
  assign n10857 = pi1154 & ~n10856;
  assign n10858 = ~n10855 & n10857;
  assign n10859 = n10737 & n10837;
  assign n10860 = ~pi1154 & ~n10711;
  assign n10861 = ~n10859 & n10860;
  assign n10862 = pi627 & ~n10861;
  assign n10863 = ~n10858 & n10862;
  assign n10864 = ~n10854 & ~n10863;
  assign n10865 = pi781 & ~n10864;
  assign n10866 = ~pi781 & ~n10844;
  assign n10867 = ~n10865 & ~n10866;
  assign n10868 = ~n10828 & ~n10843;
  assign n10869 = ~pi619 & ~n59353;
  assign n10870 = pi619 & ~n10765;
  assign n10871 = ~pi1159 & ~n10870;
  assign n10872 = ~n10869 & n10871;
  assign n10873 = n10737 & ~n59347;
  assign n10874 = pi619 & ~n7597;
  assign n10875 = n10873 & n10874;
  assign n10876 = pi1159 & ~n10711;
  assign n10877 = ~n10875 & n10876;
  assign n10878 = ~pi648 & ~n10877;
  assign n10879 = ~n10872 & n10878;
  assign n10880 = pi619 & ~n59353;
  assign n10881 = ~pi619 & ~n10765;
  assign n10882 = pi1159 & ~n10881;
  assign n10883 = ~n10880 & n10882;
  assign n10884 = ~pi619 & ~n7597;
  assign n10885 = n10873 & n10884;
  assign n10886 = ~pi1159 & ~n10711;
  assign n10887 = ~n10885 & n10886;
  assign n10888 = pi648 & ~n10887;
  assign n10889 = ~n10883 & n10888;
  assign n10890 = pi789 & ~n10889;
  assign n10891 = pi789 & ~n10879;
  assign n10892 = ~n10889 & n10891;
  assign n10893 = ~n10879 & n10890;
  assign n10894 = ~pi789 & n59353;
  assign n10895 = n59242 & ~n10894;
  assign n10896 = ~n59354 & n10895;
  assign n10897 = ~n10782 & ~n10896;
  assign n10898 = ~n10764 & ~n10897;
  assign n10899 = pi628 & pi629;
  assign n10900 = pi629 & n7961;
  assign n10901 = pi1156 & n10899;
  assign n10902 = ~pi628 & ~pi629;
  assign n10903 = ~pi629 & n7960;
  assign n10904 = ~pi1156 & n10902;
  assign n10905 = pi792 & ~n59356;
  assign n10906 = pi792 & ~n59355;
  assign n10907 = ~n59356 & n10906;
  assign n10908 = n7792 & n7959;
  assign n10909 = pi792 & ~n10908;
  assign n10910 = ~n59355 & n10905;
  assign n10911 = ~n10763 & n59357;
  assign n10912 = ~n8108 & ~n10911;
  assign n10913 = ~n10898 & n10912;
  assign n10914 = ~n59240 & n59345;
  assign n10915 = ~pi630 & ~n10914;
  assign n10916 = pi647 & ~n10915;
  assign n10917 = ~n7793 & n10753;
  assign n10918 = pi630 & n10917;
  assign n10919 = pi1157 & ~n10918;
  assign n10920 = ~n10916 & n10919;
  assign n10921 = pi630 & ~n10914;
  assign n10922 = ~pi647 & ~n10921;
  assign n10923 = ~pi630 & n10917;
  assign n10924 = ~pi1157 & ~n10923;
  assign n10925 = pi647 & ~n10923;
  assign n10926 = ~n10921 & ~n10925;
  assign n10927 = ~pi1157 & ~n10926;
  assign n10928 = ~n10922 & n10924;
  assign n10929 = ~n10920 & ~n59358;
  assign n10930 = pi787 & ~n10711;
  assign n10931 = ~n10929 & n10930;
  assign n10932 = ~n10913 & ~n10931;
  assign n10933 = pi644 & n10932;
  assign n10934 = ~n9743 & n10914;
  assign n10935 = ~n10711 & ~n10934;
  assign n10936 = ~pi644 & ~n10935;
  assign n10937 = pi715 & ~n10936;
  assign n10938 = ~n10933 & n10937;
  assign n10939 = ~n7835 & n10917;
  assign n10940 = pi644 & n10939;
  assign n10941 = ~pi715 & ~n10711;
  assign n10942 = ~n10940 & n10941;
  assign n10943 = pi1160 & ~n10942;
  assign n10944 = ~n10938 & n10943;
  assign n10945 = ~pi644 & n10932;
  assign n10946 = pi644 & ~n10935;
  assign n10947 = ~pi715 & ~n10946;
  assign n10948 = ~n10945 & n10947;
  assign n10949 = ~pi644 & n10939;
  assign n10950 = pi715 & ~n10711;
  assign n10951 = ~n10949 & n10950;
  assign n10952 = ~pi1160 & ~n10951;
  assign n10953 = ~n10948 & n10952;
  assign n10954 = ~n10944 & ~n10953;
  assign n10955 = pi790 & ~n10954;
  assign n10956 = ~pi790 & n10932;
  assign n10957 = pi832 & ~n10956;
  assign n10958 = ~n10955 & n10957;
  assign po301 = ~n10710 & ~n10958;
  assign n10960 = ~pi145 & ~n7560;
  assign n10961 = n59231 & ~n10960;
  assign n10962 = ~pi698 & n59132;
  assign n10963 = n10960 & ~n10962;
  assign n10964 = pi145 & n59251;
  assign n10965 = ~pi38 & ~n10964;
  assign n10966 = n59132 & ~n10965;
  assign n10967 = ~pi145 & n8249;
  assign n10968 = ~n10966 & ~n10967;
  assign n10969 = ~pi145 & ~n6863;
  assign n10970 = n7547 & ~n10969;
  assign n10971 = ~pi698 & ~n10970;
  assign n10972 = ~n10968 & n10971;
  assign n10973 = ~n10963 & ~n10972;
  assign n10974 = ~pi778 & n10973;
  assign n10975 = pi625 & ~n10973;
  assign n10976 = ~pi625 & n10960;
  assign n10977 = pi1153 & ~n10976;
  assign n10978 = ~n10975 & n10977;
  assign n10979 = ~pi625 & ~n10973;
  assign n10980 = pi625 & n10960;
  assign n10981 = ~pi1153 & ~n10980;
  assign n10982 = ~n10979 & n10981;
  assign n10983 = ~n10978 & ~n10982;
  assign n10984 = pi778 & ~n10983;
  assign n10985 = ~n10974 & ~n10984;
  assign n10986 = ~n59229 & n10985;
  assign n10987 = n59229 & n10960;
  assign n10988 = n59229 & ~n10960;
  assign n10989 = ~n59229 & ~n10985;
  assign n10990 = ~n10988 & ~n10989;
  assign n10991 = ~n10986 & ~n10987;
  assign n10992 = ~n59231 & ~n59359;
  assign n10993 = ~n59231 & n59359;
  assign n10994 = n59231 & n10960;
  assign n10995 = ~n10993 & ~n10994;
  assign n10996 = ~n10961 & ~n10992;
  assign n10997 = ~n7716 & ~n59360;
  assign n10998 = n7716 & n10960;
  assign n10999 = n7716 & ~n10960;
  assign n11000 = ~n7716 & n59360;
  assign n11001 = ~n10999 & ~n11000;
  assign n11002 = ~n10997 & ~n10998;
  assign n11003 = ~n7762 & n59361;
  assign n11004 = n7762 & n10960;
  assign n11005 = ~n11003 & ~n11004;
  assign n11006 = ~pi792 & n11005;
  assign n11007 = pi628 & ~n11005;
  assign n11008 = ~pi628 & n10960;
  assign n11009 = pi1156 & ~n11008;
  assign n11010 = ~n11007 & n11009;
  assign n11011 = ~pi628 & ~n11005;
  assign n11012 = pi628 & n10960;
  assign n11013 = ~pi1156 & ~n11012;
  assign n11014 = ~n11011 & n11013;
  assign n11015 = ~n11010 & ~n11014;
  assign n11016 = pi792 & ~n11015;
  assign n11017 = ~n11006 & ~n11016;
  assign n11018 = pi647 & n11017;
  assign n11019 = ~pi647 & n10960;
  assign n11020 = pi1157 & ~n11019;
  assign n11021 = pi647 & ~n11017;
  assign n11022 = ~pi647 & ~n10960;
  assign n11023 = ~n11021 & ~n11022;
  assign n11024 = pi1157 & ~n11023;
  assign n11025 = ~n11018 & n11020;
  assign n11026 = ~pi647 & n11017;
  assign n11027 = pi647 & n10960;
  assign n11028 = ~pi1157 & ~n11027;
  assign n11029 = ~n11026 & n11028;
  assign n11030 = ~pi647 & ~n11017;
  assign n11031 = pi647 & ~n10960;
  assign n11032 = ~n11030 & ~n11031;
  assign n11033 = ~pi1157 & n11032;
  assign n11034 = pi1157 & n11023;
  assign n11035 = ~n11033 & ~n11034;
  assign n11036 = ~n59362 & ~n11029;
  assign n11037 = pi787 & n59363;
  assign n11038 = ~pi787 & ~n11017;
  assign n11039 = pi787 & ~n59363;
  assign n11040 = ~pi787 & n11017;
  assign n11041 = ~n11039 & ~n11040;
  assign n11042 = ~n11037 & ~n11038;
  assign n11043 = ~pi644 & ~n59364;
  assign n11044 = pi715 & ~n11043;
  assign n11045 = pi145 & ~n59132;
  assign n11046 = ~pi767 & n6865;
  assign n11047 = ~n10969 & ~n11046;
  assign n11048 = pi38 & ~n11047;
  assign n11049 = ~pi145 & n59164;
  assign n11050 = pi145 & ~n6855;
  assign n11051 = ~pi767 & ~n11050;
  assign n11052 = ~n11049 & n11051;
  assign n11053 = ~pi145 & pi767;
  assign n11054 = ~n6656 & n11053;
  assign n11055 = ~pi145 & ~n6656;
  assign n11056 = pi767 & ~n11055;
  assign n11057 = ~pi145 & ~pi767;
  assign n11058 = n59164 & n11057;
  assign n11059 = ~n11050 & ~n11058;
  assign n11060 = ~n11056 & n11059;
  assign n11061 = ~n11052 & ~n11054;
  assign n11062 = ~pi38 & n59365;
  assign n11063 = ~pi38 & ~n59365;
  assign n11064 = pi38 & ~n10969;
  assign n11065 = ~n11046 & n11064;
  assign n11066 = ~n11063 & ~n11065;
  assign n11067 = ~n11048 & ~n11062;
  assign n11068 = n59132 & ~n59366;
  assign n11069 = ~n11045 & ~n11068;
  assign n11070 = ~n7597 & ~n11069;
  assign n11071 = n7597 & ~n10960;
  assign n11072 = ~n11070 & ~n11071;
  assign n11073 = ~pi785 & ~n11072;
  assign n11074 = ~n7598 & ~n10960;
  assign n11075 = pi609 & n11070;
  assign n11076 = ~n11074 & ~n11075;
  assign n11077 = pi1155 & ~n11076;
  assign n11078 = ~n7610 & ~n10960;
  assign n11079 = ~pi609 & n11070;
  assign n11080 = ~n11078 & ~n11079;
  assign n11081 = ~pi1155 & ~n11080;
  assign n11082 = ~n11077 & ~n11081;
  assign n11083 = pi785 & ~n11082;
  assign n11084 = ~n11073 & ~n11083;
  assign n11085 = ~pi781 & ~n11084;
  assign n11086 = pi618 & n11084;
  assign n11087 = ~pi618 & n10960;
  assign n11088 = pi1154 & ~n11087;
  assign n11089 = ~n11086 & n11088;
  assign n11090 = ~pi618 & n11084;
  assign n11091 = pi618 & n10960;
  assign n11092 = ~pi1154 & ~n11091;
  assign n11093 = ~n11090 & n11092;
  assign n11094 = ~n11089 & ~n11093;
  assign n11095 = pi781 & ~n11094;
  assign n11096 = ~n11085 & ~n11095;
  assign n11097 = ~pi789 & ~n11096;
  assign n11098 = pi619 & n11096;
  assign n11099 = ~pi619 & n10960;
  assign n11100 = pi1159 & ~n11099;
  assign n11101 = ~n11098 & n11100;
  assign n11102 = ~pi619 & n11096;
  assign n11103 = pi619 & n10960;
  assign n11104 = ~pi1159 & ~n11103;
  assign n11105 = ~n11102 & n11104;
  assign n11106 = ~n11101 & ~n11105;
  assign n11107 = pi789 & ~n11106;
  assign n11108 = ~n11097 & ~n11107;
  assign n11109 = n7913 & n11108;
  assign n11110 = ~n7913 & n10960;
  assign n11111 = pi626 & n11108;
  assign n11112 = ~pi626 & n10960;
  assign n11113 = pi1158 & ~n11112;
  assign n11114 = ~n11111 & n11113;
  assign n11115 = ~pi626 & n11108;
  assign n11116 = pi626 & n10960;
  assign n11117 = ~pi1158 & ~n11116;
  assign n11118 = ~n11115 & n11117;
  assign n11119 = ~n11114 & ~n11118;
  assign n11120 = ~n11109 & ~n11110;
  assign n11121 = pi788 & n59367;
  assign n11122 = ~pi788 & n11108;
  assign n11123 = ~pi788 & ~n11108;
  assign n11124 = pi788 & ~n59367;
  assign n11125 = ~n11123 & ~n11124;
  assign n11126 = ~n11121 & ~n11122;
  assign n11127 = ~n7793 & n59368;
  assign n11128 = n7793 & n10960;
  assign n11129 = ~n11127 & ~n11128;
  assign n11130 = ~n7835 & ~n11129;
  assign n11131 = n7835 & n10960;
  assign n11132 = n7835 & ~n10960;
  assign n11133 = ~n7835 & n11129;
  assign n11134 = ~n11132 & ~n11133;
  assign n11135 = ~n11130 & ~n11131;
  assign n11136 = pi644 & n59369;
  assign n11137 = ~pi644 & n10960;
  assign n11138 = ~pi715 & ~n11137;
  assign n11139 = ~n11136 & n11138;
  assign n11140 = pi1160 & ~n11139;
  assign n11141 = ~n11044 & n11140;
  assign n11142 = ~n7872 & n11129;
  assign n11143 = n7832 & ~n11023;
  assign n11144 = ~pi630 & n59362;
  assign n11145 = n7833 & ~n11032;
  assign n11146 = pi630 & n11029;
  assign n11147 = ~n59370 & ~n59371;
  assign n11148 = ~n11142 & n11147;
  assign n11149 = pi787 & ~n11148;
  assign n11150 = ~pi628 & pi629;
  assign n11151 = pi1156 & n11150;
  assign n11152 = pi628 & ~pi629;
  assign n11153 = ~pi1156 & n11152;
  assign n11154 = ~n11151 & ~n11153;
  assign n11155 = ~n59368 & ~n11154;
  assign n11156 = ~pi629 & n11010;
  assign n11157 = pi629 & n11014;
  assign n11158 = ~n11156 & ~n11157;
  assign n11159 = ~n11155 & n11158;
  assign n11160 = pi792 & ~n11159;
  assign n11161 = pi698 & n59366;
  assign n11162 = ~pi145 & n59177;
  assign n11163 = pi145 & n7111;
  assign n11164 = pi767 & ~n11163;
  assign n11165 = ~n11162 & n11164;
  assign n11166 = pi145 & n7188;
  assign n11167 = ~pi145 & ~n59203;
  assign n11168 = ~pi767 & ~n11167;
  assign n11169 = ~n11166 & n11168;
  assign n11170 = pi39 & ~n11169;
  assign n11171 = ~n11165 & n11170;
  assign n11172 = pi145 & n7333;
  assign n11173 = ~pi145 & n7310;
  assign n11174 = pi767 & ~n11173;
  assign n11175 = ~n11172 & n11174;
  assign n11176 = ~pi145 & ~n7339;
  assign n11177 = pi145 & ~n7347;
  assign n11178 = ~pi767 & ~n11177;
  assign n11179 = ~n11176 & n11178;
  assign n11180 = ~pi39 & ~n11179;
  assign n11181 = pi145 & ~n7333;
  assign n11182 = ~pi145 & ~n7310;
  assign n11183 = pi767 & ~n11182;
  assign n11184 = pi767 & ~n11181;
  assign n11185 = ~n11182 & n11184;
  assign n11186 = ~n11181 & n11183;
  assign n11187 = ~pi145 & n7339;
  assign n11188 = pi145 & n7347;
  assign n11189 = ~pi767 & ~n11188;
  assign n11190 = ~n11187 & n11189;
  assign n11191 = ~n59372 & ~n11190;
  assign n11192 = ~pi39 & ~n11191;
  assign n11193 = ~n11175 & n11180;
  assign n11194 = ~pi38 & ~n59373;
  assign n11195 = ~n11171 & n11194;
  assign n11196 = ~pi767 & ~n7222;
  assign n11197 = n9794 & ~n11196;
  assign n11198 = ~pi145 & ~n11197;
  assign n11199 = ~pi767 & n6822;
  assign n11200 = ~n7056 & ~n11199;
  assign n11201 = pi145 & ~n11200;
  assign n11202 = n59171 & n11201;
  assign n11203 = pi38 & ~n11202;
  assign n11204 = ~n11198 & n11203;
  assign n11205 = ~pi698 & ~n11204;
  assign n11206 = ~n11195 & n11205;
  assign n11207 = n59132 & ~n11206;
  assign n11208 = ~n11161 & n11207;
  assign n11209 = ~n11045 & ~n11208;
  assign n11210 = ~pi625 & n11209;
  assign n11211 = pi625 & n11069;
  assign n11212 = ~pi1153 & ~n11211;
  assign n11213 = ~n11210 & n11212;
  assign n11214 = ~pi608 & ~n10978;
  assign n11215 = ~n11213 & n11214;
  assign n11216 = pi625 & n11209;
  assign n11217 = ~pi625 & n11069;
  assign n11218 = pi1153 & ~n11217;
  assign n11219 = ~n11216 & n11218;
  assign n11220 = pi608 & ~n10982;
  assign n11221 = ~n11219 & n11220;
  assign n11222 = ~n11215 & ~n11221;
  assign n11223 = pi778 & ~n11222;
  assign n11224 = ~pi778 & n11209;
  assign n11225 = ~n11223 & ~n11224;
  assign n11226 = ~pi609 & ~n11225;
  assign n11227 = pi609 & n10985;
  assign n11228 = ~pi1155 & ~n11227;
  assign n11229 = ~n11226 & n11228;
  assign n11230 = ~pi660 & ~n11077;
  assign n11231 = ~n11229 & n11230;
  assign n11232 = pi609 & ~n11225;
  assign n11233 = ~pi609 & n10985;
  assign n11234 = pi1155 & ~n11233;
  assign n11235 = ~n11232 & n11234;
  assign n11236 = pi660 & ~n11081;
  assign n11237 = ~n11235 & n11236;
  assign n11238 = ~n11231 & ~n11237;
  assign n11239 = pi785 & ~n11238;
  assign n11240 = ~pi785 & ~n11225;
  assign n11241 = ~n11239 & ~n11240;
  assign n11242 = ~pi618 & ~n11241;
  assign n11243 = pi618 & n59359;
  assign n11244 = ~pi1154 & ~n11243;
  assign n11245 = ~n11242 & n11244;
  assign n11246 = ~pi627 & ~n11089;
  assign n11247 = ~n11245 & n11246;
  assign n11248 = pi618 & ~n11241;
  assign n11249 = ~pi618 & n59359;
  assign n11250 = pi1154 & ~n11249;
  assign n11251 = ~n11248 & n11250;
  assign n11252 = pi627 & ~n11093;
  assign n11253 = ~n11251 & n11252;
  assign n11254 = ~n11247 & ~n11253;
  assign n11255 = pi781 & ~n11254;
  assign n11256 = ~pi781 & ~n11241;
  assign n11257 = ~n11255 & ~n11256;
  assign n11258 = ~pi619 & ~n11257;
  assign n11259 = pi619 & ~n59360;
  assign n11260 = ~pi1159 & ~n11259;
  assign n11261 = ~n11258 & n11260;
  assign n11262 = ~pi648 & ~n11101;
  assign n11263 = ~n11261 & n11262;
  assign n11264 = pi619 & ~n11257;
  assign n11265 = ~pi619 & ~n59360;
  assign n11266 = pi1159 & ~n11265;
  assign n11267 = ~n11264 & n11266;
  assign n11268 = pi648 & ~n11105;
  assign n11269 = ~n11267 & n11268;
  assign n11270 = pi789 & ~n11269;
  assign n11271 = pi789 & ~n11263;
  assign n11272 = ~n11269 & n11271;
  assign n11273 = ~n11263 & n11270;
  assign n11274 = ~pi789 & n11257;
  assign n11275 = n59242 & ~n11274;
  assign n11276 = ~n59374 & n11275;
  assign n11277 = n7984 & n59361;
  assign n11278 = ~n7761 & n59367;
  assign n11279 = ~n11277 & ~n11278;
  assign n11280 = pi788 & ~n11279;
  assign n11281 = ~n59357 & ~n11280;
  assign n11282 = ~n11276 & n11281;
  assign n11283 = ~n11160 & ~n11282;
  assign n11284 = ~n8108 & ~n11283;
  assign n11285 = ~n11149 & ~n11284;
  assign n11286 = ~pi644 & n11285;
  assign n11287 = pi644 & ~n59364;
  assign n11288 = ~pi715 & ~n11287;
  assign n11289 = ~n11286 & n11288;
  assign n11290 = ~pi644 & n59369;
  assign n11291 = pi644 & n10960;
  assign n11292 = pi715 & ~n11291;
  assign n11293 = ~n11290 & n11292;
  assign n11294 = ~pi1160 & ~n11293;
  assign n11295 = ~n11289 & n11294;
  assign n11296 = ~n11141 & ~n11295;
  assign n11297 = pi790 & ~n11296;
  assign n11298 = pi644 & n11140;
  assign n11299 = pi790 & ~n11298;
  assign n11300 = n11285 & ~n11299;
  assign n11301 = ~n11297 & ~n11300;
  assign n11302 = n58992 & ~n11301;
  assign n11303 = ~pi145 & ~n58992;
  assign n11304 = ~pi832 & ~n11303;
  assign n11305 = ~n11302 & n11304;
  assign n11306 = ~pi145 & ~n2794;
  assign n11307 = ~n11199 & ~n11306;
  assign n11308 = ~n7875 & ~n11307;
  assign n11309 = ~pi785 & ~n11308;
  assign n11310 = ~n7880 & ~n11307;
  assign n11311 = pi1155 & ~n11310;
  assign n11312 = ~n7883 & n11308;
  assign n11313 = ~pi1155 & ~n11312;
  assign n11314 = ~n11311 & ~n11313;
  assign n11315 = pi785 & ~n11314;
  assign n11316 = ~n11309 & ~n11315;
  assign n11317 = ~pi781 & ~n11316;
  assign n11318 = ~n7890 & n11316;
  assign n11319 = pi1154 & ~n11318;
  assign n11320 = ~n7893 & n11316;
  assign n11321 = ~pi1154 & ~n11320;
  assign n11322 = ~n11319 & ~n11321;
  assign n11323 = pi781 & ~n11322;
  assign n11324 = ~n11317 & ~n11323;
  assign n11325 = ~pi789 & ~n11324;
  assign n11326 = pi619 & n11324;
  assign n11327 = ~pi619 & n11306;
  assign n11328 = pi1159 & ~n11327;
  assign n11329 = ~n11326 & n11328;
  assign n11330 = ~pi619 & n11324;
  assign n11331 = pi619 & n11306;
  assign n11332 = ~pi1159 & ~n11331;
  assign n11333 = ~n11330 & n11332;
  assign n11334 = ~n11329 & ~n11333;
  assign n11335 = pi789 & ~n11334;
  assign n11336 = ~n11325 & ~n11335;
  assign n11337 = n7913 & n11336;
  assign n11338 = ~n7913 & n11306;
  assign n11339 = pi626 & n11336;
  assign n11340 = ~pi626 & n11306;
  assign n11341 = pi1158 & ~n11340;
  assign n11342 = ~n11339 & n11341;
  assign n11343 = ~pi626 & n11336;
  assign n11344 = pi626 & n11306;
  assign n11345 = ~pi1158 & ~n11344;
  assign n11346 = ~n11343 & n11345;
  assign n11347 = ~n11342 & ~n11346;
  assign n11348 = ~n11337 & ~n11338;
  assign n11349 = pi788 & n59375;
  assign n11350 = ~pi788 & n11336;
  assign n11351 = ~pi788 & ~n11336;
  assign n11352 = pi788 & ~n59375;
  assign n11353 = ~n11351 & ~n11352;
  assign n11354 = ~n11349 & ~n11350;
  assign n11355 = ~n7793 & n59376;
  assign n11356 = n7793 & n11306;
  assign n11357 = ~n7872 & ~n11356;
  assign n11358 = ~n11355 & ~n11356;
  assign n11359 = ~n7872 & n11358;
  assign n11360 = ~n11355 & n11357;
  assign n11361 = ~pi698 & n7055;
  assign n11362 = ~n11306 & ~n11361;
  assign n11363 = ~pi778 & n11362;
  assign n11364 = ~pi625 & n11361;
  assign n11365 = ~n11362 & ~n11364;
  assign n11366 = pi1153 & ~n11365;
  assign n11367 = ~pi1153 & ~n11306;
  assign n11368 = ~n11364 & n11367;
  assign n11369 = ~n11366 & ~n11368;
  assign n11370 = pi778 & ~n11369;
  assign n11371 = ~n11363 & ~n11370;
  assign n11372 = ~n7949 & n11371;
  assign n11373 = ~n7951 & n11372;
  assign n11374 = ~n7953 & n11373;
  assign n11375 = ~n7955 & n11374;
  assign n11376 = ~n7967 & n11375;
  assign n11377 = pi647 & ~n11376;
  assign n11378 = ~pi647 & ~n11306;
  assign n11379 = ~n11377 & ~n11378;
  assign n11380 = n7832 & ~n11379;
  assign n11381 = ~pi647 & n11376;
  assign n11382 = pi647 & n11306;
  assign n11383 = ~pi1157 & ~n11382;
  assign n11384 = ~n11381 & n11383;
  assign n11385 = pi630 & n11384;
  assign n11386 = ~n11380 & ~n11385;
  assign n11387 = ~n59377 & n11386;
  assign n11388 = pi787 & ~n11387;
  assign n11389 = n7984 & n11374;
  assign n11390 = ~n7761 & n59375;
  assign n11391 = ~n11389 & ~n11390;
  assign n11392 = pi788 & ~n11391;
  assign n11393 = ~n6701 & ~n11362;
  assign n11394 = pi625 & n11393;
  assign n11395 = n11307 & ~n11393;
  assign n11396 = ~n11394 & ~n11395;
  assign n11397 = n11367 & ~n11396;
  assign n11398 = ~pi608 & ~n11366;
  assign n11399 = ~n11397 & n11398;
  assign n11400 = pi1153 & n11307;
  assign n11401 = ~n11394 & n11400;
  assign n11402 = pi608 & ~n11368;
  assign n11403 = ~n11401 & n11402;
  assign n11404 = ~n11399 & ~n11403;
  assign n11405 = pi778 & ~n11404;
  assign n11406 = ~pi778 & ~n11395;
  assign n11407 = ~n11405 & ~n11406;
  assign n11408 = ~pi609 & ~n11407;
  assign n11409 = pi609 & n11371;
  assign n11410 = ~pi1155 & ~n11409;
  assign n11411 = ~n11408 & n11410;
  assign n11412 = ~pi660 & ~n11311;
  assign n11413 = ~n11411 & n11412;
  assign n11414 = pi609 & ~n11407;
  assign n11415 = ~pi609 & n11371;
  assign n11416 = pi1155 & ~n11415;
  assign n11417 = ~n11414 & n11416;
  assign n11418 = pi660 & ~n11313;
  assign n11419 = ~n11417 & n11418;
  assign n11420 = ~n11413 & ~n11419;
  assign n11421 = pi785 & ~n11420;
  assign n11422 = ~pi785 & ~n11407;
  assign n11423 = ~n11421 & ~n11422;
  assign n11424 = ~pi618 & ~n11423;
  assign n11425 = pi618 & n11372;
  assign n11426 = ~pi1154 & ~n11425;
  assign n11427 = ~n11424 & n11426;
  assign n11428 = ~pi627 & ~n11319;
  assign n11429 = ~n11427 & n11428;
  assign n11430 = pi618 & ~n11423;
  assign n11431 = ~pi618 & n11372;
  assign n11432 = pi1154 & ~n11431;
  assign n11433 = ~n11430 & n11432;
  assign n11434 = pi627 & ~n11321;
  assign n11435 = ~n11433 & n11434;
  assign n11436 = ~n11429 & ~n11435;
  assign n11437 = pi781 & ~n11436;
  assign n11438 = ~pi781 & ~n11423;
  assign n11439 = ~n11437 & ~n11438;
  assign n11440 = ~pi619 & ~n11439;
  assign n11441 = pi619 & n11373;
  assign n11442 = ~pi1159 & ~n11441;
  assign n11443 = ~n11440 & n11442;
  assign n11444 = ~pi648 & ~n11329;
  assign n11445 = ~n11443 & n11444;
  assign n11446 = pi619 & ~n11439;
  assign n11447 = ~pi619 & n11373;
  assign n11448 = pi1159 & ~n11447;
  assign n11449 = ~n11446 & n11448;
  assign n11450 = pi648 & ~n11333;
  assign n11451 = ~n11449 & n11450;
  assign n11452 = pi789 & ~n11451;
  assign n11453 = pi789 & ~n11445;
  assign n11454 = ~n11451 & n11453;
  assign n11455 = ~n11445 & n11452;
  assign n11456 = ~pi789 & n11439;
  assign n11457 = n59242 & ~n11456;
  assign n11458 = ~n59378 & n11457;
  assign n11459 = ~n11392 & ~n11458;
  assign n11460 = ~n59357 & ~n11459;
  assign n11461 = n7957 & n59376;
  assign n11462 = n8065 & n11375;
  assign n11463 = pi629 & ~n11462;
  assign n11464 = ~n11461 & n11463;
  assign n11465 = n7958 & n59376;
  assign n11466 = n8074 & n11375;
  assign n11467 = ~pi629 & ~n11466;
  assign n11468 = ~n11465 & n11467;
  assign n11469 = pi792 & ~n11468;
  assign n11470 = ~n11465 & ~n11466;
  assign n11471 = ~pi629 & ~n11470;
  assign n11472 = ~n11461 & ~n11462;
  assign n11473 = pi629 & ~n11472;
  assign n11474 = ~n11471 & ~n11473;
  assign n11475 = pi792 & ~n11474;
  assign n11476 = pi792 & ~n11464;
  assign n11477 = ~n11468 & n11476;
  assign n11478 = ~n11464 & n11469;
  assign n11479 = ~n8108 & ~n59379;
  assign n11480 = ~n11460 & n11479;
  assign n11481 = ~n11388 & ~n11480;
  assign n11482 = pi644 & n11481;
  assign n11483 = ~pi787 & ~n11376;
  assign n11484 = pi1157 & ~n11379;
  assign n11485 = ~n11384 & ~n11484;
  assign n11486 = pi787 & ~n11485;
  assign n11487 = ~n11483 & ~n11486;
  assign n11488 = ~pi644 & n11487;
  assign n11489 = pi715 & ~n11488;
  assign n11490 = ~n11482 & n11489;
  assign n11491 = ~n7793 & ~n7835;
  assign n11492 = n11306 & ~n11491;
  assign n11493 = ~n7835 & n11355;
  assign n11494 = ~n7835 & ~n11358;
  assign n11495 = n7835 & n11306;
  assign n11496 = ~n11494 & ~n11495;
  assign n11497 = ~n11492 & ~n11493;
  assign n11498 = pi644 & ~n59380;
  assign n11499 = ~pi644 & n11306;
  assign n11500 = ~pi715 & ~n11499;
  assign n11501 = ~n11498 & n11500;
  assign n11502 = pi1160 & ~n11501;
  assign n11503 = ~n11490 & n11502;
  assign n11504 = ~pi644 & n11481;
  assign n11505 = pi644 & n11487;
  assign n11506 = ~pi715 & ~n11505;
  assign n11507 = ~n11504 & n11506;
  assign n11508 = ~pi644 & ~n59380;
  assign n11509 = pi644 & n11306;
  assign n11510 = pi715 & ~n11509;
  assign n11511 = ~n11508 & n11510;
  assign n11512 = ~pi1160 & ~n11511;
  assign n11513 = ~n11507 & n11512;
  assign n11514 = ~n11503 & ~n11513;
  assign n11515 = pi790 & ~n11514;
  assign n11516 = ~pi790 & n11481;
  assign n11517 = pi832 & ~n11516;
  assign n11518 = ~n11515 & n11517;
  assign po302 = ~n11305 & ~n11518;
  assign n11520 = ~pi173 & ~n7560;
  assign n11521 = n59231 & ~n11520;
  assign n11522 = ~pi723 & n59132;
  assign n11523 = n11520 & ~n11522;
  assign n11524 = pi173 & n59251;
  assign n11525 = ~pi38 & ~n11524;
  assign n11526 = n59132 & ~n11525;
  assign n11527 = ~pi173 & n8249;
  assign n11528 = ~n11526 & ~n11527;
  assign n11529 = ~pi173 & ~n6863;
  assign n11530 = n7547 & ~n11529;
  assign n11531 = ~pi723 & ~n11530;
  assign n11532 = ~n11528 & n11531;
  assign n11533 = ~n11523 & ~n11532;
  assign n11534 = ~pi778 & n11533;
  assign n11535 = pi625 & ~n11533;
  assign n11536 = ~pi625 & n11520;
  assign n11537 = pi1153 & ~n11536;
  assign n11538 = ~n11535 & n11537;
  assign n11539 = ~pi625 & ~n11533;
  assign n11540 = pi625 & n11520;
  assign n11541 = ~pi1153 & ~n11540;
  assign n11542 = ~n11539 & n11541;
  assign n11543 = ~n11538 & ~n11542;
  assign n11544 = pi778 & ~n11543;
  assign n11545 = ~n11534 & ~n11544;
  assign n11546 = ~n59229 & n11545;
  assign n11547 = n59229 & n11520;
  assign n11548 = n59229 & ~n11520;
  assign n11549 = ~n59229 & ~n11545;
  assign n11550 = ~n11548 & ~n11549;
  assign n11551 = ~n11546 & ~n11547;
  assign n11552 = ~n59231 & ~n59381;
  assign n11553 = ~n59231 & n59381;
  assign n11554 = n59231 & n11520;
  assign n11555 = ~n11553 & ~n11554;
  assign n11556 = ~n11521 & ~n11552;
  assign n11557 = ~n7716 & ~n59382;
  assign n11558 = n7716 & n11520;
  assign n11559 = n7716 & ~n11520;
  assign n11560 = ~n7716 & n59382;
  assign n11561 = ~n11559 & ~n11560;
  assign n11562 = ~n11557 & ~n11558;
  assign n11563 = ~n7762 & n59383;
  assign n11564 = n7762 & n11520;
  assign n11565 = ~n11563 & ~n11564;
  assign n11566 = ~pi792 & n11565;
  assign n11567 = pi628 & ~n11565;
  assign n11568 = ~pi628 & n11520;
  assign n11569 = pi1156 & ~n11568;
  assign n11570 = ~n11567 & n11569;
  assign n11571 = ~pi628 & ~n11565;
  assign n11572 = pi628 & n11520;
  assign n11573 = ~pi1156 & ~n11572;
  assign n11574 = ~n11571 & n11573;
  assign n11575 = ~n11570 & ~n11574;
  assign n11576 = pi792 & ~n11575;
  assign n11577 = ~n11566 & ~n11576;
  assign n11578 = pi647 & n11577;
  assign n11579 = ~pi647 & n11520;
  assign n11580 = pi1157 & ~n11579;
  assign n11581 = pi647 & ~n11577;
  assign n11582 = ~pi647 & ~n11520;
  assign n11583 = ~n11581 & ~n11582;
  assign n11584 = pi1157 & ~n11583;
  assign n11585 = ~n11578 & n11580;
  assign n11586 = ~pi647 & n11577;
  assign n11587 = pi647 & n11520;
  assign n11588 = ~pi1157 & ~n11587;
  assign n11589 = ~n11586 & n11588;
  assign n11590 = ~pi647 & ~n11577;
  assign n11591 = pi647 & ~n11520;
  assign n11592 = ~n11590 & ~n11591;
  assign n11593 = ~pi1157 & n11592;
  assign n11594 = pi1157 & n11583;
  assign n11595 = ~n11593 & ~n11594;
  assign n11596 = ~n59384 & ~n11589;
  assign n11597 = pi787 & n59385;
  assign n11598 = ~pi787 & ~n11577;
  assign n11599 = pi787 & ~n59385;
  assign n11600 = ~pi787 & n11577;
  assign n11601 = ~n11599 & ~n11600;
  assign n11602 = ~n11597 & ~n11598;
  assign n11603 = ~pi644 & ~n59386;
  assign n11604 = pi715 & ~n11603;
  assign n11605 = pi173 & ~n59132;
  assign n11606 = ~pi745 & n6865;
  assign n11607 = ~n11529 & ~n11606;
  assign n11608 = pi38 & ~n11607;
  assign n11609 = ~pi173 & n59164;
  assign n11610 = pi173 & ~n6855;
  assign n11611 = ~pi745 & ~n11610;
  assign n11612 = ~n11609 & n11611;
  assign n11613 = ~pi173 & pi745;
  assign n11614 = ~n6656 & n11613;
  assign n11615 = ~pi173 & ~n6656;
  assign n11616 = pi745 & ~n11615;
  assign n11617 = ~pi173 & ~pi745;
  assign n11618 = n59164 & n11617;
  assign n11619 = ~n11610 & ~n11618;
  assign n11620 = ~n11616 & n11619;
  assign n11621 = ~n11612 & ~n11614;
  assign n11622 = ~pi38 & n59387;
  assign n11623 = ~pi38 & ~n59387;
  assign n11624 = pi38 & ~n11529;
  assign n11625 = ~n11606 & n11624;
  assign n11626 = ~n11623 & ~n11625;
  assign n11627 = ~n11608 & ~n11622;
  assign n11628 = n59132 & ~n59388;
  assign n11629 = ~n11605 & ~n11628;
  assign n11630 = ~n7597 & ~n11629;
  assign n11631 = n7597 & ~n11520;
  assign n11632 = ~n11630 & ~n11631;
  assign n11633 = ~pi785 & ~n11632;
  assign n11634 = ~n7598 & ~n11520;
  assign n11635 = pi609 & n11630;
  assign n11636 = ~n11634 & ~n11635;
  assign n11637 = pi1155 & ~n11636;
  assign n11638 = ~n7610 & ~n11520;
  assign n11639 = ~pi609 & n11630;
  assign n11640 = ~n11638 & ~n11639;
  assign n11641 = ~pi1155 & ~n11640;
  assign n11642 = ~n11637 & ~n11641;
  assign n11643 = pi785 & ~n11642;
  assign n11644 = ~n11633 & ~n11643;
  assign n11645 = ~pi781 & ~n11644;
  assign n11646 = pi618 & n11644;
  assign n11647 = ~pi618 & n11520;
  assign n11648 = pi1154 & ~n11647;
  assign n11649 = ~n11646 & n11648;
  assign n11650 = ~pi618 & n11644;
  assign n11651 = pi618 & n11520;
  assign n11652 = ~pi1154 & ~n11651;
  assign n11653 = ~n11650 & n11652;
  assign n11654 = ~n11649 & ~n11653;
  assign n11655 = pi781 & ~n11654;
  assign n11656 = ~n11645 & ~n11655;
  assign n11657 = ~pi789 & ~n11656;
  assign n11658 = pi619 & n11656;
  assign n11659 = ~pi619 & n11520;
  assign n11660 = pi1159 & ~n11659;
  assign n11661 = ~n11658 & n11660;
  assign n11662 = ~pi619 & n11656;
  assign n11663 = pi619 & n11520;
  assign n11664 = ~pi1159 & ~n11663;
  assign n11665 = ~n11662 & n11664;
  assign n11666 = ~n11661 & ~n11665;
  assign n11667 = pi789 & ~n11666;
  assign n11668 = ~n11657 & ~n11667;
  assign n11669 = n7913 & n11668;
  assign n11670 = ~n7913 & n11520;
  assign n11671 = pi626 & n11668;
  assign n11672 = ~pi626 & n11520;
  assign n11673 = pi1158 & ~n11672;
  assign n11674 = ~n11671 & n11673;
  assign n11675 = ~pi626 & n11668;
  assign n11676 = pi626 & n11520;
  assign n11677 = ~pi1158 & ~n11676;
  assign n11678 = ~n11675 & n11677;
  assign n11679 = ~n11674 & ~n11678;
  assign n11680 = ~n11669 & ~n11670;
  assign n11681 = pi788 & n59389;
  assign n11682 = ~pi788 & n11668;
  assign n11683 = ~pi788 & ~n11668;
  assign n11684 = pi788 & ~n59389;
  assign n11685 = ~n11683 & ~n11684;
  assign n11686 = ~n11681 & ~n11682;
  assign n11687 = ~n7793 & n59390;
  assign n11688 = n7793 & n11520;
  assign n11689 = ~n11687 & ~n11688;
  assign n11690 = ~n7835 & ~n11689;
  assign n11691 = n7835 & n11520;
  assign n11692 = n7835 & ~n11520;
  assign n11693 = ~n7835 & n11689;
  assign n11694 = ~n11692 & ~n11693;
  assign n11695 = ~n11690 & ~n11691;
  assign n11696 = pi644 & n59391;
  assign n11697 = ~pi644 & n11520;
  assign n11698 = ~pi715 & ~n11697;
  assign n11699 = ~n11696 & n11698;
  assign n11700 = pi1160 & ~n11699;
  assign n11701 = ~n11604 & n11700;
  assign n11702 = ~n7872 & n11689;
  assign n11703 = n7832 & ~n11583;
  assign n11704 = ~pi630 & n59384;
  assign n11705 = n7833 & ~n11592;
  assign n11706 = pi630 & n11589;
  assign n11707 = ~n59392 & ~n59393;
  assign n11708 = ~n11702 & n11707;
  assign n11709 = pi787 & ~n11708;
  assign n11710 = ~n11154 & ~n59390;
  assign n11711 = ~pi629 & n11570;
  assign n11712 = pi629 & n11574;
  assign n11713 = ~n11711 & ~n11712;
  assign n11714 = ~n11710 & n11713;
  assign n11715 = pi792 & ~n11714;
  assign n11716 = pi723 & n59388;
  assign n11717 = ~pi173 & n59177;
  assign n11718 = pi173 & n7111;
  assign n11719 = pi745 & ~n11718;
  assign n11720 = ~n11717 & n11719;
  assign n11721 = pi173 & n7188;
  assign n11722 = ~pi173 & ~n59203;
  assign n11723 = ~pi745 & ~n11722;
  assign n11724 = ~n11721 & n11723;
  assign n11725 = pi39 & ~n11724;
  assign n11726 = ~n11720 & n11725;
  assign n11727 = pi173 & n7333;
  assign n11728 = ~pi173 & n7310;
  assign n11729 = pi745 & ~n11728;
  assign n11730 = ~n11727 & n11729;
  assign n11731 = ~pi173 & ~n7339;
  assign n11732 = pi173 & ~n7347;
  assign n11733 = ~pi745 & ~n11732;
  assign n11734 = ~n11731 & n11733;
  assign n11735 = ~pi39 & ~n11734;
  assign n11736 = pi173 & ~n7333;
  assign n11737 = ~pi173 & ~n7310;
  assign n11738 = pi745 & ~n11737;
  assign n11739 = pi745 & ~n11736;
  assign n11740 = ~n11737 & n11739;
  assign n11741 = ~n11736 & n11738;
  assign n11742 = ~pi173 & n7339;
  assign n11743 = pi173 & n7347;
  assign n11744 = ~pi745 & ~n11743;
  assign n11745 = ~n11742 & n11744;
  assign n11746 = ~n59394 & ~n11745;
  assign n11747 = ~pi39 & ~n11746;
  assign n11748 = ~n11730 & n11735;
  assign n11749 = ~pi38 & ~n59395;
  assign n11750 = ~n11726 & n11749;
  assign n11751 = ~pi745 & ~n7222;
  assign n11752 = n9794 & ~n11751;
  assign n11753 = ~pi173 & ~n11752;
  assign n11754 = ~pi745 & n6822;
  assign n11755 = ~n7056 & ~n11754;
  assign n11756 = pi173 & ~n11755;
  assign n11757 = n59171 & n11756;
  assign n11758 = pi38 & ~n11757;
  assign n11759 = ~n11753 & n11758;
  assign n11760 = ~pi723 & ~n11759;
  assign n11761 = ~n11750 & n11760;
  assign n11762 = n59132 & ~n11761;
  assign n11763 = ~n11716 & n11762;
  assign n11764 = ~n11605 & ~n11763;
  assign n11765 = ~pi625 & n11764;
  assign n11766 = pi625 & n11629;
  assign n11767 = ~pi1153 & ~n11766;
  assign n11768 = ~n11765 & n11767;
  assign n11769 = ~pi608 & ~n11538;
  assign n11770 = ~n11768 & n11769;
  assign n11771 = pi625 & n11764;
  assign n11772 = ~pi625 & n11629;
  assign n11773 = pi1153 & ~n11772;
  assign n11774 = ~n11771 & n11773;
  assign n11775 = pi608 & ~n11542;
  assign n11776 = ~n11774 & n11775;
  assign n11777 = ~n11770 & ~n11776;
  assign n11778 = pi778 & ~n11777;
  assign n11779 = ~pi778 & n11764;
  assign n11780 = ~n11778 & ~n11779;
  assign n11781 = ~pi609 & ~n11780;
  assign n11782 = pi609 & n11545;
  assign n11783 = ~pi1155 & ~n11782;
  assign n11784 = ~n11781 & n11783;
  assign n11785 = ~pi660 & ~n11637;
  assign n11786 = ~n11784 & n11785;
  assign n11787 = pi609 & ~n11780;
  assign n11788 = ~pi609 & n11545;
  assign n11789 = pi1155 & ~n11788;
  assign n11790 = ~n11787 & n11789;
  assign n11791 = pi660 & ~n11641;
  assign n11792 = ~n11790 & n11791;
  assign n11793 = ~n11786 & ~n11792;
  assign n11794 = pi785 & ~n11793;
  assign n11795 = ~pi785 & ~n11780;
  assign n11796 = ~n11794 & ~n11795;
  assign n11797 = ~pi618 & ~n11796;
  assign n11798 = pi618 & n59381;
  assign n11799 = ~pi1154 & ~n11798;
  assign n11800 = ~n11797 & n11799;
  assign n11801 = ~pi627 & ~n11649;
  assign n11802 = ~n11800 & n11801;
  assign n11803 = pi618 & ~n11796;
  assign n11804 = ~pi618 & n59381;
  assign n11805 = pi1154 & ~n11804;
  assign n11806 = ~n11803 & n11805;
  assign n11807 = pi627 & ~n11653;
  assign n11808 = ~n11806 & n11807;
  assign n11809 = ~n11802 & ~n11808;
  assign n11810 = pi781 & ~n11809;
  assign n11811 = ~pi781 & ~n11796;
  assign n11812 = ~n11810 & ~n11811;
  assign n11813 = ~pi619 & ~n11812;
  assign n11814 = pi619 & ~n59382;
  assign n11815 = ~pi1159 & ~n11814;
  assign n11816 = ~n11813 & n11815;
  assign n11817 = ~pi648 & ~n11661;
  assign n11818 = ~n11816 & n11817;
  assign n11819 = pi619 & ~n11812;
  assign n11820 = ~pi619 & ~n59382;
  assign n11821 = pi1159 & ~n11820;
  assign n11822 = ~n11819 & n11821;
  assign n11823 = pi648 & ~n11665;
  assign n11824 = ~n11822 & n11823;
  assign n11825 = pi789 & ~n11824;
  assign n11826 = pi789 & ~n11818;
  assign n11827 = ~n11824 & n11826;
  assign n11828 = ~n11818 & n11825;
  assign n11829 = ~pi789 & n11812;
  assign n11830 = n59242 & ~n11829;
  assign n11831 = ~n59396 & n11830;
  assign n11832 = n7984 & n59383;
  assign n11833 = ~n7761 & n59389;
  assign n11834 = ~n11832 & ~n11833;
  assign n11835 = pi788 & ~n11834;
  assign n11836 = ~n59357 & ~n11835;
  assign n11837 = ~n11831 & n11836;
  assign n11838 = ~n11715 & ~n11837;
  assign n11839 = ~n8108 & ~n11838;
  assign n11840 = ~n11709 & ~n11839;
  assign n11841 = ~pi644 & n11840;
  assign n11842 = pi644 & ~n59386;
  assign n11843 = ~pi715 & ~n11842;
  assign n11844 = ~n11841 & n11843;
  assign n11845 = ~pi644 & n59391;
  assign n11846 = pi644 & n11520;
  assign n11847 = pi715 & ~n11846;
  assign n11848 = ~n11845 & n11847;
  assign n11849 = ~pi1160 & ~n11848;
  assign n11850 = ~n11844 & n11849;
  assign n11851 = ~n11701 & ~n11850;
  assign n11852 = pi790 & ~n11851;
  assign n11853 = pi644 & n11700;
  assign n11854 = pi790 & ~n11853;
  assign n11855 = n11840 & ~n11854;
  assign n11856 = ~n11852 & ~n11855;
  assign n11857 = n58992 & ~n11856;
  assign n11858 = ~pi173 & ~n58992;
  assign n11859 = ~pi832 & ~n11858;
  assign n11860 = ~n11857 & n11859;
  assign n11861 = ~pi173 & ~n2794;
  assign n11862 = ~n11754 & ~n11861;
  assign n11863 = ~n7875 & ~n11862;
  assign n11864 = ~pi785 & ~n11863;
  assign n11865 = n7610 & n11754;
  assign n11866 = n11863 & ~n11865;
  assign n11867 = pi1155 & ~n11866;
  assign n11868 = ~pi1155 & ~n11861;
  assign n11869 = ~n11865 & n11868;
  assign n11870 = ~n11867 & ~n11869;
  assign n11871 = pi785 & ~n11870;
  assign n11872 = ~n11864 & ~n11871;
  assign n11873 = ~pi781 & ~n11872;
  assign n11874 = ~n7890 & n11872;
  assign n11875 = pi1154 & ~n11874;
  assign n11876 = ~n7893 & n11872;
  assign n11877 = ~pi1154 & ~n11876;
  assign n11878 = ~n11875 & ~n11877;
  assign n11879 = pi781 & ~n11878;
  assign n11880 = ~n11873 & ~n11879;
  assign n11881 = ~pi789 & ~n11880;
  assign n11882 = ~pi619 & n2794;
  assign n11883 = n11880 & ~n11882;
  assign n11884 = pi1159 & ~n11883;
  assign n11885 = pi619 & n2794;
  assign n11886 = n11880 & ~n11885;
  assign n11887 = ~pi1159 & ~n11886;
  assign n11888 = ~n11884 & ~n11887;
  assign n11889 = pi789 & ~n11888;
  assign n11890 = ~n11881 & ~n11889;
  assign n11891 = n7913 & n11890;
  assign n11892 = ~n7913 & n11861;
  assign n11893 = pi626 & n11890;
  assign n11894 = ~pi626 & n11861;
  assign n11895 = pi1158 & ~n11894;
  assign n11896 = ~n11893 & n11895;
  assign n11897 = ~pi626 & n11890;
  assign n11898 = pi626 & n11861;
  assign n11899 = ~pi1158 & ~n11898;
  assign n11900 = ~n11897 & n11899;
  assign n11901 = ~n11896 & ~n11900;
  assign n11902 = ~n11891 & ~n11892;
  assign n11903 = pi788 & n59397;
  assign n11904 = ~pi788 & n11890;
  assign n11905 = ~pi788 & ~n11890;
  assign n11906 = pi788 & ~n59397;
  assign n11907 = ~n11905 & ~n11906;
  assign n11908 = ~n11903 & ~n11904;
  assign n11909 = ~n7793 & n59398;
  assign n11910 = n7793 & n11861;
  assign n11911 = ~n7872 & ~n11910;
  assign n11912 = ~n11909 & ~n11910;
  assign n11913 = ~n7872 & n11912;
  assign n11914 = ~n11909 & n11911;
  assign n11915 = ~pi723 & n7055;
  assign n11916 = ~n11861 & ~n11915;
  assign n11917 = ~pi778 & ~n11916;
  assign n11918 = ~pi625 & n11915;
  assign n11919 = ~n11916 & ~n11918;
  assign n11920 = pi1153 & ~n11919;
  assign n11921 = ~pi1153 & ~n11861;
  assign n11922 = ~n11918 & n11921;
  assign n11923 = pi778 & ~n11922;
  assign n11924 = ~n11920 & n11923;
  assign n11925 = ~n11917 & ~n11924;
  assign n11926 = ~n7949 & ~n11925;
  assign n11927 = ~n7951 & n11926;
  assign n11928 = ~n7953 & n11927;
  assign n11929 = ~n7955 & n11928;
  assign n11930 = ~n7967 & n11929;
  assign n11931 = pi647 & ~n11930;
  assign n11932 = ~pi647 & ~n11861;
  assign n11933 = ~n11931 & ~n11932;
  assign n11934 = n7832 & ~n11933;
  assign n11935 = ~pi647 & n11930;
  assign n11936 = pi647 & n11861;
  assign n11937 = ~pi1157 & ~n11936;
  assign n11938 = ~n11935 & n11937;
  assign n11939 = pi630 & n11938;
  assign n11940 = ~n11934 & ~n11939;
  assign n11941 = ~n59399 & n11940;
  assign n11942 = pi787 & ~n11941;
  assign n11943 = n7984 & n11928;
  assign n11944 = ~n7761 & n59397;
  assign n11945 = ~n11943 & ~n11944;
  assign n11946 = pi788 & ~n11945;
  assign n11947 = ~n6701 & ~n11916;
  assign n11948 = pi625 & n11947;
  assign n11949 = n11862 & ~n11947;
  assign n11950 = ~n11948 & ~n11949;
  assign n11951 = n11921 & ~n11950;
  assign n11952 = ~pi608 & ~n11920;
  assign n11953 = ~n11951 & n11952;
  assign n11954 = pi1153 & n11862;
  assign n11955 = ~n11948 & n11954;
  assign n11956 = pi608 & ~n11922;
  assign n11957 = ~n11955 & n11956;
  assign n11958 = ~n11953 & ~n11957;
  assign n11959 = pi778 & ~n11958;
  assign n11960 = ~pi778 & ~n11949;
  assign n11961 = ~n11959 & ~n11960;
  assign n11962 = ~pi609 & ~n11961;
  assign n11963 = pi609 & ~n11925;
  assign n11964 = ~pi1155 & ~n11963;
  assign n11965 = ~n11962 & n11964;
  assign n11966 = ~pi660 & ~n11867;
  assign n11967 = ~n11965 & n11966;
  assign n11968 = pi609 & ~n11961;
  assign n11969 = ~pi609 & ~n11925;
  assign n11970 = pi1155 & ~n11969;
  assign n11971 = ~n11968 & n11970;
  assign n11972 = pi660 & ~n11869;
  assign n11973 = ~n11971 & n11972;
  assign n11974 = ~n11967 & ~n11973;
  assign n11975 = pi785 & ~n11974;
  assign n11976 = ~pi785 & ~n11961;
  assign n11977 = ~n11975 & ~n11976;
  assign n11978 = ~pi618 & ~n11977;
  assign n11979 = pi618 & n11926;
  assign n11980 = ~pi1154 & ~n11979;
  assign n11981 = ~n11978 & n11980;
  assign n11982 = ~pi627 & ~n11875;
  assign n11983 = ~n11981 & n11982;
  assign n11984 = pi618 & ~n11977;
  assign n11985 = ~pi618 & n11926;
  assign n11986 = pi1154 & ~n11985;
  assign n11987 = ~n11984 & n11986;
  assign n11988 = pi627 & ~n11877;
  assign n11989 = ~n11987 & n11988;
  assign n11990 = ~n11983 & ~n11989;
  assign n11991 = pi781 & ~n11990;
  assign n11992 = ~pi781 & ~n11977;
  assign n11993 = ~n11991 & ~n11992;
  assign n11994 = ~pi619 & ~n11993;
  assign n11995 = pi619 & n11927;
  assign n11996 = ~pi1159 & ~n11995;
  assign n11997 = ~n11994 & n11996;
  assign n11998 = ~pi648 & ~n11884;
  assign n11999 = ~n11997 & n11998;
  assign n12000 = pi619 & ~n11993;
  assign n12001 = ~pi619 & n11927;
  assign n12002 = pi1159 & ~n12001;
  assign n12003 = ~n12000 & n12002;
  assign n12004 = pi648 & ~n11887;
  assign n12005 = ~n12003 & n12004;
  assign n12006 = pi789 & ~n12005;
  assign n12007 = pi789 & ~n11999;
  assign n12008 = ~n12005 & n12007;
  assign n12009 = ~n11999 & n12006;
  assign n12010 = ~pi789 & n11993;
  assign n12011 = n59242 & ~n12010;
  assign n12012 = ~n59400 & n12011;
  assign n12013 = ~n11946 & ~n12012;
  assign n12014 = ~n59357 & ~n12013;
  assign n12015 = n7957 & n59398;
  assign n12016 = n8065 & n11929;
  assign n12017 = pi629 & ~n12016;
  assign n12018 = ~n12015 & n12017;
  assign n12019 = n7958 & n59398;
  assign n12020 = n8074 & n11929;
  assign n12021 = ~pi629 & ~n12020;
  assign n12022 = ~n12019 & n12021;
  assign n12023 = pi792 & ~n12022;
  assign n12024 = ~n12019 & ~n12020;
  assign n12025 = ~pi629 & ~n12024;
  assign n12026 = ~n12015 & ~n12016;
  assign n12027 = pi629 & ~n12026;
  assign n12028 = ~n12025 & ~n12027;
  assign n12029 = pi792 & ~n12028;
  assign n12030 = pi792 & ~n12018;
  assign n12031 = ~n12022 & n12030;
  assign n12032 = ~n12018 & n12023;
  assign n12033 = ~n8108 & ~n59401;
  assign n12034 = ~n12014 & n12033;
  assign n12035 = ~n11942 & ~n12034;
  assign n12036 = pi644 & n12035;
  assign n12037 = ~pi787 & ~n11930;
  assign n12038 = pi1157 & ~n11933;
  assign n12039 = ~n11938 & ~n12038;
  assign n12040 = pi787 & ~n12039;
  assign n12041 = ~n12037 & ~n12040;
  assign n12042 = ~pi644 & n12041;
  assign n12043 = pi715 & ~n12042;
  assign n12044 = ~n12036 & n12043;
  assign n12045 = ~n11491 & n11861;
  assign n12046 = ~n7835 & n11909;
  assign n12047 = ~n7835 & ~n11912;
  assign n12048 = n7835 & n11861;
  assign n12049 = ~n12047 & ~n12048;
  assign n12050 = ~n12045 & ~n12046;
  assign n12051 = pi644 & ~n59402;
  assign n12052 = ~pi644 & n11861;
  assign n12053 = ~pi715 & ~n12052;
  assign n12054 = ~n12051 & n12053;
  assign n12055 = pi1160 & ~n12054;
  assign n12056 = ~n12044 & n12055;
  assign n12057 = ~pi644 & n12035;
  assign n12058 = pi644 & n12041;
  assign n12059 = ~pi715 & ~n12058;
  assign n12060 = ~n12057 & n12059;
  assign n12061 = ~pi644 & ~n59402;
  assign n12062 = pi644 & n11861;
  assign n12063 = pi715 & ~n12062;
  assign n12064 = ~n12061 & n12063;
  assign n12065 = ~pi1160 & ~n12064;
  assign n12066 = ~n12060 & n12065;
  assign n12067 = ~n12056 & ~n12066;
  assign n12068 = pi790 & ~n12067;
  assign n12069 = ~pi790 & n12035;
  assign n12070 = pi832 & ~n12069;
  assign n12071 = ~n12068 & n12070;
  assign po330 = ~n11860 & ~n12071;
  assign n12073 = pi174 & ~n59132;
  assign n12074 = ~pi759 & ~n6654;
  assign n12075 = pi759 & n59163;
  assign n12076 = ~n12074 & ~n12075;
  assign n12077 = pi39 & ~n12076;
  assign n12078 = pi759 & n59157;
  assign n12079 = ~pi759 & n59147;
  assign n12080 = ~pi39 & ~n12079;
  assign n12081 = ~n12078 & n12080;
  assign n12082 = ~n12077 & ~n12081;
  assign n12083 = pi174 & ~n12082;
  assign n12084 = ~pi174 & pi759;
  assign n12085 = n6855 & n12084;
  assign n12086 = ~n12083 & ~n12085;
  assign n12087 = ~pi38 & ~n12086;
  assign n12088 = pi759 & n6701;
  assign n12089 = n6863 & ~n12088;
  assign n12090 = ~pi174 & ~n6863;
  assign n12091 = pi38 & ~n12090;
  assign n12092 = ~n12089 & n12091;
  assign n12093 = ~n12087 & ~n12092;
  assign n12094 = n59132 & ~n12093;
  assign n12095 = ~n12073 & ~n12094;
  assign n12096 = ~n7597 & ~n12095;
  assign n12097 = pi174 & ~n7560;
  assign n12098 = n7597 & n12097;
  assign n12099 = n7597 & ~n12097;
  assign n12100 = ~n7597 & n12095;
  assign n12101 = ~n12099 & ~n12100;
  assign n12102 = ~n12096 & ~n12098;
  assign n12103 = ~pi785 & n59403;
  assign n12104 = pi609 & ~n59403;
  assign n12105 = ~pi609 & ~n12097;
  assign n12106 = pi1155 & ~n12105;
  assign n12107 = ~n12104 & n12106;
  assign n12108 = ~pi609 & ~n59403;
  assign n12109 = pi609 & ~n12097;
  assign n12110 = ~pi1155 & ~n12109;
  assign n12111 = ~n12108 & n12110;
  assign n12112 = ~n12107 & ~n12111;
  assign n12113 = pi785 & ~n12112;
  assign n12114 = ~n12103 & ~n12113;
  assign n12115 = ~pi781 & ~n12114;
  assign n12116 = pi618 & n12114;
  assign n12117 = ~pi618 & ~n12097;
  assign n12118 = pi1154 & ~n12117;
  assign n12119 = ~n12116 & n12118;
  assign n12120 = ~pi618 & n12114;
  assign n12121 = pi618 & ~n12097;
  assign n12122 = ~pi1154 & ~n12121;
  assign n12123 = ~n12120 & n12122;
  assign n12124 = ~n12119 & ~n12123;
  assign n12125 = pi781 & ~n12124;
  assign n12126 = ~n12115 & ~n12125;
  assign n12127 = ~pi789 & ~n12126;
  assign n12128 = pi619 & n12126;
  assign n12129 = ~pi619 & ~n12097;
  assign n12130 = pi1159 & ~n12129;
  assign n12131 = ~n12128 & n12130;
  assign n12132 = ~pi619 & n12126;
  assign n12133 = pi619 & ~n12097;
  assign n12134 = ~pi1159 & ~n12133;
  assign n12135 = ~n12132 & n12134;
  assign n12136 = ~n12131 & ~n12135;
  assign n12137 = pi789 & ~n12136;
  assign n12138 = ~n12127 & ~n12137;
  assign n12139 = ~n7761 & ~n7983;
  assign n12140 = n12138 & n12139;
  assign n12141 = n59231 & ~n12097;
  assign n12142 = pi696 & n59132;
  assign n12143 = ~n12097 & ~n12142;
  assign n12144 = pi174 & ~n8249;
  assign n12145 = ~pi174 & ~n59251;
  assign n12146 = ~pi38 & ~n12145;
  assign n12147 = ~n12144 & n12146;
  assign n12148 = n10432 & ~n12090;
  assign n12149 = n12142 & ~n12148;
  assign n12150 = ~n12147 & n12149;
  assign n12151 = ~n12143 & ~n12150;
  assign n12152 = ~pi778 & n12151;
  assign n12153 = pi625 & ~n12151;
  assign n12154 = ~pi625 & ~n12097;
  assign n12155 = pi1153 & ~n12154;
  assign n12156 = ~n12153 & n12155;
  assign n12157 = ~pi625 & ~n12151;
  assign n12158 = pi625 & ~n12097;
  assign n12159 = ~pi1153 & ~n12158;
  assign n12160 = ~n12157 & n12159;
  assign n12161 = ~n12156 & ~n12160;
  assign n12162 = pi778 & ~n12161;
  assign n12163 = ~n12152 & ~n12162;
  assign n12164 = ~n59229 & ~n12163;
  assign n12165 = n59229 & n12097;
  assign n12166 = n59229 & ~n12097;
  assign n12167 = ~n59229 & n12163;
  assign n12168 = ~n12166 & ~n12167;
  assign n12169 = ~n12164 & ~n12165;
  assign n12170 = ~n59231 & ~n59404;
  assign n12171 = ~n59231 & n59404;
  assign n12172 = n59231 & n12097;
  assign n12173 = ~n12171 & ~n12172;
  assign n12174 = ~n12141 & ~n12170;
  assign n12175 = ~n7716 & ~n59405;
  assign n12176 = n7716 & n12097;
  assign n12177 = n7716 & ~n12097;
  assign n12178 = ~n7716 & n59405;
  assign n12179 = ~n12177 & ~n12178;
  assign n12180 = ~n12175 & ~n12176;
  assign n12181 = ~pi641 & n59406;
  assign n12182 = pi641 & n12097;
  assign n12183 = n7912 & ~n12182;
  assign n12184 = ~n12181 & n12183;
  assign n12185 = pi641 & n59406;
  assign n12186 = ~pi641 & n12097;
  assign n12187 = n7911 & ~n12186;
  assign n12188 = ~n12185 & n12187;
  assign n12189 = ~n12184 & ~n12188;
  assign n12190 = ~n12140 & n12189;
  assign n12191 = pi788 & ~n12190;
  assign n12192 = ~pi696 & n12087;
  assign n12193 = pi174 & ~n59177;
  assign n12194 = ~pi174 & ~n7111;
  assign n12195 = ~pi759 & ~n12194;
  assign n12196 = ~n12193 & n12195;
  assign n12197 = ~pi174 & ~n7188;
  assign n12198 = pi174 & n59203;
  assign n12199 = pi759 & ~n12198;
  assign n12200 = ~n12197 & n12199;
  assign n12201 = pi39 & ~n12200;
  assign n12202 = ~n12196 & n12201;
  assign n12203 = ~pi174 & ~n7333;
  assign n12204 = pi174 & ~n7310;
  assign n12205 = ~pi759 & ~n12204;
  assign n12206 = ~pi759 & ~n12203;
  assign n12207 = ~n12204 & n12206;
  assign n12208 = ~n12203 & n12205;
  assign n12209 = pi174 & n7339;
  assign n12210 = ~pi174 & n7347;
  assign n12211 = pi759 & ~n12210;
  assign n12212 = ~n12209 & n12211;
  assign n12213 = ~pi39 & ~n12212;
  assign n12214 = ~n59407 & n12213;
  assign n12215 = ~pi38 & ~n12214;
  assign n12216 = ~n12202 & n12215;
  assign n12217 = ~n9801 & ~n12216;
  assign n12218 = pi696 & ~n12217;
  assign n12219 = ~n12092 & ~n12218;
  assign n12220 = ~n12192 & n12219;
  assign n12221 = ~pi696 & n12093;
  assign n12222 = pi696 & ~n9801;
  assign n12223 = ~n12092 & n12222;
  assign n12224 = ~n12216 & n12223;
  assign n12225 = n59132 & ~n12224;
  assign n12226 = ~n12221 & n12225;
  assign n12227 = n59132 & ~n12220;
  assign n12228 = ~n12073 & ~n59408;
  assign n12229 = ~pi625 & n12228;
  assign n12230 = pi625 & n12095;
  assign n12231 = ~pi1153 & ~n12230;
  assign n12232 = ~n12229 & n12231;
  assign n12233 = ~pi608 & ~n12156;
  assign n12234 = ~n12232 & n12233;
  assign n12235 = pi625 & n12228;
  assign n12236 = ~pi625 & n12095;
  assign n12237 = pi1153 & ~n12236;
  assign n12238 = ~n12235 & n12237;
  assign n12239 = pi608 & ~n12160;
  assign n12240 = ~n12238 & n12239;
  assign n12241 = ~n12234 & ~n12240;
  assign n12242 = pi778 & ~n12241;
  assign n12243 = ~pi778 & n12228;
  assign n12244 = ~n12242 & ~n12243;
  assign n12245 = ~pi609 & ~n12244;
  assign n12246 = pi609 & n12163;
  assign n12247 = ~pi1155 & ~n12246;
  assign n12248 = ~n12245 & n12247;
  assign n12249 = ~pi660 & ~n12107;
  assign n12250 = ~n12248 & n12249;
  assign n12251 = pi609 & ~n12244;
  assign n12252 = ~pi609 & n12163;
  assign n12253 = pi1155 & ~n12252;
  assign n12254 = ~n12251 & n12253;
  assign n12255 = pi660 & ~n12111;
  assign n12256 = ~n12254 & n12255;
  assign n12257 = ~n12250 & ~n12256;
  assign n12258 = pi785 & ~n12257;
  assign n12259 = ~pi785 & ~n12244;
  assign n12260 = ~n12258 & ~n12259;
  assign n12261 = ~pi618 & ~n12260;
  assign n12262 = pi618 & ~n59404;
  assign n12263 = ~pi1154 & ~n12262;
  assign n12264 = ~n12261 & n12263;
  assign n12265 = ~pi627 & ~n12119;
  assign n12266 = ~n12264 & n12265;
  assign n12267 = pi618 & ~n12260;
  assign n12268 = ~pi618 & ~n59404;
  assign n12269 = pi1154 & ~n12268;
  assign n12270 = ~n12267 & n12269;
  assign n12271 = pi627 & ~n12123;
  assign n12272 = ~n12270 & n12271;
  assign n12273 = ~n12266 & ~n12272;
  assign n12274 = pi781 & ~n12273;
  assign n12275 = ~pi781 & ~n12260;
  assign n12276 = ~n12274 & ~n12275;
  assign n12277 = ~pi619 & ~n12276;
  assign n12278 = pi619 & n59405;
  assign n12279 = ~pi1159 & ~n12278;
  assign n12280 = ~n12277 & n12279;
  assign n12281 = ~pi648 & ~n12131;
  assign n12282 = ~n12280 & n12281;
  assign n12283 = pi619 & ~n12276;
  assign n12284 = ~pi619 & n59405;
  assign n12285 = pi1159 & ~n12284;
  assign n12286 = ~n12283 & n12285;
  assign n12287 = pi648 & ~n12135;
  assign n12288 = ~n12286 & n12287;
  assign n12289 = pi789 & ~n12288;
  assign n12290 = ~n12282 & n12289;
  assign n12291 = ~pi789 & n12276;
  assign n12292 = n59242 & ~n12291;
  assign n12293 = ~n12290 & n12292;
  assign n12294 = ~n12282 & ~n12288;
  assign n12295 = pi789 & ~n12294;
  assign n12296 = ~pi789 & ~n12276;
  assign n12297 = ~n12295 & ~n12296;
  assign n12298 = ~pi788 & n12297;
  assign n12299 = ~pi626 & n12297;
  assign n12300 = pi626 & n59406;
  assign n12301 = ~pi641 & ~n12300;
  assign n12302 = ~n12299 & n12301;
  assign n12303 = ~pi626 & ~n12138;
  assign n12304 = pi626 & n12097;
  assign n12305 = pi641 & ~n12304;
  assign n12306 = ~n12303 & n12305;
  assign n12307 = ~pi1158 & ~n12306;
  assign n12308 = ~n12302 & n12307;
  assign n12309 = pi626 & n12297;
  assign n12310 = ~pi626 & n59406;
  assign n12311 = pi641 & ~n12310;
  assign n12312 = ~n12309 & n12311;
  assign n12313 = pi626 & ~n12138;
  assign n12314 = ~pi626 & n12097;
  assign n12315 = ~pi641 & ~n12314;
  assign n12316 = ~n12313 & n12315;
  assign n12317 = pi1158 & ~n12316;
  assign n12318 = ~n12312 & n12317;
  assign n12319 = ~n12308 & ~n12318;
  assign n12320 = pi788 & ~n12319;
  assign n12321 = ~n12298 & ~n12320;
  assign n12322 = ~n12191 & ~n12293;
  assign n12323 = ~pi628 & n59409;
  assign n12324 = ~n8054 & ~n12138;
  assign n12325 = n8054 & n12097;
  assign n12326 = ~n12324 & ~n12325;
  assign n12327 = pi628 & n12326;
  assign n12328 = ~pi1156 & ~n12327;
  assign n12329 = ~n12323 & n12328;
  assign n12330 = n7762 & ~n12097;
  assign n12331 = ~n7762 & ~n59406;
  assign n12332 = ~n7762 & n59406;
  assign n12333 = n7762 & n12097;
  assign n12334 = ~n12332 & ~n12333;
  assign n12335 = ~n12330 & ~n12331;
  assign n12336 = pi628 & n59410;
  assign n12337 = ~pi628 & ~n12097;
  assign n12338 = pi1156 & ~n12337;
  assign n12339 = ~n12336 & n12338;
  assign n12340 = ~pi629 & ~n12339;
  assign n12341 = ~n12329 & n12340;
  assign n12342 = pi628 & n59409;
  assign n12343 = ~pi628 & n12326;
  assign n12344 = pi1156 & ~n12343;
  assign n12345 = ~n12342 & n12344;
  assign n12346 = ~pi628 & n59410;
  assign n12347 = pi628 & ~n12097;
  assign n12348 = ~pi1156 & ~n12347;
  assign n12349 = ~n12346 & n12348;
  assign n12350 = pi629 & ~n12349;
  assign n12351 = ~n12345 & n12350;
  assign n12352 = ~n12341 & ~n12351;
  assign n12353 = pi792 & ~n12352;
  assign n12354 = ~pi792 & n59409;
  assign n12355 = ~n12353 & ~n12354;
  assign n12356 = ~pi647 & ~n12355;
  assign n12357 = ~n7793 & ~n12326;
  assign n12358 = n7793 & n12097;
  assign n12359 = ~n12357 & ~n12358;
  assign n12360 = pi647 & n12359;
  assign n12361 = ~pi1157 & ~n12360;
  assign n12362 = ~n12356 & n12361;
  assign n12363 = ~pi792 & ~n59410;
  assign n12364 = ~n12339 & ~n12349;
  assign n12365 = pi792 & ~n12364;
  assign n12366 = ~n12363 & ~n12365;
  assign n12367 = pi647 & n12366;
  assign n12368 = ~pi647 & ~n12097;
  assign n12369 = pi1157 & ~n12368;
  assign n12370 = ~n12367 & n12369;
  assign n12371 = ~pi630 & ~n12370;
  assign n12372 = ~n12362 & n12371;
  assign n12373 = pi647 & ~n12355;
  assign n12374 = ~pi647 & n12359;
  assign n12375 = pi1157 & ~n12374;
  assign n12376 = ~n12373 & n12375;
  assign n12377 = ~pi647 & n12366;
  assign n12378 = pi647 & ~n12097;
  assign n12379 = ~pi1157 & ~n12378;
  assign n12380 = ~n12377 & n12379;
  assign n12381 = pi630 & ~n12380;
  assign n12382 = ~n12376 & n12381;
  assign n12383 = ~n12372 & ~n12382;
  assign n12384 = pi787 & ~n12383;
  assign n12385 = ~pi787 & ~n12355;
  assign n12386 = ~n12384 & ~n12385;
  assign n12387 = pi644 & ~n12386;
  assign n12388 = ~pi787 & ~n12366;
  assign n12389 = ~n12370 & ~n12380;
  assign n12390 = pi787 & ~n12389;
  assign n12391 = ~n12388 & ~n12390;
  assign n12392 = ~pi644 & n12391;
  assign n12393 = pi715 & ~n12392;
  assign n12394 = ~n12387 & n12393;
  assign n12395 = ~n7835 & ~n12359;
  assign n12396 = n7835 & n12097;
  assign n12397 = n7835 & ~n12097;
  assign n12398 = ~n7835 & n12359;
  assign n12399 = ~n12397 & ~n12398;
  assign n12400 = ~n12395 & ~n12396;
  assign n12401 = pi644 & ~n59411;
  assign n12402 = ~pi644 & ~n12097;
  assign n12403 = ~pi715 & ~n12402;
  assign n12404 = ~n12401 & n12403;
  assign n12405 = pi1160 & ~n12404;
  assign n12406 = ~n12394 & n12405;
  assign n12407 = ~pi644 & ~n12386;
  assign n12408 = pi644 & n12391;
  assign n12409 = ~pi715 & ~n12408;
  assign n12410 = ~n12407 & n12409;
  assign n12411 = ~pi644 & ~n59411;
  assign n12412 = pi644 & ~n12097;
  assign n12413 = pi715 & ~n12412;
  assign n12414 = ~n12411 & n12413;
  assign n12415 = ~pi1160 & ~n12414;
  assign n12416 = ~n12410 & n12415;
  assign n12417 = pi790 & ~n12416;
  assign n12418 = pi790 & ~n12406;
  assign n12419 = ~n12416 & n12418;
  assign n12420 = ~n12406 & n12417;
  assign n12421 = ~pi790 & n12386;
  assign n12422 = n4441 & ~n12421;
  assign n12423 = ~n59412 & n12422;
  assign n12424 = ~pi174 & ~n4441;
  assign n12425 = ~pi57 & ~n12424;
  assign n12426 = ~n12423 & n12425;
  assign n12427 = pi57 & pi174;
  assign n12428 = ~pi832 & ~n12427;
  assign n12429 = ~n12426 & n12428;
  assign n12430 = pi696 & n7055;
  assign n12431 = pi696 & n7056;
  assign n12432 = ~n6701 & n12430;
  assign n12433 = pi174 & ~n2794;
  assign n12434 = pi759 & n6822;
  assign n12435 = ~n12433 & ~n12434;
  assign n12436 = ~n59413 & n12435;
  assign n12437 = pi625 & n12430;
  assign n12438 = pi625 & n59413;
  assign n12439 = ~n6701 & n12437;
  assign n12440 = ~n12436 & ~n59414;
  assign n12441 = ~pi1153 & ~n12440;
  assign n12442 = pi1153 & ~n12433;
  assign n12443 = ~n12437 & n12442;
  assign n12444 = ~pi608 & ~n12443;
  assign n12445 = ~n12441 & n12444;
  assign n12446 = pi1153 & n12435;
  assign n12447 = ~n12434 & n12442;
  assign n12448 = ~n59414 & n59415;
  assign n12449 = ~n12430 & ~n12433;
  assign n12450 = ~n12437 & ~n12449;
  assign n12451 = ~pi1153 & ~n12450;
  assign n12452 = pi608 & ~n12451;
  assign n12453 = ~n12448 & n12452;
  assign n12454 = ~n12445 & ~n12453;
  assign n12455 = pi778 & ~n12454;
  assign n12456 = ~pi778 & ~n12436;
  assign n12457 = ~n12455 & ~n12456;
  assign n12458 = ~pi609 & ~n12457;
  assign n12459 = ~pi778 & n12449;
  assign n12460 = ~n12443 & ~n12451;
  assign n12461 = pi778 & ~n12460;
  assign n12462 = ~n12459 & ~n12461;
  assign n12463 = pi609 & n12462;
  assign n12464 = ~pi1155 & ~n12463;
  assign n12465 = ~n12458 & n12464;
  assign n12466 = n7598 & n12434;
  assign n12467 = pi1155 & ~n12433;
  assign n12468 = ~n12466 & n12467;
  assign n12469 = ~pi660 & ~n12468;
  assign n12470 = ~n12465 & n12469;
  assign n12471 = pi609 & ~n12457;
  assign n12472 = ~pi609 & n12462;
  assign n12473 = pi1155 & ~n12472;
  assign n12474 = ~n12471 & n12473;
  assign n12475 = n7610 & n12434;
  assign n12476 = ~pi1155 & ~n12433;
  assign n12477 = ~n12475 & n12476;
  assign n12478 = pi660 & ~n12477;
  assign n12479 = ~n12474 & n12478;
  assign n12480 = ~n12470 & ~n12479;
  assign n12481 = pi785 & ~n12480;
  assign n12482 = ~pi785 & ~n12457;
  assign n12483 = ~n12481 & ~n12482;
  assign n12484 = ~pi618 & ~n12483;
  assign n12485 = ~n59229 & n12462;
  assign n12486 = ~n12433 & ~n12485;
  assign n12487 = pi618 & ~n12486;
  assign n12488 = ~pi1154 & ~n12487;
  assign n12489 = ~n12484 & n12488;
  assign n12490 = ~n59346 & n12434;
  assign n12491 = n10835 & n12490;
  assign n12492 = pi1154 & ~n12433;
  assign n12493 = ~n12491 & n12492;
  assign n12494 = ~pi627 & ~n12493;
  assign n12495 = ~n12489 & n12494;
  assign n12496 = pi618 & ~n12483;
  assign n12497 = ~pi618 & ~n12486;
  assign n12498 = pi1154 & ~n12497;
  assign n12499 = ~n12496 & n12498;
  assign n12500 = n10837 & n12490;
  assign n12501 = ~pi1154 & ~n12433;
  assign n12502 = ~n12500 & n12501;
  assign n12503 = pi627 & ~n12502;
  assign n12504 = ~n12499 & n12503;
  assign n12505 = ~n12495 & ~n12504;
  assign n12506 = pi781 & ~n12505;
  assign n12507 = ~pi781 & ~n12483;
  assign n12508 = pi648 & n10738;
  assign n12509 = ~pi648 & n10739;
  assign n12510 = ~n12508 & ~n12509;
  assign n12511 = n7715 & n12510;
  assign n12512 = n7715 & n10740;
  assign n12513 = pi789 & ~n59416;
  assign n12514 = ~n12507 & ~n12513;
  assign n12515 = ~n12506 & n12514;
  assign n12516 = n9554 & n12462;
  assign n12517 = ~n12510 & ~n12516;
  assign n12518 = ~n59347 & n12490;
  assign n12519 = ~n7715 & ~n12518;
  assign n12520 = ~n7597 & n10740;
  assign n12521 = ~n7715 & ~n12520;
  assign n12522 = n10884 & n12518;
  assign n12523 = n7714 & ~n12522;
  assign n12524 = n10874 & n12518;
  assign n12525 = n7713 & ~n12524;
  assign n12526 = ~n12523 & ~n12525;
  assign n12527 = ~n12519 & ~n12521;
  assign n12528 = ~n12517 & n59417;
  assign n12529 = pi789 & ~n12433;
  assign n12530 = ~n12528 & n12529;
  assign n12531 = n59242 & ~n12530;
  assign n12532 = ~n12515 & n12531;
  assign n12533 = ~n7716 & n12516;
  assign n12534 = ~n12433 & ~n12533;
  assign n12535 = n7911 & ~n12534;
  assign n12536 = n59348 & n12490;
  assign n12537 = ~pi626 & n12536;
  assign n12538 = ~n12433 & ~n12537;
  assign n12539 = ~pi1158 & ~n12538;
  assign n12540 = pi641 & ~n12539;
  assign n12541 = ~n12535 & n12540;
  assign n12542 = n7912 & ~n12534;
  assign n12543 = pi626 & n12536;
  assign n12544 = ~n12433 & ~n12543;
  assign n12545 = pi1158 & ~n12544;
  assign n12546 = ~pi641 & ~n12545;
  assign n12547 = ~n12542 & n12546;
  assign n12548 = pi788 & ~n12547;
  assign n12549 = pi788 & ~n12541;
  assign n12550 = ~n12547 & n12549;
  assign n12551 = ~n12541 & n12548;
  assign n12552 = ~n59357 & ~n59418;
  assign n12553 = ~n12532 & n12552;
  assign n12554 = ~n8054 & n12536;
  assign n12555 = ~pi629 & n12554;
  assign n12556 = pi628 & ~n12555;
  assign n12557 = ~n7762 & n12533;
  assign n12558 = n9652 & n12462;
  assign n12559 = pi629 & ~n59419;
  assign n12560 = ~pi628 & n59419;
  assign n12561 = pi629 & ~n12560;
  assign n12562 = pi628 & ~n12554;
  assign n12563 = ~n12561 & ~n12562;
  assign n12564 = ~n12556 & ~n12559;
  assign n12565 = ~pi1156 & ~n59420;
  assign n12566 = pi628 & n59419;
  assign n12567 = ~pi628 & ~n12554;
  assign n12568 = pi629 & ~n12567;
  assign n12569 = pi1156 & ~n12568;
  assign n12570 = ~n12566 & n12569;
  assign n12571 = ~n12565 & ~n12570;
  assign n12572 = pi792 & ~n12433;
  assign n12573 = ~n12571 & n12572;
  assign n12574 = ~n12553 & ~n12573;
  assign n12575 = ~n8108 & ~n12574;
  assign n12576 = ~n7793 & n12554;
  assign n12577 = ~pi630 & n12576;
  assign n12578 = pi647 & ~n12577;
  assign n12579 = ~n59240 & n59419;
  assign n12580 = pi630 & ~n12579;
  assign n12581 = ~pi647 & n12579;
  assign n12582 = pi630 & ~n12581;
  assign n12583 = pi647 & ~n12576;
  assign n12584 = ~n12582 & ~n12583;
  assign n12585 = ~n12578 & ~n12580;
  assign n12586 = ~pi1157 & ~n59421;
  assign n12587 = ~pi630 & ~n12579;
  assign n12588 = pi647 & ~n12587;
  assign n12589 = pi630 & n12576;
  assign n12590 = pi1157 & ~n12589;
  assign n12591 = ~n12588 & n12590;
  assign n12592 = ~n12586 & ~n12591;
  assign n12593 = pi787 & ~n12433;
  assign n12594 = ~n12592 & n12593;
  assign n12595 = ~n12575 & ~n12594;
  assign n12596 = pi644 & n12595;
  assign n12597 = ~n9743 & n12579;
  assign n12598 = ~n12433 & ~n12597;
  assign n12599 = ~pi644 & ~n12598;
  assign n12600 = pi715 & ~n12599;
  assign n12601 = ~n12596 & n12600;
  assign n12602 = ~n8054 & n11491;
  assign n12603 = pi644 & n12602;
  assign n12604 = n11491 & n12554;
  assign n12605 = pi644 & n12604;
  assign n12606 = n12536 & n12603;
  assign n12607 = ~pi715 & ~n12433;
  assign n12608 = ~n59422 & n12607;
  assign n12609 = pi1160 & ~n12608;
  assign n12610 = ~n12601 & n12609;
  assign n12611 = ~pi644 & n12595;
  assign n12612 = pi644 & ~n12598;
  assign n12613 = ~pi715 & ~n12612;
  assign n12614 = ~n12611 & n12613;
  assign n12615 = ~pi644 & n12602;
  assign n12616 = ~pi644 & n12604;
  assign n12617 = n12536 & n12615;
  assign n12618 = pi715 & ~n12433;
  assign n12619 = ~n59423 & n12618;
  assign n12620 = ~pi1160 & ~n12619;
  assign n12621 = ~n12614 & n12620;
  assign n12622 = ~n12610 & ~n12621;
  assign n12623 = pi790 & ~n12622;
  assign n12624 = ~pi790 & n12595;
  assign n12625 = pi832 & ~n12624;
  assign n12626 = ~n12623 & n12625;
  assign po331 = ~n12429 & ~n12626;
  assign n12628 = ~pi175 & ~n2794;
  assign n12629 = pi766 & n6822;
  assign n12630 = ~n12628 & ~n12629;
  assign n12631 = ~n7875 & ~n12630;
  assign n12632 = ~pi785 & ~n12631;
  assign n12633 = n7610 & n12629;
  assign n12634 = n12631 & ~n12633;
  assign n12635 = pi1155 & ~n12634;
  assign n12636 = ~pi1155 & ~n12628;
  assign n12637 = ~n12633 & n12636;
  assign n12638 = ~n12635 & ~n12637;
  assign n12639 = pi785 & ~n12638;
  assign n12640 = ~n12632 & ~n12639;
  assign n12641 = ~pi781 & ~n12640;
  assign n12642 = ~n7890 & n12640;
  assign n12643 = pi1154 & ~n12642;
  assign n12644 = ~n7893 & n12640;
  assign n12645 = ~pi1154 & ~n12644;
  assign n12646 = ~n12643 & ~n12645;
  assign n12647 = pi781 & ~n12646;
  assign n12648 = ~n12641 & ~n12647;
  assign n12649 = ~pi789 & ~n12648;
  assign n12650 = ~n11882 & n12648;
  assign n12651 = pi1159 & ~n12650;
  assign n12652 = ~n11885 & n12648;
  assign n12653 = ~pi1159 & ~n12652;
  assign n12654 = ~n12651 & ~n12653;
  assign n12655 = pi789 & ~n12654;
  assign n12656 = ~n12649 & ~n12655;
  assign n12657 = ~n8054 & ~n12656;
  assign n12658 = n8054 & ~n12628;
  assign n12659 = ~n8054 & n12656;
  assign n12660 = n8054 & n12628;
  assign n12661 = ~n12659 & ~n12660;
  assign n12662 = ~n12657 & ~n12658;
  assign n12663 = ~n7793 & ~n59424;
  assign n12664 = n7793 & n12628;
  assign n12665 = ~n7872 & ~n12664;
  assign n12666 = ~n12663 & ~n12664;
  assign n12667 = ~n7872 & n12666;
  assign n12668 = ~n12663 & n12665;
  assign n12669 = pi700 & n7055;
  assign n12670 = ~n12628 & ~n12669;
  assign n12671 = ~pi778 & ~n12670;
  assign n12672 = ~pi625 & n12669;
  assign n12673 = ~n12670 & ~n12672;
  assign n12674 = pi1153 & ~n12673;
  assign n12675 = ~pi1153 & ~n12628;
  assign n12676 = ~n12672 & n12675;
  assign n12677 = pi778 & ~n12676;
  assign n12678 = ~n12674 & n12677;
  assign n12679 = ~n12671 & ~n12678;
  assign n12680 = ~n7949 & ~n12679;
  assign n12681 = ~n7951 & n12680;
  assign n12682 = ~n7953 & n12681;
  assign n12683 = ~n7955 & n12682;
  assign n12684 = ~n7967 & n12683;
  assign n12685 = pi647 & ~n12684;
  assign n12686 = ~pi647 & ~n12628;
  assign n12687 = ~n12685 & ~n12686;
  assign n12688 = n7832 & ~n12687;
  assign n12689 = ~pi647 & n12684;
  assign n12690 = pi647 & n12628;
  assign n12691 = ~pi1157 & ~n12690;
  assign n12692 = ~n12689 & n12691;
  assign n12693 = pi630 & n12692;
  assign n12694 = ~n12688 & ~n12693;
  assign n12695 = ~n59425 & n12694;
  assign n12696 = pi787 & ~n12695;
  assign n12697 = ~pi626 & ~n12656;
  assign n12698 = pi626 & ~n12628;
  assign n12699 = n7760 & ~n12698;
  assign n12700 = ~n12697 & n12699;
  assign n12701 = n7984 & n12682;
  assign n12702 = pi626 & ~n12656;
  assign n12703 = ~pi626 & ~n12628;
  assign n12704 = n7759 & ~n12703;
  assign n12705 = ~n12702 & n12704;
  assign n12706 = ~n12701 & ~n12705;
  assign n12707 = ~n12700 & ~n12701;
  assign n12708 = ~n12705 & n12707;
  assign n12709 = ~n12700 & n12706;
  assign n12710 = pi788 & ~n59426;
  assign n12711 = ~n6701 & ~n12670;
  assign n12712 = pi625 & n12711;
  assign n12713 = n12630 & ~n12711;
  assign n12714 = ~n12712 & ~n12713;
  assign n12715 = n12675 & ~n12714;
  assign n12716 = ~pi608 & ~n12674;
  assign n12717 = ~n12715 & n12716;
  assign n12718 = pi1153 & n12630;
  assign n12719 = ~n12712 & n12718;
  assign n12720 = pi608 & ~n12676;
  assign n12721 = ~n12719 & n12720;
  assign n12722 = ~n12717 & ~n12721;
  assign n12723 = pi778 & ~n12722;
  assign n12724 = ~pi778 & ~n12713;
  assign n12725 = ~n12723 & ~n12724;
  assign n12726 = ~pi609 & ~n12725;
  assign n12727 = pi609 & ~n12679;
  assign n12728 = ~pi1155 & ~n12727;
  assign n12729 = ~n12726 & n12728;
  assign n12730 = ~pi660 & ~n12635;
  assign n12731 = ~n12729 & n12730;
  assign n12732 = pi609 & ~n12725;
  assign n12733 = ~pi609 & ~n12679;
  assign n12734 = pi1155 & ~n12733;
  assign n12735 = ~n12732 & n12734;
  assign n12736 = pi660 & ~n12637;
  assign n12737 = ~n12735 & n12736;
  assign n12738 = ~n12731 & ~n12737;
  assign n12739 = pi785 & ~n12738;
  assign n12740 = ~pi785 & ~n12725;
  assign n12741 = ~n12739 & ~n12740;
  assign n12742 = ~pi618 & ~n12741;
  assign n12743 = pi618 & n12680;
  assign n12744 = ~pi1154 & ~n12743;
  assign n12745 = ~n12742 & n12744;
  assign n12746 = ~pi627 & ~n12643;
  assign n12747 = ~n12745 & n12746;
  assign n12748 = pi618 & ~n12741;
  assign n12749 = ~pi618 & n12680;
  assign n12750 = pi1154 & ~n12749;
  assign n12751 = ~n12748 & n12750;
  assign n12752 = pi627 & ~n12645;
  assign n12753 = ~n12751 & n12752;
  assign n12754 = ~n12747 & ~n12753;
  assign n12755 = pi781 & ~n12754;
  assign n12756 = ~pi781 & ~n12741;
  assign n12757 = ~n12755 & ~n12756;
  assign n12758 = pi619 & ~n12757;
  assign n12759 = ~pi619 & n12681;
  assign n12760 = pi1159 & ~n12759;
  assign n12761 = ~n12758 & n12760;
  assign n12762 = pi648 & ~n12653;
  assign n12763 = ~n12761 & n12762;
  assign n12764 = ~pi619 & ~n12757;
  assign n12765 = pi619 & n12681;
  assign n12766 = ~pi1159 & ~n12765;
  assign n12767 = ~n12764 & n12766;
  assign n12768 = ~pi648 & ~n12651;
  assign n12769 = ~n12767 & n12768;
  assign n12770 = pi789 & ~n12769;
  assign n12771 = pi789 & ~n12763;
  assign n12772 = ~n12769 & n12771;
  assign n12773 = ~n12763 & n12770;
  assign n12774 = ~pi789 & n12757;
  assign n12775 = n59242 & ~n12774;
  assign n12776 = ~n59427 & n12775;
  assign n12777 = ~n12710 & ~n12776;
  assign n12778 = ~n59357 & ~n12777;
  assign n12779 = n7957 & ~n59424;
  assign n12780 = n8065 & n12683;
  assign n12781 = pi629 & ~n12780;
  assign n12782 = ~n12779 & n12781;
  assign n12783 = n7958 & ~n59424;
  assign n12784 = n8074 & n12683;
  assign n12785 = ~pi629 & ~n12784;
  assign n12786 = ~n12783 & n12785;
  assign n12787 = pi792 & ~n12786;
  assign n12788 = ~n12783 & ~n12784;
  assign n12789 = ~pi629 & ~n12788;
  assign n12790 = ~n12779 & ~n12780;
  assign n12791 = pi629 & ~n12790;
  assign n12792 = ~n12789 & ~n12791;
  assign n12793 = pi792 & ~n12792;
  assign n12794 = pi792 & ~n12782;
  assign n12795 = ~n12786 & n12794;
  assign n12796 = ~n12782 & n12787;
  assign n12797 = ~n8108 & ~n59428;
  assign n12798 = ~n12778 & n12797;
  assign n12799 = ~n12696 & ~n12798;
  assign n12800 = pi644 & n12799;
  assign n12801 = ~pi787 & ~n12684;
  assign n12802 = pi1157 & ~n12687;
  assign n12803 = ~n12692 & ~n12802;
  assign n12804 = pi787 & ~n12803;
  assign n12805 = ~n12801 & ~n12804;
  assign n12806 = ~pi644 & n12805;
  assign n12807 = pi715 & ~n12806;
  assign n12808 = ~n12800 & n12807;
  assign n12809 = ~n11491 & n12628;
  assign n12810 = ~n7835 & n12663;
  assign n12811 = ~n7835 & ~n12666;
  assign n12812 = n7835 & n12628;
  assign n12813 = ~n12811 & ~n12812;
  assign n12814 = ~n12809 & ~n12810;
  assign n12815 = pi644 & ~n59429;
  assign n12816 = ~pi644 & n12628;
  assign n12817 = ~pi715 & ~n12816;
  assign n12818 = ~n12815 & n12817;
  assign n12819 = pi1160 & ~n12818;
  assign n12820 = ~n12808 & n12819;
  assign n12821 = ~pi644 & n12799;
  assign n12822 = pi644 & n12805;
  assign n12823 = ~pi715 & ~n12822;
  assign n12824 = ~n12821 & n12823;
  assign n12825 = ~pi644 & ~n59429;
  assign n12826 = pi644 & n12628;
  assign n12827 = pi715 & ~n12826;
  assign n12828 = ~n12825 & n12827;
  assign n12829 = ~pi1160 & ~n12828;
  assign n12830 = ~n12824 & n12829;
  assign n12831 = ~n12820 & ~n12830;
  assign n12832 = pi790 & ~n12831;
  assign n12833 = ~pi790 & n12799;
  assign n12834 = pi832 & ~n12833;
  assign n12835 = ~n12832 & n12834;
  assign n12836 = ~pi175 & ~n7560;
  assign n12837 = n59231 & ~n12836;
  assign n12838 = pi175 & ~n59132;
  assign n12839 = ~pi175 & n8249;
  assign n12840 = pi175 & n59251;
  assign n12841 = ~pi38 & ~n12840;
  assign n12842 = ~n12839 & n12841;
  assign n12843 = ~pi175 & ~n6863;
  assign n12844 = n7547 & ~n12843;
  assign n12845 = pi700 & ~n12844;
  assign n12846 = ~n12842 & n12845;
  assign n12847 = ~pi175 & ~pi700;
  assign n12848 = ~n7553 & n12847;
  assign n12849 = n59132 & ~n12848;
  assign n12850 = ~n12846 & n12849;
  assign n12851 = ~n12838 & ~n12850;
  assign n12852 = ~pi778 & ~n12851;
  assign n12853 = pi625 & n12851;
  assign n12854 = ~pi625 & n12836;
  assign n12855 = pi1153 & ~n12854;
  assign n12856 = ~n12853 & n12855;
  assign n12857 = ~pi625 & n12851;
  assign n12858 = pi625 & n12836;
  assign n12859 = ~pi1153 & ~n12858;
  assign n12860 = ~n12857 & n12859;
  assign n12861 = ~n12856 & ~n12860;
  assign n12862 = pi778 & ~n12861;
  assign n12863 = ~n12852 & ~n12862;
  assign n12864 = ~n59229 & n12863;
  assign n12865 = n59229 & n12836;
  assign n12866 = n59229 & ~n12836;
  assign n12867 = ~n59229 & ~n12863;
  assign n12868 = ~n12866 & ~n12867;
  assign n12869 = ~n12864 & ~n12865;
  assign n12870 = ~n59231 & ~n59430;
  assign n12871 = ~n59231 & n59430;
  assign n12872 = n59231 & n12836;
  assign n12873 = ~n12871 & ~n12872;
  assign n12874 = ~n12837 & ~n12870;
  assign n12875 = ~n7716 & ~n59431;
  assign n12876 = n7716 & n12836;
  assign n12877 = n7716 & ~n12836;
  assign n12878 = ~n7716 & n59431;
  assign n12879 = ~n12877 & ~n12878;
  assign n12880 = ~n12875 & ~n12876;
  assign n12881 = ~n7762 & n59432;
  assign n12882 = n7762 & n12836;
  assign n12883 = ~n12881 & ~n12882;
  assign n12884 = ~n59240 & ~n12883;
  assign n12885 = n59240 & n12836;
  assign n12886 = ~pi628 & ~n12883;
  assign n12887 = pi628 & n12836;
  assign n12888 = ~n12886 & ~n12887;
  assign n12889 = ~pi1156 & ~n12888;
  assign n12890 = pi628 & ~n12883;
  assign n12891 = ~pi628 & n12836;
  assign n12892 = ~n12890 & ~n12891;
  assign n12893 = pi1156 & ~n12892;
  assign n12894 = ~n12889 & ~n12893;
  assign n12895 = pi792 & ~n12894;
  assign n12896 = ~pi792 & ~n12883;
  assign n12897 = ~n12895 & ~n12896;
  assign n12898 = n59240 & ~n12836;
  assign n12899 = ~n59240 & n12883;
  assign n12900 = ~n12898 & ~n12899;
  assign n12901 = ~n12884 & ~n12885;
  assign n12902 = ~n9743 & ~n59433;
  assign n12903 = n9743 & n12836;
  assign n12904 = ~pi647 & ~n59433;
  assign n12905 = pi647 & n12836;
  assign n12906 = ~n12904 & ~n12905;
  assign n12907 = ~pi1157 & ~n12906;
  assign n12908 = pi647 & ~n59433;
  assign n12909 = ~pi647 & n12836;
  assign n12910 = ~n12908 & ~n12909;
  assign n12911 = pi1157 & ~n12910;
  assign n12912 = ~n12907 & ~n12911;
  assign n12913 = pi787 & ~n12912;
  assign n12914 = ~pi787 & ~n59433;
  assign n12915 = ~n12913 & ~n12914;
  assign n12916 = ~n12902 & ~n12903;
  assign n12917 = ~pi644 & ~n59434;
  assign n12918 = pi715 & ~n12917;
  assign n12919 = ~pi766 & n6654;
  assign n12920 = pi175 & n6853;
  assign n12921 = ~n12919 & ~n12920;
  assign n12922 = pi39 & ~n12921;
  assign n12923 = ~pi175 & pi766;
  assign n12924 = n59164 & n12923;
  assign n12925 = ~pi766 & n8180;
  assign n12926 = pi766 & ~n6799;
  assign n12927 = pi175 & ~n12926;
  assign n12928 = ~n12925 & ~n12927;
  assign n12929 = ~n12924 & n12928;
  assign n12930 = ~n12922 & n12929;
  assign n12931 = ~pi38 & ~n12930;
  assign n12932 = pi766 & n6865;
  assign n12933 = pi38 & ~n12843;
  assign n12934 = ~n12932 & n12933;
  assign n12935 = ~n12931 & ~n12934;
  assign n12936 = n59132 & ~n12935;
  assign n12937 = ~n12838 & ~n12936;
  assign n12938 = ~n7597 & ~n12937;
  assign n12939 = n7597 & ~n12836;
  assign n12940 = ~n12938 & ~n12939;
  assign n12941 = ~pi785 & ~n12940;
  assign n12942 = ~n7598 & ~n12836;
  assign n12943 = pi609 & n12938;
  assign n12944 = ~n12942 & ~n12943;
  assign n12945 = pi1155 & ~n12944;
  assign n12946 = ~n7610 & ~n12836;
  assign n12947 = ~pi609 & n12938;
  assign n12948 = ~n12946 & ~n12947;
  assign n12949 = ~pi1155 & ~n12948;
  assign n12950 = ~n12945 & ~n12949;
  assign n12951 = pi785 & ~n12950;
  assign n12952 = ~n12941 & ~n12951;
  assign n12953 = ~pi781 & ~n12952;
  assign n12954 = pi618 & n12952;
  assign n12955 = ~pi618 & n12836;
  assign n12956 = pi1154 & ~n12955;
  assign n12957 = ~n12954 & n12956;
  assign n12958 = ~pi618 & n12952;
  assign n12959 = pi618 & n12836;
  assign n12960 = ~pi1154 & ~n12959;
  assign n12961 = ~n12958 & n12960;
  assign n12962 = ~n12957 & ~n12961;
  assign n12963 = pi781 & ~n12962;
  assign n12964 = ~n12953 & ~n12963;
  assign n12965 = ~pi789 & ~n12964;
  assign n12966 = pi619 & n12964;
  assign n12967 = ~pi619 & n12836;
  assign n12968 = pi1159 & ~n12967;
  assign n12969 = ~n12966 & n12968;
  assign n12970 = ~pi619 & n12964;
  assign n12971 = pi619 & n12836;
  assign n12972 = ~pi1159 & ~n12971;
  assign n12973 = ~n12970 & n12972;
  assign n12974 = ~n12969 & ~n12973;
  assign n12975 = pi789 & ~n12974;
  assign n12976 = ~n12965 & ~n12975;
  assign n12977 = ~n8054 & n12976;
  assign n12978 = n8054 & n12836;
  assign n12979 = ~n12977 & ~n12978;
  assign n12980 = ~n7793 & ~n12979;
  assign n12981 = n7793 & n12836;
  assign n12982 = ~n12980 & ~n12981;
  assign n12983 = ~n7835 & ~n12982;
  assign n12984 = n7835 & n12836;
  assign n12985 = n7835 & ~n12836;
  assign n12986 = ~n7835 & n12982;
  assign n12987 = ~n12985 & ~n12986;
  assign n12988 = ~n12983 & ~n12984;
  assign n12989 = pi644 & n59435;
  assign n12990 = ~pi644 & n12836;
  assign n12991 = ~pi715 & ~n12990;
  assign n12992 = ~n12989 & n12991;
  assign n12993 = pi1160 & ~n12992;
  assign n12994 = ~n12918 & n12993;
  assign n12995 = pi644 & ~n59434;
  assign n12996 = ~pi715 & ~n12995;
  assign n12997 = ~pi644 & n59435;
  assign n12998 = pi644 & n12836;
  assign n12999 = pi715 & ~n12998;
  assign n13000 = ~n12997 & n12999;
  assign n13001 = ~pi1160 & ~n13000;
  assign n13002 = ~n12996 & n13001;
  assign n13003 = ~n12994 & ~n13002;
  assign n13004 = pi790 & ~n13003;
  assign n13005 = ~pi644 & n13001;
  assign n13006 = pi644 & n12993;
  assign n13007 = pi790 & ~n13006;
  assign n13008 = pi790 & ~n13005;
  assign n13009 = ~n13006 & n13008;
  assign n13010 = ~n13005 & n13007;
  assign n13011 = ~n7872 & n12982;
  assign n13012 = n7832 & ~n12909;
  assign n13013 = n7832 & n12910;
  assign n13014 = ~n12908 & n13012;
  assign n13015 = n7833 & ~n12905;
  assign n13016 = n7833 & n12906;
  assign n13017 = ~n12904 & n13015;
  assign n13018 = ~n59437 & ~n59438;
  assign n13019 = ~n13011 & ~n59438;
  assign n13020 = ~n59437 & n13019;
  assign n13021 = ~n13011 & n13018;
  assign n13022 = pi787 & ~n59439;
  assign n13023 = ~n11154 & n12979;
  assign n13024 = n7791 & ~n12887;
  assign n13025 = n7791 & n12888;
  assign n13026 = ~n12886 & n13024;
  assign n13027 = n7790 & ~n12891;
  assign n13028 = n7790 & n12892;
  assign n13029 = ~n12890 & n13027;
  assign n13030 = ~n59440 & ~n59441;
  assign n13031 = ~n13023 & n13030;
  assign n13032 = pi792 & ~n13031;
  assign n13033 = ~pi700 & n12935;
  assign n13034 = ~pi175 & n59177;
  assign n13035 = pi175 & n7111;
  assign n13036 = ~pi766 & ~n13035;
  assign n13037 = ~n13034 & n13036;
  assign n13038 = pi175 & n7188;
  assign n13039 = ~pi175 & ~n59203;
  assign n13040 = pi766 & ~n13039;
  assign n13041 = ~n13038 & n13040;
  assign n13042 = pi39 & ~n13041;
  assign n13043 = ~n13037 & n13042;
  assign n13044 = ~pi175 & n7310;
  assign n13045 = pi175 & n7333;
  assign n13046 = ~pi766 & ~n13045;
  assign n13047 = ~pi766 & ~n13044;
  assign n13048 = ~n13045 & n13047;
  assign n13049 = ~n13044 & n13046;
  assign n13050 = ~pi175 & ~n7339;
  assign n13051 = pi175 & ~n7347;
  assign n13052 = pi766 & ~n13051;
  assign n13053 = ~n13050 & n13052;
  assign n13054 = ~pi39 & ~n13053;
  assign n13055 = ~n59442 & n13054;
  assign n13056 = ~pi38 & ~n13055;
  assign n13057 = ~pi175 & n8213;
  assign n13058 = pi175 & n8217;
  assign n13059 = ~pi766 & ~n13058;
  assign n13060 = ~n13057 & n13059;
  assign n13061 = pi175 & n9808;
  assign n13062 = ~n9813 & ~n9815;
  assign n13063 = ~pi175 & ~n13062;
  assign n13064 = pi766 & ~n13063;
  assign n13065 = ~n13061 & n13064;
  assign n13066 = ~n13060 & ~n13065;
  assign n13067 = ~pi38 & ~n13066;
  assign n13068 = ~n13043 & n13056;
  assign n13069 = n6468 & ~n6873;
  assign n13070 = ~pi766 & n13069;
  assign n13071 = ~n7222 & ~n13070;
  assign n13072 = ~pi39 & ~n13071;
  assign n13073 = ~pi175 & ~n13072;
  assign n13074 = ~n7056 & ~n12629;
  assign n13075 = pi175 & ~n13074;
  assign n13076 = n59171 & n13075;
  assign n13077 = pi38 & ~n13076;
  assign n13078 = ~n13073 & n13077;
  assign n13079 = pi700 & ~n13078;
  assign n13080 = ~n59443 & n13079;
  assign n13081 = n59132 & ~n13080;
  assign n13082 = n59132 & ~n13033;
  assign n13083 = ~n13080 & n13082;
  assign n13084 = ~n13033 & n13081;
  assign n13085 = ~n12838 & ~n59444;
  assign n13086 = ~pi625 & n13085;
  assign n13087 = pi625 & n12937;
  assign n13088 = ~pi1153 & ~n13087;
  assign n13089 = ~n13086 & n13088;
  assign n13090 = ~pi608 & ~n12856;
  assign n13091 = ~n13089 & n13090;
  assign n13092 = pi625 & n13085;
  assign n13093 = ~pi625 & n12937;
  assign n13094 = pi1153 & ~n13093;
  assign n13095 = ~n13092 & n13094;
  assign n13096 = pi608 & ~n12860;
  assign n13097 = ~n13095 & n13096;
  assign n13098 = ~n13091 & ~n13097;
  assign n13099 = pi778 & ~n13098;
  assign n13100 = ~pi778 & n13085;
  assign n13101 = ~n13099 & ~n13100;
  assign n13102 = ~pi609 & ~n13101;
  assign n13103 = pi609 & n12863;
  assign n13104 = ~pi1155 & ~n13103;
  assign n13105 = ~n13102 & n13104;
  assign n13106 = ~pi660 & ~n12945;
  assign n13107 = ~n13105 & n13106;
  assign n13108 = pi609 & ~n13101;
  assign n13109 = ~pi609 & n12863;
  assign n13110 = pi1155 & ~n13109;
  assign n13111 = ~n13108 & n13110;
  assign n13112 = pi660 & ~n12949;
  assign n13113 = ~n13111 & n13112;
  assign n13114 = ~n13107 & ~n13113;
  assign n13115 = pi785 & ~n13114;
  assign n13116 = ~pi785 & ~n13101;
  assign n13117 = ~n13115 & ~n13116;
  assign n13118 = ~pi618 & ~n13117;
  assign n13119 = pi618 & n59430;
  assign n13120 = ~pi1154 & ~n13119;
  assign n13121 = ~n13118 & n13120;
  assign n13122 = ~pi627 & ~n12957;
  assign n13123 = ~n13121 & n13122;
  assign n13124 = pi618 & ~n13117;
  assign n13125 = ~pi618 & n59430;
  assign n13126 = pi1154 & ~n13125;
  assign n13127 = ~n13124 & n13126;
  assign n13128 = pi627 & ~n12961;
  assign n13129 = ~n13127 & n13128;
  assign n13130 = ~n13123 & ~n13129;
  assign n13131 = pi781 & ~n13130;
  assign n13132 = ~pi781 & ~n13117;
  assign n13133 = ~n13131 & ~n13132;
  assign n13134 = pi619 & ~n13133;
  assign n13135 = ~pi619 & ~n59431;
  assign n13136 = pi1159 & ~n13135;
  assign n13137 = ~n13134 & n13136;
  assign n13138 = pi648 & ~n12973;
  assign n13139 = ~n13137 & n13138;
  assign n13140 = ~pi619 & ~n13133;
  assign n13141 = pi619 & ~n59431;
  assign n13142 = ~pi1159 & ~n13141;
  assign n13143 = ~n13140 & n13142;
  assign n13144 = ~pi648 & ~n12969;
  assign n13145 = ~n13143 & n13144;
  assign n13146 = pi789 & ~n13145;
  assign n13147 = pi789 & ~n13139;
  assign n13148 = ~n13145 & n13147;
  assign n13149 = ~n13139 & n13146;
  assign n13150 = ~pi789 & n13133;
  assign n13151 = n59242 & ~n13150;
  assign n13152 = ~n59445 & n13151;
  assign n13153 = ~pi626 & ~n12976;
  assign n13154 = pi626 & ~n12836;
  assign n13155 = n7760 & ~n13154;
  assign n13156 = ~n13153 & n13155;
  assign n13157 = n7984 & n59432;
  assign n13158 = pi626 & ~n12976;
  assign n13159 = ~pi626 & ~n12836;
  assign n13160 = n7759 & ~n13159;
  assign n13161 = ~n13158 & n13160;
  assign n13162 = ~n13157 & ~n13161;
  assign n13163 = ~n13156 & ~n13157;
  assign n13164 = ~n13161 & n13163;
  assign n13165 = ~n13156 & n13162;
  assign n13166 = pi788 & ~n59446;
  assign n13167 = ~n59357 & ~n13166;
  assign n13168 = ~n13152 & n13167;
  assign n13169 = ~n13032 & ~n13168;
  assign n13170 = ~n8108 & ~n13169;
  assign n13171 = ~n13022 & ~n13170;
  assign n13172 = ~n59436 & n13171;
  assign n13173 = ~n13004 & ~n13172;
  assign n13174 = n58992 & ~n13173;
  assign n13175 = ~pi175 & ~n58992;
  assign n13176 = ~pi832 & ~n13175;
  assign n13177 = ~n13174 & n13176;
  assign po332 = ~n12835 & ~n13177;
  assign n13179 = ~pi176 & ~n2794;
  assign n13180 = ~pi742 & n6822;
  assign n13181 = ~n13179 & ~n13180;
  assign n13182 = ~n7875 & ~n13181;
  assign n13183 = ~pi785 & ~n13182;
  assign n13184 = ~n7880 & ~n13181;
  assign n13185 = pi1155 & ~n13184;
  assign n13186 = ~n7883 & n13182;
  assign n13187 = ~pi1155 & ~n13186;
  assign n13188 = ~n13185 & ~n13187;
  assign n13189 = pi785 & ~n13188;
  assign n13190 = ~n13183 & ~n13189;
  assign n13191 = ~pi781 & ~n13190;
  assign n13192 = ~n7890 & n13190;
  assign n13193 = pi1154 & ~n13192;
  assign n13194 = ~n7893 & n13190;
  assign n13195 = ~pi1154 & ~n13194;
  assign n13196 = ~n13193 & ~n13195;
  assign n13197 = pi781 & ~n13196;
  assign n13198 = ~n13191 & ~n13197;
  assign n13199 = ~pi789 & ~n13198;
  assign n13200 = pi619 & n13198;
  assign n13201 = ~pi619 & n13179;
  assign n13202 = pi1159 & ~n13201;
  assign n13203 = ~n13200 & n13202;
  assign n13204 = ~pi619 & n13198;
  assign n13205 = pi619 & n13179;
  assign n13206 = ~pi1159 & ~n13205;
  assign n13207 = ~n13204 & n13206;
  assign n13208 = ~n13203 & ~n13207;
  assign n13209 = pi789 & ~n13208;
  assign n13210 = ~n13199 & ~n13209;
  assign n13211 = ~n8054 & ~n13210;
  assign n13212 = n8054 & ~n13179;
  assign n13213 = ~n8054 & n13210;
  assign n13214 = n8054 & n13179;
  assign n13215 = ~n13213 & ~n13214;
  assign n13216 = ~n13211 & ~n13212;
  assign n13217 = ~n7793 & ~n59447;
  assign n13218 = n7793 & n13179;
  assign n13219 = ~n7872 & ~n13218;
  assign n13220 = ~n13217 & ~n13218;
  assign n13221 = ~n7872 & n13220;
  assign n13222 = ~n13217 & n13219;
  assign n13223 = ~pi704 & n7055;
  assign n13224 = ~n13179 & ~n13223;
  assign n13225 = ~pi778 & n13224;
  assign n13226 = ~pi625 & n13223;
  assign n13227 = ~n13224 & ~n13226;
  assign n13228 = pi1153 & ~n13227;
  assign n13229 = ~pi1153 & ~n13179;
  assign n13230 = ~n13226 & n13229;
  assign n13231 = ~n13228 & ~n13230;
  assign n13232 = pi778 & ~n13231;
  assign n13233 = ~n13225 & ~n13232;
  assign n13234 = ~n7949 & n13233;
  assign n13235 = ~n7951 & n13234;
  assign n13236 = ~n7953 & n13235;
  assign n13237 = ~n7955 & n13236;
  assign n13238 = ~n7967 & n13237;
  assign n13239 = pi647 & ~n13238;
  assign n13240 = ~pi647 & ~n13179;
  assign n13241 = ~n13239 & ~n13240;
  assign n13242 = n7832 & ~n13241;
  assign n13243 = ~pi647 & n13238;
  assign n13244 = pi647 & n13179;
  assign n13245 = ~pi1157 & ~n13244;
  assign n13246 = ~n13243 & n13245;
  assign n13247 = pi630 & n13246;
  assign n13248 = ~n13242 & ~n13247;
  assign n13249 = ~n59448 & n13248;
  assign n13250 = pi787 & ~n13249;
  assign n13251 = ~pi626 & ~n13210;
  assign n13252 = pi626 & ~n13179;
  assign n13253 = n7760 & ~n13252;
  assign n13254 = ~n13251 & n13253;
  assign n13255 = n7984 & n13236;
  assign n13256 = pi626 & ~n13210;
  assign n13257 = ~pi626 & ~n13179;
  assign n13258 = n7759 & ~n13257;
  assign n13259 = ~n13256 & n13258;
  assign n13260 = ~n13255 & ~n13259;
  assign n13261 = ~n13254 & ~n13255;
  assign n13262 = ~n13259 & n13261;
  assign n13263 = ~n13254 & n13260;
  assign n13264 = pi788 & ~n59449;
  assign n13265 = ~n6701 & ~n13224;
  assign n13266 = pi625 & n13265;
  assign n13267 = n13181 & ~n13265;
  assign n13268 = ~n13266 & ~n13267;
  assign n13269 = n13229 & ~n13268;
  assign n13270 = ~pi608 & ~n13228;
  assign n13271 = ~n13269 & n13270;
  assign n13272 = pi1153 & n13181;
  assign n13273 = ~n13266 & n13272;
  assign n13274 = pi608 & ~n13230;
  assign n13275 = ~n13273 & n13274;
  assign n13276 = ~n13271 & ~n13275;
  assign n13277 = pi778 & ~n13276;
  assign n13278 = ~pi778 & ~n13267;
  assign n13279 = ~n13277 & ~n13278;
  assign n13280 = ~pi609 & ~n13279;
  assign n13281 = pi609 & n13233;
  assign n13282 = ~pi1155 & ~n13281;
  assign n13283 = ~n13280 & n13282;
  assign n13284 = ~pi660 & ~n13185;
  assign n13285 = ~n13283 & n13284;
  assign n13286 = pi609 & ~n13279;
  assign n13287 = ~pi609 & n13233;
  assign n13288 = pi1155 & ~n13287;
  assign n13289 = ~n13286 & n13288;
  assign n13290 = pi660 & ~n13187;
  assign n13291 = ~n13289 & n13290;
  assign n13292 = ~n13285 & ~n13291;
  assign n13293 = pi785 & ~n13292;
  assign n13294 = ~pi785 & ~n13279;
  assign n13295 = ~n13293 & ~n13294;
  assign n13296 = ~pi618 & ~n13295;
  assign n13297 = pi618 & n13234;
  assign n13298 = ~pi1154 & ~n13297;
  assign n13299 = ~n13296 & n13298;
  assign n13300 = ~pi627 & ~n13193;
  assign n13301 = ~n13299 & n13300;
  assign n13302 = pi618 & ~n13295;
  assign n13303 = ~pi618 & n13234;
  assign n13304 = pi1154 & ~n13303;
  assign n13305 = ~n13302 & n13304;
  assign n13306 = pi627 & ~n13195;
  assign n13307 = ~n13305 & n13306;
  assign n13308 = ~n13301 & ~n13307;
  assign n13309 = pi781 & ~n13308;
  assign n13310 = ~pi781 & ~n13295;
  assign n13311 = ~n13309 & ~n13310;
  assign n13312 = ~pi619 & ~n13311;
  assign n13313 = pi619 & n13235;
  assign n13314 = ~pi1159 & ~n13313;
  assign n13315 = ~n13312 & n13314;
  assign n13316 = ~pi648 & ~n13203;
  assign n13317 = ~n13315 & n13316;
  assign n13318 = pi619 & ~n13311;
  assign n13319 = ~pi619 & n13235;
  assign n13320 = pi1159 & ~n13319;
  assign n13321 = ~n13318 & n13320;
  assign n13322 = pi648 & ~n13207;
  assign n13323 = ~n13321 & n13322;
  assign n13324 = pi789 & ~n13323;
  assign n13325 = pi789 & ~n13317;
  assign n13326 = ~n13323 & n13325;
  assign n13327 = ~n13317 & n13324;
  assign n13328 = ~pi789 & n13311;
  assign n13329 = n59242 & ~n13328;
  assign n13330 = ~n59450 & n13329;
  assign n13331 = ~n13264 & ~n13330;
  assign n13332 = ~n59357 & ~n13331;
  assign n13333 = n7957 & ~n59447;
  assign n13334 = n8065 & n13237;
  assign n13335 = pi629 & ~n13334;
  assign n13336 = ~n13333 & n13335;
  assign n13337 = n7958 & ~n59447;
  assign n13338 = n8074 & n13237;
  assign n13339 = ~pi629 & ~n13338;
  assign n13340 = ~n13337 & n13339;
  assign n13341 = pi792 & ~n13340;
  assign n13342 = ~n13337 & ~n13338;
  assign n13343 = ~pi629 & ~n13342;
  assign n13344 = ~n13333 & ~n13334;
  assign n13345 = pi629 & ~n13344;
  assign n13346 = ~n13343 & ~n13345;
  assign n13347 = pi792 & ~n13346;
  assign n13348 = pi792 & ~n13336;
  assign n13349 = ~n13340 & n13348;
  assign n13350 = ~n13336 & n13341;
  assign n13351 = ~n8108 & ~n59451;
  assign n13352 = ~n13332 & n13351;
  assign n13353 = ~n13250 & ~n13352;
  assign n13354 = pi644 & n13353;
  assign n13355 = ~pi787 & ~n13238;
  assign n13356 = pi1157 & ~n13241;
  assign n13357 = ~n13246 & ~n13356;
  assign n13358 = pi787 & ~n13357;
  assign n13359 = ~n13355 & ~n13358;
  assign n13360 = ~pi644 & n13359;
  assign n13361 = pi715 & ~n13360;
  assign n13362 = ~n13354 & n13361;
  assign n13363 = ~n11491 & n13179;
  assign n13364 = ~n7835 & n13217;
  assign n13365 = ~n7835 & ~n13220;
  assign n13366 = n7835 & n13179;
  assign n13367 = ~n13365 & ~n13366;
  assign n13368 = ~n13363 & ~n13364;
  assign n13369 = pi644 & ~n59452;
  assign n13370 = ~pi644 & n13179;
  assign n13371 = ~pi715 & ~n13370;
  assign n13372 = ~n13369 & n13371;
  assign n13373 = pi1160 & ~n13372;
  assign n13374 = ~n13362 & n13373;
  assign n13375 = ~pi644 & n13353;
  assign n13376 = pi644 & n13359;
  assign n13377 = ~pi715 & ~n13376;
  assign n13378 = ~n13375 & n13377;
  assign n13379 = ~pi644 & ~n59452;
  assign n13380 = pi644 & n13179;
  assign n13381 = pi715 & ~n13380;
  assign n13382 = ~n13379 & n13381;
  assign n13383 = ~pi1160 & ~n13382;
  assign n13384 = ~n13378 & n13383;
  assign n13385 = ~n13374 & ~n13384;
  assign n13386 = pi790 & ~n13385;
  assign n13387 = ~pi790 & n13353;
  assign n13388 = pi832 & ~n13387;
  assign n13389 = ~n13386 & n13388;
  assign n13390 = ~pi176 & ~n7560;
  assign n13391 = n59231 & ~n13390;
  assign n13392 = ~pi38 & ~n59251;
  assign n13393 = n59132 & ~n7547;
  assign n13394 = ~n13392 & n13393;
  assign n13395 = pi176 & ~n13394;
  assign n13396 = ~pi38 & n8249;
  assign n13397 = ~n10432 & ~n13396;
  assign n13398 = ~pi176 & n13397;
  assign n13399 = ~pi704 & ~n13398;
  assign n13400 = ~pi176 & ~n7553;
  assign n13401 = pi704 & n13400;
  assign n13402 = n59132 & ~n13401;
  assign n13403 = ~n13399 & n13402;
  assign n13404 = ~n13395 & ~n13403;
  assign n13405 = ~pi778 & ~n13404;
  assign n13406 = pi625 & n13404;
  assign n13407 = ~pi625 & n13390;
  assign n13408 = pi1153 & ~n13407;
  assign n13409 = ~n13406 & n13408;
  assign n13410 = ~pi625 & n13404;
  assign n13411 = pi625 & n13390;
  assign n13412 = ~pi1153 & ~n13411;
  assign n13413 = ~n13410 & n13412;
  assign n13414 = ~n13409 & ~n13413;
  assign n13415 = pi778 & ~n13414;
  assign n13416 = ~n13405 & ~n13415;
  assign n13417 = ~n59229 & n13416;
  assign n13418 = n59229 & n13390;
  assign n13419 = n59229 & ~n13390;
  assign n13420 = ~n59229 & ~n13416;
  assign n13421 = ~n13419 & ~n13420;
  assign n13422 = ~n13417 & ~n13418;
  assign n13423 = ~n59231 & ~n59453;
  assign n13424 = ~n59231 & n59453;
  assign n13425 = n59231 & n13390;
  assign n13426 = ~n13424 & ~n13425;
  assign n13427 = ~n13391 & ~n13423;
  assign n13428 = ~n7716 & ~n59454;
  assign n13429 = n7716 & n13390;
  assign n13430 = n7716 & ~n13390;
  assign n13431 = ~n7716 & n59454;
  assign n13432 = ~n13430 & ~n13431;
  assign n13433 = ~n13428 & ~n13429;
  assign n13434 = ~n7762 & n59455;
  assign n13435 = n7762 & n13390;
  assign n13436 = ~n13434 & ~n13435;
  assign n13437 = ~n59240 & ~n13436;
  assign n13438 = n59240 & n13390;
  assign n13439 = ~pi628 & ~n13436;
  assign n13440 = pi628 & n13390;
  assign n13441 = ~n13439 & ~n13440;
  assign n13442 = ~pi1156 & ~n13441;
  assign n13443 = pi628 & ~n13436;
  assign n13444 = ~pi628 & n13390;
  assign n13445 = ~n13443 & ~n13444;
  assign n13446 = pi1156 & ~n13445;
  assign n13447 = ~n13442 & ~n13446;
  assign n13448 = pi792 & ~n13447;
  assign n13449 = ~pi792 & ~n13436;
  assign n13450 = ~n13448 & ~n13449;
  assign n13451 = n59240 & ~n13390;
  assign n13452 = ~n59240 & n13436;
  assign n13453 = ~n13451 & ~n13452;
  assign n13454 = ~n13437 & ~n13438;
  assign n13455 = ~n9743 & ~n59456;
  assign n13456 = n9743 & n13390;
  assign n13457 = ~pi647 & ~n59456;
  assign n13458 = pi647 & n13390;
  assign n13459 = ~n13457 & ~n13458;
  assign n13460 = ~pi1157 & ~n13459;
  assign n13461 = pi647 & ~n59456;
  assign n13462 = ~pi647 & n13390;
  assign n13463 = ~n13461 & ~n13462;
  assign n13464 = pi1157 & ~n13463;
  assign n13465 = ~n13460 & ~n13464;
  assign n13466 = pi787 & ~n13465;
  assign n13467 = ~pi787 & ~n59456;
  assign n13468 = ~n13466 & ~n13467;
  assign n13469 = ~n13455 & ~n13456;
  assign n13470 = ~pi644 & ~n59457;
  assign n13471 = pi715 & ~n13470;
  assign n13472 = pi176 & ~n59132;
  assign n13473 = ~pi176 & n9787;
  assign n13474 = ~n9780 & ~n9781;
  assign n13475 = pi176 & n13474;
  assign n13476 = ~n13473 & ~n13475;
  assign n13477 = ~pi742 & ~n13476;
  assign n13478 = pi742 & ~n13400;
  assign n13479 = ~n13477 & ~n13478;
  assign n13480 = n59132 & ~n13479;
  assign n13481 = ~n13472 & ~n13480;
  assign n13482 = ~n7597 & ~n13481;
  assign n13483 = n7597 & ~n13390;
  assign n13484 = ~n13482 & ~n13483;
  assign n13485 = ~pi785 & ~n13484;
  assign n13486 = ~n7598 & ~n13390;
  assign n13487 = pi609 & n13482;
  assign n13488 = ~n13486 & ~n13487;
  assign n13489 = pi1155 & ~n13488;
  assign n13490 = ~n7610 & ~n13390;
  assign n13491 = ~pi609 & n13482;
  assign n13492 = ~n13490 & ~n13491;
  assign n13493 = ~pi1155 & ~n13492;
  assign n13494 = ~n13489 & ~n13493;
  assign n13495 = pi785 & ~n13494;
  assign n13496 = ~n13485 & ~n13495;
  assign n13497 = ~pi781 & ~n13496;
  assign n13498 = pi618 & n13496;
  assign n13499 = ~pi618 & n13390;
  assign n13500 = pi1154 & ~n13499;
  assign n13501 = ~n13498 & n13500;
  assign n13502 = ~pi618 & n13496;
  assign n13503 = pi618 & n13390;
  assign n13504 = ~pi1154 & ~n13503;
  assign n13505 = ~n13502 & n13504;
  assign n13506 = ~n13501 & ~n13505;
  assign n13507 = pi781 & ~n13506;
  assign n13508 = ~n13497 & ~n13507;
  assign n13509 = ~pi789 & ~n13508;
  assign n13510 = pi619 & n13508;
  assign n13511 = ~pi619 & n13390;
  assign n13512 = pi1159 & ~n13511;
  assign n13513 = ~n13510 & n13512;
  assign n13514 = ~pi619 & n13508;
  assign n13515 = pi619 & n13390;
  assign n13516 = ~pi1159 & ~n13515;
  assign n13517 = ~n13514 & n13516;
  assign n13518 = ~n13513 & ~n13517;
  assign n13519 = pi789 & ~n13518;
  assign n13520 = ~n13509 & ~n13519;
  assign n13521 = ~n8054 & n13520;
  assign n13522 = n8054 & n13390;
  assign n13523 = ~n13521 & ~n13522;
  assign n13524 = ~n7793 & ~n13523;
  assign n13525 = n7793 & n13390;
  assign n13526 = ~n13524 & ~n13525;
  assign n13527 = ~n7835 & ~n13526;
  assign n13528 = n7835 & n13390;
  assign n13529 = n7835 & ~n13390;
  assign n13530 = ~n7835 & n13526;
  assign n13531 = ~n13529 & ~n13530;
  assign n13532 = ~n13527 & ~n13528;
  assign n13533 = pi644 & n59458;
  assign n13534 = ~pi644 & n13390;
  assign n13535 = ~pi715 & ~n13534;
  assign n13536 = ~n13533 & n13535;
  assign n13537 = pi1160 & ~n13536;
  assign n13538 = ~n13471 & n13537;
  assign n13539 = pi644 & ~n59457;
  assign n13540 = ~pi715 & ~n13539;
  assign n13541 = ~pi644 & n59458;
  assign n13542 = pi644 & n13390;
  assign n13543 = pi715 & ~n13542;
  assign n13544 = ~n13541 & n13543;
  assign n13545 = ~pi1160 & ~n13544;
  assign n13546 = ~n13540 & n13545;
  assign n13547 = ~n13538 & ~n13546;
  assign n13548 = pi790 & ~n13547;
  assign n13549 = ~pi644 & n13545;
  assign n13550 = pi644 & n13537;
  assign n13551 = pi790 & ~n13550;
  assign n13552 = pi790 & ~n13549;
  assign n13553 = ~n13550 & n13552;
  assign n13554 = ~n13549 & n13551;
  assign n13555 = ~n7872 & n13526;
  assign n13556 = n7832 & ~n13462;
  assign n13557 = n7832 & n13463;
  assign n13558 = ~n13461 & n13556;
  assign n13559 = n7833 & ~n13458;
  assign n13560 = n7833 & n13459;
  assign n13561 = ~n13457 & n13559;
  assign n13562 = ~n59460 & ~n59461;
  assign n13563 = ~n13555 & ~n59461;
  assign n13564 = ~n59460 & n13563;
  assign n13565 = ~n13555 & n13562;
  assign n13566 = pi787 & ~n59462;
  assign n13567 = ~n11154 & n13523;
  assign n13568 = n7791 & ~n13440;
  assign n13569 = n7791 & n13441;
  assign n13570 = ~n13439 & n13568;
  assign n13571 = n7790 & ~n13444;
  assign n13572 = n7790 & n13445;
  assign n13573 = ~n13443 & n13571;
  assign n13574 = ~n59463 & ~n59464;
  assign n13575 = ~n13567 & n13574;
  assign n13576 = pi792 & ~n13575;
  assign n13577 = pi704 & n13479;
  assign n13578 = ~pi176 & n9797;
  assign n13579 = ~n9799 & ~n9801;
  assign n13580 = pi176 & ~n13579;
  assign n13581 = pi742 & ~n13580;
  assign n13582 = ~n13578 & n13581;
  assign n13583 = pi176 & n9811;
  assign n13584 = ~pi176 & ~n59320;
  assign n13585 = ~pi742 & ~n13584;
  assign n13586 = ~n13583 & n13585;
  assign n13587 = ~pi704 & ~n13586;
  assign n13588 = ~pi176 & ~n9797;
  assign n13589 = pi176 & n13579;
  assign n13590 = pi742 & ~n13589;
  assign n13591 = ~n13588 & n13590;
  assign n13592 = pi176 & ~n9811;
  assign n13593 = ~pi176 & n59320;
  assign n13594 = ~pi742 & ~n13593;
  assign n13595 = ~n13592 & n13594;
  assign n13596 = ~n13591 & ~n13595;
  assign n13597 = ~pi704 & ~n13596;
  assign n13598 = ~n13582 & n13587;
  assign n13599 = n59132 & ~n59465;
  assign n13600 = n59132 & ~n13577;
  assign n13601 = ~n59465 & n13600;
  assign n13602 = ~n13577 & n13599;
  assign n13603 = ~n13472 & ~n59466;
  assign n13604 = ~pi625 & n13603;
  assign n13605 = pi625 & n13481;
  assign n13606 = ~pi1153 & ~n13605;
  assign n13607 = ~n13604 & n13606;
  assign n13608 = ~pi608 & ~n13409;
  assign n13609 = ~n13607 & n13608;
  assign n13610 = pi625 & n13603;
  assign n13611 = ~pi625 & n13481;
  assign n13612 = pi1153 & ~n13611;
  assign n13613 = ~n13610 & n13612;
  assign n13614 = pi608 & ~n13413;
  assign n13615 = ~n13613 & n13614;
  assign n13616 = ~n13609 & ~n13615;
  assign n13617 = pi778 & ~n13616;
  assign n13618 = ~pi778 & n13603;
  assign n13619 = ~n13617 & ~n13618;
  assign n13620 = ~pi609 & ~n13619;
  assign n13621 = pi609 & n13416;
  assign n13622 = ~pi1155 & ~n13621;
  assign n13623 = ~n13620 & n13622;
  assign n13624 = ~pi660 & ~n13489;
  assign n13625 = ~n13623 & n13624;
  assign n13626 = pi609 & ~n13619;
  assign n13627 = ~pi609 & n13416;
  assign n13628 = pi1155 & ~n13627;
  assign n13629 = ~n13626 & n13628;
  assign n13630 = pi660 & ~n13493;
  assign n13631 = ~n13629 & n13630;
  assign n13632 = ~n13625 & ~n13631;
  assign n13633 = pi785 & ~n13632;
  assign n13634 = ~pi785 & ~n13619;
  assign n13635 = ~n13633 & ~n13634;
  assign n13636 = ~pi618 & ~n13635;
  assign n13637 = pi618 & n59453;
  assign n13638 = ~pi1154 & ~n13637;
  assign n13639 = ~n13636 & n13638;
  assign n13640 = ~pi627 & ~n13501;
  assign n13641 = ~n13639 & n13640;
  assign n13642 = pi618 & ~n13635;
  assign n13643 = ~pi618 & n59453;
  assign n13644 = pi1154 & ~n13643;
  assign n13645 = ~n13642 & n13644;
  assign n13646 = pi627 & ~n13505;
  assign n13647 = ~n13645 & n13646;
  assign n13648 = ~n13641 & ~n13647;
  assign n13649 = pi781 & ~n13648;
  assign n13650 = ~pi781 & ~n13635;
  assign n13651 = ~n13649 & ~n13650;
  assign n13652 = pi619 & ~n13651;
  assign n13653 = ~pi619 & ~n59454;
  assign n13654 = pi1159 & ~n13653;
  assign n13655 = ~n13652 & n13654;
  assign n13656 = pi648 & ~n13517;
  assign n13657 = ~n13655 & n13656;
  assign n13658 = ~pi619 & ~n13651;
  assign n13659 = pi619 & ~n59454;
  assign n13660 = ~pi1159 & ~n13659;
  assign n13661 = ~n13658 & n13660;
  assign n13662 = ~pi648 & ~n13513;
  assign n13663 = ~n13661 & n13662;
  assign n13664 = pi789 & ~n13663;
  assign n13665 = pi789 & ~n13657;
  assign n13666 = ~n13663 & n13665;
  assign n13667 = ~n13657 & n13664;
  assign n13668 = ~pi789 & n13651;
  assign n13669 = n59242 & ~n13668;
  assign n13670 = ~n59467 & n13669;
  assign n13671 = ~pi626 & ~n13520;
  assign n13672 = pi626 & ~n13390;
  assign n13673 = n7760 & ~n13672;
  assign n13674 = ~n13671 & n13673;
  assign n13675 = n7984 & n59455;
  assign n13676 = pi626 & ~n13520;
  assign n13677 = ~pi626 & ~n13390;
  assign n13678 = n7759 & ~n13677;
  assign n13679 = ~n13676 & n13678;
  assign n13680 = ~n13675 & ~n13679;
  assign n13681 = ~n13674 & ~n13675;
  assign n13682 = ~n13679 & n13681;
  assign n13683 = ~n13674 & n13680;
  assign n13684 = pi788 & ~n59468;
  assign n13685 = ~n59357 & ~n13684;
  assign n13686 = ~n13670 & n13685;
  assign n13687 = ~n13576 & ~n13686;
  assign n13688 = ~n13670 & ~n13684;
  assign n13689 = ~n13576 & ~n13688;
  assign n13690 = n59357 & n13575;
  assign n13691 = ~n8108 & ~n13690;
  assign n13692 = ~n13689 & n13691;
  assign n13693 = ~n8108 & ~n13687;
  assign n13694 = ~n13566 & ~n59469;
  assign n13695 = ~n59459 & n13694;
  assign n13696 = ~n13548 & ~n13695;
  assign n13697 = n58992 & ~n13696;
  assign n13698 = ~pi176 & ~n58992;
  assign n13699 = ~pi832 & ~n13698;
  assign n13700 = ~n13697 & n13699;
  assign po333 = ~n13389 & ~n13700;
  assign n13702 = ~pi177 & ~n2794;
  assign n13703 = ~pi757 & n6822;
  assign n13704 = ~n13702 & ~n13703;
  assign n13705 = ~n7875 & ~n13704;
  assign n13706 = ~pi785 & ~n13705;
  assign n13707 = ~n7880 & ~n13704;
  assign n13708 = pi1155 & ~n13707;
  assign n13709 = ~n7883 & n13705;
  assign n13710 = ~pi1155 & ~n13709;
  assign n13711 = ~n13708 & ~n13710;
  assign n13712 = pi785 & ~n13711;
  assign n13713 = ~n13706 & ~n13712;
  assign n13714 = ~pi781 & ~n13713;
  assign n13715 = ~n7890 & n13713;
  assign n13716 = pi1154 & ~n13715;
  assign n13717 = ~n7893 & n13713;
  assign n13718 = ~pi1154 & ~n13717;
  assign n13719 = ~n13716 & ~n13718;
  assign n13720 = pi781 & ~n13719;
  assign n13721 = ~n13714 & ~n13720;
  assign n13722 = ~pi789 & ~n13721;
  assign n13723 = pi619 & n13721;
  assign n13724 = ~pi619 & n13702;
  assign n13725 = pi1159 & ~n13724;
  assign n13726 = ~n13723 & n13725;
  assign n13727 = ~pi619 & n13721;
  assign n13728 = pi619 & n13702;
  assign n13729 = ~pi1159 & ~n13728;
  assign n13730 = ~n13727 & n13729;
  assign n13731 = ~n13726 & ~n13730;
  assign n13732 = pi789 & ~n13731;
  assign n13733 = ~n13722 & ~n13732;
  assign n13734 = ~n8054 & ~n13733;
  assign n13735 = n8054 & ~n13702;
  assign n13736 = ~n8054 & n13733;
  assign n13737 = n8054 & n13702;
  assign n13738 = ~n13736 & ~n13737;
  assign n13739 = ~n13734 & ~n13735;
  assign n13740 = ~n7793 & ~n59470;
  assign n13741 = n7793 & n13702;
  assign n13742 = ~n7872 & ~n13741;
  assign n13743 = ~n13740 & ~n13741;
  assign n13744 = ~n7872 & n13743;
  assign n13745 = ~n13740 & n13742;
  assign n13746 = ~pi686 & n7055;
  assign n13747 = ~n13702 & ~n13746;
  assign n13748 = ~pi778 & n13747;
  assign n13749 = ~pi625 & n13746;
  assign n13750 = ~n13747 & ~n13749;
  assign n13751 = pi1153 & ~n13750;
  assign n13752 = ~pi1153 & ~n13702;
  assign n13753 = ~n13749 & n13752;
  assign n13754 = ~n13751 & ~n13753;
  assign n13755 = pi778 & ~n13754;
  assign n13756 = ~n13748 & ~n13755;
  assign n13757 = ~n7949 & n13756;
  assign n13758 = ~n7951 & n13757;
  assign n13759 = ~n7953 & n13758;
  assign n13760 = ~n7955 & n13759;
  assign n13761 = ~n7967 & n13760;
  assign n13762 = pi647 & ~n13761;
  assign n13763 = ~pi647 & ~n13702;
  assign n13764 = ~n13762 & ~n13763;
  assign n13765 = n7832 & ~n13764;
  assign n13766 = ~pi647 & n13761;
  assign n13767 = pi647 & n13702;
  assign n13768 = ~pi1157 & ~n13767;
  assign n13769 = ~n13766 & n13768;
  assign n13770 = pi630 & n13769;
  assign n13771 = ~n13765 & ~n13770;
  assign n13772 = ~n59471 & n13771;
  assign n13773 = pi787 & ~n13772;
  assign n13774 = ~pi626 & ~n13733;
  assign n13775 = pi626 & ~n13702;
  assign n13776 = n7760 & ~n13775;
  assign n13777 = ~n13774 & n13776;
  assign n13778 = n7984 & n13759;
  assign n13779 = pi626 & ~n13733;
  assign n13780 = ~pi626 & ~n13702;
  assign n13781 = n7759 & ~n13780;
  assign n13782 = ~n13779 & n13781;
  assign n13783 = ~n13778 & ~n13782;
  assign n13784 = ~n13777 & ~n13778;
  assign n13785 = ~n13782 & n13784;
  assign n13786 = ~n13777 & n13783;
  assign n13787 = pi788 & ~n59472;
  assign n13788 = ~n6701 & ~n13747;
  assign n13789 = pi625 & n13788;
  assign n13790 = n13704 & ~n13788;
  assign n13791 = ~n13789 & ~n13790;
  assign n13792 = n13752 & ~n13791;
  assign n13793 = ~pi608 & ~n13751;
  assign n13794 = ~n13792 & n13793;
  assign n13795 = pi1153 & n13704;
  assign n13796 = ~n13789 & n13795;
  assign n13797 = pi608 & ~n13753;
  assign n13798 = ~n13796 & n13797;
  assign n13799 = ~n13794 & ~n13798;
  assign n13800 = pi778 & ~n13799;
  assign n13801 = ~pi778 & ~n13790;
  assign n13802 = ~n13800 & ~n13801;
  assign n13803 = ~pi609 & ~n13802;
  assign n13804 = pi609 & n13756;
  assign n13805 = ~pi1155 & ~n13804;
  assign n13806 = ~n13803 & n13805;
  assign n13807 = ~pi660 & ~n13708;
  assign n13808 = ~n13806 & n13807;
  assign n13809 = pi609 & ~n13802;
  assign n13810 = ~pi609 & n13756;
  assign n13811 = pi1155 & ~n13810;
  assign n13812 = ~n13809 & n13811;
  assign n13813 = pi660 & ~n13710;
  assign n13814 = ~n13812 & n13813;
  assign n13815 = ~n13808 & ~n13814;
  assign n13816 = pi785 & ~n13815;
  assign n13817 = ~pi785 & ~n13802;
  assign n13818 = ~n13816 & ~n13817;
  assign n13819 = ~pi618 & ~n13818;
  assign n13820 = pi618 & n13757;
  assign n13821 = ~pi1154 & ~n13820;
  assign n13822 = ~n13819 & n13821;
  assign n13823 = ~pi627 & ~n13716;
  assign n13824 = ~n13822 & n13823;
  assign n13825 = pi618 & ~n13818;
  assign n13826 = ~pi618 & n13757;
  assign n13827 = pi1154 & ~n13826;
  assign n13828 = ~n13825 & n13827;
  assign n13829 = pi627 & ~n13718;
  assign n13830 = ~n13828 & n13829;
  assign n13831 = ~n13824 & ~n13830;
  assign n13832 = pi781 & ~n13831;
  assign n13833 = ~pi781 & ~n13818;
  assign n13834 = ~n13832 & ~n13833;
  assign n13835 = ~pi619 & ~n13834;
  assign n13836 = pi619 & n13758;
  assign n13837 = ~pi1159 & ~n13836;
  assign n13838 = ~n13835 & n13837;
  assign n13839 = ~pi648 & ~n13726;
  assign n13840 = ~n13838 & n13839;
  assign n13841 = pi619 & ~n13834;
  assign n13842 = ~pi619 & n13758;
  assign n13843 = pi1159 & ~n13842;
  assign n13844 = ~n13841 & n13843;
  assign n13845 = pi648 & ~n13730;
  assign n13846 = ~n13844 & n13845;
  assign n13847 = pi789 & ~n13846;
  assign n13848 = pi789 & ~n13840;
  assign n13849 = ~n13846 & n13848;
  assign n13850 = ~n13840 & n13847;
  assign n13851 = ~pi789 & n13834;
  assign n13852 = n59242 & ~n13851;
  assign n13853 = ~n59473 & n13852;
  assign n13854 = ~n13787 & ~n13853;
  assign n13855 = ~n59357 & ~n13854;
  assign n13856 = n7957 & ~n59470;
  assign n13857 = n8065 & n13760;
  assign n13858 = pi629 & ~n13857;
  assign n13859 = ~n13856 & n13858;
  assign n13860 = n7958 & ~n59470;
  assign n13861 = n8074 & n13760;
  assign n13862 = ~pi629 & ~n13861;
  assign n13863 = ~n13860 & n13862;
  assign n13864 = pi792 & ~n13863;
  assign n13865 = ~n13860 & ~n13861;
  assign n13866 = ~pi629 & ~n13865;
  assign n13867 = ~n13856 & ~n13857;
  assign n13868 = pi629 & ~n13867;
  assign n13869 = ~n13866 & ~n13868;
  assign n13870 = pi792 & ~n13869;
  assign n13871 = pi792 & ~n13859;
  assign n13872 = ~n13863 & n13871;
  assign n13873 = ~n13859 & n13864;
  assign n13874 = ~n8108 & ~n59474;
  assign n13875 = ~n13855 & n13874;
  assign n13876 = ~n13773 & ~n13875;
  assign n13877 = pi644 & n13876;
  assign n13878 = ~pi787 & ~n13761;
  assign n13879 = pi1157 & ~n13764;
  assign n13880 = ~n13769 & ~n13879;
  assign n13881 = pi787 & ~n13880;
  assign n13882 = ~n13878 & ~n13881;
  assign n13883 = ~pi644 & n13882;
  assign n13884 = pi715 & ~n13883;
  assign n13885 = ~n13877 & n13884;
  assign n13886 = ~n11491 & n13702;
  assign n13887 = ~n7835 & n13740;
  assign n13888 = ~n7835 & ~n13743;
  assign n13889 = n7835 & n13702;
  assign n13890 = ~n13888 & ~n13889;
  assign n13891 = ~n13886 & ~n13887;
  assign n13892 = pi644 & ~n59475;
  assign n13893 = ~pi644 & n13702;
  assign n13894 = ~pi715 & ~n13893;
  assign n13895 = ~n13892 & n13894;
  assign n13896 = pi1160 & ~n13895;
  assign n13897 = ~n13885 & n13896;
  assign n13898 = ~pi644 & n13876;
  assign n13899 = pi644 & n13882;
  assign n13900 = ~pi715 & ~n13899;
  assign n13901 = ~n13898 & n13900;
  assign n13902 = ~pi644 & ~n59475;
  assign n13903 = pi644 & n13702;
  assign n13904 = pi715 & ~n13903;
  assign n13905 = ~n13902 & n13904;
  assign n13906 = ~pi1160 & ~n13905;
  assign n13907 = ~n13901 & n13906;
  assign n13908 = ~n13897 & ~n13907;
  assign n13909 = pi790 & ~n13908;
  assign n13910 = ~pi790 & n13876;
  assign n13911 = pi832 & ~n13910;
  assign n13912 = ~n13909 & n13911;
  assign n13913 = pi177 & ~n59132;
  assign n13914 = pi757 & ~n7553;
  assign n13915 = ~pi757 & ~n9787;
  assign n13916 = ~n13914 & ~n13915;
  assign n13917 = ~pi177 & ~n13916;
  assign n13918 = ~pi177 & ~n9780;
  assign n13919 = ~pi757 & ~n13918;
  assign n13920 = ~n13474 & n13919;
  assign n13921 = ~n13917 & ~n13920;
  assign n13922 = n59132 & n13921;
  assign n13923 = ~n13913 & ~n13922;
  assign n13924 = ~n7597 & ~n13923;
  assign n13925 = ~pi177 & ~n7560;
  assign n13926 = n7597 & ~n13925;
  assign n13927 = ~n13924 & ~n13926;
  assign n13928 = ~pi785 & ~n13927;
  assign n13929 = ~n7598 & ~n13925;
  assign n13930 = pi609 & n13924;
  assign n13931 = ~n13929 & ~n13930;
  assign n13932 = pi1155 & ~n13931;
  assign n13933 = ~n7610 & ~n13925;
  assign n13934 = ~pi609 & n13924;
  assign n13935 = ~n13933 & ~n13934;
  assign n13936 = ~pi1155 & ~n13935;
  assign n13937 = ~n13932 & ~n13936;
  assign n13938 = pi785 & ~n13937;
  assign n13939 = ~n13928 & ~n13938;
  assign n13940 = ~pi781 & ~n13939;
  assign n13941 = pi618 & n13939;
  assign n13942 = ~pi618 & n13925;
  assign n13943 = pi1154 & ~n13942;
  assign n13944 = ~n13941 & n13943;
  assign n13945 = ~pi618 & n13939;
  assign n13946 = pi618 & n13925;
  assign n13947 = ~pi1154 & ~n13946;
  assign n13948 = ~n13945 & n13947;
  assign n13949 = ~n13944 & ~n13948;
  assign n13950 = pi781 & ~n13949;
  assign n13951 = ~n13940 & ~n13950;
  assign n13952 = ~pi789 & ~n13951;
  assign n13953 = ~pi619 & n13951;
  assign n13954 = pi619 & n13925;
  assign n13955 = ~pi1159 & ~n13954;
  assign n13956 = ~n13953 & n13955;
  assign n13957 = pi619 & n13951;
  assign n13958 = ~pi619 & n13925;
  assign n13959 = pi1159 & ~n13958;
  assign n13960 = ~n13957 & n13959;
  assign n13961 = ~n13956 & ~n13960;
  assign n13962 = pi789 & ~n13961;
  assign n13963 = ~n13952 & ~n13962;
  assign n13964 = ~n8054 & n13963;
  assign n13965 = n8054 & n13925;
  assign n13966 = ~n13964 & ~n13965;
  assign n13967 = ~n11154 & n13966;
  assign n13968 = n7762 & ~n13925;
  assign n13969 = n59231 & ~n13925;
  assign n13970 = ~pi177 & n8249;
  assign n13971 = pi177 & n59251;
  assign n13972 = ~pi38 & ~n13971;
  assign n13973 = ~n13970 & n13972;
  assign n13974 = ~pi177 & ~n6863;
  assign n13975 = n7547 & ~n13974;
  assign n13976 = ~pi686 & ~n13975;
  assign n13977 = ~n13973 & n13976;
  assign n13978 = ~pi177 & pi686;
  assign n13979 = ~n7553 & n13978;
  assign n13980 = n59132 & ~n13979;
  assign n13981 = ~n13977 & n13980;
  assign n13982 = ~n13913 & ~n13981;
  assign n13983 = ~pi778 & ~n13982;
  assign n13984 = pi625 & n13982;
  assign n13985 = ~pi625 & n13925;
  assign n13986 = pi1153 & ~n13985;
  assign n13987 = ~n13984 & n13986;
  assign n13988 = ~pi625 & n13982;
  assign n13989 = pi625 & n13925;
  assign n13990 = ~pi1153 & ~n13989;
  assign n13991 = ~n13988 & n13990;
  assign n13992 = ~n13987 & ~n13991;
  assign n13993 = pi778 & ~n13992;
  assign n13994 = ~n13983 & ~n13993;
  assign n13995 = ~n59229 & n13994;
  assign n13996 = n59229 & n13925;
  assign n13997 = n59229 & ~n13925;
  assign n13998 = ~n59229 & ~n13994;
  assign n13999 = ~n13997 & ~n13998;
  assign n14000 = ~n13995 & ~n13996;
  assign n14001 = ~n59231 & ~n59476;
  assign n14002 = ~n59231 & n59476;
  assign n14003 = n59231 & n13925;
  assign n14004 = ~n14002 & ~n14003;
  assign n14005 = ~n13969 & ~n14001;
  assign n14006 = ~n7716 & ~n59477;
  assign n14007 = n7716 & n13925;
  assign n14008 = n7716 & ~n13925;
  assign n14009 = ~n7716 & n59477;
  assign n14010 = ~n14008 & ~n14009;
  assign n14011 = ~n14006 & ~n14007;
  assign n14012 = ~n7762 & ~n59478;
  assign n14013 = ~n7762 & n59478;
  assign n14014 = n7762 & n13925;
  assign n14015 = ~n14013 & ~n14014;
  assign n14016 = ~n13968 & ~n14012;
  assign n14017 = ~pi628 & ~n59479;
  assign n14018 = pi628 & n13925;
  assign n14019 = ~pi1156 & ~n14018;
  assign n14020 = ~n14017 & n14019;
  assign n14021 = pi629 & n14020;
  assign n14022 = ~pi628 & ~n13925;
  assign n14023 = pi628 & n59479;
  assign n14024 = ~n14022 & ~n14023;
  assign n14025 = n7790 & ~n14024;
  assign n14026 = ~n14021 & ~n14025;
  assign n14027 = ~n13967 & n14026;
  assign n14028 = pi792 & ~n14027;
  assign n14029 = pi619 & ~n59477;
  assign n14030 = ~pi1159 & ~n14029;
  assign n14031 = ~pi648 & ~n13960;
  assign n14032 = ~n14030 & n14031;
  assign n14033 = ~pi619 & ~n59477;
  assign n14034 = pi1159 & ~n14033;
  assign n14035 = pi648 & ~n13956;
  assign n14036 = ~n14034 & n14035;
  assign n14037 = ~n14032 & ~n14036;
  assign n14038 = pi789 & ~n14037;
  assign n14039 = pi686 & ~n13921;
  assign n14040 = ~pi177 & n8213;
  assign n14041 = pi177 & n8217;
  assign n14042 = ~pi38 & ~n14041;
  assign n14043 = ~n14040 & n14042;
  assign n14044 = n8233 & ~n13974;
  assign n14045 = pi757 & ~n14044;
  assign n14046 = ~n14043 & n14045;
  assign n14047 = pi177 & n9808;
  assign n14048 = ~pi177 & ~n13062;
  assign n14049 = ~pi38 & ~n14048;
  assign n14050 = ~n14047 & n14049;
  assign n14051 = ~pi177 & ~n59319;
  assign n14052 = pi177 & n59207;
  assign n14053 = pi38 & ~n14052;
  assign n14054 = ~n14051 & n14053;
  assign n14055 = n9810 & ~n13974;
  assign n14056 = ~pi757 & ~n59480;
  assign n14057 = ~n14050 & n14056;
  assign n14058 = ~n14046 & ~n14057;
  assign n14059 = ~pi686 & ~n14058;
  assign n14060 = n59132 & ~n14059;
  assign n14061 = ~n14039 & n14060;
  assign n14062 = ~n13913 & ~n14061;
  assign n14063 = ~pi625 & n14062;
  assign n14064 = pi625 & n13923;
  assign n14065 = ~pi1153 & ~n14064;
  assign n14066 = ~n14063 & n14065;
  assign n14067 = ~pi608 & ~n13987;
  assign n14068 = ~n14066 & n14067;
  assign n14069 = pi625 & n14062;
  assign n14070 = ~pi625 & n13923;
  assign n14071 = pi1153 & ~n14070;
  assign n14072 = ~n14069 & n14071;
  assign n14073 = pi608 & ~n13991;
  assign n14074 = ~n14072 & n14073;
  assign n14075 = ~n14068 & ~n14074;
  assign n14076 = pi778 & ~n14075;
  assign n14077 = ~pi778 & n14062;
  assign n14078 = ~pi778 & ~n14062;
  assign n14079 = pi778 & ~n14074;
  assign n14080 = ~n14068 & n14079;
  assign n14081 = ~n14078 & ~n14080;
  assign n14082 = ~n14076 & ~n14077;
  assign n14083 = ~pi609 & n59481;
  assign n14084 = pi609 & n13994;
  assign n14085 = ~pi1155 & ~n14084;
  assign n14086 = ~n14083 & n14085;
  assign n14087 = ~pi660 & ~n13932;
  assign n14088 = ~n14086 & n14087;
  assign n14089 = pi609 & n59481;
  assign n14090 = ~pi609 & n13994;
  assign n14091 = pi1155 & ~n14090;
  assign n14092 = ~n14089 & n14091;
  assign n14093 = pi660 & ~n13936;
  assign n14094 = ~n14092 & n14093;
  assign n14095 = ~n14088 & ~n14094;
  assign n14096 = pi785 & ~n14095;
  assign n14097 = ~pi785 & n59481;
  assign n14098 = ~n14096 & ~n14097;
  assign n14099 = pi618 & ~n14098;
  assign n14100 = ~pi618 & n59476;
  assign n14101 = pi1154 & ~n14100;
  assign n14102 = ~n14099 & n14101;
  assign n14103 = pi627 & ~n13948;
  assign n14104 = ~n14102 & n14103;
  assign n14105 = ~pi618 & ~n14098;
  assign n14106 = pi618 & n59476;
  assign n14107 = ~pi1154 & ~n14106;
  assign n14108 = ~n14105 & n14107;
  assign n14109 = ~pi627 & ~n13944;
  assign n14110 = ~n14108 & n14109;
  assign n14111 = pi781 & ~n14110;
  assign n14112 = ~n14104 & n14111;
  assign n14113 = ~pi619 & n14031;
  assign n14114 = pi619 & n14035;
  assign n14115 = pi789 & ~n14114;
  assign n14116 = ~n14113 & n14115;
  assign n14117 = ~pi781 & n14098;
  assign n14118 = ~n14116 & ~n14117;
  assign n14119 = ~n14112 & n14118;
  assign n14120 = ~n14104 & ~n14110;
  assign n14121 = pi781 & ~n14120;
  assign n14122 = ~pi781 & ~n14098;
  assign n14123 = ~n14121 & ~n14122;
  assign n14124 = ~pi619 & ~n14123;
  assign n14125 = n14030 & ~n14124;
  assign n14126 = n14031 & ~n14125;
  assign n14127 = pi619 & ~n14123;
  assign n14128 = n14034 & ~n14127;
  assign n14129 = n14035 & ~n14128;
  assign n14130 = ~n14126 & ~n14129;
  assign n14131 = pi789 & ~n14130;
  assign n14132 = ~pi789 & ~n14123;
  assign n14133 = ~n14131 & ~n14132;
  assign n14134 = ~n14038 & ~n14119;
  assign n14135 = n59242 & ~n59482;
  assign n14136 = n12139 & n13963;
  assign n14137 = ~pi641 & ~n59478;
  assign n14138 = pi641 & ~n13925;
  assign n14139 = n7912 & ~n14138;
  assign n14140 = ~n14137 & n14139;
  assign n14141 = pi641 & ~n59478;
  assign n14142 = ~pi641 & ~n13925;
  assign n14143 = n7911 & ~n14142;
  assign n14144 = ~n14141 & n14143;
  assign n14145 = ~n14140 & ~n14144;
  assign n14146 = ~n14136 & n14145;
  assign n14147 = pi788 & ~n14146;
  assign n14148 = ~n59357 & ~n14147;
  assign n14149 = ~n14135 & n14148;
  assign n14150 = ~pi788 & n59482;
  assign n14151 = ~pi626 & n59482;
  assign n14152 = pi626 & ~n59478;
  assign n14153 = ~pi641 & ~n14152;
  assign n14154 = ~n14151 & n14153;
  assign n14155 = ~pi626 & ~n13963;
  assign n14156 = pi626 & ~n13925;
  assign n14157 = pi641 & ~n14156;
  assign n14158 = ~n14155 & n14157;
  assign n14159 = ~pi1158 & ~n14158;
  assign n14160 = ~n14154 & n14159;
  assign n14161 = pi626 & n59482;
  assign n14162 = ~pi626 & ~n59478;
  assign n14163 = pi641 & ~n14162;
  assign n14164 = ~n14161 & n14163;
  assign n14165 = pi626 & ~n13963;
  assign n14166 = ~pi626 & ~n13925;
  assign n14167 = ~pi641 & ~n14166;
  assign n14168 = ~n14165 & n14167;
  assign n14169 = pi1158 & ~n14168;
  assign n14170 = ~n14164 & n14169;
  assign n14171 = ~n14160 & ~n14170;
  assign n14172 = pi788 & ~n14171;
  assign n14173 = ~n14150 & ~n14172;
  assign n14174 = ~pi628 & n14173;
  assign n14175 = pi628 & ~n13966;
  assign n14176 = ~pi1156 & ~n14175;
  assign n14177 = ~n14174 & n14176;
  assign n14178 = pi628 & ~n59479;
  assign n14179 = ~pi628 & n13925;
  assign n14180 = pi1156 & ~n14179;
  assign n14181 = pi1156 & ~n14024;
  assign n14182 = ~n14178 & n14180;
  assign n14183 = ~pi629 & ~n59483;
  assign n14184 = ~n14177 & n14183;
  assign n14185 = pi628 & n14173;
  assign n14186 = ~pi628 & ~n13966;
  assign n14187 = pi1156 & ~n14186;
  assign n14188 = ~n14185 & n14187;
  assign n14189 = pi629 & ~n14020;
  assign n14190 = ~n14188 & n14189;
  assign n14191 = ~n14184 & ~n14190;
  assign n14192 = pi792 & ~n14191;
  assign n14193 = ~pi792 & n14173;
  assign n14194 = ~n14192 & ~n14193;
  assign n14195 = ~n14028 & ~n14149;
  assign n14196 = n59244 & n59484;
  assign n14197 = ~n7793 & ~n13966;
  assign n14198 = n7793 & n13925;
  assign n14199 = ~n14197 & ~n14198;
  assign n14200 = ~n7872 & n14199;
  assign n14201 = ~pi792 & n59479;
  assign n14202 = ~n14020 & ~n59483;
  assign n14203 = pi792 & ~n14202;
  assign n14204 = ~n14201 & ~n14203;
  assign n14205 = ~pi647 & n14204;
  assign n14206 = pi647 & n13925;
  assign n14207 = ~pi1157 & ~n14206;
  assign n14208 = ~n14205 & n14207;
  assign n14209 = pi630 & n14208;
  assign n14210 = ~pi647 & ~n13925;
  assign n14211 = pi647 & ~n14204;
  assign n14212 = ~n14210 & ~n14211;
  assign n14213 = n7832 & ~n14212;
  assign n14214 = ~n14209 & ~n14213;
  assign n14215 = ~n14200 & n14214;
  assign n14216 = ~pi647 & ~n59484;
  assign n14217 = pi647 & ~n14199;
  assign n14218 = ~pi1157 & ~n14217;
  assign n14219 = ~n14216 & n14218;
  assign n14220 = pi647 & n14204;
  assign n14221 = ~pi647 & n13925;
  assign n14222 = pi1157 & ~n14221;
  assign n14223 = pi1157 & ~n14212;
  assign n14224 = ~n14220 & n14222;
  assign n14225 = ~pi630 & ~n59485;
  assign n14226 = ~n14219 & n14225;
  assign n14227 = pi647 & ~n59484;
  assign n14228 = ~pi647 & ~n14199;
  assign n14229 = pi1157 & ~n14228;
  assign n14230 = ~n14227 & n14229;
  assign n14231 = pi630 & ~n14208;
  assign n14232 = ~n14230 & n14231;
  assign n14233 = ~n14226 & ~n14232;
  assign n14234 = ~n14196 & n14215;
  assign n14235 = pi787 & n59486;
  assign n14236 = ~pi787 & n59484;
  assign n14237 = pi787 & ~n59486;
  assign n14238 = ~pi787 & ~n59484;
  assign n14239 = ~n14237 & ~n14238;
  assign n14240 = ~n14235 & ~n14236;
  assign n14241 = pi644 & ~n59487;
  assign n14242 = ~pi787 & ~n14204;
  assign n14243 = ~n14208 & ~n59485;
  assign n14244 = pi787 & ~n14243;
  assign n14245 = ~n14242 & ~n14244;
  assign n14246 = ~pi644 & n14245;
  assign n14247 = pi715 & ~n14246;
  assign n14248 = ~n14241 & n14247;
  assign n14249 = ~n7835 & ~n14199;
  assign n14250 = n7835 & n13925;
  assign n14251 = n7835 & ~n13925;
  assign n14252 = ~n7835 & n14199;
  assign n14253 = ~n14251 & ~n14252;
  assign n14254 = ~n14249 & ~n14250;
  assign n14255 = pi644 & n59488;
  assign n14256 = ~pi644 & n13925;
  assign n14257 = ~pi715 & ~n14256;
  assign n14258 = ~n14255 & n14257;
  assign n14259 = pi1160 & ~n14258;
  assign n14260 = ~n14248 & n14259;
  assign n14261 = ~pi644 & n59488;
  assign n14262 = pi644 & n13925;
  assign n14263 = pi715 & ~n14262;
  assign n14264 = ~n14261 & n14263;
  assign n14265 = ~pi1160 & ~n14264;
  assign n14266 = pi644 & n14245;
  assign n14267 = ~pi715 & ~n14266;
  assign n14268 = ~pi644 & ~n59487;
  assign n14269 = n14267 & ~n14268;
  assign n14270 = n14265 & ~n14269;
  assign n14271 = pi790 & ~n14270;
  assign n14272 = pi790 & ~n14260;
  assign n14273 = ~n14270 & n14272;
  assign n14274 = ~n14260 & n14271;
  assign n14275 = ~pi790 & n59487;
  assign n14276 = n58992 & ~n14275;
  assign n14277 = n14265 & ~n14267;
  assign n14278 = ~n14260 & ~n14277;
  assign n14279 = pi790 & ~n14278;
  assign n14280 = ~pi644 & n14265;
  assign n14281 = pi790 & ~n14280;
  assign n14282 = ~n59487 & ~n14281;
  assign n14283 = ~n14279 & ~n14282;
  assign n14284 = n58992 & ~n14283;
  assign n14285 = ~n59489 & n14276;
  assign n14286 = ~pi177 & ~n58992;
  assign n14287 = ~pi832 & ~n14286;
  assign n14288 = ~n59490 & n14287;
  assign po334 = ~n13912 & ~n14288;
  assign n14290 = ~pi178 & ~n2794;
  assign n14291 = ~pi760 & n6822;
  assign n14292 = ~n14290 & ~n14291;
  assign n14293 = ~n7875 & ~n14292;
  assign n14294 = ~pi785 & ~n14293;
  assign n14295 = n7610 & n14291;
  assign n14296 = n14293 & ~n14295;
  assign n14297 = pi1155 & ~n14296;
  assign n14298 = ~pi1155 & ~n14290;
  assign n14299 = ~n14295 & n14298;
  assign n14300 = ~n14297 & ~n14299;
  assign n14301 = pi785 & ~n14300;
  assign n14302 = ~n14294 & ~n14301;
  assign n14303 = ~pi781 & ~n14302;
  assign n14304 = ~n7890 & n14302;
  assign n14305 = pi1154 & ~n14304;
  assign n14306 = ~n7893 & n14302;
  assign n14307 = ~pi1154 & ~n14306;
  assign n14308 = ~n14305 & ~n14307;
  assign n14309 = pi781 & ~n14308;
  assign n14310 = ~n14303 & ~n14309;
  assign n14311 = ~pi789 & ~n14310;
  assign n14312 = ~n11882 & n14310;
  assign n14313 = pi1159 & ~n14312;
  assign n14314 = ~n11885 & n14310;
  assign n14315 = ~pi1159 & ~n14314;
  assign n14316 = ~n14313 & ~n14315;
  assign n14317 = pi789 & ~n14316;
  assign n14318 = ~n14311 & ~n14317;
  assign n14319 = ~n8054 & ~n14318;
  assign n14320 = n8054 & ~n14290;
  assign n14321 = ~n8054 & n14318;
  assign n14322 = n8054 & n14290;
  assign n14323 = ~n14321 & ~n14322;
  assign n14324 = ~n14319 & ~n14320;
  assign n14325 = ~n7793 & ~n59491;
  assign n14326 = n7793 & n14290;
  assign n14327 = ~n7872 & ~n14326;
  assign n14328 = ~n14325 & ~n14326;
  assign n14329 = ~n7872 & n14328;
  assign n14330 = ~n14325 & n14327;
  assign n14331 = ~pi688 & n7055;
  assign n14332 = ~n14290 & ~n14331;
  assign n14333 = ~pi778 & ~n14332;
  assign n14334 = ~pi625 & n14331;
  assign n14335 = ~n14332 & ~n14334;
  assign n14336 = pi1153 & ~n14335;
  assign n14337 = ~pi1153 & ~n14290;
  assign n14338 = ~n14334 & n14337;
  assign n14339 = pi778 & ~n14338;
  assign n14340 = ~n14336 & n14339;
  assign n14341 = ~n14333 & ~n14340;
  assign n14342 = ~n7949 & ~n14341;
  assign n14343 = ~n7951 & n14342;
  assign n14344 = ~n7953 & n14343;
  assign n14345 = ~n7955 & n14344;
  assign n14346 = ~n7967 & n14345;
  assign n14347 = pi647 & ~n14346;
  assign n14348 = ~pi647 & ~n14290;
  assign n14349 = ~n14347 & ~n14348;
  assign n14350 = n7832 & ~n14349;
  assign n14351 = ~pi647 & n14346;
  assign n14352 = pi647 & n14290;
  assign n14353 = ~pi1157 & ~n14352;
  assign n14354 = ~n14351 & n14353;
  assign n14355 = pi630 & n14354;
  assign n14356 = ~n14350 & ~n14355;
  assign n14357 = ~n59492 & n14356;
  assign n14358 = pi787 & ~n14357;
  assign n14359 = ~pi626 & ~n14318;
  assign n14360 = pi626 & ~n14290;
  assign n14361 = n7760 & ~n14360;
  assign n14362 = ~n14359 & n14361;
  assign n14363 = n7984 & n14344;
  assign n14364 = pi626 & ~n14318;
  assign n14365 = ~pi626 & ~n14290;
  assign n14366 = n7759 & ~n14365;
  assign n14367 = ~n14364 & n14366;
  assign n14368 = ~n14363 & ~n14367;
  assign n14369 = ~n14362 & ~n14363;
  assign n14370 = ~n14367 & n14369;
  assign n14371 = ~n14362 & n14368;
  assign n14372 = pi788 & ~n59493;
  assign n14373 = ~n6701 & ~n14332;
  assign n14374 = pi625 & n14373;
  assign n14375 = n14292 & ~n14373;
  assign n14376 = ~n14374 & ~n14375;
  assign n14377 = n14337 & ~n14376;
  assign n14378 = ~pi608 & ~n14336;
  assign n14379 = ~n14377 & n14378;
  assign n14380 = pi1153 & n14292;
  assign n14381 = ~n14374 & n14380;
  assign n14382 = pi608 & ~n14338;
  assign n14383 = ~n14381 & n14382;
  assign n14384 = ~n14379 & ~n14383;
  assign n14385 = pi778 & ~n14384;
  assign n14386 = ~pi778 & ~n14375;
  assign n14387 = ~n14385 & ~n14386;
  assign n14388 = ~pi609 & ~n14387;
  assign n14389 = pi609 & ~n14341;
  assign n14390 = ~pi1155 & ~n14389;
  assign n14391 = ~n14388 & n14390;
  assign n14392 = ~pi660 & ~n14297;
  assign n14393 = ~n14391 & n14392;
  assign n14394 = pi609 & ~n14387;
  assign n14395 = ~pi609 & ~n14341;
  assign n14396 = pi1155 & ~n14395;
  assign n14397 = ~n14394 & n14396;
  assign n14398 = pi660 & ~n14299;
  assign n14399 = ~n14397 & n14398;
  assign n14400 = ~n14393 & ~n14399;
  assign n14401 = pi785 & ~n14400;
  assign n14402 = ~pi785 & ~n14387;
  assign n14403 = ~n14401 & ~n14402;
  assign n14404 = ~pi618 & ~n14403;
  assign n14405 = pi618 & n14342;
  assign n14406 = ~pi1154 & ~n14405;
  assign n14407 = ~n14404 & n14406;
  assign n14408 = ~pi627 & ~n14305;
  assign n14409 = ~n14407 & n14408;
  assign n14410 = pi618 & ~n14403;
  assign n14411 = ~pi618 & n14342;
  assign n14412 = pi1154 & ~n14411;
  assign n14413 = ~n14410 & n14412;
  assign n14414 = pi627 & ~n14307;
  assign n14415 = ~n14413 & n14414;
  assign n14416 = ~n14409 & ~n14415;
  assign n14417 = pi781 & ~n14416;
  assign n14418 = ~pi781 & ~n14403;
  assign n14419 = ~n14417 & ~n14418;
  assign n14420 = pi619 & ~n14419;
  assign n14421 = ~pi619 & n14343;
  assign n14422 = pi1159 & ~n14421;
  assign n14423 = ~n14420 & n14422;
  assign n14424 = pi648 & ~n14315;
  assign n14425 = ~n14423 & n14424;
  assign n14426 = ~pi619 & ~n14419;
  assign n14427 = pi619 & n14343;
  assign n14428 = ~pi1159 & ~n14427;
  assign n14429 = ~n14426 & n14428;
  assign n14430 = ~pi648 & ~n14313;
  assign n14431 = ~n14429 & n14430;
  assign n14432 = pi789 & ~n14431;
  assign n14433 = pi789 & ~n14425;
  assign n14434 = ~n14431 & n14433;
  assign n14435 = ~n14425 & n14432;
  assign n14436 = ~pi789 & n14419;
  assign n14437 = n59242 & ~n14436;
  assign n14438 = ~n59494 & n14437;
  assign n14439 = ~n14372 & ~n14438;
  assign n14440 = ~n59357 & ~n14439;
  assign n14441 = n7957 & ~n59491;
  assign n14442 = n8065 & n14345;
  assign n14443 = pi629 & ~n14442;
  assign n14444 = ~n14441 & n14443;
  assign n14445 = n7958 & ~n59491;
  assign n14446 = n8074 & n14345;
  assign n14447 = ~pi629 & ~n14446;
  assign n14448 = ~n14445 & n14447;
  assign n14449 = pi792 & ~n14448;
  assign n14450 = ~n14445 & ~n14446;
  assign n14451 = ~pi629 & ~n14450;
  assign n14452 = ~n14441 & ~n14442;
  assign n14453 = pi629 & ~n14452;
  assign n14454 = ~n14451 & ~n14453;
  assign n14455 = pi792 & ~n14454;
  assign n14456 = pi792 & ~n14444;
  assign n14457 = ~n14448 & n14456;
  assign n14458 = ~n14444 & n14449;
  assign n14459 = ~n8108 & ~n59495;
  assign n14460 = ~n14440 & n14459;
  assign n14461 = ~n14358 & ~n14460;
  assign n14462 = pi644 & n14461;
  assign n14463 = ~pi787 & ~n14346;
  assign n14464 = pi1157 & ~n14349;
  assign n14465 = ~n14354 & ~n14464;
  assign n14466 = pi787 & ~n14465;
  assign n14467 = ~n14463 & ~n14466;
  assign n14468 = ~pi644 & n14467;
  assign n14469 = pi715 & ~n14468;
  assign n14470 = ~n14462 & n14469;
  assign n14471 = ~n11491 & n14290;
  assign n14472 = ~n7835 & n14325;
  assign n14473 = ~n7835 & ~n14328;
  assign n14474 = n7835 & n14290;
  assign n14475 = ~n14473 & ~n14474;
  assign n14476 = ~n14471 & ~n14472;
  assign n14477 = pi644 & ~n59496;
  assign n14478 = ~pi644 & n14290;
  assign n14479 = ~pi715 & ~n14478;
  assign n14480 = ~n14477 & n14479;
  assign n14481 = pi1160 & ~n14480;
  assign n14482 = ~n14470 & n14481;
  assign n14483 = ~pi644 & n14461;
  assign n14484 = pi644 & n14467;
  assign n14485 = ~pi715 & ~n14484;
  assign n14486 = ~n14483 & n14485;
  assign n14487 = ~pi644 & ~n59496;
  assign n14488 = pi644 & n14290;
  assign n14489 = pi715 & ~n14488;
  assign n14490 = ~n14487 & n14489;
  assign n14491 = ~pi1160 & ~n14490;
  assign n14492 = ~n14486 & n14491;
  assign n14493 = ~n14482 & ~n14492;
  assign n14494 = pi790 & ~n14493;
  assign n14495 = ~pi790 & n14461;
  assign n14496 = pi832 & ~n14495;
  assign n14497 = ~n14494 & n14496;
  assign n14498 = ~pi178 & ~n7560;
  assign n14499 = n59231 & ~n14498;
  assign n14500 = ~pi688 & n59132;
  assign n14501 = n14498 & ~n14500;
  assign n14502 = pi178 & n59251;
  assign n14503 = ~pi38 & ~n14502;
  assign n14504 = n59132 & ~n14503;
  assign n14505 = ~pi178 & n8249;
  assign n14506 = ~n14504 & ~n14505;
  assign n14507 = ~pi178 & ~n6863;
  assign n14508 = n7547 & ~n14507;
  assign n14509 = ~pi688 & ~n14508;
  assign n14510 = ~n14506 & n14509;
  assign n14511 = ~n14501 & ~n14510;
  assign n14512 = ~pi778 & n14511;
  assign n14513 = pi625 & ~n14511;
  assign n14514 = ~pi625 & n14498;
  assign n14515 = pi1153 & ~n14514;
  assign n14516 = ~n14513 & n14515;
  assign n14517 = ~pi625 & ~n14511;
  assign n14518 = pi625 & n14498;
  assign n14519 = ~pi1153 & ~n14518;
  assign n14520 = ~n14517 & n14519;
  assign n14521 = ~n14516 & ~n14520;
  assign n14522 = pi778 & ~n14521;
  assign n14523 = ~n14512 & ~n14522;
  assign n14524 = ~n59229 & n14523;
  assign n14525 = n59229 & n14498;
  assign n14526 = n59229 & ~n14498;
  assign n14527 = ~n59229 & ~n14523;
  assign n14528 = ~n14526 & ~n14527;
  assign n14529 = ~n14524 & ~n14525;
  assign n14530 = ~n59231 & ~n59497;
  assign n14531 = ~n59231 & n59497;
  assign n14532 = n59231 & n14498;
  assign n14533 = ~n14531 & ~n14532;
  assign n14534 = ~n14499 & ~n14530;
  assign n14535 = ~n7716 & ~n59498;
  assign n14536 = n7716 & n14498;
  assign n14537 = n7716 & ~n14498;
  assign n14538 = ~n7716 & n59498;
  assign n14539 = ~n14537 & ~n14538;
  assign n14540 = ~n14535 & ~n14536;
  assign n14541 = ~n7762 & n59499;
  assign n14542 = n7762 & n14498;
  assign n14543 = ~n14541 & ~n14542;
  assign n14544 = ~pi792 & n14543;
  assign n14545 = pi628 & ~n14543;
  assign n14546 = ~pi628 & n14498;
  assign n14547 = pi1156 & ~n14546;
  assign n14548 = ~n14545 & n14547;
  assign n14549 = ~pi628 & ~n14543;
  assign n14550 = pi628 & n14498;
  assign n14551 = ~pi1156 & ~n14550;
  assign n14552 = ~n14549 & n14551;
  assign n14553 = ~n14548 & ~n14552;
  assign n14554 = pi792 & ~n14553;
  assign n14555 = ~n14544 & ~n14554;
  assign n14556 = pi647 & n14555;
  assign n14557 = ~pi647 & n14498;
  assign n14558 = pi647 & ~n14555;
  assign n14559 = ~pi647 & ~n14498;
  assign n14560 = ~n14558 & ~n14559;
  assign n14561 = ~n14556 & ~n14557;
  assign n14562 = pi1157 & ~n59500;
  assign n14563 = ~pi647 & n14555;
  assign n14564 = pi647 & n14498;
  assign n14565 = ~pi1157 & ~n14564;
  assign n14566 = ~n14563 & n14565;
  assign n14567 = ~pi647 & ~n14555;
  assign n14568 = pi647 & ~n14498;
  assign n14569 = ~n14567 & ~n14568;
  assign n14570 = ~pi1157 & n14569;
  assign n14571 = pi1157 & n59500;
  assign n14572 = ~n14570 & ~n14571;
  assign n14573 = ~n14562 & ~n14566;
  assign n14574 = pi787 & n59501;
  assign n14575 = ~pi787 & ~n14555;
  assign n14576 = pi787 & ~n59501;
  assign n14577 = ~pi787 & n14555;
  assign n14578 = ~n14576 & ~n14577;
  assign n14579 = ~n14574 & ~n14575;
  assign n14580 = ~pi644 & ~n59502;
  assign n14581 = pi715 & ~n14580;
  assign n14582 = pi178 & ~n59132;
  assign n14583 = ~pi760 & n6865;
  assign n14584 = ~n14507 & ~n14583;
  assign n14585 = pi38 & ~n14584;
  assign n14586 = ~pi178 & n59164;
  assign n14587 = pi178 & ~n6855;
  assign n14588 = ~pi760 & ~n14587;
  assign n14589 = ~n14586 & n14588;
  assign n14590 = ~pi178 & pi760;
  assign n14591 = ~n6656 & n14590;
  assign n14592 = pi760 & ~n6656;
  assign n14593 = ~pi760 & ~n14586;
  assign n14594 = ~n14592 & ~n14593;
  assign n14595 = ~pi178 & ~n14594;
  assign n14596 = n6855 & n14593;
  assign n14597 = ~n14595 & ~n14596;
  assign n14598 = ~n14589 & ~n14591;
  assign n14599 = ~pi38 & ~n59503;
  assign n14600 = ~n14585 & ~n14599;
  assign n14601 = n59132 & n14600;
  assign n14602 = ~n14582 & ~n14601;
  assign n14603 = ~n7597 & ~n14602;
  assign n14604 = n7597 & ~n14498;
  assign n14605 = ~n14603 & ~n14604;
  assign n14606 = ~pi785 & ~n14605;
  assign n14607 = ~n7598 & ~n14498;
  assign n14608 = pi609 & n14603;
  assign n14609 = ~n14607 & ~n14608;
  assign n14610 = pi1155 & ~n14609;
  assign n14611 = ~n7610 & ~n14498;
  assign n14612 = ~pi609 & n14603;
  assign n14613 = ~n14611 & ~n14612;
  assign n14614 = ~pi1155 & ~n14613;
  assign n14615 = ~n14610 & ~n14614;
  assign n14616 = pi785 & ~n14615;
  assign n14617 = ~n14606 & ~n14616;
  assign n14618 = ~pi781 & ~n14617;
  assign n14619 = pi618 & n14617;
  assign n14620 = ~pi618 & n14498;
  assign n14621 = pi1154 & ~n14620;
  assign n14622 = ~n14619 & n14621;
  assign n14623 = ~pi618 & n14617;
  assign n14624 = pi618 & n14498;
  assign n14625 = ~pi1154 & ~n14624;
  assign n14626 = ~n14623 & n14625;
  assign n14627 = ~n14622 & ~n14626;
  assign n14628 = pi781 & ~n14627;
  assign n14629 = ~n14618 & ~n14628;
  assign n14630 = ~pi789 & ~n14629;
  assign n14631 = pi619 & n14629;
  assign n14632 = ~pi619 & n14498;
  assign n14633 = pi1159 & ~n14632;
  assign n14634 = ~n14631 & n14633;
  assign n14635 = ~pi619 & n14629;
  assign n14636 = pi619 & n14498;
  assign n14637 = ~pi1159 & ~n14636;
  assign n14638 = ~n14635 & n14637;
  assign n14639 = ~n14634 & ~n14638;
  assign n14640 = pi789 & ~n14639;
  assign n14641 = ~n14630 & ~n14640;
  assign n14642 = ~n8054 & n14641;
  assign n14643 = n8054 & n14498;
  assign n14644 = ~n14642 & ~n14643;
  assign n14645 = ~n7793 & ~n14644;
  assign n14646 = n7793 & n14498;
  assign n14647 = ~n14645 & ~n14646;
  assign n14648 = ~n7835 & ~n14647;
  assign n14649 = n7835 & n14498;
  assign n14650 = n7835 & ~n14498;
  assign n14651 = ~n7835 & n14647;
  assign n14652 = ~n14650 & ~n14651;
  assign n14653 = ~n14648 & ~n14649;
  assign n14654 = pi644 & n59504;
  assign n14655 = ~pi644 & n14498;
  assign n14656 = ~pi715 & ~n14655;
  assign n14657 = ~n14654 & n14656;
  assign n14658 = pi1160 & ~n14657;
  assign n14659 = ~n14581 & n14658;
  assign n14660 = pi644 & ~n59502;
  assign n14661 = ~pi715 & ~n14660;
  assign n14662 = ~pi644 & n59504;
  assign n14663 = pi644 & n14498;
  assign n14664 = pi715 & ~n14663;
  assign n14665 = ~n14662 & n14664;
  assign n14666 = ~pi1160 & ~n14665;
  assign n14667 = ~n14661 & n14666;
  assign n14668 = ~n14659 & ~n14667;
  assign n14669 = pi790 & ~n14668;
  assign n14670 = ~pi644 & n14666;
  assign n14671 = pi644 & n14658;
  assign n14672 = pi790 & ~n14671;
  assign n14673 = pi790 & ~n14670;
  assign n14674 = ~n14671 & n14673;
  assign n14675 = ~n14670 & n14672;
  assign n14676 = ~n7872 & n14647;
  assign n14677 = n7832 & ~n59500;
  assign n14678 = n7833 & ~n14569;
  assign n14679 = pi630 & n14566;
  assign n14680 = ~n14677 & ~n59506;
  assign n14681 = ~n14676 & n14680;
  assign n14682 = pi787 & ~n14681;
  assign n14683 = ~n11154 & n14644;
  assign n14684 = ~pi629 & n14548;
  assign n14685 = pi629 & n14552;
  assign n14686 = ~n14684 & ~n14685;
  assign n14687 = ~n14683 & n14686;
  assign n14688 = pi792 & ~n14687;
  assign n14689 = pi688 & ~n14600;
  assign n14690 = ~pi178 & n59177;
  assign n14691 = pi178 & n7111;
  assign n14692 = pi760 & ~n14691;
  assign n14693 = ~n14690 & n14692;
  assign n14694 = pi178 & n7188;
  assign n14695 = ~pi178 & ~n59203;
  assign n14696 = ~pi760 & ~n14695;
  assign n14697 = ~n14694 & n14696;
  assign n14698 = pi39 & ~n14697;
  assign n14699 = ~n14693 & n14698;
  assign n14700 = pi178 & n7333;
  assign n14701 = ~pi178 & n7310;
  assign n14702 = pi760 & ~n14701;
  assign n14703 = ~n14700 & n14702;
  assign n14704 = ~pi178 & ~n7339;
  assign n14705 = pi178 & ~n7347;
  assign n14706 = ~pi760 & ~n14705;
  assign n14707 = ~n14704 & n14706;
  assign n14708 = ~pi39 & ~n14707;
  assign n14709 = pi178 & ~n7333;
  assign n14710 = ~pi178 & ~n7310;
  assign n14711 = pi760 & ~n14710;
  assign n14712 = pi760 & ~n14709;
  assign n14713 = ~n14710 & n14712;
  assign n14714 = ~n14709 & n14711;
  assign n14715 = ~pi178 & n7339;
  assign n14716 = pi178 & n7347;
  assign n14717 = ~pi760 & ~n14716;
  assign n14718 = ~n14715 & n14717;
  assign n14719 = ~n59507 & ~n14718;
  assign n14720 = ~pi39 & ~n14719;
  assign n14721 = ~n14703 & n14708;
  assign n14722 = ~pi38 & ~n59508;
  assign n14723 = ~n14699 & n14722;
  assign n14724 = ~pi760 & ~n7222;
  assign n14725 = n9794 & ~n14724;
  assign n14726 = ~pi178 & ~n14725;
  assign n14727 = ~n7056 & ~n14291;
  assign n14728 = pi178 & ~n14727;
  assign n14729 = n59171 & n14728;
  assign n14730 = pi38 & ~n14729;
  assign n14731 = ~n14726 & n14730;
  assign n14732 = ~pi688 & ~n14731;
  assign n14733 = ~n14723 & n14732;
  assign n14734 = n59132 & ~n14733;
  assign n14735 = ~n14689 & n14734;
  assign n14736 = ~n14582 & ~n14735;
  assign n14737 = ~pi625 & n14736;
  assign n14738 = pi625 & n14602;
  assign n14739 = ~pi1153 & ~n14738;
  assign n14740 = ~n14737 & n14739;
  assign n14741 = ~pi608 & ~n14516;
  assign n14742 = ~n14740 & n14741;
  assign n14743 = pi625 & n14736;
  assign n14744 = ~pi625 & n14602;
  assign n14745 = pi1153 & ~n14744;
  assign n14746 = ~n14743 & n14745;
  assign n14747 = pi608 & ~n14520;
  assign n14748 = ~n14746 & n14747;
  assign n14749 = ~n14742 & ~n14748;
  assign n14750 = pi778 & ~n14749;
  assign n14751 = ~pi778 & n14736;
  assign n14752 = ~n14750 & ~n14751;
  assign n14753 = ~pi609 & ~n14752;
  assign n14754 = pi609 & n14523;
  assign n14755 = ~pi1155 & ~n14754;
  assign n14756 = ~n14753 & n14755;
  assign n14757 = ~pi660 & ~n14610;
  assign n14758 = ~n14756 & n14757;
  assign n14759 = pi609 & ~n14752;
  assign n14760 = ~pi609 & n14523;
  assign n14761 = pi1155 & ~n14760;
  assign n14762 = ~n14759 & n14761;
  assign n14763 = pi660 & ~n14614;
  assign n14764 = ~n14762 & n14763;
  assign n14765 = ~n14758 & ~n14764;
  assign n14766 = pi785 & ~n14765;
  assign n14767 = ~pi785 & ~n14752;
  assign n14768 = ~n14766 & ~n14767;
  assign n14769 = ~pi618 & ~n14768;
  assign n14770 = pi618 & n59497;
  assign n14771 = ~pi1154 & ~n14770;
  assign n14772 = ~n14769 & n14771;
  assign n14773 = ~pi627 & ~n14622;
  assign n14774 = ~n14772 & n14773;
  assign n14775 = pi618 & ~n14768;
  assign n14776 = ~pi618 & n59497;
  assign n14777 = pi1154 & ~n14776;
  assign n14778 = ~n14775 & n14777;
  assign n14779 = pi627 & ~n14626;
  assign n14780 = ~n14778 & n14779;
  assign n14781 = ~n14774 & ~n14780;
  assign n14782 = pi781 & ~n14781;
  assign n14783 = ~pi781 & ~n14768;
  assign n14784 = ~n14782 & ~n14783;
  assign n14785 = pi619 & ~n14784;
  assign n14786 = ~pi619 & ~n59498;
  assign n14787 = pi1159 & ~n14786;
  assign n14788 = ~n14785 & n14787;
  assign n14789 = pi648 & ~n14638;
  assign n14790 = ~n14788 & n14789;
  assign n14791 = ~pi619 & ~n14784;
  assign n14792 = pi619 & ~n59498;
  assign n14793 = ~pi1159 & ~n14792;
  assign n14794 = ~n14791 & n14793;
  assign n14795 = ~pi648 & ~n14634;
  assign n14796 = ~n14794 & n14795;
  assign n14797 = pi789 & ~n14796;
  assign n14798 = pi789 & ~n14790;
  assign n14799 = ~n14796 & n14798;
  assign n14800 = ~n14790 & n14797;
  assign n14801 = ~pi789 & n14784;
  assign n14802 = n59242 & ~n14801;
  assign n14803 = ~n59509 & n14802;
  assign n14804 = ~pi626 & ~n14641;
  assign n14805 = pi626 & ~n14498;
  assign n14806 = n7760 & ~n14805;
  assign n14807 = ~n14804 & n14806;
  assign n14808 = n7984 & n59499;
  assign n14809 = pi626 & ~n14641;
  assign n14810 = ~pi626 & ~n14498;
  assign n14811 = n7759 & ~n14810;
  assign n14812 = ~n14809 & n14811;
  assign n14813 = ~n14808 & ~n14812;
  assign n14814 = ~n14807 & ~n14808;
  assign n14815 = ~n14812 & n14814;
  assign n14816 = ~n14807 & n14813;
  assign n14817 = pi788 & ~n59510;
  assign n14818 = ~n59357 & ~n14817;
  assign n14819 = ~n14803 & n14818;
  assign n14820 = ~n14688 & ~n14819;
  assign n14821 = ~n8108 & ~n14820;
  assign n14822 = ~n14682 & ~n14821;
  assign n14823 = ~n59505 & n14822;
  assign n14824 = ~n14669 & ~n14823;
  assign n14825 = n58992 & ~n14824;
  assign n14826 = ~pi178 & ~n58992;
  assign n14827 = ~pi832 & ~n14826;
  assign n14828 = ~n14825 & n14827;
  assign po335 = ~n14497 & ~n14828;
  assign n14830 = ~pi179 & ~n2794;
  assign n14831 = ~pi741 & n6822;
  assign n14832 = ~n14830 & ~n14831;
  assign n14833 = ~n7875 & ~n14832;
  assign n14834 = ~pi785 & ~n14833;
  assign n14835 = ~n7880 & ~n14832;
  assign n14836 = pi1155 & ~n14835;
  assign n14837 = ~n7883 & n14833;
  assign n14838 = ~pi1155 & ~n14837;
  assign n14839 = ~n14836 & ~n14838;
  assign n14840 = pi785 & ~n14839;
  assign n14841 = ~n14834 & ~n14840;
  assign n14842 = ~pi781 & ~n14841;
  assign n14843 = ~n7890 & n14841;
  assign n14844 = pi1154 & ~n14843;
  assign n14845 = ~n7893 & n14841;
  assign n14846 = ~pi1154 & ~n14845;
  assign n14847 = ~n14844 & ~n14846;
  assign n14848 = pi781 & ~n14847;
  assign n14849 = ~n14842 & ~n14848;
  assign n14850 = ~pi789 & ~n14849;
  assign n14851 = pi619 & n14849;
  assign n14852 = ~pi619 & n14830;
  assign n14853 = pi1159 & ~n14852;
  assign n14854 = ~n14851 & n14853;
  assign n14855 = ~pi619 & n14849;
  assign n14856 = pi619 & n14830;
  assign n14857 = ~pi1159 & ~n14856;
  assign n14858 = ~n14855 & n14857;
  assign n14859 = ~n14854 & ~n14858;
  assign n14860 = pi789 & ~n14859;
  assign n14861 = ~n14850 & ~n14860;
  assign n14862 = ~n8054 & ~n14861;
  assign n14863 = n8054 & ~n14830;
  assign n14864 = ~n8054 & n14861;
  assign n14865 = n8054 & n14830;
  assign n14866 = ~n14864 & ~n14865;
  assign n14867 = ~n14862 & ~n14863;
  assign n14868 = ~n7793 & ~n59511;
  assign n14869 = n7793 & n14830;
  assign n14870 = ~n7872 & ~n14869;
  assign n14871 = ~n14868 & ~n14869;
  assign n14872 = ~n7872 & n14871;
  assign n14873 = ~n14868 & n14870;
  assign n14874 = ~pi724 & n7055;
  assign n14875 = ~n14830 & ~n14874;
  assign n14876 = ~pi778 & n14875;
  assign n14877 = ~pi625 & n14874;
  assign n14878 = ~n14875 & ~n14877;
  assign n14879 = pi1153 & ~n14878;
  assign n14880 = ~pi1153 & ~n14830;
  assign n14881 = ~n14877 & n14880;
  assign n14882 = ~n14879 & ~n14881;
  assign n14883 = pi778 & ~n14882;
  assign n14884 = ~n14876 & ~n14883;
  assign n14885 = ~n7949 & n14884;
  assign n14886 = ~n7951 & n14885;
  assign n14887 = ~n7953 & n14886;
  assign n14888 = ~n7955 & n14887;
  assign n14889 = ~n7967 & n14888;
  assign n14890 = pi647 & ~n14889;
  assign n14891 = ~pi647 & ~n14830;
  assign n14892 = ~n14890 & ~n14891;
  assign n14893 = n7832 & ~n14892;
  assign n14894 = ~pi647 & n14889;
  assign n14895 = pi647 & n14830;
  assign n14896 = ~pi1157 & ~n14895;
  assign n14897 = ~n14894 & n14896;
  assign n14898 = pi630 & n14897;
  assign n14899 = ~n14893 & ~n14898;
  assign n14900 = ~n59512 & n14899;
  assign n14901 = pi787 & ~n14900;
  assign n14902 = ~pi626 & ~n14861;
  assign n14903 = pi626 & ~n14830;
  assign n14904 = n7760 & ~n14903;
  assign n14905 = ~n14902 & n14904;
  assign n14906 = n7984 & n14887;
  assign n14907 = pi626 & ~n14861;
  assign n14908 = ~pi626 & ~n14830;
  assign n14909 = n7759 & ~n14908;
  assign n14910 = ~n14907 & n14909;
  assign n14911 = ~n14906 & ~n14910;
  assign n14912 = ~n14905 & ~n14906;
  assign n14913 = ~n14910 & n14912;
  assign n14914 = ~n14905 & n14911;
  assign n14915 = pi788 & ~n59513;
  assign n14916 = ~n6701 & ~n14875;
  assign n14917 = pi625 & n14916;
  assign n14918 = n14832 & ~n14916;
  assign n14919 = ~n14917 & ~n14918;
  assign n14920 = n14880 & ~n14919;
  assign n14921 = ~pi608 & ~n14879;
  assign n14922 = ~n14920 & n14921;
  assign n14923 = pi1153 & n14832;
  assign n14924 = ~n14917 & n14923;
  assign n14925 = pi608 & ~n14881;
  assign n14926 = ~n14924 & n14925;
  assign n14927 = ~n14922 & ~n14926;
  assign n14928 = pi778 & ~n14927;
  assign n14929 = ~pi778 & ~n14918;
  assign n14930 = ~n14928 & ~n14929;
  assign n14931 = ~pi609 & ~n14930;
  assign n14932 = pi609 & n14884;
  assign n14933 = ~pi1155 & ~n14932;
  assign n14934 = ~n14931 & n14933;
  assign n14935 = ~pi660 & ~n14836;
  assign n14936 = ~n14934 & n14935;
  assign n14937 = pi609 & ~n14930;
  assign n14938 = ~pi609 & n14884;
  assign n14939 = pi1155 & ~n14938;
  assign n14940 = ~n14937 & n14939;
  assign n14941 = pi660 & ~n14838;
  assign n14942 = ~n14940 & n14941;
  assign n14943 = ~n14936 & ~n14942;
  assign n14944 = pi785 & ~n14943;
  assign n14945 = ~pi785 & ~n14930;
  assign n14946 = ~n14944 & ~n14945;
  assign n14947 = ~pi618 & ~n14946;
  assign n14948 = pi618 & n14885;
  assign n14949 = ~pi1154 & ~n14948;
  assign n14950 = ~n14947 & n14949;
  assign n14951 = ~pi627 & ~n14844;
  assign n14952 = ~n14950 & n14951;
  assign n14953 = pi618 & ~n14946;
  assign n14954 = ~pi618 & n14885;
  assign n14955 = pi1154 & ~n14954;
  assign n14956 = ~n14953 & n14955;
  assign n14957 = pi627 & ~n14846;
  assign n14958 = ~n14956 & n14957;
  assign n14959 = ~n14952 & ~n14958;
  assign n14960 = pi781 & ~n14959;
  assign n14961 = ~pi781 & ~n14946;
  assign n14962 = ~n14960 & ~n14961;
  assign n14963 = ~pi619 & ~n14962;
  assign n14964 = pi619 & n14886;
  assign n14965 = ~pi1159 & ~n14964;
  assign n14966 = ~n14963 & n14965;
  assign n14967 = ~pi648 & ~n14854;
  assign n14968 = ~n14966 & n14967;
  assign n14969 = pi619 & ~n14962;
  assign n14970 = ~pi619 & n14886;
  assign n14971 = pi1159 & ~n14970;
  assign n14972 = ~n14969 & n14971;
  assign n14973 = pi648 & ~n14858;
  assign n14974 = ~n14972 & n14973;
  assign n14975 = pi789 & ~n14974;
  assign n14976 = pi789 & ~n14968;
  assign n14977 = ~n14974 & n14976;
  assign n14978 = ~n14968 & n14975;
  assign n14979 = ~pi789 & n14962;
  assign n14980 = n59242 & ~n14979;
  assign n14981 = ~n59514 & n14980;
  assign n14982 = ~n14915 & ~n14981;
  assign n14983 = ~n59357 & ~n14982;
  assign n14984 = n7957 & ~n59511;
  assign n14985 = n8065 & n14888;
  assign n14986 = pi629 & ~n14985;
  assign n14987 = ~n14984 & n14986;
  assign n14988 = n7958 & ~n59511;
  assign n14989 = n8074 & n14888;
  assign n14990 = ~pi629 & ~n14989;
  assign n14991 = ~n14988 & n14990;
  assign n14992 = pi792 & ~n14991;
  assign n14993 = ~n14988 & ~n14989;
  assign n14994 = ~pi629 & ~n14993;
  assign n14995 = ~n14984 & ~n14985;
  assign n14996 = pi629 & ~n14995;
  assign n14997 = ~n14994 & ~n14996;
  assign n14998 = pi792 & ~n14997;
  assign n14999 = pi792 & ~n14987;
  assign n15000 = ~n14991 & n14999;
  assign n15001 = ~n14987 & n14992;
  assign n15002 = ~n8108 & ~n59515;
  assign n15003 = ~n14983 & n15002;
  assign n15004 = ~n14901 & ~n15003;
  assign n15005 = pi644 & n15004;
  assign n15006 = ~pi787 & ~n14889;
  assign n15007 = pi1157 & ~n14892;
  assign n15008 = ~n14897 & ~n15007;
  assign n15009 = pi787 & ~n15008;
  assign n15010 = ~n15006 & ~n15009;
  assign n15011 = ~pi644 & n15010;
  assign n15012 = pi715 & ~n15011;
  assign n15013 = ~n15005 & n15012;
  assign n15014 = ~n11491 & n14830;
  assign n15015 = ~n7835 & n14868;
  assign n15016 = ~n7835 & ~n14871;
  assign n15017 = n7835 & n14830;
  assign n15018 = ~n15016 & ~n15017;
  assign n15019 = ~n15014 & ~n15015;
  assign n15020 = pi644 & ~n59516;
  assign n15021 = ~pi644 & n14830;
  assign n15022 = ~pi715 & ~n15021;
  assign n15023 = ~n15020 & n15022;
  assign n15024 = pi1160 & ~n15023;
  assign n15025 = ~n15013 & n15024;
  assign n15026 = ~pi644 & n15004;
  assign n15027 = pi644 & n15010;
  assign n15028 = ~pi715 & ~n15027;
  assign n15029 = ~n15026 & n15028;
  assign n15030 = ~pi644 & ~n59516;
  assign n15031 = pi644 & n14830;
  assign n15032 = pi715 & ~n15031;
  assign n15033 = ~n15030 & n15032;
  assign n15034 = ~pi1160 & ~n15033;
  assign n15035 = ~n15029 & n15034;
  assign n15036 = ~n15025 & ~n15035;
  assign n15037 = pi790 & ~n15036;
  assign n15038 = ~pi790 & n15004;
  assign n15039 = pi832 & ~n15038;
  assign n15040 = ~n15037 & n15039;
  assign n15041 = ~pi179 & ~n7560;
  assign n15042 = n7762 & ~n15041;
  assign n15043 = n59231 & ~n15041;
  assign n15044 = ~pi724 & n59132;
  assign n15045 = n15041 & ~n15044;
  assign n15046 = ~pi179 & n8249;
  assign n15047 = pi179 & n59251;
  assign n15048 = ~pi38 & ~n15047;
  assign n15049 = n59132 & ~n15048;
  assign n15050 = ~n15046 & ~n15049;
  assign n15051 = ~pi179 & ~n6863;
  assign n15052 = n7547 & ~n15051;
  assign n15053 = ~pi724 & ~n15052;
  assign n15054 = ~n15050 & n15053;
  assign n15055 = ~n15045 & ~n15054;
  assign n15056 = ~pi778 & n15055;
  assign n15057 = ~pi625 & ~n15055;
  assign n15058 = pi625 & n15041;
  assign n15059 = ~pi1153 & ~n15058;
  assign n15060 = ~n15057 & n15059;
  assign n15061 = pi625 & ~n15055;
  assign n15062 = ~pi625 & n15041;
  assign n15063 = pi1153 & ~n15062;
  assign n15064 = ~n15061 & n15063;
  assign n15065 = ~n15060 & ~n15064;
  assign n15066 = pi778 & ~n15065;
  assign n15067 = ~n15056 & ~n15066;
  assign n15068 = ~n59229 & n15067;
  assign n15069 = n59229 & n15041;
  assign n15070 = n59229 & ~n15041;
  assign n15071 = ~n59229 & ~n15067;
  assign n15072 = ~n15070 & ~n15071;
  assign n15073 = ~n15068 & ~n15069;
  assign n15074 = ~n59231 & ~n59517;
  assign n15075 = ~n59231 & n59517;
  assign n15076 = n59231 & n15041;
  assign n15077 = ~n15075 & ~n15076;
  assign n15078 = ~n15043 & ~n15074;
  assign n15079 = ~n7716 & ~n59518;
  assign n15080 = n7716 & n15041;
  assign n15081 = n7716 & ~n15041;
  assign n15082 = ~n7716 & n59518;
  assign n15083 = ~n15081 & ~n15082;
  assign n15084 = ~n15079 & ~n15080;
  assign n15085 = ~n7762 & ~n59519;
  assign n15086 = ~n7762 & n59519;
  assign n15087 = n7762 & n15041;
  assign n15088 = ~n15086 & ~n15087;
  assign n15089 = ~n15042 & ~n15085;
  assign n15090 = pi628 & ~n59520;
  assign n15091 = ~pi628 & n15041;
  assign n15092 = pi1156 & ~n15091;
  assign n15093 = ~n15090 & n15092;
  assign n15094 = ~pi628 & ~n59520;
  assign n15095 = pi628 & n15041;
  assign n15096 = ~pi1156 & ~n15095;
  assign n15097 = ~n15094 & n15096;
  assign n15098 = pi628 & ~n15041;
  assign n15099 = ~pi628 & n59520;
  assign n15100 = ~n15098 & ~n15099;
  assign n15101 = ~pi1156 & n15100;
  assign n15102 = ~pi628 & ~n15041;
  assign n15103 = pi628 & n59520;
  assign n15104 = ~n15102 & ~n15103;
  assign n15105 = pi1156 & n15104;
  assign n15106 = ~n15101 & ~n15105;
  assign n15107 = ~n15093 & ~n15097;
  assign n15108 = pi792 & ~n59521;
  assign n15109 = ~pi792 & ~n59520;
  assign n15110 = ~pi792 & n59520;
  assign n15111 = pi792 & n59521;
  assign n15112 = ~n15110 & ~n15111;
  assign n15113 = ~n15108 & ~n15109;
  assign n15114 = pi647 & n59522;
  assign n15115 = ~pi647 & n15041;
  assign n15116 = ~n15114 & ~n15115;
  assign n15117 = n7832 & n15116;
  assign n15118 = ~pi647 & n59522;
  assign n15119 = pi647 & n15041;
  assign n15120 = ~pi1157 & ~n15119;
  assign n15121 = ~n15118 & n15120;
  assign n15122 = pi630 & n15121;
  assign n15123 = pi179 & ~n59132;
  assign n15124 = pi741 & n7553;
  assign n15125 = ~pi179 & ~pi741;
  assign n15126 = ~n9780 & n15125;
  assign n15127 = n9787 & n15126;
  assign n15128 = n9787 & n15125;
  assign n15129 = ~pi741 & ~n13474;
  assign n15130 = pi179 & ~n15129;
  assign n15131 = ~n59523 & ~n15130;
  assign n15132 = ~n15124 & n15131;
  assign n15133 = n59132 & ~n15132;
  assign n15134 = ~n15123 & ~n15133;
  assign n15135 = ~n7597 & ~n15134;
  assign n15136 = n7597 & ~n15041;
  assign n15137 = ~n15135 & ~n15136;
  assign n15138 = ~pi785 & ~n15137;
  assign n15139 = ~n7598 & ~n15041;
  assign n15140 = pi609 & n15135;
  assign n15141 = ~n15139 & ~n15140;
  assign n15142 = pi1155 & ~n15141;
  assign n15143 = ~n7610 & ~n15041;
  assign n15144 = ~pi609 & n15135;
  assign n15145 = ~n15143 & ~n15144;
  assign n15146 = ~pi1155 & ~n15145;
  assign n15147 = ~n15142 & ~n15146;
  assign n15148 = pi785 & ~n15147;
  assign n15149 = ~n15138 & ~n15148;
  assign n15150 = ~pi781 & ~n15149;
  assign n15151 = pi618 & n15149;
  assign n15152 = ~pi618 & n15041;
  assign n15153 = pi1154 & ~n15152;
  assign n15154 = ~n15151 & n15153;
  assign n15155 = ~pi618 & n15149;
  assign n15156 = pi618 & n15041;
  assign n15157 = ~pi1154 & ~n15156;
  assign n15158 = ~n15155 & n15157;
  assign n15159 = ~n15154 & ~n15158;
  assign n15160 = pi781 & ~n15159;
  assign n15161 = ~n15150 & ~n15160;
  assign n15162 = ~pi789 & ~n15161;
  assign n15163 = ~pi619 & n15161;
  assign n15164 = pi619 & n15041;
  assign n15165 = ~pi1159 & ~n15164;
  assign n15166 = ~n15163 & n15165;
  assign n15167 = pi619 & n15161;
  assign n15168 = ~pi619 & n15041;
  assign n15169 = pi1159 & ~n15168;
  assign n15170 = ~n15167 & n15169;
  assign n15171 = ~n15166 & ~n15170;
  assign n15172 = pi789 & ~n15171;
  assign n15173 = ~n15162 & ~n15172;
  assign n15174 = ~n8054 & n15173;
  assign n15175 = n8054 & n15041;
  assign n15176 = ~n15174 & ~n15175;
  assign n15177 = ~n7793 & ~n15176;
  assign n15178 = n7793 & n15041;
  assign n15179 = ~n15177 & ~n15178;
  assign n15180 = ~n7872 & n15179;
  assign n15181 = ~n15122 & ~n15180;
  assign n15182 = ~n15117 & n15181;
  assign n15183 = pi787 & ~n15182;
  assign n15184 = n12139 & n15173;
  assign n15185 = ~pi641 & ~n59519;
  assign n15186 = pi641 & ~n15041;
  assign n15187 = n7912 & ~n15186;
  assign n15188 = ~n15185 & n15187;
  assign n15189 = pi641 & ~n59519;
  assign n15190 = ~pi641 & ~n15041;
  assign n15191 = n7911 & ~n15190;
  assign n15192 = ~n15189 & n15191;
  assign n15193 = ~n15188 & ~n15192;
  assign n15194 = ~n15184 & n15193;
  assign n15195 = pi788 & ~n15194;
  assign n15196 = pi619 & ~n59518;
  assign n15197 = ~pi1159 & ~n15196;
  assign n15198 = ~pi648 & ~n15170;
  assign n15199 = ~n15197 & n15198;
  assign n15200 = ~pi619 & ~n59518;
  assign n15201 = pi1159 & ~n15200;
  assign n15202 = pi648 & ~n15166;
  assign n15203 = ~n15201 & n15202;
  assign n15204 = ~n15199 & ~n15203;
  assign n15205 = pi789 & ~n15204;
  assign n15206 = pi618 & n59517;
  assign n15207 = ~pi1154 & ~n15206;
  assign n15208 = ~pi627 & ~n15154;
  assign n15209 = ~n15207 & n15208;
  assign n15210 = n8233 & ~n15051;
  assign n15211 = ~pi179 & n8213;
  assign n15212 = pi179 & n8217;
  assign n15213 = ~pi38 & ~n15212;
  assign n15214 = ~pi179 & n59177;
  assign n15215 = pi179 & n7111;
  assign n15216 = pi39 & ~n15215;
  assign n15217 = ~n15214 & n15216;
  assign n15218 = ~pi179 & n7310;
  assign n15219 = pi179 & n7333;
  assign n15220 = ~pi39 & ~n15219;
  assign n15221 = ~pi39 & ~n15218;
  assign n15222 = ~n15219 & n15221;
  assign n15223 = ~n15218 & n15220;
  assign n15224 = ~n15217 & ~n59524;
  assign n15225 = ~pi38 & ~n15224;
  assign n15226 = ~n15211 & n15213;
  assign n15227 = ~n15210 & ~n59525;
  assign n15228 = pi741 & ~n15227;
  assign n15229 = pi179 & n9811;
  assign n15230 = ~pi179 & ~n59320;
  assign n15231 = ~pi741 & ~n15230;
  assign n15232 = ~n15229 & n15231;
  assign n15233 = ~pi724 & ~n15232;
  assign n15234 = ~n15228 & n15233;
  assign n15235 = pi724 & n15132;
  assign n15236 = n59132 & ~n15235;
  assign n15237 = ~n15234 & n15236;
  assign n15238 = ~n15123 & ~n15237;
  assign n15239 = pi625 & n15238;
  assign n15240 = ~pi625 & n15134;
  assign n15241 = pi1153 & ~n15240;
  assign n15242 = ~n15239 & n15241;
  assign n15243 = pi608 & ~n15060;
  assign n15244 = ~n15242 & n15243;
  assign n15245 = ~pi625 & n15238;
  assign n15246 = pi625 & n15134;
  assign n15247 = ~pi1153 & ~n15246;
  assign n15248 = ~n15245 & n15247;
  assign n15249 = ~pi608 & ~n15064;
  assign n15250 = ~n15248 & n15249;
  assign n15251 = ~n15244 & ~n15250;
  assign n15252 = pi778 & ~n15251;
  assign n15253 = ~pi778 & n15238;
  assign n15254 = ~pi778 & ~n15238;
  assign n15255 = pi778 & ~n15250;
  assign n15256 = ~n15244 & n15255;
  assign n15257 = ~n15254 & ~n15256;
  assign n15258 = ~n15252 & ~n15253;
  assign n15259 = ~pi609 & n59526;
  assign n15260 = pi609 & n15067;
  assign n15261 = ~pi1155 & ~n15260;
  assign n15262 = ~n15259 & n15261;
  assign n15263 = ~pi660 & ~n15142;
  assign n15264 = ~n15262 & n15263;
  assign n15265 = pi609 & n59526;
  assign n15266 = ~pi609 & n15067;
  assign n15267 = pi1155 & ~n15266;
  assign n15268 = ~n15265 & n15267;
  assign n15269 = pi660 & ~n15146;
  assign n15270 = ~n15268 & n15269;
  assign n15271 = ~n15264 & ~n15270;
  assign n15272 = pi785 & ~n15271;
  assign n15273 = ~pi785 & n59526;
  assign n15274 = ~n15272 & ~n15273;
  assign n15275 = pi618 & ~n15274;
  assign n15276 = ~pi618 & n59517;
  assign n15277 = pi1154 & ~n15276;
  assign n15278 = ~n15275 & n15277;
  assign n15279 = pi627 & ~n15158;
  assign n15280 = ~n15278 & n15279;
  assign n15281 = ~n15209 & ~n15280;
  assign n15282 = pi781 & ~n15281;
  assign n15283 = ~pi618 & n15208;
  assign n15284 = pi781 & ~n15283;
  assign n15285 = ~n15274 & ~n15284;
  assign n15286 = ~pi618 & ~n15274;
  assign n15287 = n15207 & ~n15286;
  assign n15288 = n15208 & ~n15287;
  assign n15289 = ~n15280 & ~n15288;
  assign n15290 = pi781 & ~n15289;
  assign n15291 = ~pi781 & ~n15274;
  assign n15292 = ~n15290 & ~n15291;
  assign n15293 = ~n15282 & ~n15285;
  assign n15294 = ~pi619 & n15198;
  assign n15295 = pi619 & n15202;
  assign n15296 = pi789 & ~n15295;
  assign n15297 = ~n15294 & n15296;
  assign n15298 = ~n59527 & ~n15297;
  assign n15299 = ~pi619 & ~n59527;
  assign n15300 = n15197 & ~n15299;
  assign n15301 = n15198 & ~n15300;
  assign n15302 = pi619 & ~n59527;
  assign n15303 = n15201 & ~n15302;
  assign n15304 = n15202 & ~n15303;
  assign n15305 = ~n15301 & ~n15304;
  assign n15306 = pi789 & ~n15305;
  assign n15307 = ~pi789 & ~n59527;
  assign n15308 = ~n15306 & ~n15307;
  assign n15309 = ~n15205 & ~n15298;
  assign n15310 = n59242 & ~n59528;
  assign n15311 = ~pi788 & n59528;
  assign n15312 = ~pi626 & n59528;
  assign n15313 = pi626 & ~n59519;
  assign n15314 = ~pi641 & ~n15313;
  assign n15315 = ~n15312 & n15314;
  assign n15316 = ~pi626 & ~n15173;
  assign n15317 = pi626 & ~n15041;
  assign n15318 = pi641 & ~n15317;
  assign n15319 = ~n15316 & n15318;
  assign n15320 = ~pi1158 & ~n15319;
  assign n15321 = ~n15315 & n15320;
  assign n15322 = pi626 & n59528;
  assign n15323 = ~pi626 & ~n59519;
  assign n15324 = pi641 & ~n15323;
  assign n15325 = ~n15322 & n15324;
  assign n15326 = pi626 & ~n15173;
  assign n15327 = ~pi626 & ~n15041;
  assign n15328 = ~pi641 & ~n15327;
  assign n15329 = ~n15326 & n15328;
  assign n15330 = pi1158 & ~n15329;
  assign n15331 = ~n15325 & n15330;
  assign n15332 = ~n15321 & ~n15331;
  assign n15333 = pi788 & ~n15332;
  assign n15334 = ~n15311 & ~n15333;
  assign n15335 = ~n15195 & ~n15310;
  assign n15336 = ~n11154 & n15176;
  assign n15337 = n7791 & ~n15100;
  assign n15338 = n7790 & ~n15104;
  assign n15339 = ~n15337 & ~n15338;
  assign n15340 = ~n15336 & n15339;
  assign n15341 = pi792 & ~n15340;
  assign n15342 = n59529 & ~n15341;
  assign n15343 = n59357 & n15340;
  assign n15344 = ~n8108 & ~n15343;
  assign n15345 = ~n15342 & n15344;
  assign n15346 = ~pi628 & n59529;
  assign n15347 = pi628 & ~n15176;
  assign n15348 = ~pi1156 & ~n15347;
  assign n15349 = ~n15346 & n15348;
  assign n15350 = ~pi629 & ~n15093;
  assign n15351 = ~n15349 & n15350;
  assign n15352 = pi628 & n59529;
  assign n15353 = ~pi628 & ~n15176;
  assign n15354 = pi1156 & ~n15353;
  assign n15355 = ~n15352 & n15354;
  assign n15356 = pi629 & ~n15097;
  assign n15357 = ~n15355 & n15356;
  assign n15358 = ~n15351 & ~n15357;
  assign n15359 = pi792 & ~n15358;
  assign n15360 = ~pi792 & n59529;
  assign n15361 = ~n15359 & ~n15360;
  assign n15362 = ~pi647 & ~n15361;
  assign n15363 = pi647 & ~n15179;
  assign n15364 = ~pi1157 & ~n15363;
  assign n15365 = ~n15362 & n15364;
  assign n15366 = pi1157 & ~n15115;
  assign n15367 = pi1157 & n15116;
  assign n15368 = ~n15114 & n15366;
  assign n15369 = ~pi630 & ~n59530;
  assign n15370 = ~n15365 & n15369;
  assign n15371 = pi647 & ~n15361;
  assign n15372 = ~pi647 & ~n15179;
  assign n15373 = pi1157 & ~n15372;
  assign n15374 = ~n15371 & n15373;
  assign n15375 = pi630 & ~n15121;
  assign n15376 = ~n15374 & n15375;
  assign n15377 = ~n15370 & ~n15376;
  assign n15378 = pi787 & ~n15377;
  assign n15379 = ~pi787 & ~n15361;
  assign n15380 = ~n15378 & ~n15379;
  assign n15381 = ~n15183 & ~n15345;
  assign n15382 = pi644 & ~n59531;
  assign n15383 = ~pi787 & ~n59522;
  assign n15384 = ~n15121 & ~n59530;
  assign n15385 = pi787 & ~n15384;
  assign n15386 = ~n15383 & ~n15385;
  assign n15387 = ~pi644 & n15386;
  assign n15388 = pi715 & ~n15387;
  assign n15389 = ~n15382 & n15388;
  assign n15390 = ~n7835 & ~n15179;
  assign n15391 = n7835 & n15041;
  assign n15392 = n7835 & ~n15041;
  assign n15393 = ~n7835 & n15179;
  assign n15394 = ~n15392 & ~n15393;
  assign n15395 = ~n15390 & ~n15391;
  assign n15396 = pi644 & n59532;
  assign n15397 = ~pi644 & n15041;
  assign n15398 = ~pi715 & ~n15397;
  assign n15399 = ~n15396 & n15398;
  assign n15400 = pi1160 & ~n15399;
  assign n15401 = ~n15389 & n15400;
  assign n15402 = ~pi644 & n59532;
  assign n15403 = pi644 & n15041;
  assign n15404 = pi715 & ~n15403;
  assign n15405 = ~n15402 & n15404;
  assign n15406 = ~pi1160 & ~n15405;
  assign n15407 = pi644 & n15386;
  assign n15408 = ~pi715 & ~n15407;
  assign n15409 = ~pi644 & ~n59531;
  assign n15410 = n15408 & ~n15409;
  assign n15411 = n15406 & ~n15410;
  assign n15412 = pi790 & ~n15411;
  assign n15413 = pi790 & ~n15401;
  assign n15414 = ~n15411 & n15413;
  assign n15415 = ~n15401 & n15412;
  assign n15416 = ~pi790 & n59531;
  assign n15417 = n58992 & ~n15416;
  assign n15418 = n15406 & ~n15408;
  assign n15419 = ~n15401 & ~n15418;
  assign n15420 = pi790 & ~n15419;
  assign n15421 = ~pi644 & n15406;
  assign n15422 = pi790 & ~n15421;
  assign n15423 = ~n59531 & ~n15422;
  assign n15424 = ~n15420 & ~n15423;
  assign n15425 = n58992 & ~n15424;
  assign n15426 = ~n59533 & n15417;
  assign n15427 = ~pi179 & ~n58992;
  assign n15428 = ~pi832 & ~n15427;
  assign n15429 = ~n59534 & n15428;
  assign po336 = ~n15040 & ~n15429;
  assign n15431 = ~pi180 & ~n2794;
  assign n15432 = ~pi753 & n6822;
  assign n15433 = ~n15431 & ~n15432;
  assign n15434 = ~n7875 & ~n15433;
  assign n15435 = ~pi785 & ~n15434;
  assign n15436 = n7610 & n15432;
  assign n15437 = n15434 & ~n15436;
  assign n15438 = pi1155 & ~n15437;
  assign n15439 = ~pi1155 & ~n15431;
  assign n15440 = ~n15436 & n15439;
  assign n15441 = ~n15438 & ~n15440;
  assign n15442 = pi785 & ~n15441;
  assign n15443 = ~n15435 & ~n15442;
  assign n15444 = ~pi781 & ~n15443;
  assign n15445 = ~n7890 & n15443;
  assign n15446 = pi1154 & ~n15445;
  assign n15447 = ~n7893 & n15443;
  assign n15448 = ~pi1154 & ~n15447;
  assign n15449 = ~n15446 & ~n15448;
  assign n15450 = pi781 & ~n15449;
  assign n15451 = ~n15444 & ~n15450;
  assign n15452 = ~pi789 & ~n15451;
  assign n15453 = ~n11882 & n15451;
  assign n15454 = pi1159 & ~n15453;
  assign n15455 = ~n11885 & n15451;
  assign n15456 = ~pi1159 & ~n15455;
  assign n15457 = ~n15454 & ~n15456;
  assign n15458 = pi789 & ~n15457;
  assign n15459 = ~n15452 & ~n15458;
  assign n15460 = ~n8054 & ~n15459;
  assign n15461 = n8054 & ~n15431;
  assign n15462 = ~n8054 & n15459;
  assign n15463 = n8054 & n15431;
  assign n15464 = ~n15462 & ~n15463;
  assign n15465 = ~n15460 & ~n15461;
  assign n15466 = ~n7793 & ~n59535;
  assign n15467 = n7793 & n15431;
  assign n15468 = ~n7872 & ~n15467;
  assign n15469 = ~n15466 & ~n15467;
  assign n15470 = ~n7872 & n15469;
  assign n15471 = ~n15466 & n15468;
  assign n15472 = ~pi702 & n7055;
  assign n15473 = ~n15431 & ~n15472;
  assign n15474 = ~pi778 & ~n15473;
  assign n15475 = ~pi625 & n15472;
  assign n15476 = ~n15473 & ~n15475;
  assign n15477 = pi1153 & ~n15476;
  assign n15478 = ~pi1153 & ~n15431;
  assign n15479 = ~n15475 & n15478;
  assign n15480 = pi778 & ~n15479;
  assign n15481 = ~n15477 & n15480;
  assign n15482 = ~n15474 & ~n15481;
  assign n15483 = ~n7949 & ~n15482;
  assign n15484 = ~n7951 & n15483;
  assign n15485 = ~n7953 & n15484;
  assign n15486 = ~n7955 & n15485;
  assign n15487 = ~n7967 & n15486;
  assign n15488 = pi647 & ~n15487;
  assign n15489 = ~pi647 & ~n15431;
  assign n15490 = ~n15488 & ~n15489;
  assign n15491 = n7832 & ~n15490;
  assign n15492 = ~pi647 & n15487;
  assign n15493 = pi647 & n15431;
  assign n15494 = ~pi1157 & ~n15493;
  assign n15495 = ~n15492 & n15494;
  assign n15496 = pi630 & n15495;
  assign n15497 = ~n15491 & ~n15496;
  assign n15498 = ~n59536 & n15497;
  assign n15499 = pi787 & ~n15498;
  assign n15500 = ~pi626 & ~n15459;
  assign n15501 = pi626 & ~n15431;
  assign n15502 = n7760 & ~n15501;
  assign n15503 = ~n15500 & n15502;
  assign n15504 = n7984 & n15485;
  assign n15505 = pi626 & ~n15459;
  assign n15506 = ~pi626 & ~n15431;
  assign n15507 = n7759 & ~n15506;
  assign n15508 = ~n15505 & n15507;
  assign n15509 = ~n15504 & ~n15508;
  assign n15510 = ~n15503 & ~n15504;
  assign n15511 = ~n15508 & n15510;
  assign n15512 = ~n15503 & n15509;
  assign n15513 = pi788 & ~n59537;
  assign n15514 = ~n6701 & ~n15473;
  assign n15515 = pi625 & n15514;
  assign n15516 = n15433 & ~n15514;
  assign n15517 = ~n15515 & ~n15516;
  assign n15518 = n15478 & ~n15517;
  assign n15519 = ~pi608 & ~n15477;
  assign n15520 = ~n15518 & n15519;
  assign n15521 = pi1153 & n15433;
  assign n15522 = ~n15515 & n15521;
  assign n15523 = pi608 & ~n15479;
  assign n15524 = ~n15522 & n15523;
  assign n15525 = ~n15520 & ~n15524;
  assign n15526 = pi778 & ~n15525;
  assign n15527 = ~pi778 & ~n15516;
  assign n15528 = ~n15526 & ~n15527;
  assign n15529 = ~pi609 & ~n15528;
  assign n15530 = pi609 & ~n15482;
  assign n15531 = ~pi1155 & ~n15530;
  assign n15532 = ~n15529 & n15531;
  assign n15533 = ~pi660 & ~n15438;
  assign n15534 = ~n15532 & n15533;
  assign n15535 = pi609 & ~n15528;
  assign n15536 = ~pi609 & ~n15482;
  assign n15537 = pi1155 & ~n15536;
  assign n15538 = ~n15535 & n15537;
  assign n15539 = pi660 & ~n15440;
  assign n15540 = ~n15538 & n15539;
  assign n15541 = ~n15534 & ~n15540;
  assign n15542 = pi785 & ~n15541;
  assign n15543 = ~pi785 & ~n15528;
  assign n15544 = ~n15542 & ~n15543;
  assign n15545 = ~pi618 & ~n15544;
  assign n15546 = pi618 & n15483;
  assign n15547 = ~pi1154 & ~n15546;
  assign n15548 = ~n15545 & n15547;
  assign n15549 = ~pi627 & ~n15446;
  assign n15550 = ~n15548 & n15549;
  assign n15551 = pi618 & ~n15544;
  assign n15552 = ~pi618 & n15483;
  assign n15553 = pi1154 & ~n15552;
  assign n15554 = ~n15551 & n15553;
  assign n15555 = pi627 & ~n15448;
  assign n15556 = ~n15554 & n15555;
  assign n15557 = ~n15550 & ~n15556;
  assign n15558 = pi781 & ~n15557;
  assign n15559 = ~pi781 & ~n15544;
  assign n15560 = ~n15558 & ~n15559;
  assign n15561 = pi619 & ~n15560;
  assign n15562 = ~pi619 & n15484;
  assign n15563 = pi1159 & ~n15562;
  assign n15564 = ~n15561 & n15563;
  assign n15565 = pi648 & ~n15456;
  assign n15566 = ~n15564 & n15565;
  assign n15567 = ~pi619 & ~n15560;
  assign n15568 = pi619 & n15484;
  assign n15569 = ~pi1159 & ~n15568;
  assign n15570 = ~n15567 & n15569;
  assign n15571 = ~pi648 & ~n15454;
  assign n15572 = ~n15570 & n15571;
  assign n15573 = pi789 & ~n15572;
  assign n15574 = pi789 & ~n15566;
  assign n15575 = ~n15572 & n15574;
  assign n15576 = ~n15566 & n15573;
  assign n15577 = ~pi789 & n15560;
  assign n15578 = n59242 & ~n15577;
  assign n15579 = ~n59538 & n15578;
  assign n15580 = ~n15513 & ~n15579;
  assign n15581 = ~n59357 & ~n15580;
  assign n15582 = n7957 & ~n59535;
  assign n15583 = n8065 & n15486;
  assign n15584 = pi629 & ~n15583;
  assign n15585 = ~n15582 & n15584;
  assign n15586 = n7958 & ~n59535;
  assign n15587 = n8074 & n15486;
  assign n15588 = ~pi629 & ~n15587;
  assign n15589 = ~n15586 & n15588;
  assign n15590 = pi792 & ~n15589;
  assign n15591 = ~n15586 & ~n15587;
  assign n15592 = ~pi629 & ~n15591;
  assign n15593 = ~n15582 & ~n15583;
  assign n15594 = pi629 & ~n15593;
  assign n15595 = ~n15592 & ~n15594;
  assign n15596 = pi792 & ~n15595;
  assign n15597 = pi792 & ~n15585;
  assign n15598 = ~n15589 & n15597;
  assign n15599 = ~n15585 & n15590;
  assign n15600 = ~n8108 & ~n59539;
  assign n15601 = ~n15581 & n15600;
  assign n15602 = ~n15499 & ~n15601;
  assign n15603 = pi644 & n15602;
  assign n15604 = ~pi787 & ~n15487;
  assign n15605 = pi1157 & ~n15490;
  assign n15606 = ~n15495 & ~n15605;
  assign n15607 = pi787 & ~n15606;
  assign n15608 = ~n15604 & ~n15607;
  assign n15609 = ~pi644 & n15608;
  assign n15610 = pi715 & ~n15609;
  assign n15611 = ~n15603 & n15610;
  assign n15612 = ~n11491 & n15431;
  assign n15613 = ~n7835 & n15466;
  assign n15614 = ~n7835 & ~n15469;
  assign n15615 = n7835 & n15431;
  assign n15616 = ~n15614 & ~n15615;
  assign n15617 = ~n15612 & ~n15613;
  assign n15618 = pi644 & ~n59540;
  assign n15619 = ~pi644 & n15431;
  assign n15620 = ~pi715 & ~n15619;
  assign n15621 = ~n15618 & n15620;
  assign n15622 = pi1160 & ~n15621;
  assign n15623 = ~n15611 & n15622;
  assign n15624 = ~pi644 & n15602;
  assign n15625 = pi644 & n15608;
  assign n15626 = ~pi715 & ~n15625;
  assign n15627 = ~n15624 & n15626;
  assign n15628 = ~pi644 & ~n59540;
  assign n15629 = pi644 & n15431;
  assign n15630 = pi715 & ~n15629;
  assign n15631 = ~n15628 & n15630;
  assign n15632 = ~pi1160 & ~n15631;
  assign n15633 = ~n15627 & n15632;
  assign n15634 = ~n15623 & ~n15633;
  assign n15635 = pi790 & ~n15634;
  assign n15636 = ~pi790 & n15602;
  assign n15637 = pi832 & ~n15636;
  assign n15638 = ~n15635 & n15637;
  assign n15639 = ~pi180 & ~n7560;
  assign n15640 = n59231 & ~n15639;
  assign n15641 = ~pi702 & n59132;
  assign n15642 = n15639 & ~n15641;
  assign n15643 = pi180 & n59251;
  assign n15644 = ~pi38 & ~n15643;
  assign n15645 = n59132 & ~n15644;
  assign n15646 = ~pi180 & n8249;
  assign n15647 = ~n15645 & ~n15646;
  assign n15648 = ~pi180 & ~n6863;
  assign n15649 = n7547 & ~n15648;
  assign n15650 = ~pi702 & ~n15649;
  assign n15651 = ~n15647 & n15650;
  assign n15652 = ~n15642 & ~n15651;
  assign n15653 = ~pi778 & n15652;
  assign n15654 = pi625 & ~n15652;
  assign n15655 = ~pi625 & n15639;
  assign n15656 = pi1153 & ~n15655;
  assign n15657 = ~n15654 & n15656;
  assign n15658 = ~pi625 & ~n15652;
  assign n15659 = pi625 & n15639;
  assign n15660 = ~pi1153 & ~n15659;
  assign n15661 = ~n15658 & n15660;
  assign n15662 = ~n15657 & ~n15661;
  assign n15663 = pi778 & ~n15662;
  assign n15664 = ~n15653 & ~n15663;
  assign n15665 = ~n59229 & n15664;
  assign n15666 = n59229 & n15639;
  assign n15667 = n59229 & ~n15639;
  assign n15668 = ~n59229 & ~n15664;
  assign n15669 = ~n15667 & ~n15668;
  assign n15670 = ~n15665 & ~n15666;
  assign n15671 = ~n59231 & ~n59541;
  assign n15672 = ~n59231 & n59541;
  assign n15673 = n59231 & n15639;
  assign n15674 = ~n15672 & ~n15673;
  assign n15675 = ~n15640 & ~n15671;
  assign n15676 = ~n7716 & ~n59542;
  assign n15677 = n7716 & n15639;
  assign n15678 = n7716 & ~n15639;
  assign n15679 = ~n7716 & n59542;
  assign n15680 = ~n15678 & ~n15679;
  assign n15681 = ~n15676 & ~n15677;
  assign n15682 = ~n7762 & n59543;
  assign n15683 = n7762 & n15639;
  assign n15684 = ~n15682 & ~n15683;
  assign n15685 = ~pi792 & n15684;
  assign n15686 = pi628 & ~n15684;
  assign n15687 = ~pi628 & n15639;
  assign n15688 = pi1156 & ~n15687;
  assign n15689 = ~n15686 & n15688;
  assign n15690 = ~pi628 & ~n15684;
  assign n15691 = pi628 & n15639;
  assign n15692 = ~pi1156 & ~n15691;
  assign n15693 = ~n15690 & n15692;
  assign n15694 = ~n15689 & ~n15693;
  assign n15695 = pi792 & ~n15694;
  assign n15696 = ~n15685 & ~n15695;
  assign n15697 = pi647 & n15696;
  assign n15698 = ~pi647 & n15639;
  assign n15699 = pi647 & ~n15696;
  assign n15700 = ~pi647 & ~n15639;
  assign n15701 = ~n15699 & ~n15700;
  assign n15702 = ~n15697 & ~n15698;
  assign n15703 = pi1157 & ~n59544;
  assign n15704 = ~pi647 & n15696;
  assign n15705 = pi647 & n15639;
  assign n15706 = ~pi1157 & ~n15705;
  assign n15707 = ~n15704 & n15706;
  assign n15708 = ~pi647 & ~n15696;
  assign n15709 = pi647 & ~n15639;
  assign n15710 = ~n15708 & ~n15709;
  assign n15711 = ~pi1157 & n15710;
  assign n15712 = pi1157 & n59544;
  assign n15713 = ~n15711 & ~n15712;
  assign n15714 = ~n15703 & ~n15707;
  assign n15715 = pi787 & n59545;
  assign n15716 = ~pi787 & ~n15696;
  assign n15717 = pi787 & ~n59545;
  assign n15718 = ~pi787 & n15696;
  assign n15719 = ~n15717 & ~n15718;
  assign n15720 = ~n15715 & ~n15716;
  assign n15721 = ~pi644 & ~n59546;
  assign n15722 = pi715 & ~n15721;
  assign n15723 = pi180 & ~n59132;
  assign n15724 = pi753 & n6654;
  assign n15725 = pi180 & n6853;
  assign n15726 = ~n15724 & ~n15725;
  assign n15727 = pi39 & ~n15726;
  assign n15728 = ~pi180 & ~pi753;
  assign n15729 = n59164 & n15728;
  assign n15730 = pi180 & pi753;
  assign n15731 = pi753 & n59147;
  assign n15732 = pi180 & ~n6798;
  assign n15733 = ~n15731 & ~n15732;
  assign n15734 = ~pi39 & ~n15733;
  assign n15735 = ~n15730 & ~n15734;
  assign n15736 = ~n15729 & n15735;
  assign n15737 = ~n15727 & n15736;
  assign n15738 = ~pi38 & ~n15737;
  assign n15739 = ~pi753 & n6865;
  assign n15740 = pi38 & ~n15648;
  assign n15741 = ~n15739 & n15740;
  assign n15742 = ~n15738 & ~n15741;
  assign n15743 = n59132 & ~n15742;
  assign n15744 = ~n15723 & ~n15743;
  assign n15745 = ~n7597 & ~n15744;
  assign n15746 = n7597 & ~n15639;
  assign n15747 = ~n15745 & ~n15746;
  assign n15748 = ~pi785 & ~n15747;
  assign n15749 = ~n7598 & ~n15639;
  assign n15750 = pi609 & n15745;
  assign n15751 = ~n15749 & ~n15750;
  assign n15752 = pi1155 & ~n15751;
  assign n15753 = ~n7610 & ~n15639;
  assign n15754 = ~pi609 & n15745;
  assign n15755 = ~n15753 & ~n15754;
  assign n15756 = ~pi1155 & ~n15755;
  assign n15757 = ~n15752 & ~n15756;
  assign n15758 = pi785 & ~n15757;
  assign n15759 = ~n15748 & ~n15758;
  assign n15760 = ~pi781 & ~n15759;
  assign n15761 = pi618 & n15759;
  assign n15762 = ~pi618 & n15639;
  assign n15763 = pi1154 & ~n15762;
  assign n15764 = ~n15761 & n15763;
  assign n15765 = ~pi618 & n15759;
  assign n15766 = pi618 & n15639;
  assign n15767 = ~pi1154 & ~n15766;
  assign n15768 = ~n15765 & n15767;
  assign n15769 = ~n15764 & ~n15768;
  assign n15770 = pi781 & ~n15769;
  assign n15771 = ~n15760 & ~n15770;
  assign n15772 = ~pi789 & ~n15771;
  assign n15773 = pi619 & n15771;
  assign n15774 = ~pi619 & n15639;
  assign n15775 = pi1159 & ~n15774;
  assign n15776 = ~n15773 & n15775;
  assign n15777 = ~pi619 & n15771;
  assign n15778 = pi619 & n15639;
  assign n15779 = ~pi1159 & ~n15778;
  assign n15780 = ~n15777 & n15779;
  assign n15781 = ~n15776 & ~n15780;
  assign n15782 = pi789 & ~n15781;
  assign n15783 = ~n15772 & ~n15782;
  assign n15784 = ~n8054 & n15783;
  assign n15785 = n8054 & n15639;
  assign n15786 = ~n15784 & ~n15785;
  assign n15787 = ~n7793 & ~n15786;
  assign n15788 = n7793 & n15639;
  assign n15789 = ~n15787 & ~n15788;
  assign n15790 = ~n7835 & ~n15789;
  assign n15791 = n7835 & n15639;
  assign n15792 = n7835 & ~n15639;
  assign n15793 = ~n7835 & n15789;
  assign n15794 = ~n15792 & ~n15793;
  assign n15795 = ~n15790 & ~n15791;
  assign n15796 = pi644 & n59547;
  assign n15797 = ~pi644 & n15639;
  assign n15798 = ~pi715 & ~n15797;
  assign n15799 = ~n15796 & n15798;
  assign n15800 = pi1160 & ~n15799;
  assign n15801 = ~n15722 & n15800;
  assign n15802 = pi644 & ~n59546;
  assign n15803 = ~pi715 & ~n15802;
  assign n15804 = ~pi644 & n59547;
  assign n15805 = pi644 & n15639;
  assign n15806 = pi715 & ~n15805;
  assign n15807 = ~n15804 & n15806;
  assign n15808 = ~pi1160 & ~n15807;
  assign n15809 = ~n15803 & n15808;
  assign n15810 = ~n15801 & ~n15809;
  assign n15811 = pi790 & ~n15810;
  assign n15812 = ~pi644 & n15808;
  assign n15813 = pi644 & n15800;
  assign n15814 = pi790 & ~n15813;
  assign n15815 = pi790 & ~n15812;
  assign n15816 = ~n15813 & n15815;
  assign n15817 = ~n15812 & n15814;
  assign n15818 = ~n7872 & n15789;
  assign n15819 = n7832 & ~n59544;
  assign n15820 = n7833 & ~n15710;
  assign n15821 = pi630 & n15707;
  assign n15822 = ~n15819 & ~n59549;
  assign n15823 = ~n15818 & n15822;
  assign n15824 = pi787 & ~n15823;
  assign n15825 = ~n11154 & n15786;
  assign n15826 = ~pi629 & n15689;
  assign n15827 = pi629 & n15693;
  assign n15828 = ~n15826 & ~n15827;
  assign n15829 = ~n15825 & n15828;
  assign n15830 = pi792 & ~n15829;
  assign n15831 = pi702 & n15742;
  assign n15832 = ~pi180 & n59177;
  assign n15833 = pi180 & n7111;
  assign n15834 = pi753 & ~n15833;
  assign n15835 = ~n15832 & n15834;
  assign n15836 = pi180 & n7188;
  assign n15837 = ~pi180 & ~n59203;
  assign n15838 = ~pi753 & ~n15837;
  assign n15839 = ~n15836 & n15838;
  assign n15840 = pi39 & ~n15839;
  assign n15841 = ~n15835 & n15840;
  assign n15842 = pi180 & n7333;
  assign n15843 = ~pi180 & n7310;
  assign n15844 = pi753 & ~n15843;
  assign n15845 = ~n15842 & n15844;
  assign n15846 = ~pi180 & ~n7339;
  assign n15847 = pi180 & ~n7347;
  assign n15848 = ~pi753 & ~n15847;
  assign n15849 = ~n15846 & n15848;
  assign n15850 = ~pi39 & ~n15849;
  assign n15851 = pi180 & ~n7333;
  assign n15852 = ~pi180 & ~n7310;
  assign n15853 = pi753 & ~n15852;
  assign n15854 = pi753 & ~n15851;
  assign n15855 = ~n15852 & n15854;
  assign n15856 = ~n15851 & n15853;
  assign n15857 = ~pi180 & n7339;
  assign n15858 = pi180 & n7347;
  assign n15859 = ~pi753 & ~n15858;
  assign n15860 = ~n15857 & n15859;
  assign n15861 = ~n59550 & ~n15860;
  assign n15862 = ~pi39 & ~n15861;
  assign n15863 = ~n15845 & n15850;
  assign n15864 = ~pi38 & ~n59551;
  assign n15865 = ~n15841 & n15864;
  assign n15866 = ~pi753 & ~n7222;
  assign n15867 = n9794 & ~n15866;
  assign n15868 = ~pi180 & ~n15867;
  assign n15869 = ~n7056 & ~n15432;
  assign n15870 = pi180 & ~n15869;
  assign n15871 = n59171 & n15870;
  assign n15872 = pi38 & ~n15871;
  assign n15873 = ~n15868 & n15872;
  assign n15874 = ~pi702 & ~n15873;
  assign n15875 = ~n15865 & n15874;
  assign n15876 = n59132 & ~n15875;
  assign n15877 = ~n15831 & n15876;
  assign n15878 = ~n15723 & ~n15877;
  assign n15879 = ~pi625 & n15878;
  assign n15880 = pi625 & n15744;
  assign n15881 = ~pi1153 & ~n15880;
  assign n15882 = ~n15879 & n15881;
  assign n15883 = ~pi608 & ~n15657;
  assign n15884 = ~n15882 & n15883;
  assign n15885 = pi625 & n15878;
  assign n15886 = ~pi625 & n15744;
  assign n15887 = pi1153 & ~n15886;
  assign n15888 = ~n15885 & n15887;
  assign n15889 = pi608 & ~n15661;
  assign n15890 = ~n15888 & n15889;
  assign n15891 = ~n15884 & ~n15890;
  assign n15892 = pi778 & ~n15891;
  assign n15893 = ~pi778 & n15878;
  assign n15894 = ~n15892 & ~n15893;
  assign n15895 = ~pi609 & ~n15894;
  assign n15896 = pi609 & n15664;
  assign n15897 = ~pi1155 & ~n15896;
  assign n15898 = ~n15895 & n15897;
  assign n15899 = ~pi660 & ~n15752;
  assign n15900 = ~n15898 & n15899;
  assign n15901 = pi609 & ~n15894;
  assign n15902 = ~pi609 & n15664;
  assign n15903 = pi1155 & ~n15902;
  assign n15904 = ~n15901 & n15903;
  assign n15905 = pi660 & ~n15756;
  assign n15906 = ~n15904 & n15905;
  assign n15907 = ~n15900 & ~n15906;
  assign n15908 = pi785 & ~n15907;
  assign n15909 = ~pi785 & ~n15894;
  assign n15910 = ~n15908 & ~n15909;
  assign n15911 = ~pi618 & ~n15910;
  assign n15912 = pi618 & n59541;
  assign n15913 = ~pi1154 & ~n15912;
  assign n15914 = ~n15911 & n15913;
  assign n15915 = ~pi627 & ~n15764;
  assign n15916 = ~n15914 & n15915;
  assign n15917 = pi618 & ~n15910;
  assign n15918 = ~pi618 & n59541;
  assign n15919 = pi1154 & ~n15918;
  assign n15920 = ~n15917 & n15919;
  assign n15921 = pi627 & ~n15768;
  assign n15922 = ~n15920 & n15921;
  assign n15923 = ~n15916 & ~n15922;
  assign n15924 = pi781 & ~n15923;
  assign n15925 = ~pi781 & ~n15910;
  assign n15926 = ~n15924 & ~n15925;
  assign n15927 = pi619 & ~n15926;
  assign n15928 = ~pi619 & ~n59542;
  assign n15929 = pi1159 & ~n15928;
  assign n15930 = ~n15927 & n15929;
  assign n15931 = pi648 & ~n15780;
  assign n15932 = ~n15930 & n15931;
  assign n15933 = ~pi619 & ~n15926;
  assign n15934 = pi619 & ~n59542;
  assign n15935 = ~pi1159 & ~n15934;
  assign n15936 = ~n15933 & n15935;
  assign n15937 = ~pi648 & ~n15776;
  assign n15938 = ~n15936 & n15937;
  assign n15939 = pi789 & ~n15938;
  assign n15940 = pi789 & ~n15932;
  assign n15941 = ~n15938 & n15940;
  assign n15942 = ~n15932 & n15939;
  assign n15943 = ~pi789 & n15926;
  assign n15944 = n59242 & ~n15943;
  assign n15945 = ~n59552 & n15944;
  assign n15946 = ~pi626 & ~n15783;
  assign n15947 = pi626 & ~n15639;
  assign n15948 = n7760 & ~n15947;
  assign n15949 = ~n15946 & n15948;
  assign n15950 = n7984 & n59543;
  assign n15951 = pi626 & ~n15783;
  assign n15952 = ~pi626 & ~n15639;
  assign n15953 = n7759 & ~n15952;
  assign n15954 = ~n15951 & n15953;
  assign n15955 = ~n15950 & ~n15954;
  assign n15956 = ~n15949 & ~n15950;
  assign n15957 = ~n15954 & n15956;
  assign n15958 = ~n15949 & n15955;
  assign n15959 = pi788 & ~n59553;
  assign n15960 = ~n59357 & ~n15959;
  assign n15961 = ~n15945 & n15960;
  assign n15962 = ~n15830 & ~n15961;
  assign n15963 = ~n8108 & ~n15962;
  assign n15964 = ~n15824 & ~n15963;
  assign n15965 = ~n59548 & n15964;
  assign n15966 = ~n15811 & ~n15965;
  assign n15967 = n58992 & ~n15966;
  assign n15968 = ~pi180 & ~n58992;
  assign n15969 = ~pi832 & ~n15968;
  assign n15970 = ~n15967 & n15969;
  assign po337 = ~n15638 & ~n15970;
  assign n15972 = ~pi181 & ~n2794;
  assign n15973 = ~pi754 & n6822;
  assign n15974 = ~n15972 & ~n15973;
  assign n15975 = ~n7875 & ~n15974;
  assign n15976 = ~pi785 & ~n15975;
  assign n15977 = n7610 & n15973;
  assign n15978 = n15975 & ~n15977;
  assign n15979 = pi1155 & ~n15978;
  assign n15980 = ~pi1155 & ~n15972;
  assign n15981 = ~n15977 & n15980;
  assign n15982 = ~n15979 & ~n15981;
  assign n15983 = pi785 & ~n15982;
  assign n15984 = ~n15976 & ~n15983;
  assign n15985 = ~pi781 & ~n15984;
  assign n15986 = ~n7890 & n15984;
  assign n15987 = pi1154 & ~n15986;
  assign n15988 = ~n7893 & n15984;
  assign n15989 = ~pi1154 & ~n15988;
  assign n15990 = ~n15987 & ~n15989;
  assign n15991 = pi781 & ~n15990;
  assign n15992 = ~n15985 & ~n15991;
  assign n15993 = ~pi789 & ~n15992;
  assign n15994 = ~n11882 & n15992;
  assign n15995 = pi1159 & ~n15994;
  assign n15996 = ~n11885 & n15992;
  assign n15997 = ~pi1159 & ~n15996;
  assign n15998 = ~n15995 & ~n15997;
  assign n15999 = pi789 & ~n15998;
  assign n16000 = ~n15993 & ~n15999;
  assign n16001 = ~n8054 & ~n16000;
  assign n16002 = n8054 & ~n15972;
  assign n16003 = ~n8054 & n16000;
  assign n16004 = n8054 & n15972;
  assign n16005 = ~n16003 & ~n16004;
  assign n16006 = ~n16001 & ~n16002;
  assign n16007 = ~n7793 & ~n59554;
  assign n16008 = n7793 & n15972;
  assign n16009 = ~n7872 & ~n16008;
  assign n16010 = ~n16007 & ~n16008;
  assign n16011 = ~n7872 & n16010;
  assign n16012 = ~n16007 & n16009;
  assign n16013 = ~pi709 & n7055;
  assign n16014 = ~n15972 & ~n16013;
  assign n16015 = ~pi778 & ~n16014;
  assign n16016 = ~pi625 & n16013;
  assign n16017 = ~n16014 & ~n16016;
  assign n16018 = pi1153 & ~n16017;
  assign n16019 = ~pi1153 & ~n15972;
  assign n16020 = ~n16016 & n16019;
  assign n16021 = pi778 & ~n16020;
  assign n16022 = ~n16018 & n16021;
  assign n16023 = ~n16015 & ~n16022;
  assign n16024 = ~n7949 & ~n16023;
  assign n16025 = ~n7951 & n16024;
  assign n16026 = ~n7953 & n16025;
  assign n16027 = ~n7955 & n16026;
  assign n16028 = ~n7967 & n16027;
  assign n16029 = pi647 & ~n16028;
  assign n16030 = ~pi647 & ~n15972;
  assign n16031 = ~n16029 & ~n16030;
  assign n16032 = n7832 & ~n16031;
  assign n16033 = ~pi647 & n16028;
  assign n16034 = pi647 & n15972;
  assign n16035 = ~pi1157 & ~n16034;
  assign n16036 = ~n16033 & n16035;
  assign n16037 = pi630 & n16036;
  assign n16038 = ~n16032 & ~n16037;
  assign n16039 = ~n59555 & n16038;
  assign n16040 = pi787 & ~n16039;
  assign n16041 = ~pi626 & ~n16000;
  assign n16042 = pi626 & ~n15972;
  assign n16043 = n7760 & ~n16042;
  assign n16044 = ~n16041 & n16043;
  assign n16045 = n7984 & n16026;
  assign n16046 = pi626 & ~n16000;
  assign n16047 = ~pi626 & ~n15972;
  assign n16048 = n7759 & ~n16047;
  assign n16049 = ~n16046 & n16048;
  assign n16050 = ~n16045 & ~n16049;
  assign n16051 = ~n16044 & ~n16045;
  assign n16052 = ~n16049 & n16051;
  assign n16053 = ~n16044 & n16050;
  assign n16054 = pi788 & ~n59556;
  assign n16055 = ~n6701 & ~n16014;
  assign n16056 = pi625 & n16055;
  assign n16057 = n15974 & ~n16055;
  assign n16058 = ~n16056 & ~n16057;
  assign n16059 = n16019 & ~n16058;
  assign n16060 = ~pi608 & ~n16018;
  assign n16061 = ~n16059 & n16060;
  assign n16062 = pi1153 & n15974;
  assign n16063 = ~n16056 & n16062;
  assign n16064 = pi608 & ~n16020;
  assign n16065 = ~n16063 & n16064;
  assign n16066 = ~n16061 & ~n16065;
  assign n16067 = pi778 & ~n16066;
  assign n16068 = ~pi778 & ~n16057;
  assign n16069 = ~n16067 & ~n16068;
  assign n16070 = ~pi609 & ~n16069;
  assign n16071 = pi609 & ~n16023;
  assign n16072 = ~pi1155 & ~n16071;
  assign n16073 = ~n16070 & n16072;
  assign n16074 = ~pi660 & ~n15979;
  assign n16075 = ~n16073 & n16074;
  assign n16076 = pi609 & ~n16069;
  assign n16077 = ~pi609 & ~n16023;
  assign n16078 = pi1155 & ~n16077;
  assign n16079 = ~n16076 & n16078;
  assign n16080 = pi660 & ~n15981;
  assign n16081 = ~n16079 & n16080;
  assign n16082 = ~n16075 & ~n16081;
  assign n16083 = pi785 & ~n16082;
  assign n16084 = ~pi785 & ~n16069;
  assign n16085 = ~n16083 & ~n16084;
  assign n16086 = ~pi618 & ~n16085;
  assign n16087 = pi618 & n16024;
  assign n16088 = ~pi1154 & ~n16087;
  assign n16089 = ~n16086 & n16088;
  assign n16090 = ~pi627 & ~n15987;
  assign n16091 = ~n16089 & n16090;
  assign n16092 = pi618 & ~n16085;
  assign n16093 = ~pi618 & n16024;
  assign n16094 = pi1154 & ~n16093;
  assign n16095 = ~n16092 & n16094;
  assign n16096 = pi627 & ~n15989;
  assign n16097 = ~n16095 & n16096;
  assign n16098 = ~n16091 & ~n16097;
  assign n16099 = pi781 & ~n16098;
  assign n16100 = ~pi781 & ~n16085;
  assign n16101 = ~n16099 & ~n16100;
  assign n16102 = pi619 & ~n16101;
  assign n16103 = ~pi619 & n16025;
  assign n16104 = pi1159 & ~n16103;
  assign n16105 = ~n16102 & n16104;
  assign n16106 = pi648 & ~n15997;
  assign n16107 = ~n16105 & n16106;
  assign n16108 = ~pi619 & ~n16101;
  assign n16109 = pi619 & n16025;
  assign n16110 = ~pi1159 & ~n16109;
  assign n16111 = ~n16108 & n16110;
  assign n16112 = ~pi648 & ~n15995;
  assign n16113 = ~n16111 & n16112;
  assign n16114 = pi789 & ~n16113;
  assign n16115 = pi789 & ~n16107;
  assign n16116 = ~n16113 & n16115;
  assign n16117 = ~n16107 & n16114;
  assign n16118 = ~pi789 & n16101;
  assign n16119 = n59242 & ~n16118;
  assign n16120 = ~n59557 & n16119;
  assign n16121 = ~n16054 & ~n16120;
  assign n16122 = ~n59357 & ~n16121;
  assign n16123 = n7957 & ~n59554;
  assign n16124 = n8065 & n16027;
  assign n16125 = pi629 & ~n16124;
  assign n16126 = ~n16123 & n16125;
  assign n16127 = n7958 & ~n59554;
  assign n16128 = n8074 & n16027;
  assign n16129 = ~pi629 & ~n16128;
  assign n16130 = ~n16127 & n16129;
  assign n16131 = pi792 & ~n16130;
  assign n16132 = ~n16127 & ~n16128;
  assign n16133 = ~pi629 & ~n16132;
  assign n16134 = ~n16123 & ~n16124;
  assign n16135 = pi629 & ~n16134;
  assign n16136 = ~n16133 & ~n16135;
  assign n16137 = pi792 & ~n16136;
  assign n16138 = pi792 & ~n16126;
  assign n16139 = ~n16130 & n16138;
  assign n16140 = ~n16126 & n16131;
  assign n16141 = ~n8108 & ~n59558;
  assign n16142 = ~n16122 & n16141;
  assign n16143 = ~n16040 & ~n16142;
  assign n16144 = pi644 & n16143;
  assign n16145 = ~pi787 & ~n16028;
  assign n16146 = pi1157 & ~n16031;
  assign n16147 = ~n16036 & ~n16146;
  assign n16148 = pi787 & ~n16147;
  assign n16149 = ~n16145 & ~n16148;
  assign n16150 = ~pi644 & n16149;
  assign n16151 = pi715 & ~n16150;
  assign n16152 = ~n16144 & n16151;
  assign n16153 = ~n11491 & n15972;
  assign n16154 = ~n7835 & n16007;
  assign n16155 = ~n7835 & ~n16010;
  assign n16156 = n7835 & n15972;
  assign n16157 = ~n16155 & ~n16156;
  assign n16158 = ~n16153 & ~n16154;
  assign n16159 = pi644 & ~n59559;
  assign n16160 = ~pi644 & n15972;
  assign n16161 = ~pi715 & ~n16160;
  assign n16162 = ~n16159 & n16161;
  assign n16163 = pi1160 & ~n16162;
  assign n16164 = ~n16152 & n16163;
  assign n16165 = ~pi644 & n16143;
  assign n16166 = pi644 & n16149;
  assign n16167 = ~pi715 & ~n16166;
  assign n16168 = ~n16165 & n16167;
  assign n16169 = ~pi644 & ~n59559;
  assign n16170 = pi644 & n15972;
  assign n16171 = pi715 & ~n16170;
  assign n16172 = ~n16169 & n16171;
  assign n16173 = ~pi1160 & ~n16172;
  assign n16174 = ~n16168 & n16173;
  assign n16175 = ~n16164 & ~n16174;
  assign n16176 = pi790 & ~n16175;
  assign n16177 = ~pi790 & n16143;
  assign n16178 = pi832 & ~n16177;
  assign n16179 = ~n16176 & n16178;
  assign n16180 = ~pi181 & ~n7560;
  assign n16181 = n59231 & ~n16180;
  assign n16182 = ~pi709 & n59132;
  assign n16183 = n16180 & ~n16182;
  assign n16184 = pi181 & n59251;
  assign n16185 = ~pi38 & ~n16184;
  assign n16186 = n59132 & ~n16185;
  assign n16187 = ~pi181 & n8249;
  assign n16188 = ~n16186 & ~n16187;
  assign n16189 = ~pi181 & ~n6863;
  assign n16190 = n7547 & ~n16189;
  assign n16191 = ~pi709 & ~n16190;
  assign n16192 = ~n16188 & n16191;
  assign n16193 = ~n16183 & ~n16192;
  assign n16194 = ~pi778 & n16193;
  assign n16195 = pi625 & ~n16193;
  assign n16196 = ~pi625 & n16180;
  assign n16197 = pi1153 & ~n16196;
  assign n16198 = ~n16195 & n16197;
  assign n16199 = ~pi625 & ~n16193;
  assign n16200 = pi625 & n16180;
  assign n16201 = ~pi1153 & ~n16200;
  assign n16202 = ~n16199 & n16201;
  assign n16203 = ~n16198 & ~n16202;
  assign n16204 = pi778 & ~n16203;
  assign n16205 = ~n16194 & ~n16204;
  assign n16206 = ~n59229 & n16205;
  assign n16207 = n59229 & n16180;
  assign n16208 = n59229 & ~n16180;
  assign n16209 = ~n59229 & ~n16205;
  assign n16210 = ~n16208 & ~n16209;
  assign n16211 = ~n16206 & ~n16207;
  assign n16212 = ~n59231 & ~n59560;
  assign n16213 = ~n59231 & n59560;
  assign n16214 = n59231 & n16180;
  assign n16215 = ~n16213 & ~n16214;
  assign n16216 = ~n16181 & ~n16212;
  assign n16217 = ~n7716 & ~n59561;
  assign n16218 = n7716 & n16180;
  assign n16219 = n7716 & ~n16180;
  assign n16220 = ~n7716 & n59561;
  assign n16221 = ~n16219 & ~n16220;
  assign n16222 = ~n16217 & ~n16218;
  assign n16223 = ~n7762 & n59562;
  assign n16224 = n7762 & n16180;
  assign n16225 = ~n16223 & ~n16224;
  assign n16226 = ~pi792 & n16225;
  assign n16227 = pi628 & ~n16225;
  assign n16228 = ~pi628 & n16180;
  assign n16229 = pi1156 & ~n16228;
  assign n16230 = ~n16227 & n16229;
  assign n16231 = ~pi628 & ~n16225;
  assign n16232 = pi628 & n16180;
  assign n16233 = ~pi1156 & ~n16232;
  assign n16234 = ~n16231 & n16233;
  assign n16235 = ~n16230 & ~n16234;
  assign n16236 = pi792 & ~n16235;
  assign n16237 = ~n16226 & ~n16236;
  assign n16238 = pi647 & n16237;
  assign n16239 = ~pi647 & n16180;
  assign n16240 = pi647 & ~n16237;
  assign n16241 = ~pi647 & ~n16180;
  assign n16242 = ~n16240 & ~n16241;
  assign n16243 = ~n16238 & ~n16239;
  assign n16244 = pi1157 & ~n59563;
  assign n16245 = ~pi647 & n16237;
  assign n16246 = pi647 & n16180;
  assign n16247 = ~pi1157 & ~n16246;
  assign n16248 = ~n16245 & n16247;
  assign n16249 = ~pi647 & ~n16237;
  assign n16250 = pi647 & ~n16180;
  assign n16251 = ~n16249 & ~n16250;
  assign n16252 = ~pi1157 & n16251;
  assign n16253 = pi1157 & n59563;
  assign n16254 = ~n16252 & ~n16253;
  assign n16255 = ~n16244 & ~n16248;
  assign n16256 = pi787 & n59564;
  assign n16257 = ~pi787 & ~n16237;
  assign n16258 = pi787 & ~n59564;
  assign n16259 = ~pi787 & n16237;
  assign n16260 = ~n16258 & ~n16259;
  assign n16261 = ~n16256 & ~n16257;
  assign n16262 = ~pi644 & ~n59565;
  assign n16263 = pi715 & ~n16262;
  assign n16264 = pi181 & ~n59132;
  assign n16265 = pi754 & n6654;
  assign n16266 = pi181 & n6853;
  assign n16267 = ~n16265 & ~n16266;
  assign n16268 = pi39 & ~n16267;
  assign n16269 = ~pi181 & ~pi754;
  assign n16270 = n59164 & n16269;
  assign n16271 = pi181 & pi754;
  assign n16272 = pi754 & n59147;
  assign n16273 = pi181 & ~n6798;
  assign n16274 = ~n16272 & ~n16273;
  assign n16275 = ~pi39 & ~n16274;
  assign n16276 = ~n16271 & ~n16275;
  assign n16277 = ~n16270 & n16276;
  assign n16278 = ~n16268 & n16277;
  assign n16279 = ~pi38 & ~n16278;
  assign n16280 = ~pi754 & n6865;
  assign n16281 = pi38 & ~n16189;
  assign n16282 = ~n16280 & n16281;
  assign n16283 = ~n16279 & ~n16282;
  assign n16284 = n59132 & ~n16283;
  assign n16285 = ~n16264 & ~n16284;
  assign n16286 = ~n7597 & ~n16285;
  assign n16287 = n7597 & ~n16180;
  assign n16288 = ~n16286 & ~n16287;
  assign n16289 = ~pi785 & ~n16288;
  assign n16290 = ~n7598 & ~n16180;
  assign n16291 = pi609 & n16286;
  assign n16292 = ~n16290 & ~n16291;
  assign n16293 = pi1155 & ~n16292;
  assign n16294 = ~n7610 & ~n16180;
  assign n16295 = ~pi609 & n16286;
  assign n16296 = ~n16294 & ~n16295;
  assign n16297 = ~pi1155 & ~n16296;
  assign n16298 = ~n16293 & ~n16297;
  assign n16299 = pi785 & ~n16298;
  assign n16300 = ~n16289 & ~n16299;
  assign n16301 = ~pi781 & ~n16300;
  assign n16302 = pi618 & n16300;
  assign n16303 = ~pi618 & n16180;
  assign n16304 = pi1154 & ~n16303;
  assign n16305 = ~n16302 & n16304;
  assign n16306 = ~pi618 & n16300;
  assign n16307 = pi618 & n16180;
  assign n16308 = ~pi1154 & ~n16307;
  assign n16309 = ~n16306 & n16308;
  assign n16310 = ~n16305 & ~n16309;
  assign n16311 = pi781 & ~n16310;
  assign n16312 = ~n16301 & ~n16311;
  assign n16313 = ~pi789 & ~n16312;
  assign n16314 = pi619 & n16312;
  assign n16315 = ~pi619 & n16180;
  assign n16316 = pi1159 & ~n16315;
  assign n16317 = ~n16314 & n16316;
  assign n16318 = ~pi619 & n16312;
  assign n16319 = pi619 & n16180;
  assign n16320 = ~pi1159 & ~n16319;
  assign n16321 = ~n16318 & n16320;
  assign n16322 = ~n16317 & ~n16321;
  assign n16323 = pi789 & ~n16322;
  assign n16324 = ~n16313 & ~n16323;
  assign n16325 = ~n8054 & n16324;
  assign n16326 = n8054 & n16180;
  assign n16327 = ~n16325 & ~n16326;
  assign n16328 = ~n7793 & ~n16327;
  assign n16329 = n7793 & n16180;
  assign n16330 = ~n16328 & ~n16329;
  assign n16331 = ~n7835 & ~n16330;
  assign n16332 = n7835 & n16180;
  assign n16333 = n7835 & ~n16180;
  assign n16334 = ~n7835 & n16330;
  assign n16335 = ~n16333 & ~n16334;
  assign n16336 = ~n16331 & ~n16332;
  assign n16337 = pi644 & n59566;
  assign n16338 = ~pi644 & n16180;
  assign n16339 = ~pi715 & ~n16338;
  assign n16340 = ~n16337 & n16339;
  assign n16341 = pi1160 & ~n16340;
  assign n16342 = ~n16263 & n16341;
  assign n16343 = pi644 & ~n59565;
  assign n16344 = ~pi715 & ~n16343;
  assign n16345 = ~pi644 & n59566;
  assign n16346 = pi644 & n16180;
  assign n16347 = pi715 & ~n16346;
  assign n16348 = ~n16345 & n16347;
  assign n16349 = ~pi1160 & ~n16348;
  assign n16350 = ~n16344 & n16349;
  assign n16351 = ~n16342 & ~n16350;
  assign n16352 = pi790 & ~n16351;
  assign n16353 = ~pi644 & n16349;
  assign n16354 = pi644 & n16341;
  assign n16355 = pi790 & ~n16354;
  assign n16356 = pi790 & ~n16353;
  assign n16357 = ~n16354 & n16356;
  assign n16358 = ~n16353 & n16355;
  assign n16359 = ~n7872 & n16330;
  assign n16360 = n7832 & ~n59563;
  assign n16361 = n7833 & ~n16251;
  assign n16362 = pi630 & n16248;
  assign n16363 = ~n16360 & ~n59568;
  assign n16364 = ~n16359 & n16363;
  assign n16365 = pi787 & ~n16364;
  assign n16366 = ~n11154 & n16327;
  assign n16367 = ~pi629 & n16230;
  assign n16368 = pi629 & n16234;
  assign n16369 = ~n16367 & ~n16368;
  assign n16370 = ~n16366 & n16369;
  assign n16371 = pi792 & ~n16370;
  assign n16372 = pi709 & n16283;
  assign n16373 = ~pi181 & n59177;
  assign n16374 = pi181 & n7111;
  assign n16375 = pi754 & ~n16374;
  assign n16376 = ~n16373 & n16375;
  assign n16377 = pi181 & n7188;
  assign n16378 = ~pi181 & ~n59203;
  assign n16379 = ~pi754 & ~n16378;
  assign n16380 = ~n16377 & n16379;
  assign n16381 = pi39 & ~n16380;
  assign n16382 = ~n16376 & n16381;
  assign n16383 = pi181 & n7333;
  assign n16384 = ~pi181 & n7310;
  assign n16385 = pi754 & ~n16384;
  assign n16386 = ~n16383 & n16385;
  assign n16387 = ~pi181 & ~n7339;
  assign n16388 = pi181 & ~n7347;
  assign n16389 = ~pi754 & ~n16388;
  assign n16390 = ~n16387 & n16389;
  assign n16391 = ~pi39 & ~n16390;
  assign n16392 = pi181 & ~n7333;
  assign n16393 = ~pi181 & ~n7310;
  assign n16394 = pi754 & ~n16393;
  assign n16395 = pi754 & ~n16392;
  assign n16396 = ~n16393 & n16395;
  assign n16397 = ~n16392 & n16394;
  assign n16398 = ~pi181 & n7339;
  assign n16399 = pi181 & n7347;
  assign n16400 = ~pi754 & ~n16399;
  assign n16401 = ~n16398 & n16400;
  assign n16402 = ~n59569 & ~n16401;
  assign n16403 = ~pi39 & ~n16402;
  assign n16404 = ~n16386 & n16391;
  assign n16405 = ~pi38 & ~n59570;
  assign n16406 = ~n16382 & n16405;
  assign n16407 = ~pi754 & ~n7222;
  assign n16408 = n9794 & ~n16407;
  assign n16409 = ~pi181 & ~n16408;
  assign n16410 = ~n7056 & ~n15973;
  assign n16411 = pi181 & ~n16410;
  assign n16412 = n59171 & n16411;
  assign n16413 = pi38 & ~n16412;
  assign n16414 = ~n16409 & n16413;
  assign n16415 = ~pi709 & ~n16414;
  assign n16416 = ~n16406 & n16415;
  assign n16417 = n59132 & ~n16416;
  assign n16418 = ~n16372 & n16417;
  assign n16419 = ~n16264 & ~n16418;
  assign n16420 = ~pi625 & n16419;
  assign n16421 = pi625 & n16285;
  assign n16422 = ~pi1153 & ~n16421;
  assign n16423 = ~n16420 & n16422;
  assign n16424 = ~pi608 & ~n16198;
  assign n16425 = ~n16423 & n16424;
  assign n16426 = pi625 & n16419;
  assign n16427 = ~pi625 & n16285;
  assign n16428 = pi1153 & ~n16427;
  assign n16429 = ~n16426 & n16428;
  assign n16430 = pi608 & ~n16202;
  assign n16431 = ~n16429 & n16430;
  assign n16432 = ~n16425 & ~n16431;
  assign n16433 = pi778 & ~n16432;
  assign n16434 = ~pi778 & n16419;
  assign n16435 = ~n16433 & ~n16434;
  assign n16436 = ~pi609 & ~n16435;
  assign n16437 = pi609 & n16205;
  assign n16438 = ~pi1155 & ~n16437;
  assign n16439 = ~n16436 & n16438;
  assign n16440 = ~pi660 & ~n16293;
  assign n16441 = ~n16439 & n16440;
  assign n16442 = pi609 & ~n16435;
  assign n16443 = ~pi609 & n16205;
  assign n16444 = pi1155 & ~n16443;
  assign n16445 = ~n16442 & n16444;
  assign n16446 = pi660 & ~n16297;
  assign n16447 = ~n16445 & n16446;
  assign n16448 = ~n16441 & ~n16447;
  assign n16449 = pi785 & ~n16448;
  assign n16450 = ~pi785 & ~n16435;
  assign n16451 = ~n16449 & ~n16450;
  assign n16452 = ~pi618 & ~n16451;
  assign n16453 = pi618 & n59560;
  assign n16454 = ~pi1154 & ~n16453;
  assign n16455 = ~n16452 & n16454;
  assign n16456 = ~pi627 & ~n16305;
  assign n16457 = ~n16455 & n16456;
  assign n16458 = pi618 & ~n16451;
  assign n16459 = ~pi618 & n59560;
  assign n16460 = pi1154 & ~n16459;
  assign n16461 = ~n16458 & n16460;
  assign n16462 = pi627 & ~n16309;
  assign n16463 = ~n16461 & n16462;
  assign n16464 = ~n16457 & ~n16463;
  assign n16465 = pi781 & ~n16464;
  assign n16466 = ~pi781 & ~n16451;
  assign n16467 = ~n16465 & ~n16466;
  assign n16468 = pi619 & ~n16467;
  assign n16469 = ~pi619 & ~n59561;
  assign n16470 = pi1159 & ~n16469;
  assign n16471 = ~n16468 & n16470;
  assign n16472 = pi648 & ~n16321;
  assign n16473 = ~n16471 & n16472;
  assign n16474 = ~pi619 & ~n16467;
  assign n16475 = pi619 & ~n59561;
  assign n16476 = ~pi1159 & ~n16475;
  assign n16477 = ~n16474 & n16476;
  assign n16478 = ~pi648 & ~n16317;
  assign n16479 = ~n16477 & n16478;
  assign n16480 = pi789 & ~n16479;
  assign n16481 = pi789 & ~n16473;
  assign n16482 = ~n16479 & n16481;
  assign n16483 = ~n16473 & n16480;
  assign n16484 = ~pi789 & n16467;
  assign n16485 = n59242 & ~n16484;
  assign n16486 = ~n59571 & n16485;
  assign n16487 = ~pi626 & ~n16324;
  assign n16488 = pi626 & ~n16180;
  assign n16489 = n7760 & ~n16488;
  assign n16490 = ~n16487 & n16489;
  assign n16491 = n7984 & n59562;
  assign n16492 = pi626 & ~n16324;
  assign n16493 = ~pi626 & ~n16180;
  assign n16494 = n7759 & ~n16493;
  assign n16495 = ~n16492 & n16494;
  assign n16496 = ~n16491 & ~n16495;
  assign n16497 = ~n16490 & ~n16491;
  assign n16498 = ~n16495 & n16497;
  assign n16499 = ~n16490 & n16496;
  assign n16500 = pi788 & ~n59572;
  assign n16501 = ~n59357 & ~n16500;
  assign n16502 = ~n16486 & n16501;
  assign n16503 = ~n16371 & ~n16502;
  assign n16504 = ~n8108 & ~n16503;
  assign n16505 = ~n16365 & ~n16504;
  assign n16506 = ~n59567 & n16505;
  assign n16507 = ~n16352 & ~n16506;
  assign n16508 = n58992 & ~n16507;
  assign n16509 = ~pi181 & ~n58992;
  assign n16510 = ~pi832 & ~n16509;
  assign n16511 = ~n16508 & n16510;
  assign po338 = ~n16179 & ~n16511;
  assign n16513 = ~pi182 & ~n2794;
  assign n16514 = ~pi756 & n6822;
  assign n16515 = ~n16513 & ~n16514;
  assign n16516 = ~n7875 & ~n16515;
  assign n16517 = ~pi785 & ~n16516;
  assign n16518 = n7610 & n16514;
  assign n16519 = n16516 & ~n16518;
  assign n16520 = pi1155 & ~n16519;
  assign n16521 = ~pi1155 & ~n16513;
  assign n16522 = ~n16518 & n16521;
  assign n16523 = ~n16520 & ~n16522;
  assign n16524 = pi785 & ~n16523;
  assign n16525 = ~n16517 & ~n16524;
  assign n16526 = ~pi781 & ~n16525;
  assign n16527 = ~n7890 & n16525;
  assign n16528 = pi1154 & ~n16527;
  assign n16529 = ~n7893 & n16525;
  assign n16530 = ~pi1154 & ~n16529;
  assign n16531 = ~n16528 & ~n16530;
  assign n16532 = pi781 & ~n16531;
  assign n16533 = ~n16526 & ~n16532;
  assign n16534 = ~pi789 & ~n16533;
  assign n16535 = ~n11882 & n16533;
  assign n16536 = pi1159 & ~n16535;
  assign n16537 = ~n11885 & n16533;
  assign n16538 = ~pi1159 & ~n16537;
  assign n16539 = ~n16536 & ~n16538;
  assign n16540 = pi789 & ~n16539;
  assign n16541 = ~n16534 & ~n16540;
  assign n16542 = ~n8054 & ~n16541;
  assign n16543 = n8054 & ~n16513;
  assign n16544 = ~n8054 & n16541;
  assign n16545 = n8054 & n16513;
  assign n16546 = ~n16544 & ~n16545;
  assign n16547 = ~n16542 & ~n16543;
  assign n16548 = ~n7793 & ~n59573;
  assign n16549 = n7793 & n16513;
  assign n16550 = ~n7872 & ~n16549;
  assign n16551 = ~n16548 & ~n16549;
  assign n16552 = ~n7872 & n16551;
  assign n16553 = ~n16548 & n16550;
  assign n16554 = ~pi734 & n7055;
  assign n16555 = ~n16513 & ~n16554;
  assign n16556 = ~pi778 & ~n16555;
  assign n16557 = ~pi625 & n16554;
  assign n16558 = ~n16555 & ~n16557;
  assign n16559 = pi1153 & ~n16558;
  assign n16560 = ~pi1153 & ~n16513;
  assign n16561 = ~n16557 & n16560;
  assign n16562 = pi778 & ~n16561;
  assign n16563 = ~n16559 & n16562;
  assign n16564 = ~n16556 & ~n16563;
  assign n16565 = ~n7949 & ~n16564;
  assign n16566 = ~n7951 & n16565;
  assign n16567 = ~n7953 & n16566;
  assign n16568 = ~n7955 & n16567;
  assign n16569 = ~n7967 & n16568;
  assign n16570 = pi647 & ~n16569;
  assign n16571 = ~pi647 & ~n16513;
  assign n16572 = ~n16570 & ~n16571;
  assign n16573 = n7832 & ~n16572;
  assign n16574 = ~pi647 & n16569;
  assign n16575 = pi647 & n16513;
  assign n16576 = ~pi1157 & ~n16575;
  assign n16577 = ~n16574 & n16576;
  assign n16578 = pi630 & n16577;
  assign n16579 = ~n16573 & ~n16578;
  assign n16580 = ~n59574 & n16579;
  assign n16581 = pi787 & ~n16580;
  assign n16582 = ~pi626 & ~n16541;
  assign n16583 = pi626 & ~n16513;
  assign n16584 = n7760 & ~n16583;
  assign n16585 = ~n16582 & n16584;
  assign n16586 = n7984 & n16567;
  assign n16587 = pi626 & ~n16541;
  assign n16588 = ~pi626 & ~n16513;
  assign n16589 = n7759 & ~n16588;
  assign n16590 = ~n16587 & n16589;
  assign n16591 = ~n16586 & ~n16590;
  assign n16592 = ~n16585 & ~n16586;
  assign n16593 = ~n16590 & n16592;
  assign n16594 = ~n16585 & n16591;
  assign n16595 = pi788 & ~n59575;
  assign n16596 = ~n6701 & ~n16555;
  assign n16597 = pi625 & n16596;
  assign n16598 = n16515 & ~n16596;
  assign n16599 = ~n16597 & ~n16598;
  assign n16600 = n16560 & ~n16599;
  assign n16601 = ~pi608 & ~n16559;
  assign n16602 = ~n16600 & n16601;
  assign n16603 = pi1153 & n16515;
  assign n16604 = ~n16597 & n16603;
  assign n16605 = pi608 & ~n16561;
  assign n16606 = ~n16604 & n16605;
  assign n16607 = ~n16602 & ~n16606;
  assign n16608 = pi778 & ~n16607;
  assign n16609 = ~pi778 & ~n16598;
  assign n16610 = ~n16608 & ~n16609;
  assign n16611 = ~pi609 & ~n16610;
  assign n16612 = pi609 & ~n16564;
  assign n16613 = ~pi1155 & ~n16612;
  assign n16614 = ~n16611 & n16613;
  assign n16615 = ~pi660 & ~n16520;
  assign n16616 = ~n16614 & n16615;
  assign n16617 = pi609 & ~n16610;
  assign n16618 = ~pi609 & ~n16564;
  assign n16619 = pi1155 & ~n16618;
  assign n16620 = ~n16617 & n16619;
  assign n16621 = pi660 & ~n16522;
  assign n16622 = ~n16620 & n16621;
  assign n16623 = ~n16616 & ~n16622;
  assign n16624 = pi785 & ~n16623;
  assign n16625 = ~pi785 & ~n16610;
  assign n16626 = ~n16624 & ~n16625;
  assign n16627 = ~pi618 & ~n16626;
  assign n16628 = pi618 & n16565;
  assign n16629 = ~pi1154 & ~n16628;
  assign n16630 = ~n16627 & n16629;
  assign n16631 = ~pi627 & ~n16528;
  assign n16632 = ~n16630 & n16631;
  assign n16633 = pi618 & ~n16626;
  assign n16634 = ~pi618 & n16565;
  assign n16635 = pi1154 & ~n16634;
  assign n16636 = ~n16633 & n16635;
  assign n16637 = pi627 & ~n16530;
  assign n16638 = ~n16636 & n16637;
  assign n16639 = ~n16632 & ~n16638;
  assign n16640 = pi781 & ~n16639;
  assign n16641 = ~pi781 & ~n16626;
  assign n16642 = ~n16640 & ~n16641;
  assign n16643 = pi619 & ~n16642;
  assign n16644 = ~pi619 & n16566;
  assign n16645 = pi1159 & ~n16644;
  assign n16646 = ~n16643 & n16645;
  assign n16647 = pi648 & ~n16538;
  assign n16648 = ~n16646 & n16647;
  assign n16649 = ~pi619 & ~n16642;
  assign n16650 = pi619 & n16566;
  assign n16651 = ~pi1159 & ~n16650;
  assign n16652 = ~n16649 & n16651;
  assign n16653 = ~pi648 & ~n16536;
  assign n16654 = ~n16652 & n16653;
  assign n16655 = pi789 & ~n16654;
  assign n16656 = pi789 & ~n16648;
  assign n16657 = ~n16654 & n16656;
  assign n16658 = ~n16648 & n16655;
  assign n16659 = ~pi789 & n16642;
  assign n16660 = n59242 & ~n16659;
  assign n16661 = ~n59576 & n16660;
  assign n16662 = ~n16595 & ~n16661;
  assign n16663 = ~n59357 & ~n16662;
  assign n16664 = n7957 & ~n59573;
  assign n16665 = n8065 & n16568;
  assign n16666 = pi629 & ~n16665;
  assign n16667 = ~n16664 & n16666;
  assign n16668 = n7958 & ~n59573;
  assign n16669 = n8074 & n16568;
  assign n16670 = ~pi629 & ~n16669;
  assign n16671 = ~n16668 & n16670;
  assign n16672 = pi792 & ~n16671;
  assign n16673 = ~n16668 & ~n16669;
  assign n16674 = ~pi629 & ~n16673;
  assign n16675 = ~n16664 & ~n16665;
  assign n16676 = pi629 & ~n16675;
  assign n16677 = ~n16674 & ~n16676;
  assign n16678 = pi792 & ~n16677;
  assign n16679 = pi792 & ~n16667;
  assign n16680 = ~n16671 & n16679;
  assign n16681 = ~n16667 & n16672;
  assign n16682 = ~n8108 & ~n59577;
  assign n16683 = ~n16663 & n16682;
  assign n16684 = ~n16581 & ~n16683;
  assign n16685 = pi644 & n16684;
  assign n16686 = ~pi787 & ~n16569;
  assign n16687 = pi1157 & ~n16572;
  assign n16688 = ~n16577 & ~n16687;
  assign n16689 = pi787 & ~n16688;
  assign n16690 = ~n16686 & ~n16689;
  assign n16691 = ~pi644 & n16690;
  assign n16692 = pi715 & ~n16691;
  assign n16693 = ~n16685 & n16692;
  assign n16694 = ~n11491 & n16513;
  assign n16695 = ~n7835 & n16548;
  assign n16696 = ~n7835 & ~n16551;
  assign n16697 = n7835 & n16513;
  assign n16698 = ~n16696 & ~n16697;
  assign n16699 = ~n16694 & ~n16695;
  assign n16700 = pi644 & ~n59578;
  assign n16701 = ~pi644 & n16513;
  assign n16702 = ~pi715 & ~n16701;
  assign n16703 = ~n16700 & n16702;
  assign n16704 = pi1160 & ~n16703;
  assign n16705 = ~n16693 & n16704;
  assign n16706 = ~pi644 & n16684;
  assign n16707 = pi644 & n16690;
  assign n16708 = ~pi715 & ~n16707;
  assign n16709 = ~n16706 & n16708;
  assign n16710 = ~pi644 & ~n59578;
  assign n16711 = pi644 & n16513;
  assign n16712 = pi715 & ~n16711;
  assign n16713 = ~n16710 & n16712;
  assign n16714 = ~pi1160 & ~n16713;
  assign n16715 = ~n16709 & n16714;
  assign n16716 = ~n16705 & ~n16715;
  assign n16717 = pi790 & ~n16716;
  assign n16718 = ~pi790 & n16684;
  assign n16719 = pi832 & ~n16718;
  assign n16720 = ~n16717 & n16719;
  assign n16721 = ~pi182 & ~n7560;
  assign n16722 = n59231 & ~n16721;
  assign n16723 = ~pi734 & n59132;
  assign n16724 = n16721 & ~n16723;
  assign n16725 = pi182 & n59251;
  assign n16726 = ~pi38 & ~n16725;
  assign n16727 = n59132 & ~n16726;
  assign n16728 = ~pi182 & n8249;
  assign n16729 = ~n16727 & ~n16728;
  assign n16730 = ~pi182 & ~n6863;
  assign n16731 = n7547 & ~n16730;
  assign n16732 = ~pi734 & ~n16731;
  assign n16733 = ~n16729 & n16732;
  assign n16734 = ~n16724 & ~n16733;
  assign n16735 = ~pi778 & n16734;
  assign n16736 = pi625 & ~n16734;
  assign n16737 = ~pi625 & n16721;
  assign n16738 = pi1153 & ~n16737;
  assign n16739 = ~n16736 & n16738;
  assign n16740 = ~pi625 & ~n16734;
  assign n16741 = pi625 & n16721;
  assign n16742 = ~pi1153 & ~n16741;
  assign n16743 = ~n16740 & n16742;
  assign n16744 = ~n16739 & ~n16743;
  assign n16745 = pi778 & ~n16744;
  assign n16746 = ~n16735 & ~n16745;
  assign n16747 = ~n59229 & n16746;
  assign n16748 = n59229 & n16721;
  assign n16749 = n59229 & ~n16721;
  assign n16750 = ~n59229 & ~n16746;
  assign n16751 = ~n16749 & ~n16750;
  assign n16752 = ~n16747 & ~n16748;
  assign n16753 = ~n59231 & ~n59579;
  assign n16754 = ~n59231 & n59579;
  assign n16755 = n59231 & n16721;
  assign n16756 = ~n16754 & ~n16755;
  assign n16757 = ~n16722 & ~n16753;
  assign n16758 = ~n7716 & ~n59580;
  assign n16759 = n7716 & n16721;
  assign n16760 = n7716 & ~n16721;
  assign n16761 = ~n7716 & n59580;
  assign n16762 = ~n16760 & ~n16761;
  assign n16763 = ~n16758 & ~n16759;
  assign n16764 = ~n7762 & n59581;
  assign n16765 = n7762 & n16721;
  assign n16766 = ~n16764 & ~n16765;
  assign n16767 = ~pi792 & n16766;
  assign n16768 = pi628 & ~n16766;
  assign n16769 = ~pi628 & n16721;
  assign n16770 = pi1156 & ~n16769;
  assign n16771 = ~n16768 & n16770;
  assign n16772 = ~pi628 & ~n16766;
  assign n16773 = pi628 & n16721;
  assign n16774 = ~pi1156 & ~n16773;
  assign n16775 = ~n16772 & n16774;
  assign n16776 = ~n16771 & ~n16775;
  assign n16777 = pi792 & ~n16776;
  assign n16778 = ~n16767 & ~n16777;
  assign n16779 = pi647 & n16778;
  assign n16780 = ~pi647 & n16721;
  assign n16781 = pi647 & ~n16778;
  assign n16782 = ~pi647 & ~n16721;
  assign n16783 = ~n16781 & ~n16782;
  assign n16784 = ~n16779 & ~n16780;
  assign n16785 = pi1157 & ~n59582;
  assign n16786 = ~pi647 & n16778;
  assign n16787 = pi647 & n16721;
  assign n16788 = ~pi1157 & ~n16787;
  assign n16789 = ~n16786 & n16788;
  assign n16790 = ~pi647 & ~n16778;
  assign n16791 = pi647 & ~n16721;
  assign n16792 = ~n16790 & ~n16791;
  assign n16793 = ~pi1157 & n16792;
  assign n16794 = pi1157 & n59582;
  assign n16795 = ~n16793 & ~n16794;
  assign n16796 = ~n16785 & ~n16789;
  assign n16797 = pi787 & n59583;
  assign n16798 = ~pi787 & ~n16778;
  assign n16799 = pi787 & ~n59583;
  assign n16800 = ~pi787 & n16778;
  assign n16801 = ~n16799 & ~n16800;
  assign n16802 = ~n16797 & ~n16798;
  assign n16803 = ~pi644 & ~n59584;
  assign n16804 = pi715 & ~n16803;
  assign n16805 = pi182 & ~n59132;
  assign n16806 = ~pi756 & n6865;
  assign n16807 = ~n16730 & ~n16806;
  assign n16808 = pi38 & ~n16807;
  assign n16809 = ~pi182 & n59164;
  assign n16810 = pi182 & ~n6855;
  assign n16811 = ~pi756 & ~n16810;
  assign n16812 = ~n16809 & n16811;
  assign n16813 = ~pi182 & pi756;
  assign n16814 = ~n6656 & n16813;
  assign n16815 = pi756 & ~n6656;
  assign n16816 = ~pi756 & ~n16809;
  assign n16817 = ~n16815 & ~n16816;
  assign n16818 = ~pi182 & ~n16817;
  assign n16819 = n6855 & n16816;
  assign n16820 = ~n16818 & ~n16819;
  assign n16821 = ~n16812 & ~n16814;
  assign n16822 = ~pi38 & ~n59585;
  assign n16823 = ~n16808 & ~n16822;
  assign n16824 = n59132 & n16823;
  assign n16825 = ~n16805 & ~n16824;
  assign n16826 = ~n7597 & ~n16825;
  assign n16827 = n7597 & ~n16721;
  assign n16828 = ~n16826 & ~n16827;
  assign n16829 = ~pi785 & ~n16828;
  assign n16830 = ~n7598 & ~n16721;
  assign n16831 = pi609 & n16826;
  assign n16832 = ~n16830 & ~n16831;
  assign n16833 = pi1155 & ~n16832;
  assign n16834 = ~n7610 & ~n16721;
  assign n16835 = ~pi609 & n16826;
  assign n16836 = ~n16834 & ~n16835;
  assign n16837 = ~pi1155 & ~n16836;
  assign n16838 = ~n16833 & ~n16837;
  assign n16839 = pi785 & ~n16838;
  assign n16840 = ~n16829 & ~n16839;
  assign n16841 = ~pi781 & ~n16840;
  assign n16842 = pi618 & n16840;
  assign n16843 = ~pi618 & n16721;
  assign n16844 = pi1154 & ~n16843;
  assign n16845 = ~n16842 & n16844;
  assign n16846 = ~pi618 & n16840;
  assign n16847 = pi618 & n16721;
  assign n16848 = ~pi1154 & ~n16847;
  assign n16849 = ~n16846 & n16848;
  assign n16850 = ~n16845 & ~n16849;
  assign n16851 = pi781 & ~n16850;
  assign n16852 = ~n16841 & ~n16851;
  assign n16853 = ~pi789 & ~n16852;
  assign n16854 = pi619 & n16852;
  assign n16855 = ~pi619 & n16721;
  assign n16856 = pi1159 & ~n16855;
  assign n16857 = ~n16854 & n16856;
  assign n16858 = ~pi619 & n16852;
  assign n16859 = pi619 & n16721;
  assign n16860 = ~pi1159 & ~n16859;
  assign n16861 = ~n16858 & n16860;
  assign n16862 = ~n16857 & ~n16861;
  assign n16863 = pi789 & ~n16862;
  assign n16864 = ~n16853 & ~n16863;
  assign n16865 = ~n8054 & n16864;
  assign n16866 = n8054 & n16721;
  assign n16867 = ~n16865 & ~n16866;
  assign n16868 = ~n7793 & ~n16867;
  assign n16869 = n7793 & n16721;
  assign n16870 = ~n16868 & ~n16869;
  assign n16871 = ~n7835 & ~n16870;
  assign n16872 = n7835 & n16721;
  assign n16873 = n7835 & ~n16721;
  assign n16874 = ~n7835 & n16870;
  assign n16875 = ~n16873 & ~n16874;
  assign n16876 = ~n16871 & ~n16872;
  assign n16877 = pi644 & n59586;
  assign n16878 = ~pi644 & n16721;
  assign n16879 = ~pi715 & ~n16878;
  assign n16880 = ~n16877 & n16879;
  assign n16881 = pi1160 & ~n16880;
  assign n16882 = ~n16804 & n16881;
  assign n16883 = pi644 & ~n59584;
  assign n16884 = ~pi715 & ~n16883;
  assign n16885 = ~pi644 & n59586;
  assign n16886 = pi644 & n16721;
  assign n16887 = pi715 & ~n16886;
  assign n16888 = ~n16885 & n16887;
  assign n16889 = ~pi1160 & ~n16888;
  assign n16890 = ~n16884 & n16889;
  assign n16891 = ~n16882 & ~n16890;
  assign n16892 = pi790 & ~n16891;
  assign n16893 = ~pi644 & n16889;
  assign n16894 = pi644 & n16881;
  assign n16895 = pi790 & ~n16894;
  assign n16896 = pi790 & ~n16893;
  assign n16897 = ~n16894 & n16896;
  assign n16898 = ~n16893 & n16895;
  assign n16899 = ~n7872 & n16870;
  assign n16900 = n7832 & ~n59582;
  assign n16901 = n7833 & ~n16792;
  assign n16902 = pi630 & n16789;
  assign n16903 = ~n16900 & ~n59588;
  assign n16904 = ~n16899 & n16903;
  assign n16905 = pi787 & ~n16904;
  assign n16906 = ~n11154 & n16867;
  assign n16907 = ~pi629 & n16771;
  assign n16908 = pi629 & n16775;
  assign n16909 = ~n16907 & ~n16908;
  assign n16910 = ~n16906 & n16909;
  assign n16911 = pi792 & ~n16910;
  assign n16912 = pi734 & ~n16823;
  assign n16913 = ~pi182 & n59177;
  assign n16914 = pi182 & n7111;
  assign n16915 = pi756 & ~n16914;
  assign n16916 = ~n16913 & n16915;
  assign n16917 = pi182 & n7188;
  assign n16918 = ~pi182 & ~n59203;
  assign n16919 = ~pi756 & ~n16918;
  assign n16920 = ~n16917 & n16919;
  assign n16921 = pi39 & ~n16920;
  assign n16922 = ~n16916 & n16921;
  assign n16923 = pi182 & n7333;
  assign n16924 = ~pi182 & n7310;
  assign n16925 = pi756 & ~n16924;
  assign n16926 = ~n16923 & n16925;
  assign n16927 = ~pi182 & ~n7339;
  assign n16928 = pi182 & ~n7347;
  assign n16929 = ~pi756 & ~n16928;
  assign n16930 = ~n16927 & n16929;
  assign n16931 = ~pi39 & ~n16930;
  assign n16932 = pi182 & ~n7333;
  assign n16933 = ~pi182 & ~n7310;
  assign n16934 = pi756 & ~n16933;
  assign n16935 = pi756 & ~n16932;
  assign n16936 = ~n16933 & n16935;
  assign n16937 = ~n16932 & n16934;
  assign n16938 = ~pi182 & n7339;
  assign n16939 = pi182 & n7347;
  assign n16940 = ~pi756 & ~n16939;
  assign n16941 = ~n16938 & n16940;
  assign n16942 = ~n59589 & ~n16941;
  assign n16943 = ~pi39 & ~n16942;
  assign n16944 = ~n16926 & n16931;
  assign n16945 = ~pi38 & ~n59590;
  assign n16946 = ~n16922 & n16945;
  assign n16947 = ~pi756 & ~n7222;
  assign n16948 = n9794 & ~n16947;
  assign n16949 = ~pi182 & ~n16948;
  assign n16950 = ~n7056 & ~n16514;
  assign n16951 = pi182 & ~n16950;
  assign n16952 = n59171 & n16951;
  assign n16953 = pi38 & ~n16952;
  assign n16954 = ~n16949 & n16953;
  assign n16955 = ~pi734 & ~n16954;
  assign n16956 = ~n16946 & n16955;
  assign n16957 = n59132 & ~n16956;
  assign n16958 = ~n16912 & n16957;
  assign n16959 = ~n16805 & ~n16958;
  assign n16960 = ~pi625 & n16959;
  assign n16961 = pi625 & n16825;
  assign n16962 = ~pi1153 & ~n16961;
  assign n16963 = ~n16960 & n16962;
  assign n16964 = ~pi608 & ~n16739;
  assign n16965 = ~n16963 & n16964;
  assign n16966 = pi625 & n16959;
  assign n16967 = ~pi625 & n16825;
  assign n16968 = pi1153 & ~n16967;
  assign n16969 = ~n16966 & n16968;
  assign n16970 = pi608 & ~n16743;
  assign n16971 = ~n16969 & n16970;
  assign n16972 = ~n16965 & ~n16971;
  assign n16973 = pi778 & ~n16972;
  assign n16974 = ~pi778 & n16959;
  assign n16975 = ~n16973 & ~n16974;
  assign n16976 = ~pi609 & ~n16975;
  assign n16977 = pi609 & n16746;
  assign n16978 = ~pi1155 & ~n16977;
  assign n16979 = ~n16976 & n16978;
  assign n16980 = ~pi660 & ~n16833;
  assign n16981 = ~n16979 & n16980;
  assign n16982 = pi609 & ~n16975;
  assign n16983 = ~pi609 & n16746;
  assign n16984 = pi1155 & ~n16983;
  assign n16985 = ~n16982 & n16984;
  assign n16986 = pi660 & ~n16837;
  assign n16987 = ~n16985 & n16986;
  assign n16988 = ~n16981 & ~n16987;
  assign n16989 = pi785 & ~n16988;
  assign n16990 = ~pi785 & ~n16975;
  assign n16991 = ~n16989 & ~n16990;
  assign n16992 = ~pi618 & ~n16991;
  assign n16993 = pi618 & n59579;
  assign n16994 = ~pi1154 & ~n16993;
  assign n16995 = ~n16992 & n16994;
  assign n16996 = ~pi627 & ~n16845;
  assign n16997 = ~n16995 & n16996;
  assign n16998 = pi618 & ~n16991;
  assign n16999 = ~pi618 & n59579;
  assign n17000 = pi1154 & ~n16999;
  assign n17001 = ~n16998 & n17000;
  assign n17002 = pi627 & ~n16849;
  assign n17003 = ~n17001 & n17002;
  assign n17004 = ~n16997 & ~n17003;
  assign n17005 = pi781 & ~n17004;
  assign n17006 = ~pi781 & ~n16991;
  assign n17007 = ~n17005 & ~n17006;
  assign n17008 = pi619 & ~n17007;
  assign n17009 = ~pi619 & ~n59580;
  assign n17010 = pi1159 & ~n17009;
  assign n17011 = ~n17008 & n17010;
  assign n17012 = pi648 & ~n16861;
  assign n17013 = ~n17011 & n17012;
  assign n17014 = ~pi619 & ~n17007;
  assign n17015 = pi619 & ~n59580;
  assign n17016 = ~pi1159 & ~n17015;
  assign n17017 = ~n17014 & n17016;
  assign n17018 = ~pi648 & ~n16857;
  assign n17019 = ~n17017 & n17018;
  assign n17020 = pi789 & ~n17019;
  assign n17021 = pi789 & ~n17013;
  assign n17022 = ~n17019 & n17021;
  assign n17023 = ~n17013 & n17020;
  assign n17024 = ~pi789 & n17007;
  assign n17025 = n59242 & ~n17024;
  assign n17026 = ~n59591 & n17025;
  assign n17027 = ~pi626 & ~n16864;
  assign n17028 = pi626 & ~n16721;
  assign n17029 = n7760 & ~n17028;
  assign n17030 = ~n17027 & n17029;
  assign n17031 = n7984 & n59581;
  assign n17032 = pi626 & ~n16864;
  assign n17033 = ~pi626 & ~n16721;
  assign n17034 = n7759 & ~n17033;
  assign n17035 = ~n17032 & n17034;
  assign n17036 = ~n17031 & ~n17035;
  assign n17037 = ~n17030 & ~n17031;
  assign n17038 = ~n17035 & n17037;
  assign n17039 = ~n17030 & n17036;
  assign n17040 = pi788 & ~n59592;
  assign n17041 = ~n59357 & ~n17040;
  assign n17042 = ~n17026 & n17041;
  assign n17043 = ~n16911 & ~n17042;
  assign n17044 = ~n8108 & ~n17043;
  assign n17045 = ~n16905 & ~n17044;
  assign n17046 = ~n59587 & n17045;
  assign n17047 = ~n16892 & ~n17046;
  assign n17048 = n58992 & ~n17047;
  assign n17049 = ~pi182 & ~n58992;
  assign n17050 = ~pi832 & ~n17049;
  assign n17051 = ~n17048 & n17050;
  assign po339 = ~n16720 & ~n17051;
  assign n17053 = ~pi183 & ~n2794;
  assign n17054 = ~pi755 & n6822;
  assign n17055 = ~n17053 & ~n17054;
  assign n17056 = ~n7875 & ~n17055;
  assign n17057 = ~pi785 & ~n17056;
  assign n17058 = n7610 & n17054;
  assign n17059 = n17056 & ~n17058;
  assign n17060 = pi1155 & ~n17059;
  assign n17061 = ~pi1155 & ~n17053;
  assign n17062 = ~n17058 & n17061;
  assign n17063 = ~n17060 & ~n17062;
  assign n17064 = pi785 & ~n17063;
  assign n17065 = ~n17057 & ~n17064;
  assign n17066 = ~pi781 & ~n17065;
  assign n17067 = ~n7890 & n17065;
  assign n17068 = pi1154 & ~n17067;
  assign n17069 = ~n7893 & n17065;
  assign n17070 = ~pi1154 & ~n17069;
  assign n17071 = ~n17068 & ~n17070;
  assign n17072 = pi781 & ~n17071;
  assign n17073 = ~n17066 & ~n17072;
  assign n17074 = ~pi789 & ~n17073;
  assign n17075 = ~n11882 & n17073;
  assign n17076 = pi1159 & ~n17075;
  assign n17077 = ~n11885 & n17073;
  assign n17078 = ~pi1159 & ~n17077;
  assign n17079 = ~n17076 & ~n17078;
  assign n17080 = pi789 & ~n17079;
  assign n17081 = ~n17074 & ~n17080;
  assign n17082 = ~n8054 & ~n17081;
  assign n17083 = n8054 & ~n17053;
  assign n17084 = ~n8054 & n17081;
  assign n17085 = n8054 & n17053;
  assign n17086 = ~n17084 & ~n17085;
  assign n17087 = ~n17082 & ~n17083;
  assign n17088 = ~n7793 & ~n59593;
  assign n17089 = n7793 & n17053;
  assign n17090 = ~n7872 & ~n17089;
  assign n17091 = ~n17088 & ~n17089;
  assign n17092 = ~n7872 & n17091;
  assign n17093 = ~n17088 & n17090;
  assign n17094 = ~pi725 & n7055;
  assign n17095 = ~n17053 & ~n17094;
  assign n17096 = ~pi778 & ~n17095;
  assign n17097 = ~pi625 & n17094;
  assign n17098 = ~n17095 & ~n17097;
  assign n17099 = pi1153 & ~n17098;
  assign n17100 = ~pi1153 & ~n17053;
  assign n17101 = ~n17097 & n17100;
  assign n17102 = pi778 & ~n17101;
  assign n17103 = ~n17099 & n17102;
  assign n17104 = ~n17096 & ~n17103;
  assign n17105 = ~n7949 & ~n17104;
  assign n17106 = ~n7951 & n17105;
  assign n17107 = ~n7953 & n17106;
  assign n17108 = ~n7955 & n17107;
  assign n17109 = ~n7967 & n17108;
  assign n17110 = pi647 & ~n17109;
  assign n17111 = ~pi647 & ~n17053;
  assign n17112 = ~n17110 & ~n17111;
  assign n17113 = n7832 & ~n17112;
  assign n17114 = ~pi647 & n17109;
  assign n17115 = pi647 & n17053;
  assign n17116 = ~pi1157 & ~n17115;
  assign n17117 = ~n17114 & n17116;
  assign n17118 = pi630 & n17117;
  assign n17119 = ~n17113 & ~n17118;
  assign n17120 = ~n59594 & n17119;
  assign n17121 = pi787 & ~n17120;
  assign n17122 = ~pi626 & ~n17081;
  assign n17123 = pi626 & ~n17053;
  assign n17124 = n7760 & ~n17123;
  assign n17125 = ~n17122 & n17124;
  assign n17126 = n7984 & n17107;
  assign n17127 = pi626 & ~n17081;
  assign n17128 = ~pi626 & ~n17053;
  assign n17129 = n7759 & ~n17128;
  assign n17130 = ~n17127 & n17129;
  assign n17131 = ~n17126 & ~n17130;
  assign n17132 = ~n17125 & ~n17126;
  assign n17133 = ~n17130 & n17132;
  assign n17134 = ~n17125 & n17131;
  assign n17135 = pi788 & ~n59595;
  assign n17136 = ~n6701 & ~n17095;
  assign n17137 = pi625 & n17136;
  assign n17138 = n17055 & ~n17136;
  assign n17139 = ~n17137 & ~n17138;
  assign n17140 = n17100 & ~n17139;
  assign n17141 = ~pi608 & ~n17099;
  assign n17142 = ~n17140 & n17141;
  assign n17143 = pi1153 & n17055;
  assign n17144 = ~n17137 & n17143;
  assign n17145 = pi608 & ~n17101;
  assign n17146 = ~n17144 & n17145;
  assign n17147 = ~n17142 & ~n17146;
  assign n17148 = pi778 & ~n17147;
  assign n17149 = ~pi778 & ~n17138;
  assign n17150 = ~n17148 & ~n17149;
  assign n17151 = ~pi609 & ~n17150;
  assign n17152 = pi609 & ~n17104;
  assign n17153 = ~pi1155 & ~n17152;
  assign n17154 = ~n17151 & n17153;
  assign n17155 = ~pi660 & ~n17060;
  assign n17156 = ~n17154 & n17155;
  assign n17157 = pi609 & ~n17150;
  assign n17158 = ~pi609 & ~n17104;
  assign n17159 = pi1155 & ~n17158;
  assign n17160 = ~n17157 & n17159;
  assign n17161 = pi660 & ~n17062;
  assign n17162 = ~n17160 & n17161;
  assign n17163 = ~n17156 & ~n17162;
  assign n17164 = pi785 & ~n17163;
  assign n17165 = ~pi785 & ~n17150;
  assign n17166 = ~n17164 & ~n17165;
  assign n17167 = ~pi618 & ~n17166;
  assign n17168 = pi618 & n17105;
  assign n17169 = ~pi1154 & ~n17168;
  assign n17170 = ~n17167 & n17169;
  assign n17171 = ~pi627 & ~n17068;
  assign n17172 = ~n17170 & n17171;
  assign n17173 = pi618 & ~n17166;
  assign n17174 = ~pi618 & n17105;
  assign n17175 = pi1154 & ~n17174;
  assign n17176 = ~n17173 & n17175;
  assign n17177 = pi627 & ~n17070;
  assign n17178 = ~n17176 & n17177;
  assign n17179 = ~n17172 & ~n17178;
  assign n17180 = pi781 & ~n17179;
  assign n17181 = ~pi781 & ~n17166;
  assign n17182 = ~n17180 & ~n17181;
  assign n17183 = pi619 & ~n17182;
  assign n17184 = ~pi619 & n17106;
  assign n17185 = pi1159 & ~n17184;
  assign n17186 = ~n17183 & n17185;
  assign n17187 = pi648 & ~n17078;
  assign n17188 = ~n17186 & n17187;
  assign n17189 = ~pi619 & ~n17182;
  assign n17190 = pi619 & n17106;
  assign n17191 = ~pi1159 & ~n17190;
  assign n17192 = ~n17189 & n17191;
  assign n17193 = ~pi648 & ~n17076;
  assign n17194 = ~n17192 & n17193;
  assign n17195 = pi789 & ~n17194;
  assign n17196 = pi789 & ~n17188;
  assign n17197 = ~n17194 & n17196;
  assign n17198 = ~n17188 & n17195;
  assign n17199 = ~pi789 & n17182;
  assign n17200 = n59242 & ~n17199;
  assign n17201 = ~n59596 & n17200;
  assign n17202 = ~n17135 & ~n17201;
  assign n17203 = ~n59357 & ~n17202;
  assign n17204 = n7957 & ~n59593;
  assign n17205 = n8065 & n17108;
  assign n17206 = pi629 & ~n17205;
  assign n17207 = ~n17204 & n17206;
  assign n17208 = n7958 & ~n59593;
  assign n17209 = n8074 & n17108;
  assign n17210 = ~pi629 & ~n17209;
  assign n17211 = ~n17208 & n17210;
  assign n17212 = pi792 & ~n17211;
  assign n17213 = ~n17208 & ~n17209;
  assign n17214 = ~pi629 & ~n17213;
  assign n17215 = ~n17204 & ~n17205;
  assign n17216 = pi629 & ~n17215;
  assign n17217 = ~n17214 & ~n17216;
  assign n17218 = pi792 & ~n17217;
  assign n17219 = pi792 & ~n17207;
  assign n17220 = ~n17211 & n17219;
  assign n17221 = ~n17207 & n17212;
  assign n17222 = ~n8108 & ~n59597;
  assign n17223 = ~n17203 & n17222;
  assign n17224 = ~n17121 & ~n17223;
  assign n17225 = pi644 & n17224;
  assign n17226 = ~pi787 & ~n17109;
  assign n17227 = pi1157 & ~n17112;
  assign n17228 = ~n17117 & ~n17227;
  assign n17229 = pi787 & ~n17228;
  assign n17230 = ~n17226 & ~n17229;
  assign n17231 = ~pi644 & n17230;
  assign n17232 = pi715 & ~n17231;
  assign n17233 = ~n17225 & n17232;
  assign n17234 = ~n11491 & n17053;
  assign n17235 = ~n7835 & n17088;
  assign n17236 = ~n7835 & ~n17091;
  assign n17237 = n7835 & n17053;
  assign n17238 = ~n17236 & ~n17237;
  assign n17239 = ~n17234 & ~n17235;
  assign n17240 = pi644 & ~n59598;
  assign n17241 = ~pi644 & n17053;
  assign n17242 = ~pi715 & ~n17241;
  assign n17243 = ~n17240 & n17242;
  assign n17244 = pi1160 & ~n17243;
  assign n17245 = ~n17233 & n17244;
  assign n17246 = ~pi644 & n17224;
  assign n17247 = pi644 & n17230;
  assign n17248 = ~pi715 & ~n17247;
  assign n17249 = ~n17246 & n17248;
  assign n17250 = ~pi644 & ~n59598;
  assign n17251 = pi644 & n17053;
  assign n17252 = pi715 & ~n17251;
  assign n17253 = ~n17250 & n17252;
  assign n17254 = ~pi1160 & ~n17253;
  assign n17255 = ~n17249 & n17254;
  assign n17256 = ~n17245 & ~n17255;
  assign n17257 = pi790 & ~n17256;
  assign n17258 = ~pi790 & n17224;
  assign n17259 = pi832 & ~n17258;
  assign n17260 = ~n17257 & n17259;
  assign n17261 = ~pi183 & ~n7560;
  assign n17262 = n59231 & ~n17261;
  assign n17263 = ~pi725 & n59132;
  assign n17264 = n17261 & ~n17263;
  assign n17265 = pi183 & n59251;
  assign n17266 = ~pi38 & ~n17265;
  assign n17267 = n59132 & ~n17266;
  assign n17268 = ~pi183 & n8249;
  assign n17269 = ~n17267 & ~n17268;
  assign n17270 = ~pi183 & ~n6863;
  assign n17271 = n7547 & ~n17270;
  assign n17272 = ~pi725 & ~n17271;
  assign n17273 = ~n17269 & n17272;
  assign n17274 = ~n17264 & ~n17273;
  assign n17275 = ~pi778 & n17274;
  assign n17276 = pi625 & ~n17274;
  assign n17277 = ~pi625 & n17261;
  assign n17278 = pi1153 & ~n17277;
  assign n17279 = ~n17276 & n17278;
  assign n17280 = ~pi625 & ~n17274;
  assign n17281 = pi625 & n17261;
  assign n17282 = ~pi1153 & ~n17281;
  assign n17283 = ~n17280 & n17282;
  assign n17284 = ~n17279 & ~n17283;
  assign n17285 = pi778 & ~n17284;
  assign n17286 = ~n17275 & ~n17285;
  assign n17287 = ~n59229 & n17286;
  assign n17288 = n59229 & n17261;
  assign n17289 = n59229 & ~n17261;
  assign n17290 = ~n59229 & ~n17286;
  assign n17291 = ~n17289 & ~n17290;
  assign n17292 = ~n17287 & ~n17288;
  assign n17293 = ~n59231 & ~n59599;
  assign n17294 = ~n59231 & n59599;
  assign n17295 = n59231 & n17261;
  assign n17296 = ~n17294 & ~n17295;
  assign n17297 = ~n17262 & ~n17293;
  assign n17298 = ~n7716 & ~n59600;
  assign n17299 = n7716 & n17261;
  assign n17300 = n7716 & ~n17261;
  assign n17301 = ~n7716 & n59600;
  assign n17302 = ~n17300 & ~n17301;
  assign n17303 = ~n17298 & ~n17299;
  assign n17304 = ~n7762 & n59601;
  assign n17305 = n7762 & n17261;
  assign n17306 = ~n17304 & ~n17305;
  assign n17307 = ~pi792 & n17306;
  assign n17308 = pi628 & ~n17306;
  assign n17309 = ~pi628 & n17261;
  assign n17310 = pi1156 & ~n17309;
  assign n17311 = ~n17308 & n17310;
  assign n17312 = ~pi628 & ~n17306;
  assign n17313 = pi628 & n17261;
  assign n17314 = ~pi1156 & ~n17313;
  assign n17315 = ~n17312 & n17314;
  assign n17316 = ~n17311 & ~n17315;
  assign n17317 = pi792 & ~n17316;
  assign n17318 = ~n17307 & ~n17317;
  assign n17319 = pi647 & n17318;
  assign n17320 = ~pi647 & n17261;
  assign n17321 = pi647 & ~n17318;
  assign n17322 = ~pi647 & ~n17261;
  assign n17323 = ~n17321 & ~n17322;
  assign n17324 = ~n17319 & ~n17320;
  assign n17325 = pi1157 & ~n59602;
  assign n17326 = ~pi647 & n17318;
  assign n17327 = pi647 & n17261;
  assign n17328 = ~pi1157 & ~n17327;
  assign n17329 = ~n17326 & n17328;
  assign n17330 = ~pi647 & ~n17318;
  assign n17331 = pi647 & ~n17261;
  assign n17332 = ~n17330 & ~n17331;
  assign n17333 = ~pi1157 & n17332;
  assign n17334 = pi1157 & n59602;
  assign n17335 = ~n17333 & ~n17334;
  assign n17336 = ~n17325 & ~n17329;
  assign n17337 = pi787 & n59603;
  assign n17338 = ~pi787 & ~n17318;
  assign n17339 = pi787 & ~n59603;
  assign n17340 = ~pi787 & n17318;
  assign n17341 = ~n17339 & ~n17340;
  assign n17342 = ~n17337 & ~n17338;
  assign n17343 = ~pi644 & ~n59604;
  assign n17344 = pi715 & ~n17343;
  assign n17345 = pi183 & ~n59132;
  assign n17346 = ~pi755 & n6865;
  assign n17347 = ~n17270 & ~n17346;
  assign n17348 = pi38 & ~n17347;
  assign n17349 = ~pi183 & n59164;
  assign n17350 = pi183 & ~n6855;
  assign n17351 = ~pi755 & ~n17350;
  assign n17352 = ~n17349 & n17351;
  assign n17353 = ~pi183 & pi755;
  assign n17354 = ~n6656 & n17353;
  assign n17355 = pi755 & ~n6656;
  assign n17356 = ~pi755 & ~n17349;
  assign n17357 = ~n17355 & ~n17356;
  assign n17358 = ~pi183 & ~n17357;
  assign n17359 = n6855 & n17356;
  assign n17360 = ~n17358 & ~n17359;
  assign n17361 = ~n17352 & ~n17354;
  assign n17362 = ~pi38 & ~n59605;
  assign n17363 = ~n17348 & ~n17362;
  assign n17364 = n59132 & n17363;
  assign n17365 = ~n17345 & ~n17364;
  assign n17366 = ~n7597 & ~n17365;
  assign n17367 = n7597 & ~n17261;
  assign n17368 = ~n17366 & ~n17367;
  assign n17369 = ~pi785 & ~n17368;
  assign n17370 = ~n7598 & ~n17261;
  assign n17371 = pi609 & n17366;
  assign n17372 = ~n17370 & ~n17371;
  assign n17373 = pi1155 & ~n17372;
  assign n17374 = ~n7610 & ~n17261;
  assign n17375 = ~pi609 & n17366;
  assign n17376 = ~n17374 & ~n17375;
  assign n17377 = ~pi1155 & ~n17376;
  assign n17378 = ~n17373 & ~n17377;
  assign n17379 = pi785 & ~n17378;
  assign n17380 = ~n17369 & ~n17379;
  assign n17381 = ~pi781 & ~n17380;
  assign n17382 = pi618 & n17380;
  assign n17383 = ~pi618 & n17261;
  assign n17384 = pi1154 & ~n17383;
  assign n17385 = ~n17382 & n17384;
  assign n17386 = ~pi618 & n17380;
  assign n17387 = pi618 & n17261;
  assign n17388 = ~pi1154 & ~n17387;
  assign n17389 = ~n17386 & n17388;
  assign n17390 = ~n17385 & ~n17389;
  assign n17391 = pi781 & ~n17390;
  assign n17392 = ~n17381 & ~n17391;
  assign n17393 = ~pi789 & ~n17392;
  assign n17394 = pi619 & n17392;
  assign n17395 = ~pi619 & n17261;
  assign n17396 = pi1159 & ~n17395;
  assign n17397 = ~n17394 & n17396;
  assign n17398 = ~pi619 & n17392;
  assign n17399 = pi619 & n17261;
  assign n17400 = ~pi1159 & ~n17399;
  assign n17401 = ~n17398 & n17400;
  assign n17402 = ~n17397 & ~n17401;
  assign n17403 = pi789 & ~n17402;
  assign n17404 = ~n17393 & ~n17403;
  assign n17405 = ~n8054 & n17404;
  assign n17406 = n8054 & n17261;
  assign n17407 = ~n17405 & ~n17406;
  assign n17408 = ~n7793 & ~n17407;
  assign n17409 = n7793 & n17261;
  assign n17410 = ~n17408 & ~n17409;
  assign n17411 = ~n7835 & ~n17410;
  assign n17412 = n7835 & n17261;
  assign n17413 = n7835 & ~n17261;
  assign n17414 = ~n7835 & n17410;
  assign n17415 = ~n17413 & ~n17414;
  assign n17416 = ~n17411 & ~n17412;
  assign n17417 = pi644 & n59606;
  assign n17418 = ~pi644 & n17261;
  assign n17419 = ~pi715 & ~n17418;
  assign n17420 = ~n17417 & n17419;
  assign n17421 = pi1160 & ~n17420;
  assign n17422 = ~n17344 & n17421;
  assign n17423 = pi644 & ~n59604;
  assign n17424 = ~pi715 & ~n17423;
  assign n17425 = ~pi644 & n59606;
  assign n17426 = pi644 & n17261;
  assign n17427 = pi715 & ~n17426;
  assign n17428 = ~n17425 & n17427;
  assign n17429 = ~pi1160 & ~n17428;
  assign n17430 = ~n17424 & n17429;
  assign n17431 = ~n17422 & ~n17430;
  assign n17432 = pi790 & ~n17431;
  assign n17433 = ~pi644 & n17429;
  assign n17434 = pi644 & n17421;
  assign n17435 = pi790 & ~n17434;
  assign n17436 = pi790 & ~n17433;
  assign n17437 = ~n17434 & n17436;
  assign n17438 = ~n17433 & n17435;
  assign n17439 = ~n7872 & n17410;
  assign n17440 = n7832 & ~n59602;
  assign n17441 = n7833 & ~n17332;
  assign n17442 = pi630 & n17329;
  assign n17443 = ~n17440 & ~n59608;
  assign n17444 = ~n17439 & n17443;
  assign n17445 = pi787 & ~n17444;
  assign n17446 = ~n11154 & n17407;
  assign n17447 = ~pi629 & n17311;
  assign n17448 = pi629 & n17315;
  assign n17449 = ~n17447 & ~n17448;
  assign n17450 = ~n17446 & n17449;
  assign n17451 = pi792 & ~n17450;
  assign n17452 = pi725 & ~n17363;
  assign n17453 = ~pi183 & n59177;
  assign n17454 = pi183 & n7111;
  assign n17455 = pi755 & ~n17454;
  assign n17456 = ~n17453 & n17455;
  assign n17457 = pi183 & n7188;
  assign n17458 = ~pi183 & ~n59203;
  assign n17459 = ~pi755 & ~n17458;
  assign n17460 = ~n17457 & n17459;
  assign n17461 = pi39 & ~n17460;
  assign n17462 = ~n17456 & n17461;
  assign n17463 = pi183 & n7333;
  assign n17464 = ~pi183 & n7310;
  assign n17465 = pi755 & ~n17464;
  assign n17466 = ~n17463 & n17465;
  assign n17467 = ~pi183 & ~n7339;
  assign n17468 = pi183 & ~n7347;
  assign n17469 = ~pi755 & ~n17468;
  assign n17470 = ~n17467 & n17469;
  assign n17471 = ~pi39 & ~n17470;
  assign n17472 = pi183 & ~n7333;
  assign n17473 = ~pi183 & ~n7310;
  assign n17474 = pi755 & ~n17473;
  assign n17475 = pi755 & ~n17472;
  assign n17476 = ~n17473 & n17475;
  assign n17477 = ~n17472 & n17474;
  assign n17478 = ~pi183 & n7339;
  assign n17479 = pi183 & n7347;
  assign n17480 = ~pi755 & ~n17479;
  assign n17481 = ~n17478 & n17480;
  assign n17482 = ~n59609 & ~n17481;
  assign n17483 = ~pi39 & ~n17482;
  assign n17484 = ~n17466 & n17471;
  assign n17485 = ~pi38 & ~n59610;
  assign n17486 = ~n17462 & n17485;
  assign n17487 = ~pi755 & ~n7222;
  assign n17488 = n9794 & ~n17487;
  assign n17489 = ~pi183 & ~n17488;
  assign n17490 = ~n7056 & ~n17054;
  assign n17491 = pi183 & ~n17490;
  assign n17492 = n59171 & n17491;
  assign n17493 = pi38 & ~n17492;
  assign n17494 = ~n17489 & n17493;
  assign n17495 = ~pi725 & ~n17494;
  assign n17496 = ~n17486 & n17495;
  assign n17497 = n59132 & ~n17496;
  assign n17498 = ~n17452 & n17497;
  assign n17499 = ~n17345 & ~n17498;
  assign n17500 = ~pi625 & n17499;
  assign n17501 = pi625 & n17365;
  assign n17502 = ~pi1153 & ~n17501;
  assign n17503 = ~n17500 & n17502;
  assign n17504 = ~pi608 & ~n17279;
  assign n17505 = ~n17503 & n17504;
  assign n17506 = pi625 & n17499;
  assign n17507 = ~pi625 & n17365;
  assign n17508 = pi1153 & ~n17507;
  assign n17509 = ~n17506 & n17508;
  assign n17510 = pi608 & ~n17283;
  assign n17511 = ~n17509 & n17510;
  assign n17512 = ~n17505 & ~n17511;
  assign n17513 = pi778 & ~n17512;
  assign n17514 = ~pi778 & n17499;
  assign n17515 = ~n17513 & ~n17514;
  assign n17516 = ~pi609 & ~n17515;
  assign n17517 = pi609 & n17286;
  assign n17518 = ~pi1155 & ~n17517;
  assign n17519 = ~n17516 & n17518;
  assign n17520 = ~pi660 & ~n17373;
  assign n17521 = ~n17519 & n17520;
  assign n17522 = pi609 & ~n17515;
  assign n17523 = ~pi609 & n17286;
  assign n17524 = pi1155 & ~n17523;
  assign n17525 = ~n17522 & n17524;
  assign n17526 = pi660 & ~n17377;
  assign n17527 = ~n17525 & n17526;
  assign n17528 = ~n17521 & ~n17527;
  assign n17529 = pi785 & ~n17528;
  assign n17530 = ~pi785 & ~n17515;
  assign n17531 = ~n17529 & ~n17530;
  assign n17532 = ~pi618 & ~n17531;
  assign n17533 = pi618 & n59599;
  assign n17534 = ~pi1154 & ~n17533;
  assign n17535 = ~n17532 & n17534;
  assign n17536 = ~pi627 & ~n17385;
  assign n17537 = ~n17535 & n17536;
  assign n17538 = pi618 & ~n17531;
  assign n17539 = ~pi618 & n59599;
  assign n17540 = pi1154 & ~n17539;
  assign n17541 = ~n17538 & n17540;
  assign n17542 = pi627 & ~n17389;
  assign n17543 = ~n17541 & n17542;
  assign n17544 = ~n17537 & ~n17543;
  assign n17545 = pi781 & ~n17544;
  assign n17546 = ~pi781 & ~n17531;
  assign n17547 = ~n17545 & ~n17546;
  assign n17548 = pi619 & ~n17547;
  assign n17549 = ~pi619 & ~n59600;
  assign n17550 = pi1159 & ~n17549;
  assign n17551 = ~n17548 & n17550;
  assign n17552 = pi648 & ~n17401;
  assign n17553 = ~n17551 & n17552;
  assign n17554 = ~pi619 & ~n17547;
  assign n17555 = pi619 & ~n59600;
  assign n17556 = ~pi1159 & ~n17555;
  assign n17557 = ~n17554 & n17556;
  assign n17558 = ~pi648 & ~n17397;
  assign n17559 = ~n17557 & n17558;
  assign n17560 = pi789 & ~n17559;
  assign n17561 = pi789 & ~n17553;
  assign n17562 = ~n17559 & n17561;
  assign n17563 = ~n17553 & n17560;
  assign n17564 = ~pi789 & n17547;
  assign n17565 = n59242 & ~n17564;
  assign n17566 = ~n59611 & n17565;
  assign n17567 = ~pi626 & ~n17404;
  assign n17568 = pi626 & ~n17261;
  assign n17569 = n7760 & ~n17568;
  assign n17570 = ~n17567 & n17569;
  assign n17571 = n7984 & n59601;
  assign n17572 = pi626 & ~n17404;
  assign n17573 = ~pi626 & ~n17261;
  assign n17574 = n7759 & ~n17573;
  assign n17575 = ~n17572 & n17574;
  assign n17576 = ~n17571 & ~n17575;
  assign n17577 = ~n17570 & ~n17571;
  assign n17578 = ~n17575 & n17577;
  assign n17579 = ~n17570 & n17576;
  assign n17580 = pi788 & ~n59612;
  assign n17581 = ~n59357 & ~n17580;
  assign n17582 = ~n17566 & n17581;
  assign n17583 = ~n17451 & ~n17582;
  assign n17584 = ~n8108 & ~n17583;
  assign n17585 = ~n17445 & ~n17584;
  assign n17586 = ~n59607 & n17585;
  assign n17587 = ~n17432 & ~n17586;
  assign n17588 = n58992 & ~n17587;
  assign n17589 = ~pi183 & ~n58992;
  assign n17590 = ~pi832 & ~n17589;
  assign n17591 = ~n17588 & n17590;
  assign po340 = ~n17260 & ~n17591;
  assign n17593 = ~pi184 & ~n2794;
  assign n17594 = ~pi777 & n6822;
  assign n17595 = ~n17593 & ~n17594;
  assign n17596 = ~n7875 & ~n17595;
  assign n17597 = ~pi785 & ~n17596;
  assign n17598 = n7610 & n17594;
  assign n17599 = n17596 & ~n17598;
  assign n17600 = pi1155 & ~n17599;
  assign n17601 = ~pi1155 & ~n17593;
  assign n17602 = ~n17598 & n17601;
  assign n17603 = ~n17600 & ~n17602;
  assign n17604 = pi785 & ~n17603;
  assign n17605 = ~n17597 & ~n17604;
  assign n17606 = ~pi781 & ~n17605;
  assign n17607 = ~n7890 & n17605;
  assign n17608 = pi1154 & ~n17607;
  assign n17609 = ~n7893 & n17605;
  assign n17610 = ~pi1154 & ~n17609;
  assign n17611 = ~n17608 & ~n17610;
  assign n17612 = pi781 & ~n17611;
  assign n17613 = ~n17606 & ~n17612;
  assign n17614 = ~pi789 & ~n17613;
  assign n17615 = ~n11882 & n17613;
  assign n17616 = pi1159 & ~n17615;
  assign n17617 = ~n11885 & n17613;
  assign n17618 = ~pi1159 & ~n17617;
  assign n17619 = ~n17616 & ~n17618;
  assign n17620 = pi789 & ~n17619;
  assign n17621 = ~n17614 & ~n17620;
  assign n17622 = ~n8054 & ~n17621;
  assign n17623 = n8054 & ~n17593;
  assign n17624 = ~n8054 & n17621;
  assign n17625 = n8054 & n17593;
  assign n17626 = ~n17624 & ~n17625;
  assign n17627 = ~n17622 & ~n17623;
  assign n17628 = ~n7793 & ~n59613;
  assign n17629 = n7793 & n17593;
  assign n17630 = ~n7872 & ~n17629;
  assign n17631 = ~n17628 & ~n17629;
  assign n17632 = ~n7872 & n17631;
  assign n17633 = ~n17628 & n17630;
  assign n17634 = ~pi737 & n7055;
  assign n17635 = ~n17593 & ~n17634;
  assign n17636 = ~pi778 & ~n17635;
  assign n17637 = ~pi625 & n17634;
  assign n17638 = ~n17635 & ~n17637;
  assign n17639 = pi1153 & ~n17638;
  assign n17640 = ~pi1153 & ~n17593;
  assign n17641 = ~n17637 & n17640;
  assign n17642 = pi778 & ~n17641;
  assign n17643 = ~n17639 & n17642;
  assign n17644 = ~n17636 & ~n17643;
  assign n17645 = ~n7949 & ~n17644;
  assign n17646 = ~n7951 & n17645;
  assign n17647 = ~n7953 & n17646;
  assign n17648 = ~n7955 & n17647;
  assign n17649 = ~n7967 & n17648;
  assign n17650 = pi647 & ~n17649;
  assign n17651 = ~pi647 & ~n17593;
  assign n17652 = ~n17650 & ~n17651;
  assign n17653 = n7832 & ~n17652;
  assign n17654 = ~pi647 & n17649;
  assign n17655 = pi647 & n17593;
  assign n17656 = ~pi1157 & ~n17655;
  assign n17657 = ~n17654 & n17656;
  assign n17658 = pi630 & n17657;
  assign n17659 = ~n17653 & ~n17658;
  assign n17660 = ~n59614 & n17659;
  assign n17661 = pi787 & ~n17660;
  assign n17662 = ~pi626 & ~n17621;
  assign n17663 = pi626 & ~n17593;
  assign n17664 = n7760 & ~n17663;
  assign n17665 = ~n17662 & n17664;
  assign n17666 = n7984 & n17647;
  assign n17667 = pi626 & ~n17621;
  assign n17668 = ~pi626 & ~n17593;
  assign n17669 = n7759 & ~n17668;
  assign n17670 = ~n17667 & n17669;
  assign n17671 = ~n17666 & ~n17670;
  assign n17672 = ~n17665 & ~n17666;
  assign n17673 = ~n17670 & n17672;
  assign n17674 = ~n17665 & n17671;
  assign n17675 = pi788 & ~n59615;
  assign n17676 = ~n6701 & ~n17635;
  assign n17677 = pi625 & n17676;
  assign n17678 = n17595 & ~n17676;
  assign n17679 = ~n17677 & ~n17678;
  assign n17680 = n17640 & ~n17679;
  assign n17681 = ~pi608 & ~n17639;
  assign n17682 = ~n17680 & n17681;
  assign n17683 = pi1153 & n17595;
  assign n17684 = ~n17677 & n17683;
  assign n17685 = pi608 & ~n17641;
  assign n17686 = ~n17684 & n17685;
  assign n17687 = ~n17682 & ~n17686;
  assign n17688 = pi778 & ~n17687;
  assign n17689 = ~pi778 & ~n17678;
  assign n17690 = ~n17688 & ~n17689;
  assign n17691 = ~pi609 & ~n17690;
  assign n17692 = pi609 & ~n17644;
  assign n17693 = ~pi1155 & ~n17692;
  assign n17694 = ~n17691 & n17693;
  assign n17695 = ~pi660 & ~n17600;
  assign n17696 = ~n17694 & n17695;
  assign n17697 = pi609 & ~n17690;
  assign n17698 = ~pi609 & ~n17644;
  assign n17699 = pi1155 & ~n17698;
  assign n17700 = ~n17697 & n17699;
  assign n17701 = pi660 & ~n17602;
  assign n17702 = ~n17700 & n17701;
  assign n17703 = ~n17696 & ~n17702;
  assign n17704 = pi785 & ~n17703;
  assign n17705 = ~pi785 & ~n17690;
  assign n17706 = ~n17704 & ~n17705;
  assign n17707 = ~pi618 & ~n17706;
  assign n17708 = pi618 & n17645;
  assign n17709 = ~pi1154 & ~n17708;
  assign n17710 = ~n17707 & n17709;
  assign n17711 = ~pi627 & ~n17608;
  assign n17712 = ~n17710 & n17711;
  assign n17713 = pi618 & ~n17706;
  assign n17714 = ~pi618 & n17645;
  assign n17715 = pi1154 & ~n17714;
  assign n17716 = ~n17713 & n17715;
  assign n17717 = pi627 & ~n17610;
  assign n17718 = ~n17716 & n17717;
  assign n17719 = ~n17712 & ~n17718;
  assign n17720 = pi781 & ~n17719;
  assign n17721 = ~pi781 & ~n17706;
  assign n17722 = ~n17720 & ~n17721;
  assign n17723 = pi619 & ~n17722;
  assign n17724 = ~pi619 & n17646;
  assign n17725 = pi1159 & ~n17724;
  assign n17726 = ~n17723 & n17725;
  assign n17727 = pi648 & ~n17618;
  assign n17728 = ~n17726 & n17727;
  assign n17729 = ~pi619 & ~n17722;
  assign n17730 = pi619 & n17646;
  assign n17731 = ~pi1159 & ~n17730;
  assign n17732 = ~n17729 & n17731;
  assign n17733 = ~pi648 & ~n17616;
  assign n17734 = ~n17732 & n17733;
  assign n17735 = pi789 & ~n17734;
  assign n17736 = pi789 & ~n17728;
  assign n17737 = ~n17734 & n17736;
  assign n17738 = ~n17728 & n17735;
  assign n17739 = ~pi789 & n17722;
  assign n17740 = n59242 & ~n17739;
  assign n17741 = ~n59616 & n17740;
  assign n17742 = ~n17675 & ~n17741;
  assign n17743 = ~n59357 & ~n17742;
  assign n17744 = n7957 & ~n59613;
  assign n17745 = n8065 & n17648;
  assign n17746 = pi629 & ~n17745;
  assign n17747 = ~n17744 & n17746;
  assign n17748 = n7958 & ~n59613;
  assign n17749 = n8074 & n17648;
  assign n17750 = ~pi629 & ~n17749;
  assign n17751 = ~n17748 & n17750;
  assign n17752 = pi792 & ~n17751;
  assign n17753 = ~n17748 & ~n17749;
  assign n17754 = ~pi629 & ~n17753;
  assign n17755 = ~n17744 & ~n17745;
  assign n17756 = pi629 & ~n17755;
  assign n17757 = ~n17754 & ~n17756;
  assign n17758 = pi792 & ~n17757;
  assign n17759 = pi792 & ~n17747;
  assign n17760 = ~n17751 & n17759;
  assign n17761 = ~n17747 & n17752;
  assign n17762 = ~n8108 & ~n59617;
  assign n17763 = ~n17743 & n17762;
  assign n17764 = ~n17661 & ~n17763;
  assign n17765 = pi644 & n17764;
  assign n17766 = ~pi787 & ~n17649;
  assign n17767 = pi1157 & ~n17652;
  assign n17768 = ~n17657 & ~n17767;
  assign n17769 = pi787 & ~n17768;
  assign n17770 = ~n17766 & ~n17769;
  assign n17771 = ~pi644 & n17770;
  assign n17772 = pi715 & ~n17771;
  assign n17773 = ~n17765 & n17772;
  assign n17774 = ~n11491 & n17593;
  assign n17775 = ~n7835 & n17628;
  assign n17776 = ~n7835 & ~n17631;
  assign n17777 = n7835 & n17593;
  assign n17778 = ~n17776 & ~n17777;
  assign n17779 = ~n17774 & ~n17775;
  assign n17780 = pi644 & ~n59618;
  assign n17781 = ~pi644 & n17593;
  assign n17782 = ~pi715 & ~n17781;
  assign n17783 = ~n17780 & n17782;
  assign n17784 = pi1160 & ~n17783;
  assign n17785 = ~n17773 & n17784;
  assign n17786 = ~pi644 & n17764;
  assign n17787 = pi644 & n17770;
  assign n17788 = ~pi715 & ~n17787;
  assign n17789 = ~n17786 & n17788;
  assign n17790 = ~pi644 & ~n59618;
  assign n17791 = pi644 & n17593;
  assign n17792 = pi715 & ~n17791;
  assign n17793 = ~n17790 & n17792;
  assign n17794 = ~pi1160 & ~n17793;
  assign n17795 = ~n17789 & n17794;
  assign n17796 = ~n17785 & ~n17795;
  assign n17797 = pi790 & ~n17796;
  assign n17798 = ~pi790 & n17764;
  assign n17799 = pi832 & ~n17798;
  assign n17800 = ~n17797 & n17799;
  assign n17801 = ~pi184 & ~n7560;
  assign n17802 = n59231 & ~n17801;
  assign n17803 = ~pi737 & n59132;
  assign n17804 = n17801 & ~n17803;
  assign n17805 = pi184 & n59251;
  assign n17806 = ~pi38 & ~n17805;
  assign n17807 = n59132 & ~n17806;
  assign n17808 = ~pi184 & n8249;
  assign n17809 = ~n17807 & ~n17808;
  assign n17810 = ~pi184 & ~n6863;
  assign n17811 = n7547 & ~n17810;
  assign n17812 = ~pi737 & ~n17811;
  assign n17813 = ~n17809 & n17812;
  assign n17814 = ~n17804 & ~n17813;
  assign n17815 = ~pi778 & n17814;
  assign n17816 = pi625 & ~n17814;
  assign n17817 = ~pi625 & n17801;
  assign n17818 = pi1153 & ~n17817;
  assign n17819 = ~n17816 & n17818;
  assign n17820 = ~pi625 & ~n17814;
  assign n17821 = pi625 & n17801;
  assign n17822 = ~pi1153 & ~n17821;
  assign n17823 = ~n17820 & n17822;
  assign n17824 = ~n17819 & ~n17823;
  assign n17825 = pi778 & ~n17824;
  assign n17826 = ~n17815 & ~n17825;
  assign n17827 = ~n59229 & n17826;
  assign n17828 = n59229 & n17801;
  assign n17829 = n59229 & ~n17801;
  assign n17830 = ~n59229 & ~n17826;
  assign n17831 = ~n17829 & ~n17830;
  assign n17832 = ~n17827 & ~n17828;
  assign n17833 = ~n59231 & ~n59619;
  assign n17834 = ~n59231 & n59619;
  assign n17835 = n59231 & n17801;
  assign n17836 = ~n17834 & ~n17835;
  assign n17837 = ~n17802 & ~n17833;
  assign n17838 = ~n7716 & ~n59620;
  assign n17839 = n7716 & n17801;
  assign n17840 = n7716 & ~n17801;
  assign n17841 = ~n7716 & n59620;
  assign n17842 = ~n17840 & ~n17841;
  assign n17843 = ~n17838 & ~n17839;
  assign n17844 = ~n7762 & n59621;
  assign n17845 = n7762 & n17801;
  assign n17846 = ~n17844 & ~n17845;
  assign n17847 = ~pi792 & n17846;
  assign n17848 = pi628 & ~n17846;
  assign n17849 = ~pi628 & n17801;
  assign n17850 = pi1156 & ~n17849;
  assign n17851 = ~n17848 & n17850;
  assign n17852 = ~pi628 & ~n17846;
  assign n17853 = pi628 & n17801;
  assign n17854 = ~pi1156 & ~n17853;
  assign n17855 = ~n17852 & n17854;
  assign n17856 = ~n17851 & ~n17855;
  assign n17857 = pi792 & ~n17856;
  assign n17858 = ~n17847 & ~n17857;
  assign n17859 = pi647 & n17858;
  assign n17860 = ~pi647 & n17801;
  assign n17861 = pi647 & ~n17858;
  assign n17862 = ~pi647 & ~n17801;
  assign n17863 = ~n17861 & ~n17862;
  assign n17864 = ~n17859 & ~n17860;
  assign n17865 = pi1157 & ~n59622;
  assign n17866 = ~pi647 & n17858;
  assign n17867 = pi647 & n17801;
  assign n17868 = ~pi1157 & ~n17867;
  assign n17869 = ~n17866 & n17868;
  assign n17870 = ~pi647 & ~n17858;
  assign n17871 = pi647 & ~n17801;
  assign n17872 = ~n17870 & ~n17871;
  assign n17873 = ~pi1157 & n17872;
  assign n17874 = pi1157 & n59622;
  assign n17875 = ~n17873 & ~n17874;
  assign n17876 = ~n17865 & ~n17869;
  assign n17877 = pi787 & n59623;
  assign n17878 = ~pi787 & ~n17858;
  assign n17879 = pi787 & ~n59623;
  assign n17880 = ~pi787 & n17858;
  assign n17881 = ~n17879 & ~n17880;
  assign n17882 = ~n17877 & ~n17878;
  assign n17883 = ~pi644 & ~n59624;
  assign n17884 = pi715 & ~n17883;
  assign n17885 = pi184 & ~n59132;
  assign n17886 = ~pi777 & n6865;
  assign n17887 = ~n17810 & ~n17886;
  assign n17888 = pi38 & ~n17887;
  assign n17889 = ~pi184 & n59164;
  assign n17890 = pi184 & ~n6855;
  assign n17891 = ~pi777 & ~n17890;
  assign n17892 = ~n17889 & n17891;
  assign n17893 = ~pi184 & pi777;
  assign n17894 = ~n6656 & n17893;
  assign n17895 = pi777 & ~n6656;
  assign n17896 = ~pi777 & ~n17889;
  assign n17897 = ~n17895 & ~n17896;
  assign n17898 = ~pi184 & ~n17897;
  assign n17899 = n6855 & n17896;
  assign n17900 = ~n17898 & ~n17899;
  assign n17901 = ~n17892 & ~n17894;
  assign n17902 = ~pi38 & ~n59625;
  assign n17903 = ~n17888 & ~n17902;
  assign n17904 = n59132 & n17903;
  assign n17905 = ~n17885 & ~n17904;
  assign n17906 = ~n7597 & ~n17905;
  assign n17907 = n7597 & ~n17801;
  assign n17908 = ~n17906 & ~n17907;
  assign n17909 = ~pi785 & ~n17908;
  assign n17910 = ~n7598 & ~n17801;
  assign n17911 = pi609 & n17906;
  assign n17912 = ~n17910 & ~n17911;
  assign n17913 = pi1155 & ~n17912;
  assign n17914 = ~n7610 & ~n17801;
  assign n17915 = ~pi609 & n17906;
  assign n17916 = ~n17914 & ~n17915;
  assign n17917 = ~pi1155 & ~n17916;
  assign n17918 = ~n17913 & ~n17917;
  assign n17919 = pi785 & ~n17918;
  assign n17920 = ~n17909 & ~n17919;
  assign n17921 = ~pi781 & ~n17920;
  assign n17922 = pi618 & n17920;
  assign n17923 = ~pi618 & n17801;
  assign n17924 = pi1154 & ~n17923;
  assign n17925 = ~n17922 & n17924;
  assign n17926 = ~pi618 & n17920;
  assign n17927 = pi618 & n17801;
  assign n17928 = ~pi1154 & ~n17927;
  assign n17929 = ~n17926 & n17928;
  assign n17930 = ~n17925 & ~n17929;
  assign n17931 = pi781 & ~n17930;
  assign n17932 = ~n17921 & ~n17931;
  assign n17933 = ~pi789 & ~n17932;
  assign n17934 = pi619 & n17932;
  assign n17935 = ~pi619 & n17801;
  assign n17936 = pi1159 & ~n17935;
  assign n17937 = ~n17934 & n17936;
  assign n17938 = ~pi619 & n17932;
  assign n17939 = pi619 & n17801;
  assign n17940 = ~pi1159 & ~n17939;
  assign n17941 = ~n17938 & n17940;
  assign n17942 = ~n17937 & ~n17941;
  assign n17943 = pi789 & ~n17942;
  assign n17944 = ~n17933 & ~n17943;
  assign n17945 = ~n8054 & n17944;
  assign n17946 = n8054 & n17801;
  assign n17947 = ~n17945 & ~n17946;
  assign n17948 = ~n7793 & ~n17947;
  assign n17949 = n7793 & n17801;
  assign n17950 = ~n17948 & ~n17949;
  assign n17951 = ~n7835 & ~n17950;
  assign n17952 = n7835 & n17801;
  assign n17953 = n7835 & ~n17801;
  assign n17954 = ~n7835 & n17950;
  assign n17955 = ~n17953 & ~n17954;
  assign n17956 = ~n17951 & ~n17952;
  assign n17957 = pi644 & n59626;
  assign n17958 = ~pi644 & n17801;
  assign n17959 = ~pi715 & ~n17958;
  assign n17960 = ~n17957 & n17959;
  assign n17961 = pi1160 & ~n17960;
  assign n17962 = ~n17884 & n17961;
  assign n17963 = pi644 & ~n59624;
  assign n17964 = ~pi715 & ~n17963;
  assign n17965 = ~pi644 & n59626;
  assign n17966 = pi644 & n17801;
  assign n17967 = pi715 & ~n17966;
  assign n17968 = ~n17965 & n17967;
  assign n17969 = ~pi1160 & ~n17968;
  assign n17970 = ~n17964 & n17969;
  assign n17971 = ~n17962 & ~n17970;
  assign n17972 = pi790 & ~n17971;
  assign n17973 = ~pi644 & n17969;
  assign n17974 = pi644 & n17961;
  assign n17975 = pi790 & ~n17974;
  assign n17976 = pi790 & ~n17973;
  assign n17977 = ~n17974 & n17976;
  assign n17978 = ~n17973 & n17975;
  assign n17979 = ~n7872 & n17950;
  assign n17980 = n7832 & ~n59622;
  assign n17981 = n7833 & ~n17872;
  assign n17982 = pi630 & n17869;
  assign n17983 = ~n17980 & ~n59628;
  assign n17984 = ~n17979 & n17983;
  assign n17985 = pi787 & ~n17984;
  assign n17986 = ~n11154 & n17947;
  assign n17987 = ~pi629 & n17851;
  assign n17988 = pi629 & n17855;
  assign n17989 = ~n17987 & ~n17988;
  assign n17990 = ~n17986 & n17989;
  assign n17991 = pi792 & ~n17990;
  assign n17992 = pi737 & ~n17903;
  assign n17993 = ~pi184 & n59177;
  assign n17994 = pi184 & n7111;
  assign n17995 = pi777 & ~n17994;
  assign n17996 = ~n17993 & n17995;
  assign n17997 = pi184 & n7188;
  assign n17998 = ~pi184 & ~n59203;
  assign n17999 = ~pi777 & ~n17998;
  assign n18000 = ~n17997 & n17999;
  assign n18001 = pi39 & ~n18000;
  assign n18002 = ~n17996 & n18001;
  assign n18003 = pi184 & n7333;
  assign n18004 = ~pi184 & n7310;
  assign n18005 = pi777 & ~n18004;
  assign n18006 = ~n18003 & n18005;
  assign n18007 = ~pi184 & ~n7339;
  assign n18008 = pi184 & ~n7347;
  assign n18009 = ~pi777 & ~n18008;
  assign n18010 = ~n18007 & n18009;
  assign n18011 = ~pi39 & ~n18010;
  assign n18012 = pi184 & ~n7333;
  assign n18013 = ~pi184 & ~n7310;
  assign n18014 = pi777 & ~n18013;
  assign n18015 = pi777 & ~n18012;
  assign n18016 = ~n18013 & n18015;
  assign n18017 = ~n18012 & n18014;
  assign n18018 = ~pi184 & n7339;
  assign n18019 = pi184 & n7347;
  assign n18020 = ~pi777 & ~n18019;
  assign n18021 = ~n18018 & n18020;
  assign n18022 = ~n59629 & ~n18021;
  assign n18023 = ~pi39 & ~n18022;
  assign n18024 = ~n18006 & n18011;
  assign n18025 = ~pi38 & ~n59630;
  assign n18026 = ~n18002 & n18025;
  assign n18027 = ~pi777 & ~n7222;
  assign n18028 = n9794 & ~n18027;
  assign n18029 = ~pi184 & ~n18028;
  assign n18030 = ~n7056 & ~n17594;
  assign n18031 = pi184 & ~n18030;
  assign n18032 = n59171 & n18031;
  assign n18033 = pi38 & ~n18032;
  assign n18034 = ~n18029 & n18033;
  assign n18035 = ~pi737 & ~n18034;
  assign n18036 = ~n18026 & n18035;
  assign n18037 = n59132 & ~n18036;
  assign n18038 = ~n17992 & n18037;
  assign n18039 = ~n17885 & ~n18038;
  assign n18040 = ~pi625 & n18039;
  assign n18041 = pi625 & n17905;
  assign n18042 = ~pi1153 & ~n18041;
  assign n18043 = ~n18040 & n18042;
  assign n18044 = ~pi608 & ~n17819;
  assign n18045 = ~n18043 & n18044;
  assign n18046 = pi625 & n18039;
  assign n18047 = ~pi625 & n17905;
  assign n18048 = pi1153 & ~n18047;
  assign n18049 = ~n18046 & n18048;
  assign n18050 = pi608 & ~n17823;
  assign n18051 = ~n18049 & n18050;
  assign n18052 = ~n18045 & ~n18051;
  assign n18053 = pi778 & ~n18052;
  assign n18054 = ~pi778 & n18039;
  assign n18055 = ~n18053 & ~n18054;
  assign n18056 = ~pi609 & ~n18055;
  assign n18057 = pi609 & n17826;
  assign n18058 = ~pi1155 & ~n18057;
  assign n18059 = ~n18056 & n18058;
  assign n18060 = ~pi660 & ~n17913;
  assign n18061 = ~n18059 & n18060;
  assign n18062 = pi609 & ~n18055;
  assign n18063 = ~pi609 & n17826;
  assign n18064 = pi1155 & ~n18063;
  assign n18065 = ~n18062 & n18064;
  assign n18066 = pi660 & ~n17917;
  assign n18067 = ~n18065 & n18066;
  assign n18068 = ~n18061 & ~n18067;
  assign n18069 = pi785 & ~n18068;
  assign n18070 = ~pi785 & ~n18055;
  assign n18071 = ~n18069 & ~n18070;
  assign n18072 = ~pi618 & ~n18071;
  assign n18073 = pi618 & n59619;
  assign n18074 = ~pi1154 & ~n18073;
  assign n18075 = ~n18072 & n18074;
  assign n18076 = ~pi627 & ~n17925;
  assign n18077 = ~n18075 & n18076;
  assign n18078 = pi618 & ~n18071;
  assign n18079 = ~pi618 & n59619;
  assign n18080 = pi1154 & ~n18079;
  assign n18081 = ~n18078 & n18080;
  assign n18082 = pi627 & ~n17929;
  assign n18083 = ~n18081 & n18082;
  assign n18084 = ~n18077 & ~n18083;
  assign n18085 = pi781 & ~n18084;
  assign n18086 = ~pi781 & ~n18071;
  assign n18087 = ~n18085 & ~n18086;
  assign n18088 = pi619 & ~n18087;
  assign n18089 = ~pi619 & ~n59620;
  assign n18090 = pi1159 & ~n18089;
  assign n18091 = ~n18088 & n18090;
  assign n18092 = pi648 & ~n17941;
  assign n18093 = ~n18091 & n18092;
  assign n18094 = ~pi619 & ~n18087;
  assign n18095 = pi619 & ~n59620;
  assign n18096 = ~pi1159 & ~n18095;
  assign n18097 = ~n18094 & n18096;
  assign n18098 = ~pi648 & ~n17937;
  assign n18099 = ~n18097 & n18098;
  assign n18100 = pi789 & ~n18099;
  assign n18101 = pi789 & ~n18093;
  assign n18102 = ~n18099 & n18101;
  assign n18103 = ~n18093 & n18100;
  assign n18104 = ~pi789 & n18087;
  assign n18105 = n59242 & ~n18104;
  assign n18106 = ~n59631 & n18105;
  assign n18107 = ~pi626 & ~n17944;
  assign n18108 = pi626 & ~n17801;
  assign n18109 = n7760 & ~n18108;
  assign n18110 = ~n18107 & n18109;
  assign n18111 = n7984 & n59621;
  assign n18112 = pi626 & ~n17944;
  assign n18113 = ~pi626 & ~n17801;
  assign n18114 = n7759 & ~n18113;
  assign n18115 = ~n18112 & n18114;
  assign n18116 = ~n18111 & ~n18115;
  assign n18117 = ~n18110 & ~n18111;
  assign n18118 = ~n18115 & n18117;
  assign n18119 = ~n18110 & n18116;
  assign n18120 = pi788 & ~n59632;
  assign n18121 = ~n59357 & ~n18120;
  assign n18122 = ~n18106 & n18121;
  assign n18123 = ~n17991 & ~n18122;
  assign n18124 = ~n8108 & ~n18123;
  assign n18125 = ~n17985 & ~n18124;
  assign n18126 = ~n59627 & n18125;
  assign n18127 = ~n17972 & ~n18126;
  assign n18128 = n58992 & ~n18127;
  assign n18129 = ~pi184 & ~n58992;
  assign n18130 = ~pi832 & ~n18129;
  assign n18131 = ~n18128 & n18130;
  assign po341 = ~n17800 & ~n18131;
  assign n18133 = ~pi185 & ~n2794;
  assign n18134 = ~pi751 & n6822;
  assign n18135 = ~n18133 & ~n18134;
  assign n18136 = ~n7875 & ~n18135;
  assign n18137 = ~pi785 & ~n18136;
  assign n18138 = n7610 & n18134;
  assign n18139 = n18136 & ~n18138;
  assign n18140 = pi1155 & ~n18139;
  assign n18141 = ~pi1155 & ~n18133;
  assign n18142 = ~n18138 & n18141;
  assign n18143 = ~n18140 & ~n18142;
  assign n18144 = pi785 & ~n18143;
  assign n18145 = ~n18137 & ~n18144;
  assign n18146 = ~pi781 & ~n18145;
  assign n18147 = ~n7890 & n18145;
  assign n18148 = pi1154 & ~n18147;
  assign n18149 = ~n7893 & n18145;
  assign n18150 = ~pi1154 & ~n18149;
  assign n18151 = ~n18148 & ~n18150;
  assign n18152 = pi781 & ~n18151;
  assign n18153 = ~n18146 & ~n18152;
  assign n18154 = ~pi789 & ~n18153;
  assign n18155 = ~n11882 & n18153;
  assign n18156 = pi1159 & ~n18155;
  assign n18157 = ~n11885 & n18153;
  assign n18158 = ~pi1159 & ~n18157;
  assign n18159 = ~n18156 & ~n18158;
  assign n18160 = pi789 & ~n18159;
  assign n18161 = ~n18154 & ~n18160;
  assign n18162 = ~n8054 & ~n18161;
  assign n18163 = n8054 & ~n18133;
  assign n18164 = ~n8054 & n18161;
  assign n18165 = n8054 & n18133;
  assign n18166 = ~n18164 & ~n18165;
  assign n18167 = ~n18162 & ~n18163;
  assign n18168 = ~n7793 & ~n59633;
  assign n18169 = n7793 & n18133;
  assign n18170 = ~n7872 & ~n18169;
  assign n18171 = ~n18168 & ~n18169;
  assign n18172 = ~n7872 & n18171;
  assign n18173 = ~n18168 & n18170;
  assign n18174 = ~pi701 & n7055;
  assign n18175 = ~n18133 & ~n18174;
  assign n18176 = ~pi778 & ~n18175;
  assign n18177 = ~pi625 & n18174;
  assign n18178 = ~n18175 & ~n18177;
  assign n18179 = pi1153 & ~n18178;
  assign n18180 = ~pi1153 & ~n18133;
  assign n18181 = ~n18177 & n18180;
  assign n18182 = pi778 & ~n18181;
  assign n18183 = ~n18179 & n18182;
  assign n18184 = ~n18176 & ~n18183;
  assign n18185 = ~n7949 & ~n18184;
  assign n18186 = ~n7951 & n18185;
  assign n18187 = ~n7953 & n18186;
  assign n18188 = ~n7955 & n18187;
  assign n18189 = ~n7967 & n18188;
  assign n18190 = pi647 & ~n18189;
  assign n18191 = ~pi647 & ~n18133;
  assign n18192 = ~n18190 & ~n18191;
  assign n18193 = n7832 & ~n18192;
  assign n18194 = ~pi647 & n18189;
  assign n18195 = pi647 & n18133;
  assign n18196 = ~pi1157 & ~n18195;
  assign n18197 = ~n18194 & n18196;
  assign n18198 = pi630 & n18197;
  assign n18199 = ~n18193 & ~n18198;
  assign n18200 = ~n59634 & n18199;
  assign n18201 = pi787 & ~n18200;
  assign n18202 = ~pi626 & ~n18161;
  assign n18203 = pi626 & ~n18133;
  assign n18204 = n7760 & ~n18203;
  assign n18205 = ~n18202 & n18204;
  assign n18206 = n7984 & n18187;
  assign n18207 = pi626 & ~n18161;
  assign n18208 = ~pi626 & ~n18133;
  assign n18209 = n7759 & ~n18208;
  assign n18210 = ~n18207 & n18209;
  assign n18211 = ~n18206 & ~n18210;
  assign n18212 = ~n18205 & ~n18206;
  assign n18213 = ~n18210 & n18212;
  assign n18214 = ~n18205 & n18211;
  assign n18215 = pi788 & ~n59635;
  assign n18216 = ~n6701 & ~n18175;
  assign n18217 = pi625 & n18216;
  assign n18218 = n18135 & ~n18216;
  assign n18219 = ~n18217 & ~n18218;
  assign n18220 = n18180 & ~n18219;
  assign n18221 = ~pi608 & ~n18179;
  assign n18222 = ~n18220 & n18221;
  assign n18223 = pi1153 & n18135;
  assign n18224 = ~n18217 & n18223;
  assign n18225 = pi608 & ~n18181;
  assign n18226 = ~n18224 & n18225;
  assign n18227 = ~n18222 & ~n18226;
  assign n18228 = pi778 & ~n18227;
  assign n18229 = ~pi778 & ~n18218;
  assign n18230 = ~n18228 & ~n18229;
  assign n18231 = ~pi609 & ~n18230;
  assign n18232 = pi609 & ~n18184;
  assign n18233 = ~pi1155 & ~n18232;
  assign n18234 = ~n18231 & n18233;
  assign n18235 = ~pi660 & ~n18140;
  assign n18236 = ~n18234 & n18235;
  assign n18237 = pi609 & ~n18230;
  assign n18238 = ~pi609 & ~n18184;
  assign n18239 = pi1155 & ~n18238;
  assign n18240 = ~n18237 & n18239;
  assign n18241 = pi660 & ~n18142;
  assign n18242 = ~n18240 & n18241;
  assign n18243 = ~n18236 & ~n18242;
  assign n18244 = pi785 & ~n18243;
  assign n18245 = ~pi785 & ~n18230;
  assign n18246 = ~n18244 & ~n18245;
  assign n18247 = ~pi618 & ~n18246;
  assign n18248 = pi618 & n18185;
  assign n18249 = ~pi1154 & ~n18248;
  assign n18250 = ~n18247 & n18249;
  assign n18251 = ~pi627 & ~n18148;
  assign n18252 = ~n18250 & n18251;
  assign n18253 = pi618 & ~n18246;
  assign n18254 = ~pi618 & n18185;
  assign n18255 = pi1154 & ~n18254;
  assign n18256 = ~n18253 & n18255;
  assign n18257 = pi627 & ~n18150;
  assign n18258 = ~n18256 & n18257;
  assign n18259 = ~n18252 & ~n18258;
  assign n18260 = pi781 & ~n18259;
  assign n18261 = ~pi781 & ~n18246;
  assign n18262 = ~n18260 & ~n18261;
  assign n18263 = pi619 & ~n18262;
  assign n18264 = ~pi619 & n18186;
  assign n18265 = pi1159 & ~n18264;
  assign n18266 = ~n18263 & n18265;
  assign n18267 = pi648 & ~n18158;
  assign n18268 = ~n18266 & n18267;
  assign n18269 = ~pi619 & ~n18262;
  assign n18270 = pi619 & n18186;
  assign n18271 = ~pi1159 & ~n18270;
  assign n18272 = ~n18269 & n18271;
  assign n18273 = ~pi648 & ~n18156;
  assign n18274 = ~n18272 & n18273;
  assign n18275 = pi789 & ~n18274;
  assign n18276 = pi789 & ~n18268;
  assign n18277 = ~n18274 & n18276;
  assign n18278 = ~n18268 & n18275;
  assign n18279 = ~pi789 & n18262;
  assign n18280 = n59242 & ~n18279;
  assign n18281 = ~n59636 & n18280;
  assign n18282 = ~n18215 & ~n18281;
  assign n18283 = ~n59357 & ~n18282;
  assign n18284 = n7957 & ~n59633;
  assign n18285 = n8065 & n18188;
  assign n18286 = pi629 & ~n18285;
  assign n18287 = ~n18284 & n18286;
  assign n18288 = n7958 & ~n59633;
  assign n18289 = n8074 & n18188;
  assign n18290 = ~pi629 & ~n18289;
  assign n18291 = ~n18288 & n18290;
  assign n18292 = pi792 & ~n18291;
  assign n18293 = ~n18288 & ~n18289;
  assign n18294 = ~pi629 & ~n18293;
  assign n18295 = ~n18284 & ~n18285;
  assign n18296 = pi629 & ~n18295;
  assign n18297 = ~n18294 & ~n18296;
  assign n18298 = pi792 & ~n18297;
  assign n18299 = pi792 & ~n18287;
  assign n18300 = ~n18291 & n18299;
  assign n18301 = ~n18287 & n18292;
  assign n18302 = ~n8108 & ~n59637;
  assign n18303 = ~n18283 & n18302;
  assign n18304 = ~n18201 & ~n18303;
  assign n18305 = pi644 & n18304;
  assign n18306 = ~pi787 & ~n18189;
  assign n18307 = pi1157 & ~n18192;
  assign n18308 = ~n18197 & ~n18307;
  assign n18309 = pi787 & ~n18308;
  assign n18310 = ~n18306 & ~n18309;
  assign n18311 = ~pi644 & n18310;
  assign n18312 = pi715 & ~n18311;
  assign n18313 = ~n18305 & n18312;
  assign n18314 = ~n11491 & n18133;
  assign n18315 = ~n7835 & n18168;
  assign n18316 = ~n7835 & ~n18171;
  assign n18317 = n7835 & n18133;
  assign n18318 = ~n18316 & ~n18317;
  assign n18319 = ~n18314 & ~n18315;
  assign n18320 = pi644 & ~n59638;
  assign n18321 = ~pi644 & n18133;
  assign n18322 = ~pi715 & ~n18321;
  assign n18323 = ~n18320 & n18322;
  assign n18324 = pi1160 & ~n18323;
  assign n18325 = ~n18313 & n18324;
  assign n18326 = ~pi644 & n18304;
  assign n18327 = pi644 & n18310;
  assign n18328 = ~pi715 & ~n18327;
  assign n18329 = ~n18326 & n18328;
  assign n18330 = ~pi644 & ~n59638;
  assign n18331 = pi644 & n18133;
  assign n18332 = pi715 & ~n18331;
  assign n18333 = ~n18330 & n18332;
  assign n18334 = ~pi1160 & ~n18333;
  assign n18335 = ~n18329 & n18334;
  assign n18336 = ~n18325 & ~n18335;
  assign n18337 = pi790 & ~n18336;
  assign n18338 = ~pi790 & n18304;
  assign n18339 = pi832 & ~n18338;
  assign n18340 = ~n18337 & n18339;
  assign n18341 = ~pi185 & ~n7560;
  assign n18342 = n59231 & ~n18341;
  assign n18343 = ~pi701 & n59132;
  assign n18344 = n18341 & ~n18343;
  assign n18345 = pi185 & n59251;
  assign n18346 = ~pi38 & ~n18345;
  assign n18347 = n59132 & ~n18346;
  assign n18348 = ~pi185 & n8249;
  assign n18349 = ~n18347 & ~n18348;
  assign n18350 = ~pi185 & ~n6863;
  assign n18351 = n7547 & ~n18350;
  assign n18352 = ~pi701 & ~n18351;
  assign n18353 = ~n18349 & n18352;
  assign n18354 = ~n18344 & ~n18353;
  assign n18355 = ~pi778 & n18354;
  assign n18356 = pi625 & ~n18354;
  assign n18357 = ~pi625 & n18341;
  assign n18358 = pi1153 & ~n18357;
  assign n18359 = ~n18356 & n18358;
  assign n18360 = ~pi625 & ~n18354;
  assign n18361 = pi625 & n18341;
  assign n18362 = ~pi1153 & ~n18361;
  assign n18363 = ~n18360 & n18362;
  assign n18364 = ~n18359 & ~n18363;
  assign n18365 = pi778 & ~n18364;
  assign n18366 = ~n18355 & ~n18365;
  assign n18367 = ~n59229 & n18366;
  assign n18368 = n59229 & n18341;
  assign n18369 = n59229 & ~n18341;
  assign n18370 = ~n59229 & ~n18366;
  assign n18371 = ~n18369 & ~n18370;
  assign n18372 = ~n18367 & ~n18368;
  assign n18373 = ~n59231 & ~n59639;
  assign n18374 = ~n59231 & n59639;
  assign n18375 = n59231 & n18341;
  assign n18376 = ~n18374 & ~n18375;
  assign n18377 = ~n18342 & ~n18373;
  assign n18378 = ~n7716 & ~n59640;
  assign n18379 = n7716 & n18341;
  assign n18380 = n7716 & ~n18341;
  assign n18381 = ~n7716 & n59640;
  assign n18382 = ~n18380 & ~n18381;
  assign n18383 = ~n18378 & ~n18379;
  assign n18384 = ~n7762 & n59641;
  assign n18385 = n7762 & n18341;
  assign n18386 = ~n18384 & ~n18385;
  assign n18387 = ~pi792 & n18386;
  assign n18388 = pi628 & ~n18386;
  assign n18389 = ~pi628 & n18341;
  assign n18390 = pi1156 & ~n18389;
  assign n18391 = ~n18388 & n18390;
  assign n18392 = ~pi628 & ~n18386;
  assign n18393 = pi628 & n18341;
  assign n18394 = ~pi1156 & ~n18393;
  assign n18395 = ~n18392 & n18394;
  assign n18396 = ~n18391 & ~n18395;
  assign n18397 = pi792 & ~n18396;
  assign n18398 = ~n18387 & ~n18397;
  assign n18399 = pi647 & n18398;
  assign n18400 = ~pi647 & n18341;
  assign n18401 = pi647 & ~n18398;
  assign n18402 = ~pi647 & ~n18341;
  assign n18403 = ~n18401 & ~n18402;
  assign n18404 = ~n18399 & ~n18400;
  assign n18405 = pi1157 & ~n59642;
  assign n18406 = ~pi647 & n18398;
  assign n18407 = pi647 & n18341;
  assign n18408 = ~pi1157 & ~n18407;
  assign n18409 = ~n18406 & n18408;
  assign n18410 = ~pi647 & ~n18398;
  assign n18411 = pi647 & ~n18341;
  assign n18412 = ~n18410 & ~n18411;
  assign n18413 = ~pi1157 & n18412;
  assign n18414 = pi1157 & n59642;
  assign n18415 = ~n18413 & ~n18414;
  assign n18416 = ~n18405 & ~n18409;
  assign n18417 = pi787 & n59643;
  assign n18418 = ~pi787 & ~n18398;
  assign n18419 = pi787 & ~n59643;
  assign n18420 = ~pi787 & n18398;
  assign n18421 = ~n18419 & ~n18420;
  assign n18422 = ~n18417 & ~n18418;
  assign n18423 = ~pi644 & ~n59644;
  assign n18424 = pi715 & ~n18423;
  assign n18425 = pi185 & ~n59132;
  assign n18426 = pi751 & n6654;
  assign n18427 = pi185 & n6853;
  assign n18428 = ~n18426 & ~n18427;
  assign n18429 = pi39 & ~n18428;
  assign n18430 = ~pi185 & ~pi751;
  assign n18431 = n59164 & n18430;
  assign n18432 = pi185 & pi751;
  assign n18433 = pi751 & n59147;
  assign n18434 = pi185 & ~n6798;
  assign n18435 = ~n18433 & ~n18434;
  assign n18436 = ~pi39 & ~n18435;
  assign n18437 = ~n18432 & ~n18436;
  assign n18438 = ~n18431 & n18437;
  assign n18439 = ~n18429 & n18438;
  assign n18440 = ~pi38 & ~n18439;
  assign n18441 = ~pi751 & n6865;
  assign n18442 = pi38 & ~n18350;
  assign n18443 = ~n18441 & n18442;
  assign n18444 = ~n18440 & ~n18443;
  assign n18445 = n59132 & ~n18444;
  assign n18446 = ~n18425 & ~n18445;
  assign n18447 = ~n7597 & ~n18446;
  assign n18448 = n7597 & ~n18341;
  assign n18449 = ~n18447 & ~n18448;
  assign n18450 = ~pi785 & ~n18449;
  assign n18451 = ~n7598 & ~n18341;
  assign n18452 = pi609 & n18447;
  assign n18453 = ~n18451 & ~n18452;
  assign n18454 = pi1155 & ~n18453;
  assign n18455 = ~n7610 & ~n18341;
  assign n18456 = ~pi609 & n18447;
  assign n18457 = ~n18455 & ~n18456;
  assign n18458 = ~pi1155 & ~n18457;
  assign n18459 = ~n18454 & ~n18458;
  assign n18460 = pi785 & ~n18459;
  assign n18461 = ~n18450 & ~n18460;
  assign n18462 = ~pi781 & ~n18461;
  assign n18463 = pi618 & n18461;
  assign n18464 = ~pi618 & n18341;
  assign n18465 = pi1154 & ~n18464;
  assign n18466 = ~n18463 & n18465;
  assign n18467 = ~pi618 & n18461;
  assign n18468 = pi618 & n18341;
  assign n18469 = ~pi1154 & ~n18468;
  assign n18470 = ~n18467 & n18469;
  assign n18471 = ~n18466 & ~n18470;
  assign n18472 = pi781 & ~n18471;
  assign n18473 = ~n18462 & ~n18472;
  assign n18474 = ~pi789 & ~n18473;
  assign n18475 = pi619 & n18473;
  assign n18476 = ~pi619 & n18341;
  assign n18477 = pi1159 & ~n18476;
  assign n18478 = ~n18475 & n18477;
  assign n18479 = ~pi619 & n18473;
  assign n18480 = pi619 & n18341;
  assign n18481 = ~pi1159 & ~n18480;
  assign n18482 = ~n18479 & n18481;
  assign n18483 = ~n18478 & ~n18482;
  assign n18484 = pi789 & ~n18483;
  assign n18485 = ~n18474 & ~n18484;
  assign n18486 = ~n8054 & n18485;
  assign n18487 = n8054 & n18341;
  assign n18488 = ~n18486 & ~n18487;
  assign n18489 = ~n7793 & ~n18488;
  assign n18490 = n7793 & n18341;
  assign n18491 = ~n18489 & ~n18490;
  assign n18492 = ~n7835 & ~n18491;
  assign n18493 = n7835 & n18341;
  assign n18494 = n7835 & ~n18341;
  assign n18495 = ~n7835 & n18491;
  assign n18496 = ~n18494 & ~n18495;
  assign n18497 = ~n18492 & ~n18493;
  assign n18498 = pi644 & n59645;
  assign n18499 = ~pi644 & n18341;
  assign n18500 = ~pi715 & ~n18499;
  assign n18501 = ~n18498 & n18500;
  assign n18502 = pi1160 & ~n18501;
  assign n18503 = ~n18424 & n18502;
  assign n18504 = pi644 & ~n59644;
  assign n18505 = ~pi715 & ~n18504;
  assign n18506 = ~pi644 & n59645;
  assign n18507 = pi644 & n18341;
  assign n18508 = pi715 & ~n18507;
  assign n18509 = ~n18506 & n18508;
  assign n18510 = ~pi1160 & ~n18509;
  assign n18511 = ~n18505 & n18510;
  assign n18512 = ~n18503 & ~n18511;
  assign n18513 = pi790 & ~n18512;
  assign n18514 = ~pi644 & n18510;
  assign n18515 = pi644 & n18502;
  assign n18516 = pi790 & ~n18515;
  assign n18517 = pi790 & ~n18514;
  assign n18518 = ~n18515 & n18517;
  assign n18519 = ~n18514 & n18516;
  assign n18520 = ~n7872 & n18491;
  assign n18521 = n7832 & ~n59642;
  assign n18522 = n7833 & ~n18412;
  assign n18523 = pi630 & n18409;
  assign n18524 = ~n18521 & ~n59647;
  assign n18525 = ~n18520 & n18524;
  assign n18526 = pi787 & ~n18525;
  assign n18527 = ~n11154 & n18488;
  assign n18528 = ~pi629 & n18391;
  assign n18529 = pi629 & n18395;
  assign n18530 = ~n18528 & ~n18529;
  assign n18531 = ~n18527 & n18530;
  assign n18532 = pi792 & ~n18531;
  assign n18533 = pi701 & n18444;
  assign n18534 = ~pi185 & n59177;
  assign n18535 = pi185 & n7111;
  assign n18536 = pi751 & ~n18535;
  assign n18537 = ~n18534 & n18536;
  assign n18538 = pi185 & n7188;
  assign n18539 = ~pi185 & ~n59203;
  assign n18540 = ~pi751 & ~n18539;
  assign n18541 = ~n18538 & n18540;
  assign n18542 = pi39 & ~n18541;
  assign n18543 = ~n18537 & n18542;
  assign n18544 = pi185 & n7333;
  assign n18545 = ~pi185 & n7310;
  assign n18546 = pi751 & ~n18545;
  assign n18547 = ~n18544 & n18546;
  assign n18548 = ~pi185 & ~n7339;
  assign n18549 = pi185 & ~n7347;
  assign n18550 = ~pi751 & ~n18549;
  assign n18551 = ~n18548 & n18550;
  assign n18552 = ~pi39 & ~n18551;
  assign n18553 = pi185 & ~n7333;
  assign n18554 = ~pi185 & ~n7310;
  assign n18555 = pi751 & ~n18554;
  assign n18556 = pi751 & ~n18553;
  assign n18557 = ~n18554 & n18556;
  assign n18558 = ~n18553 & n18555;
  assign n18559 = ~pi185 & n7339;
  assign n18560 = pi185 & n7347;
  assign n18561 = ~pi751 & ~n18560;
  assign n18562 = ~n18559 & n18561;
  assign n18563 = ~n59648 & ~n18562;
  assign n18564 = ~pi39 & ~n18563;
  assign n18565 = ~n18547 & n18552;
  assign n18566 = ~pi38 & ~n59649;
  assign n18567 = ~n18543 & n18566;
  assign n18568 = ~pi751 & ~n7222;
  assign n18569 = n9794 & ~n18568;
  assign n18570 = ~pi185 & ~n18569;
  assign n18571 = ~n7056 & ~n18134;
  assign n18572 = pi185 & ~n18571;
  assign n18573 = n59171 & n18572;
  assign n18574 = pi38 & ~n18573;
  assign n18575 = ~n18570 & n18574;
  assign n18576 = ~pi701 & ~n18575;
  assign n18577 = ~n18567 & n18576;
  assign n18578 = n59132 & ~n18577;
  assign n18579 = ~n18533 & n18578;
  assign n18580 = ~n18425 & ~n18579;
  assign n18581 = ~pi625 & n18580;
  assign n18582 = pi625 & n18446;
  assign n18583 = ~pi1153 & ~n18582;
  assign n18584 = ~n18581 & n18583;
  assign n18585 = ~pi608 & ~n18359;
  assign n18586 = ~n18584 & n18585;
  assign n18587 = pi625 & n18580;
  assign n18588 = ~pi625 & n18446;
  assign n18589 = pi1153 & ~n18588;
  assign n18590 = ~n18587 & n18589;
  assign n18591 = pi608 & ~n18363;
  assign n18592 = ~n18590 & n18591;
  assign n18593 = ~n18586 & ~n18592;
  assign n18594 = pi778 & ~n18593;
  assign n18595 = ~pi778 & n18580;
  assign n18596 = ~n18594 & ~n18595;
  assign n18597 = ~pi609 & ~n18596;
  assign n18598 = pi609 & n18366;
  assign n18599 = ~pi1155 & ~n18598;
  assign n18600 = ~n18597 & n18599;
  assign n18601 = ~pi660 & ~n18454;
  assign n18602 = ~n18600 & n18601;
  assign n18603 = pi609 & ~n18596;
  assign n18604 = ~pi609 & n18366;
  assign n18605 = pi1155 & ~n18604;
  assign n18606 = ~n18603 & n18605;
  assign n18607 = pi660 & ~n18458;
  assign n18608 = ~n18606 & n18607;
  assign n18609 = ~n18602 & ~n18608;
  assign n18610 = pi785 & ~n18609;
  assign n18611 = ~pi785 & ~n18596;
  assign n18612 = ~n18610 & ~n18611;
  assign n18613 = ~pi618 & ~n18612;
  assign n18614 = pi618 & n59639;
  assign n18615 = ~pi1154 & ~n18614;
  assign n18616 = ~n18613 & n18615;
  assign n18617 = ~pi627 & ~n18466;
  assign n18618 = ~n18616 & n18617;
  assign n18619 = pi618 & ~n18612;
  assign n18620 = ~pi618 & n59639;
  assign n18621 = pi1154 & ~n18620;
  assign n18622 = ~n18619 & n18621;
  assign n18623 = pi627 & ~n18470;
  assign n18624 = ~n18622 & n18623;
  assign n18625 = ~n18618 & ~n18624;
  assign n18626 = pi781 & ~n18625;
  assign n18627 = ~pi781 & ~n18612;
  assign n18628 = ~n18626 & ~n18627;
  assign n18629 = pi619 & ~n18628;
  assign n18630 = ~pi619 & ~n59640;
  assign n18631 = pi1159 & ~n18630;
  assign n18632 = ~n18629 & n18631;
  assign n18633 = pi648 & ~n18482;
  assign n18634 = ~n18632 & n18633;
  assign n18635 = ~pi619 & ~n18628;
  assign n18636 = pi619 & ~n59640;
  assign n18637 = ~pi1159 & ~n18636;
  assign n18638 = ~n18635 & n18637;
  assign n18639 = ~pi648 & ~n18478;
  assign n18640 = ~n18638 & n18639;
  assign n18641 = pi789 & ~n18640;
  assign n18642 = pi789 & ~n18634;
  assign n18643 = ~n18640 & n18642;
  assign n18644 = ~n18634 & n18641;
  assign n18645 = ~pi789 & n18628;
  assign n18646 = n59242 & ~n18645;
  assign n18647 = ~n59650 & n18646;
  assign n18648 = ~pi626 & ~n18485;
  assign n18649 = pi626 & ~n18341;
  assign n18650 = n7760 & ~n18649;
  assign n18651 = ~n18648 & n18650;
  assign n18652 = n7984 & n59641;
  assign n18653 = pi626 & ~n18485;
  assign n18654 = ~pi626 & ~n18341;
  assign n18655 = n7759 & ~n18654;
  assign n18656 = ~n18653 & n18655;
  assign n18657 = ~n18652 & ~n18656;
  assign n18658 = ~n18651 & ~n18652;
  assign n18659 = ~n18656 & n18658;
  assign n18660 = ~n18651 & n18657;
  assign n18661 = pi788 & ~n59651;
  assign n18662 = ~n59357 & ~n18661;
  assign n18663 = ~n18647 & n18662;
  assign n18664 = ~n18532 & ~n18663;
  assign n18665 = ~n8108 & ~n18664;
  assign n18666 = ~n18526 & ~n18665;
  assign n18667 = ~n59646 & n18666;
  assign n18668 = ~n18513 & ~n18667;
  assign n18669 = n58992 & ~n18668;
  assign n18670 = ~pi185 & ~n58992;
  assign n18671 = ~pi832 & ~n18670;
  assign n18672 = ~n18669 & n18671;
  assign po342 = ~n18340 & ~n18672;
  assign n18674 = ~pi186 & ~n2794;
  assign n18675 = ~pi752 & n6822;
  assign n18676 = ~n18674 & ~n18675;
  assign n18677 = ~n7875 & ~n18676;
  assign n18678 = ~pi785 & ~n18677;
  assign n18679 = ~n7880 & ~n18676;
  assign n18680 = pi1155 & ~n18679;
  assign n18681 = ~n7883 & n18677;
  assign n18682 = ~pi1155 & ~n18681;
  assign n18683 = ~n18680 & ~n18682;
  assign n18684 = pi785 & ~n18683;
  assign n18685 = ~n18678 & ~n18684;
  assign n18686 = ~pi781 & ~n18685;
  assign n18687 = ~n7890 & n18685;
  assign n18688 = pi1154 & ~n18687;
  assign n18689 = ~n7893 & n18685;
  assign n18690 = ~pi1154 & ~n18689;
  assign n18691 = ~n18688 & ~n18690;
  assign n18692 = pi781 & ~n18691;
  assign n18693 = ~n18686 & ~n18692;
  assign n18694 = ~pi789 & ~n18693;
  assign n18695 = pi619 & n18693;
  assign n18696 = ~pi619 & n18674;
  assign n18697 = pi1159 & ~n18696;
  assign n18698 = ~n18695 & n18697;
  assign n18699 = ~pi619 & n18693;
  assign n18700 = pi619 & n18674;
  assign n18701 = ~pi1159 & ~n18700;
  assign n18702 = ~n18699 & n18701;
  assign n18703 = ~n18698 & ~n18702;
  assign n18704 = pi789 & ~n18703;
  assign n18705 = ~n18694 & ~n18704;
  assign n18706 = ~n8054 & ~n18705;
  assign n18707 = n8054 & ~n18674;
  assign n18708 = ~n8054 & n18705;
  assign n18709 = n8054 & n18674;
  assign n18710 = ~n18708 & ~n18709;
  assign n18711 = ~n18706 & ~n18707;
  assign n18712 = ~n7793 & ~n59652;
  assign n18713 = n7793 & n18674;
  assign n18714 = ~n7872 & ~n18713;
  assign n18715 = ~n18712 & ~n18713;
  assign n18716 = ~n7872 & n18715;
  assign n18717 = ~n18712 & n18714;
  assign n18718 = pi703 & n7055;
  assign n18719 = ~n18674 & ~n18718;
  assign n18720 = ~pi778 & n18719;
  assign n18721 = ~pi625 & n18718;
  assign n18722 = ~n18719 & ~n18721;
  assign n18723 = pi1153 & ~n18722;
  assign n18724 = ~pi1153 & ~n18674;
  assign n18725 = ~n18721 & n18724;
  assign n18726 = ~n18723 & ~n18725;
  assign n18727 = pi778 & ~n18726;
  assign n18728 = ~n18720 & ~n18727;
  assign n18729 = ~n7949 & n18728;
  assign n18730 = ~n7951 & n18729;
  assign n18731 = ~n7953 & n18730;
  assign n18732 = ~n7955 & n18731;
  assign n18733 = ~n7967 & n18732;
  assign n18734 = pi647 & ~n18733;
  assign n18735 = ~pi647 & ~n18674;
  assign n18736 = ~n18734 & ~n18735;
  assign n18737 = n7832 & ~n18736;
  assign n18738 = ~pi647 & n18733;
  assign n18739 = pi647 & n18674;
  assign n18740 = ~pi1157 & ~n18739;
  assign n18741 = ~n18738 & n18740;
  assign n18742 = pi630 & n18741;
  assign n18743 = ~n18737 & ~n18742;
  assign n18744 = ~n59653 & n18743;
  assign n18745 = pi787 & ~n18744;
  assign n18746 = ~pi626 & ~n18705;
  assign n18747 = pi626 & ~n18674;
  assign n18748 = n7760 & ~n18747;
  assign n18749 = ~n18746 & n18748;
  assign n18750 = n7984 & n18731;
  assign n18751 = pi626 & ~n18705;
  assign n18752 = ~pi626 & ~n18674;
  assign n18753 = n7759 & ~n18752;
  assign n18754 = ~n18751 & n18753;
  assign n18755 = ~n18750 & ~n18754;
  assign n18756 = ~n18749 & ~n18750;
  assign n18757 = ~n18754 & n18756;
  assign n18758 = ~n18749 & n18755;
  assign n18759 = pi788 & ~n59654;
  assign n18760 = ~n6701 & ~n18719;
  assign n18761 = pi625 & n18760;
  assign n18762 = n18676 & ~n18760;
  assign n18763 = ~n18761 & ~n18762;
  assign n18764 = n18724 & ~n18763;
  assign n18765 = ~pi608 & ~n18723;
  assign n18766 = ~n18764 & n18765;
  assign n18767 = pi1153 & n18676;
  assign n18768 = ~n18761 & n18767;
  assign n18769 = pi608 & ~n18725;
  assign n18770 = ~n18768 & n18769;
  assign n18771 = ~n18766 & ~n18770;
  assign n18772 = pi778 & ~n18771;
  assign n18773 = ~pi778 & ~n18762;
  assign n18774 = ~n18772 & ~n18773;
  assign n18775 = ~pi609 & ~n18774;
  assign n18776 = pi609 & n18728;
  assign n18777 = ~pi1155 & ~n18776;
  assign n18778 = ~n18775 & n18777;
  assign n18779 = ~pi660 & ~n18680;
  assign n18780 = ~n18778 & n18779;
  assign n18781 = pi609 & ~n18774;
  assign n18782 = ~pi609 & n18728;
  assign n18783 = pi1155 & ~n18782;
  assign n18784 = ~n18781 & n18783;
  assign n18785 = pi660 & ~n18682;
  assign n18786 = ~n18784 & n18785;
  assign n18787 = ~n18780 & ~n18786;
  assign n18788 = pi785 & ~n18787;
  assign n18789 = ~pi785 & ~n18774;
  assign n18790 = ~n18788 & ~n18789;
  assign n18791 = ~pi618 & ~n18790;
  assign n18792 = pi618 & n18729;
  assign n18793 = ~pi1154 & ~n18792;
  assign n18794 = ~n18791 & n18793;
  assign n18795 = ~pi627 & ~n18688;
  assign n18796 = ~n18794 & n18795;
  assign n18797 = pi618 & ~n18790;
  assign n18798 = ~pi618 & n18729;
  assign n18799 = pi1154 & ~n18798;
  assign n18800 = ~n18797 & n18799;
  assign n18801 = pi627 & ~n18690;
  assign n18802 = ~n18800 & n18801;
  assign n18803 = ~n18796 & ~n18802;
  assign n18804 = pi781 & ~n18803;
  assign n18805 = ~pi781 & ~n18790;
  assign n18806 = ~n18804 & ~n18805;
  assign n18807 = ~pi619 & ~n18806;
  assign n18808 = pi619 & n18730;
  assign n18809 = ~pi1159 & ~n18808;
  assign n18810 = ~n18807 & n18809;
  assign n18811 = ~pi648 & ~n18698;
  assign n18812 = ~n18810 & n18811;
  assign n18813 = pi619 & ~n18806;
  assign n18814 = ~pi619 & n18730;
  assign n18815 = pi1159 & ~n18814;
  assign n18816 = ~n18813 & n18815;
  assign n18817 = pi648 & ~n18702;
  assign n18818 = ~n18816 & n18817;
  assign n18819 = pi789 & ~n18818;
  assign n18820 = pi789 & ~n18812;
  assign n18821 = ~n18818 & n18820;
  assign n18822 = ~n18812 & n18819;
  assign n18823 = ~pi789 & n18806;
  assign n18824 = n59242 & ~n18823;
  assign n18825 = ~n59655 & n18824;
  assign n18826 = ~n18759 & ~n18825;
  assign n18827 = ~n59357 & ~n18826;
  assign n18828 = n7957 & ~n59652;
  assign n18829 = n8065 & n18732;
  assign n18830 = pi629 & ~n18829;
  assign n18831 = ~n18828 & n18830;
  assign n18832 = n7958 & ~n59652;
  assign n18833 = n8074 & n18732;
  assign n18834 = ~pi629 & ~n18833;
  assign n18835 = ~n18832 & n18834;
  assign n18836 = pi792 & ~n18835;
  assign n18837 = ~n18832 & ~n18833;
  assign n18838 = ~pi629 & ~n18837;
  assign n18839 = ~n18828 & ~n18829;
  assign n18840 = pi629 & ~n18839;
  assign n18841 = ~n18838 & ~n18840;
  assign n18842 = pi792 & ~n18841;
  assign n18843 = pi792 & ~n18831;
  assign n18844 = ~n18835 & n18843;
  assign n18845 = ~n18831 & n18836;
  assign n18846 = ~n8108 & ~n59656;
  assign n18847 = ~n18827 & n18846;
  assign n18848 = ~n18745 & ~n18847;
  assign n18849 = pi644 & n18848;
  assign n18850 = ~pi787 & ~n18733;
  assign n18851 = pi1157 & ~n18736;
  assign n18852 = ~n18741 & ~n18851;
  assign n18853 = pi787 & ~n18852;
  assign n18854 = ~n18850 & ~n18853;
  assign n18855 = ~pi644 & n18854;
  assign n18856 = pi715 & ~n18855;
  assign n18857 = ~n18849 & n18856;
  assign n18858 = ~n11491 & n18674;
  assign n18859 = ~n7835 & n18712;
  assign n18860 = ~n7835 & ~n18715;
  assign n18861 = n7835 & n18674;
  assign n18862 = ~n18860 & ~n18861;
  assign n18863 = ~n18858 & ~n18859;
  assign n18864 = pi644 & ~n59657;
  assign n18865 = ~pi644 & n18674;
  assign n18866 = ~pi715 & ~n18865;
  assign n18867 = ~n18864 & n18866;
  assign n18868 = pi1160 & ~n18867;
  assign n18869 = ~n18857 & n18868;
  assign n18870 = ~pi644 & n18848;
  assign n18871 = pi644 & n18854;
  assign n18872 = ~pi715 & ~n18871;
  assign n18873 = ~n18870 & n18872;
  assign n18874 = ~pi644 & ~n59657;
  assign n18875 = pi644 & n18674;
  assign n18876 = pi715 & ~n18875;
  assign n18877 = ~n18874 & n18876;
  assign n18878 = ~pi1160 & ~n18877;
  assign n18879 = ~n18873 & n18878;
  assign n18880 = ~n18869 & ~n18879;
  assign n18881 = pi790 & ~n18880;
  assign n18882 = ~pi790 & n18848;
  assign n18883 = pi832 & ~n18882;
  assign n18884 = ~n18881 & n18883;
  assign n18885 = pi186 & ~n59132;
  assign n18886 = ~pi186 & ~n7553;
  assign n18887 = pi752 & ~n18886;
  assign n18888 = pi186 & ~n9781;
  assign n18889 = ~pi186 & ~pi752;
  assign n18890 = n9787 & n18889;
  assign n18891 = ~n18888 & ~n18890;
  assign n18892 = ~n9780 & ~n18891;
  assign n18893 = ~n18887 & ~n18892;
  assign n18894 = n59132 & ~n18893;
  assign n18895 = ~n18885 & ~n18894;
  assign n18896 = ~n7597 & ~n18895;
  assign n18897 = ~pi186 & ~n7560;
  assign n18898 = n7597 & ~n18897;
  assign n18899 = ~n18896 & ~n18898;
  assign n18900 = ~pi785 & ~n18899;
  assign n18901 = ~n7598 & ~n18897;
  assign n18902 = pi609 & n18896;
  assign n18903 = ~n18901 & ~n18902;
  assign n18904 = pi1155 & ~n18903;
  assign n18905 = ~n7610 & ~n18897;
  assign n18906 = ~pi609 & n18896;
  assign n18907 = ~n18905 & ~n18906;
  assign n18908 = ~pi1155 & ~n18907;
  assign n18909 = ~n18904 & ~n18908;
  assign n18910 = pi785 & ~n18909;
  assign n18911 = ~n18900 & ~n18910;
  assign n18912 = ~pi781 & ~n18911;
  assign n18913 = pi618 & n18911;
  assign n18914 = ~pi618 & n18897;
  assign n18915 = pi1154 & ~n18914;
  assign n18916 = ~n18913 & n18915;
  assign n18917 = ~pi618 & n18911;
  assign n18918 = pi618 & n18897;
  assign n18919 = ~pi1154 & ~n18918;
  assign n18920 = ~n18917 & n18919;
  assign n18921 = ~n18916 & ~n18920;
  assign n18922 = pi781 & ~n18921;
  assign n18923 = ~n18912 & ~n18922;
  assign n18924 = ~pi789 & ~n18923;
  assign n18925 = ~pi619 & n18923;
  assign n18926 = pi619 & n18897;
  assign n18927 = ~pi1159 & ~n18926;
  assign n18928 = ~n18925 & n18927;
  assign n18929 = pi619 & n18923;
  assign n18930 = ~pi619 & n18897;
  assign n18931 = pi1159 & ~n18930;
  assign n18932 = ~n18929 & n18931;
  assign n18933 = ~n18928 & ~n18932;
  assign n18934 = pi789 & ~n18933;
  assign n18935 = ~n18924 & ~n18934;
  assign n18936 = ~n8054 & n18935;
  assign n18937 = n8054 & n18897;
  assign n18938 = ~n18936 & ~n18937;
  assign n18939 = ~n11154 & n18938;
  assign n18940 = n7762 & ~n18897;
  assign n18941 = n59231 & ~n18897;
  assign n18942 = ~pi186 & n8249;
  assign n18943 = pi186 & n59251;
  assign n18944 = ~pi38 & ~n18943;
  assign n18945 = ~n18942 & n18944;
  assign n18946 = ~pi186 & ~n6863;
  assign n18947 = n7547 & ~n18946;
  assign n18948 = pi703 & ~n18947;
  assign n18949 = ~n18945 & n18948;
  assign n18950 = ~pi703 & n18886;
  assign n18951 = n59132 & ~n18950;
  assign n18952 = ~n18949 & n18951;
  assign n18953 = ~n18885 & ~n18952;
  assign n18954 = ~pi778 & ~n18953;
  assign n18955 = ~pi625 & n18953;
  assign n18956 = pi625 & n18897;
  assign n18957 = ~pi1153 & ~n18956;
  assign n18958 = ~n18955 & n18957;
  assign n18959 = pi625 & n18953;
  assign n18960 = ~pi625 & n18897;
  assign n18961 = pi1153 & ~n18960;
  assign n18962 = ~n18959 & n18961;
  assign n18963 = ~n18958 & ~n18962;
  assign n18964 = pi778 & ~n18963;
  assign n18965 = ~n18954 & ~n18964;
  assign n18966 = ~n59229 & n18965;
  assign n18967 = n59229 & n18897;
  assign n18968 = n59229 & ~n18897;
  assign n18969 = ~n59229 & ~n18965;
  assign n18970 = ~n18968 & ~n18969;
  assign n18971 = ~n18966 & ~n18967;
  assign n18972 = ~n59231 & ~n59658;
  assign n18973 = ~n59231 & n59658;
  assign n18974 = n59231 & n18897;
  assign n18975 = ~n18973 & ~n18974;
  assign n18976 = ~n18941 & ~n18972;
  assign n18977 = ~n7716 & ~n59659;
  assign n18978 = n7716 & n18897;
  assign n18979 = n7716 & ~n18897;
  assign n18980 = ~n7716 & n59659;
  assign n18981 = ~n18979 & ~n18980;
  assign n18982 = ~n18977 & ~n18978;
  assign n18983 = ~n7762 & ~n59660;
  assign n18984 = ~n7762 & n59660;
  assign n18985 = n7762 & n18897;
  assign n18986 = ~n18984 & ~n18985;
  assign n18987 = ~n18940 & ~n18983;
  assign n18988 = ~pi628 & ~n59661;
  assign n18989 = pi628 & n18897;
  assign n18990 = ~pi1156 & ~n18989;
  assign n18991 = ~n18988 & n18990;
  assign n18992 = pi629 & n18991;
  assign n18993 = ~pi628 & ~n18897;
  assign n18994 = pi628 & n59661;
  assign n18995 = ~n18993 & ~n18994;
  assign n18996 = n7790 & ~n18995;
  assign n18997 = ~n18992 & ~n18996;
  assign n18998 = ~n18939 & n18997;
  assign n18999 = pi792 & ~n18998;
  assign n19000 = pi619 & ~n59659;
  assign n19001 = ~pi1159 & ~n19000;
  assign n19002 = ~pi648 & ~n18932;
  assign n19003 = ~n19001 & n19002;
  assign n19004 = ~pi619 & ~n59659;
  assign n19005 = pi1159 & ~n19004;
  assign n19006 = pi648 & ~n18928;
  assign n19007 = ~n19005 & n19006;
  assign n19008 = ~n19003 & ~n19007;
  assign n19009 = pi789 & ~n19008;
  assign n19010 = pi618 & n59658;
  assign n19011 = ~pi1154 & ~n19010;
  assign n19012 = ~pi627 & ~n18916;
  assign n19013 = ~n19011 & n19012;
  assign n19014 = ~pi703 & n18893;
  assign n19015 = ~pi186 & n9797;
  assign n19016 = pi186 & n9799;
  assign n19017 = pi752 & ~n9801;
  assign n19018 = ~n19016 & n19017;
  assign n19019 = ~n19015 & n19018;
  assign n19020 = pi186 & n9811;
  assign n19021 = ~pi186 & ~n59320;
  assign n19022 = ~pi752 & ~n19021;
  assign n19023 = ~n19020 & n19022;
  assign n19024 = pi703 & ~n19023;
  assign n19025 = ~n19019 & n19024;
  assign n19026 = n59132 & ~n19025;
  assign n19027 = n59132 & ~n19014;
  assign n19028 = ~n19025 & n19027;
  assign n19029 = ~n19014 & n19026;
  assign n19030 = ~n18885 & ~n59662;
  assign n19031 = pi625 & n19030;
  assign n19032 = ~pi625 & n18895;
  assign n19033 = pi1153 & ~n19032;
  assign n19034 = ~n19031 & n19033;
  assign n19035 = pi608 & ~n18958;
  assign n19036 = ~n19034 & n19035;
  assign n19037 = ~pi625 & n19030;
  assign n19038 = pi625 & n18895;
  assign n19039 = ~pi1153 & ~n19038;
  assign n19040 = ~n19037 & n19039;
  assign n19041 = ~pi608 & ~n18962;
  assign n19042 = ~n19040 & n19041;
  assign n19043 = ~n19036 & ~n19042;
  assign n19044 = pi778 & ~n19043;
  assign n19045 = ~pi778 & n19030;
  assign n19046 = ~pi778 & ~n19030;
  assign n19047 = pi778 & ~n19042;
  assign n19048 = ~n19036 & n19047;
  assign n19049 = ~n19046 & ~n19048;
  assign n19050 = ~n19044 & ~n19045;
  assign n19051 = ~pi609 & n59663;
  assign n19052 = pi609 & n18965;
  assign n19053 = ~pi1155 & ~n19052;
  assign n19054 = ~n19051 & n19053;
  assign n19055 = ~pi660 & ~n18904;
  assign n19056 = ~n19054 & n19055;
  assign n19057 = pi609 & n59663;
  assign n19058 = ~pi609 & n18965;
  assign n19059 = pi1155 & ~n19058;
  assign n19060 = ~n19057 & n19059;
  assign n19061 = pi660 & ~n18908;
  assign n19062 = ~n19060 & n19061;
  assign n19063 = ~n19056 & ~n19062;
  assign n19064 = pi785 & ~n19063;
  assign n19065 = ~pi785 & n59663;
  assign n19066 = ~n19064 & ~n19065;
  assign n19067 = pi618 & ~n19066;
  assign n19068 = ~pi618 & n59658;
  assign n19069 = pi1154 & ~n19068;
  assign n19070 = ~n19067 & n19069;
  assign n19071 = pi627 & ~n18920;
  assign n19072 = ~n19070 & n19071;
  assign n19073 = ~n19013 & ~n19072;
  assign n19074 = pi781 & ~n19073;
  assign n19075 = ~pi618 & n19012;
  assign n19076 = pi781 & ~n19075;
  assign n19077 = ~n19066 & ~n19076;
  assign n19078 = ~pi618 & ~n19066;
  assign n19079 = n19011 & ~n19078;
  assign n19080 = n19012 & ~n19079;
  assign n19081 = ~n19072 & ~n19080;
  assign n19082 = pi781 & ~n19081;
  assign n19083 = ~pi781 & ~n19066;
  assign n19084 = ~n19082 & ~n19083;
  assign n19085 = ~n19074 & ~n19077;
  assign n19086 = ~pi619 & n19002;
  assign n19087 = pi619 & n19006;
  assign n19088 = pi789 & ~n19087;
  assign n19089 = ~n19086 & n19088;
  assign n19090 = ~n59664 & ~n19089;
  assign n19091 = ~pi619 & ~n59664;
  assign n19092 = n19001 & ~n19091;
  assign n19093 = n19002 & ~n19092;
  assign n19094 = pi619 & ~n59664;
  assign n19095 = n19005 & ~n19094;
  assign n19096 = n19006 & ~n19095;
  assign n19097 = ~n19093 & ~n19096;
  assign n19098 = pi789 & ~n19097;
  assign n19099 = ~pi789 & ~n59664;
  assign n19100 = ~n19098 & ~n19099;
  assign n19101 = ~n19009 & ~n19090;
  assign n19102 = n59242 & ~n59665;
  assign n19103 = n12139 & n18935;
  assign n19104 = ~pi641 & ~n59660;
  assign n19105 = pi641 & ~n18897;
  assign n19106 = n7912 & ~n19105;
  assign n19107 = ~n19104 & n19106;
  assign n19108 = pi641 & ~n59660;
  assign n19109 = ~pi641 & ~n18897;
  assign n19110 = n7911 & ~n19109;
  assign n19111 = ~n19108 & n19110;
  assign n19112 = ~n19107 & ~n19111;
  assign n19113 = ~n19103 & n19112;
  assign n19114 = pi788 & ~n19113;
  assign n19115 = ~n59357 & ~n19114;
  assign n19116 = ~n19102 & n19115;
  assign n19117 = ~pi788 & n59665;
  assign n19118 = ~pi626 & n59665;
  assign n19119 = pi626 & ~n59660;
  assign n19120 = ~pi641 & ~n19119;
  assign n19121 = ~n19118 & n19120;
  assign n19122 = ~pi626 & ~n18935;
  assign n19123 = pi626 & ~n18897;
  assign n19124 = pi641 & ~n19123;
  assign n19125 = ~n19122 & n19124;
  assign n19126 = ~pi1158 & ~n19125;
  assign n19127 = ~n19121 & n19126;
  assign n19128 = pi626 & n59665;
  assign n19129 = ~pi626 & ~n59660;
  assign n19130 = pi641 & ~n19129;
  assign n19131 = ~n19128 & n19130;
  assign n19132 = pi626 & ~n18935;
  assign n19133 = ~pi626 & ~n18897;
  assign n19134 = ~pi641 & ~n19133;
  assign n19135 = ~n19132 & n19134;
  assign n19136 = pi1158 & ~n19135;
  assign n19137 = ~n19131 & n19136;
  assign n19138 = ~n19127 & ~n19137;
  assign n19139 = pi788 & ~n19138;
  assign n19140 = ~n19117 & ~n19139;
  assign n19141 = ~pi628 & n19140;
  assign n19142 = pi628 & ~n18938;
  assign n19143 = ~pi1156 & ~n19142;
  assign n19144 = ~n19141 & n19143;
  assign n19145 = pi628 & ~n59661;
  assign n19146 = ~pi628 & n18897;
  assign n19147 = pi1156 & ~n19146;
  assign n19148 = pi1156 & ~n18995;
  assign n19149 = ~n19145 & n19147;
  assign n19150 = ~pi629 & ~n59666;
  assign n19151 = ~n19144 & n19150;
  assign n19152 = pi628 & n19140;
  assign n19153 = ~pi628 & ~n18938;
  assign n19154 = pi1156 & ~n19153;
  assign n19155 = ~n19152 & n19154;
  assign n19156 = pi629 & ~n18991;
  assign n19157 = ~n19155 & n19156;
  assign n19158 = ~n19151 & ~n19157;
  assign n19159 = pi792 & ~n19158;
  assign n19160 = ~pi792 & n19140;
  assign n19161 = ~n19159 & ~n19160;
  assign n19162 = ~n18999 & ~n19116;
  assign n19163 = n59244 & n59667;
  assign n19164 = ~pi647 & ~n18897;
  assign n19165 = ~pi792 & n59661;
  assign n19166 = ~n18991 & ~n59666;
  assign n19167 = pi792 & ~n19166;
  assign n19168 = ~n19165 & ~n19167;
  assign n19169 = pi647 & ~n19168;
  assign n19170 = ~n19164 & ~n19169;
  assign n19171 = n7832 & ~n19170;
  assign n19172 = ~pi647 & n19168;
  assign n19173 = pi647 & n18897;
  assign n19174 = ~pi1157 & ~n19173;
  assign n19175 = ~n19172 & n19174;
  assign n19176 = pi630 & n19175;
  assign n19177 = ~n7793 & ~n18938;
  assign n19178 = n7793 & n18897;
  assign n19179 = ~n19177 & ~n19178;
  assign n19180 = ~n7872 & n19179;
  assign n19181 = ~n19176 & ~n19180;
  assign n19182 = ~n19171 & n19181;
  assign n19183 = ~pi647 & ~n59667;
  assign n19184 = pi647 & ~n19179;
  assign n19185 = ~pi1157 & ~n19184;
  assign n19186 = ~n19183 & n19185;
  assign n19187 = pi647 & n19168;
  assign n19188 = ~pi647 & n18897;
  assign n19189 = pi1157 & ~n19188;
  assign n19190 = pi1157 & ~n19170;
  assign n19191 = ~n19187 & n19189;
  assign n19192 = ~pi630 & ~n59668;
  assign n19193 = ~n19186 & n19192;
  assign n19194 = pi647 & ~n59667;
  assign n19195 = ~pi647 & ~n19179;
  assign n19196 = pi1157 & ~n19195;
  assign n19197 = ~n19194 & n19196;
  assign n19198 = pi630 & ~n19175;
  assign n19199 = ~n19197 & n19198;
  assign n19200 = ~n19193 & ~n19199;
  assign n19201 = ~n19163 & n19182;
  assign n19202 = pi787 & n59669;
  assign n19203 = ~pi787 & n59667;
  assign n19204 = pi787 & ~n59669;
  assign n19205 = ~pi787 & ~n59667;
  assign n19206 = ~n19204 & ~n19205;
  assign n19207 = ~n19202 & ~n19203;
  assign n19208 = pi644 & ~n59670;
  assign n19209 = ~pi787 & ~n19168;
  assign n19210 = ~n19175 & ~n59668;
  assign n19211 = pi787 & ~n19210;
  assign n19212 = ~n19209 & ~n19211;
  assign n19213 = ~pi644 & n19212;
  assign n19214 = pi715 & ~n19213;
  assign n19215 = ~n19208 & n19214;
  assign n19216 = ~n7835 & ~n19179;
  assign n19217 = n7835 & n18897;
  assign n19218 = n7835 & ~n18897;
  assign n19219 = ~n7835 & n19179;
  assign n19220 = ~n19218 & ~n19219;
  assign n19221 = ~n19216 & ~n19217;
  assign n19222 = pi644 & n59671;
  assign n19223 = ~pi644 & n18897;
  assign n19224 = ~pi715 & ~n19223;
  assign n19225 = ~n19222 & n19224;
  assign n19226 = pi1160 & ~n19225;
  assign n19227 = ~n19215 & n19226;
  assign n19228 = ~pi644 & n59671;
  assign n19229 = pi644 & n18897;
  assign n19230 = pi715 & ~n19229;
  assign n19231 = ~n19228 & n19230;
  assign n19232 = ~pi1160 & ~n19231;
  assign n19233 = pi644 & n19212;
  assign n19234 = ~pi715 & ~n19233;
  assign n19235 = ~pi644 & ~n59670;
  assign n19236 = n19234 & ~n19235;
  assign n19237 = n19232 & ~n19236;
  assign n19238 = pi790 & ~n19237;
  assign n19239 = pi790 & ~n19227;
  assign n19240 = ~n19237 & n19239;
  assign n19241 = ~n19227 & n19238;
  assign n19242 = ~pi790 & n59670;
  assign n19243 = n58992 & ~n19242;
  assign n19244 = n19232 & ~n19234;
  assign n19245 = ~n19227 & ~n19244;
  assign n19246 = pi790 & ~n19245;
  assign n19247 = ~pi644 & n19232;
  assign n19248 = pi790 & ~n19247;
  assign n19249 = ~n59670 & ~n19248;
  assign n19250 = ~n19246 & ~n19249;
  assign n19251 = n58992 & ~n19250;
  assign n19252 = ~n59672 & n19243;
  assign n19253 = ~pi186 & ~n58992;
  assign n19254 = ~pi832 & ~n19253;
  assign n19255 = ~n59673 & n19254;
  assign po343 = ~n18884 & ~n19255;
  assign n19257 = ~pi187 & ~n2794;
  assign n19258 = ~pi770 & n6822;
  assign n19259 = ~n19257 & ~n19258;
  assign n19260 = ~n7875 & ~n19259;
  assign n19261 = ~pi785 & ~n19260;
  assign n19262 = ~n7880 & ~n19259;
  assign n19263 = pi1155 & ~n19262;
  assign n19264 = ~n7883 & n19260;
  assign n19265 = ~pi1155 & ~n19264;
  assign n19266 = ~n19263 & ~n19265;
  assign n19267 = pi785 & ~n19266;
  assign n19268 = ~n19261 & ~n19267;
  assign n19269 = ~pi781 & ~n19268;
  assign n19270 = ~n7890 & n19268;
  assign n19271 = pi1154 & ~n19270;
  assign n19272 = ~n7893 & n19268;
  assign n19273 = ~pi1154 & ~n19272;
  assign n19274 = ~n19271 & ~n19273;
  assign n19275 = pi781 & ~n19274;
  assign n19276 = ~n19269 & ~n19275;
  assign n19277 = ~pi789 & ~n19276;
  assign n19278 = pi619 & n19276;
  assign n19279 = ~pi619 & n19257;
  assign n19280 = pi1159 & ~n19279;
  assign n19281 = ~n19278 & n19280;
  assign n19282 = ~pi619 & n19276;
  assign n19283 = pi619 & n19257;
  assign n19284 = ~pi1159 & ~n19283;
  assign n19285 = ~n19282 & n19284;
  assign n19286 = ~n19281 & ~n19285;
  assign n19287 = pi789 & ~n19286;
  assign n19288 = ~n19277 & ~n19287;
  assign n19289 = ~n8054 & ~n19288;
  assign n19290 = n8054 & ~n19257;
  assign n19291 = ~n8054 & n19288;
  assign n19292 = n8054 & n19257;
  assign n19293 = ~n19291 & ~n19292;
  assign n19294 = ~n19289 & ~n19290;
  assign n19295 = ~n7793 & ~n59674;
  assign n19296 = n7793 & n19257;
  assign n19297 = ~n7872 & ~n19296;
  assign n19298 = ~n19295 & ~n19296;
  assign n19299 = ~n7872 & n19298;
  assign n19300 = ~n19295 & n19297;
  assign n19301 = pi726 & n7055;
  assign n19302 = ~n19257 & ~n19301;
  assign n19303 = ~pi778 & n19302;
  assign n19304 = ~pi625 & n19301;
  assign n19305 = ~n19302 & ~n19304;
  assign n19306 = pi1153 & ~n19305;
  assign n19307 = ~pi1153 & ~n19257;
  assign n19308 = ~n19304 & n19307;
  assign n19309 = ~n19306 & ~n19308;
  assign n19310 = pi778 & ~n19309;
  assign n19311 = ~n19303 & ~n19310;
  assign n19312 = ~n7949 & n19311;
  assign n19313 = ~n7951 & n19312;
  assign n19314 = ~n7953 & n19313;
  assign n19315 = ~n7955 & n19314;
  assign n19316 = ~n7967 & n19315;
  assign n19317 = pi647 & ~n19316;
  assign n19318 = ~pi647 & ~n19257;
  assign n19319 = ~n19317 & ~n19318;
  assign n19320 = n7832 & ~n19319;
  assign n19321 = ~pi647 & n19316;
  assign n19322 = pi647 & n19257;
  assign n19323 = ~pi1157 & ~n19322;
  assign n19324 = ~n19321 & n19323;
  assign n19325 = pi630 & n19324;
  assign n19326 = ~n19320 & ~n19325;
  assign n19327 = ~n59675 & n19326;
  assign n19328 = pi787 & ~n19327;
  assign n19329 = ~pi626 & ~n19288;
  assign n19330 = pi626 & ~n19257;
  assign n19331 = n7760 & ~n19330;
  assign n19332 = ~n19329 & n19331;
  assign n19333 = n7984 & n19314;
  assign n19334 = pi626 & ~n19288;
  assign n19335 = ~pi626 & ~n19257;
  assign n19336 = n7759 & ~n19335;
  assign n19337 = ~n19334 & n19336;
  assign n19338 = ~n19333 & ~n19337;
  assign n19339 = ~n19332 & ~n19333;
  assign n19340 = ~n19337 & n19339;
  assign n19341 = ~n19332 & n19338;
  assign n19342 = pi788 & ~n59676;
  assign n19343 = ~n6701 & ~n19302;
  assign n19344 = pi625 & n19343;
  assign n19345 = n19259 & ~n19343;
  assign n19346 = ~n19344 & ~n19345;
  assign n19347 = n19307 & ~n19346;
  assign n19348 = ~pi608 & ~n19306;
  assign n19349 = ~n19347 & n19348;
  assign n19350 = pi1153 & n19259;
  assign n19351 = ~n19344 & n19350;
  assign n19352 = pi608 & ~n19308;
  assign n19353 = ~n19351 & n19352;
  assign n19354 = ~n19349 & ~n19353;
  assign n19355 = pi778 & ~n19354;
  assign n19356 = ~pi778 & ~n19345;
  assign n19357 = ~n19355 & ~n19356;
  assign n19358 = ~pi609 & ~n19357;
  assign n19359 = pi609 & n19311;
  assign n19360 = ~pi1155 & ~n19359;
  assign n19361 = ~n19358 & n19360;
  assign n19362 = ~pi660 & ~n19263;
  assign n19363 = ~n19361 & n19362;
  assign n19364 = pi609 & ~n19357;
  assign n19365 = ~pi609 & n19311;
  assign n19366 = pi1155 & ~n19365;
  assign n19367 = ~n19364 & n19366;
  assign n19368 = pi660 & ~n19265;
  assign n19369 = ~n19367 & n19368;
  assign n19370 = ~n19363 & ~n19369;
  assign n19371 = pi785 & ~n19370;
  assign n19372 = ~pi785 & ~n19357;
  assign n19373 = ~n19371 & ~n19372;
  assign n19374 = ~pi618 & ~n19373;
  assign n19375 = pi618 & n19312;
  assign n19376 = ~pi1154 & ~n19375;
  assign n19377 = ~n19374 & n19376;
  assign n19378 = ~pi627 & ~n19271;
  assign n19379 = ~n19377 & n19378;
  assign n19380 = pi618 & ~n19373;
  assign n19381 = ~pi618 & n19312;
  assign n19382 = pi1154 & ~n19381;
  assign n19383 = ~n19380 & n19382;
  assign n19384 = pi627 & ~n19273;
  assign n19385 = ~n19383 & n19384;
  assign n19386 = ~n19379 & ~n19385;
  assign n19387 = pi781 & ~n19386;
  assign n19388 = ~pi781 & ~n19373;
  assign n19389 = ~n19387 & ~n19388;
  assign n19390 = ~pi619 & ~n19389;
  assign n19391 = pi619 & n19313;
  assign n19392 = ~pi1159 & ~n19391;
  assign n19393 = ~n19390 & n19392;
  assign n19394 = ~pi648 & ~n19281;
  assign n19395 = ~n19393 & n19394;
  assign n19396 = pi619 & ~n19389;
  assign n19397 = ~pi619 & n19313;
  assign n19398 = pi1159 & ~n19397;
  assign n19399 = ~n19396 & n19398;
  assign n19400 = pi648 & ~n19285;
  assign n19401 = ~n19399 & n19400;
  assign n19402 = pi789 & ~n19401;
  assign n19403 = pi789 & ~n19395;
  assign n19404 = ~n19401 & n19403;
  assign n19405 = ~n19395 & n19402;
  assign n19406 = ~pi789 & n19389;
  assign n19407 = n59242 & ~n19406;
  assign n19408 = ~n59677 & n19407;
  assign n19409 = ~n19342 & ~n19408;
  assign n19410 = ~n59357 & ~n19409;
  assign n19411 = n7957 & ~n59674;
  assign n19412 = n8065 & n19315;
  assign n19413 = pi629 & ~n19412;
  assign n19414 = ~n19411 & n19413;
  assign n19415 = n7958 & ~n59674;
  assign n19416 = n8074 & n19315;
  assign n19417 = ~pi629 & ~n19416;
  assign n19418 = ~n19415 & n19417;
  assign n19419 = pi792 & ~n19418;
  assign n19420 = ~n19415 & ~n19416;
  assign n19421 = ~pi629 & ~n19420;
  assign n19422 = ~n19411 & ~n19412;
  assign n19423 = pi629 & ~n19422;
  assign n19424 = ~n19421 & ~n19423;
  assign n19425 = pi792 & ~n19424;
  assign n19426 = pi792 & ~n19414;
  assign n19427 = ~n19418 & n19426;
  assign n19428 = ~n19414 & n19419;
  assign n19429 = ~n8108 & ~n59678;
  assign n19430 = ~n19410 & n19429;
  assign n19431 = ~n19328 & ~n19430;
  assign n19432 = pi644 & n19431;
  assign n19433 = ~pi787 & ~n19316;
  assign n19434 = pi1157 & ~n19319;
  assign n19435 = ~n19324 & ~n19434;
  assign n19436 = pi787 & ~n19435;
  assign n19437 = ~n19433 & ~n19436;
  assign n19438 = ~pi644 & n19437;
  assign n19439 = pi715 & ~n19438;
  assign n19440 = ~n19432 & n19439;
  assign n19441 = ~n11491 & n19257;
  assign n19442 = ~n7835 & n19295;
  assign n19443 = ~n7835 & ~n19298;
  assign n19444 = n7835 & n19257;
  assign n19445 = ~n19443 & ~n19444;
  assign n19446 = ~n19441 & ~n19442;
  assign n19447 = pi644 & ~n59679;
  assign n19448 = ~pi644 & n19257;
  assign n19449 = ~pi715 & ~n19448;
  assign n19450 = ~n19447 & n19449;
  assign n19451 = pi1160 & ~n19450;
  assign n19452 = ~n19440 & n19451;
  assign n19453 = ~pi644 & n19431;
  assign n19454 = pi644 & n19437;
  assign n19455 = ~pi715 & ~n19454;
  assign n19456 = ~n19453 & n19455;
  assign n19457 = ~pi644 & ~n59679;
  assign n19458 = pi644 & n19257;
  assign n19459 = pi715 & ~n19458;
  assign n19460 = ~n19457 & n19459;
  assign n19461 = ~pi1160 & ~n19460;
  assign n19462 = ~n19456 & n19461;
  assign n19463 = ~n19452 & ~n19462;
  assign n19464 = pi790 & ~n19463;
  assign n19465 = ~pi790 & n19431;
  assign n19466 = pi832 & ~n19465;
  assign n19467 = ~n19464 & n19466;
  assign n19468 = pi187 & ~n59132;
  assign n19469 = pi770 & n7553;
  assign n19470 = ~pi187 & ~pi770;
  assign n19471 = n9787 & n19470;
  assign n19472 = ~pi770 & ~n13474;
  assign n19473 = pi187 & ~n19472;
  assign n19474 = ~n19471 & ~n19473;
  assign n19475 = pi770 & ~n7553;
  assign n19476 = ~pi770 & ~n9787;
  assign n19477 = ~n19475 & ~n19476;
  assign n19478 = ~pi187 & ~n19477;
  assign n19479 = ~pi187 & ~n9780;
  assign n19480 = ~pi770 & ~n19479;
  assign n19481 = ~n13474 & n19480;
  assign n19482 = ~n19478 & ~n19481;
  assign n19483 = ~n19469 & n19474;
  assign n19484 = n59132 & n59680;
  assign n19485 = ~n19468 & ~n19484;
  assign n19486 = ~n7597 & ~n19485;
  assign n19487 = ~pi187 & ~n7560;
  assign n19488 = n7597 & ~n19487;
  assign n19489 = ~n19486 & ~n19488;
  assign n19490 = ~pi785 & ~n19489;
  assign n19491 = ~n7598 & ~n19487;
  assign n19492 = pi609 & n19486;
  assign n19493 = ~n19491 & ~n19492;
  assign n19494 = pi1155 & ~n19493;
  assign n19495 = ~n7610 & ~n19487;
  assign n19496 = ~pi609 & n19486;
  assign n19497 = ~n19495 & ~n19496;
  assign n19498 = ~pi1155 & ~n19497;
  assign n19499 = ~n19494 & ~n19498;
  assign n19500 = pi785 & ~n19499;
  assign n19501 = ~n19490 & ~n19500;
  assign n19502 = ~pi781 & ~n19501;
  assign n19503 = pi618 & n19501;
  assign n19504 = ~pi618 & n19487;
  assign n19505 = pi1154 & ~n19504;
  assign n19506 = ~n19503 & n19505;
  assign n19507 = ~pi618 & n19501;
  assign n19508 = pi618 & n19487;
  assign n19509 = ~pi1154 & ~n19508;
  assign n19510 = ~n19507 & n19509;
  assign n19511 = ~n19506 & ~n19510;
  assign n19512 = pi781 & ~n19511;
  assign n19513 = ~n19502 & ~n19512;
  assign n19514 = ~pi789 & ~n19513;
  assign n19515 = ~pi619 & n19513;
  assign n19516 = pi619 & n19487;
  assign n19517 = ~pi1159 & ~n19516;
  assign n19518 = ~n19515 & n19517;
  assign n19519 = pi619 & n19513;
  assign n19520 = ~pi619 & n19487;
  assign n19521 = pi1159 & ~n19520;
  assign n19522 = ~n19519 & n19521;
  assign n19523 = ~n19518 & ~n19522;
  assign n19524 = pi789 & ~n19523;
  assign n19525 = ~n19514 & ~n19524;
  assign n19526 = ~n8054 & n19525;
  assign n19527 = n8054 & n19487;
  assign n19528 = ~n19526 & ~n19527;
  assign n19529 = ~n11154 & n19528;
  assign n19530 = n7762 & ~n19487;
  assign n19531 = n59231 & ~n19487;
  assign n19532 = ~pi187 & n8249;
  assign n19533 = pi187 & n59251;
  assign n19534 = ~pi38 & ~n19533;
  assign n19535 = ~n19532 & n19534;
  assign n19536 = ~pi187 & ~n6863;
  assign n19537 = n7547 & ~n19536;
  assign n19538 = pi726 & ~n19537;
  assign n19539 = ~n19535 & n19538;
  assign n19540 = ~pi187 & ~pi726;
  assign n19541 = ~n7553 & n19540;
  assign n19542 = n59132 & ~n19541;
  assign n19543 = ~n19539 & n19542;
  assign n19544 = ~n19468 & ~n19543;
  assign n19545 = ~pi778 & ~n19544;
  assign n19546 = pi625 & n19544;
  assign n19547 = ~pi625 & n19487;
  assign n19548 = pi1153 & ~n19547;
  assign n19549 = ~n19546 & n19548;
  assign n19550 = ~pi625 & n19544;
  assign n19551 = pi625 & n19487;
  assign n19552 = ~pi1153 & ~n19551;
  assign n19553 = ~n19550 & n19552;
  assign n19554 = ~n19549 & ~n19553;
  assign n19555 = pi778 & ~n19554;
  assign n19556 = ~n19545 & ~n19555;
  assign n19557 = ~n59229 & n19556;
  assign n19558 = n59229 & n19487;
  assign n19559 = n59229 & ~n19487;
  assign n19560 = ~n59229 & ~n19556;
  assign n19561 = ~n19559 & ~n19560;
  assign n19562 = ~n19557 & ~n19558;
  assign n19563 = ~n59231 & ~n59681;
  assign n19564 = ~n59231 & n59681;
  assign n19565 = n59231 & n19487;
  assign n19566 = ~n19564 & ~n19565;
  assign n19567 = ~n19531 & ~n19563;
  assign n19568 = ~n7716 & ~n59682;
  assign n19569 = n7716 & n19487;
  assign n19570 = n7716 & ~n19487;
  assign n19571 = ~n7716 & n59682;
  assign n19572 = ~n19570 & ~n19571;
  assign n19573 = ~n19568 & ~n19569;
  assign n19574 = ~n7762 & ~n59683;
  assign n19575 = ~n7762 & n59683;
  assign n19576 = n7762 & n19487;
  assign n19577 = ~n19575 & ~n19576;
  assign n19578 = ~n19530 & ~n19574;
  assign n19579 = ~pi628 & ~n59684;
  assign n19580 = pi628 & n19487;
  assign n19581 = ~pi1156 & ~n19580;
  assign n19582 = ~n19579 & n19581;
  assign n19583 = pi629 & n19582;
  assign n19584 = ~pi628 & ~n19487;
  assign n19585 = pi628 & n59684;
  assign n19586 = ~n19584 & ~n19585;
  assign n19587 = n7790 & ~n19586;
  assign n19588 = ~n19583 & ~n19587;
  assign n19589 = ~n19529 & n19588;
  assign n19590 = pi792 & ~n19589;
  assign n19591 = pi619 & ~n59682;
  assign n19592 = ~pi1159 & ~n19591;
  assign n19593 = ~pi648 & ~n19522;
  assign n19594 = ~n19592 & n19593;
  assign n19595 = ~pi619 & ~n59682;
  assign n19596 = pi1159 & ~n19595;
  assign n19597 = pi648 & ~n19518;
  assign n19598 = ~n19596 & n19597;
  assign n19599 = ~n19594 & ~n19598;
  assign n19600 = pi789 & ~n19599;
  assign n19601 = pi618 & n59681;
  assign n19602 = ~pi1154 & ~n19601;
  assign n19603 = ~pi627 & ~n19506;
  assign n19604 = ~n19602 & n19603;
  assign n19605 = ~pi187 & n9797;
  assign n19606 = pi187 & n9799;
  assign n19607 = pi770 & ~n9801;
  assign n19608 = ~n19606 & n19607;
  assign n19609 = ~n19605 & n19608;
  assign n19610 = pi187 & n9811;
  assign n19611 = ~pi187 & ~n59320;
  assign n19612 = ~pi770 & ~n19611;
  assign n19613 = ~n19610 & n19612;
  assign n19614 = pi726 & ~n19613;
  assign n19615 = ~n19609 & n19614;
  assign n19616 = ~pi726 & ~n59680;
  assign n19617 = n59132 & ~n19616;
  assign n19618 = n59132 & ~n19615;
  assign n19619 = ~n19616 & n19618;
  assign n19620 = ~n19615 & n19617;
  assign n19621 = ~n19468 & ~n59685;
  assign n19622 = ~pi625 & n19621;
  assign n19623 = pi625 & n19485;
  assign n19624 = ~pi1153 & ~n19623;
  assign n19625 = ~n19622 & n19624;
  assign n19626 = ~pi608 & ~n19549;
  assign n19627 = ~n19625 & n19626;
  assign n19628 = pi625 & n19621;
  assign n19629 = ~pi625 & n19485;
  assign n19630 = pi1153 & ~n19629;
  assign n19631 = ~n19628 & n19630;
  assign n19632 = pi608 & ~n19553;
  assign n19633 = ~n19631 & n19632;
  assign n19634 = ~n19627 & ~n19633;
  assign n19635 = pi778 & ~n19634;
  assign n19636 = ~pi778 & n19621;
  assign n19637 = ~pi778 & ~n19621;
  assign n19638 = pi778 & ~n19633;
  assign n19639 = ~n19627 & n19638;
  assign n19640 = ~n19637 & ~n19639;
  assign n19641 = ~n19635 & ~n19636;
  assign n19642 = ~pi609 & n59686;
  assign n19643 = pi609 & n19556;
  assign n19644 = ~pi1155 & ~n19643;
  assign n19645 = ~n19642 & n19644;
  assign n19646 = ~pi660 & ~n19494;
  assign n19647 = ~n19645 & n19646;
  assign n19648 = pi609 & n59686;
  assign n19649 = ~pi609 & n19556;
  assign n19650 = pi1155 & ~n19649;
  assign n19651 = ~n19648 & n19650;
  assign n19652 = pi660 & ~n19498;
  assign n19653 = ~n19651 & n19652;
  assign n19654 = ~n19647 & ~n19653;
  assign n19655 = pi785 & ~n19654;
  assign n19656 = ~pi785 & n59686;
  assign n19657 = ~n19655 & ~n19656;
  assign n19658 = pi618 & ~n19657;
  assign n19659 = ~pi618 & n59681;
  assign n19660 = pi1154 & ~n19659;
  assign n19661 = ~n19658 & n19660;
  assign n19662 = pi627 & ~n19510;
  assign n19663 = ~n19661 & n19662;
  assign n19664 = ~n19604 & ~n19663;
  assign n19665 = pi781 & ~n19664;
  assign n19666 = ~pi618 & n19603;
  assign n19667 = pi781 & ~n19666;
  assign n19668 = ~n19657 & ~n19667;
  assign n19669 = ~pi618 & ~n19657;
  assign n19670 = n19602 & ~n19669;
  assign n19671 = n19603 & ~n19670;
  assign n19672 = ~n19663 & ~n19671;
  assign n19673 = pi781 & ~n19672;
  assign n19674 = ~pi781 & ~n19657;
  assign n19675 = ~n19673 & ~n19674;
  assign n19676 = ~n19665 & ~n19668;
  assign n19677 = ~pi619 & n19593;
  assign n19678 = pi619 & n19597;
  assign n19679 = pi789 & ~n19678;
  assign n19680 = ~n19677 & n19679;
  assign n19681 = ~n59687 & ~n19680;
  assign n19682 = ~pi619 & ~n59687;
  assign n19683 = n19592 & ~n19682;
  assign n19684 = n19593 & ~n19683;
  assign n19685 = pi619 & ~n59687;
  assign n19686 = n19596 & ~n19685;
  assign n19687 = n19597 & ~n19686;
  assign n19688 = ~n19684 & ~n19687;
  assign n19689 = pi789 & ~n19688;
  assign n19690 = ~pi789 & ~n59687;
  assign n19691 = ~n19689 & ~n19690;
  assign n19692 = ~n19600 & ~n19681;
  assign n19693 = n59242 & ~n59688;
  assign n19694 = n12139 & n19525;
  assign n19695 = ~pi641 & ~n59683;
  assign n19696 = pi641 & ~n19487;
  assign n19697 = n7912 & ~n19696;
  assign n19698 = ~n19695 & n19697;
  assign n19699 = pi641 & ~n59683;
  assign n19700 = ~pi641 & ~n19487;
  assign n19701 = n7911 & ~n19700;
  assign n19702 = ~n19699 & n19701;
  assign n19703 = ~n19698 & ~n19702;
  assign n19704 = ~n19694 & n19703;
  assign n19705 = pi788 & ~n19704;
  assign n19706 = ~n59357 & ~n19705;
  assign n19707 = ~n19693 & n19706;
  assign n19708 = ~pi788 & n59688;
  assign n19709 = ~pi626 & n59688;
  assign n19710 = pi626 & ~n59683;
  assign n19711 = ~pi641 & ~n19710;
  assign n19712 = ~n19709 & n19711;
  assign n19713 = ~pi626 & ~n19525;
  assign n19714 = pi626 & ~n19487;
  assign n19715 = pi641 & ~n19714;
  assign n19716 = ~n19713 & n19715;
  assign n19717 = ~pi1158 & ~n19716;
  assign n19718 = ~n19712 & n19717;
  assign n19719 = pi626 & n59688;
  assign n19720 = ~pi626 & ~n59683;
  assign n19721 = pi641 & ~n19720;
  assign n19722 = ~n19719 & n19721;
  assign n19723 = pi626 & ~n19525;
  assign n19724 = ~pi626 & ~n19487;
  assign n19725 = ~pi641 & ~n19724;
  assign n19726 = ~n19723 & n19725;
  assign n19727 = pi1158 & ~n19726;
  assign n19728 = ~n19722 & n19727;
  assign n19729 = ~n19718 & ~n19728;
  assign n19730 = pi788 & ~n19729;
  assign n19731 = ~n19708 & ~n19730;
  assign n19732 = ~pi628 & n19731;
  assign n19733 = pi628 & ~n19528;
  assign n19734 = ~pi1156 & ~n19733;
  assign n19735 = ~n19732 & n19734;
  assign n19736 = pi628 & ~n59684;
  assign n19737 = ~pi628 & n19487;
  assign n19738 = pi1156 & ~n19737;
  assign n19739 = pi1156 & ~n19586;
  assign n19740 = ~n19736 & n19738;
  assign n19741 = ~pi629 & ~n59689;
  assign n19742 = ~n19735 & n19741;
  assign n19743 = pi628 & n19731;
  assign n19744 = ~pi628 & ~n19528;
  assign n19745 = pi1156 & ~n19744;
  assign n19746 = ~n19743 & n19745;
  assign n19747 = pi629 & ~n19582;
  assign n19748 = ~n19746 & n19747;
  assign n19749 = ~n19742 & ~n19748;
  assign n19750 = pi792 & ~n19749;
  assign n19751 = ~pi792 & n19731;
  assign n19752 = ~n19750 & ~n19751;
  assign n19753 = ~n19590 & ~n19707;
  assign n19754 = n59244 & n59690;
  assign n19755 = ~pi647 & ~n19487;
  assign n19756 = ~pi792 & n59684;
  assign n19757 = ~n19582 & ~n59689;
  assign n19758 = pi792 & ~n19757;
  assign n19759 = ~n19756 & ~n19758;
  assign n19760 = pi647 & ~n19759;
  assign n19761 = ~n19755 & ~n19760;
  assign n19762 = n7832 & ~n19761;
  assign n19763 = ~pi647 & n19759;
  assign n19764 = pi647 & n19487;
  assign n19765 = ~pi1157 & ~n19764;
  assign n19766 = ~n19763 & n19765;
  assign n19767 = pi630 & n19766;
  assign n19768 = ~n7793 & ~n19528;
  assign n19769 = n7793 & n19487;
  assign n19770 = ~n19768 & ~n19769;
  assign n19771 = ~n7872 & n19770;
  assign n19772 = ~n19767 & ~n19771;
  assign n19773 = ~n19762 & n19772;
  assign n19774 = ~pi647 & ~n59690;
  assign n19775 = pi647 & ~n19770;
  assign n19776 = ~pi1157 & ~n19775;
  assign n19777 = ~n19774 & n19776;
  assign n19778 = pi647 & n19759;
  assign n19779 = ~pi647 & n19487;
  assign n19780 = pi1157 & ~n19779;
  assign n19781 = pi1157 & ~n19761;
  assign n19782 = ~n19778 & n19780;
  assign n19783 = ~pi630 & ~n59691;
  assign n19784 = ~n19777 & n19783;
  assign n19785 = pi647 & ~n59690;
  assign n19786 = ~pi647 & ~n19770;
  assign n19787 = pi1157 & ~n19786;
  assign n19788 = ~n19785 & n19787;
  assign n19789 = pi630 & ~n19766;
  assign n19790 = ~n19788 & n19789;
  assign n19791 = ~n19784 & ~n19790;
  assign n19792 = ~n19754 & n19773;
  assign n19793 = pi787 & n59692;
  assign n19794 = ~pi787 & n59690;
  assign n19795 = pi787 & ~n59692;
  assign n19796 = ~pi787 & ~n59690;
  assign n19797 = ~n19795 & ~n19796;
  assign n19798 = ~n19793 & ~n19794;
  assign n19799 = pi644 & ~n59693;
  assign n19800 = ~pi787 & ~n19759;
  assign n19801 = ~n19766 & ~n59691;
  assign n19802 = pi787 & ~n19801;
  assign n19803 = ~n19800 & ~n19802;
  assign n19804 = ~pi644 & n19803;
  assign n19805 = pi715 & ~n19804;
  assign n19806 = ~n19799 & n19805;
  assign n19807 = ~n7835 & ~n19770;
  assign n19808 = n7835 & n19487;
  assign n19809 = n7835 & ~n19487;
  assign n19810 = ~n7835 & n19770;
  assign n19811 = ~n19809 & ~n19810;
  assign n19812 = ~n19807 & ~n19808;
  assign n19813 = pi644 & n59694;
  assign n19814 = ~pi644 & n19487;
  assign n19815 = ~pi715 & ~n19814;
  assign n19816 = ~n19813 & n19815;
  assign n19817 = pi1160 & ~n19816;
  assign n19818 = ~n19806 & n19817;
  assign n19819 = ~pi644 & n59694;
  assign n19820 = pi644 & n19487;
  assign n19821 = pi715 & ~n19820;
  assign n19822 = ~n19819 & n19821;
  assign n19823 = ~pi1160 & ~n19822;
  assign n19824 = pi644 & n19803;
  assign n19825 = ~pi715 & ~n19824;
  assign n19826 = ~pi644 & ~n59693;
  assign n19827 = n19825 & ~n19826;
  assign n19828 = n19823 & ~n19827;
  assign n19829 = pi790 & ~n19828;
  assign n19830 = pi790 & ~n19818;
  assign n19831 = ~n19828 & n19830;
  assign n19832 = ~n19818 & n19829;
  assign n19833 = ~pi790 & n59693;
  assign n19834 = n58992 & ~n19833;
  assign n19835 = n19823 & ~n19825;
  assign n19836 = ~n19818 & ~n19835;
  assign n19837 = pi790 & ~n19836;
  assign n19838 = ~pi644 & n19823;
  assign n19839 = pi790 & ~n19838;
  assign n19840 = ~n59693 & ~n19839;
  assign n19841 = ~n19837 & ~n19840;
  assign n19842 = n58992 & ~n19841;
  assign n19843 = ~n59695 & n19834;
  assign n19844 = ~pi187 & ~n58992;
  assign n19845 = ~pi832 & ~n19844;
  assign n19846 = ~n59696 & n19845;
  assign po344 = ~n19467 & ~n19846;
  assign n19848 = ~pi188 & ~n2794;
  assign n19849 = ~pi768 & n6822;
  assign n19850 = ~n19848 & ~n19849;
  assign n19851 = ~n7875 & ~n19850;
  assign n19852 = ~pi785 & ~n19851;
  assign n19853 = ~n7880 & ~n19850;
  assign n19854 = pi1155 & ~n19853;
  assign n19855 = ~n7883 & n19851;
  assign n19856 = ~pi1155 & ~n19855;
  assign n19857 = ~n19854 & ~n19856;
  assign n19858 = pi785 & ~n19857;
  assign n19859 = ~n19852 & ~n19858;
  assign n19860 = ~pi781 & ~n19859;
  assign n19861 = ~n7890 & n19859;
  assign n19862 = pi1154 & ~n19861;
  assign n19863 = ~n7893 & n19859;
  assign n19864 = ~pi1154 & ~n19863;
  assign n19865 = ~n19862 & ~n19864;
  assign n19866 = pi781 & ~n19865;
  assign n19867 = ~n19860 & ~n19866;
  assign n19868 = ~pi789 & ~n19867;
  assign n19869 = pi619 & n19867;
  assign n19870 = ~pi619 & n19848;
  assign n19871 = pi1159 & ~n19870;
  assign n19872 = ~n19869 & n19871;
  assign n19873 = ~pi619 & n19867;
  assign n19874 = pi619 & n19848;
  assign n19875 = ~pi1159 & ~n19874;
  assign n19876 = ~n19873 & n19875;
  assign n19877 = ~n19872 & ~n19876;
  assign n19878 = pi789 & ~n19877;
  assign n19879 = ~n19868 & ~n19878;
  assign n19880 = ~n8054 & ~n19879;
  assign n19881 = n8054 & ~n19848;
  assign n19882 = ~n8054 & n19879;
  assign n19883 = n8054 & n19848;
  assign n19884 = ~n19882 & ~n19883;
  assign n19885 = ~n19880 & ~n19881;
  assign n19886 = ~n7793 & ~n59697;
  assign n19887 = n7793 & n19848;
  assign n19888 = ~n7872 & ~n19887;
  assign n19889 = ~n19886 & ~n19887;
  assign n19890 = ~n7872 & n19889;
  assign n19891 = ~n19886 & n19888;
  assign n19892 = pi705 & n7055;
  assign n19893 = ~n19848 & ~n19892;
  assign n19894 = ~pi778 & n19893;
  assign n19895 = ~pi625 & n19892;
  assign n19896 = ~n19893 & ~n19895;
  assign n19897 = pi1153 & ~n19896;
  assign n19898 = ~pi1153 & ~n19848;
  assign n19899 = ~n19895 & n19898;
  assign n19900 = ~n19897 & ~n19899;
  assign n19901 = pi778 & ~n19900;
  assign n19902 = ~n19894 & ~n19901;
  assign n19903 = ~n7949 & n19902;
  assign n19904 = ~n7951 & n19903;
  assign n19905 = ~n7953 & n19904;
  assign n19906 = ~n7955 & n19905;
  assign n19907 = ~n7967 & n19906;
  assign n19908 = pi647 & ~n19907;
  assign n19909 = ~pi647 & ~n19848;
  assign n19910 = ~n19908 & ~n19909;
  assign n19911 = n7832 & ~n19910;
  assign n19912 = ~pi647 & n19907;
  assign n19913 = pi647 & n19848;
  assign n19914 = ~pi1157 & ~n19913;
  assign n19915 = ~n19912 & n19914;
  assign n19916 = pi630 & n19915;
  assign n19917 = ~n19911 & ~n19916;
  assign n19918 = ~n59698 & n19917;
  assign n19919 = pi787 & ~n19918;
  assign n19920 = ~pi626 & ~n19879;
  assign n19921 = pi626 & ~n19848;
  assign n19922 = n7760 & ~n19921;
  assign n19923 = ~n19920 & n19922;
  assign n19924 = n7984 & n19905;
  assign n19925 = pi626 & ~n19879;
  assign n19926 = ~pi626 & ~n19848;
  assign n19927 = n7759 & ~n19926;
  assign n19928 = ~n19925 & n19927;
  assign n19929 = ~n19924 & ~n19928;
  assign n19930 = ~n19923 & ~n19924;
  assign n19931 = ~n19928 & n19930;
  assign n19932 = ~n19923 & n19929;
  assign n19933 = pi788 & ~n59699;
  assign n19934 = ~n6701 & ~n19893;
  assign n19935 = pi625 & n19934;
  assign n19936 = n19850 & ~n19934;
  assign n19937 = ~n19935 & ~n19936;
  assign n19938 = n19898 & ~n19937;
  assign n19939 = ~pi608 & ~n19897;
  assign n19940 = ~n19938 & n19939;
  assign n19941 = pi1153 & n19850;
  assign n19942 = ~n19935 & n19941;
  assign n19943 = pi608 & ~n19899;
  assign n19944 = ~n19942 & n19943;
  assign n19945 = ~n19940 & ~n19944;
  assign n19946 = pi778 & ~n19945;
  assign n19947 = ~pi778 & ~n19936;
  assign n19948 = ~n19946 & ~n19947;
  assign n19949 = ~pi609 & ~n19948;
  assign n19950 = pi609 & n19902;
  assign n19951 = ~pi1155 & ~n19950;
  assign n19952 = ~n19949 & n19951;
  assign n19953 = ~pi660 & ~n19854;
  assign n19954 = ~n19952 & n19953;
  assign n19955 = pi609 & ~n19948;
  assign n19956 = ~pi609 & n19902;
  assign n19957 = pi1155 & ~n19956;
  assign n19958 = ~n19955 & n19957;
  assign n19959 = pi660 & ~n19856;
  assign n19960 = ~n19958 & n19959;
  assign n19961 = ~n19954 & ~n19960;
  assign n19962 = pi785 & ~n19961;
  assign n19963 = ~pi785 & ~n19948;
  assign n19964 = ~n19962 & ~n19963;
  assign n19965 = ~pi618 & ~n19964;
  assign n19966 = pi618 & n19903;
  assign n19967 = ~pi1154 & ~n19966;
  assign n19968 = ~n19965 & n19967;
  assign n19969 = ~pi627 & ~n19862;
  assign n19970 = ~n19968 & n19969;
  assign n19971 = pi618 & ~n19964;
  assign n19972 = ~pi618 & n19903;
  assign n19973 = pi1154 & ~n19972;
  assign n19974 = ~n19971 & n19973;
  assign n19975 = pi627 & ~n19864;
  assign n19976 = ~n19974 & n19975;
  assign n19977 = ~n19970 & ~n19976;
  assign n19978 = pi781 & ~n19977;
  assign n19979 = ~pi781 & ~n19964;
  assign n19980 = ~n19978 & ~n19979;
  assign n19981 = ~pi619 & ~n19980;
  assign n19982 = pi619 & n19904;
  assign n19983 = ~pi1159 & ~n19982;
  assign n19984 = ~n19981 & n19983;
  assign n19985 = ~pi648 & ~n19872;
  assign n19986 = ~n19984 & n19985;
  assign n19987 = pi619 & ~n19980;
  assign n19988 = ~pi619 & n19904;
  assign n19989 = pi1159 & ~n19988;
  assign n19990 = ~n19987 & n19989;
  assign n19991 = pi648 & ~n19876;
  assign n19992 = ~n19990 & n19991;
  assign n19993 = pi789 & ~n19992;
  assign n19994 = pi789 & ~n19986;
  assign n19995 = ~n19992 & n19994;
  assign n19996 = ~n19986 & n19993;
  assign n19997 = ~pi789 & n19980;
  assign n19998 = n59242 & ~n19997;
  assign n19999 = ~n59700 & n19998;
  assign n20000 = ~n19933 & ~n19999;
  assign n20001 = ~n59357 & ~n20000;
  assign n20002 = n7957 & ~n59697;
  assign n20003 = n8065 & n19906;
  assign n20004 = pi629 & ~n20003;
  assign n20005 = ~n20002 & n20004;
  assign n20006 = n7958 & ~n59697;
  assign n20007 = n8074 & n19906;
  assign n20008 = ~pi629 & ~n20007;
  assign n20009 = ~n20006 & n20008;
  assign n20010 = pi792 & ~n20009;
  assign n20011 = ~n20006 & ~n20007;
  assign n20012 = ~pi629 & ~n20011;
  assign n20013 = ~n20002 & ~n20003;
  assign n20014 = pi629 & ~n20013;
  assign n20015 = ~n20012 & ~n20014;
  assign n20016 = pi792 & ~n20015;
  assign n20017 = pi792 & ~n20005;
  assign n20018 = ~n20009 & n20017;
  assign n20019 = ~n20005 & n20010;
  assign n20020 = ~n8108 & ~n59701;
  assign n20021 = ~n20001 & n20020;
  assign n20022 = ~n19919 & ~n20021;
  assign n20023 = pi644 & n20022;
  assign n20024 = ~pi787 & ~n19907;
  assign n20025 = pi1157 & ~n19910;
  assign n20026 = ~n19915 & ~n20025;
  assign n20027 = pi787 & ~n20026;
  assign n20028 = ~n20024 & ~n20027;
  assign n20029 = ~pi644 & n20028;
  assign n20030 = pi715 & ~n20029;
  assign n20031 = ~n20023 & n20030;
  assign n20032 = ~n11491 & n19848;
  assign n20033 = ~n7835 & n19886;
  assign n20034 = ~n7835 & ~n19889;
  assign n20035 = n7835 & n19848;
  assign n20036 = ~n20034 & ~n20035;
  assign n20037 = ~n20032 & ~n20033;
  assign n20038 = pi644 & ~n59702;
  assign n20039 = ~pi644 & n19848;
  assign n20040 = ~pi715 & ~n20039;
  assign n20041 = ~n20038 & n20040;
  assign n20042 = pi1160 & ~n20041;
  assign n20043 = ~n20031 & n20042;
  assign n20044 = ~pi644 & n20022;
  assign n20045 = pi644 & n20028;
  assign n20046 = ~pi715 & ~n20045;
  assign n20047 = ~n20044 & n20046;
  assign n20048 = ~pi644 & ~n59702;
  assign n20049 = pi644 & n19848;
  assign n20050 = pi715 & ~n20049;
  assign n20051 = ~n20048 & n20050;
  assign n20052 = ~pi1160 & ~n20051;
  assign n20053 = ~n20047 & n20052;
  assign n20054 = ~n20043 & ~n20053;
  assign n20055 = pi790 & ~n20054;
  assign n20056 = ~pi790 & n20022;
  assign n20057 = pi832 & ~n20056;
  assign n20058 = ~n20055 & n20057;
  assign n20059 = pi188 & ~n59132;
  assign n20060 = pi768 & n7553;
  assign n20061 = ~pi768 & ~n13474;
  assign n20062 = pi188 & ~n20061;
  assign n20063 = ~pi188 & ~pi768;
  assign n20064 = n9787 & n20063;
  assign n20065 = ~n20062 & ~n20064;
  assign n20066 = pi768 & ~n7553;
  assign n20067 = ~pi768 & ~n9787;
  assign n20068 = ~n20066 & ~n20067;
  assign n20069 = ~pi188 & ~n20068;
  assign n20070 = ~pi188 & ~n9780;
  assign n20071 = ~pi768 & ~n20070;
  assign n20072 = ~n13474 & n20071;
  assign n20073 = ~n20069 & ~n20072;
  assign n20074 = ~n20060 & n20065;
  assign n20075 = n59132 & n59703;
  assign n20076 = ~n20059 & ~n20075;
  assign n20077 = ~n7597 & ~n20076;
  assign n20078 = ~pi188 & ~n7560;
  assign n20079 = n7597 & ~n20078;
  assign n20080 = ~n20077 & ~n20079;
  assign n20081 = ~pi785 & ~n20080;
  assign n20082 = ~n7598 & ~n20078;
  assign n20083 = pi609 & n20077;
  assign n20084 = ~n20082 & ~n20083;
  assign n20085 = pi1155 & ~n20084;
  assign n20086 = ~n7610 & ~n20078;
  assign n20087 = ~pi609 & n20077;
  assign n20088 = ~n20086 & ~n20087;
  assign n20089 = ~pi1155 & ~n20088;
  assign n20090 = ~n20085 & ~n20089;
  assign n20091 = pi785 & ~n20090;
  assign n20092 = ~n20081 & ~n20091;
  assign n20093 = ~pi781 & ~n20092;
  assign n20094 = pi618 & n20092;
  assign n20095 = ~pi618 & n20078;
  assign n20096 = pi1154 & ~n20095;
  assign n20097 = ~n20094 & n20096;
  assign n20098 = ~pi618 & n20092;
  assign n20099 = pi618 & n20078;
  assign n20100 = ~pi1154 & ~n20099;
  assign n20101 = ~n20098 & n20100;
  assign n20102 = ~n20097 & ~n20101;
  assign n20103 = pi781 & ~n20102;
  assign n20104 = ~n20093 & ~n20103;
  assign n20105 = ~pi789 & ~n20104;
  assign n20106 = ~pi619 & n20104;
  assign n20107 = pi619 & n20078;
  assign n20108 = ~pi1159 & ~n20107;
  assign n20109 = ~n20106 & n20108;
  assign n20110 = pi619 & n20104;
  assign n20111 = ~pi619 & n20078;
  assign n20112 = pi1159 & ~n20111;
  assign n20113 = ~n20110 & n20112;
  assign n20114 = ~n20109 & ~n20113;
  assign n20115 = pi789 & ~n20114;
  assign n20116 = ~n20105 & ~n20115;
  assign n20117 = ~n8054 & n20116;
  assign n20118 = n8054 & n20078;
  assign n20119 = ~n20117 & ~n20118;
  assign n20120 = ~n11154 & n20119;
  assign n20121 = n7762 & ~n20078;
  assign n20122 = n59231 & ~n20078;
  assign n20123 = ~pi188 & n8249;
  assign n20124 = pi188 & n59251;
  assign n20125 = ~pi38 & ~n20124;
  assign n20126 = ~n20123 & n20125;
  assign n20127 = ~pi188 & ~n6863;
  assign n20128 = n7547 & ~n20127;
  assign n20129 = pi705 & ~n20128;
  assign n20130 = ~n20126 & n20129;
  assign n20131 = ~pi188 & ~pi705;
  assign n20132 = ~n7553 & n20131;
  assign n20133 = n59132 & ~n20132;
  assign n20134 = ~n20130 & n20133;
  assign n20135 = ~n20059 & ~n20134;
  assign n20136 = ~pi778 & ~n20135;
  assign n20137 = pi625 & n20135;
  assign n20138 = ~pi625 & n20078;
  assign n20139 = pi1153 & ~n20138;
  assign n20140 = ~n20137 & n20139;
  assign n20141 = ~pi625 & n20135;
  assign n20142 = pi625 & n20078;
  assign n20143 = ~pi1153 & ~n20142;
  assign n20144 = ~n20141 & n20143;
  assign n20145 = ~n20140 & ~n20144;
  assign n20146 = pi778 & ~n20145;
  assign n20147 = ~n20136 & ~n20146;
  assign n20148 = ~n59229 & n20147;
  assign n20149 = n59229 & n20078;
  assign n20150 = n59229 & ~n20078;
  assign n20151 = ~n59229 & ~n20147;
  assign n20152 = ~n20150 & ~n20151;
  assign n20153 = ~n20148 & ~n20149;
  assign n20154 = ~n59231 & ~n59704;
  assign n20155 = ~n59231 & n59704;
  assign n20156 = n59231 & n20078;
  assign n20157 = ~n20155 & ~n20156;
  assign n20158 = ~n20122 & ~n20154;
  assign n20159 = ~n7716 & ~n59705;
  assign n20160 = n7716 & n20078;
  assign n20161 = n7716 & ~n20078;
  assign n20162 = ~n7716 & n59705;
  assign n20163 = ~n20161 & ~n20162;
  assign n20164 = ~n20159 & ~n20160;
  assign n20165 = ~n7762 & ~n59706;
  assign n20166 = ~n7762 & n59706;
  assign n20167 = n7762 & n20078;
  assign n20168 = ~n20166 & ~n20167;
  assign n20169 = ~n20121 & ~n20165;
  assign n20170 = ~pi628 & ~n59707;
  assign n20171 = pi628 & n20078;
  assign n20172 = ~pi1156 & ~n20171;
  assign n20173 = ~n20170 & n20172;
  assign n20174 = pi629 & n20173;
  assign n20175 = ~pi628 & ~n20078;
  assign n20176 = pi628 & n59707;
  assign n20177 = ~n20175 & ~n20176;
  assign n20178 = n7790 & ~n20177;
  assign n20179 = ~n20174 & ~n20178;
  assign n20180 = ~n20120 & n20179;
  assign n20181 = pi792 & ~n20180;
  assign n20182 = pi619 & ~n59705;
  assign n20183 = ~pi1159 & ~n20182;
  assign n20184 = ~pi648 & ~n20113;
  assign n20185 = ~n20183 & n20184;
  assign n20186 = ~pi619 & ~n59705;
  assign n20187 = pi1159 & ~n20186;
  assign n20188 = pi648 & ~n20109;
  assign n20189 = ~n20187 & n20188;
  assign n20190 = ~n20185 & ~n20189;
  assign n20191 = pi789 & ~n20190;
  assign n20192 = pi618 & n59704;
  assign n20193 = ~pi1154 & ~n20192;
  assign n20194 = ~pi627 & ~n20097;
  assign n20195 = ~n20193 & n20194;
  assign n20196 = ~pi188 & n9797;
  assign n20197 = pi188 & n9799;
  assign n20198 = pi768 & ~n9801;
  assign n20199 = ~n20197 & n20198;
  assign n20200 = ~n20196 & n20199;
  assign n20201 = pi188 & n9811;
  assign n20202 = ~pi188 & ~n59320;
  assign n20203 = ~pi768 & ~n20202;
  assign n20204 = ~n20201 & n20203;
  assign n20205 = pi705 & ~n20204;
  assign n20206 = ~n20200 & n20205;
  assign n20207 = ~pi705 & ~n59703;
  assign n20208 = n59132 & ~n20207;
  assign n20209 = n59132 & ~n20206;
  assign n20210 = ~n20207 & n20209;
  assign n20211 = ~n20206 & n20208;
  assign n20212 = ~n20059 & ~n59708;
  assign n20213 = ~pi625 & n20212;
  assign n20214 = pi625 & n20076;
  assign n20215 = ~pi1153 & ~n20214;
  assign n20216 = ~n20213 & n20215;
  assign n20217 = ~pi608 & ~n20140;
  assign n20218 = ~n20216 & n20217;
  assign n20219 = pi625 & n20212;
  assign n20220 = ~pi625 & n20076;
  assign n20221 = pi1153 & ~n20220;
  assign n20222 = ~n20219 & n20221;
  assign n20223 = pi608 & ~n20144;
  assign n20224 = ~n20222 & n20223;
  assign n20225 = ~n20218 & ~n20224;
  assign n20226 = pi778 & ~n20225;
  assign n20227 = ~pi778 & n20212;
  assign n20228 = ~pi778 & ~n20212;
  assign n20229 = pi778 & ~n20224;
  assign n20230 = ~n20218 & n20229;
  assign n20231 = ~n20228 & ~n20230;
  assign n20232 = ~n20226 & ~n20227;
  assign n20233 = ~pi609 & n59709;
  assign n20234 = pi609 & n20147;
  assign n20235 = ~pi1155 & ~n20234;
  assign n20236 = ~n20233 & n20235;
  assign n20237 = ~pi660 & ~n20085;
  assign n20238 = ~n20236 & n20237;
  assign n20239 = pi609 & n59709;
  assign n20240 = ~pi609 & n20147;
  assign n20241 = pi1155 & ~n20240;
  assign n20242 = ~n20239 & n20241;
  assign n20243 = pi660 & ~n20089;
  assign n20244 = ~n20242 & n20243;
  assign n20245 = ~n20238 & ~n20244;
  assign n20246 = pi785 & ~n20245;
  assign n20247 = ~pi785 & n59709;
  assign n20248 = ~n20246 & ~n20247;
  assign n20249 = pi618 & ~n20248;
  assign n20250 = ~pi618 & n59704;
  assign n20251 = pi1154 & ~n20250;
  assign n20252 = ~n20249 & n20251;
  assign n20253 = pi627 & ~n20101;
  assign n20254 = ~n20252 & n20253;
  assign n20255 = ~n20195 & ~n20254;
  assign n20256 = pi781 & ~n20255;
  assign n20257 = ~pi618 & n20194;
  assign n20258 = pi781 & ~n20257;
  assign n20259 = ~n20248 & ~n20258;
  assign n20260 = ~pi618 & ~n20248;
  assign n20261 = n20193 & ~n20260;
  assign n20262 = n20194 & ~n20261;
  assign n20263 = ~n20254 & ~n20262;
  assign n20264 = pi781 & ~n20263;
  assign n20265 = ~pi781 & ~n20248;
  assign n20266 = ~n20264 & ~n20265;
  assign n20267 = ~n20256 & ~n20259;
  assign n20268 = ~pi619 & n20184;
  assign n20269 = pi619 & n20188;
  assign n20270 = pi789 & ~n20269;
  assign n20271 = ~n20268 & n20270;
  assign n20272 = ~n59710 & ~n20271;
  assign n20273 = ~pi619 & ~n59710;
  assign n20274 = n20183 & ~n20273;
  assign n20275 = n20184 & ~n20274;
  assign n20276 = pi619 & ~n59710;
  assign n20277 = n20187 & ~n20276;
  assign n20278 = n20188 & ~n20277;
  assign n20279 = ~n20275 & ~n20278;
  assign n20280 = pi789 & ~n20279;
  assign n20281 = ~pi789 & ~n59710;
  assign n20282 = ~n20280 & ~n20281;
  assign n20283 = ~n20191 & ~n20272;
  assign n20284 = n59242 & ~n59711;
  assign n20285 = n12139 & n20116;
  assign n20286 = ~pi641 & ~n59706;
  assign n20287 = pi641 & ~n20078;
  assign n20288 = n7912 & ~n20287;
  assign n20289 = ~n20286 & n20288;
  assign n20290 = pi641 & ~n59706;
  assign n20291 = ~pi641 & ~n20078;
  assign n20292 = n7911 & ~n20291;
  assign n20293 = ~n20290 & n20292;
  assign n20294 = ~n20289 & ~n20293;
  assign n20295 = ~n20285 & n20294;
  assign n20296 = pi788 & ~n20295;
  assign n20297 = ~n59357 & ~n20296;
  assign n20298 = ~n20284 & n20297;
  assign n20299 = ~pi788 & n59711;
  assign n20300 = ~pi626 & n59711;
  assign n20301 = pi626 & ~n59706;
  assign n20302 = ~pi641 & ~n20301;
  assign n20303 = ~n20300 & n20302;
  assign n20304 = ~pi626 & ~n20116;
  assign n20305 = pi626 & ~n20078;
  assign n20306 = pi641 & ~n20305;
  assign n20307 = ~n20304 & n20306;
  assign n20308 = ~pi1158 & ~n20307;
  assign n20309 = ~n20303 & n20308;
  assign n20310 = pi626 & n59711;
  assign n20311 = ~pi626 & ~n59706;
  assign n20312 = pi641 & ~n20311;
  assign n20313 = ~n20310 & n20312;
  assign n20314 = pi626 & ~n20116;
  assign n20315 = ~pi626 & ~n20078;
  assign n20316 = ~pi641 & ~n20315;
  assign n20317 = ~n20314 & n20316;
  assign n20318 = pi1158 & ~n20317;
  assign n20319 = ~n20313 & n20318;
  assign n20320 = ~n20309 & ~n20319;
  assign n20321 = pi788 & ~n20320;
  assign n20322 = ~n20299 & ~n20321;
  assign n20323 = ~pi628 & n20322;
  assign n20324 = pi628 & ~n20119;
  assign n20325 = ~pi1156 & ~n20324;
  assign n20326 = ~n20323 & n20325;
  assign n20327 = pi628 & ~n59707;
  assign n20328 = ~pi628 & n20078;
  assign n20329 = pi1156 & ~n20328;
  assign n20330 = pi1156 & ~n20177;
  assign n20331 = ~n20327 & n20329;
  assign n20332 = ~pi629 & ~n59712;
  assign n20333 = ~n20326 & n20332;
  assign n20334 = pi628 & n20322;
  assign n20335 = ~pi628 & ~n20119;
  assign n20336 = pi1156 & ~n20335;
  assign n20337 = ~n20334 & n20336;
  assign n20338 = pi629 & ~n20173;
  assign n20339 = ~n20337 & n20338;
  assign n20340 = ~n20333 & ~n20339;
  assign n20341 = pi792 & ~n20340;
  assign n20342 = ~pi792 & n20322;
  assign n20343 = ~n20341 & ~n20342;
  assign n20344 = ~n20181 & ~n20298;
  assign n20345 = n59244 & n59713;
  assign n20346 = ~pi647 & ~n20078;
  assign n20347 = ~pi792 & n59707;
  assign n20348 = ~n20173 & ~n59712;
  assign n20349 = pi792 & ~n20348;
  assign n20350 = ~n20347 & ~n20349;
  assign n20351 = pi647 & ~n20350;
  assign n20352 = ~n20346 & ~n20351;
  assign n20353 = n7832 & ~n20352;
  assign n20354 = ~pi647 & n20350;
  assign n20355 = pi647 & n20078;
  assign n20356 = ~pi1157 & ~n20355;
  assign n20357 = ~n20354 & n20356;
  assign n20358 = pi630 & n20357;
  assign n20359 = ~n7793 & ~n20119;
  assign n20360 = n7793 & n20078;
  assign n20361 = ~n20359 & ~n20360;
  assign n20362 = ~n7872 & n20361;
  assign n20363 = ~n20358 & ~n20362;
  assign n20364 = ~n20353 & n20363;
  assign n20365 = ~pi647 & ~n59713;
  assign n20366 = pi647 & ~n20361;
  assign n20367 = ~pi1157 & ~n20366;
  assign n20368 = ~n20365 & n20367;
  assign n20369 = pi647 & n20350;
  assign n20370 = ~pi647 & n20078;
  assign n20371 = pi1157 & ~n20370;
  assign n20372 = pi1157 & ~n20352;
  assign n20373 = ~n20369 & n20371;
  assign n20374 = ~pi630 & ~n59714;
  assign n20375 = ~n20368 & n20374;
  assign n20376 = pi647 & ~n59713;
  assign n20377 = ~pi647 & ~n20361;
  assign n20378 = pi1157 & ~n20377;
  assign n20379 = ~n20376 & n20378;
  assign n20380 = pi630 & ~n20357;
  assign n20381 = ~n20379 & n20380;
  assign n20382 = ~n20375 & ~n20381;
  assign n20383 = ~n20345 & n20364;
  assign n20384 = pi787 & n59715;
  assign n20385 = ~pi787 & n59713;
  assign n20386 = pi787 & ~n59715;
  assign n20387 = ~pi787 & ~n59713;
  assign n20388 = ~n20386 & ~n20387;
  assign n20389 = ~n20384 & ~n20385;
  assign n20390 = pi644 & ~n59716;
  assign n20391 = ~pi787 & ~n20350;
  assign n20392 = ~n20357 & ~n59714;
  assign n20393 = pi787 & ~n20392;
  assign n20394 = ~n20391 & ~n20393;
  assign n20395 = ~pi644 & n20394;
  assign n20396 = pi715 & ~n20395;
  assign n20397 = ~n20390 & n20396;
  assign n20398 = ~n7835 & ~n20361;
  assign n20399 = n7835 & n20078;
  assign n20400 = n7835 & ~n20078;
  assign n20401 = ~n7835 & n20361;
  assign n20402 = ~n20400 & ~n20401;
  assign n20403 = ~n20398 & ~n20399;
  assign n20404 = pi644 & n59717;
  assign n20405 = ~pi644 & n20078;
  assign n20406 = ~pi715 & ~n20405;
  assign n20407 = ~n20404 & n20406;
  assign n20408 = pi1160 & ~n20407;
  assign n20409 = ~n20397 & n20408;
  assign n20410 = ~pi644 & n59717;
  assign n20411 = pi644 & n20078;
  assign n20412 = pi715 & ~n20411;
  assign n20413 = ~n20410 & n20412;
  assign n20414 = ~pi1160 & ~n20413;
  assign n20415 = pi644 & n20394;
  assign n20416 = ~pi715 & ~n20415;
  assign n20417 = ~pi644 & ~n59716;
  assign n20418 = n20416 & ~n20417;
  assign n20419 = n20414 & ~n20418;
  assign n20420 = pi790 & ~n20419;
  assign n20421 = pi790 & ~n20409;
  assign n20422 = ~n20419 & n20421;
  assign n20423 = ~n20409 & n20420;
  assign n20424 = ~pi790 & n59716;
  assign n20425 = n58992 & ~n20424;
  assign n20426 = n20414 & ~n20416;
  assign n20427 = ~n20409 & ~n20426;
  assign n20428 = pi790 & ~n20427;
  assign n20429 = ~pi644 & n20414;
  assign n20430 = pi790 & ~n20429;
  assign n20431 = ~n59716 & ~n20430;
  assign n20432 = ~n20428 & ~n20431;
  assign n20433 = n58992 & ~n20432;
  assign n20434 = ~n59718 & n20425;
  assign n20435 = ~pi188 & ~n58992;
  assign n20436 = ~pi832 & ~n20435;
  assign n20437 = ~n59719 & n20436;
  assign po345 = ~n20058 & ~n20437;
  assign n20439 = pi727 & n7055;
  assign n20440 = pi727 & n7056;
  assign n20441 = ~n6701 & n20439;
  assign n20442 = pi189 & ~n2794;
  assign n20443 = pi772 & n6822;
  assign n20444 = ~n20442 & ~n20443;
  assign n20445 = ~n59720 & n20444;
  assign n20446 = pi625 & n20439;
  assign n20447 = pi625 & n59720;
  assign n20448 = ~n6701 & n20446;
  assign n20449 = ~n20445 & ~n59721;
  assign n20450 = ~pi1153 & ~n20449;
  assign n20451 = pi1153 & ~n20442;
  assign n20452 = ~n20446 & n20451;
  assign n20453 = ~pi608 & ~n20452;
  assign n20454 = ~n20450 & n20453;
  assign n20455 = pi1153 & n20444;
  assign n20456 = ~n20443 & n20451;
  assign n20457 = ~n59721 & n59722;
  assign n20458 = ~n20439 & ~n20442;
  assign n20459 = ~n20446 & ~n20458;
  assign n20460 = ~pi1153 & ~n20459;
  assign n20461 = pi608 & ~n20460;
  assign n20462 = ~n20457 & n20461;
  assign n20463 = ~n20454 & ~n20462;
  assign n20464 = pi778 & ~n20463;
  assign n20465 = ~pi778 & ~n20445;
  assign n20466 = ~n20464 & ~n20465;
  assign n20467 = ~pi609 & ~n20466;
  assign n20468 = ~pi778 & n20458;
  assign n20469 = ~n20452 & ~n20460;
  assign n20470 = pi778 & ~n20469;
  assign n20471 = ~n20468 & ~n20470;
  assign n20472 = pi609 & n20471;
  assign n20473 = ~pi1155 & ~n20472;
  assign n20474 = ~n20467 & n20473;
  assign n20475 = n7598 & n20443;
  assign n20476 = pi1155 & ~n20442;
  assign n20477 = ~n20475 & n20476;
  assign n20478 = ~pi660 & ~n20477;
  assign n20479 = ~n20474 & n20478;
  assign n20480 = pi609 & ~n20466;
  assign n20481 = ~pi609 & n20471;
  assign n20482 = pi1155 & ~n20481;
  assign n20483 = ~n20480 & n20482;
  assign n20484 = n7610 & n20443;
  assign n20485 = ~pi1155 & ~n20442;
  assign n20486 = ~n20484 & n20485;
  assign n20487 = pi660 & ~n20486;
  assign n20488 = ~n20483 & n20487;
  assign n20489 = ~n20479 & ~n20488;
  assign n20490 = pi785 & ~n20489;
  assign n20491 = ~pi785 & ~n20466;
  assign n20492 = ~n20490 & ~n20491;
  assign n20493 = pi618 & ~n20492;
  assign n20494 = ~n59229 & n20471;
  assign n20495 = ~n20442 & ~n20494;
  assign n20496 = ~pi618 & ~n20495;
  assign n20497 = pi1154 & ~n20496;
  assign n20498 = ~n20493 & n20497;
  assign n20499 = ~n59346 & n20443;
  assign n20500 = n10837 & n20499;
  assign n20501 = ~pi1154 & ~n20442;
  assign n20502 = ~n20500 & n20501;
  assign n20503 = pi627 & ~n20502;
  assign n20504 = ~n20498 & n20503;
  assign n20505 = ~pi618 & ~n20492;
  assign n20506 = pi618 & ~n20495;
  assign n20507 = ~pi1154 & ~n20506;
  assign n20508 = ~n20505 & n20507;
  assign n20509 = n10835 & n20499;
  assign n20510 = pi1154 & ~n20442;
  assign n20511 = ~n20509 & n20510;
  assign n20512 = ~pi627 & ~n20511;
  assign n20513 = ~n20508 & n20512;
  assign n20514 = ~n20504 & ~n20513;
  assign n20515 = pi781 & ~n20514;
  assign n20516 = ~pi781 & ~n20492;
  assign n20517 = ~n12513 & ~n20516;
  assign n20518 = ~n20515 & n20517;
  assign n20519 = n9554 & n20471;
  assign n20520 = ~n12510 & ~n20519;
  assign n20521 = ~n59347 & n20499;
  assign n20522 = ~n7715 & ~n20521;
  assign n20523 = n10884 & n20521;
  assign n20524 = n7714 & ~n20523;
  assign n20525 = n10874 & n20521;
  assign n20526 = n7713 & ~n20525;
  assign n20527 = ~n20524 & ~n20526;
  assign n20528 = ~n12521 & ~n20522;
  assign n20529 = ~n20520 & n59723;
  assign n20530 = pi789 & ~n20442;
  assign n20531 = ~n20529 & n20530;
  assign n20532 = n59242 & ~n20531;
  assign n20533 = ~n20518 & n20532;
  assign n20534 = ~n7716 & n20519;
  assign n20535 = ~n20442 & ~n20534;
  assign n20536 = n7911 & ~n20535;
  assign n20537 = n59348 & n20499;
  assign n20538 = ~pi626 & n20537;
  assign n20539 = ~n20442 & ~n20538;
  assign n20540 = ~pi1158 & ~n20539;
  assign n20541 = pi641 & ~n20540;
  assign n20542 = ~n20536 & n20541;
  assign n20543 = n7912 & ~n20535;
  assign n20544 = pi626 & n20537;
  assign n20545 = ~n20442 & ~n20544;
  assign n20546 = pi1158 & ~n20545;
  assign n20547 = ~pi641 & ~n20546;
  assign n20548 = ~n20543 & n20547;
  assign n20549 = pi788 & ~n20548;
  assign n20550 = pi788 & ~n20542;
  assign n20551 = ~n20548 & n20550;
  assign n20552 = ~n20542 & n20549;
  assign n20553 = ~n59357 & ~n59724;
  assign n20554 = ~n20533 & n20553;
  assign n20555 = ~n8054 & n20537;
  assign n20556 = ~pi629 & n20555;
  assign n20557 = pi628 & ~n20556;
  assign n20558 = ~n7762 & n20534;
  assign n20559 = n9652 & n20471;
  assign n20560 = pi629 & ~n59725;
  assign n20561 = ~pi628 & n59725;
  assign n20562 = pi629 & ~n20561;
  assign n20563 = pi628 & ~n20555;
  assign n20564 = ~n20562 & ~n20563;
  assign n20565 = ~n20557 & ~n20560;
  assign n20566 = ~pi1156 & ~n59726;
  assign n20567 = pi628 & n59725;
  assign n20568 = ~pi628 & ~n20555;
  assign n20569 = pi629 & ~n20568;
  assign n20570 = pi1156 & ~n20569;
  assign n20571 = ~n20567 & n20570;
  assign n20572 = ~n20566 & ~n20571;
  assign n20573 = pi792 & ~n20442;
  assign n20574 = ~n20572 & n20573;
  assign n20575 = ~n20554 & ~n20574;
  assign n20576 = ~n8108 & ~n20575;
  assign n20577 = ~n59240 & n59725;
  assign n20578 = ~pi630 & ~n20577;
  assign n20579 = pi647 & ~n20578;
  assign n20580 = ~n7793 & n20555;
  assign n20581 = pi630 & n20580;
  assign n20582 = pi1157 & ~n20581;
  assign n20583 = ~n20579 & n20582;
  assign n20584 = pi630 & ~n20577;
  assign n20585 = ~pi647 & ~n20584;
  assign n20586 = ~pi630 & n20580;
  assign n20587 = ~pi1157 & ~n20586;
  assign n20588 = pi647 & ~n20586;
  assign n20589 = ~n20584 & ~n20588;
  assign n20590 = ~pi1157 & ~n20589;
  assign n20591 = ~n20585 & n20587;
  assign n20592 = ~n20583 & ~n59727;
  assign n20593 = pi787 & ~n20442;
  assign n20594 = ~n20592 & n20593;
  assign n20595 = ~n20576 & ~n20594;
  assign n20596 = pi644 & n20595;
  assign n20597 = ~n9743 & n20577;
  assign n20598 = ~n20442 & ~n20597;
  assign n20599 = ~pi644 & ~n20598;
  assign n20600 = pi715 & ~n20599;
  assign n20601 = ~n20596 & n20600;
  assign n20602 = n12602 & n20537;
  assign n20603 = pi644 & n20602;
  assign n20604 = ~pi715 & ~n20442;
  assign n20605 = ~n20603 & n20604;
  assign n20606 = pi1160 & ~n20605;
  assign n20607 = ~n20601 & n20606;
  assign n20608 = ~pi644 & n20595;
  assign n20609 = pi644 & ~n20598;
  assign n20610 = ~pi715 & ~n20609;
  assign n20611 = ~n20608 & n20610;
  assign n20612 = ~pi644 & n20602;
  assign n20613 = pi715 & ~n20442;
  assign n20614 = ~n20612 & n20613;
  assign n20615 = ~pi1160 & ~n20614;
  assign n20616 = ~n20611 & n20615;
  assign n20617 = ~n20607 & ~n20616;
  assign n20618 = pi790 & ~n20617;
  assign n20619 = ~pi790 & n20595;
  assign n20620 = pi832 & ~n20619;
  assign n20621 = ~n20618 & n20620;
  assign n20622 = pi189 & ~n59132;
  assign n20623 = ~pi772 & ~n6654;
  assign n20624 = pi772 & n59163;
  assign n20625 = ~n20623 & ~n20624;
  assign n20626 = pi39 & ~n20625;
  assign n20627 = pi772 & n59157;
  assign n20628 = ~pi772 & n59147;
  assign n20629 = ~pi39 & ~n20628;
  assign n20630 = ~n20627 & n20629;
  assign n20631 = ~n20626 & ~n20630;
  assign n20632 = pi189 & ~n20631;
  assign n20633 = ~pi189 & pi772;
  assign n20634 = n6855 & n20633;
  assign n20635 = ~n20632 & ~n20634;
  assign n20636 = ~pi38 & ~n20635;
  assign n20637 = pi772 & n6701;
  assign n20638 = n6863 & ~n20637;
  assign n20639 = ~pi189 & ~n6863;
  assign n20640 = pi38 & ~n20639;
  assign n20641 = ~n20638 & n20640;
  assign n20642 = ~n20636 & ~n20641;
  assign n20643 = n59132 & ~n20642;
  assign n20644 = ~n20622 & ~n20643;
  assign n20645 = ~n7597 & ~n20644;
  assign n20646 = pi189 & ~n7560;
  assign n20647 = n7597 & n20646;
  assign n20648 = n7597 & ~n20646;
  assign n20649 = ~n7597 & n20644;
  assign n20650 = ~n20648 & ~n20649;
  assign n20651 = ~n20645 & ~n20647;
  assign n20652 = ~pi785 & n59728;
  assign n20653 = pi609 & ~n59728;
  assign n20654 = ~pi609 & ~n20646;
  assign n20655 = pi1155 & ~n20654;
  assign n20656 = ~n20653 & n20655;
  assign n20657 = ~pi609 & ~n59728;
  assign n20658 = pi609 & ~n20646;
  assign n20659 = ~pi1155 & ~n20658;
  assign n20660 = ~n20657 & n20659;
  assign n20661 = ~n20656 & ~n20660;
  assign n20662 = pi785 & ~n20661;
  assign n20663 = ~n20652 & ~n20662;
  assign n20664 = ~pi781 & ~n20663;
  assign n20665 = pi618 & n20663;
  assign n20666 = ~pi618 & ~n20646;
  assign n20667 = pi1154 & ~n20666;
  assign n20668 = ~n20665 & n20667;
  assign n20669 = ~pi618 & n20663;
  assign n20670 = pi618 & ~n20646;
  assign n20671 = ~pi1154 & ~n20670;
  assign n20672 = ~n20669 & n20671;
  assign n20673 = ~n20668 & ~n20672;
  assign n20674 = pi781 & ~n20673;
  assign n20675 = ~n20664 & ~n20674;
  assign n20676 = ~pi789 & ~n20675;
  assign n20677 = pi619 & n20675;
  assign n20678 = ~pi619 & ~n20646;
  assign n20679 = pi1159 & ~n20678;
  assign n20680 = ~n20677 & n20679;
  assign n20681 = ~pi619 & n20675;
  assign n20682 = pi619 & ~n20646;
  assign n20683 = ~pi1159 & ~n20682;
  assign n20684 = ~n20681 & n20683;
  assign n20685 = ~n20680 & ~n20684;
  assign n20686 = pi789 & ~n20685;
  assign n20687 = ~n20676 & ~n20686;
  assign n20688 = ~n8054 & ~n20687;
  assign n20689 = n8054 & n20646;
  assign n20690 = ~n20688 & ~n20689;
  assign n20691 = ~n11154 & ~n20690;
  assign n20692 = n7762 & ~n20646;
  assign n20693 = n59231 & ~n20646;
  assign n20694 = pi727 & n59132;
  assign n20695 = ~n20646 & ~n20694;
  assign n20696 = pi189 & ~n8249;
  assign n20697 = ~pi189 & ~n59251;
  assign n20698 = ~pi38 & ~n20697;
  assign n20699 = ~n20696 & n20698;
  assign n20700 = n10432 & ~n20639;
  assign n20701 = n20694 & ~n20700;
  assign n20702 = ~n20699 & n20701;
  assign n20703 = ~n20695 & ~n20702;
  assign n20704 = ~pi778 & n20703;
  assign n20705 = pi625 & ~n20703;
  assign n20706 = ~pi625 & ~n20646;
  assign n20707 = pi1153 & ~n20706;
  assign n20708 = ~n20705 & n20707;
  assign n20709 = ~pi625 & ~n20703;
  assign n20710 = pi625 & ~n20646;
  assign n20711 = ~pi1153 & ~n20710;
  assign n20712 = ~n20709 & n20711;
  assign n20713 = ~n20708 & ~n20712;
  assign n20714 = pi778 & ~n20713;
  assign n20715 = ~n20704 & ~n20714;
  assign n20716 = ~n59229 & ~n20715;
  assign n20717 = n59229 & n20646;
  assign n20718 = n59229 & ~n20646;
  assign n20719 = ~n59229 & n20715;
  assign n20720 = ~n20718 & ~n20719;
  assign n20721 = ~n20716 & ~n20717;
  assign n20722 = ~n59231 & ~n59729;
  assign n20723 = ~n59231 & n59729;
  assign n20724 = n59231 & n20646;
  assign n20725 = ~n20723 & ~n20724;
  assign n20726 = ~n20693 & ~n20722;
  assign n20727 = ~n7716 & ~n59730;
  assign n20728 = n7716 & n20646;
  assign n20729 = n7716 & ~n20646;
  assign n20730 = ~n7716 & n59730;
  assign n20731 = ~n20729 & ~n20730;
  assign n20732 = ~n20727 & ~n20728;
  assign n20733 = ~n7762 & ~n59731;
  assign n20734 = ~n7762 & n59731;
  assign n20735 = n7762 & n20646;
  assign n20736 = ~n20734 & ~n20735;
  assign n20737 = ~n20692 & ~n20733;
  assign n20738 = ~pi628 & n59732;
  assign n20739 = pi628 & ~n20646;
  assign n20740 = ~pi1156 & ~n20739;
  assign n20741 = ~n20738 & n20740;
  assign n20742 = pi629 & n20741;
  assign n20743 = pi628 & ~n59732;
  assign n20744 = ~pi628 & n20646;
  assign n20745 = ~n20743 & ~n20744;
  assign n20746 = n7790 & ~n20745;
  assign n20747 = ~n20742 & ~n20746;
  assign n20748 = ~n20691 & n20747;
  assign n20749 = pi792 & ~n20748;
  assign n20750 = pi619 & n59730;
  assign n20751 = ~pi1159 & ~n20750;
  assign n20752 = ~pi648 & ~n20680;
  assign n20753 = ~n20751 & n20752;
  assign n20754 = ~pi619 & n59730;
  assign n20755 = pi1159 & ~n20754;
  assign n20756 = pi648 & ~n20684;
  assign n20757 = ~n20755 & n20756;
  assign n20758 = ~n20753 & ~n20757;
  assign n20759 = pi789 & ~n20758;
  assign n20760 = ~pi727 & n20636;
  assign n20761 = pi189 & ~n59177;
  assign n20762 = ~pi189 & ~n7111;
  assign n20763 = ~pi772 & ~n20762;
  assign n20764 = ~n20761 & n20763;
  assign n20765 = ~pi189 & ~n7188;
  assign n20766 = pi189 & n59203;
  assign n20767 = pi772 & ~n20766;
  assign n20768 = ~n20765 & n20767;
  assign n20769 = pi39 & ~n20768;
  assign n20770 = ~n20764 & n20769;
  assign n20771 = ~pi189 & ~n7333;
  assign n20772 = pi189 & ~n7310;
  assign n20773 = ~pi772 & ~n20772;
  assign n20774 = ~pi772 & ~n20771;
  assign n20775 = ~n20772 & n20774;
  assign n20776 = ~n20771 & n20773;
  assign n20777 = pi189 & n7339;
  assign n20778 = ~pi189 & n7347;
  assign n20779 = pi772 & ~n20778;
  assign n20780 = ~n20777 & n20779;
  assign n20781 = ~pi39 & ~n20780;
  assign n20782 = ~n59733 & n20781;
  assign n20783 = ~pi38 & ~n20782;
  assign n20784 = ~n20770 & n20783;
  assign n20785 = ~n9801 & ~n20784;
  assign n20786 = pi727 & ~n20785;
  assign n20787 = ~n20641 & ~n20786;
  assign n20788 = ~n20760 & n20787;
  assign n20789 = ~pi727 & n20642;
  assign n20790 = pi727 & ~n9801;
  assign n20791 = ~n20641 & n20790;
  assign n20792 = ~n20784 & n20791;
  assign n20793 = n59132 & ~n20792;
  assign n20794 = ~n20789 & n20793;
  assign n20795 = n59132 & ~n20788;
  assign n20796 = ~n20622 & ~n59734;
  assign n20797 = ~pi625 & n20796;
  assign n20798 = pi625 & n20644;
  assign n20799 = ~pi1153 & ~n20798;
  assign n20800 = ~n20797 & n20799;
  assign n20801 = ~pi608 & ~n20708;
  assign n20802 = ~n20800 & n20801;
  assign n20803 = pi625 & n20796;
  assign n20804 = ~pi625 & n20644;
  assign n20805 = pi1153 & ~n20804;
  assign n20806 = ~n20803 & n20805;
  assign n20807 = pi608 & ~n20712;
  assign n20808 = ~n20806 & n20807;
  assign n20809 = ~n20802 & ~n20808;
  assign n20810 = pi778 & ~n20809;
  assign n20811 = ~pi778 & n20796;
  assign n20812 = ~n20810 & ~n20811;
  assign n20813 = ~pi609 & ~n20812;
  assign n20814 = pi609 & n20715;
  assign n20815 = ~pi1155 & ~n20814;
  assign n20816 = ~n20813 & n20815;
  assign n20817 = ~pi660 & ~n20656;
  assign n20818 = ~n20816 & n20817;
  assign n20819 = pi609 & ~n20812;
  assign n20820 = ~pi609 & n20715;
  assign n20821 = pi1155 & ~n20820;
  assign n20822 = ~n20819 & n20821;
  assign n20823 = pi660 & ~n20660;
  assign n20824 = ~n20822 & n20823;
  assign n20825 = ~n20818 & ~n20824;
  assign n20826 = pi785 & ~n20825;
  assign n20827 = ~pi785 & ~n20812;
  assign n20828 = ~n20826 & ~n20827;
  assign n20829 = pi618 & ~n20828;
  assign n20830 = ~pi618 & ~n59729;
  assign n20831 = pi1154 & ~n20830;
  assign n20832 = ~n20829 & n20831;
  assign n20833 = pi627 & ~n20672;
  assign n20834 = ~n20832 & n20833;
  assign n20835 = ~pi618 & ~n20828;
  assign n20836 = pi618 & ~n59729;
  assign n20837 = ~pi1154 & ~n20836;
  assign n20838 = ~n20835 & n20837;
  assign n20839 = ~pi627 & ~n20668;
  assign n20840 = ~n20838 & n20839;
  assign n20841 = pi781 & ~n20840;
  assign n20842 = ~n20834 & n20841;
  assign n20843 = ~pi619 & n20752;
  assign n20844 = pi619 & n20756;
  assign n20845 = pi789 & ~n20844;
  assign n20846 = ~n20843 & n20845;
  assign n20847 = ~pi781 & n20828;
  assign n20848 = ~n20846 & ~n20847;
  assign n20849 = ~n20842 & n20848;
  assign n20850 = ~n20834 & ~n20840;
  assign n20851 = pi781 & ~n20850;
  assign n20852 = ~pi781 & ~n20828;
  assign n20853 = ~n20851 & ~n20852;
  assign n20854 = ~pi619 & ~n20853;
  assign n20855 = n20751 & ~n20854;
  assign n20856 = n20752 & ~n20855;
  assign n20857 = pi619 & ~n20853;
  assign n20858 = n20755 & ~n20857;
  assign n20859 = n20756 & ~n20858;
  assign n20860 = ~n20856 & ~n20859;
  assign n20861 = pi789 & ~n20860;
  assign n20862 = ~pi789 & ~n20853;
  assign n20863 = ~n20861 & ~n20862;
  assign n20864 = ~n20759 & ~n20849;
  assign n20865 = n59242 & ~n59735;
  assign n20866 = n12139 & n20687;
  assign n20867 = ~pi641 & n59731;
  assign n20868 = pi641 & n20646;
  assign n20869 = n7912 & ~n20868;
  assign n20870 = ~n20867 & n20869;
  assign n20871 = pi641 & n59731;
  assign n20872 = ~pi641 & n20646;
  assign n20873 = n7911 & ~n20872;
  assign n20874 = ~n20871 & n20873;
  assign n20875 = ~n20870 & ~n20874;
  assign n20876 = ~n20866 & n20875;
  assign n20877 = pi788 & ~n20876;
  assign n20878 = ~n59357 & ~n20877;
  assign n20879 = ~n20865 & n20878;
  assign n20880 = ~pi788 & n59735;
  assign n20881 = ~pi626 & n59735;
  assign n20882 = pi626 & n59731;
  assign n20883 = ~pi641 & ~n20882;
  assign n20884 = ~n20881 & n20883;
  assign n20885 = ~pi626 & ~n20687;
  assign n20886 = pi626 & n20646;
  assign n20887 = pi641 & ~n20886;
  assign n20888 = ~n20885 & n20887;
  assign n20889 = ~pi1158 & ~n20888;
  assign n20890 = ~n20884 & n20889;
  assign n20891 = pi626 & n59735;
  assign n20892 = ~pi626 & n59731;
  assign n20893 = pi641 & ~n20892;
  assign n20894 = ~n20891 & n20893;
  assign n20895 = pi626 & ~n20687;
  assign n20896 = ~pi626 & n20646;
  assign n20897 = ~pi641 & ~n20896;
  assign n20898 = ~n20895 & n20897;
  assign n20899 = pi1158 & ~n20898;
  assign n20900 = ~n20894 & n20899;
  assign n20901 = ~n20890 & ~n20900;
  assign n20902 = pi788 & ~n20901;
  assign n20903 = ~n20880 & ~n20902;
  assign n20904 = ~pi628 & n20903;
  assign n20905 = pi628 & n20690;
  assign n20906 = ~pi1156 & ~n20905;
  assign n20907 = ~n20904 & n20906;
  assign n20908 = pi628 & n59732;
  assign n20909 = ~pi628 & ~n20646;
  assign n20910 = pi1156 & ~n20909;
  assign n20911 = pi1156 & ~n20745;
  assign n20912 = ~n20908 & n20910;
  assign n20913 = ~pi629 & ~n59736;
  assign n20914 = ~n20907 & n20913;
  assign n20915 = pi628 & n20903;
  assign n20916 = ~pi628 & n20690;
  assign n20917 = pi1156 & ~n20916;
  assign n20918 = ~n20915 & n20917;
  assign n20919 = pi629 & ~n20741;
  assign n20920 = ~n20918 & n20919;
  assign n20921 = ~n20914 & ~n20920;
  assign n20922 = pi792 & ~n20921;
  assign n20923 = ~pi792 & n20903;
  assign n20924 = ~n20922 & ~n20923;
  assign n20925 = ~n20749 & ~n20879;
  assign n20926 = ~n8108 & n59737;
  assign n20927 = ~n7793 & ~n20690;
  assign n20928 = n7793 & n20646;
  assign n20929 = ~n20927 & ~n20928;
  assign n20930 = ~n7872 & ~n20929;
  assign n20931 = ~pi792 & ~n59732;
  assign n20932 = ~n20741 & ~n59736;
  assign n20933 = pi792 & ~n20932;
  assign n20934 = ~n20931 & ~n20933;
  assign n20935 = pi647 & n20934;
  assign n20936 = ~pi647 & ~n20646;
  assign n20937 = pi1157 & ~n20936;
  assign n20938 = ~n20935 & n20937;
  assign n20939 = ~pi630 & n20938;
  assign n20940 = pi647 & ~n20646;
  assign n20941 = ~pi647 & n20934;
  assign n20942 = ~n20940 & ~n20941;
  assign n20943 = n7833 & n20942;
  assign n20944 = ~n20939 & ~n20943;
  assign n20945 = ~n20930 & n20944;
  assign n20946 = pi787 & ~n20945;
  assign n20947 = ~pi647 & ~n59737;
  assign n20948 = pi647 & n20929;
  assign n20949 = ~pi1157 & ~n20948;
  assign n20950 = ~n20947 & n20949;
  assign n20951 = ~pi630 & ~n20938;
  assign n20952 = ~n20950 & n20951;
  assign n20953 = pi647 & ~n59737;
  assign n20954 = ~pi647 & n20929;
  assign n20955 = pi1157 & ~n20954;
  assign n20956 = ~n20953 & n20955;
  assign n20957 = ~pi1157 & ~n20940;
  assign n20958 = ~pi1157 & n20942;
  assign n20959 = ~n20941 & n20957;
  assign n20960 = pi630 & ~n59738;
  assign n20961 = ~n20956 & n20960;
  assign n20962 = ~n20952 & ~n20961;
  assign n20963 = pi787 & ~n20962;
  assign n20964 = ~pi787 & ~n59737;
  assign n20965 = ~n20963 & ~n20964;
  assign n20966 = ~n20926 & ~n20946;
  assign n20967 = pi644 & ~n59739;
  assign n20968 = ~pi787 & ~n20934;
  assign n20969 = ~n20938 & ~n59738;
  assign n20970 = pi787 & ~n20969;
  assign n20971 = ~n20968 & ~n20970;
  assign n20972 = ~pi644 & n20971;
  assign n20973 = pi715 & ~n20972;
  assign n20974 = ~n20967 & n20973;
  assign n20975 = ~n7835 & ~n20929;
  assign n20976 = n7835 & n20646;
  assign n20977 = n7835 & ~n20646;
  assign n20978 = ~n7835 & n20929;
  assign n20979 = ~n20977 & ~n20978;
  assign n20980 = ~n20975 & ~n20976;
  assign n20981 = pi644 & ~n59740;
  assign n20982 = ~pi644 & ~n20646;
  assign n20983 = ~pi715 & ~n20982;
  assign n20984 = ~n20981 & n20983;
  assign n20985 = pi1160 & ~n20984;
  assign n20986 = ~n20974 & n20985;
  assign n20987 = ~pi644 & ~n59740;
  assign n20988 = pi644 & ~n20646;
  assign n20989 = pi715 & ~n20988;
  assign n20990 = ~n20987 & n20989;
  assign n20991 = ~pi1160 & ~n20990;
  assign n20992 = pi644 & n20971;
  assign n20993 = ~pi715 & ~n20992;
  assign n20994 = ~pi644 & ~n59739;
  assign n20995 = n20993 & ~n20994;
  assign n20996 = n20991 & ~n20995;
  assign n20997 = pi790 & ~n20996;
  assign n20998 = pi790 & ~n20986;
  assign n20999 = ~n20996 & n20998;
  assign n21000 = ~n20986 & n20997;
  assign n21001 = ~pi790 & n59739;
  assign n21002 = n4441 & ~n21001;
  assign n21003 = n20991 & ~n20993;
  assign n21004 = ~n20986 & ~n21003;
  assign n21005 = pi790 & ~n21004;
  assign n21006 = ~pi644 & n20991;
  assign n21007 = pi790 & ~n21006;
  assign n21008 = ~n59739 & ~n21007;
  assign n21009 = ~n21005 & ~n21008;
  assign n21010 = n4441 & ~n21009;
  assign n21011 = ~n59741 & n21002;
  assign n21012 = ~pi189 & ~n4441;
  assign n21013 = ~pi57 & ~n21012;
  assign n21014 = ~n59742 & n21013;
  assign n21015 = pi57 & pi189;
  assign n21016 = ~pi832 & ~n21015;
  assign n21017 = ~n21014 & n21016;
  assign po346 = ~n20621 & ~n21017;
  assign n21019 = ~pi190 & ~n2794;
  assign n21020 = pi763 & n6822;
  assign n21021 = ~n21019 & ~n21020;
  assign n21022 = ~n7875 & ~n21021;
  assign n21023 = ~pi785 & ~n21022;
  assign n21024 = n7610 & n21020;
  assign n21025 = n21022 & ~n21024;
  assign n21026 = pi1155 & ~n21025;
  assign n21027 = ~pi1155 & ~n21019;
  assign n21028 = ~n21024 & n21027;
  assign n21029 = ~n21026 & ~n21028;
  assign n21030 = pi785 & ~n21029;
  assign n21031 = ~n21023 & ~n21030;
  assign n21032 = ~pi781 & ~n21031;
  assign n21033 = ~n7890 & n21031;
  assign n21034 = pi1154 & ~n21033;
  assign n21035 = ~n7893 & n21031;
  assign n21036 = ~pi1154 & ~n21035;
  assign n21037 = ~n21034 & ~n21036;
  assign n21038 = pi781 & ~n21037;
  assign n21039 = ~n21032 & ~n21038;
  assign n21040 = ~pi789 & ~n21039;
  assign n21041 = ~n11882 & n21039;
  assign n21042 = pi1159 & ~n21041;
  assign n21043 = ~n11885 & n21039;
  assign n21044 = ~pi1159 & ~n21043;
  assign n21045 = ~n21042 & ~n21044;
  assign n21046 = pi789 & ~n21045;
  assign n21047 = ~n21040 & ~n21046;
  assign n21048 = ~n8054 & ~n21047;
  assign n21049 = n8054 & ~n21019;
  assign n21050 = ~n8054 & n21047;
  assign n21051 = n8054 & n21019;
  assign n21052 = ~n21050 & ~n21051;
  assign n21053 = ~n21048 & ~n21049;
  assign n21054 = ~n7793 & ~n59743;
  assign n21055 = n7793 & n21019;
  assign n21056 = ~n7872 & ~n21055;
  assign n21057 = ~n21054 & ~n21055;
  assign n21058 = ~n7872 & n21057;
  assign n21059 = ~n21054 & n21056;
  assign n21060 = pi699 & n7055;
  assign n21061 = ~n21019 & ~n21060;
  assign n21062 = ~pi778 & ~n21061;
  assign n21063 = ~pi625 & n21060;
  assign n21064 = ~n21061 & ~n21063;
  assign n21065 = pi1153 & ~n21064;
  assign n21066 = ~pi1153 & ~n21019;
  assign n21067 = ~n21063 & n21066;
  assign n21068 = pi778 & ~n21067;
  assign n21069 = ~n21065 & n21068;
  assign n21070 = ~n21062 & ~n21069;
  assign n21071 = ~n7949 & ~n21070;
  assign n21072 = ~n7951 & n21071;
  assign n21073 = ~n7953 & n21072;
  assign n21074 = ~n7955 & n21073;
  assign n21075 = ~n7967 & n21074;
  assign n21076 = pi647 & ~n21075;
  assign n21077 = ~pi647 & ~n21019;
  assign n21078 = ~n21076 & ~n21077;
  assign n21079 = n7832 & ~n21078;
  assign n21080 = ~pi647 & n21075;
  assign n21081 = pi647 & n21019;
  assign n21082 = ~pi1157 & ~n21081;
  assign n21083 = ~n21080 & n21082;
  assign n21084 = pi630 & n21083;
  assign n21085 = ~n21079 & ~n21084;
  assign n21086 = ~n59744 & n21085;
  assign n21087 = pi787 & ~n21086;
  assign n21088 = ~pi626 & ~n21047;
  assign n21089 = pi626 & ~n21019;
  assign n21090 = n7760 & ~n21089;
  assign n21091 = ~n21088 & n21090;
  assign n21092 = n7984 & n21073;
  assign n21093 = pi626 & ~n21047;
  assign n21094 = ~pi626 & ~n21019;
  assign n21095 = n7759 & ~n21094;
  assign n21096 = ~n21093 & n21095;
  assign n21097 = ~n21092 & ~n21096;
  assign n21098 = ~n21091 & ~n21092;
  assign n21099 = ~n21096 & n21098;
  assign n21100 = ~n21091 & n21097;
  assign n21101 = pi788 & ~n59745;
  assign n21102 = ~n6701 & ~n21061;
  assign n21103 = pi625 & n21102;
  assign n21104 = n21021 & ~n21102;
  assign n21105 = ~n21103 & ~n21104;
  assign n21106 = n21066 & ~n21105;
  assign n21107 = ~pi608 & ~n21065;
  assign n21108 = ~n21106 & n21107;
  assign n21109 = pi1153 & n21021;
  assign n21110 = ~n21103 & n21109;
  assign n21111 = pi608 & ~n21067;
  assign n21112 = ~n21110 & n21111;
  assign n21113 = ~n21108 & ~n21112;
  assign n21114 = pi778 & ~n21113;
  assign n21115 = ~pi778 & ~n21104;
  assign n21116 = ~n21114 & ~n21115;
  assign n21117 = ~pi609 & ~n21116;
  assign n21118 = pi609 & ~n21070;
  assign n21119 = ~pi1155 & ~n21118;
  assign n21120 = ~n21117 & n21119;
  assign n21121 = ~pi660 & ~n21026;
  assign n21122 = ~n21120 & n21121;
  assign n21123 = pi609 & ~n21116;
  assign n21124 = ~pi609 & ~n21070;
  assign n21125 = pi1155 & ~n21124;
  assign n21126 = ~n21123 & n21125;
  assign n21127 = pi660 & ~n21028;
  assign n21128 = ~n21126 & n21127;
  assign n21129 = ~n21122 & ~n21128;
  assign n21130 = pi785 & ~n21129;
  assign n21131 = ~pi785 & ~n21116;
  assign n21132 = ~n21130 & ~n21131;
  assign n21133 = ~pi618 & ~n21132;
  assign n21134 = pi618 & n21071;
  assign n21135 = ~pi1154 & ~n21134;
  assign n21136 = ~n21133 & n21135;
  assign n21137 = ~pi627 & ~n21034;
  assign n21138 = ~n21136 & n21137;
  assign n21139 = pi618 & ~n21132;
  assign n21140 = ~pi618 & n21071;
  assign n21141 = pi1154 & ~n21140;
  assign n21142 = ~n21139 & n21141;
  assign n21143 = pi627 & ~n21036;
  assign n21144 = ~n21142 & n21143;
  assign n21145 = ~n21138 & ~n21144;
  assign n21146 = pi781 & ~n21145;
  assign n21147 = ~pi781 & ~n21132;
  assign n21148 = ~n21146 & ~n21147;
  assign n21149 = pi619 & ~n21148;
  assign n21150 = ~pi619 & n21072;
  assign n21151 = pi1159 & ~n21150;
  assign n21152 = ~n21149 & n21151;
  assign n21153 = pi648 & ~n21044;
  assign n21154 = ~n21152 & n21153;
  assign n21155 = ~pi619 & ~n21148;
  assign n21156 = pi619 & n21072;
  assign n21157 = ~pi1159 & ~n21156;
  assign n21158 = ~n21155 & n21157;
  assign n21159 = ~pi648 & ~n21042;
  assign n21160 = ~n21158 & n21159;
  assign n21161 = pi789 & ~n21160;
  assign n21162 = pi789 & ~n21154;
  assign n21163 = ~n21160 & n21162;
  assign n21164 = ~n21154 & n21161;
  assign n21165 = ~pi789 & n21148;
  assign n21166 = n59242 & ~n21165;
  assign n21167 = ~n59746 & n21166;
  assign n21168 = ~n21101 & ~n21167;
  assign n21169 = ~n59357 & ~n21168;
  assign n21170 = n7957 & ~n59743;
  assign n21171 = n8065 & n21074;
  assign n21172 = pi629 & ~n21171;
  assign n21173 = ~n21170 & n21172;
  assign n21174 = n7958 & ~n59743;
  assign n21175 = n8074 & n21074;
  assign n21176 = ~pi629 & ~n21175;
  assign n21177 = ~n21174 & n21176;
  assign n21178 = pi792 & ~n21177;
  assign n21179 = ~n21174 & ~n21175;
  assign n21180 = ~pi629 & ~n21179;
  assign n21181 = ~n21170 & ~n21171;
  assign n21182 = pi629 & ~n21181;
  assign n21183 = ~n21180 & ~n21182;
  assign n21184 = pi792 & ~n21183;
  assign n21185 = pi792 & ~n21173;
  assign n21186 = ~n21177 & n21185;
  assign n21187 = ~n21173 & n21178;
  assign n21188 = ~n8108 & ~n59747;
  assign n21189 = ~n21169 & n21188;
  assign n21190 = ~n21087 & ~n21189;
  assign n21191 = pi644 & n21190;
  assign n21192 = ~pi787 & ~n21075;
  assign n21193 = pi1157 & ~n21078;
  assign n21194 = ~n21083 & ~n21193;
  assign n21195 = pi787 & ~n21194;
  assign n21196 = ~n21192 & ~n21195;
  assign n21197 = ~pi644 & n21196;
  assign n21198 = pi715 & ~n21197;
  assign n21199 = ~n21191 & n21198;
  assign n21200 = ~n11491 & n21019;
  assign n21201 = ~n7835 & n21054;
  assign n21202 = ~n7835 & ~n21057;
  assign n21203 = n7835 & n21019;
  assign n21204 = ~n21202 & ~n21203;
  assign n21205 = ~n21200 & ~n21201;
  assign n21206 = pi644 & ~n59748;
  assign n21207 = ~pi644 & n21019;
  assign n21208 = ~pi715 & ~n21207;
  assign n21209 = ~n21206 & n21208;
  assign n21210 = pi1160 & ~n21209;
  assign n21211 = ~n21199 & n21210;
  assign n21212 = ~pi644 & n21190;
  assign n21213 = pi644 & n21196;
  assign n21214 = ~pi715 & ~n21213;
  assign n21215 = ~n21212 & n21214;
  assign n21216 = ~pi644 & ~n59748;
  assign n21217 = pi644 & n21019;
  assign n21218 = pi715 & ~n21217;
  assign n21219 = ~n21216 & n21218;
  assign n21220 = ~pi1160 & ~n21219;
  assign n21221 = ~n21215 & n21220;
  assign n21222 = ~n21211 & ~n21221;
  assign n21223 = pi790 & ~n21222;
  assign n21224 = ~pi790 & n21190;
  assign n21225 = pi832 & ~n21224;
  assign n21226 = ~n21223 & n21225;
  assign n21227 = ~pi190 & ~n7560;
  assign n21228 = n59231 & ~n21227;
  assign n21229 = pi190 & ~n59132;
  assign n21230 = ~pi190 & n8249;
  assign n21231 = pi190 & n59251;
  assign n21232 = ~pi38 & ~n21231;
  assign n21233 = ~n21230 & n21232;
  assign n21234 = ~pi190 & ~n6863;
  assign n21235 = n7547 & ~n21234;
  assign n21236 = pi699 & ~n21235;
  assign n21237 = ~n21233 & n21236;
  assign n21238 = ~pi190 & ~pi699;
  assign n21239 = ~n7553 & n21238;
  assign n21240 = n59132 & ~n21239;
  assign n21241 = ~n21237 & n21240;
  assign n21242 = ~n21229 & ~n21241;
  assign n21243 = ~pi778 & ~n21242;
  assign n21244 = pi625 & n21242;
  assign n21245 = ~pi625 & n21227;
  assign n21246 = pi1153 & ~n21245;
  assign n21247 = ~n21244 & n21246;
  assign n21248 = ~pi625 & n21242;
  assign n21249 = pi625 & n21227;
  assign n21250 = ~pi1153 & ~n21249;
  assign n21251 = ~n21248 & n21250;
  assign n21252 = ~n21247 & ~n21251;
  assign n21253 = pi778 & ~n21252;
  assign n21254 = ~n21243 & ~n21253;
  assign n21255 = ~n59229 & n21254;
  assign n21256 = n59229 & n21227;
  assign n21257 = n59229 & ~n21227;
  assign n21258 = ~n59229 & ~n21254;
  assign n21259 = ~n21257 & ~n21258;
  assign n21260 = ~n21255 & ~n21256;
  assign n21261 = ~n59231 & ~n59749;
  assign n21262 = ~n59231 & n59749;
  assign n21263 = n59231 & n21227;
  assign n21264 = ~n21262 & ~n21263;
  assign n21265 = ~n21228 & ~n21261;
  assign n21266 = ~n7716 & ~n59750;
  assign n21267 = n7716 & n21227;
  assign n21268 = n7716 & ~n21227;
  assign n21269 = ~n7716 & n59750;
  assign n21270 = ~n21268 & ~n21269;
  assign n21271 = ~n21266 & ~n21267;
  assign n21272 = ~n7762 & n59751;
  assign n21273 = n7762 & n21227;
  assign n21274 = ~n21272 & ~n21273;
  assign n21275 = ~n59240 & ~n21274;
  assign n21276 = n59240 & n21227;
  assign n21277 = ~pi628 & ~n21274;
  assign n21278 = pi628 & n21227;
  assign n21279 = ~n21277 & ~n21278;
  assign n21280 = ~pi1156 & ~n21279;
  assign n21281 = pi628 & ~n21274;
  assign n21282 = ~pi628 & n21227;
  assign n21283 = ~n21281 & ~n21282;
  assign n21284 = pi1156 & ~n21283;
  assign n21285 = ~n21280 & ~n21284;
  assign n21286 = pi792 & ~n21285;
  assign n21287 = ~pi792 & ~n21274;
  assign n21288 = ~n21286 & ~n21287;
  assign n21289 = n59240 & ~n21227;
  assign n21290 = ~n59240 & n21274;
  assign n21291 = ~n21289 & ~n21290;
  assign n21292 = ~n21275 & ~n21276;
  assign n21293 = ~n9743 & ~n59752;
  assign n21294 = n9743 & n21227;
  assign n21295 = ~pi647 & ~n59752;
  assign n21296 = pi647 & n21227;
  assign n21297 = ~n21295 & ~n21296;
  assign n21298 = ~pi1157 & ~n21297;
  assign n21299 = pi647 & ~n59752;
  assign n21300 = ~pi647 & n21227;
  assign n21301 = ~n21299 & ~n21300;
  assign n21302 = pi1157 & ~n21301;
  assign n21303 = ~n21298 & ~n21302;
  assign n21304 = pi787 & ~n21303;
  assign n21305 = ~pi787 & ~n59752;
  assign n21306 = ~n21304 & ~n21305;
  assign n21307 = ~n21293 & ~n21294;
  assign n21308 = ~pi644 & ~n59753;
  assign n21309 = pi715 & ~n21308;
  assign n21310 = ~pi763 & n6654;
  assign n21311 = pi190 & n6853;
  assign n21312 = ~n21310 & ~n21311;
  assign n21313 = pi39 & ~n21312;
  assign n21314 = ~pi190 & pi763;
  assign n21315 = n59164 & n21314;
  assign n21316 = ~pi763 & n8180;
  assign n21317 = pi763 & ~n6799;
  assign n21318 = pi190 & ~n21317;
  assign n21319 = ~n21316 & ~n21318;
  assign n21320 = ~n21315 & n21319;
  assign n21321 = ~n21313 & n21320;
  assign n21322 = ~pi38 & ~n21321;
  assign n21323 = pi763 & n6865;
  assign n21324 = pi38 & ~n21234;
  assign n21325 = ~n21323 & n21324;
  assign n21326 = ~n21322 & ~n21325;
  assign n21327 = n59132 & ~n21326;
  assign n21328 = ~n21229 & ~n21327;
  assign n21329 = ~n7597 & ~n21328;
  assign n21330 = n7597 & ~n21227;
  assign n21331 = ~n21329 & ~n21330;
  assign n21332 = ~pi785 & ~n21331;
  assign n21333 = ~n7598 & ~n21227;
  assign n21334 = pi609 & n21329;
  assign n21335 = ~n21333 & ~n21334;
  assign n21336 = pi1155 & ~n21335;
  assign n21337 = ~n7610 & ~n21227;
  assign n21338 = ~pi609 & n21329;
  assign n21339 = ~n21337 & ~n21338;
  assign n21340 = ~pi1155 & ~n21339;
  assign n21341 = ~n21336 & ~n21340;
  assign n21342 = pi785 & ~n21341;
  assign n21343 = ~n21332 & ~n21342;
  assign n21344 = ~pi781 & ~n21343;
  assign n21345 = pi618 & n21343;
  assign n21346 = ~pi618 & n21227;
  assign n21347 = pi1154 & ~n21346;
  assign n21348 = ~n21345 & n21347;
  assign n21349 = ~pi618 & n21343;
  assign n21350 = pi618 & n21227;
  assign n21351 = ~pi1154 & ~n21350;
  assign n21352 = ~n21349 & n21351;
  assign n21353 = ~n21348 & ~n21352;
  assign n21354 = pi781 & ~n21353;
  assign n21355 = ~n21344 & ~n21354;
  assign n21356 = ~pi789 & ~n21355;
  assign n21357 = pi619 & n21355;
  assign n21358 = ~pi619 & n21227;
  assign n21359 = pi1159 & ~n21358;
  assign n21360 = ~n21357 & n21359;
  assign n21361 = ~pi619 & n21355;
  assign n21362 = pi619 & n21227;
  assign n21363 = ~pi1159 & ~n21362;
  assign n21364 = ~n21361 & n21363;
  assign n21365 = ~n21360 & ~n21364;
  assign n21366 = pi789 & ~n21365;
  assign n21367 = ~n21356 & ~n21366;
  assign n21368 = ~n8054 & n21367;
  assign n21369 = n8054 & n21227;
  assign n21370 = ~n21368 & ~n21369;
  assign n21371 = ~n7793 & ~n21370;
  assign n21372 = n7793 & n21227;
  assign n21373 = ~n21371 & ~n21372;
  assign n21374 = ~n7835 & ~n21373;
  assign n21375 = n7835 & n21227;
  assign n21376 = n7835 & ~n21227;
  assign n21377 = ~n7835 & n21373;
  assign n21378 = ~n21376 & ~n21377;
  assign n21379 = ~n21374 & ~n21375;
  assign n21380 = pi644 & n59754;
  assign n21381 = ~pi644 & n21227;
  assign n21382 = ~pi715 & ~n21381;
  assign n21383 = ~n21380 & n21382;
  assign n21384 = pi1160 & ~n21383;
  assign n21385 = ~n21309 & n21384;
  assign n21386 = pi644 & ~n59753;
  assign n21387 = ~pi715 & ~n21386;
  assign n21388 = ~pi644 & n59754;
  assign n21389 = pi644 & n21227;
  assign n21390 = pi715 & ~n21389;
  assign n21391 = ~n21388 & n21390;
  assign n21392 = ~pi1160 & ~n21391;
  assign n21393 = ~n21387 & n21392;
  assign n21394 = ~n21385 & ~n21393;
  assign n21395 = pi790 & ~n21394;
  assign n21396 = ~pi644 & n21392;
  assign n21397 = pi644 & n21384;
  assign n21398 = pi790 & ~n21397;
  assign n21399 = pi790 & ~n21396;
  assign n21400 = ~n21397 & n21399;
  assign n21401 = ~n21396 & n21398;
  assign n21402 = ~n7872 & n21373;
  assign n21403 = n7832 & ~n21300;
  assign n21404 = n7832 & n21301;
  assign n21405 = ~n21299 & n21403;
  assign n21406 = n7833 & ~n21296;
  assign n21407 = n7833 & n21297;
  assign n21408 = ~n21295 & n21406;
  assign n21409 = ~n59756 & ~n59757;
  assign n21410 = ~n21402 & ~n59757;
  assign n21411 = ~n59756 & n21410;
  assign n21412 = ~n21402 & n21409;
  assign n21413 = pi787 & ~n59758;
  assign n21414 = ~n11154 & n21370;
  assign n21415 = n7791 & ~n21278;
  assign n21416 = n7791 & n21279;
  assign n21417 = ~n21277 & n21415;
  assign n21418 = n7790 & ~n21282;
  assign n21419 = n7790 & n21283;
  assign n21420 = ~n21281 & n21418;
  assign n21421 = ~n59759 & ~n59760;
  assign n21422 = ~n21414 & n21421;
  assign n21423 = pi792 & ~n21422;
  assign n21424 = ~pi699 & n21326;
  assign n21425 = ~pi190 & n59177;
  assign n21426 = pi190 & n7111;
  assign n21427 = ~pi763 & ~n21426;
  assign n21428 = ~n21425 & n21427;
  assign n21429 = pi190 & n7188;
  assign n21430 = ~pi190 & ~n59203;
  assign n21431 = pi763 & ~n21430;
  assign n21432 = ~n21429 & n21431;
  assign n21433 = pi39 & ~n21432;
  assign n21434 = ~n21428 & n21433;
  assign n21435 = ~pi190 & n7310;
  assign n21436 = pi190 & n7333;
  assign n21437 = ~pi763 & ~n21436;
  assign n21438 = ~pi763 & ~n21435;
  assign n21439 = ~n21436 & n21438;
  assign n21440 = ~n21435 & n21437;
  assign n21441 = ~pi190 & ~n7339;
  assign n21442 = pi190 & ~n7347;
  assign n21443 = pi763 & ~n21442;
  assign n21444 = ~n21441 & n21443;
  assign n21445 = ~pi39 & ~n21444;
  assign n21446 = ~n59761 & n21445;
  assign n21447 = ~pi38 & ~n21446;
  assign n21448 = ~pi190 & n8213;
  assign n21449 = pi190 & n8217;
  assign n21450 = ~pi763 & ~n21449;
  assign n21451 = ~n21448 & n21450;
  assign n21452 = pi190 & n9808;
  assign n21453 = ~pi190 & ~n13062;
  assign n21454 = pi763 & ~n21453;
  assign n21455 = ~n21452 & n21454;
  assign n21456 = ~n21451 & ~n21455;
  assign n21457 = ~pi38 & ~n21456;
  assign n21458 = ~n21434 & n21447;
  assign n21459 = ~pi763 & n13069;
  assign n21460 = ~n7222 & ~n21459;
  assign n21461 = ~pi39 & ~n21460;
  assign n21462 = ~pi190 & ~n21461;
  assign n21463 = ~n7056 & ~n21020;
  assign n21464 = pi190 & ~n21463;
  assign n21465 = n59171 & n21464;
  assign n21466 = pi38 & ~n21465;
  assign n21467 = ~n21462 & n21466;
  assign n21468 = pi699 & ~n21467;
  assign n21469 = ~n59762 & n21468;
  assign n21470 = n59132 & ~n21469;
  assign n21471 = n59132 & ~n21424;
  assign n21472 = ~n21469 & n21471;
  assign n21473 = ~n21424 & n21470;
  assign n21474 = ~n21229 & ~n59763;
  assign n21475 = ~pi625 & n21474;
  assign n21476 = pi625 & n21328;
  assign n21477 = ~pi1153 & ~n21476;
  assign n21478 = ~n21475 & n21477;
  assign n21479 = ~pi608 & ~n21247;
  assign n21480 = ~n21478 & n21479;
  assign n21481 = pi625 & n21474;
  assign n21482 = ~pi625 & n21328;
  assign n21483 = pi1153 & ~n21482;
  assign n21484 = ~n21481 & n21483;
  assign n21485 = pi608 & ~n21251;
  assign n21486 = ~n21484 & n21485;
  assign n21487 = ~n21480 & ~n21486;
  assign n21488 = pi778 & ~n21487;
  assign n21489 = ~pi778 & n21474;
  assign n21490 = ~n21488 & ~n21489;
  assign n21491 = ~pi609 & ~n21490;
  assign n21492 = pi609 & n21254;
  assign n21493 = ~pi1155 & ~n21492;
  assign n21494 = ~n21491 & n21493;
  assign n21495 = ~pi660 & ~n21336;
  assign n21496 = ~n21494 & n21495;
  assign n21497 = pi609 & ~n21490;
  assign n21498 = ~pi609 & n21254;
  assign n21499 = pi1155 & ~n21498;
  assign n21500 = ~n21497 & n21499;
  assign n21501 = pi660 & ~n21340;
  assign n21502 = ~n21500 & n21501;
  assign n21503 = ~n21496 & ~n21502;
  assign n21504 = pi785 & ~n21503;
  assign n21505 = ~pi785 & ~n21490;
  assign n21506 = ~n21504 & ~n21505;
  assign n21507 = ~pi618 & ~n21506;
  assign n21508 = pi618 & n59749;
  assign n21509 = ~pi1154 & ~n21508;
  assign n21510 = ~n21507 & n21509;
  assign n21511 = ~pi627 & ~n21348;
  assign n21512 = ~n21510 & n21511;
  assign n21513 = pi618 & ~n21506;
  assign n21514 = ~pi618 & n59749;
  assign n21515 = pi1154 & ~n21514;
  assign n21516 = ~n21513 & n21515;
  assign n21517 = pi627 & ~n21352;
  assign n21518 = ~n21516 & n21517;
  assign n21519 = ~n21512 & ~n21518;
  assign n21520 = pi781 & ~n21519;
  assign n21521 = ~pi781 & ~n21506;
  assign n21522 = ~n21520 & ~n21521;
  assign n21523 = pi619 & ~n21522;
  assign n21524 = ~pi619 & ~n59750;
  assign n21525 = pi1159 & ~n21524;
  assign n21526 = ~n21523 & n21525;
  assign n21527 = pi648 & ~n21364;
  assign n21528 = ~n21526 & n21527;
  assign n21529 = ~pi619 & ~n21522;
  assign n21530 = pi619 & ~n59750;
  assign n21531 = ~pi1159 & ~n21530;
  assign n21532 = ~n21529 & n21531;
  assign n21533 = ~pi648 & ~n21360;
  assign n21534 = ~n21532 & n21533;
  assign n21535 = pi789 & ~n21534;
  assign n21536 = pi789 & ~n21528;
  assign n21537 = ~n21534 & n21536;
  assign n21538 = ~n21528 & n21535;
  assign n21539 = ~pi789 & n21522;
  assign n21540 = n59242 & ~n21539;
  assign n21541 = ~n59764 & n21540;
  assign n21542 = ~pi626 & ~n21367;
  assign n21543 = pi626 & ~n21227;
  assign n21544 = n7760 & ~n21543;
  assign n21545 = ~n21542 & n21544;
  assign n21546 = n7984 & n59751;
  assign n21547 = pi626 & ~n21367;
  assign n21548 = ~pi626 & ~n21227;
  assign n21549 = n7759 & ~n21548;
  assign n21550 = ~n21547 & n21549;
  assign n21551 = ~n21546 & ~n21550;
  assign n21552 = ~n21545 & ~n21546;
  assign n21553 = ~n21550 & n21552;
  assign n21554 = ~n21545 & n21551;
  assign n21555 = pi788 & ~n59765;
  assign n21556 = ~n59357 & ~n21555;
  assign n21557 = ~n21541 & n21556;
  assign n21558 = ~n21423 & ~n21557;
  assign n21559 = ~n8108 & ~n21558;
  assign n21560 = ~n21413 & ~n21559;
  assign n21561 = ~n59755 & n21560;
  assign n21562 = ~n21395 & ~n21561;
  assign n21563 = n58992 & ~n21562;
  assign n21564 = ~pi190 & ~n58992;
  assign n21565 = ~pi832 & ~n21564;
  assign n21566 = ~n21563 & n21565;
  assign po347 = ~n21226 & ~n21566;
  assign n21568 = ~pi191 & ~n2794;
  assign n21569 = pi746 & n6822;
  assign n21570 = ~n21568 & ~n21569;
  assign n21571 = ~n7875 & ~n21570;
  assign n21572 = ~pi785 & ~n21571;
  assign n21573 = n7610 & n21569;
  assign n21574 = n21571 & ~n21573;
  assign n21575 = pi1155 & ~n21574;
  assign n21576 = ~pi1155 & ~n21568;
  assign n21577 = ~n21573 & n21576;
  assign n21578 = ~n21575 & ~n21577;
  assign n21579 = pi785 & ~n21578;
  assign n21580 = ~n21572 & ~n21579;
  assign n21581 = ~pi781 & ~n21580;
  assign n21582 = ~n7890 & n21580;
  assign n21583 = pi1154 & ~n21582;
  assign n21584 = ~n7893 & n21580;
  assign n21585 = ~pi1154 & ~n21584;
  assign n21586 = ~n21583 & ~n21585;
  assign n21587 = pi781 & ~n21586;
  assign n21588 = ~n21581 & ~n21587;
  assign n21589 = ~pi789 & ~n21588;
  assign n21590 = ~n11882 & n21588;
  assign n21591 = pi1159 & ~n21590;
  assign n21592 = ~n11885 & n21588;
  assign n21593 = ~pi1159 & ~n21592;
  assign n21594 = ~n21591 & ~n21593;
  assign n21595 = pi789 & ~n21594;
  assign n21596 = ~n21589 & ~n21595;
  assign n21597 = ~n8054 & ~n21596;
  assign n21598 = n8054 & ~n21568;
  assign n21599 = ~n8054 & n21596;
  assign n21600 = n8054 & n21568;
  assign n21601 = ~n21599 & ~n21600;
  assign n21602 = ~n21597 & ~n21598;
  assign n21603 = ~n7793 & ~n59766;
  assign n21604 = n7793 & n21568;
  assign n21605 = ~n7872 & ~n21604;
  assign n21606 = ~n21603 & ~n21604;
  assign n21607 = ~n7872 & n21606;
  assign n21608 = ~n21603 & n21605;
  assign n21609 = pi729 & n7055;
  assign n21610 = ~n21568 & ~n21609;
  assign n21611 = ~pi778 & ~n21610;
  assign n21612 = ~pi625 & n21609;
  assign n21613 = ~n21610 & ~n21612;
  assign n21614 = pi1153 & ~n21613;
  assign n21615 = ~pi1153 & ~n21568;
  assign n21616 = ~n21612 & n21615;
  assign n21617 = pi778 & ~n21616;
  assign n21618 = ~n21614 & n21617;
  assign n21619 = ~n21611 & ~n21618;
  assign n21620 = ~n7949 & ~n21619;
  assign n21621 = ~n7951 & n21620;
  assign n21622 = ~n7953 & n21621;
  assign n21623 = ~n7955 & n21622;
  assign n21624 = ~n7967 & n21623;
  assign n21625 = pi647 & ~n21624;
  assign n21626 = ~pi647 & ~n21568;
  assign n21627 = ~n21625 & ~n21626;
  assign n21628 = n7832 & ~n21627;
  assign n21629 = ~pi647 & n21624;
  assign n21630 = pi647 & n21568;
  assign n21631 = ~pi1157 & ~n21630;
  assign n21632 = ~n21629 & n21631;
  assign n21633 = pi630 & n21632;
  assign n21634 = ~n21628 & ~n21633;
  assign n21635 = ~n59767 & n21634;
  assign n21636 = pi787 & ~n21635;
  assign n21637 = ~pi626 & ~n21596;
  assign n21638 = pi626 & ~n21568;
  assign n21639 = n7760 & ~n21638;
  assign n21640 = ~n21637 & n21639;
  assign n21641 = n7984 & n21622;
  assign n21642 = pi626 & ~n21596;
  assign n21643 = ~pi626 & ~n21568;
  assign n21644 = n7759 & ~n21643;
  assign n21645 = ~n21642 & n21644;
  assign n21646 = ~n21641 & ~n21645;
  assign n21647 = ~n21640 & ~n21641;
  assign n21648 = ~n21645 & n21647;
  assign n21649 = ~n21640 & n21646;
  assign n21650 = pi788 & ~n59768;
  assign n21651 = ~n6701 & ~n21610;
  assign n21652 = pi625 & n21651;
  assign n21653 = n21570 & ~n21651;
  assign n21654 = ~n21652 & ~n21653;
  assign n21655 = n21615 & ~n21654;
  assign n21656 = ~pi608 & ~n21614;
  assign n21657 = ~n21655 & n21656;
  assign n21658 = pi1153 & n21570;
  assign n21659 = ~n21652 & n21658;
  assign n21660 = pi608 & ~n21616;
  assign n21661 = ~n21659 & n21660;
  assign n21662 = ~n21657 & ~n21661;
  assign n21663 = pi778 & ~n21662;
  assign n21664 = ~pi778 & ~n21653;
  assign n21665 = ~n21663 & ~n21664;
  assign n21666 = ~pi609 & ~n21665;
  assign n21667 = pi609 & ~n21619;
  assign n21668 = ~pi1155 & ~n21667;
  assign n21669 = ~n21666 & n21668;
  assign n21670 = ~pi660 & ~n21575;
  assign n21671 = ~n21669 & n21670;
  assign n21672 = pi609 & ~n21665;
  assign n21673 = ~pi609 & ~n21619;
  assign n21674 = pi1155 & ~n21673;
  assign n21675 = ~n21672 & n21674;
  assign n21676 = pi660 & ~n21577;
  assign n21677 = ~n21675 & n21676;
  assign n21678 = ~n21671 & ~n21677;
  assign n21679 = pi785 & ~n21678;
  assign n21680 = ~pi785 & ~n21665;
  assign n21681 = ~n21679 & ~n21680;
  assign n21682 = ~pi618 & ~n21681;
  assign n21683 = pi618 & n21620;
  assign n21684 = ~pi1154 & ~n21683;
  assign n21685 = ~n21682 & n21684;
  assign n21686 = ~pi627 & ~n21583;
  assign n21687 = ~n21685 & n21686;
  assign n21688 = pi618 & ~n21681;
  assign n21689 = ~pi618 & n21620;
  assign n21690 = pi1154 & ~n21689;
  assign n21691 = ~n21688 & n21690;
  assign n21692 = pi627 & ~n21585;
  assign n21693 = ~n21691 & n21692;
  assign n21694 = ~n21687 & ~n21693;
  assign n21695 = pi781 & ~n21694;
  assign n21696 = ~pi781 & ~n21681;
  assign n21697 = ~n21695 & ~n21696;
  assign n21698 = pi619 & ~n21697;
  assign n21699 = ~pi619 & n21621;
  assign n21700 = pi1159 & ~n21699;
  assign n21701 = ~n21698 & n21700;
  assign n21702 = pi648 & ~n21593;
  assign n21703 = ~n21701 & n21702;
  assign n21704 = ~pi619 & ~n21697;
  assign n21705 = pi619 & n21621;
  assign n21706 = ~pi1159 & ~n21705;
  assign n21707 = ~n21704 & n21706;
  assign n21708 = ~pi648 & ~n21591;
  assign n21709 = ~n21707 & n21708;
  assign n21710 = pi789 & ~n21709;
  assign n21711 = pi789 & ~n21703;
  assign n21712 = ~n21709 & n21711;
  assign n21713 = ~n21703 & n21710;
  assign n21714 = ~pi789 & n21697;
  assign n21715 = n59242 & ~n21714;
  assign n21716 = ~n59769 & n21715;
  assign n21717 = ~n21650 & ~n21716;
  assign n21718 = ~n59357 & ~n21717;
  assign n21719 = n7957 & ~n59766;
  assign n21720 = n8065 & n21623;
  assign n21721 = pi629 & ~n21720;
  assign n21722 = ~n21719 & n21721;
  assign n21723 = n7958 & ~n59766;
  assign n21724 = n8074 & n21623;
  assign n21725 = ~pi629 & ~n21724;
  assign n21726 = ~n21723 & n21725;
  assign n21727 = pi792 & ~n21726;
  assign n21728 = ~n21723 & ~n21724;
  assign n21729 = ~pi629 & ~n21728;
  assign n21730 = ~n21719 & ~n21720;
  assign n21731 = pi629 & ~n21730;
  assign n21732 = ~n21729 & ~n21731;
  assign n21733 = pi792 & ~n21732;
  assign n21734 = pi792 & ~n21722;
  assign n21735 = ~n21726 & n21734;
  assign n21736 = ~n21722 & n21727;
  assign n21737 = ~n8108 & ~n59770;
  assign n21738 = ~n21718 & n21737;
  assign n21739 = ~n21636 & ~n21738;
  assign n21740 = pi644 & n21739;
  assign n21741 = ~pi787 & ~n21624;
  assign n21742 = pi1157 & ~n21627;
  assign n21743 = ~n21632 & ~n21742;
  assign n21744 = pi787 & ~n21743;
  assign n21745 = ~n21741 & ~n21744;
  assign n21746 = ~pi644 & n21745;
  assign n21747 = pi715 & ~n21746;
  assign n21748 = ~n21740 & n21747;
  assign n21749 = ~n11491 & n21568;
  assign n21750 = ~n7835 & n21603;
  assign n21751 = ~n7835 & ~n21606;
  assign n21752 = n7835 & n21568;
  assign n21753 = ~n21751 & ~n21752;
  assign n21754 = ~n21749 & ~n21750;
  assign n21755 = pi644 & ~n59771;
  assign n21756 = ~pi644 & n21568;
  assign n21757 = ~pi715 & ~n21756;
  assign n21758 = ~n21755 & n21757;
  assign n21759 = pi1160 & ~n21758;
  assign n21760 = ~n21748 & n21759;
  assign n21761 = ~pi644 & n21739;
  assign n21762 = pi644 & n21745;
  assign n21763 = ~pi715 & ~n21762;
  assign n21764 = ~n21761 & n21763;
  assign n21765 = ~pi644 & ~n59771;
  assign n21766 = pi644 & n21568;
  assign n21767 = pi715 & ~n21766;
  assign n21768 = ~n21765 & n21767;
  assign n21769 = ~pi1160 & ~n21768;
  assign n21770 = ~n21764 & n21769;
  assign n21771 = ~n21760 & ~n21770;
  assign n21772 = pi790 & ~n21771;
  assign n21773 = ~pi790 & n21739;
  assign n21774 = pi832 & ~n21773;
  assign n21775 = ~n21772 & n21774;
  assign n21776 = ~pi191 & ~n7560;
  assign n21777 = n59231 & ~n21776;
  assign n21778 = pi191 & ~n59132;
  assign n21779 = ~pi191 & n8249;
  assign n21780 = pi191 & n59251;
  assign n21781 = ~pi38 & ~n21780;
  assign n21782 = ~n21779 & n21781;
  assign n21783 = ~pi191 & ~n6863;
  assign n21784 = n7547 & ~n21783;
  assign n21785 = pi729 & ~n21784;
  assign n21786 = ~n21782 & n21785;
  assign n21787 = ~pi191 & ~pi729;
  assign n21788 = ~n7553 & n21787;
  assign n21789 = n59132 & ~n21788;
  assign n21790 = ~n21786 & n21789;
  assign n21791 = ~n21778 & ~n21790;
  assign n21792 = ~pi778 & ~n21791;
  assign n21793 = pi625 & n21791;
  assign n21794 = ~pi625 & n21776;
  assign n21795 = pi1153 & ~n21794;
  assign n21796 = ~n21793 & n21795;
  assign n21797 = ~pi625 & n21791;
  assign n21798 = pi625 & n21776;
  assign n21799 = ~pi1153 & ~n21798;
  assign n21800 = ~n21797 & n21799;
  assign n21801 = ~n21796 & ~n21800;
  assign n21802 = pi778 & ~n21801;
  assign n21803 = ~n21792 & ~n21802;
  assign n21804 = ~n59229 & n21803;
  assign n21805 = n59229 & n21776;
  assign n21806 = n59229 & ~n21776;
  assign n21807 = ~n59229 & ~n21803;
  assign n21808 = ~n21806 & ~n21807;
  assign n21809 = ~n21804 & ~n21805;
  assign n21810 = ~n59231 & ~n59772;
  assign n21811 = ~n59231 & n59772;
  assign n21812 = n59231 & n21776;
  assign n21813 = ~n21811 & ~n21812;
  assign n21814 = ~n21777 & ~n21810;
  assign n21815 = ~n7716 & ~n59773;
  assign n21816 = n7716 & n21776;
  assign n21817 = n7716 & ~n21776;
  assign n21818 = ~n7716 & n59773;
  assign n21819 = ~n21817 & ~n21818;
  assign n21820 = ~n21815 & ~n21816;
  assign n21821 = ~n7762 & n59774;
  assign n21822 = n7762 & n21776;
  assign n21823 = ~n21821 & ~n21822;
  assign n21824 = ~n59240 & ~n21823;
  assign n21825 = n59240 & n21776;
  assign n21826 = ~pi628 & ~n21823;
  assign n21827 = pi628 & n21776;
  assign n21828 = ~n21826 & ~n21827;
  assign n21829 = ~pi1156 & ~n21828;
  assign n21830 = pi628 & ~n21823;
  assign n21831 = ~pi628 & n21776;
  assign n21832 = ~n21830 & ~n21831;
  assign n21833 = pi1156 & ~n21832;
  assign n21834 = ~n21829 & ~n21833;
  assign n21835 = pi792 & ~n21834;
  assign n21836 = ~pi792 & ~n21823;
  assign n21837 = ~n21835 & ~n21836;
  assign n21838 = n59240 & ~n21776;
  assign n21839 = ~n59240 & n21823;
  assign n21840 = ~n21838 & ~n21839;
  assign n21841 = ~n21824 & ~n21825;
  assign n21842 = ~n9743 & ~n59775;
  assign n21843 = n9743 & n21776;
  assign n21844 = ~pi647 & ~n59775;
  assign n21845 = pi647 & n21776;
  assign n21846 = ~n21844 & ~n21845;
  assign n21847 = ~pi1157 & ~n21846;
  assign n21848 = pi647 & ~n59775;
  assign n21849 = ~pi647 & n21776;
  assign n21850 = ~n21848 & ~n21849;
  assign n21851 = pi1157 & ~n21850;
  assign n21852 = ~n21847 & ~n21851;
  assign n21853 = pi787 & ~n21852;
  assign n21854 = ~pi787 & ~n59775;
  assign n21855 = ~n21853 & ~n21854;
  assign n21856 = ~n21842 & ~n21843;
  assign n21857 = ~pi644 & ~n59776;
  assign n21858 = pi715 & ~n21857;
  assign n21859 = ~pi746 & n6654;
  assign n21860 = pi191 & n6853;
  assign n21861 = ~n21859 & ~n21860;
  assign n21862 = pi39 & ~n21861;
  assign n21863 = ~pi191 & pi746;
  assign n21864 = n59164 & n21863;
  assign n21865 = ~pi746 & n8180;
  assign n21866 = pi746 & ~n6799;
  assign n21867 = pi191 & ~n21866;
  assign n21868 = ~n21865 & ~n21867;
  assign n21869 = ~n21864 & n21868;
  assign n21870 = ~n21862 & n21869;
  assign n21871 = ~pi38 & ~n21870;
  assign n21872 = pi746 & n6865;
  assign n21873 = pi38 & ~n21783;
  assign n21874 = ~n21872 & n21873;
  assign n21875 = ~n21871 & ~n21874;
  assign n21876 = n59132 & ~n21875;
  assign n21877 = ~n21778 & ~n21876;
  assign n21878 = ~n7597 & ~n21877;
  assign n21879 = n7597 & ~n21776;
  assign n21880 = ~n21878 & ~n21879;
  assign n21881 = ~pi785 & ~n21880;
  assign n21882 = ~n7598 & ~n21776;
  assign n21883 = pi609 & n21878;
  assign n21884 = ~n21882 & ~n21883;
  assign n21885 = pi1155 & ~n21884;
  assign n21886 = ~n7610 & ~n21776;
  assign n21887 = ~pi609 & n21878;
  assign n21888 = ~n21886 & ~n21887;
  assign n21889 = ~pi1155 & ~n21888;
  assign n21890 = ~n21885 & ~n21889;
  assign n21891 = pi785 & ~n21890;
  assign n21892 = ~n21881 & ~n21891;
  assign n21893 = ~pi781 & ~n21892;
  assign n21894 = pi618 & n21892;
  assign n21895 = ~pi618 & n21776;
  assign n21896 = pi1154 & ~n21895;
  assign n21897 = ~n21894 & n21896;
  assign n21898 = ~pi618 & n21892;
  assign n21899 = pi618 & n21776;
  assign n21900 = ~pi1154 & ~n21899;
  assign n21901 = ~n21898 & n21900;
  assign n21902 = ~n21897 & ~n21901;
  assign n21903 = pi781 & ~n21902;
  assign n21904 = ~n21893 & ~n21903;
  assign n21905 = ~pi789 & ~n21904;
  assign n21906 = pi619 & n21904;
  assign n21907 = ~pi619 & n21776;
  assign n21908 = pi1159 & ~n21907;
  assign n21909 = ~n21906 & n21908;
  assign n21910 = ~pi619 & n21904;
  assign n21911 = pi619 & n21776;
  assign n21912 = ~pi1159 & ~n21911;
  assign n21913 = ~n21910 & n21912;
  assign n21914 = ~n21909 & ~n21913;
  assign n21915 = pi789 & ~n21914;
  assign n21916 = ~n21905 & ~n21915;
  assign n21917 = ~n8054 & n21916;
  assign n21918 = n8054 & n21776;
  assign n21919 = ~n21917 & ~n21918;
  assign n21920 = ~n7793 & ~n21919;
  assign n21921 = n7793 & n21776;
  assign n21922 = ~n21920 & ~n21921;
  assign n21923 = ~n7835 & ~n21922;
  assign n21924 = n7835 & n21776;
  assign n21925 = n7835 & ~n21776;
  assign n21926 = ~n7835 & n21922;
  assign n21927 = ~n21925 & ~n21926;
  assign n21928 = ~n21923 & ~n21924;
  assign n21929 = pi644 & n59777;
  assign n21930 = ~pi644 & n21776;
  assign n21931 = ~pi715 & ~n21930;
  assign n21932 = ~n21929 & n21931;
  assign n21933 = pi1160 & ~n21932;
  assign n21934 = ~n21858 & n21933;
  assign n21935 = pi644 & ~n59776;
  assign n21936 = ~pi715 & ~n21935;
  assign n21937 = ~pi644 & n59777;
  assign n21938 = pi644 & n21776;
  assign n21939 = pi715 & ~n21938;
  assign n21940 = ~n21937 & n21939;
  assign n21941 = ~pi1160 & ~n21940;
  assign n21942 = ~n21936 & n21941;
  assign n21943 = ~n21934 & ~n21942;
  assign n21944 = pi790 & ~n21943;
  assign n21945 = ~pi644 & n21941;
  assign n21946 = pi644 & n21933;
  assign n21947 = pi790 & ~n21946;
  assign n21948 = pi790 & ~n21945;
  assign n21949 = ~n21946 & n21948;
  assign n21950 = ~n21945 & n21947;
  assign n21951 = ~n7872 & n21922;
  assign n21952 = n7832 & ~n21849;
  assign n21953 = n7832 & n21850;
  assign n21954 = ~n21848 & n21952;
  assign n21955 = n7833 & ~n21845;
  assign n21956 = n7833 & n21846;
  assign n21957 = ~n21844 & n21955;
  assign n21958 = ~n59779 & ~n59780;
  assign n21959 = ~n21951 & ~n59780;
  assign n21960 = ~n59779 & n21959;
  assign n21961 = ~n21951 & n21958;
  assign n21962 = pi787 & ~n59781;
  assign n21963 = ~n11154 & n21919;
  assign n21964 = n7791 & ~n21827;
  assign n21965 = n7791 & n21828;
  assign n21966 = ~n21826 & n21964;
  assign n21967 = n7790 & ~n21831;
  assign n21968 = n7790 & n21832;
  assign n21969 = ~n21830 & n21967;
  assign n21970 = ~n59782 & ~n59783;
  assign n21971 = ~n21963 & n21970;
  assign n21972 = pi792 & ~n21971;
  assign n21973 = ~pi729 & n21875;
  assign n21974 = ~pi191 & n59177;
  assign n21975 = pi191 & n7111;
  assign n21976 = ~pi746 & ~n21975;
  assign n21977 = ~n21974 & n21976;
  assign n21978 = pi191 & n7188;
  assign n21979 = ~pi191 & ~n59203;
  assign n21980 = pi746 & ~n21979;
  assign n21981 = ~n21978 & n21980;
  assign n21982 = pi39 & ~n21981;
  assign n21983 = ~n21977 & n21982;
  assign n21984 = ~pi191 & n7310;
  assign n21985 = pi191 & n7333;
  assign n21986 = ~pi746 & ~n21985;
  assign n21987 = ~pi746 & ~n21984;
  assign n21988 = ~n21985 & n21987;
  assign n21989 = ~n21984 & n21986;
  assign n21990 = ~pi191 & ~n7339;
  assign n21991 = pi191 & ~n7347;
  assign n21992 = pi746 & ~n21991;
  assign n21993 = ~n21990 & n21992;
  assign n21994 = ~pi39 & ~n21993;
  assign n21995 = ~n59784 & n21994;
  assign n21996 = ~pi38 & ~n21995;
  assign n21997 = ~pi191 & n8213;
  assign n21998 = pi191 & n8217;
  assign n21999 = ~pi746 & ~n21998;
  assign n22000 = ~n21997 & n21999;
  assign n22001 = pi191 & n9808;
  assign n22002 = ~pi191 & ~n13062;
  assign n22003 = pi746 & ~n22002;
  assign n22004 = ~n22001 & n22003;
  assign n22005 = ~n22000 & ~n22004;
  assign n22006 = ~pi38 & ~n22005;
  assign n22007 = ~n21983 & n21996;
  assign n22008 = ~pi746 & n13069;
  assign n22009 = ~n7222 & ~n22008;
  assign n22010 = ~pi39 & ~n22009;
  assign n22011 = ~pi191 & ~n22010;
  assign n22012 = ~n7056 & ~n21569;
  assign n22013 = pi191 & ~n22012;
  assign n22014 = n59171 & n22013;
  assign n22015 = pi38 & ~n22014;
  assign n22016 = ~n22011 & n22015;
  assign n22017 = pi729 & ~n22016;
  assign n22018 = ~n59785 & n22017;
  assign n22019 = n59132 & ~n22018;
  assign n22020 = n59132 & ~n21973;
  assign n22021 = ~n22018 & n22020;
  assign n22022 = ~n21973 & n22019;
  assign n22023 = ~n21778 & ~n59786;
  assign n22024 = ~pi625 & n22023;
  assign n22025 = pi625 & n21877;
  assign n22026 = ~pi1153 & ~n22025;
  assign n22027 = ~n22024 & n22026;
  assign n22028 = ~pi608 & ~n21796;
  assign n22029 = ~n22027 & n22028;
  assign n22030 = pi625 & n22023;
  assign n22031 = ~pi625 & n21877;
  assign n22032 = pi1153 & ~n22031;
  assign n22033 = ~n22030 & n22032;
  assign n22034 = pi608 & ~n21800;
  assign n22035 = ~n22033 & n22034;
  assign n22036 = ~n22029 & ~n22035;
  assign n22037 = pi778 & ~n22036;
  assign n22038 = ~pi778 & n22023;
  assign n22039 = ~n22037 & ~n22038;
  assign n22040 = ~pi609 & ~n22039;
  assign n22041 = pi609 & n21803;
  assign n22042 = ~pi1155 & ~n22041;
  assign n22043 = ~n22040 & n22042;
  assign n22044 = ~pi660 & ~n21885;
  assign n22045 = ~n22043 & n22044;
  assign n22046 = pi609 & ~n22039;
  assign n22047 = ~pi609 & n21803;
  assign n22048 = pi1155 & ~n22047;
  assign n22049 = ~n22046 & n22048;
  assign n22050 = pi660 & ~n21889;
  assign n22051 = ~n22049 & n22050;
  assign n22052 = ~n22045 & ~n22051;
  assign n22053 = pi785 & ~n22052;
  assign n22054 = ~pi785 & ~n22039;
  assign n22055 = ~n22053 & ~n22054;
  assign n22056 = ~pi618 & ~n22055;
  assign n22057 = pi618 & n59772;
  assign n22058 = ~pi1154 & ~n22057;
  assign n22059 = ~n22056 & n22058;
  assign n22060 = ~pi627 & ~n21897;
  assign n22061 = ~n22059 & n22060;
  assign n22062 = pi618 & ~n22055;
  assign n22063 = ~pi618 & n59772;
  assign n22064 = pi1154 & ~n22063;
  assign n22065 = ~n22062 & n22064;
  assign n22066 = pi627 & ~n21901;
  assign n22067 = ~n22065 & n22066;
  assign n22068 = ~n22061 & ~n22067;
  assign n22069 = pi781 & ~n22068;
  assign n22070 = ~pi781 & ~n22055;
  assign n22071 = ~n22069 & ~n22070;
  assign n22072 = pi619 & ~n22071;
  assign n22073 = ~pi619 & ~n59773;
  assign n22074 = pi1159 & ~n22073;
  assign n22075 = ~n22072 & n22074;
  assign n22076 = pi648 & ~n21913;
  assign n22077 = ~n22075 & n22076;
  assign n22078 = ~pi619 & ~n22071;
  assign n22079 = pi619 & ~n59773;
  assign n22080 = ~pi1159 & ~n22079;
  assign n22081 = ~n22078 & n22080;
  assign n22082 = ~pi648 & ~n21909;
  assign n22083 = ~n22081 & n22082;
  assign n22084 = pi789 & ~n22083;
  assign n22085 = pi789 & ~n22077;
  assign n22086 = ~n22083 & n22085;
  assign n22087 = ~n22077 & n22084;
  assign n22088 = ~pi789 & n22071;
  assign n22089 = n59242 & ~n22088;
  assign n22090 = ~n59787 & n22089;
  assign n22091 = ~pi626 & ~n21916;
  assign n22092 = pi626 & ~n21776;
  assign n22093 = n7760 & ~n22092;
  assign n22094 = ~n22091 & n22093;
  assign n22095 = n7984 & n59774;
  assign n22096 = pi626 & ~n21916;
  assign n22097 = ~pi626 & ~n21776;
  assign n22098 = n7759 & ~n22097;
  assign n22099 = ~n22096 & n22098;
  assign n22100 = ~n22095 & ~n22099;
  assign n22101 = ~n22094 & ~n22095;
  assign n22102 = ~n22099 & n22101;
  assign n22103 = ~n22094 & n22100;
  assign n22104 = pi788 & ~n59788;
  assign n22105 = ~n59357 & ~n22104;
  assign n22106 = ~n22090 & n22105;
  assign n22107 = ~n21972 & ~n22106;
  assign n22108 = ~n8108 & ~n22107;
  assign n22109 = ~n21962 & ~n22108;
  assign n22110 = ~n59778 & n22109;
  assign n22111 = ~n21944 & ~n22110;
  assign n22112 = n58992 & ~n22111;
  assign n22113 = ~pi191 & ~n58992;
  assign n22114 = ~pi832 & ~n22113;
  assign n22115 = ~n22112 & n22114;
  assign po348 = ~n21775 & ~n22115;
  assign n22117 = ~pi192 & ~n2794;
  assign n22118 = pi764 & n6822;
  assign n22119 = ~n22117 & ~n22118;
  assign n22120 = ~n7875 & ~n22119;
  assign n22121 = ~pi785 & ~n22120;
  assign n22122 = n7610 & n22118;
  assign n22123 = n22120 & ~n22122;
  assign n22124 = pi1155 & ~n22123;
  assign n22125 = ~pi1155 & ~n22117;
  assign n22126 = ~n22122 & n22125;
  assign n22127 = ~n22124 & ~n22126;
  assign n22128 = pi785 & ~n22127;
  assign n22129 = ~n22121 & ~n22128;
  assign n22130 = ~pi781 & ~n22129;
  assign n22131 = ~n7890 & n22129;
  assign n22132 = pi1154 & ~n22131;
  assign n22133 = ~n7893 & n22129;
  assign n22134 = ~pi1154 & ~n22133;
  assign n22135 = ~n22132 & ~n22134;
  assign n22136 = pi781 & ~n22135;
  assign n22137 = ~n22130 & ~n22136;
  assign n22138 = ~pi789 & ~n22137;
  assign n22139 = ~n11882 & n22137;
  assign n22140 = pi1159 & ~n22139;
  assign n22141 = ~n11885 & n22137;
  assign n22142 = ~pi1159 & ~n22141;
  assign n22143 = ~n22140 & ~n22142;
  assign n22144 = pi789 & ~n22143;
  assign n22145 = ~n22138 & ~n22144;
  assign n22146 = ~n8054 & ~n22145;
  assign n22147 = n8054 & ~n22117;
  assign n22148 = ~n8054 & n22145;
  assign n22149 = n8054 & n22117;
  assign n22150 = ~n22148 & ~n22149;
  assign n22151 = ~n22146 & ~n22147;
  assign n22152 = ~n7793 & ~n59789;
  assign n22153 = n7793 & n22117;
  assign n22154 = ~n7872 & ~n22153;
  assign n22155 = ~n22152 & ~n22153;
  assign n22156 = ~n7872 & n22155;
  assign n22157 = ~n22152 & n22154;
  assign n22158 = pi691 & n7055;
  assign n22159 = ~n22117 & ~n22158;
  assign n22160 = ~pi778 & ~n22159;
  assign n22161 = ~pi625 & n22158;
  assign n22162 = ~n22159 & ~n22161;
  assign n22163 = pi1153 & ~n22162;
  assign n22164 = ~pi1153 & ~n22117;
  assign n22165 = ~n22161 & n22164;
  assign n22166 = pi778 & ~n22165;
  assign n22167 = ~n22163 & n22166;
  assign n22168 = ~n22160 & ~n22167;
  assign n22169 = ~n7949 & ~n22168;
  assign n22170 = ~n7951 & n22169;
  assign n22171 = ~n7953 & n22170;
  assign n22172 = ~n7955 & n22171;
  assign n22173 = ~n7967 & n22172;
  assign n22174 = pi647 & ~n22173;
  assign n22175 = ~pi647 & ~n22117;
  assign n22176 = ~n22174 & ~n22175;
  assign n22177 = n7832 & ~n22176;
  assign n22178 = ~pi647 & n22173;
  assign n22179 = pi647 & n22117;
  assign n22180 = ~pi1157 & ~n22179;
  assign n22181 = ~n22178 & n22180;
  assign n22182 = pi630 & n22181;
  assign n22183 = ~n22177 & ~n22182;
  assign n22184 = ~n59790 & n22183;
  assign n22185 = pi787 & ~n22184;
  assign n22186 = ~pi626 & ~n22145;
  assign n22187 = pi626 & ~n22117;
  assign n22188 = n7760 & ~n22187;
  assign n22189 = ~n22186 & n22188;
  assign n22190 = n7984 & n22171;
  assign n22191 = pi626 & ~n22145;
  assign n22192 = ~pi626 & ~n22117;
  assign n22193 = n7759 & ~n22192;
  assign n22194 = ~n22191 & n22193;
  assign n22195 = ~n22190 & ~n22194;
  assign n22196 = ~n22189 & ~n22190;
  assign n22197 = ~n22194 & n22196;
  assign n22198 = ~n22189 & n22195;
  assign n22199 = pi788 & ~n59791;
  assign n22200 = ~n6701 & ~n22159;
  assign n22201 = pi625 & n22200;
  assign n22202 = n22119 & ~n22200;
  assign n22203 = ~n22201 & ~n22202;
  assign n22204 = n22164 & ~n22203;
  assign n22205 = ~pi608 & ~n22163;
  assign n22206 = ~n22204 & n22205;
  assign n22207 = pi1153 & n22119;
  assign n22208 = ~n22201 & n22207;
  assign n22209 = pi608 & ~n22165;
  assign n22210 = ~n22208 & n22209;
  assign n22211 = ~n22206 & ~n22210;
  assign n22212 = pi778 & ~n22211;
  assign n22213 = ~pi778 & ~n22202;
  assign n22214 = ~n22212 & ~n22213;
  assign n22215 = ~pi609 & ~n22214;
  assign n22216 = pi609 & ~n22168;
  assign n22217 = ~pi1155 & ~n22216;
  assign n22218 = ~n22215 & n22217;
  assign n22219 = ~pi660 & ~n22124;
  assign n22220 = ~n22218 & n22219;
  assign n22221 = pi609 & ~n22214;
  assign n22222 = ~pi609 & ~n22168;
  assign n22223 = pi1155 & ~n22222;
  assign n22224 = ~n22221 & n22223;
  assign n22225 = pi660 & ~n22126;
  assign n22226 = ~n22224 & n22225;
  assign n22227 = ~n22220 & ~n22226;
  assign n22228 = pi785 & ~n22227;
  assign n22229 = ~pi785 & ~n22214;
  assign n22230 = ~n22228 & ~n22229;
  assign n22231 = ~pi618 & ~n22230;
  assign n22232 = pi618 & n22169;
  assign n22233 = ~pi1154 & ~n22232;
  assign n22234 = ~n22231 & n22233;
  assign n22235 = ~pi627 & ~n22132;
  assign n22236 = ~n22234 & n22235;
  assign n22237 = pi618 & ~n22230;
  assign n22238 = ~pi618 & n22169;
  assign n22239 = pi1154 & ~n22238;
  assign n22240 = ~n22237 & n22239;
  assign n22241 = pi627 & ~n22134;
  assign n22242 = ~n22240 & n22241;
  assign n22243 = ~n22236 & ~n22242;
  assign n22244 = pi781 & ~n22243;
  assign n22245 = ~pi781 & ~n22230;
  assign n22246 = ~n22244 & ~n22245;
  assign n22247 = pi619 & ~n22246;
  assign n22248 = ~pi619 & n22170;
  assign n22249 = pi1159 & ~n22248;
  assign n22250 = ~n22247 & n22249;
  assign n22251 = pi648 & ~n22142;
  assign n22252 = ~n22250 & n22251;
  assign n22253 = ~pi619 & ~n22246;
  assign n22254 = pi619 & n22170;
  assign n22255 = ~pi1159 & ~n22254;
  assign n22256 = ~n22253 & n22255;
  assign n22257 = ~pi648 & ~n22140;
  assign n22258 = ~n22256 & n22257;
  assign n22259 = pi789 & ~n22258;
  assign n22260 = pi789 & ~n22252;
  assign n22261 = ~n22258 & n22260;
  assign n22262 = ~n22252 & n22259;
  assign n22263 = ~pi789 & n22246;
  assign n22264 = n59242 & ~n22263;
  assign n22265 = ~n59792 & n22264;
  assign n22266 = ~n22199 & ~n22265;
  assign n22267 = ~n59357 & ~n22266;
  assign n22268 = n7957 & ~n59789;
  assign n22269 = n8065 & n22172;
  assign n22270 = pi629 & ~n22269;
  assign n22271 = ~n22268 & n22270;
  assign n22272 = n7958 & ~n59789;
  assign n22273 = n8074 & n22172;
  assign n22274 = ~pi629 & ~n22273;
  assign n22275 = ~n22272 & n22274;
  assign n22276 = pi792 & ~n22275;
  assign n22277 = ~n22272 & ~n22273;
  assign n22278 = ~pi629 & ~n22277;
  assign n22279 = ~n22268 & ~n22269;
  assign n22280 = pi629 & ~n22279;
  assign n22281 = ~n22278 & ~n22280;
  assign n22282 = pi792 & ~n22281;
  assign n22283 = pi792 & ~n22271;
  assign n22284 = ~n22275 & n22283;
  assign n22285 = ~n22271 & n22276;
  assign n22286 = ~n8108 & ~n59793;
  assign n22287 = ~n22267 & n22286;
  assign n22288 = ~n22185 & ~n22287;
  assign n22289 = pi644 & n22288;
  assign n22290 = ~pi787 & ~n22173;
  assign n22291 = pi1157 & ~n22176;
  assign n22292 = ~n22181 & ~n22291;
  assign n22293 = pi787 & ~n22292;
  assign n22294 = ~n22290 & ~n22293;
  assign n22295 = ~pi644 & n22294;
  assign n22296 = pi715 & ~n22295;
  assign n22297 = ~n22289 & n22296;
  assign n22298 = ~n11491 & n22117;
  assign n22299 = ~n7835 & n22152;
  assign n22300 = ~n7835 & ~n22155;
  assign n22301 = n7835 & n22117;
  assign n22302 = ~n22300 & ~n22301;
  assign n22303 = ~n22298 & ~n22299;
  assign n22304 = pi644 & ~n59794;
  assign n22305 = ~pi644 & n22117;
  assign n22306 = ~pi715 & ~n22305;
  assign n22307 = ~n22304 & n22306;
  assign n22308 = pi1160 & ~n22307;
  assign n22309 = ~n22297 & n22308;
  assign n22310 = ~pi644 & n22288;
  assign n22311 = pi644 & n22294;
  assign n22312 = ~pi715 & ~n22311;
  assign n22313 = ~n22310 & n22312;
  assign n22314 = ~pi644 & ~n59794;
  assign n22315 = pi644 & n22117;
  assign n22316 = pi715 & ~n22315;
  assign n22317 = ~n22314 & n22316;
  assign n22318 = ~pi1160 & ~n22317;
  assign n22319 = ~n22313 & n22318;
  assign n22320 = ~n22309 & ~n22319;
  assign n22321 = pi790 & ~n22320;
  assign n22322 = ~pi790 & n22288;
  assign n22323 = pi832 & ~n22322;
  assign n22324 = ~n22321 & n22323;
  assign n22325 = ~pi192 & ~n7560;
  assign n22326 = n59231 & ~n22325;
  assign n22327 = pi192 & ~n59132;
  assign n22328 = ~pi192 & n8249;
  assign n22329 = pi192 & n59251;
  assign n22330 = ~pi38 & ~n22329;
  assign n22331 = ~n22328 & n22330;
  assign n22332 = ~pi192 & ~n6863;
  assign n22333 = n7547 & ~n22332;
  assign n22334 = pi691 & ~n22333;
  assign n22335 = ~n22331 & n22334;
  assign n22336 = ~pi192 & ~pi691;
  assign n22337 = ~n7553 & n22336;
  assign n22338 = n59132 & ~n22337;
  assign n22339 = ~n22335 & n22338;
  assign n22340 = ~n22327 & ~n22339;
  assign n22341 = ~pi778 & ~n22340;
  assign n22342 = pi625 & n22340;
  assign n22343 = ~pi625 & n22325;
  assign n22344 = pi1153 & ~n22343;
  assign n22345 = ~n22342 & n22344;
  assign n22346 = ~pi625 & n22340;
  assign n22347 = pi625 & n22325;
  assign n22348 = ~pi1153 & ~n22347;
  assign n22349 = ~n22346 & n22348;
  assign n22350 = ~n22345 & ~n22349;
  assign n22351 = pi778 & ~n22350;
  assign n22352 = ~n22341 & ~n22351;
  assign n22353 = ~n59229 & n22352;
  assign n22354 = n59229 & n22325;
  assign n22355 = n59229 & ~n22325;
  assign n22356 = ~n59229 & ~n22352;
  assign n22357 = ~n22355 & ~n22356;
  assign n22358 = ~n22353 & ~n22354;
  assign n22359 = ~n59231 & ~n59795;
  assign n22360 = ~n59231 & n59795;
  assign n22361 = n59231 & n22325;
  assign n22362 = ~n22360 & ~n22361;
  assign n22363 = ~n22326 & ~n22359;
  assign n22364 = ~n7716 & ~n59796;
  assign n22365 = n7716 & n22325;
  assign n22366 = n7716 & ~n22325;
  assign n22367 = ~n7716 & n59796;
  assign n22368 = ~n22366 & ~n22367;
  assign n22369 = ~n22364 & ~n22365;
  assign n22370 = ~n7762 & n59797;
  assign n22371 = n7762 & n22325;
  assign n22372 = ~n22370 & ~n22371;
  assign n22373 = ~n59240 & ~n22372;
  assign n22374 = n59240 & n22325;
  assign n22375 = ~pi628 & ~n22372;
  assign n22376 = pi628 & n22325;
  assign n22377 = ~n22375 & ~n22376;
  assign n22378 = ~pi1156 & ~n22377;
  assign n22379 = pi628 & ~n22372;
  assign n22380 = ~pi628 & n22325;
  assign n22381 = ~n22379 & ~n22380;
  assign n22382 = pi1156 & ~n22381;
  assign n22383 = ~n22378 & ~n22382;
  assign n22384 = pi792 & ~n22383;
  assign n22385 = ~pi792 & ~n22372;
  assign n22386 = ~n22384 & ~n22385;
  assign n22387 = n59240 & ~n22325;
  assign n22388 = ~n59240 & n22372;
  assign n22389 = ~n22387 & ~n22388;
  assign n22390 = ~n22373 & ~n22374;
  assign n22391 = ~n9743 & ~n59798;
  assign n22392 = n9743 & n22325;
  assign n22393 = ~pi647 & ~n59798;
  assign n22394 = pi647 & n22325;
  assign n22395 = ~n22393 & ~n22394;
  assign n22396 = ~pi1157 & ~n22395;
  assign n22397 = pi647 & ~n59798;
  assign n22398 = ~pi647 & n22325;
  assign n22399 = ~n22397 & ~n22398;
  assign n22400 = pi1157 & ~n22399;
  assign n22401 = ~n22396 & ~n22400;
  assign n22402 = pi787 & ~n22401;
  assign n22403 = ~pi787 & ~n59798;
  assign n22404 = ~n22402 & ~n22403;
  assign n22405 = ~n22391 & ~n22392;
  assign n22406 = ~pi644 & ~n59799;
  assign n22407 = pi715 & ~n22406;
  assign n22408 = ~pi764 & n6654;
  assign n22409 = pi192 & n6853;
  assign n22410 = ~n22408 & ~n22409;
  assign n22411 = pi39 & ~n22410;
  assign n22412 = ~pi192 & pi764;
  assign n22413 = n59164 & n22412;
  assign n22414 = ~pi764 & n8180;
  assign n22415 = pi764 & ~n6799;
  assign n22416 = pi192 & ~n22415;
  assign n22417 = ~n22414 & ~n22416;
  assign n22418 = ~n22413 & n22417;
  assign n22419 = ~n22411 & n22418;
  assign n22420 = ~pi38 & ~n22419;
  assign n22421 = pi764 & n6865;
  assign n22422 = pi38 & ~n22332;
  assign n22423 = ~n22421 & n22422;
  assign n22424 = ~n22420 & ~n22423;
  assign n22425 = n59132 & ~n22424;
  assign n22426 = ~n22327 & ~n22425;
  assign n22427 = ~n7597 & ~n22426;
  assign n22428 = n7597 & ~n22325;
  assign n22429 = ~n22427 & ~n22428;
  assign n22430 = ~pi785 & ~n22429;
  assign n22431 = ~n7598 & ~n22325;
  assign n22432 = pi609 & n22427;
  assign n22433 = ~n22431 & ~n22432;
  assign n22434 = pi1155 & ~n22433;
  assign n22435 = ~n7610 & ~n22325;
  assign n22436 = ~pi609 & n22427;
  assign n22437 = ~n22435 & ~n22436;
  assign n22438 = ~pi1155 & ~n22437;
  assign n22439 = ~n22434 & ~n22438;
  assign n22440 = pi785 & ~n22439;
  assign n22441 = ~n22430 & ~n22440;
  assign n22442 = ~pi781 & ~n22441;
  assign n22443 = pi618 & n22441;
  assign n22444 = ~pi618 & n22325;
  assign n22445 = pi1154 & ~n22444;
  assign n22446 = ~n22443 & n22445;
  assign n22447 = ~pi618 & n22441;
  assign n22448 = pi618 & n22325;
  assign n22449 = ~pi1154 & ~n22448;
  assign n22450 = ~n22447 & n22449;
  assign n22451 = ~n22446 & ~n22450;
  assign n22452 = pi781 & ~n22451;
  assign n22453 = ~n22442 & ~n22452;
  assign n22454 = ~pi789 & ~n22453;
  assign n22455 = pi619 & n22453;
  assign n22456 = ~pi619 & n22325;
  assign n22457 = pi1159 & ~n22456;
  assign n22458 = ~n22455 & n22457;
  assign n22459 = ~pi619 & n22453;
  assign n22460 = pi619 & n22325;
  assign n22461 = ~pi1159 & ~n22460;
  assign n22462 = ~n22459 & n22461;
  assign n22463 = ~n22458 & ~n22462;
  assign n22464 = pi789 & ~n22463;
  assign n22465 = ~n22454 & ~n22464;
  assign n22466 = ~n8054 & n22465;
  assign n22467 = n8054 & n22325;
  assign n22468 = ~n22466 & ~n22467;
  assign n22469 = ~n7793 & ~n22468;
  assign n22470 = n7793 & n22325;
  assign n22471 = ~n22469 & ~n22470;
  assign n22472 = ~n7835 & ~n22471;
  assign n22473 = n7835 & n22325;
  assign n22474 = n7835 & ~n22325;
  assign n22475 = ~n7835 & n22471;
  assign n22476 = ~n22474 & ~n22475;
  assign n22477 = ~n22472 & ~n22473;
  assign n22478 = pi644 & n59800;
  assign n22479 = ~pi644 & n22325;
  assign n22480 = ~pi715 & ~n22479;
  assign n22481 = ~n22478 & n22480;
  assign n22482 = pi1160 & ~n22481;
  assign n22483 = ~n22407 & n22482;
  assign n22484 = pi644 & ~n59799;
  assign n22485 = ~pi715 & ~n22484;
  assign n22486 = ~pi644 & n59800;
  assign n22487 = pi644 & n22325;
  assign n22488 = pi715 & ~n22487;
  assign n22489 = ~n22486 & n22488;
  assign n22490 = ~pi1160 & ~n22489;
  assign n22491 = ~n22485 & n22490;
  assign n22492 = ~n22483 & ~n22491;
  assign n22493 = pi790 & ~n22492;
  assign n22494 = ~pi644 & n22490;
  assign n22495 = pi644 & n22482;
  assign n22496 = pi790 & ~n22495;
  assign n22497 = pi790 & ~n22494;
  assign n22498 = ~n22495 & n22497;
  assign n22499 = ~n22494 & n22496;
  assign n22500 = ~n7872 & n22471;
  assign n22501 = n7832 & ~n22398;
  assign n22502 = n7832 & n22399;
  assign n22503 = ~n22397 & n22501;
  assign n22504 = n7833 & ~n22394;
  assign n22505 = n7833 & n22395;
  assign n22506 = ~n22393 & n22504;
  assign n22507 = ~n59802 & ~n59803;
  assign n22508 = ~n22500 & ~n59803;
  assign n22509 = ~n59802 & n22508;
  assign n22510 = ~n22500 & n22507;
  assign n22511 = pi787 & ~n59804;
  assign n22512 = ~n11154 & n22468;
  assign n22513 = n7791 & ~n22376;
  assign n22514 = n7791 & n22377;
  assign n22515 = ~n22375 & n22513;
  assign n22516 = n7790 & ~n22380;
  assign n22517 = n7790 & n22381;
  assign n22518 = ~n22379 & n22516;
  assign n22519 = ~n59805 & ~n59806;
  assign n22520 = ~n22512 & n22519;
  assign n22521 = pi792 & ~n22520;
  assign n22522 = ~pi691 & n22424;
  assign n22523 = ~pi192 & n59177;
  assign n22524 = pi192 & n7111;
  assign n22525 = ~pi764 & ~n22524;
  assign n22526 = ~n22523 & n22525;
  assign n22527 = pi192 & n7188;
  assign n22528 = ~pi192 & ~n59203;
  assign n22529 = pi764 & ~n22528;
  assign n22530 = ~n22527 & n22529;
  assign n22531 = pi39 & ~n22530;
  assign n22532 = ~n22526 & n22531;
  assign n22533 = ~pi192 & n7310;
  assign n22534 = pi192 & n7333;
  assign n22535 = ~pi764 & ~n22534;
  assign n22536 = ~pi764 & ~n22533;
  assign n22537 = ~n22534 & n22536;
  assign n22538 = ~n22533 & n22535;
  assign n22539 = ~pi192 & ~n7339;
  assign n22540 = pi192 & ~n7347;
  assign n22541 = pi764 & ~n22540;
  assign n22542 = ~n22539 & n22541;
  assign n22543 = ~pi39 & ~n22542;
  assign n22544 = ~n59807 & n22543;
  assign n22545 = ~pi38 & ~n22544;
  assign n22546 = ~pi192 & n8213;
  assign n22547 = pi192 & n8217;
  assign n22548 = ~pi764 & ~n22547;
  assign n22549 = ~n22546 & n22548;
  assign n22550 = pi192 & n9808;
  assign n22551 = ~pi192 & ~n13062;
  assign n22552 = pi764 & ~n22551;
  assign n22553 = ~n22550 & n22552;
  assign n22554 = ~n22549 & ~n22553;
  assign n22555 = ~pi38 & ~n22554;
  assign n22556 = ~n22532 & n22545;
  assign n22557 = ~pi764 & n13069;
  assign n22558 = ~n7222 & ~n22557;
  assign n22559 = ~pi39 & ~n22558;
  assign n22560 = ~pi192 & ~n22559;
  assign n22561 = ~n7056 & ~n22118;
  assign n22562 = pi192 & ~n22561;
  assign n22563 = n59171 & n22562;
  assign n22564 = pi38 & ~n22563;
  assign n22565 = ~n22560 & n22564;
  assign n22566 = pi691 & ~n22565;
  assign n22567 = ~n59808 & n22566;
  assign n22568 = n59132 & ~n22567;
  assign n22569 = n59132 & ~n22522;
  assign n22570 = ~n22567 & n22569;
  assign n22571 = ~n22522 & n22568;
  assign n22572 = ~n22327 & ~n59809;
  assign n22573 = ~pi625 & n22572;
  assign n22574 = pi625 & n22426;
  assign n22575 = ~pi1153 & ~n22574;
  assign n22576 = ~n22573 & n22575;
  assign n22577 = ~pi608 & ~n22345;
  assign n22578 = ~n22576 & n22577;
  assign n22579 = pi625 & n22572;
  assign n22580 = ~pi625 & n22426;
  assign n22581 = pi1153 & ~n22580;
  assign n22582 = ~n22579 & n22581;
  assign n22583 = pi608 & ~n22349;
  assign n22584 = ~n22582 & n22583;
  assign n22585 = ~n22578 & ~n22584;
  assign n22586 = pi778 & ~n22585;
  assign n22587 = ~pi778 & n22572;
  assign n22588 = ~n22586 & ~n22587;
  assign n22589 = ~pi609 & ~n22588;
  assign n22590 = pi609 & n22352;
  assign n22591 = ~pi1155 & ~n22590;
  assign n22592 = ~n22589 & n22591;
  assign n22593 = ~pi660 & ~n22434;
  assign n22594 = ~n22592 & n22593;
  assign n22595 = pi609 & ~n22588;
  assign n22596 = ~pi609 & n22352;
  assign n22597 = pi1155 & ~n22596;
  assign n22598 = ~n22595 & n22597;
  assign n22599 = pi660 & ~n22438;
  assign n22600 = ~n22598 & n22599;
  assign n22601 = ~n22594 & ~n22600;
  assign n22602 = pi785 & ~n22601;
  assign n22603 = ~pi785 & ~n22588;
  assign n22604 = ~n22602 & ~n22603;
  assign n22605 = ~pi618 & ~n22604;
  assign n22606 = pi618 & n59795;
  assign n22607 = ~pi1154 & ~n22606;
  assign n22608 = ~n22605 & n22607;
  assign n22609 = ~pi627 & ~n22446;
  assign n22610 = ~n22608 & n22609;
  assign n22611 = pi618 & ~n22604;
  assign n22612 = ~pi618 & n59795;
  assign n22613 = pi1154 & ~n22612;
  assign n22614 = ~n22611 & n22613;
  assign n22615 = pi627 & ~n22450;
  assign n22616 = ~n22614 & n22615;
  assign n22617 = ~n22610 & ~n22616;
  assign n22618 = pi781 & ~n22617;
  assign n22619 = ~pi781 & ~n22604;
  assign n22620 = ~n22618 & ~n22619;
  assign n22621 = pi619 & ~n22620;
  assign n22622 = ~pi619 & ~n59796;
  assign n22623 = pi1159 & ~n22622;
  assign n22624 = ~n22621 & n22623;
  assign n22625 = pi648 & ~n22462;
  assign n22626 = ~n22624 & n22625;
  assign n22627 = ~pi619 & ~n22620;
  assign n22628 = pi619 & ~n59796;
  assign n22629 = ~pi1159 & ~n22628;
  assign n22630 = ~n22627 & n22629;
  assign n22631 = ~pi648 & ~n22458;
  assign n22632 = ~n22630 & n22631;
  assign n22633 = pi789 & ~n22632;
  assign n22634 = pi789 & ~n22626;
  assign n22635 = ~n22632 & n22634;
  assign n22636 = ~n22626 & n22633;
  assign n22637 = ~pi789 & n22620;
  assign n22638 = n59242 & ~n22637;
  assign n22639 = ~n59810 & n22638;
  assign n22640 = ~pi626 & ~n22465;
  assign n22641 = pi626 & ~n22325;
  assign n22642 = n7760 & ~n22641;
  assign n22643 = ~n22640 & n22642;
  assign n22644 = n7984 & n59797;
  assign n22645 = pi626 & ~n22465;
  assign n22646 = ~pi626 & ~n22325;
  assign n22647 = n7759 & ~n22646;
  assign n22648 = ~n22645 & n22647;
  assign n22649 = ~n22644 & ~n22648;
  assign n22650 = ~n22643 & ~n22644;
  assign n22651 = ~n22648 & n22650;
  assign n22652 = ~n22643 & n22649;
  assign n22653 = pi788 & ~n59811;
  assign n22654 = ~n59357 & ~n22653;
  assign n22655 = ~n22639 & n22654;
  assign n22656 = ~n22521 & ~n22655;
  assign n22657 = ~n8108 & ~n22656;
  assign n22658 = ~n22511 & ~n22657;
  assign n22659 = ~n59801 & n22658;
  assign n22660 = ~n22493 & ~n22659;
  assign n22661 = n58992 & ~n22660;
  assign n22662 = ~pi192 & ~n58992;
  assign n22663 = ~pi832 & ~n22662;
  assign n22664 = ~n22661 & n22663;
  assign po349 = ~n22324 & ~n22664;
  assign n22666 = ~pi193 & ~n2794;
  assign n22667 = pi739 & n6822;
  assign n22668 = ~n22666 & ~n22667;
  assign n22669 = ~n7875 & ~n22668;
  assign n22670 = ~pi785 & ~n22669;
  assign n22671 = n7610 & n22667;
  assign n22672 = n22669 & ~n22671;
  assign n22673 = pi1155 & ~n22672;
  assign n22674 = ~pi1155 & ~n22666;
  assign n22675 = ~n22671 & n22674;
  assign n22676 = ~n22673 & ~n22675;
  assign n22677 = pi785 & ~n22676;
  assign n22678 = ~n22670 & ~n22677;
  assign n22679 = ~pi781 & ~n22678;
  assign n22680 = ~n7890 & n22678;
  assign n22681 = pi1154 & ~n22680;
  assign n22682 = ~n7893 & n22678;
  assign n22683 = ~pi1154 & ~n22682;
  assign n22684 = ~n22681 & ~n22683;
  assign n22685 = pi781 & ~n22684;
  assign n22686 = ~n22679 & ~n22685;
  assign n22687 = ~pi789 & ~n22686;
  assign n22688 = ~n11882 & n22686;
  assign n22689 = pi1159 & ~n22688;
  assign n22690 = ~n11885 & n22686;
  assign n22691 = ~pi1159 & ~n22690;
  assign n22692 = ~n22689 & ~n22691;
  assign n22693 = pi789 & ~n22692;
  assign n22694 = ~n22687 & ~n22693;
  assign n22695 = ~n8054 & ~n22694;
  assign n22696 = n8054 & ~n22666;
  assign n22697 = ~n8054 & n22694;
  assign n22698 = n8054 & n22666;
  assign n22699 = ~n22697 & ~n22698;
  assign n22700 = ~n22695 & ~n22696;
  assign n22701 = ~n7793 & ~n59812;
  assign n22702 = n7793 & n22666;
  assign n22703 = ~n7872 & ~n22702;
  assign n22704 = ~n22701 & ~n22702;
  assign n22705 = ~n7872 & n22704;
  assign n22706 = ~n22701 & n22703;
  assign n22707 = pi690 & n7055;
  assign n22708 = ~n22666 & ~n22707;
  assign n22709 = ~pi778 & ~n22708;
  assign n22710 = ~pi625 & n22707;
  assign n22711 = ~n22708 & ~n22710;
  assign n22712 = pi1153 & ~n22711;
  assign n22713 = ~pi1153 & ~n22666;
  assign n22714 = ~n22710 & n22713;
  assign n22715 = pi778 & ~n22714;
  assign n22716 = ~n22712 & n22715;
  assign n22717 = ~n22709 & ~n22716;
  assign n22718 = ~n7949 & ~n22717;
  assign n22719 = ~n7951 & n22718;
  assign n22720 = ~n7953 & n22719;
  assign n22721 = ~n7955 & n22720;
  assign n22722 = ~n7967 & n22721;
  assign n22723 = pi647 & ~n22722;
  assign n22724 = ~pi647 & ~n22666;
  assign n22725 = ~n22723 & ~n22724;
  assign n22726 = n7832 & ~n22725;
  assign n22727 = ~pi647 & n22722;
  assign n22728 = pi647 & n22666;
  assign n22729 = ~pi1157 & ~n22728;
  assign n22730 = ~n22727 & n22729;
  assign n22731 = pi630 & n22730;
  assign n22732 = ~n22726 & ~n22731;
  assign n22733 = ~n59813 & n22732;
  assign n22734 = pi787 & ~n22733;
  assign n22735 = ~pi626 & ~n22694;
  assign n22736 = pi626 & ~n22666;
  assign n22737 = n7760 & ~n22736;
  assign n22738 = ~n22735 & n22737;
  assign n22739 = n7984 & n22720;
  assign n22740 = pi626 & ~n22694;
  assign n22741 = ~pi626 & ~n22666;
  assign n22742 = n7759 & ~n22741;
  assign n22743 = ~n22740 & n22742;
  assign n22744 = ~n22739 & ~n22743;
  assign n22745 = ~n22738 & ~n22739;
  assign n22746 = ~n22743 & n22745;
  assign n22747 = ~n22738 & n22744;
  assign n22748 = pi788 & ~n59814;
  assign n22749 = ~n6701 & ~n22708;
  assign n22750 = pi625 & n22749;
  assign n22751 = n22668 & ~n22749;
  assign n22752 = ~n22750 & ~n22751;
  assign n22753 = n22713 & ~n22752;
  assign n22754 = ~pi608 & ~n22712;
  assign n22755 = ~n22753 & n22754;
  assign n22756 = pi1153 & n22668;
  assign n22757 = ~n22750 & n22756;
  assign n22758 = pi608 & ~n22714;
  assign n22759 = ~n22757 & n22758;
  assign n22760 = ~n22755 & ~n22759;
  assign n22761 = pi778 & ~n22760;
  assign n22762 = ~pi778 & ~n22751;
  assign n22763 = ~n22761 & ~n22762;
  assign n22764 = ~pi609 & ~n22763;
  assign n22765 = pi609 & ~n22717;
  assign n22766 = ~pi1155 & ~n22765;
  assign n22767 = ~n22764 & n22766;
  assign n22768 = ~pi660 & ~n22673;
  assign n22769 = ~n22767 & n22768;
  assign n22770 = pi609 & ~n22763;
  assign n22771 = ~pi609 & ~n22717;
  assign n22772 = pi1155 & ~n22771;
  assign n22773 = ~n22770 & n22772;
  assign n22774 = pi660 & ~n22675;
  assign n22775 = ~n22773 & n22774;
  assign n22776 = ~n22769 & ~n22775;
  assign n22777 = pi785 & ~n22776;
  assign n22778 = ~pi785 & ~n22763;
  assign n22779 = ~n22777 & ~n22778;
  assign n22780 = ~pi618 & ~n22779;
  assign n22781 = pi618 & n22718;
  assign n22782 = ~pi1154 & ~n22781;
  assign n22783 = ~n22780 & n22782;
  assign n22784 = ~pi627 & ~n22681;
  assign n22785 = ~n22783 & n22784;
  assign n22786 = pi618 & ~n22779;
  assign n22787 = ~pi618 & n22718;
  assign n22788 = pi1154 & ~n22787;
  assign n22789 = ~n22786 & n22788;
  assign n22790 = pi627 & ~n22683;
  assign n22791 = ~n22789 & n22790;
  assign n22792 = ~n22785 & ~n22791;
  assign n22793 = pi781 & ~n22792;
  assign n22794 = ~pi781 & ~n22779;
  assign n22795 = ~n22793 & ~n22794;
  assign n22796 = pi619 & ~n22795;
  assign n22797 = ~pi619 & n22719;
  assign n22798 = pi1159 & ~n22797;
  assign n22799 = ~n22796 & n22798;
  assign n22800 = pi648 & ~n22691;
  assign n22801 = ~n22799 & n22800;
  assign n22802 = ~pi619 & ~n22795;
  assign n22803 = pi619 & n22719;
  assign n22804 = ~pi1159 & ~n22803;
  assign n22805 = ~n22802 & n22804;
  assign n22806 = ~pi648 & ~n22689;
  assign n22807 = ~n22805 & n22806;
  assign n22808 = pi789 & ~n22807;
  assign n22809 = pi789 & ~n22801;
  assign n22810 = ~n22807 & n22809;
  assign n22811 = ~n22801 & n22808;
  assign n22812 = ~pi789 & n22795;
  assign n22813 = n59242 & ~n22812;
  assign n22814 = ~n59815 & n22813;
  assign n22815 = ~n22748 & ~n22814;
  assign n22816 = ~n59357 & ~n22815;
  assign n22817 = n7957 & ~n59812;
  assign n22818 = n8065 & n22721;
  assign n22819 = pi629 & ~n22818;
  assign n22820 = ~n22817 & n22819;
  assign n22821 = n7958 & ~n59812;
  assign n22822 = n8074 & n22721;
  assign n22823 = ~pi629 & ~n22822;
  assign n22824 = ~n22821 & n22823;
  assign n22825 = pi792 & ~n22824;
  assign n22826 = ~n22821 & ~n22822;
  assign n22827 = ~pi629 & ~n22826;
  assign n22828 = ~n22817 & ~n22818;
  assign n22829 = pi629 & ~n22828;
  assign n22830 = ~n22827 & ~n22829;
  assign n22831 = pi792 & ~n22830;
  assign n22832 = pi792 & ~n22820;
  assign n22833 = ~n22824 & n22832;
  assign n22834 = ~n22820 & n22825;
  assign n22835 = ~n8108 & ~n59816;
  assign n22836 = ~n22816 & n22835;
  assign n22837 = ~n22734 & ~n22836;
  assign n22838 = pi644 & n22837;
  assign n22839 = ~pi787 & ~n22722;
  assign n22840 = pi1157 & ~n22725;
  assign n22841 = ~n22730 & ~n22840;
  assign n22842 = pi787 & ~n22841;
  assign n22843 = ~n22839 & ~n22842;
  assign n22844 = ~pi644 & n22843;
  assign n22845 = pi715 & ~n22844;
  assign n22846 = ~n22838 & n22845;
  assign n22847 = ~n11491 & n22666;
  assign n22848 = ~n7835 & n22701;
  assign n22849 = ~n7835 & ~n22704;
  assign n22850 = n7835 & n22666;
  assign n22851 = ~n22849 & ~n22850;
  assign n22852 = ~n22847 & ~n22848;
  assign n22853 = pi644 & ~n59817;
  assign n22854 = ~pi644 & n22666;
  assign n22855 = ~pi715 & ~n22854;
  assign n22856 = ~n22853 & n22855;
  assign n22857 = pi1160 & ~n22856;
  assign n22858 = ~n22846 & n22857;
  assign n22859 = ~pi644 & n22837;
  assign n22860 = pi644 & n22843;
  assign n22861 = ~pi715 & ~n22860;
  assign n22862 = ~n22859 & n22861;
  assign n22863 = ~pi644 & ~n59817;
  assign n22864 = pi644 & n22666;
  assign n22865 = pi715 & ~n22864;
  assign n22866 = ~n22863 & n22865;
  assign n22867 = ~pi1160 & ~n22866;
  assign n22868 = ~n22862 & n22867;
  assign n22869 = ~n22858 & ~n22868;
  assign n22870 = pi790 & ~n22869;
  assign n22871 = ~pi790 & n22837;
  assign n22872 = pi832 & ~n22871;
  assign n22873 = ~n22870 & n22872;
  assign n22874 = ~pi193 & ~n7560;
  assign n22875 = n59231 & ~n22874;
  assign n22876 = pi690 & n59132;
  assign n22877 = n22874 & ~n22876;
  assign n22878 = pi193 & n59251;
  assign n22879 = ~pi38 & ~n22878;
  assign n22880 = n59132 & ~n22879;
  assign n22881 = ~pi193 & n8249;
  assign n22882 = ~n22880 & ~n22881;
  assign n22883 = ~pi193 & ~n6863;
  assign n22884 = n7547 & ~n22883;
  assign n22885 = pi690 & ~n22884;
  assign n22886 = ~n22882 & n22885;
  assign n22887 = ~n22877 & ~n22886;
  assign n22888 = ~pi778 & n22887;
  assign n22889 = pi625 & ~n22887;
  assign n22890 = ~pi625 & n22874;
  assign n22891 = pi1153 & ~n22890;
  assign n22892 = ~n22889 & n22891;
  assign n22893 = ~pi625 & ~n22887;
  assign n22894 = pi625 & n22874;
  assign n22895 = ~pi1153 & ~n22894;
  assign n22896 = ~n22893 & n22895;
  assign n22897 = ~n22892 & ~n22896;
  assign n22898 = pi778 & ~n22897;
  assign n22899 = ~n22888 & ~n22898;
  assign n22900 = ~n59229 & n22899;
  assign n22901 = n59229 & n22874;
  assign n22902 = n59229 & ~n22874;
  assign n22903 = ~n59229 & ~n22899;
  assign n22904 = ~n22902 & ~n22903;
  assign n22905 = ~n22900 & ~n22901;
  assign n22906 = ~n59231 & ~n59818;
  assign n22907 = ~n59231 & n59818;
  assign n22908 = n59231 & n22874;
  assign n22909 = ~n22907 & ~n22908;
  assign n22910 = ~n22875 & ~n22906;
  assign n22911 = ~n7716 & ~n59819;
  assign n22912 = n7716 & n22874;
  assign n22913 = n7716 & ~n22874;
  assign n22914 = ~n7716 & n59819;
  assign n22915 = ~n22913 & ~n22914;
  assign n22916 = ~n22911 & ~n22912;
  assign n22917 = ~n7762 & n59820;
  assign n22918 = n7762 & n22874;
  assign n22919 = ~n22917 & ~n22918;
  assign n22920 = ~pi792 & n22919;
  assign n22921 = pi628 & ~n22919;
  assign n22922 = ~pi628 & n22874;
  assign n22923 = pi1156 & ~n22922;
  assign n22924 = ~n22921 & n22923;
  assign n22925 = ~pi628 & ~n22919;
  assign n22926 = pi628 & n22874;
  assign n22927 = ~pi1156 & ~n22926;
  assign n22928 = ~n22925 & n22927;
  assign n22929 = ~n22924 & ~n22928;
  assign n22930 = pi792 & ~n22929;
  assign n22931 = ~n22920 & ~n22930;
  assign n22932 = pi647 & n22931;
  assign n22933 = ~pi647 & n22874;
  assign n22934 = pi647 & ~n22931;
  assign n22935 = ~pi647 & ~n22874;
  assign n22936 = ~n22934 & ~n22935;
  assign n22937 = ~n22932 & ~n22933;
  assign n22938 = pi1157 & ~n59821;
  assign n22939 = ~pi647 & n22931;
  assign n22940 = pi647 & n22874;
  assign n22941 = ~pi1157 & ~n22940;
  assign n22942 = ~n22939 & n22941;
  assign n22943 = ~pi647 & ~n22931;
  assign n22944 = pi647 & ~n22874;
  assign n22945 = ~n22943 & ~n22944;
  assign n22946 = ~pi1157 & n22945;
  assign n22947 = pi1157 & n59821;
  assign n22948 = ~n22946 & ~n22947;
  assign n22949 = ~n22938 & ~n22942;
  assign n22950 = pi787 & n59822;
  assign n22951 = ~pi787 & ~n22931;
  assign n22952 = pi787 & ~n59822;
  assign n22953 = ~pi787 & n22931;
  assign n22954 = ~n22952 & ~n22953;
  assign n22955 = ~n22950 & ~n22951;
  assign n22956 = ~pi644 & ~n59823;
  assign n22957 = pi715 & ~n22956;
  assign n22958 = pi193 & ~n59132;
  assign n22959 = pi739 & n6865;
  assign n22960 = ~n22883 & ~n22959;
  assign n22961 = pi38 & ~n22960;
  assign n22962 = ~pi193 & n59164;
  assign n22963 = pi193 & ~n6855;
  assign n22964 = pi739 & ~n22963;
  assign n22965 = ~n22962 & n22964;
  assign n22966 = ~pi193 & ~pi739;
  assign n22967 = ~n6656 & n22966;
  assign n22968 = ~n22965 & ~n22967;
  assign n22969 = ~pi38 & ~n22968;
  assign n22970 = ~n22961 & ~n22969;
  assign n22971 = n59132 & n22970;
  assign n22972 = ~n22958 & ~n22971;
  assign n22973 = ~n7597 & ~n22972;
  assign n22974 = n7597 & ~n22874;
  assign n22975 = ~n22973 & ~n22974;
  assign n22976 = ~pi785 & ~n22975;
  assign n22977 = ~n7598 & ~n22874;
  assign n22978 = pi609 & n22973;
  assign n22979 = ~n22977 & ~n22978;
  assign n22980 = pi1155 & ~n22979;
  assign n22981 = ~n7610 & ~n22874;
  assign n22982 = ~pi609 & n22973;
  assign n22983 = ~n22981 & ~n22982;
  assign n22984 = ~pi1155 & ~n22983;
  assign n22985 = ~n22980 & ~n22984;
  assign n22986 = pi785 & ~n22985;
  assign n22987 = ~n22976 & ~n22986;
  assign n22988 = ~pi781 & ~n22987;
  assign n22989 = pi618 & n22987;
  assign n22990 = ~pi618 & n22874;
  assign n22991 = pi1154 & ~n22990;
  assign n22992 = ~n22989 & n22991;
  assign n22993 = ~pi618 & n22987;
  assign n22994 = pi618 & n22874;
  assign n22995 = ~pi1154 & ~n22994;
  assign n22996 = ~n22993 & n22995;
  assign n22997 = ~n22992 & ~n22996;
  assign n22998 = pi781 & ~n22997;
  assign n22999 = ~n22988 & ~n22998;
  assign n23000 = ~pi789 & ~n22999;
  assign n23001 = pi619 & n22999;
  assign n23002 = ~pi619 & n22874;
  assign n23003 = pi1159 & ~n23002;
  assign n23004 = ~n23001 & n23003;
  assign n23005 = ~pi619 & n22999;
  assign n23006 = pi619 & n22874;
  assign n23007 = ~pi1159 & ~n23006;
  assign n23008 = ~n23005 & n23007;
  assign n23009 = ~n23004 & ~n23008;
  assign n23010 = pi789 & ~n23009;
  assign n23011 = ~n23000 & ~n23010;
  assign n23012 = ~n8054 & n23011;
  assign n23013 = n8054 & n22874;
  assign n23014 = ~n23012 & ~n23013;
  assign n23015 = ~n7793 & ~n23014;
  assign n23016 = n7793 & n22874;
  assign n23017 = ~n23015 & ~n23016;
  assign n23018 = ~n7835 & ~n23017;
  assign n23019 = n7835 & n22874;
  assign n23020 = n7835 & ~n22874;
  assign n23021 = ~n7835 & n23017;
  assign n23022 = ~n23020 & ~n23021;
  assign n23023 = ~n23018 & ~n23019;
  assign n23024 = pi644 & n59824;
  assign n23025 = ~pi644 & n22874;
  assign n23026 = ~pi715 & ~n23025;
  assign n23027 = ~n23024 & n23026;
  assign n23028 = pi1160 & ~n23027;
  assign n23029 = ~n22957 & n23028;
  assign n23030 = pi644 & ~n59823;
  assign n23031 = ~pi715 & ~n23030;
  assign n23032 = ~pi644 & n59824;
  assign n23033 = pi644 & n22874;
  assign n23034 = pi715 & ~n23033;
  assign n23035 = ~n23032 & n23034;
  assign n23036 = ~pi1160 & ~n23035;
  assign n23037 = ~n23031 & n23036;
  assign n23038 = ~n23029 & ~n23037;
  assign n23039 = pi790 & ~n23038;
  assign n23040 = ~pi644 & n23036;
  assign n23041 = pi644 & n23028;
  assign n23042 = pi790 & ~n23041;
  assign n23043 = pi790 & ~n23040;
  assign n23044 = ~n23041 & n23043;
  assign n23045 = ~n23040 & n23042;
  assign n23046 = ~n7872 & n23017;
  assign n23047 = n7832 & ~n59821;
  assign n23048 = n7833 & ~n22945;
  assign n23049 = pi630 & n22942;
  assign n23050 = ~n23047 & ~n59826;
  assign n23051 = ~n23046 & n23050;
  assign n23052 = pi787 & ~n23051;
  assign n23053 = ~n11154 & n23014;
  assign n23054 = ~pi629 & n22924;
  assign n23055 = pi629 & n22928;
  assign n23056 = ~n23054 & ~n23055;
  assign n23057 = ~n23053 & n23056;
  assign n23058 = pi792 & ~n23057;
  assign n23059 = ~pi690 & ~n22970;
  assign n23060 = ~pi193 & n59177;
  assign n23061 = pi193 & n7111;
  assign n23062 = ~pi739 & ~n23061;
  assign n23063 = ~n23060 & n23062;
  assign n23064 = pi193 & n7188;
  assign n23065 = ~pi193 & ~n59203;
  assign n23066 = pi739 & ~n23065;
  assign n23067 = ~n23064 & n23066;
  assign n23068 = pi39 & ~n23067;
  assign n23069 = ~n23063 & n23068;
  assign n23070 = pi193 & n7333;
  assign n23071 = ~pi193 & n7310;
  assign n23072 = ~pi739 & ~n23071;
  assign n23073 = ~n23070 & n23072;
  assign n23074 = ~pi193 & ~n7339;
  assign n23075 = pi193 & ~n7347;
  assign n23076 = pi739 & ~n23075;
  assign n23077 = ~n23074 & n23076;
  assign n23078 = ~pi39 & ~n23077;
  assign n23079 = ~pi193 & n7339;
  assign n23080 = pi193 & n7347;
  assign n23081 = pi739 & ~n23080;
  assign n23082 = ~n23079 & n23081;
  assign n23083 = pi193 & ~n7333;
  assign n23084 = ~pi193 & ~n7310;
  assign n23085 = ~pi739 & ~n23084;
  assign n23086 = ~pi739 & ~n23083;
  assign n23087 = ~n23084 & n23086;
  assign n23088 = ~n23083 & n23085;
  assign n23089 = ~n23082 & ~n59827;
  assign n23090 = ~pi39 & ~n23089;
  assign n23091 = ~n23073 & n23078;
  assign n23092 = ~pi38 & ~n59828;
  assign n23093 = ~n23069 & n23092;
  assign n23094 = ~pi739 & n13069;
  assign n23095 = ~n7222 & ~n23094;
  assign n23096 = ~pi39 & ~n23095;
  assign n23097 = ~pi193 & ~n23096;
  assign n23098 = ~n7056 & ~n22667;
  assign n23099 = pi193 & ~n23098;
  assign n23100 = n59171 & n23099;
  assign n23101 = pi38 & ~n23100;
  assign n23102 = ~n23097 & n23101;
  assign n23103 = pi690 & ~n23102;
  assign n23104 = ~n23093 & n23103;
  assign n23105 = n59132 & ~n23104;
  assign n23106 = ~n23059 & n23105;
  assign n23107 = ~n22958 & ~n23106;
  assign n23108 = ~pi625 & n23107;
  assign n23109 = pi625 & n22972;
  assign n23110 = ~pi1153 & ~n23109;
  assign n23111 = ~n23108 & n23110;
  assign n23112 = ~pi608 & ~n22892;
  assign n23113 = ~n23111 & n23112;
  assign n23114 = pi625 & n23107;
  assign n23115 = ~pi625 & n22972;
  assign n23116 = pi1153 & ~n23115;
  assign n23117 = ~n23114 & n23116;
  assign n23118 = pi608 & ~n22896;
  assign n23119 = ~n23117 & n23118;
  assign n23120 = ~n23113 & ~n23119;
  assign n23121 = pi778 & ~n23120;
  assign n23122 = ~pi778 & n23107;
  assign n23123 = ~n23121 & ~n23122;
  assign n23124 = ~pi609 & ~n23123;
  assign n23125 = pi609 & n22899;
  assign n23126 = ~pi1155 & ~n23125;
  assign n23127 = ~n23124 & n23126;
  assign n23128 = ~pi660 & ~n22980;
  assign n23129 = ~n23127 & n23128;
  assign n23130 = pi609 & ~n23123;
  assign n23131 = ~pi609 & n22899;
  assign n23132 = pi1155 & ~n23131;
  assign n23133 = ~n23130 & n23132;
  assign n23134 = pi660 & ~n22984;
  assign n23135 = ~n23133 & n23134;
  assign n23136 = ~n23129 & ~n23135;
  assign n23137 = pi785 & ~n23136;
  assign n23138 = ~pi785 & ~n23123;
  assign n23139 = ~n23137 & ~n23138;
  assign n23140 = ~pi618 & ~n23139;
  assign n23141 = pi618 & n59818;
  assign n23142 = ~pi1154 & ~n23141;
  assign n23143 = ~n23140 & n23142;
  assign n23144 = ~pi627 & ~n22992;
  assign n23145 = ~n23143 & n23144;
  assign n23146 = pi618 & ~n23139;
  assign n23147 = ~pi618 & n59818;
  assign n23148 = pi1154 & ~n23147;
  assign n23149 = ~n23146 & n23148;
  assign n23150 = pi627 & ~n22996;
  assign n23151 = ~n23149 & n23150;
  assign n23152 = ~n23145 & ~n23151;
  assign n23153 = pi781 & ~n23152;
  assign n23154 = ~pi781 & ~n23139;
  assign n23155 = ~n23153 & ~n23154;
  assign n23156 = pi619 & ~n23155;
  assign n23157 = ~pi619 & ~n59819;
  assign n23158 = pi1159 & ~n23157;
  assign n23159 = ~n23156 & n23158;
  assign n23160 = pi648 & ~n23008;
  assign n23161 = ~n23159 & n23160;
  assign n23162 = ~pi619 & ~n23155;
  assign n23163 = pi619 & ~n59819;
  assign n23164 = ~pi1159 & ~n23163;
  assign n23165 = ~n23162 & n23164;
  assign n23166 = ~pi648 & ~n23004;
  assign n23167 = ~n23165 & n23166;
  assign n23168 = pi789 & ~n23167;
  assign n23169 = pi789 & ~n23161;
  assign n23170 = ~n23167 & n23169;
  assign n23171 = ~n23161 & n23168;
  assign n23172 = ~pi789 & n23155;
  assign n23173 = n59242 & ~n23172;
  assign n23174 = ~n59829 & n23173;
  assign n23175 = ~pi626 & ~n23011;
  assign n23176 = pi626 & ~n22874;
  assign n23177 = n7760 & ~n23176;
  assign n23178 = ~n23175 & n23177;
  assign n23179 = n7984 & n59820;
  assign n23180 = pi626 & ~n23011;
  assign n23181 = ~pi626 & ~n22874;
  assign n23182 = n7759 & ~n23181;
  assign n23183 = ~n23180 & n23182;
  assign n23184 = ~n23179 & ~n23183;
  assign n23185 = ~n23178 & ~n23179;
  assign n23186 = ~n23183 & n23185;
  assign n23187 = ~n23178 & n23184;
  assign n23188 = pi788 & ~n59830;
  assign n23189 = ~n59357 & ~n23188;
  assign n23190 = ~n23174 & n23189;
  assign n23191 = ~n23058 & ~n23190;
  assign n23192 = ~n8108 & ~n23191;
  assign n23193 = ~n23052 & ~n23192;
  assign n23194 = ~n59825 & n23193;
  assign n23195 = ~n23039 & ~n23194;
  assign n23196 = n58992 & ~n23195;
  assign n23197 = ~pi193 & ~n58992;
  assign n23198 = ~pi832 & ~n23197;
  assign n23199 = ~n23196 & n23198;
  assign po350 = ~n22873 & ~n23199;
  assign n23201 = ~pi194 & ~n7560;
  assign n23202 = n7762 & ~n23201;
  assign n23203 = n59231 & ~n23201;
  assign n23204 = pi194 & ~n13394;
  assign n23205 = ~pi194 & n13397;
  assign n23206 = pi730 & ~n23205;
  assign n23207 = ~pi194 & ~n7553;
  assign n23208 = ~pi730 & n23207;
  assign n23209 = n59132 & ~n23208;
  assign n23210 = ~n23206 & n23209;
  assign n23211 = ~n23204 & ~n23210;
  assign n23212 = ~pi778 & ~n23211;
  assign n23213 = pi625 & n23211;
  assign n23214 = ~pi625 & n23201;
  assign n23215 = pi1153 & ~n23214;
  assign n23216 = ~n23213 & n23215;
  assign n23217 = ~pi625 & n23211;
  assign n23218 = pi625 & n23201;
  assign n23219 = ~pi1153 & ~n23218;
  assign n23220 = ~n23217 & n23219;
  assign n23221 = ~n23216 & ~n23220;
  assign n23222 = pi778 & ~n23221;
  assign n23223 = ~n23212 & ~n23222;
  assign n23224 = ~n59229 & n23223;
  assign n23225 = n59229 & n23201;
  assign n23226 = n59229 & ~n23201;
  assign n23227 = ~n59229 & ~n23223;
  assign n23228 = ~n23226 & ~n23227;
  assign n23229 = ~n23224 & ~n23225;
  assign n23230 = ~n59231 & ~n59831;
  assign n23231 = ~n59231 & n59831;
  assign n23232 = n59231 & n23201;
  assign n23233 = ~n23231 & ~n23232;
  assign n23234 = ~n23203 & ~n23230;
  assign n23235 = ~n7716 & ~n59832;
  assign n23236 = n7716 & n23201;
  assign n23237 = n7716 & ~n23201;
  assign n23238 = ~n7716 & n59832;
  assign n23239 = ~n23237 & ~n23238;
  assign n23240 = ~n23235 & ~n23236;
  assign n23241 = ~n7762 & ~n59833;
  assign n23242 = ~n7762 & n59833;
  assign n23243 = n7762 & n23201;
  assign n23244 = ~n23242 & ~n23243;
  assign n23245 = ~n23202 & ~n23241;
  assign n23246 = pi628 & ~n59834;
  assign n23247 = ~pi628 & n23201;
  assign n23248 = pi1156 & ~n23247;
  assign n23249 = ~n23246 & n23248;
  assign n23250 = ~pi628 & ~n59834;
  assign n23251 = pi628 & n23201;
  assign n23252 = ~pi1156 & ~n23251;
  assign n23253 = ~n23250 & n23252;
  assign n23254 = pi628 & ~n23201;
  assign n23255 = ~pi628 & n59834;
  assign n23256 = ~n23254 & ~n23255;
  assign n23257 = ~pi1156 & n23256;
  assign n23258 = ~pi628 & ~n23201;
  assign n23259 = pi628 & n59834;
  assign n23260 = ~n23258 & ~n23259;
  assign n23261 = pi1156 & n23260;
  assign n23262 = ~n23257 & ~n23261;
  assign n23263 = ~n23249 & ~n23253;
  assign n23264 = pi792 & ~n59835;
  assign n23265 = ~pi792 & ~n59834;
  assign n23266 = ~pi792 & n59834;
  assign n23267 = pi792 & n59835;
  assign n23268 = ~n23266 & ~n23267;
  assign n23269 = ~n23264 & ~n23265;
  assign n23270 = pi647 & n59836;
  assign n23271 = ~pi647 & n23201;
  assign n23272 = ~n23270 & ~n23271;
  assign n23273 = n7832 & n23272;
  assign n23274 = ~pi647 & n59836;
  assign n23275 = pi647 & n23201;
  assign n23276 = ~n23274 & ~n23275;
  assign n23277 = n7833 & n23276;
  assign n23278 = pi194 & ~n59132;
  assign n23279 = ~pi194 & n9787;
  assign n23280 = pi194 & n13474;
  assign n23281 = ~n23279 & ~n23280;
  assign n23282 = pi748 & ~n23281;
  assign n23283 = ~pi748 & ~n23207;
  assign n23284 = ~n23282 & ~n23283;
  assign n23285 = n59132 & ~n23284;
  assign n23286 = ~n23278 & ~n23285;
  assign n23287 = ~n7597 & ~n23286;
  assign n23288 = n7597 & ~n23201;
  assign n23289 = ~n23287 & ~n23288;
  assign n23290 = ~pi785 & ~n23289;
  assign n23291 = ~n7598 & ~n23201;
  assign n23292 = pi609 & n23287;
  assign n23293 = ~n23291 & ~n23292;
  assign n23294 = pi1155 & ~n23293;
  assign n23295 = ~n7610 & ~n23201;
  assign n23296 = ~pi609 & n23287;
  assign n23297 = ~n23295 & ~n23296;
  assign n23298 = ~pi1155 & ~n23297;
  assign n23299 = ~n23294 & ~n23298;
  assign n23300 = pi785 & ~n23299;
  assign n23301 = ~n23290 & ~n23300;
  assign n23302 = ~pi781 & ~n23301;
  assign n23303 = pi618 & n23301;
  assign n23304 = ~pi618 & n23201;
  assign n23305 = pi1154 & ~n23304;
  assign n23306 = ~n23303 & n23305;
  assign n23307 = ~pi618 & n23301;
  assign n23308 = pi618 & n23201;
  assign n23309 = ~pi1154 & ~n23308;
  assign n23310 = ~n23307 & n23309;
  assign n23311 = ~n23306 & ~n23310;
  assign n23312 = pi781 & ~n23311;
  assign n23313 = ~n23302 & ~n23312;
  assign n23314 = ~pi789 & ~n23313;
  assign n23315 = ~pi619 & n23313;
  assign n23316 = pi619 & n23201;
  assign n23317 = ~pi1159 & ~n23316;
  assign n23318 = ~n23315 & n23317;
  assign n23319 = pi619 & n23313;
  assign n23320 = ~pi619 & n23201;
  assign n23321 = pi1159 & ~n23320;
  assign n23322 = ~n23319 & n23321;
  assign n23323 = ~n23318 & ~n23322;
  assign n23324 = pi789 & ~n23323;
  assign n23325 = ~n23314 & ~n23324;
  assign n23326 = ~n8054 & n23325;
  assign n23327 = n8054 & n23201;
  assign n23328 = ~n23326 & ~n23327;
  assign n23329 = ~n7793 & ~n23328;
  assign n23330 = n7793 & n23201;
  assign n23331 = ~n23329 & ~n23330;
  assign n23332 = ~n7872 & n23331;
  assign n23333 = ~n23277 & ~n23332;
  assign n23334 = ~n23273 & n23333;
  assign n23335 = pi787 & ~n23334;
  assign n23336 = n12139 & n23325;
  assign n23337 = ~pi641 & ~n59833;
  assign n23338 = pi641 & ~n23201;
  assign n23339 = n7912 & ~n23338;
  assign n23340 = ~n23337 & n23339;
  assign n23341 = pi641 & ~n59833;
  assign n23342 = ~pi641 & ~n23201;
  assign n23343 = n7911 & ~n23342;
  assign n23344 = ~n23341 & n23343;
  assign n23345 = ~n23340 & ~n23344;
  assign n23346 = ~n23336 & n23345;
  assign n23347 = pi788 & ~n23346;
  assign n23348 = pi619 & ~n59832;
  assign n23349 = ~pi1159 & ~n23348;
  assign n23350 = ~pi648 & ~n23322;
  assign n23351 = ~n23349 & n23350;
  assign n23352 = ~pi619 & ~n59832;
  assign n23353 = pi1159 & ~n23352;
  assign n23354 = pi648 & ~n23318;
  assign n23355 = ~n23353 & n23354;
  assign n23356 = ~n23351 & ~n23355;
  assign n23357 = pi789 & ~n23356;
  assign n23358 = pi618 & n59831;
  assign n23359 = ~pi1154 & ~n23358;
  assign n23360 = ~pi627 & ~n23306;
  assign n23361 = ~n23359 & n23360;
  assign n23362 = ~pi730 & n23284;
  assign n23363 = ~pi194 & n9797;
  assign n23364 = pi194 & ~n13579;
  assign n23365 = ~pi748 & ~n23364;
  assign n23366 = ~n23363 & n23365;
  assign n23367 = pi194 & n9811;
  assign n23368 = ~pi194 & ~n59320;
  assign n23369 = pi748 & ~n23368;
  assign n23370 = ~n23367 & n23369;
  assign n23371 = pi730 & ~n23370;
  assign n23372 = pi194 & ~n9811;
  assign n23373 = ~pi194 & n59320;
  assign n23374 = pi748 & ~n23373;
  assign n23375 = ~n23372 & n23374;
  assign n23376 = ~pi194 & ~n9797;
  assign n23377 = pi194 & n13579;
  assign n23378 = ~pi748 & ~n23377;
  assign n23379 = ~n23376 & n23378;
  assign n23380 = ~n23375 & ~n23379;
  assign n23381 = pi730 & ~n23380;
  assign n23382 = ~n23366 & n23371;
  assign n23383 = n59132 & ~n59837;
  assign n23384 = n59132 & ~n23362;
  assign n23385 = ~n59837 & n23384;
  assign n23386 = ~n23362 & n23383;
  assign n23387 = ~n23278 & ~n59838;
  assign n23388 = ~pi625 & n23387;
  assign n23389 = pi625 & n23286;
  assign n23390 = ~pi1153 & ~n23389;
  assign n23391 = ~n23388 & n23390;
  assign n23392 = ~pi608 & ~n23216;
  assign n23393 = ~n23391 & n23392;
  assign n23394 = pi625 & n23387;
  assign n23395 = ~pi625 & n23286;
  assign n23396 = pi1153 & ~n23395;
  assign n23397 = ~n23394 & n23396;
  assign n23398 = pi608 & ~n23220;
  assign n23399 = ~n23397 & n23398;
  assign n23400 = ~n23393 & ~n23399;
  assign n23401 = pi778 & ~n23400;
  assign n23402 = ~pi778 & n23387;
  assign n23403 = ~pi778 & ~n23387;
  assign n23404 = pi778 & ~n23399;
  assign n23405 = ~n23393 & n23404;
  assign n23406 = ~n23403 & ~n23405;
  assign n23407 = ~n23401 & ~n23402;
  assign n23408 = ~pi609 & n59839;
  assign n23409 = pi609 & n23223;
  assign n23410 = ~pi1155 & ~n23409;
  assign n23411 = ~n23408 & n23410;
  assign n23412 = ~pi660 & ~n23294;
  assign n23413 = ~n23411 & n23412;
  assign n23414 = pi609 & n59839;
  assign n23415 = ~pi609 & n23223;
  assign n23416 = pi1155 & ~n23415;
  assign n23417 = ~n23414 & n23416;
  assign n23418 = pi660 & ~n23298;
  assign n23419 = ~n23417 & n23418;
  assign n23420 = ~n23413 & ~n23419;
  assign n23421 = pi785 & ~n23420;
  assign n23422 = ~pi785 & n59839;
  assign n23423 = ~n23421 & ~n23422;
  assign n23424 = pi618 & ~n23423;
  assign n23425 = ~pi618 & n59831;
  assign n23426 = pi1154 & ~n23425;
  assign n23427 = ~n23424 & n23426;
  assign n23428 = pi627 & ~n23310;
  assign n23429 = ~n23427 & n23428;
  assign n23430 = ~n23361 & ~n23429;
  assign n23431 = pi781 & ~n23430;
  assign n23432 = ~pi618 & n23360;
  assign n23433 = pi781 & ~n23432;
  assign n23434 = ~n23423 & ~n23433;
  assign n23435 = ~pi618 & ~n23423;
  assign n23436 = n23359 & ~n23435;
  assign n23437 = n23360 & ~n23436;
  assign n23438 = ~n23429 & ~n23437;
  assign n23439 = pi781 & ~n23438;
  assign n23440 = ~pi781 & ~n23423;
  assign n23441 = ~n23439 & ~n23440;
  assign n23442 = ~n23431 & ~n23434;
  assign n23443 = ~pi619 & n23350;
  assign n23444 = pi619 & n23354;
  assign n23445 = pi789 & ~n23444;
  assign n23446 = ~n23443 & n23445;
  assign n23447 = ~n59840 & ~n23446;
  assign n23448 = ~pi619 & ~n59840;
  assign n23449 = n23349 & ~n23448;
  assign n23450 = n23350 & ~n23449;
  assign n23451 = pi619 & ~n59840;
  assign n23452 = n23353 & ~n23451;
  assign n23453 = n23354 & ~n23452;
  assign n23454 = ~n23450 & ~n23453;
  assign n23455 = pi789 & ~n23454;
  assign n23456 = ~pi789 & ~n59840;
  assign n23457 = ~n23455 & ~n23456;
  assign n23458 = ~n23357 & ~n23447;
  assign n23459 = n59242 & ~n59841;
  assign n23460 = ~pi788 & n59841;
  assign n23461 = ~pi626 & n59841;
  assign n23462 = pi626 & ~n59833;
  assign n23463 = ~pi641 & ~n23462;
  assign n23464 = ~n23461 & n23463;
  assign n23465 = ~pi626 & ~n23325;
  assign n23466 = pi626 & ~n23201;
  assign n23467 = pi641 & ~n23466;
  assign n23468 = ~n23465 & n23467;
  assign n23469 = ~pi1158 & ~n23468;
  assign n23470 = ~n23464 & n23469;
  assign n23471 = pi626 & n59841;
  assign n23472 = ~pi626 & ~n59833;
  assign n23473 = pi641 & ~n23472;
  assign n23474 = ~n23471 & n23473;
  assign n23475 = pi626 & ~n23325;
  assign n23476 = ~pi626 & ~n23201;
  assign n23477 = ~pi641 & ~n23476;
  assign n23478 = ~n23475 & n23477;
  assign n23479 = pi1158 & ~n23478;
  assign n23480 = ~n23474 & n23479;
  assign n23481 = ~n23470 & ~n23480;
  assign n23482 = pi788 & ~n23481;
  assign n23483 = ~n23460 & ~n23482;
  assign n23484 = ~n23347 & ~n23459;
  assign n23485 = ~n11154 & n23328;
  assign n23486 = n7791 & ~n23256;
  assign n23487 = n7790 & ~n23260;
  assign n23488 = ~n23486 & ~n23487;
  assign n23489 = ~n23485 & n23488;
  assign n23490 = pi792 & ~n23489;
  assign n23491 = n59842 & ~n23490;
  assign n23492 = n59357 & n23489;
  assign n23493 = ~n8108 & ~n23492;
  assign n23494 = ~n23491 & n23493;
  assign n23495 = ~pi628 & n59842;
  assign n23496 = pi628 & ~n23328;
  assign n23497 = ~pi1156 & ~n23496;
  assign n23498 = ~n23495 & n23497;
  assign n23499 = ~pi629 & ~n23249;
  assign n23500 = ~n23498 & n23499;
  assign n23501 = pi628 & n59842;
  assign n23502 = ~pi628 & ~n23328;
  assign n23503 = pi1156 & ~n23502;
  assign n23504 = ~n23501 & n23503;
  assign n23505 = pi629 & ~n23253;
  assign n23506 = ~n23504 & n23505;
  assign n23507 = ~n23500 & ~n23506;
  assign n23508 = pi792 & ~n23507;
  assign n23509 = ~pi792 & n59842;
  assign n23510 = ~n23508 & ~n23509;
  assign n23511 = ~pi647 & ~n23510;
  assign n23512 = pi647 & ~n23331;
  assign n23513 = ~pi1157 & ~n23512;
  assign n23514 = ~n23511 & n23513;
  assign n23515 = pi1157 & ~n23271;
  assign n23516 = ~n23270 & n23515;
  assign n23517 = ~pi630 & ~n23516;
  assign n23518 = ~n23514 & n23517;
  assign n23519 = pi647 & ~n23510;
  assign n23520 = ~pi647 & ~n23331;
  assign n23521 = pi1157 & ~n23520;
  assign n23522 = ~n23519 & n23521;
  assign n23523 = ~pi1157 & ~n23275;
  assign n23524 = ~n23274 & n23523;
  assign n23525 = pi630 & ~n23524;
  assign n23526 = ~n23522 & n23525;
  assign n23527 = ~n23518 & ~n23526;
  assign n23528 = pi787 & ~n23527;
  assign n23529 = ~pi787 & ~n23510;
  assign n23530 = ~n23528 & ~n23529;
  assign n23531 = ~n23335 & ~n23494;
  assign n23532 = ~pi715 & ~pi1160;
  assign n23533 = ~pi644 & n23532;
  assign n23534 = pi715 & pi1160;
  assign n23535 = pi644 & n23534;
  assign n23536 = ~n23533 & ~n23535;
  assign n23537 = pi790 & n23536;
  assign n23538 = n59843 & ~n23537;
  assign n23539 = ~pi1157 & ~n23276;
  assign n23540 = pi1157 & ~n23272;
  assign n23541 = ~n23539 & ~n23540;
  assign n23542 = ~n23516 & ~n23524;
  assign n23543 = pi787 & ~n59844;
  assign n23544 = ~pi787 & n59836;
  assign n23545 = pi644 & n23532;
  assign n23546 = ~pi644 & n23534;
  assign n23547 = ~n23545 & ~n23546;
  assign n23548 = ~n23544 & ~n23547;
  assign n23549 = ~n23543 & n23548;
  assign n23550 = ~n7835 & ~n23331;
  assign n23551 = n7835 & n23201;
  assign n23552 = n7835 & ~n23201;
  assign n23553 = ~n7835 & n23331;
  assign n23554 = ~n23552 & ~n23553;
  assign n23555 = ~n23550 & ~n23551;
  assign n23556 = pi644 & n59845;
  assign n23557 = ~pi715 & pi1160;
  assign n23558 = ~pi644 & n23201;
  assign n23559 = n23557 & ~n23558;
  assign n23560 = ~n23556 & n23559;
  assign n23561 = ~pi644 & n59845;
  assign n23562 = pi715 & ~pi1160;
  assign n23563 = pi644 & n23201;
  assign n23564 = n23562 & ~n23563;
  assign n23565 = ~n23561 & n23564;
  assign n23566 = ~n23560 & ~n23565;
  assign n23567 = ~n23549 & n23566;
  assign n23568 = pi790 & ~n23567;
  assign n23569 = n58992 & ~n23568;
  assign n23570 = pi644 & ~n59843;
  assign n23571 = ~pi787 & ~n59836;
  assign n23572 = pi787 & n59844;
  assign n23573 = ~n23571 & ~n23572;
  assign n23574 = ~pi644 & n23573;
  assign n23575 = pi715 & ~n23574;
  assign n23576 = ~n23570 & n23575;
  assign n23577 = ~pi715 & ~n23558;
  assign n23578 = ~n23556 & n23577;
  assign n23579 = pi1160 & ~n23578;
  assign n23580 = ~n23576 & n23579;
  assign n23581 = ~pi644 & ~n59843;
  assign n23582 = pi644 & n23573;
  assign n23583 = ~pi715 & ~n23582;
  assign n23584 = ~n23581 & n23583;
  assign n23585 = pi715 & ~n23563;
  assign n23586 = ~n23561 & n23585;
  assign n23587 = ~pi1160 & ~n23586;
  assign n23588 = ~n23584 & n23587;
  assign n23589 = pi790 & ~n23588;
  assign n23590 = pi790 & ~n23580;
  assign n23591 = ~n23588 & n23590;
  assign n23592 = ~n23580 & n23589;
  assign n23593 = ~pi790 & n59843;
  assign n23594 = n58992 & ~n23593;
  assign n23595 = ~n59846 & n23594;
  assign n23596 = ~n23538 & n23569;
  assign n23597 = ~pi194 & ~n58992;
  assign n23598 = ~pi832 & ~n23597;
  assign n23599 = ~n59847 & n23598;
  assign n23600 = ~pi194 & ~n2794;
  assign n23601 = pi748 & n6822;
  assign n23602 = ~n23600 & ~n23601;
  assign n23603 = ~n7875 & ~n23602;
  assign n23604 = ~pi785 & ~n23603;
  assign n23605 = ~n7880 & ~n23602;
  assign n23606 = pi1155 & ~n23605;
  assign n23607 = ~n7883 & n23603;
  assign n23608 = ~pi1155 & ~n23607;
  assign n23609 = ~n23606 & ~n23608;
  assign n23610 = pi785 & ~n23609;
  assign n23611 = ~n23604 & ~n23610;
  assign n23612 = ~pi781 & ~n23611;
  assign n23613 = ~n7890 & n23611;
  assign n23614 = pi1154 & ~n23613;
  assign n23615 = ~n7893 & n23611;
  assign n23616 = ~pi1154 & ~n23615;
  assign n23617 = ~n23614 & ~n23616;
  assign n23618 = pi781 & ~n23617;
  assign n23619 = ~n23612 & ~n23618;
  assign n23620 = ~pi789 & ~n23619;
  assign n23621 = pi619 & n23619;
  assign n23622 = ~pi619 & n23600;
  assign n23623 = pi1159 & ~n23622;
  assign n23624 = ~n23621 & n23623;
  assign n23625 = ~pi619 & n23619;
  assign n23626 = pi619 & n23600;
  assign n23627 = ~pi1159 & ~n23626;
  assign n23628 = ~n23625 & n23627;
  assign n23629 = ~n23624 & ~n23628;
  assign n23630 = pi789 & ~n23629;
  assign n23631 = ~n23620 & ~n23630;
  assign n23632 = ~n8054 & ~n23631;
  assign n23633 = n8054 & ~n23600;
  assign n23634 = ~n8054 & n23631;
  assign n23635 = n8054 & n23600;
  assign n23636 = ~n23634 & ~n23635;
  assign n23637 = ~n23632 & ~n23633;
  assign n23638 = ~n7793 & ~n59848;
  assign n23639 = n7793 & n23600;
  assign n23640 = ~n7872 & ~n23639;
  assign n23641 = ~n23638 & ~n23639;
  assign n23642 = ~n7872 & n23641;
  assign n23643 = ~n23638 & n23640;
  assign n23644 = pi730 & n7055;
  assign n23645 = ~n23600 & ~n23644;
  assign n23646 = ~pi778 & n23645;
  assign n23647 = ~pi625 & n23644;
  assign n23648 = ~n23645 & ~n23647;
  assign n23649 = pi1153 & ~n23648;
  assign n23650 = ~pi1153 & ~n23600;
  assign n23651 = ~n23647 & n23650;
  assign n23652 = ~n23649 & ~n23651;
  assign n23653 = pi778 & ~n23652;
  assign n23654 = ~n23646 & ~n23653;
  assign n23655 = ~n7949 & n23654;
  assign n23656 = ~n7951 & n23655;
  assign n23657 = ~n7953 & n23656;
  assign n23658 = ~n7955 & n23657;
  assign n23659 = ~n7967 & n23658;
  assign n23660 = pi647 & ~n23659;
  assign n23661 = ~pi647 & ~n23600;
  assign n23662 = ~n23660 & ~n23661;
  assign n23663 = n7832 & ~n23662;
  assign n23664 = ~pi647 & n23659;
  assign n23665 = pi647 & n23600;
  assign n23666 = ~pi1157 & ~n23665;
  assign n23667 = ~n23664 & n23666;
  assign n23668 = pi630 & n23667;
  assign n23669 = ~n23663 & ~n23668;
  assign n23670 = ~n59849 & n23669;
  assign n23671 = pi787 & ~n23670;
  assign n23672 = ~pi626 & ~n23631;
  assign n23673 = pi626 & ~n23600;
  assign n23674 = n7760 & ~n23673;
  assign n23675 = ~n23672 & n23674;
  assign n23676 = n7984 & n23657;
  assign n23677 = pi626 & ~n23631;
  assign n23678 = ~pi626 & ~n23600;
  assign n23679 = n7759 & ~n23678;
  assign n23680 = ~n23677 & n23679;
  assign n23681 = ~n23676 & ~n23680;
  assign n23682 = ~n23675 & ~n23676;
  assign n23683 = ~n23680 & n23682;
  assign n23684 = ~n23675 & n23681;
  assign n23685 = pi788 & ~n59850;
  assign n23686 = ~n6701 & ~n23645;
  assign n23687 = pi625 & n23686;
  assign n23688 = n23602 & ~n23686;
  assign n23689 = ~n23687 & ~n23688;
  assign n23690 = n23650 & ~n23689;
  assign n23691 = ~pi608 & ~n23649;
  assign n23692 = ~n23690 & n23691;
  assign n23693 = pi1153 & n23602;
  assign n23694 = ~n23687 & n23693;
  assign n23695 = pi608 & ~n23651;
  assign n23696 = ~n23694 & n23695;
  assign n23697 = ~n23692 & ~n23696;
  assign n23698 = pi778 & ~n23697;
  assign n23699 = ~pi778 & ~n23688;
  assign n23700 = ~n23698 & ~n23699;
  assign n23701 = ~pi609 & ~n23700;
  assign n23702 = pi609 & n23654;
  assign n23703 = ~pi1155 & ~n23702;
  assign n23704 = ~n23701 & n23703;
  assign n23705 = ~pi660 & ~n23606;
  assign n23706 = ~n23704 & n23705;
  assign n23707 = pi609 & ~n23700;
  assign n23708 = ~pi609 & n23654;
  assign n23709 = pi1155 & ~n23708;
  assign n23710 = ~n23707 & n23709;
  assign n23711 = pi660 & ~n23608;
  assign n23712 = ~n23710 & n23711;
  assign n23713 = ~n23706 & ~n23712;
  assign n23714 = pi785 & ~n23713;
  assign n23715 = ~pi785 & ~n23700;
  assign n23716 = ~n23714 & ~n23715;
  assign n23717 = ~pi618 & ~n23716;
  assign n23718 = pi618 & n23655;
  assign n23719 = ~pi1154 & ~n23718;
  assign n23720 = ~n23717 & n23719;
  assign n23721 = ~pi627 & ~n23614;
  assign n23722 = ~n23720 & n23721;
  assign n23723 = pi618 & ~n23716;
  assign n23724 = ~pi618 & n23655;
  assign n23725 = pi1154 & ~n23724;
  assign n23726 = ~n23723 & n23725;
  assign n23727 = pi627 & ~n23616;
  assign n23728 = ~n23726 & n23727;
  assign n23729 = ~n23722 & ~n23728;
  assign n23730 = pi781 & ~n23729;
  assign n23731 = ~pi781 & ~n23716;
  assign n23732 = ~n23730 & ~n23731;
  assign n23733 = ~pi619 & ~n23732;
  assign n23734 = pi619 & n23656;
  assign n23735 = ~pi1159 & ~n23734;
  assign n23736 = ~n23733 & n23735;
  assign n23737 = ~pi648 & ~n23624;
  assign n23738 = ~n23736 & n23737;
  assign n23739 = pi619 & ~n23732;
  assign n23740 = ~pi619 & n23656;
  assign n23741 = pi1159 & ~n23740;
  assign n23742 = ~n23739 & n23741;
  assign n23743 = pi648 & ~n23628;
  assign n23744 = ~n23742 & n23743;
  assign n23745 = pi789 & ~n23744;
  assign n23746 = pi789 & ~n23738;
  assign n23747 = ~n23744 & n23746;
  assign n23748 = ~n23738 & n23745;
  assign n23749 = ~pi789 & n23732;
  assign n23750 = n59242 & ~n23749;
  assign n23751 = ~n59851 & n23750;
  assign n23752 = ~n23685 & ~n23751;
  assign n23753 = ~n59357 & ~n23752;
  assign n23754 = n7957 & ~n59848;
  assign n23755 = n8065 & n23658;
  assign n23756 = pi629 & ~n23755;
  assign n23757 = ~n23754 & n23756;
  assign n23758 = n7958 & ~n59848;
  assign n23759 = n8074 & n23658;
  assign n23760 = ~pi629 & ~n23759;
  assign n23761 = ~n23758 & n23760;
  assign n23762 = pi792 & ~n23761;
  assign n23763 = ~n23758 & ~n23759;
  assign n23764 = ~pi629 & ~n23763;
  assign n23765 = ~n23754 & ~n23755;
  assign n23766 = pi629 & ~n23765;
  assign n23767 = ~n23764 & ~n23766;
  assign n23768 = pi792 & ~n23767;
  assign n23769 = pi792 & ~n23757;
  assign n23770 = ~n23761 & n23769;
  assign n23771 = ~n23757 & n23762;
  assign n23772 = ~n8108 & ~n59852;
  assign n23773 = ~n23753 & n23772;
  assign n23774 = ~n23671 & ~n23773;
  assign n23775 = pi644 & n23774;
  assign n23776 = ~pi787 & ~n23659;
  assign n23777 = pi1157 & ~n23662;
  assign n23778 = ~n23667 & ~n23777;
  assign n23779 = pi787 & ~n23778;
  assign n23780 = ~n23776 & ~n23779;
  assign n23781 = ~pi644 & n23780;
  assign n23782 = pi715 & ~n23781;
  assign n23783 = ~n23775 & n23782;
  assign n23784 = ~n11491 & n23600;
  assign n23785 = ~n7835 & n23638;
  assign n23786 = ~n7835 & ~n23641;
  assign n23787 = n7835 & n23600;
  assign n23788 = ~n23786 & ~n23787;
  assign n23789 = ~n23784 & ~n23785;
  assign n23790 = pi644 & ~n59853;
  assign n23791 = ~pi644 & n23600;
  assign n23792 = ~pi715 & ~n23791;
  assign n23793 = ~n23790 & n23792;
  assign n23794 = pi1160 & ~n23793;
  assign n23795 = ~n23783 & n23794;
  assign n23796 = ~pi644 & n23774;
  assign n23797 = pi644 & n23780;
  assign n23798 = ~pi715 & ~n23797;
  assign n23799 = ~n23796 & n23798;
  assign n23800 = ~pi644 & ~n59853;
  assign n23801 = pi644 & n23600;
  assign n23802 = pi715 & ~n23801;
  assign n23803 = ~n23800 & n23802;
  assign n23804 = ~pi1160 & ~n23803;
  assign n23805 = ~n23799 & n23804;
  assign n23806 = ~n23795 & ~n23805;
  assign n23807 = pi790 & ~n23806;
  assign n23808 = ~pi790 & n23774;
  assign n23809 = pi832 & ~n23808;
  assign n23810 = ~n23807 & n23809;
  assign po351 = ~n23599 & ~n23810;
  assign n23812 = pi199 & ~n7560;
  assign n23813 = n7762 & ~n23812;
  assign n23814 = n59231 & ~n23812;
  assign n23815 = ~pi637 & ~n23812;
  assign n23816 = ~pi199 & ~n6863;
  assign n23817 = n10432 & ~n23816;
  assign n23818 = pi199 & ~n59220;
  assign n23819 = ~pi199 & ~n7537;
  assign n23820 = pi39 & ~n23819;
  assign n23821 = ~n23818 & n23820;
  assign n23822 = ~pi199 & n7345;
  assign n23823 = pi199 & ~n7308;
  assign n23824 = ~pi39 & ~n23823;
  assign n23825 = ~n23822 & n23824;
  assign n23826 = ~pi38 & ~n23825;
  assign n23827 = ~n23821 & n23826;
  assign n23828 = ~n23817 & ~n23827;
  assign n23829 = n59132 & ~n23828;
  assign n23830 = pi199 & ~n59132;
  assign n23831 = pi637 & ~n23830;
  assign n23832 = ~n23829 & n23831;
  assign n23833 = ~n23815 & ~n23832;
  assign n23834 = ~pi778 & n23833;
  assign n23835 = pi625 & ~n23833;
  assign n23836 = ~pi625 & ~n23812;
  assign n23837 = pi1153 & ~n23836;
  assign n23838 = ~n23835 & n23837;
  assign n23839 = ~pi625 & ~n23833;
  assign n23840 = pi625 & ~n23812;
  assign n23841 = ~pi1153 & ~n23840;
  assign n23842 = ~n23839 & n23841;
  assign n23843 = ~n23838 & ~n23842;
  assign n23844 = pi778 & ~n23843;
  assign n23845 = ~n23834 & ~n23844;
  assign n23846 = ~n59229 & ~n23845;
  assign n23847 = n59229 & n23812;
  assign n23848 = n59229 & ~n23812;
  assign n23849 = ~n59229 & n23845;
  assign n23850 = ~n23848 & ~n23849;
  assign n23851 = ~n23846 & ~n23847;
  assign n23852 = ~n59231 & ~n59854;
  assign n23853 = ~n59231 & n59854;
  assign n23854 = n59231 & n23812;
  assign n23855 = ~n23853 & ~n23854;
  assign n23856 = ~n23814 & ~n23852;
  assign n23857 = ~n7716 & ~n59855;
  assign n23858 = n7716 & n23812;
  assign n23859 = n7716 & ~n23812;
  assign n23860 = ~n7716 & n59855;
  assign n23861 = ~n23859 & ~n23860;
  assign n23862 = ~n23857 & ~n23858;
  assign n23863 = ~n7762 & ~n59856;
  assign n23864 = ~n7762 & n59856;
  assign n23865 = n7762 & n23812;
  assign n23866 = ~n23864 & ~n23865;
  assign n23867 = ~n23813 & ~n23863;
  assign n23868 = pi628 & n59857;
  assign n23869 = ~pi628 & ~n23812;
  assign n23870 = pi1156 & ~n23869;
  assign n23871 = ~n23868 & n23870;
  assign n23872 = ~pi628 & n59857;
  assign n23873 = pi628 & ~n23812;
  assign n23874 = ~pi1156 & ~n23873;
  assign n23875 = ~n23872 & n23874;
  assign n23876 = ~n23872 & ~n23873;
  assign n23877 = ~pi1156 & ~n23876;
  assign n23878 = pi628 & ~n59857;
  assign n23879 = ~pi628 & n23812;
  assign n23880 = ~n23878 & ~n23879;
  assign n23881 = pi1156 & n23880;
  assign n23882 = ~n23877 & ~n23881;
  assign n23883 = ~n23871 & ~n23875;
  assign n23884 = pi792 & ~n59858;
  assign n23885 = ~pi792 & n59857;
  assign n23886 = ~pi792 & ~n59857;
  assign n23887 = pi792 & n59858;
  assign n23888 = ~n23886 & ~n23887;
  assign n23889 = ~n23884 & ~n23885;
  assign n23890 = pi647 & ~n59859;
  assign n23891 = ~pi647 & n23812;
  assign n23892 = ~n23890 & ~n23891;
  assign n23893 = n7832 & ~n23892;
  assign n23894 = ~pi647 & n59859;
  assign n23895 = pi647 & ~n23812;
  assign n23896 = ~pi1157 & ~n23895;
  assign n23897 = ~n23894 & n23896;
  assign n23898 = pi630 & n23897;
  assign n23899 = ~pi617 & ~n23812;
  assign n23900 = ~pi199 & ~n6865;
  assign n23901 = n9786 & ~n23900;
  assign n23902 = pi199 & n59164;
  assign n23903 = ~pi199 & ~n6855;
  assign n23904 = ~pi38 & ~n23903;
  assign n23905 = ~n23902 & n23904;
  assign n23906 = ~n23901 & ~n23905;
  assign n23907 = n59132 & ~n23906;
  assign n23908 = pi617 & ~n23830;
  assign n23909 = ~n23907 & n23908;
  assign n23910 = ~n23899 & ~n23909;
  assign n23911 = ~n7597 & n23910;
  assign n23912 = n7597 & n23812;
  assign n23913 = ~n7597 & ~n23910;
  assign n23914 = n7597 & ~n23812;
  assign n23915 = ~n23913 & ~n23914;
  assign n23916 = ~n23911 & ~n23912;
  assign n23917 = ~pi785 & n59860;
  assign n23918 = pi609 & ~n59860;
  assign n23919 = ~pi609 & ~n23812;
  assign n23920 = pi1155 & ~n23919;
  assign n23921 = ~n23918 & n23920;
  assign n23922 = ~pi609 & ~n59860;
  assign n23923 = pi609 & ~n23812;
  assign n23924 = ~pi1155 & ~n23923;
  assign n23925 = ~n23922 & n23924;
  assign n23926 = ~n23921 & ~n23925;
  assign n23927 = pi785 & ~n23926;
  assign n23928 = ~n23917 & ~n23927;
  assign n23929 = ~pi781 & ~n23928;
  assign n23930 = pi618 & n23928;
  assign n23931 = ~pi618 & ~n23812;
  assign n23932 = pi1154 & ~n23931;
  assign n23933 = ~n23930 & n23932;
  assign n23934 = ~pi618 & n23928;
  assign n23935 = pi618 & ~n23812;
  assign n23936 = ~pi1154 & ~n23935;
  assign n23937 = ~n23934 & n23936;
  assign n23938 = ~n23933 & ~n23937;
  assign n23939 = pi781 & ~n23938;
  assign n23940 = ~n23929 & ~n23939;
  assign n23941 = ~pi789 & ~n23940;
  assign n23942 = ~pi619 & n23940;
  assign n23943 = pi619 & ~n23812;
  assign n23944 = ~pi1159 & ~n23943;
  assign n23945 = ~n23942 & n23944;
  assign n23946 = pi619 & n23940;
  assign n23947 = ~pi619 & ~n23812;
  assign n23948 = pi1159 & ~n23947;
  assign n23949 = ~n23946 & n23948;
  assign n23950 = ~n23945 & ~n23949;
  assign n23951 = pi789 & ~n23950;
  assign n23952 = ~n23941 & ~n23951;
  assign n23953 = ~n8054 & ~n23952;
  assign n23954 = n8054 & n23812;
  assign n23955 = ~n23953 & ~n23954;
  assign n23956 = ~n7793 & ~n23955;
  assign n23957 = n7793 & n23812;
  assign n23958 = ~n23956 & ~n23957;
  assign n23959 = ~n7872 & ~n23958;
  assign n23960 = ~n23898 & ~n23959;
  assign n23961 = ~n23893 & n23960;
  assign n23962 = pi787 & ~n23961;
  assign n23963 = pi619 & n59855;
  assign n23964 = ~pi1159 & ~n23963;
  assign n23965 = ~pi648 & ~n23949;
  assign n23966 = ~n23964 & n23965;
  assign n23967 = ~pi619 & n59855;
  assign n23968 = pi1159 & ~n23967;
  assign n23969 = pi648 & ~n23945;
  assign n23970 = ~n23968 & n23969;
  assign n23971 = ~n23966 & ~n23970;
  assign n23972 = pi789 & ~n23971;
  assign n23973 = ~pi637 & n23910;
  assign n23974 = pi199 & n9796;
  assign n23975 = n59132 & ~n13579;
  assign n23976 = ~pi199 & ~n23975;
  assign n23977 = ~pi617 & ~n9795;
  assign n23978 = ~n23976 & n23977;
  assign n23979 = ~n23974 & n23977;
  assign n23980 = ~n23976 & n23979;
  assign n23981 = ~n23974 & n23978;
  assign n23982 = n59132 & n9811;
  assign n23983 = ~pi199 & ~n23982;
  assign n23984 = pi199 & n59320;
  assign n23985 = pi617 & ~n23984;
  assign n23986 = ~n23983 & n23985;
  assign n23987 = ~n23830 & ~n23986;
  assign n23988 = ~n59861 & n23987;
  assign n23989 = pi637 & ~n23988;
  assign n23990 = ~n23973 & ~n23989;
  assign n23991 = ~pi625 & n23990;
  assign n23992 = pi625 & ~n23910;
  assign n23993 = ~pi1153 & ~n23992;
  assign n23994 = ~n23991 & n23993;
  assign n23995 = ~pi608 & ~n23838;
  assign n23996 = ~n23994 & n23995;
  assign n23997 = pi625 & n23990;
  assign n23998 = ~pi625 & ~n23910;
  assign n23999 = pi1153 & ~n23998;
  assign n24000 = ~n23997 & n23999;
  assign n24001 = pi608 & ~n23842;
  assign n24002 = ~n24000 & n24001;
  assign n24003 = ~n23996 & ~n24002;
  assign n24004 = pi778 & ~n24003;
  assign n24005 = ~pi778 & n23990;
  assign n24006 = ~n24004 & ~n24005;
  assign n24007 = ~pi609 & ~n24006;
  assign n24008 = pi609 & n23845;
  assign n24009 = ~pi1155 & ~n24008;
  assign n24010 = ~n24007 & n24009;
  assign n24011 = ~pi660 & ~n23921;
  assign n24012 = ~n24010 & n24011;
  assign n24013 = pi609 & ~n24006;
  assign n24014 = ~pi609 & n23845;
  assign n24015 = pi1155 & ~n24014;
  assign n24016 = ~n24013 & n24015;
  assign n24017 = pi660 & ~n23925;
  assign n24018 = ~n24016 & n24017;
  assign n24019 = ~n24012 & ~n24018;
  assign n24020 = pi785 & ~n24019;
  assign n24021 = ~pi785 & ~n24006;
  assign n24022 = ~n24020 & ~n24021;
  assign n24023 = pi618 & ~n24022;
  assign n24024 = ~pi618 & ~n59854;
  assign n24025 = pi1154 & ~n24024;
  assign n24026 = ~n24023 & n24025;
  assign n24027 = pi627 & ~n23937;
  assign n24028 = ~n24026 & n24027;
  assign n24029 = ~pi618 & ~n24022;
  assign n24030 = pi618 & ~n59854;
  assign n24031 = ~pi1154 & ~n24030;
  assign n24032 = ~n24029 & n24031;
  assign n24033 = ~pi627 & ~n23933;
  assign n24034 = ~n24032 & n24033;
  assign n24035 = pi781 & ~n24034;
  assign n24036 = ~n24028 & n24035;
  assign n24037 = ~pi619 & n23965;
  assign n24038 = pi619 & n23969;
  assign n24039 = pi789 & ~n24038;
  assign n24040 = ~n24037 & n24039;
  assign n24041 = ~pi781 & n24022;
  assign n24042 = ~n24040 & ~n24041;
  assign n24043 = ~n24036 & n24042;
  assign n24044 = ~n24028 & ~n24034;
  assign n24045 = pi781 & ~n24044;
  assign n24046 = ~pi781 & ~n24022;
  assign n24047 = ~n24045 & ~n24046;
  assign n24048 = ~pi619 & ~n24047;
  assign n24049 = n23964 & ~n24048;
  assign n24050 = n23965 & ~n24049;
  assign n24051 = pi619 & ~n24047;
  assign n24052 = n23968 & ~n24051;
  assign n24053 = n23969 & ~n24052;
  assign n24054 = ~n24050 & ~n24053;
  assign n24055 = pi789 & ~n24054;
  assign n24056 = ~pi789 & ~n24047;
  assign n24057 = ~n24055 & ~n24056;
  assign n24058 = ~n23972 & ~n24043;
  assign n24059 = n59242 & ~n59862;
  assign n24060 = n12139 & n23952;
  assign n24061 = ~pi641 & n59856;
  assign n24062 = pi641 & n23812;
  assign n24063 = n7912 & ~n24062;
  assign n24064 = ~n24061 & n24063;
  assign n24065 = pi641 & n59856;
  assign n24066 = ~pi641 & n23812;
  assign n24067 = n7911 & ~n24066;
  assign n24068 = ~n24065 & n24067;
  assign n24069 = ~n24064 & ~n24068;
  assign n24070 = ~n24060 & n24069;
  assign n24071 = pi788 & ~n24070;
  assign n24072 = ~pi788 & n59862;
  assign n24073 = ~pi626 & n59862;
  assign n24074 = pi626 & n59856;
  assign n24075 = ~pi641 & ~n24074;
  assign n24076 = ~n24073 & n24075;
  assign n24077 = ~pi626 & ~n23952;
  assign n24078 = pi626 & n23812;
  assign n24079 = pi641 & ~n24078;
  assign n24080 = ~n24077 & n24079;
  assign n24081 = ~pi1158 & ~n24080;
  assign n24082 = ~n24076 & n24081;
  assign n24083 = pi626 & n59862;
  assign n24084 = ~pi626 & n59856;
  assign n24085 = pi641 & ~n24084;
  assign n24086 = ~n24083 & n24085;
  assign n24087 = pi626 & ~n23952;
  assign n24088 = ~pi626 & n23812;
  assign n24089 = ~pi641 & ~n24088;
  assign n24090 = ~n24087 & n24089;
  assign n24091 = pi1158 & ~n24090;
  assign n24092 = ~n24086 & n24091;
  assign n24093 = ~n24082 & ~n24092;
  assign n24094 = pi788 & ~n24093;
  assign n24095 = ~n24072 & ~n24094;
  assign n24096 = ~n24059 & ~n24071;
  assign n24097 = ~n11154 & ~n23955;
  assign n24098 = n7791 & n23876;
  assign n24099 = n7790 & ~n23880;
  assign n24100 = ~n24098 & ~n24099;
  assign n24101 = ~n24097 & n24100;
  assign n24102 = pi792 & ~n24101;
  assign n24103 = n59863 & ~n24102;
  assign n24104 = n59357 & n24101;
  assign n24105 = ~n8108 & ~n24104;
  assign n24106 = ~n24103 & n24105;
  assign n24107 = ~pi628 & n59863;
  assign n24108 = pi628 & n23955;
  assign n24109 = ~pi1156 & ~n24108;
  assign n24110 = ~n24107 & n24109;
  assign n24111 = ~pi629 & ~n23871;
  assign n24112 = ~n24110 & n24111;
  assign n24113 = pi628 & n59863;
  assign n24114 = ~pi628 & n23955;
  assign n24115 = pi1156 & ~n24114;
  assign n24116 = ~n24113 & n24115;
  assign n24117 = pi629 & ~n23875;
  assign n24118 = ~n24116 & n24117;
  assign n24119 = ~n24112 & ~n24118;
  assign n24120 = pi792 & ~n24119;
  assign n24121 = ~pi792 & n59863;
  assign n24122 = ~n24120 & ~n24121;
  assign n24123 = ~pi647 & ~n24122;
  assign n24124 = pi647 & n23958;
  assign n24125 = ~pi1157 & ~n24124;
  assign n24126 = ~n24123 & n24125;
  assign n24127 = pi647 & n59859;
  assign n24128 = ~pi647 & ~n23812;
  assign n24129 = pi1157 & ~n24128;
  assign n24130 = pi1157 & ~n23892;
  assign n24131 = ~n24127 & n24129;
  assign n24132 = ~pi630 & ~n59864;
  assign n24133 = ~n24126 & n24132;
  assign n24134 = pi647 & ~n24122;
  assign n24135 = ~pi647 & n23958;
  assign n24136 = pi1157 & ~n24135;
  assign n24137 = ~n24134 & n24136;
  assign n24138 = pi630 & ~n23897;
  assign n24139 = ~n24137 & n24138;
  assign n24140 = ~n24133 & ~n24139;
  assign n24141 = pi787 & ~n24140;
  assign n24142 = ~pi787 & ~n24122;
  assign n24143 = ~n24141 & ~n24142;
  assign n24144 = ~n23962 & ~n24106;
  assign n24145 = ~pi644 & ~n59865;
  assign n24146 = ~pi787 & ~n59859;
  assign n24147 = ~n23897 & ~n59864;
  assign n24148 = pi787 & ~n24147;
  assign n24149 = ~n24146 & ~n24148;
  assign n24150 = pi644 & n24149;
  assign n24151 = ~pi715 & ~n24150;
  assign n24152 = ~n24145 & n24151;
  assign n24153 = ~n7835 & ~n23958;
  assign n24154 = n7835 & n23812;
  assign n24155 = n7835 & ~n23812;
  assign n24156 = ~n7835 & n23958;
  assign n24157 = ~n24155 & ~n24156;
  assign n24158 = ~n24153 & ~n24154;
  assign n24159 = ~pi644 & ~n59866;
  assign n24160 = pi644 & ~n23812;
  assign n24161 = pi715 & ~n24160;
  assign n24162 = ~n24159 & n24161;
  assign n24163 = ~pi1160 & ~n24162;
  assign n24164 = ~n24152 & n24163;
  assign n24165 = pi644 & ~n59865;
  assign n24166 = ~pi644 & n24149;
  assign n24167 = pi715 & ~n24166;
  assign n24168 = ~n24165 & n24167;
  assign n24169 = pi644 & ~n59866;
  assign n24170 = ~pi644 & ~n23812;
  assign n24171 = ~pi715 & ~n24170;
  assign n24172 = ~n24169 & n24171;
  assign n24173 = pi1160 & ~n24172;
  assign n24174 = ~n24168 & n24173;
  assign n24175 = ~n24164 & ~n24174;
  assign n24176 = pi790 & ~n24175;
  assign n24177 = ~pi790 & ~n59865;
  assign n24178 = ~pi790 & n59865;
  assign n24179 = pi790 & ~n24164;
  assign n24180 = pi790 & ~n24174;
  assign n24181 = ~n24164 & n24180;
  assign n24182 = ~n24174 & n24179;
  assign n24183 = ~n24178 & ~n59867;
  assign n24184 = ~n24176 & ~n24177;
  assign n24185 = n58992 & n59868;
  assign n24186 = ~pi199 & ~n58992;
  assign n24187 = n58992 & ~n59868;
  assign n24188 = pi199 & ~n58992;
  assign n24189 = ~n24187 & ~n24188;
  assign n24190 = ~n24185 & ~n24186;
  assign n24191 = pi200 & ~n58992;
  assign n24192 = pi200 & ~n7560;
  assign n24193 = n59231 & ~n24192;
  assign n24194 = ~pi643 & ~n24192;
  assign n24195 = ~pi200 & ~n6863;
  assign n24196 = n10432 & ~n24195;
  assign n24197 = pi200 & ~n59219;
  assign n24198 = ~pi200 & n7511;
  assign n24199 = ~pi299 & ~n24198;
  assign n24200 = ~n24197 & n24199;
  assign n24201 = pi200 & ~n59216;
  assign n24202 = ~pi200 & n7535;
  assign n24203 = pi299 & ~n24202;
  assign n24204 = ~n24201 & n24203;
  assign n24205 = ~n24200 & ~n24204;
  assign n24206 = pi39 & ~n24205;
  assign n24207 = ~pi200 & ~n7345;
  assign n24208 = pi200 & n7308;
  assign n24209 = ~pi39 & ~n24208;
  assign n24210 = ~pi39 & ~n24207;
  assign n24211 = ~n24208 & n24210;
  assign n24212 = ~n24207 & n24209;
  assign n24213 = ~n24206 & ~n59870;
  assign n24214 = ~pi38 & ~n24213;
  assign n24215 = ~n24196 & ~n24214;
  assign n24216 = n59132 & ~n24215;
  assign n24217 = pi200 & ~n59132;
  assign n24218 = pi643 & ~n24217;
  assign n24219 = ~n24216 & n24218;
  assign n24220 = ~n24194 & ~n24219;
  assign n24221 = ~pi778 & n24220;
  assign n24222 = pi625 & ~n24220;
  assign n24223 = ~pi625 & ~n24192;
  assign n24224 = pi1153 & ~n24223;
  assign n24225 = ~n24222 & n24224;
  assign n24226 = ~pi625 & ~n24220;
  assign n24227 = pi625 & ~n24192;
  assign n24228 = ~pi1153 & ~n24227;
  assign n24229 = ~n24226 & n24228;
  assign n24230 = ~n24225 & ~n24229;
  assign n24231 = pi778 & ~n24230;
  assign n24232 = ~n24221 & ~n24231;
  assign n24233 = ~n59229 & ~n24232;
  assign n24234 = n59229 & n24192;
  assign n24235 = n59229 & ~n24192;
  assign n24236 = ~n59229 & n24232;
  assign n24237 = ~n24235 & ~n24236;
  assign n24238 = ~n24233 & ~n24234;
  assign n24239 = ~n59231 & ~n59871;
  assign n24240 = ~n59231 & n59871;
  assign n24241 = n59231 & n24192;
  assign n24242 = ~n24240 & ~n24241;
  assign n24243 = ~n24193 & ~n24239;
  assign n24244 = ~n7716 & ~n59872;
  assign n24245 = n7716 & n24192;
  assign n24246 = n7716 & ~n24192;
  assign n24247 = ~n7716 & n59872;
  assign n24248 = ~n24246 & ~n24247;
  assign n24249 = ~n24244 & ~n24245;
  assign n24250 = ~n7762 & n59873;
  assign n24251 = n7762 & n24192;
  assign n24252 = ~n24250 & ~n24251;
  assign n24253 = ~pi792 & ~n24252;
  assign n24254 = pi628 & n24252;
  assign n24255 = ~pi628 & ~n24192;
  assign n24256 = pi1156 & ~n24255;
  assign n24257 = ~n24254 & n24256;
  assign n24258 = ~pi628 & n24252;
  assign n24259 = pi628 & ~n24192;
  assign n24260 = ~pi1156 & ~n24259;
  assign n24261 = ~n24258 & n24260;
  assign n24262 = ~n24257 & ~n24261;
  assign n24263 = pi792 & ~n24262;
  assign n24264 = ~n24253 & ~n24263;
  assign n24265 = pi647 & ~n24264;
  assign n24266 = ~pi647 & n24192;
  assign n24267 = ~n24265 & ~n24266;
  assign n24268 = pi1157 & ~n24267;
  assign n24269 = ~pi647 & n24264;
  assign n24270 = pi647 & ~n24192;
  assign n24271 = ~pi1157 & ~n24270;
  assign n24272 = ~n24269 & n24271;
  assign n24273 = pi787 & ~n24272;
  assign n24274 = ~n24268 & n24273;
  assign n24275 = ~pi787 & n24264;
  assign n24276 = ~n23547 & ~n24275;
  assign n24277 = ~n24274 & n24276;
  assign n24278 = ~pi606 & ~n24192;
  assign n24279 = ~pi200 & ~n6865;
  assign n24280 = n9786 & ~n24279;
  assign n24281 = pi200 & n59164;
  assign n24282 = ~pi200 & ~n6855;
  assign n24283 = ~pi38 & ~n24282;
  assign n24284 = ~n24281 & n24283;
  assign n24285 = ~n24280 & ~n24284;
  assign n24286 = n59132 & ~n24285;
  assign n24287 = pi606 & ~n24217;
  assign n24288 = ~n24286 & n24287;
  assign n24289 = ~n24278 & ~n24288;
  assign n24290 = ~n7597 & n24289;
  assign n24291 = n7597 & n24192;
  assign n24292 = ~n7597 & ~n24289;
  assign n24293 = n7597 & ~n24192;
  assign n24294 = ~n24292 & ~n24293;
  assign n24295 = ~n24290 & ~n24291;
  assign n24296 = ~pi785 & n59874;
  assign n24297 = pi609 & ~n59874;
  assign n24298 = ~pi609 & ~n24192;
  assign n24299 = pi1155 & ~n24298;
  assign n24300 = ~n24297 & n24299;
  assign n24301 = ~pi609 & ~n59874;
  assign n24302 = pi609 & ~n24192;
  assign n24303 = ~pi1155 & ~n24302;
  assign n24304 = ~n24301 & n24303;
  assign n24305 = ~n24300 & ~n24304;
  assign n24306 = pi785 & ~n24305;
  assign n24307 = ~n24296 & ~n24306;
  assign n24308 = ~pi781 & ~n24307;
  assign n24309 = pi618 & n24307;
  assign n24310 = ~pi618 & ~n24192;
  assign n24311 = pi1154 & ~n24310;
  assign n24312 = ~n24309 & n24311;
  assign n24313 = ~pi618 & n24307;
  assign n24314 = pi618 & ~n24192;
  assign n24315 = ~pi1154 & ~n24314;
  assign n24316 = ~n24313 & n24315;
  assign n24317 = ~n24312 & ~n24316;
  assign n24318 = pi781 & ~n24317;
  assign n24319 = ~n24308 & ~n24318;
  assign n24320 = ~pi789 & ~n24319;
  assign n24321 = pi619 & n24319;
  assign n24322 = ~pi619 & ~n24192;
  assign n24323 = pi1159 & ~n24322;
  assign n24324 = ~n24321 & n24323;
  assign n24325 = ~pi619 & n24319;
  assign n24326 = pi619 & ~n24192;
  assign n24327 = ~pi1159 & ~n24326;
  assign n24328 = ~n24325 & n24327;
  assign n24329 = ~n24324 & ~n24328;
  assign n24330 = pi789 & ~n24329;
  assign n24331 = ~n24320 & ~n24330;
  assign n24332 = ~n8054 & ~n24331;
  assign n24333 = n8054 & n24192;
  assign n24334 = ~n24332 & ~n24333;
  assign n24335 = ~n7793 & ~n24334;
  assign n24336 = n7793 & n24192;
  assign n24337 = ~n24335 & ~n24336;
  assign n24338 = ~n7835 & ~n24337;
  assign n24339 = n7835 & n24192;
  assign n24340 = n7835 & ~n24192;
  assign n24341 = ~n7835 & n24337;
  assign n24342 = ~n24340 & ~n24341;
  assign n24343 = ~n24338 & ~n24339;
  assign n24344 = pi644 & ~n59875;
  assign n24345 = ~pi644 & ~n24192;
  assign n24346 = n23557 & ~n24345;
  assign n24347 = ~n24344 & n24346;
  assign n24348 = ~pi644 & ~n59875;
  assign n24349 = pi644 & ~n24192;
  assign n24350 = n23562 & ~n24349;
  assign n24351 = ~n24348 & n24350;
  assign n24352 = ~n24347 & ~n24351;
  assign n24353 = ~n24277 & n24352;
  assign n24354 = pi790 & ~n24353;
  assign n24355 = n7832 & ~n24267;
  assign n24356 = ~n7872 & ~n24337;
  assign n24357 = pi630 & n24272;
  assign n24358 = ~n24356 & ~n24357;
  assign n24359 = ~n24355 & ~n24356;
  assign n24360 = ~n24357 & n24359;
  assign n24361 = ~n24355 & n24358;
  assign n24362 = pi787 & ~n59876;
  assign n24363 = ~n11154 & ~n24334;
  assign n24364 = ~pi629 & n24257;
  assign n24365 = pi629 & n24261;
  assign n24366 = ~n24364 & ~n24365;
  assign n24367 = ~n24363 & n24366;
  assign n24368 = pi792 & ~n24367;
  assign n24369 = ~pi643 & n24289;
  assign n24370 = ~n6914 & ~n7547;
  assign n24371 = n24196 & ~n24370;
  assign n24372 = pi200 & ~n8213;
  assign n24373 = ~pi200 & ~n8217;
  assign n24374 = ~pi38 & ~n24373;
  assign n24375 = ~n24372 & n24374;
  assign n24376 = ~n24371 & ~n24375;
  assign n24377 = ~pi606 & n59132;
  assign n24378 = ~n24376 & n24377;
  assign n24379 = pi200 & ~n13062;
  assign n24380 = ~pi200 & ~n59317;
  assign n24381 = ~pi38 & ~n24380;
  assign n24382 = ~n24379 & n24381;
  assign n24383 = ~n9805 & ~n9810;
  assign n24384 = ~pi200 & ~n24383;
  assign n24385 = pi38 & ~pi39;
  assign n24386 = pi200 & n24385;
  assign n24387 = pi38 & pi200;
  assign n24388 = n59319 & n24387;
  assign n24389 = n7222 & n24386;
  assign n24390 = pi606 & n59132;
  assign n24391 = ~n59877 & n24390;
  assign n24392 = ~n24384 & n24391;
  assign n24393 = ~n24382 & n24392;
  assign n24394 = ~n24217 & ~n24393;
  assign n24395 = ~n24378 & n24394;
  assign n24396 = pi643 & ~n24395;
  assign n24397 = ~n24369 & ~n24396;
  assign n24398 = ~pi625 & n24397;
  assign n24399 = pi625 & ~n24289;
  assign n24400 = ~pi1153 & ~n24399;
  assign n24401 = ~n24398 & n24400;
  assign n24402 = ~pi608 & ~n24225;
  assign n24403 = ~n24401 & n24402;
  assign n24404 = pi625 & n24397;
  assign n24405 = ~pi625 & ~n24289;
  assign n24406 = pi1153 & ~n24405;
  assign n24407 = ~n24404 & n24406;
  assign n24408 = pi608 & ~n24229;
  assign n24409 = ~n24407 & n24408;
  assign n24410 = ~n24403 & ~n24409;
  assign n24411 = pi778 & ~n24410;
  assign n24412 = ~pi778 & n24397;
  assign n24413 = ~n24411 & ~n24412;
  assign n24414 = ~pi609 & ~n24413;
  assign n24415 = pi609 & n24232;
  assign n24416 = ~pi1155 & ~n24415;
  assign n24417 = ~n24414 & n24416;
  assign n24418 = ~pi660 & ~n24300;
  assign n24419 = ~n24417 & n24418;
  assign n24420 = pi609 & ~n24413;
  assign n24421 = ~pi609 & n24232;
  assign n24422 = pi1155 & ~n24421;
  assign n24423 = ~n24420 & n24422;
  assign n24424 = pi660 & ~n24304;
  assign n24425 = ~n24423 & n24424;
  assign n24426 = ~n24419 & ~n24425;
  assign n24427 = pi785 & ~n24426;
  assign n24428 = ~pi785 & ~n24413;
  assign n24429 = ~n24427 & ~n24428;
  assign n24430 = ~pi618 & ~n24429;
  assign n24431 = pi618 & ~n59871;
  assign n24432 = ~pi1154 & ~n24431;
  assign n24433 = ~n24430 & n24432;
  assign n24434 = ~pi627 & ~n24312;
  assign n24435 = ~n24433 & n24434;
  assign n24436 = pi618 & ~n24429;
  assign n24437 = ~pi618 & ~n59871;
  assign n24438 = pi1154 & ~n24437;
  assign n24439 = ~n24436 & n24438;
  assign n24440 = pi627 & ~n24316;
  assign n24441 = ~n24439 & n24440;
  assign n24442 = ~n24435 & ~n24441;
  assign n24443 = pi781 & ~n24442;
  assign n24444 = ~pi781 & ~n24429;
  assign n24445 = ~n24443 & ~n24444;
  assign n24446 = ~pi619 & ~n24445;
  assign n24447 = pi619 & n59872;
  assign n24448 = ~pi1159 & ~n24447;
  assign n24449 = ~n24446 & n24448;
  assign n24450 = ~pi648 & ~n24324;
  assign n24451 = ~n24449 & n24450;
  assign n24452 = pi619 & ~n24445;
  assign n24453 = ~pi619 & n59872;
  assign n24454 = pi1159 & ~n24453;
  assign n24455 = ~n24452 & n24454;
  assign n24456 = pi648 & ~n24328;
  assign n24457 = ~n24455 & n24456;
  assign n24458 = pi789 & ~n24457;
  assign n24459 = pi789 & ~n24451;
  assign n24460 = ~n24457 & n24459;
  assign n24461 = ~n24451 & n24458;
  assign n24462 = ~pi789 & n24445;
  assign n24463 = n59242 & ~n24462;
  assign n24464 = ~n59878 & n24463;
  assign n24465 = ~pi626 & ~n24331;
  assign n24466 = pi626 & n24192;
  assign n24467 = n7760 & ~n24466;
  assign n24468 = ~n24465 & n24467;
  assign n24469 = n7984 & ~n59873;
  assign n24470 = pi626 & ~n24331;
  assign n24471 = ~pi626 & n24192;
  assign n24472 = n7759 & ~n24471;
  assign n24473 = ~n24470 & n24472;
  assign n24474 = ~n24469 & ~n24473;
  assign n24475 = ~n24468 & ~n24469;
  assign n24476 = ~n24473 & n24475;
  assign n24477 = ~n24468 & n24474;
  assign n24478 = pi788 & ~n59879;
  assign n24479 = ~n59357 & ~n24478;
  assign n24480 = ~n24464 & n24479;
  assign n24481 = ~n24368 & ~n24480;
  assign n24482 = ~n8108 & ~n24481;
  assign n24483 = ~n24362 & ~n24482;
  assign n24484 = ~n23537 & ~n24483;
  assign n24485 = ~pi644 & n24483;
  assign n24486 = ~pi787 & ~n24264;
  assign n24487 = ~n24268 & ~n24272;
  assign n24488 = pi787 & ~n24487;
  assign n24489 = ~n24486 & ~n24488;
  assign n24490 = pi644 & n24489;
  assign n24491 = ~pi715 & ~n24490;
  assign n24492 = ~n24485 & n24491;
  assign n24493 = pi715 & ~n24349;
  assign n24494 = ~n24348 & n24493;
  assign n24495 = ~pi1160 & ~n24494;
  assign n24496 = ~n24492 & n24495;
  assign n24497 = pi644 & n24483;
  assign n24498 = ~pi644 & n24489;
  assign n24499 = pi715 & ~n24498;
  assign n24500 = ~n24497 & n24499;
  assign n24501 = ~pi715 & ~n24345;
  assign n24502 = ~n24344 & n24501;
  assign n24503 = pi1160 & ~n24502;
  assign n24504 = ~n24500 & n24503;
  assign n24505 = ~n24496 & ~n24504;
  assign n24506 = pi790 & ~n24505;
  assign n24507 = ~pi790 & n24483;
  assign n24508 = ~n24506 & ~n24507;
  assign n24509 = ~n24354 & ~n24484;
  assign n24510 = n58992 & n59880;
  assign n24511 = n58992 & ~n59880;
  assign n24512 = ~pi200 & ~n58992;
  assign n24513 = ~n24511 & ~n24512;
  assign n24514 = ~n24191 & ~n24510;
  assign n24515 = ~n59304 & n13394;
  assign n24516 = n9554 & n24515;
  assign n24517 = ~n7716 & n24516;
  assign n24518 = ~n7762 & n24517;
  assign n24519 = n9652 & n24515;
  assign n24520 = ~n59240 & n59882;
  assign n24521 = pi207 & ~n24520;
  assign n24522 = ~n7560 & n7762;
  assign n24523 = ~n7560 & n59231;
  assign n24524 = n59132 & n13397;
  assign n24525 = ~pi778 & ~n24524;
  assign n24526 = ~pi625 & ~n7560;
  assign n24527 = pi625 & ~n24524;
  assign n24528 = ~n24526 & ~n24527;
  assign n24529 = pi1153 & ~n24528;
  assign n24530 = pi625 & ~n7560;
  assign n24531 = ~pi625 & ~n24524;
  assign n24532 = ~n24530 & ~n24531;
  assign n24533 = ~pi1153 & ~n24532;
  assign n24534 = ~n24529 & ~n24533;
  assign n24535 = pi778 & ~n24534;
  assign n24536 = ~n24525 & ~n24535;
  assign n24537 = ~n59229 & n24536;
  assign n24538 = n7560 & n59229;
  assign n24539 = ~n7560 & n59229;
  assign n24540 = ~n59229 & ~n24536;
  assign n24541 = ~n24539 & ~n24540;
  assign n24542 = ~n24537 & ~n24538;
  assign n24543 = ~n59231 & ~n59883;
  assign n24544 = ~n59231 & n59883;
  assign n24545 = n7560 & n59231;
  assign n24546 = ~n24544 & ~n24545;
  assign n24547 = ~n24523 & ~n24543;
  assign n24548 = ~n7716 & ~n59884;
  assign n24549 = n7560 & n7716;
  assign n24550 = ~n7560 & n7716;
  assign n24551 = ~n7716 & n59884;
  assign n24552 = ~n24550 & ~n24551;
  assign n24553 = ~n24548 & ~n24549;
  assign n24554 = ~n7762 & ~n59885;
  assign n24555 = ~n7762 & n59885;
  assign n24556 = n7560 & n7762;
  assign n24557 = ~n24555 & ~n24556;
  assign n24558 = ~n24522 & ~n24554;
  assign n24559 = ~n59240 & n59886;
  assign n24560 = ~n7560 & n59240;
  assign n24561 = ~n59240 & ~n59886;
  assign n24562 = n7560 & n59240;
  assign n24563 = ~n24561 & ~n24562;
  assign n24564 = ~n24559 & ~n24560;
  assign n24565 = ~pi207 & ~n59887;
  assign n24566 = ~n24521 & ~n24565;
  assign n24567 = pi710 & ~n24566;
  assign n24568 = ~pi207 & ~n7560;
  assign n24569 = ~pi710 & ~n24568;
  assign n24570 = ~n24567 & ~n24569;
  assign n24571 = ~pi647 & n24570;
  assign n24572 = pi647 & n24568;
  assign n24573 = ~pi1157 & ~n24572;
  assign n24574 = ~n24571 & n24573;
  assign n24575 = pi630 & n24574;
  assign n24576 = pi647 & n24570;
  assign n24577 = ~pi647 & n24568;
  assign n24578 = pi1157 & ~n24577;
  assign n24579 = ~n24576 & n24578;
  assign n24580 = ~pi630 & n24579;
  assign n24581 = ~n7560 & n7597;
  assign n24582 = n59132 & n9787;
  assign n24583 = ~n7597 & ~n24582;
  assign n24584 = ~n24581 & ~n24583;
  assign n24585 = ~pi785 & ~n24584;
  assign n24586 = ~n7560 & ~n7610;
  assign n24587 = ~pi609 & n24583;
  assign n24588 = ~n24586 & ~n24587;
  assign n24589 = ~pi1155 & ~n24588;
  assign n24590 = ~n7560 & ~n7598;
  assign n24591 = pi609 & n24583;
  assign n24592 = ~n24590 & ~n24591;
  assign n24593 = pi1155 & ~n24592;
  assign n24594 = ~n24589 & ~n24593;
  assign n24595 = pi785 & ~n24594;
  assign n24596 = ~n24585 & ~n24595;
  assign n24597 = ~pi781 & ~n24596;
  assign n24598 = ~pi618 & n24596;
  assign n24599 = pi618 & n7560;
  assign n24600 = ~pi1154 & ~n24599;
  assign n24601 = ~n24598 & n24600;
  assign n24602 = pi618 & n24596;
  assign n24603 = ~pi618 & n7560;
  assign n24604 = pi1154 & ~n24603;
  assign n24605 = ~n24602 & n24604;
  assign n24606 = ~n24601 & ~n24605;
  assign n24607 = pi781 & ~n24606;
  assign n24608 = ~n24597 & ~n24607;
  assign n24609 = ~pi789 & ~n24608;
  assign n24610 = ~pi619 & n24608;
  assign n24611 = pi619 & n7560;
  assign n24612 = ~pi1159 & ~n24611;
  assign n24613 = ~n24610 & n24612;
  assign n24614 = pi619 & n24608;
  assign n24615 = ~pi619 & n7560;
  assign n24616 = pi1159 & ~n24615;
  assign n24617 = ~n24614 & n24616;
  assign n24618 = ~n24613 & ~n24617;
  assign n24619 = pi789 & ~n24618;
  assign n24620 = ~n24609 & ~n24619;
  assign n24621 = ~n8054 & n24620;
  assign n24622 = n7560 & n8054;
  assign n24623 = ~n24621 & ~n24622;
  assign n24624 = ~n7793 & ~n24623;
  assign n24625 = n7560 & n7793;
  assign n24626 = ~n24624 & ~n24625;
  assign n24627 = ~pi207 & ~n24626;
  assign n24628 = n59132 & ~n13474;
  assign n24629 = ~n7597 & n24628;
  assign n24630 = ~n59346 & n24629;
  assign n24631 = ~n59347 & n24630;
  assign n24632 = ~n10741 & n24631;
  assign n24633 = ~n8054 & n24632;
  assign n24634 = ~n7793 & n24633;
  assign n24635 = pi207 & ~n24634;
  assign n24636 = pi623 & ~n24635;
  assign n24637 = ~pi207 & n24626;
  assign n24638 = pi207 & n24634;
  assign n24639 = ~n24637 & ~n24638;
  assign n24640 = pi623 & ~n24639;
  assign n24641 = ~n24627 & n24636;
  assign n24642 = ~pi623 & n24568;
  assign n24643 = ~n59888 & ~n24642;
  assign n24644 = ~n7872 & n24643;
  assign n24645 = ~n24580 & ~n24644;
  assign n24646 = ~n24575 & ~n24580;
  assign n24647 = ~n24644 & n24646;
  assign n24648 = ~n24575 & n24645;
  assign n24649 = pi787 & ~n59889;
  assign n24650 = pi641 & ~n7560;
  assign n24651 = ~pi1158 & ~n24650;
  assign n24652 = pi619 & n59884;
  assign n24653 = pi618 & ~n59883;
  assign n24654 = pi609 & ~n24536;
  assign n24655 = n59132 & ~n9797;
  assign n24656 = ~pi778 & ~n24655;
  assign n24657 = ~pi608 & ~n24529;
  assign n24658 = ~pi625 & ~n24655;
  assign n24659 = ~n24530 & ~n24658;
  assign n24660 = ~pi1153 & ~n24659;
  assign n24661 = n24657 & ~n24660;
  assign n24662 = pi608 & ~n24533;
  assign n24663 = pi625 & ~n24655;
  assign n24664 = ~n24526 & ~n24663;
  assign n24665 = pi1153 & ~n24664;
  assign n24666 = n24662 & ~n24665;
  assign n24667 = pi778 & ~n24666;
  assign n24668 = pi778 & ~n24661;
  assign n24669 = ~n24666 & n24668;
  assign n24670 = ~n24661 & n24667;
  assign n24671 = ~n24656 & ~n59890;
  assign n24672 = ~pi609 & ~n24671;
  assign n24673 = ~n24654 & ~n24672;
  assign n24674 = ~pi1155 & ~n24673;
  assign n24675 = pi1155 & ~n7560;
  assign n24676 = ~pi660 & ~n24675;
  assign n24677 = ~n24674 & n24676;
  assign n24678 = ~pi609 & ~n24536;
  assign n24679 = pi609 & ~n24671;
  assign n24680 = ~n24678 & ~n24679;
  assign n24681 = pi1155 & ~n24680;
  assign n24682 = ~pi1155 & ~n7560;
  assign n24683 = pi660 & ~n24682;
  assign n24684 = ~n24681 & n24683;
  assign n24685 = ~n24677 & ~n24684;
  assign n24686 = pi785 & ~n24685;
  assign n24687 = ~pi785 & n24671;
  assign n24688 = ~n24686 & ~n24687;
  assign n24689 = ~pi618 & n24688;
  assign n24690 = ~n24653 & ~n24689;
  assign n24691 = ~pi1154 & ~n24690;
  assign n24692 = pi1154 & ~n7560;
  assign n24693 = ~pi627 & ~n24692;
  assign n24694 = ~n24691 & n24693;
  assign n24695 = ~pi618 & ~n59883;
  assign n24696 = pi618 & n24688;
  assign n24697 = ~n24695 & ~n24696;
  assign n24698 = pi1154 & ~n24697;
  assign n24699 = ~pi1154 & ~n7560;
  assign n24700 = pi627 & ~n24699;
  assign n24701 = ~n24698 & n24700;
  assign n24702 = ~n24694 & ~n24701;
  assign n24703 = pi781 & ~n24702;
  assign n24704 = ~pi781 & ~n24688;
  assign n24705 = ~n24703 & ~n24704;
  assign n24706 = ~pi619 & n24705;
  assign n24707 = ~n24652 & ~n24706;
  assign n24708 = ~pi1159 & ~n24707;
  assign n24709 = pi1159 & ~n7560;
  assign n24710 = ~pi648 & ~n24709;
  assign n24711 = ~n24708 & n24710;
  assign n24712 = ~pi619 & n59884;
  assign n24713 = pi619 & n24705;
  assign n24714 = ~n24712 & ~n24713;
  assign n24715 = pi1159 & ~n24714;
  assign n24716 = ~pi1159 & ~n7560;
  assign n24717 = pi648 & ~n24716;
  assign n24718 = ~n24715 & n24717;
  assign n24719 = ~n24711 & ~n24718;
  assign n24720 = pi789 & ~n24719;
  assign n24721 = ~pi789 & ~n24705;
  assign n24722 = ~n24720 & ~n24721;
  assign n24723 = ~pi626 & ~n24722;
  assign n24724 = pi626 & n59885;
  assign n24725 = ~pi641 & ~n24724;
  assign n24726 = ~n24723 & n24725;
  assign n24727 = n24651 & ~n24726;
  assign n24728 = ~pi641 & ~n7560;
  assign n24729 = pi1158 & ~n24728;
  assign n24730 = pi626 & ~n24722;
  assign n24731 = ~pi626 & n59885;
  assign n24732 = pi641 & ~n24731;
  assign n24733 = ~n24730 & n24732;
  assign n24734 = n24729 & ~n24733;
  assign n24735 = ~n24727 & ~n24734;
  assign n24736 = pi788 & ~n24735;
  assign n24737 = ~pi788 & ~n24722;
  assign n24738 = ~n59357 & ~n24737;
  assign n24739 = ~n24736 & n24738;
  assign n24740 = ~pi628 & ~n7560;
  assign n24741 = pi628 & n59886;
  assign n24742 = ~n24740 & ~n24741;
  assign n24743 = ~pi629 & ~n24742;
  assign n24744 = ~n24740 & ~n24743;
  assign n24745 = pi1156 & ~n24744;
  assign n24746 = ~pi628 & ~n59886;
  assign n24747 = pi628 & n7560;
  assign n24748 = n7791 & ~n24747;
  assign n24749 = pi628 & ~n7560;
  assign n24750 = ~pi628 & n59886;
  assign n24751 = ~n24749 & ~n24750;
  assign n24752 = n7791 & ~n24751;
  assign n24753 = ~n24746 & n24748;
  assign n24754 = ~pi1156 & n24749;
  assign n24755 = n7958 & ~n24747;
  assign n24756 = ~n59891 & ~n59892;
  assign n24757 = ~n24745 & n24756;
  assign n24758 = pi792 & ~n24757;
  assign n24759 = ~n24739 & ~n24758;
  assign n24760 = ~pi207 & ~n24759;
  assign n24761 = ~pi609 & ~n24515;
  assign n24762 = pi1155 & ~n24761;
  assign n24763 = pi660 & n24762;
  assign n24764 = n7626 & ~n24761;
  assign n24765 = ~pi609 & ~n59893;
  assign n24766 = pi609 & ~n24515;
  assign n24767 = ~pi1155 & ~n24766;
  assign n24768 = ~pi660 & n24767;
  assign n24769 = n7625 & ~n24766;
  assign n24770 = pi609 & ~n59894;
  assign n24771 = pi785 & ~n24770;
  assign n24772 = ~n24765 & n24771;
  assign n24773 = pi625 & n13394;
  assign n24774 = pi1153 & ~n24773;
  assign n24775 = ~pi608 & ~n24774;
  assign n24776 = ~pi625 & n23975;
  assign n24777 = ~pi1153 & ~n24776;
  assign n24778 = n24775 & ~n24777;
  assign n24779 = ~pi625 & n13394;
  assign n24780 = ~pi1153 & ~n24779;
  assign n24781 = pi608 & ~n24780;
  assign n24782 = pi625 & n23975;
  assign n24783 = pi1153 & ~n24782;
  assign n24784 = n24781 & ~n24783;
  assign n24785 = pi778 & ~n24784;
  assign n24786 = pi778 & ~n24778;
  assign n24787 = ~n24784 & n24786;
  assign n24788 = ~n24778 & n24785;
  assign n24789 = ~pi778 & ~n23975;
  assign n24790 = pi785 & ~n59894;
  assign n24791 = ~n59893 & n24790;
  assign n24792 = ~n24789 & ~n24791;
  assign n24793 = ~n59895 & n24792;
  assign n24794 = ~n59895 & ~n24789;
  assign n24795 = ~pi609 & ~n24794;
  assign n24796 = n59894 & ~n24795;
  assign n24797 = pi609 & ~n24794;
  assign n24798 = n59893 & ~n24797;
  assign n24799 = ~n24796 & ~n24798;
  assign n24800 = pi785 & ~n24799;
  assign n24801 = ~pi785 & n24794;
  assign n24802 = ~n24800 & ~n24801;
  assign n24803 = ~n24772 & ~n24793;
  assign n24804 = ~n10826 & ~n59896;
  assign n24805 = ~n59229 & n24515;
  assign n24806 = pi781 & ~n10832;
  assign n24807 = n24805 & n24806;
  assign n24808 = ~n24804 & ~n24807;
  assign n24809 = ~pi618 & n59896;
  assign n24810 = pi618 & ~n24805;
  assign n24811 = n7671 & ~n24810;
  assign n24812 = ~n24809 & n24811;
  assign n24813 = pi618 & n59896;
  assign n24814 = ~pi618 & ~n24805;
  assign n24815 = n7672 & ~n24814;
  assign n24816 = ~n24813 & n24815;
  assign n24817 = pi781 & ~n24816;
  assign n24818 = pi781 & ~n24812;
  assign n24819 = ~n24816 & n24818;
  assign n24820 = ~n24812 & n24817;
  assign n24821 = ~pi781 & n59896;
  assign n24822 = ~n12513 & ~n24821;
  assign n24823 = ~n59897 & n24822;
  assign n24824 = ~n12513 & ~n24808;
  assign n24825 = n7715 & n10741;
  assign n24826 = n24516 & n24825;
  assign n24827 = ~n59898 & ~n24826;
  assign n24828 = n59242 & ~n24827;
  assign n24829 = ~n7983 & n8054;
  assign n24830 = n24517 & n24829;
  assign n24831 = ~n24828 & ~n24830;
  assign n24832 = ~pi626 & n24827;
  assign n24833 = pi626 & ~n24517;
  assign n24834 = ~pi641 & ~n24833;
  assign n24835 = ~pi1158 & n24834;
  assign n24836 = ~n24832 & n24835;
  assign n24837 = pi626 & n24827;
  assign n24838 = ~pi626 & ~n24517;
  assign n24839 = pi641 & ~n24838;
  assign n24840 = pi1158 & n24839;
  assign n24841 = ~n24837 & n24840;
  assign n24842 = pi788 & ~n24841;
  assign n24843 = pi788 & ~n24836;
  assign n24844 = ~n24841 & n24843;
  assign n24845 = ~n24836 & n24842;
  assign n24846 = ~pi788 & n24827;
  assign n24847 = ~n59357 & ~n24846;
  assign n24848 = ~n59899 & n24847;
  assign n24849 = ~n59357 & ~n24831;
  assign n24850 = n7793 & n7959;
  assign n24851 = n59882 & n24850;
  assign n24852 = ~n59900 & ~n24851;
  assign n24853 = pi207 & ~n24852;
  assign n24854 = ~pi623 & ~n24853;
  assign n24855 = ~n24760 & n24854;
  assign n24856 = pi1156 & n24743;
  assign n24857 = ~n11154 & n24623;
  assign n24858 = ~n59891 & ~n24857;
  assign n24859 = ~n24856 & n24858;
  assign n24860 = pi792 & ~n24859;
  assign n24861 = n59132 & n59320;
  assign n24862 = ~pi778 & ~n24861;
  assign n24863 = pi625 & n24861;
  assign n24864 = ~pi625 & n24582;
  assign n24865 = pi1153 & ~n24864;
  assign n24866 = pi1153 & ~n24863;
  assign n24867 = ~n24864 & n24866;
  assign n24868 = ~n24863 & n24865;
  assign n24869 = n24662 & ~n59901;
  assign n24870 = pi625 & n24582;
  assign n24871 = ~pi625 & n24861;
  assign n24872 = ~pi1153 & ~n24871;
  assign n24873 = ~n24870 & n24872;
  assign n24874 = n24657 & ~n24873;
  assign n24875 = pi778 & ~n24874;
  assign n24876 = pi778 & ~n24869;
  assign n24877 = ~n24874 & n24876;
  assign n24878 = ~n24869 & n24875;
  assign n24879 = ~n24862 & ~n59902;
  assign n24880 = ~pi609 & ~n24879;
  assign n24881 = ~n24654 & ~n24880;
  assign n24882 = ~pi1155 & ~n24881;
  assign n24883 = ~pi660 & ~n24593;
  assign n24884 = ~n24882 & n24883;
  assign n24885 = pi609 & ~n24879;
  assign n24886 = ~n24678 & ~n24885;
  assign n24887 = pi1155 & ~n24886;
  assign n24888 = pi660 & ~n24589;
  assign n24889 = ~n24887 & n24888;
  assign n24890 = ~n24884 & ~n24889;
  assign n24891 = pi785 & ~n24890;
  assign n24892 = ~pi785 & n24879;
  assign n24893 = ~n24891 & ~n24892;
  assign n24894 = ~pi618 & n24893;
  assign n24895 = ~n24653 & ~n24894;
  assign n24896 = ~pi1154 & ~n24895;
  assign n24897 = ~pi627 & ~n24605;
  assign n24898 = ~n24896 & n24897;
  assign n24899 = pi618 & n24893;
  assign n24900 = ~n24695 & ~n24899;
  assign n24901 = pi1154 & ~n24900;
  assign n24902 = pi627 & ~n24601;
  assign n24903 = ~n24901 & n24902;
  assign n24904 = ~n24898 & ~n24903;
  assign n24905 = pi781 & ~n24904;
  assign n24906 = ~pi781 & ~n24893;
  assign n24907 = ~n24905 & ~n24906;
  assign n24908 = ~pi619 & n24907;
  assign n24909 = ~n24652 & ~n24908;
  assign n24910 = ~pi1159 & ~n24909;
  assign n24911 = ~pi648 & ~n24617;
  assign n24912 = ~n24910 & n24911;
  assign n24913 = pi619 & n24907;
  assign n24914 = ~n24712 & ~n24913;
  assign n24915 = pi1159 & ~n24914;
  assign n24916 = pi648 & ~n24613;
  assign n24917 = ~n24915 & n24916;
  assign n24918 = pi789 & ~n24917;
  assign n24919 = pi789 & ~n24912;
  assign n24920 = ~n24917 & n24919;
  assign n24921 = ~n24912 & n24918;
  assign n24922 = ~pi789 & n24907;
  assign n24923 = n59242 & ~n24922;
  assign n24924 = ~n59903 & n24923;
  assign n24925 = n12139 & n24620;
  assign n24926 = pi641 & ~n59885;
  assign n24927 = ~pi626 & n24729;
  assign n24928 = n7911 & ~n24728;
  assign n24929 = ~n24926 & n59904;
  assign n24930 = ~pi641 & ~n59885;
  assign n24931 = pi626 & n24651;
  assign n24932 = n7912 & ~n24650;
  assign n24933 = ~n24930 & n59905;
  assign n24934 = ~n24929 & ~n24933;
  assign n24935 = ~n24925 & n24934;
  assign n24936 = pi788 & ~n24935;
  assign n24937 = ~n59357 & ~n24936;
  assign n24938 = ~n24924 & n24937;
  assign n24939 = ~n24860 & ~n24938;
  assign n24940 = ~pi207 & ~n24939;
  assign n24941 = ~pi778 & ~n23982;
  assign n24942 = ~pi625 & n23982;
  assign n24943 = pi625 & n24628;
  assign n24944 = ~pi1153 & ~n24943;
  assign n24945 = ~n24942 & n24944;
  assign n24946 = n24775 & ~n24945;
  assign n24947 = pi625 & n23982;
  assign n24948 = ~pi625 & n24628;
  assign n24949 = pi1153 & ~n24948;
  assign n24950 = ~n24947 & n24949;
  assign n24951 = n24781 & ~n24950;
  assign n24952 = pi778 & ~n24951;
  assign n24953 = pi778 & ~n24946;
  assign n24954 = ~n24951 & n24953;
  assign n24955 = ~n24946 & n24952;
  assign n24956 = ~n24941 & ~n59906;
  assign n24957 = ~pi785 & ~n24956;
  assign n24958 = ~pi609 & ~n24956;
  assign n24959 = n24767 & ~n24958;
  assign n24960 = n10731 & n24629;
  assign n24961 = ~pi660 & ~n24960;
  assign n24962 = ~n24959 & n24961;
  assign n24963 = pi609 & ~n24956;
  assign n24964 = n24762 & ~n24963;
  assign n24965 = n10730 & n24629;
  assign n24966 = pi660 & ~n24965;
  assign n24967 = ~n24964 & n24966;
  assign n24968 = ~n24962 & ~n24967;
  assign n24969 = pi785 & ~n24968;
  assign n24970 = ~n24957 & ~n24969;
  assign n24971 = pi618 & ~n24970;
  assign n24972 = pi1154 & ~n24814;
  assign n24973 = ~n24971 & n24972;
  assign n24974 = n10742 & n24630;
  assign n24975 = pi627 & ~n24974;
  assign n24976 = ~n24973 & n24975;
  assign n24977 = ~pi1154 & ~n24810;
  assign n24978 = n10743 & n24630;
  assign n24979 = ~pi627 & ~n24978;
  assign n24980 = ~n24977 & n24979;
  assign n24981 = ~n24976 & ~n24980;
  assign n24982 = pi781 & ~n24981;
  assign n24983 = ~pi618 & ~pi627;
  assign n24984 = pi781 & ~n24983;
  assign n24985 = ~n24970 & ~n24984;
  assign n24986 = pi1159 & ~n24631;
  assign n24987 = ~pi1159 & ~n24516;
  assign n24988 = pi619 & ~pi648;
  assign n24989 = ~n24987 & n24988;
  assign n24990 = ~n24986 & n24988;
  assign n24991 = ~n24987 & n24990;
  assign n24992 = ~n24986 & n24989;
  assign n24993 = ~pi1159 & ~n24631;
  assign n24994 = pi1159 & ~n24516;
  assign n24995 = ~pi619 & pi648;
  assign n24996 = ~n24994 & n24995;
  assign n24997 = ~n24993 & n24995;
  assign n24998 = ~n24994 & n24997;
  assign n24999 = ~n24993 & n24996;
  assign n25000 = pi789 & ~n59908;
  assign n25001 = ~n59907 & n25000;
  assign n25002 = ~n59416 & n25001;
  assign n25003 = ~n24985 & ~n25002;
  assign n25004 = ~n59907 & ~n59908;
  assign n25005 = pi789 & ~n25001;
  assign n25006 = pi789 & ~n25004;
  assign n25007 = ~n12513 & ~n24985;
  assign n25008 = ~n24982 & n25007;
  assign n25009 = ~n59909 & ~n25008;
  assign n25010 = ~n24982 & n25003;
  assign n25011 = n59242 & ~n59910;
  assign n25012 = n7982 & n24632;
  assign n25013 = n7981 & n24517;
  assign n25014 = pi1158 & ~n25013;
  assign n25015 = ~n25012 & n25014;
  assign n25016 = n7981 & n24632;
  assign n25017 = n7982 & n24517;
  assign n25018 = ~pi1158 & ~n25017;
  assign n25019 = ~n25016 & n25018;
  assign n25020 = pi788 & ~n25019;
  assign n25021 = ~n25015 & n25020;
  assign n25022 = ~n25011 & ~n25021;
  assign n25023 = ~pi626 & n59910;
  assign n25024 = n24834 & ~n25023;
  assign n25025 = ~pi1158 & ~n25016;
  assign n25026 = ~n25024 & n25025;
  assign n25027 = pi626 & n59910;
  assign n25028 = n24839 & ~n25027;
  assign n25029 = pi1158 & ~n25012;
  assign n25030 = ~n25028 & n25029;
  assign n25031 = ~n25026 & ~n25030;
  assign n25032 = pi788 & ~n25031;
  assign n25033 = ~pi788 & n59910;
  assign n25034 = ~n59357 & ~n25033;
  assign n25035 = ~n25032 & n25034;
  assign n25036 = ~n59357 & ~n25022;
  assign n25037 = n11150 & n24633;
  assign n25038 = n11152 & n59882;
  assign n25039 = pi1156 & ~n25038;
  assign n25040 = ~n25037 & n25039;
  assign n25041 = n11152 & n24633;
  assign n25042 = n11150 & n59882;
  assign n25043 = ~pi1156 & ~n25042;
  assign n25044 = ~n25041 & n25043;
  assign n25045 = pi792 & ~n25044;
  assign n25046 = pi1156 & ~n24633;
  assign n25047 = ~pi1156 & ~n59882;
  assign n25048 = n11150 & ~n25047;
  assign n25049 = n11150 & ~n25046;
  assign n25050 = ~n25047 & n25049;
  assign n25051 = ~n25046 & n25048;
  assign n25052 = ~pi1156 & ~n24633;
  assign n25053 = pi1156 & ~n59882;
  assign n25054 = n11152 & ~n25053;
  assign n25055 = n11152 & ~n25052;
  assign n25056 = ~n25053 & n25055;
  assign n25057 = ~n25052 & n25054;
  assign n25058 = ~n59912 & ~n59913;
  assign n25059 = pi792 & ~n25058;
  assign n25060 = ~n25040 & n25045;
  assign n25061 = ~n59911 & ~n59914;
  assign n25062 = pi207 & ~n25061;
  assign n25063 = pi623 & ~n25062;
  assign n25064 = ~n24940 & n25063;
  assign n25065 = pi710 & ~n25064;
  assign n25066 = ~n24855 & n25065;
  assign n25067 = ~pi710 & ~n24643;
  assign n25068 = ~n8108 & ~n25067;
  assign n25069 = ~n25066 & n25068;
  assign n25070 = ~n24649 & ~n25069;
  assign n25071 = ~pi790 & ~n25070;
  assign n25072 = ~pi644 & n25070;
  assign n25073 = ~pi787 & ~n24570;
  assign n25074 = ~n24574 & ~n24579;
  assign n25075 = pi787 & ~n25074;
  assign n25076 = ~n25073 & ~n25075;
  assign n25077 = pi644 & n25076;
  assign n25078 = ~pi715 & ~n25077;
  assign n25079 = ~n25072 & n25078;
  assign n25080 = ~n7835 & ~n24643;
  assign n25081 = n7835 & n24568;
  assign n25082 = n7835 & ~n24568;
  assign n25083 = ~n7835 & n24643;
  assign n25084 = ~n25082 & ~n25083;
  assign n25085 = ~n25080 & ~n25081;
  assign n25086 = ~pi644 & n59915;
  assign n25087 = pi644 & n24568;
  assign n25088 = pi715 & ~n25087;
  assign n25089 = ~n25086 & n25088;
  assign n25090 = ~pi1160 & ~n25089;
  assign n25091 = ~n25079 & n25090;
  assign n25092 = pi644 & n25070;
  assign n25093 = ~pi644 & n25076;
  assign n25094 = pi715 & ~n25093;
  assign n25095 = ~n25092 & n25094;
  assign n25096 = pi644 & n59915;
  assign n25097 = ~pi644 & n24568;
  assign n25098 = ~pi715 & ~n25097;
  assign n25099 = ~n25096 & n25098;
  assign n25100 = pi1160 & ~n25099;
  assign n25101 = ~n25095 & n25100;
  assign n25102 = pi790 & ~n25101;
  assign n25103 = pi790 & ~n25091;
  assign n25104 = ~n25101 & n25103;
  assign n25105 = ~n25091 & n25102;
  assign n25106 = ~n25091 & ~n25101;
  assign n25107 = pi790 & ~n25106;
  assign n25108 = ~pi790 & n25070;
  assign n25109 = ~n25107 & ~n25108;
  assign n25110 = ~n25071 & ~n59916;
  assign n25111 = n58992 & n59917;
  assign n25112 = pi207 & ~n58992;
  assign n25113 = n58992 & ~n59917;
  assign n25114 = ~pi207 & ~n58992;
  assign n25115 = ~n25113 & ~n25114;
  assign n25116 = ~n25111 & ~n25112;
  assign n25117 = pi208 & ~n24520;
  assign n25118 = ~pi208 & ~n59887;
  assign n25119 = ~n25117 & ~n25118;
  assign n25120 = pi638 & ~n25119;
  assign n25121 = ~pi208 & ~n7560;
  assign n25122 = ~pi638 & ~n25121;
  assign n25123 = ~n25120 & ~n25122;
  assign n25124 = ~pi647 & n25123;
  assign n25125 = pi647 & n25121;
  assign n25126 = ~pi1157 & ~n25125;
  assign n25127 = ~n25124 & n25126;
  assign n25128 = pi630 & n25127;
  assign n25129 = pi647 & n25123;
  assign n25130 = ~pi647 & n25121;
  assign n25131 = pi1157 & ~n25130;
  assign n25132 = ~n25129 & n25131;
  assign n25133 = ~pi630 & n25132;
  assign n25134 = ~pi208 & ~n24626;
  assign n25135 = pi208 & ~n24634;
  assign n25136 = pi607 & ~n25135;
  assign n25137 = ~pi208 & n24626;
  assign n25138 = pi208 & n24634;
  assign n25139 = ~n25137 & ~n25138;
  assign n25140 = pi607 & ~n25139;
  assign n25141 = ~n25134 & n25136;
  assign n25142 = ~pi607 & n25121;
  assign n25143 = ~n59919 & ~n25142;
  assign n25144 = ~n7872 & n25143;
  assign n25145 = ~n25133 & ~n25144;
  assign n25146 = ~n25128 & ~n25133;
  assign n25147 = ~n25144 & n25146;
  assign n25148 = ~n25128 & n25145;
  assign n25149 = pi787 & ~n59920;
  assign n25150 = ~pi208 & ~n24759;
  assign n25151 = pi208 & ~n24852;
  assign n25152 = ~pi607 & ~n25151;
  assign n25153 = ~n25150 & n25152;
  assign n25154 = ~pi208 & ~n24939;
  assign n25155 = pi208 & ~n25061;
  assign n25156 = pi607 & ~n25155;
  assign n25157 = ~n25154 & n25156;
  assign n25158 = pi638 & ~n25157;
  assign n25159 = ~n25153 & n25158;
  assign n25160 = ~pi638 & ~n25143;
  assign n25161 = ~n8108 & ~n25160;
  assign n25162 = ~n25159 & n25161;
  assign n25163 = ~n25149 & ~n25162;
  assign n25164 = ~pi790 & ~n25163;
  assign n25165 = ~pi644 & n25163;
  assign n25166 = ~pi787 & ~n25123;
  assign n25167 = ~n25127 & ~n25132;
  assign n25168 = pi787 & ~n25167;
  assign n25169 = ~n25166 & ~n25168;
  assign n25170 = pi644 & n25169;
  assign n25171 = ~pi715 & ~n25170;
  assign n25172 = ~n25165 & n25171;
  assign n25173 = ~n7835 & ~n25143;
  assign n25174 = n7835 & n25121;
  assign n25175 = n7835 & ~n25121;
  assign n25176 = ~n7835 & n25143;
  assign n25177 = ~n25175 & ~n25176;
  assign n25178 = ~n25173 & ~n25174;
  assign n25179 = ~pi644 & n59921;
  assign n25180 = pi644 & n25121;
  assign n25181 = pi715 & ~n25180;
  assign n25182 = ~n25179 & n25181;
  assign n25183 = ~pi1160 & ~n25182;
  assign n25184 = ~n25172 & n25183;
  assign n25185 = pi644 & n25163;
  assign n25186 = ~pi644 & n25169;
  assign n25187 = pi715 & ~n25186;
  assign n25188 = ~n25185 & n25187;
  assign n25189 = pi644 & n59921;
  assign n25190 = ~pi644 & n25121;
  assign n25191 = ~pi715 & ~n25190;
  assign n25192 = ~n25189 & n25191;
  assign n25193 = pi1160 & ~n25192;
  assign n25194 = ~n25188 & n25193;
  assign n25195 = pi790 & ~n25194;
  assign n25196 = pi790 & ~n25184;
  assign n25197 = ~n25194 & n25196;
  assign n25198 = ~n25184 & n25195;
  assign n25199 = ~n25184 & ~n25194;
  assign n25200 = pi790 & ~n25199;
  assign n25201 = ~pi790 & n25163;
  assign n25202 = ~n25200 & ~n25201;
  assign n25203 = ~n25164 & ~n59922;
  assign n25204 = n58992 & n59923;
  assign n25205 = pi208 & ~n58992;
  assign n25206 = n58992 & ~n59923;
  assign n25207 = ~pi208 & ~n58992;
  assign n25208 = ~n25206 & ~n25207;
  assign n25209 = ~n25204 & ~n25205;
  assign n25210 = ~n8108 & ~n24759;
  assign n25211 = ~pi647 & ~n7560;
  assign n25212 = pi647 & n59887;
  assign n25213 = ~n25211 & ~n25212;
  assign n25214 = ~pi630 & ~n25213;
  assign n25215 = ~n25211 & ~n25214;
  assign n25216 = pi1157 & ~n25215;
  assign n25217 = pi647 & n7560;
  assign n25218 = pi647 & ~n7560;
  assign n25219 = ~pi1157 & n25218;
  assign n25220 = n8104 & ~n25217;
  assign n25221 = ~pi647 & ~n59887;
  assign n25222 = n7833 & ~n25217;
  assign n25223 = ~pi647 & n59887;
  assign n25224 = ~n25218 & ~n25223;
  assign n25225 = n7833 & ~n25224;
  assign n25226 = ~n25221 & n25222;
  assign n25227 = ~n59925 & ~n59926;
  assign n25228 = ~n25216 & n25227;
  assign n25229 = pi787 & ~n25228;
  assign n25230 = ~n25210 & ~n25229;
  assign n25231 = ~pi644 & ~n25230;
  assign n25232 = ~n9743 & ~n59887;
  assign n25233 = n7560 & n9743;
  assign n25234 = ~n9743 & n59887;
  assign n25235 = ~n7560 & n9743;
  assign n25236 = ~n25234 & ~n25235;
  assign n25237 = ~n25232 & ~n25233;
  assign n25238 = pi644 & ~n59927;
  assign n25239 = ~pi715 & ~n25238;
  assign n25240 = ~n25231 & n25239;
  assign n25241 = pi715 & n7560;
  assign n25242 = ~pi1160 & ~n25241;
  assign n25243 = ~n25240 & n25242;
  assign n25244 = pi644 & ~n25230;
  assign n25245 = ~pi644 & ~n59927;
  assign n25246 = pi715 & ~n25245;
  assign n25247 = ~n25244 & n25246;
  assign n25248 = ~pi715 & n7560;
  assign n25249 = pi1160 & ~n25248;
  assign n25250 = ~n25247 & n25249;
  assign n25251 = ~n25243 & ~n25250;
  assign n25252 = pi790 & ~n25251;
  assign n25253 = ~pi790 & ~n25230;
  assign n25254 = n58992 & ~n25253;
  assign n25255 = ~n25252 & n25254;
  assign n25256 = pi639 & n25255;
  assign n25257 = n4441 & n59132;
  assign n25258 = ~pi57 & n25257;
  assign n25259 = n58992 & n59132;
  assign n25260 = n58992 & n7560;
  assign n25261 = n7553 & n59928;
  assign n25262 = ~pi639 & n59929;
  assign n25263 = ~pi622 & ~n25262;
  assign n25264 = ~n25256 & n25263;
  assign n25265 = ~n8108 & ~n24939;
  assign n25266 = pi1157 & n25214;
  assign n25267 = ~n7872 & n24626;
  assign n25268 = ~n59926 & ~n25267;
  assign n25269 = ~n25266 & n25268;
  assign n25270 = pi787 & ~n25269;
  assign n25271 = ~n25265 & ~n25270;
  assign n25272 = ~pi644 & ~n25271;
  assign n25273 = n25239 & ~n25272;
  assign n25274 = ~n7835 & ~n24626;
  assign n25275 = n7560 & n7835;
  assign n25276 = ~n7560 & n7835;
  assign n25277 = ~n7835 & n24626;
  assign n25278 = ~n25276 & ~n25277;
  assign n25279 = ~n25274 & ~n25275;
  assign n25280 = ~pi644 & n59930;
  assign n25281 = pi644 & n7560;
  assign n25282 = pi644 & ~n7560;
  assign n25283 = ~pi644 & ~n59930;
  assign n25284 = ~n25282 & ~n25283;
  assign n25285 = ~n25280 & ~n25281;
  assign n25286 = pi715 & n59931;
  assign n25287 = ~pi1160 & ~n25286;
  assign n25288 = ~n25273 & n25287;
  assign n25289 = pi644 & ~n25271;
  assign n25290 = n25246 & ~n25289;
  assign n25291 = pi644 & n59930;
  assign n25292 = ~pi644 & n7560;
  assign n25293 = ~pi644 & ~n7560;
  assign n25294 = pi644 & ~n59930;
  assign n25295 = ~n25293 & ~n25294;
  assign n25296 = ~n25291 & ~n25292;
  assign n25297 = ~pi715 & n59932;
  assign n25298 = pi1160 & ~n25297;
  assign n25299 = ~n25290 & n25298;
  assign n25300 = ~n25288 & ~n25299;
  assign n25301 = pi790 & ~n25300;
  assign n25302 = ~pi790 & ~n25271;
  assign n25303 = n58992 & ~n25302;
  assign n25304 = ~n25301 & n25303;
  assign n25305 = pi639 & n25304;
  assign n25306 = ~pi1160 & n59931;
  assign n25307 = pi1160 & n59932;
  assign n25308 = pi790 & ~n25307;
  assign n25309 = pi790 & ~n25306;
  assign n25310 = ~n25307 & n25309;
  assign n25311 = ~n25306 & n25308;
  assign n25312 = ~pi790 & ~n59930;
  assign n25313 = n58992 & ~n25312;
  assign n25314 = ~n59933 & n25313;
  assign n25315 = ~pi639 & n25314;
  assign n25316 = pi622 & ~n25315;
  assign n25317 = ~n25305 & n25316;
  assign n25318 = ~n25264 & ~n25317;
  assign n25319 = ~pi209 & ~n25318;
  assign n25320 = pi1157 & ~n24634;
  assign n25321 = ~pi1157 & ~n24520;
  assign n25322 = n7868 & ~n25321;
  assign n25323 = ~n25320 & n25322;
  assign n25324 = ~pi1157 & ~n24634;
  assign n25325 = pi1157 & ~n24520;
  assign n25326 = n7870 & ~n25325;
  assign n25327 = ~n25324 & n25326;
  assign n25328 = ~n25323 & ~n25327;
  assign n25329 = pi787 & ~n25328;
  assign n25330 = ~n8108 & ~n25061;
  assign n25331 = ~pi647 & ~n25061;
  assign n25332 = pi647 & n24634;
  assign n25333 = ~pi1157 & ~n25332;
  assign n25334 = ~n25331 & n25333;
  assign n25335 = pi647 & n24520;
  assign n25336 = pi1157 & ~n25335;
  assign n25337 = ~pi630 & ~n25336;
  assign n25338 = ~n25334 & n25337;
  assign n25339 = pi647 & ~n25061;
  assign n25340 = ~pi647 & n24634;
  assign n25341 = pi1157 & ~n25340;
  assign n25342 = ~n25339 & n25341;
  assign n25343 = ~pi647 & n24520;
  assign n25344 = ~pi1157 & ~n25343;
  assign n25345 = pi630 & ~n25344;
  assign n25346 = ~n25342 & n25345;
  assign n25347 = ~n25338 & ~n25346;
  assign n25348 = pi787 & ~n25347;
  assign n25349 = ~pi787 & ~n25061;
  assign n25350 = ~n25348 & ~n25349;
  assign n25351 = ~n25329 & ~n25330;
  assign n25352 = ~pi644 & n59934;
  assign n25353 = ~n9743 & n24520;
  assign n25354 = pi644 & ~n25353;
  assign n25355 = ~pi715 & ~n25354;
  assign n25356 = ~n25352 & n25355;
  assign n25357 = pi715 & n12615;
  assign n25358 = n11491 & n24633;
  assign n25359 = ~pi644 & pi715;
  assign n25360 = n25358 & n25359;
  assign n25361 = n24632 & n25357;
  assign n25362 = ~pi1160 & ~n59935;
  assign n25363 = ~n25356 & n25362;
  assign n25364 = pi644 & n59934;
  assign n25365 = ~pi644 & ~n25353;
  assign n25366 = pi715 & ~n25365;
  assign n25367 = ~n25364 & n25366;
  assign n25368 = ~pi715 & n12603;
  assign n25369 = pi644 & ~pi715;
  assign n25370 = n25358 & n25369;
  assign n25371 = n24632 & n25368;
  assign n25372 = pi1160 & ~n59936;
  assign n25373 = ~n25367 & n25372;
  assign n25374 = ~n25363 & ~n25373;
  assign n25375 = pi790 & ~n25374;
  assign n25376 = ~pi790 & n59934;
  assign n25377 = n58992 & ~n25376;
  assign n25378 = ~n25375 & n25377;
  assign n25379 = pi622 & pi639;
  assign n25380 = ~n25378 & n25379;
  assign n25381 = ~n8108 & ~n24852;
  assign n25382 = n7835 & n8105;
  assign n25383 = n24520 & n25382;
  assign n25384 = ~n25381 & ~n25383;
  assign n25385 = ~n23537 & ~n25384;
  assign n25386 = pi790 & ~n23547;
  assign n25387 = n25353 & n25386;
  assign n25388 = ~n25385 & ~n25387;
  assign n25389 = pi644 & n25384;
  assign n25390 = pi1160 & n25366;
  assign n25391 = ~n25389 & n25390;
  assign n25392 = ~pi644 & n25384;
  assign n25393 = ~pi1160 & n25355;
  assign n25394 = ~n25392 & n25393;
  assign n25395 = pi790 & ~n25394;
  assign n25396 = pi790 & ~n25391;
  assign n25397 = ~n25394 & n25396;
  assign n25398 = ~n25391 & n25395;
  assign n25399 = ~pi790 & n25384;
  assign n25400 = n58992 & ~n25399;
  assign n25401 = ~n59937 & n25400;
  assign n25402 = n58992 & ~n25388;
  assign n25403 = ~pi622 & ~n59938;
  assign n25404 = pi644 & ~pi1160;
  assign n25405 = ~pi644 & pi1160;
  assign n25406 = ~n25404 & ~n25405;
  assign n25407 = pi790 & ~n25406;
  assign n25408 = n58992 & ~n25407;
  assign n25409 = n12602 & n25408;
  assign n25410 = n25358 & n25408;
  assign n25411 = n24632 & n25409;
  assign n25412 = pi622 & n59939;
  assign n25413 = ~pi639 & ~n25412;
  assign n25414 = pi209 & ~n25413;
  assign n25415 = pi639 & ~n25403;
  assign n25416 = ~n25412 & ~n25415;
  assign n25417 = pi209 & ~n25416;
  assign n25418 = ~n25403 & n25414;
  assign n25419 = ~n25380 & n59940;
  assign n25420 = ~n25319 & ~n25419;
  assign n25421 = ~pi695 & ~n25255;
  assign n25422 = pi695 & ~n59929;
  assign n25423 = ~pi217 & ~n25422;
  assign n25424 = ~n25421 & n25423;
  assign n25425 = ~pi695 & n59938;
  assign n25426 = pi217 & ~n25425;
  assign n25427 = ~pi612 & ~n25426;
  assign n25428 = ~n25424 & n25427;
  assign n25429 = ~pi695 & ~n25304;
  assign n25430 = pi695 & ~n25314;
  assign n25431 = ~pi217 & ~n25430;
  assign n25432 = ~n25429 & n25431;
  assign n25433 = ~pi695 & n25378;
  assign n25434 = pi695 & n59939;
  assign n25435 = pi217 & ~n25434;
  assign n25436 = ~n25433 & n25435;
  assign n25437 = pi612 & ~n25436;
  assign n25438 = ~n25432 & n25437;
  assign n25439 = ~n25428 & ~n25438;
  assign n25440 = n2634 & ~n59147;
  assign n25441 = n9184 & ~n25440;
  assign n25442 = pi198 & ~n25441;
  assign n25443 = pi198 & ~n59152;
  assign n25444 = ~n58846 & n25443;
  assign n25445 = pi198 & ~n6464;
  assign n25446 = n2782 & ~n25445;
  assign n25447 = pi198 & ~n6587;
  assign n25448 = ~n2782 & ~n25447;
  assign n25449 = ~n25446 & ~n25448;
  assign n25450 = n58846 & n25449;
  assign n25451 = ~n6629 & ~n25450;
  assign n25452 = ~n25444 & n25451;
  assign n25453 = n6629 & ~n25445;
  assign n25454 = ~pi215 & ~n25453;
  assign n25455 = ~n25452 & n25454;
  assign n25456 = pi198 & ~n6490;
  assign n25457 = ~n25446 & n25456;
  assign n25458 = ~n2778 & ~n6486;
  assign n25459 = n2778 & ~n6484;
  assign n25460 = pi198 & ~n25459;
  assign n25461 = ~n25458 & n25460;
  assign n25462 = ~n58846 & n25461;
  assign n25463 = ~n25457 & ~n25462;
  assign n25464 = pi215 & ~n25463;
  assign n25465 = pi299 & ~n25464;
  assign n25466 = ~n25455 & n25465;
  assign n25467 = ~n2790 & n25443;
  assign n25468 = n2790 & n25449;
  assign n25469 = ~n6544 & ~n25468;
  assign n25470 = ~n25467 & n25469;
  assign n25471 = n6544 & ~n25445;
  assign n25472 = ~pi223 & ~n25471;
  assign n25473 = ~n25470 & n25472;
  assign n25474 = ~n2790 & n25461;
  assign n25475 = ~n25457 & ~n25474;
  assign n25476 = pi223 & ~n25475;
  assign n25477 = ~pi299 & ~n25476;
  assign n25478 = ~n25473 & n25477;
  assign n25479 = ~pi38 & pi39;
  assign n25480 = pi39 & n59292;
  assign n25481 = n59132 & n25479;
  assign n25482 = ~n25478 & n59941;
  assign n25483 = ~n25466 & n59941;
  assign n25484 = ~n25478 & n25483;
  assign n25485 = ~n25466 & n25482;
  assign n25486 = ~n25442 & ~n59942;
  assign n25487 = n8054 & n25486;
  assign n25488 = pi198 & ~n59132;
  assign n25489 = pi633 & n6464;
  assign n25490 = ~n6684 & n25489;
  assign n25491 = ~n25445 & ~n25490;
  assign n25492 = pi603 & ~n25491;
  assign n25493 = ~pi603 & n25445;
  assign n25494 = ~n25492 & ~n25493;
  assign n25495 = ~n6700 & n25494;
  assign n25496 = n2680 & ~n25491;
  assign n25497 = ~n6484 & n25490;
  assign n25498 = ~n25456 & ~n25497;
  assign n25499 = ~n25496 & n25498;
  assign n25500 = pi603 & ~n25499;
  assign n25501 = n6700 & ~n25493;
  assign n25502 = ~n25500 & n25501;
  assign n25503 = ~n25495 & ~n25502;
  assign n25504 = ~n2781 & n25503;
  assign n25505 = ~n25456 & ~n25500;
  assign n25506 = n2781 & ~n25505;
  assign n25507 = ~n25504 & ~n25506;
  assign n25508 = n58846 & n25507;
  assign n25509 = pi633 & n6830;
  assign n25510 = ~n25461 & ~n25509;
  assign n25511 = ~n2781 & ~n25510;
  assign n25512 = pi198 & n6484;
  assign n25513 = ~n25497 & ~n25512;
  assign n25514 = n59159 & ~n25513;
  assign n25515 = ~n25511 & ~n25514;
  assign n25516 = ~n58846 & n25515;
  assign n25517 = pi215 & ~n25516;
  assign n25518 = ~n25508 & n25517;
  assign n25519 = pi198 & n6566;
  assign n25520 = pi633 & n6687;
  assign n25521 = ~n25519 & ~n25520;
  assign n25522 = ~n2680 & ~n25521;
  assign n25523 = ~n25496 & ~n25522;
  assign n25524 = pi603 & ~n25523;
  assign n25525 = ~pi642 & ~n25524;
  assign n25526 = pi642 & ~n25492;
  assign n25527 = n2777 & ~n25526;
  assign n25528 = ~n25525 & n25527;
  assign n25529 = ~n2777 & n25492;
  assign n25530 = ~n25493 & ~n25529;
  assign n25531 = ~n25528 & n25530;
  assign n25532 = ~n2781 & n25531;
  assign n25533 = ~pi603 & n25447;
  assign n25534 = n2781 & ~n25533;
  assign n25535 = ~n25524 & n25534;
  assign n25536 = ~n25532 & ~n25535;
  assign n25537 = n58846 & n25536;
  assign n25538 = n2680 & n25521;
  assign n25539 = ~n2680 & n25491;
  assign n25540 = pi603 & ~n6700;
  assign n25541 = ~n25539 & n25540;
  assign n25542 = ~n25538 & n25541;
  assign n25543 = pi603 & ~n25521;
  assign n25544 = n6700 & n25543;
  assign n25545 = pi198 & n7005;
  assign n25546 = ~n25544 & ~n25545;
  assign n25547 = ~n25542 & n25546;
  assign n25548 = ~n2781 & n25547;
  assign n25549 = n2781 & ~n25519;
  assign n25550 = ~n25543 & n25549;
  assign n25551 = ~n25548 & ~n25550;
  assign n25552 = ~n58846 & n25551;
  assign n25553 = ~n6629 & ~n25552;
  assign n25554 = ~n25537 & n25553;
  assign n25555 = n6629 & n25494;
  assign n25556 = ~pi215 & ~n25555;
  assign n25557 = ~n25554 & n25556;
  assign n25558 = ~n25518 & ~n25557;
  assign n25559 = pi299 & ~n25558;
  assign n25560 = n2790 & n25507;
  assign n25561 = ~n2790 & n25515;
  assign n25562 = pi223 & ~n25561;
  assign n25563 = ~n25560 & n25562;
  assign n25564 = n2790 & n25536;
  assign n25565 = ~n2790 & n25551;
  assign n25566 = ~n6544 & ~n25565;
  assign n25567 = ~n25564 & n25566;
  assign n25568 = n6544 & n25494;
  assign n25569 = ~pi223 & ~n25568;
  assign n25570 = ~n25567 & n25569;
  assign n25571 = ~n25563 & ~n25570;
  assign n25572 = ~pi299 & ~n25571;
  assign n25573 = pi39 & ~n25572;
  assign n25574 = pi39 & ~n25559;
  assign n25575 = ~n25572 & n25574;
  assign n25576 = ~n25559 & n25573;
  assign n25577 = pi198 & ~n6453;
  assign n25578 = pi603 & pi633;
  assign n25579 = ~n25577 & ~n25578;
  assign n25580 = pi198 & ~n6675;
  assign n25581 = ~pi198 & n6795;
  assign n25582 = ~pi198 & ~n6795;
  assign n25583 = pi198 & n6675;
  assign n25584 = ~n25582 & ~n25583;
  assign n25585 = ~n25580 & ~n25581;
  assign n25586 = n25578 & ~n59944;
  assign n25587 = ~n25579 & ~n25586;
  assign n25588 = pi299 & n25587;
  assign n25589 = ~n6661 & ~n6665;
  assign n25590 = pi633 & ~n25589;
  assign n25591 = ~n6448 & ~n25590;
  assign n25592 = ~n6670 & ~n25591;
  assign n25593 = ~pi299 & n25592;
  assign n25594 = ~pi39 & ~n25593;
  assign n25595 = ~n25588 & n25594;
  assign n25596 = ~n59943 & ~n25595;
  assign n25597 = ~pi38 & ~n25596;
  assign n25598 = pi39 & pi198;
  assign n25599 = pi38 & ~n25598;
  assign n25600 = pi198 & ~n6468;
  assign n25601 = pi633 & n6701;
  assign n25602 = n6468 & n25601;
  assign n25603 = ~n25600 & ~n25602;
  assign n25604 = ~pi39 & ~n25603;
  assign n25605 = n25599 & ~n25604;
  assign n25606 = n59132 & ~n25605;
  assign n25607 = ~n25597 & n25606;
  assign n25608 = ~n25488 & ~n25607;
  assign n25609 = ~n7597 & ~n25608;
  assign n25610 = n7597 & ~n25486;
  assign n25611 = ~n25609 & ~n25610;
  assign n25612 = ~pi785 & ~n25611;
  assign n25613 = ~n7598 & ~n25486;
  assign n25614 = pi609 & n25609;
  assign n25615 = ~n25613 & ~n25614;
  assign n25616 = pi1155 & ~n25615;
  assign n25617 = ~n7610 & ~n25486;
  assign n25618 = ~pi609 & n25609;
  assign n25619 = ~n25617 & ~n25618;
  assign n25620 = ~pi1155 & ~n25619;
  assign n25621 = ~n25616 & ~n25620;
  assign n25622 = pi785 & ~n25621;
  assign n25623 = ~n25612 & ~n25622;
  assign n25624 = ~pi781 & ~n25623;
  assign n25625 = pi618 & n25623;
  assign n25626 = ~pi618 & n25486;
  assign n25627 = pi1154 & ~n25626;
  assign n25628 = ~n25625 & n25627;
  assign n25629 = ~pi618 & n25623;
  assign n25630 = pi618 & n25486;
  assign n25631 = ~pi1154 & ~n25630;
  assign n25632 = ~n25629 & n25631;
  assign n25633 = ~n25628 & ~n25632;
  assign n25634 = pi781 & ~n25633;
  assign n25635 = ~n25624 & ~n25634;
  assign n25636 = ~pi789 & ~n25635;
  assign n25637 = pi619 & n25635;
  assign n25638 = ~pi619 & n25486;
  assign n25639 = pi1159 & ~n25638;
  assign n25640 = ~n25637 & n25639;
  assign n25641 = ~pi619 & n25635;
  assign n25642 = pi619 & n25486;
  assign n25643 = ~pi1159 & ~n25642;
  assign n25644 = ~n25641 & n25643;
  assign n25645 = ~n25640 & ~n25644;
  assign n25646 = pi789 & ~n25645;
  assign n25647 = ~n25636 & ~n25646;
  assign n25648 = ~n8054 & n25647;
  assign n25649 = ~n25487 & ~n25648;
  assign n25650 = ~n7793 & ~n25649;
  assign n25651 = n7793 & n25486;
  assign n25652 = ~n7872 & ~n25651;
  assign n25653 = n7793 & ~n25486;
  assign n25654 = ~n7793 & n25649;
  assign n25655 = ~n25653 & ~n25654;
  assign n25656 = ~n7872 & ~n25655;
  assign n25657 = ~n25650 & n25652;
  assign n25658 = ~n9651 & n25486;
  assign n25659 = ~n7035 & ~n25445;
  assign n25660 = pi634 & ~n25659;
  assign n25661 = ~n25445 & ~n25660;
  assign n25662 = ~n2680 & n25661;
  assign n25663 = pi634 & ~n6484;
  assign n25664 = n7035 & n25663;
  assign n25665 = ~n25512 & ~n25664;
  assign n25666 = n2680 & n25665;
  assign n25667 = ~n25662 & ~n25666;
  assign n25668 = ~n2778 & ~n25667;
  assign n25669 = n2778 & n25665;
  assign n25670 = n6871 & ~n25669;
  assign n25671 = ~n25668 & n25670;
  assign n25672 = ~pi680 & n25461;
  assign n25673 = n2781 & ~n25665;
  assign n25674 = ~n25672 & ~n25673;
  assign n25675 = ~n25671 & n25674;
  assign n25676 = ~n58846 & n25675;
  assign n25677 = n2680 & ~n25661;
  assign n25678 = ~n2680 & ~n25665;
  assign n25679 = ~n25677 & ~n25678;
  assign n25680 = n2778 & n25679;
  assign n25681 = ~n2778 & n25661;
  assign n25682 = n6871 & ~n25681;
  assign n25683 = ~n25680 & n25682;
  assign n25684 = n25456 & n25672;
  assign n25685 = n2781 & ~n25679;
  assign n25686 = ~n25684 & ~n25685;
  assign n25687 = ~n25683 & n25686;
  assign n25688 = n58846 & n25687;
  assign n25689 = pi215 & ~n25688;
  assign n25690 = pi215 & ~n25676;
  assign n25691 = ~n25688 & n25690;
  assign n25692 = ~n25676 & n25689;
  assign n25693 = pi634 & ~n59178;
  assign n25694 = ~n25519 & ~n25693;
  assign n25695 = n2680 & n25694;
  assign n25696 = ~n25662 & ~n25695;
  assign n25697 = ~n2778 & ~n25696;
  assign n25698 = n2778 & n25694;
  assign n25699 = n6871 & ~n25698;
  assign n25700 = ~n25697 & n25699;
  assign n25701 = pi198 & n6903;
  assign n25702 = n2781 & ~n25694;
  assign n25703 = ~n25701 & ~n25702;
  assign n25704 = ~n25700 & n25703;
  assign n25705 = ~n58846 & ~n25704;
  assign n25706 = ~n2680 & ~n25694;
  assign n25707 = ~n25677 & ~n25706;
  assign n25708 = n2778 & n25707;
  assign n25709 = n25682 & ~n25708;
  assign n25710 = n2781 & ~n25707;
  assign n25711 = n2778 & ~n25447;
  assign n25712 = ~n2778 & ~n25445;
  assign n25713 = ~pi680 & ~n25712;
  assign n25714 = ~n25711 & n25713;
  assign n25715 = ~n25710 & ~n25714;
  assign n25716 = ~n25709 & n25715;
  assign n25717 = n58846 & ~n25716;
  assign n25718 = ~n6629 & ~n25717;
  assign n25719 = ~n6629 & ~n25705;
  assign n25720 = ~n25717 & n25719;
  assign n25721 = ~n25705 & n25718;
  assign n25722 = pi634 & n6464;
  assign n25723 = n7054 & n25722;
  assign n25724 = pi634 & pi680;
  assign n25725 = pi680 & n25660;
  assign n25726 = ~n25659 & n25724;
  assign n25727 = ~n25445 & ~n59948;
  assign n25728 = n6629 & n25727;
  assign n25729 = n25453 & ~n25723;
  assign n25730 = ~pi215 & ~n59949;
  assign n25731 = ~n59947 & n25730;
  assign n25732 = ~n59946 & ~n25731;
  assign n25733 = pi39 & ~n25732;
  assign n25734 = ~pi198 & n7327;
  assign n25735 = pi198 & ~n7304;
  assign n25736 = ~n25734 & ~n25735;
  assign n25737 = n25724 & n25736;
  assign n25738 = ~n25577 & ~n25724;
  assign n25739 = ~pi39 & ~n25738;
  assign n25740 = ~n25737 & n25739;
  assign n25741 = ~n25733 & ~n25740;
  assign n25742 = pi299 & ~n25741;
  assign n25743 = n2790 & ~n25716;
  assign n25744 = ~n2790 & ~n25704;
  assign n25745 = ~n6544 & ~n25744;
  assign n25746 = ~n6544 & ~n25743;
  assign n25747 = ~n25744 & n25746;
  assign n25748 = ~n25743 & n25745;
  assign n25749 = n6544 & n25727;
  assign n25750 = n25471 & ~n25723;
  assign n25751 = ~pi223 & ~n59951;
  assign n25752 = ~n59950 & n25751;
  assign n25753 = ~n2790 & n25675;
  assign n25754 = n2790 & n25687;
  assign n25755 = pi223 & ~n25754;
  assign n25756 = pi223 & ~n25753;
  assign n25757 = ~n25754 & n25756;
  assign n25758 = ~n25753 & n25755;
  assign n25759 = pi39 & ~n59952;
  assign n25760 = ~n25752 & n25759;
  assign n25761 = pi198 & n7294;
  assign n25762 = ~n7314 & n25724;
  assign n25763 = ~n25761 & n25762;
  assign n25764 = ~n6448 & ~n25763;
  assign n25765 = ~pi39 & n25764;
  assign n25766 = ~pi299 & ~n25765;
  assign n25767 = ~n25760 & n25766;
  assign n25768 = ~pi38 & ~n25767;
  assign n25769 = ~pi299 & ~n59952;
  assign n25770 = ~n25752 & n25769;
  assign n25771 = pi299 & ~n59946;
  assign n25772 = ~n25731 & n25771;
  assign n25773 = ~n25770 & ~n25772;
  assign n25774 = pi39 & ~n25773;
  assign n25775 = pi299 & ~n25738;
  assign n25776 = n25724 & ~n25736;
  assign n25777 = n25577 & ~n25724;
  assign n25778 = ~n25776 & ~n25777;
  assign n25779 = pi299 & ~n25778;
  assign n25780 = ~n25737 & n25775;
  assign n25781 = ~pi299 & ~n25764;
  assign n25782 = ~pi39 & ~n25781;
  assign n25783 = ~n59953 & n25782;
  assign n25784 = ~n25774 & ~n25783;
  assign n25785 = ~pi38 & ~n25784;
  assign n25786 = ~n25742 & n25768;
  assign n25787 = pi634 & n7054;
  assign n25788 = n6468 & n25787;
  assign n25789 = ~n25600 & ~n25788;
  assign n25790 = ~pi39 & ~n25789;
  assign n25791 = n25599 & ~n25790;
  assign n25792 = n59132 & ~n25791;
  assign n25793 = ~n59954 & n25792;
  assign n25794 = ~n25488 & ~n25793;
  assign n25795 = ~pi778 & ~n25794;
  assign n25796 = pi625 & n25794;
  assign n25797 = ~pi625 & n25486;
  assign n25798 = pi1153 & ~n25797;
  assign n25799 = ~n25796 & n25798;
  assign n25800 = ~pi625 & n25794;
  assign n25801 = pi625 & n25486;
  assign n25802 = ~pi1153 & ~n25801;
  assign n25803 = ~n25800 & n25802;
  assign n25804 = ~n25799 & ~n25803;
  assign n25805 = pi778 & ~n25804;
  assign n25806 = ~n25795 & ~n25805;
  assign n25807 = ~n59229 & ~n25806;
  assign n25808 = n59229 & ~n25486;
  assign n25809 = ~n59229 & n25806;
  assign n25810 = n59229 & n25486;
  assign n25811 = ~n25809 & ~n25810;
  assign n25812 = ~n25807 & ~n25808;
  assign n25813 = ~n59231 & ~n59955;
  assign n25814 = n59231 & n25486;
  assign n25815 = n59231 & ~n25486;
  assign n25816 = ~n59231 & n59955;
  assign n25817 = ~n25815 & ~n25816;
  assign n25818 = ~n25813 & ~n25814;
  assign n25819 = ~n7716 & n59956;
  assign n25820 = ~n7762 & n25819;
  assign n25821 = ~n25658 & ~n25820;
  assign n25822 = ~pi792 & n25821;
  assign n25823 = pi628 & ~n25821;
  assign n25824 = ~pi628 & n25486;
  assign n25825 = pi1156 & ~n25824;
  assign n25826 = ~n25823 & ~n25824;
  assign n25827 = pi1156 & n25826;
  assign n25828 = ~n25823 & n25825;
  assign n25829 = ~pi628 & ~n25821;
  assign n25830 = pi628 & n25486;
  assign n25831 = ~pi1156 & ~n25830;
  assign n25832 = ~n25829 & n25831;
  assign n25833 = ~n59957 & ~n25832;
  assign n25834 = pi792 & ~n25833;
  assign n25835 = ~n25822 & ~n25834;
  assign n25836 = pi647 & ~n25835;
  assign n25837 = ~pi647 & ~n25486;
  assign n25838 = ~n25836 & ~n25837;
  assign n25839 = n7832 & ~n25838;
  assign n25840 = ~pi647 & n25835;
  assign n25841 = pi647 & n25486;
  assign n25842 = ~pi1157 & ~n25841;
  assign n25843 = ~n25840 & n25842;
  assign n25844 = pi630 & n25843;
  assign n25845 = ~n25839 & ~n25844;
  assign n25846 = ~n59945 & n25845;
  assign n25847 = pi787 & ~n25846;
  assign n25848 = ~n11154 & n25649;
  assign n25849 = n7790 & n25826;
  assign n25850 = ~pi629 & n59957;
  assign n25851 = pi629 & n25832;
  assign n25852 = ~n59958 & ~n25851;
  assign n25853 = ~n25848 & n25852;
  assign n25854 = pi792 & ~n25853;
  assign n25855 = ~pi626 & ~n25647;
  assign n25856 = pi626 & ~n25486;
  assign n25857 = n7760 & ~n25856;
  assign n25858 = ~n25855 & n25857;
  assign n25859 = n7716 & n25486;
  assign n25860 = ~n25819 & ~n25859;
  assign n25861 = n7984 & ~n25860;
  assign n25862 = pi626 & ~n25647;
  assign n25863 = ~pi626 & ~n25486;
  assign n25864 = n7759 & ~n25863;
  assign n25865 = ~n25862 & n25864;
  assign n25866 = ~n25861 & ~n25865;
  assign n25867 = ~n25858 & ~n25861;
  assign n25868 = ~n25865 & n25867;
  assign n25869 = ~n25858 & n25866;
  assign n25870 = pi788 & ~n59959;
  assign n25871 = ~n6667 & n7295;
  assign n25872 = pi634 & ~n25871;
  assign n25873 = ~pi634 & ~n6448;
  assign n25874 = ~pi633 & ~n25873;
  assign n25875 = ~pi634 & n6448;
  assign n25876 = pi634 & n7295;
  assign n25877 = ~n6667 & n25876;
  assign n25878 = ~n25875 & ~n25877;
  assign n25879 = ~pi633 & ~n25878;
  assign n25880 = ~n25872 & n25874;
  assign n25881 = pi634 & ~pi665;
  assign n25882 = pi198 & ~pi633;
  assign n25883 = n25881 & ~n25882;
  assign n25884 = ~n6659 & n25883;
  assign n25885 = pi603 & ~n25884;
  assign n25886 = ~n25590 & n25885;
  assign n25887 = ~n59960 & n25886;
  assign n25888 = ~pi603 & n25764;
  assign n25889 = pi680 & ~n25888;
  assign n25890 = ~n25590 & ~n25884;
  assign n25891 = ~n59960 & n25890;
  assign n25892 = pi603 & ~n25891;
  assign n25893 = ~pi603 & ~n25764;
  assign n25894 = ~n25892 & ~n25893;
  assign n25895 = pi680 & ~n25894;
  assign n25896 = ~n25887 & n25889;
  assign n25897 = ~pi680 & n25592;
  assign n25898 = ~pi299 & ~n25897;
  assign n25899 = ~n59961 & n25898;
  assign n25900 = ~n6795 & n25735;
  assign n25901 = ~pi198 & ~pi665;
  assign n25902 = n6675 & n25901;
  assign n25903 = ~pi633 & ~n25902;
  assign n25904 = ~n25900 & n25903;
  assign n25905 = pi198 & ~pi665;
  assign n25906 = pi633 & ~n25905;
  assign n25907 = ~n25734 & n25906;
  assign n25908 = ~n59944 & n25907;
  assign n25909 = ~n25904 & ~n25908;
  assign n25910 = pi603 & ~n25909;
  assign n25911 = ~pi603 & n25736;
  assign n25912 = n25724 & ~n25911;
  assign n25913 = ~pi603 & ~n25736;
  assign n25914 = pi603 & ~n25904;
  assign n25915 = ~n25908 & n25914;
  assign n25916 = ~n25913 & ~n25915;
  assign n25917 = n25724 & ~n25916;
  assign n25918 = ~n25910 & n25912;
  assign n25919 = n25587 & ~n25724;
  assign n25920 = pi299 & ~n25919;
  assign n25921 = ~n59962 & n25920;
  assign n25922 = ~n25899 & ~n25921;
  assign n25923 = ~pi39 & ~n25922;
  assign n25924 = ~pi680 & n25531;
  assign n25925 = n6692 & n25881;
  assign n25926 = n25491 & ~n25925;
  assign n25927 = n2680 & ~n25926;
  assign n25928 = pi634 & n59180;
  assign n25929 = n25521 & ~n25928;
  assign n25930 = ~n2680 & ~n25929;
  assign n25931 = ~n25927 & ~n25930;
  assign n25932 = pi603 & ~n25931;
  assign n25933 = ~pi642 & n25932;
  assign n25934 = ~pi603 & ~n25661;
  assign n25935 = pi603 & ~n25926;
  assign n25936 = pi642 & n25935;
  assign n25937 = ~n25934 & ~n25936;
  assign n25938 = ~n25933 & n25937;
  assign n25939 = n2777 & ~n25938;
  assign n25940 = ~n25934 & ~n25935;
  assign n25941 = ~n2777 & ~n25940;
  assign n25942 = ~n6518 & ~n25941;
  assign n25943 = ~n25939 & n25942;
  assign n25944 = ~pi603 & ~n25707;
  assign n25945 = n6518 & ~n25944;
  assign n25946 = ~n25932 & n25945;
  assign n25947 = ~n25943 & ~n25946;
  assign n25948 = pi680 & ~n25947;
  assign n25949 = ~n25924 & ~n25948;
  assign n25950 = n58846 & n25949;
  assign n25951 = ~pi603 & n25696;
  assign n25952 = ~n6700 & n25935;
  assign n25953 = ~n25541 & ~n25952;
  assign n25954 = ~n2778 & n25953;
  assign n25955 = ~n2680 & ~n25953;
  assign n25956 = n25929 & ~n25955;
  assign n25957 = ~n25954 & ~n25956;
  assign n25958 = ~n25951 & ~n25957;
  assign n25959 = n6871 & ~n25958;
  assign n25960 = ~pi680 & ~n25547;
  assign n25961 = ~n6701 & ~n25694;
  assign n25962 = ~n25543 & ~n25961;
  assign n25963 = n2781 & ~n25962;
  assign n25964 = ~n25960 & ~n25963;
  assign n25965 = ~n25959 & n25964;
  assign n25966 = ~n58846 & ~n25965;
  assign n25967 = ~n6629 & ~n25966;
  assign n25968 = ~n25950 & n25967;
  assign n25969 = n6914 & n25660;
  assign n25970 = n25494 & ~n25969;
  assign n25971 = n6629 & n25970;
  assign n25972 = ~pi215 & ~n25971;
  assign n25973 = ~n25968 & n25972;
  assign n25974 = n6721 & n25901;
  assign n25975 = n6684 & n25905;
  assign n25976 = ~n25512 & ~n25975;
  assign n25977 = ~n25974 & n25976;
  assign n25978 = pi634 & ~n25977;
  assign n25979 = ~pi634 & n25512;
  assign n25980 = ~n25497 & ~n25979;
  assign n25981 = ~n25978 & n25980;
  assign n25982 = ~n2680 & ~n25981;
  assign n25983 = ~n25927 & ~n25982;
  assign n25984 = pi603 & ~n25983;
  assign n25985 = n6700 & ~n25934;
  assign n25986 = ~n25984 & n25985;
  assign n25987 = ~n6700 & n25940;
  assign n25988 = n6871 & ~n25987;
  assign n25989 = ~n25986 & n25988;
  assign n25990 = ~pi680 & n25503;
  assign n25991 = ~pi603 & ~n25679;
  assign n25992 = ~n25984 & ~n25991;
  assign n25993 = n2781 & ~n25992;
  assign n25994 = ~n25990 & ~n25993;
  assign n25995 = ~n25989 & n25994;
  assign n25996 = n58846 & n25995;
  assign n25997 = pi603 & ~n25981;
  assign n25998 = n6700 & n25997;
  assign n25999 = ~n25953 & ~n25981;
  assign n26000 = ~n25998 & ~n25999;
  assign n26001 = ~n25954 & ~n25981;
  assign n26002 = ~pi603 & n25667;
  assign n26003 = ~n25955 & ~n26002;
  assign n26004 = n59963 & n26003;
  assign n26005 = n6871 & ~n26004;
  assign n26006 = ~pi680 & ~n25510;
  assign n26007 = pi603 & n25981;
  assign n26008 = ~pi603 & n25665;
  assign n26009 = n2781 & ~n26008;
  assign n26010 = ~pi603 & ~n25665;
  assign n26011 = ~n25997 & ~n26010;
  assign n26012 = n2781 & ~n26011;
  assign n26013 = ~n26007 & n26009;
  assign n26014 = ~n26006 & ~n59964;
  assign n26015 = ~n26005 & n26014;
  assign n26016 = ~n58846 & n26015;
  assign n26017 = pi215 & ~n26016;
  assign n26018 = ~n25996 & n26017;
  assign n26019 = ~n25973 & ~n26018;
  assign n26020 = pi299 & ~n26019;
  assign n26021 = n2790 & n25949;
  assign n26022 = ~n2790 & ~n25965;
  assign n26023 = ~n6544 & ~n26022;
  assign n26024 = ~n26021 & n26023;
  assign n26025 = n6544 & n25970;
  assign n26026 = ~pi223 & ~n26025;
  assign n26027 = ~n26024 & n26026;
  assign n26028 = n2790 & n25995;
  assign n26029 = ~n2790 & n26015;
  assign n26030 = pi223 & ~n26029;
  assign n26031 = ~n26028 & n26030;
  assign n26032 = ~n26027 & ~n26031;
  assign n26033 = ~pi299 & ~n26032;
  assign n26034 = pi39 & ~n26033;
  assign n26035 = pi39 & ~n26020;
  assign n26036 = ~n26033 & n26035;
  assign n26037 = ~n26020 & n26034;
  assign n26038 = ~n25923 & ~n59965;
  assign n26039 = ~pi38 & ~n26038;
  assign n26040 = pi634 & n59208;
  assign n26041 = n25603 & ~n26040;
  assign n26042 = ~pi39 & ~n26041;
  assign n26043 = n25599 & ~n26042;
  assign n26044 = n59132 & ~n26043;
  assign n26045 = ~n26039 & n26044;
  assign n26046 = ~n25488 & ~n26045;
  assign n26047 = ~pi625 & n26046;
  assign n26048 = pi625 & n25608;
  assign n26049 = ~pi1153 & ~n26048;
  assign n26050 = ~n26047 & n26049;
  assign n26051 = ~pi608 & ~n25799;
  assign n26052 = ~n26050 & n26051;
  assign n26053 = pi625 & n26046;
  assign n26054 = ~pi625 & n25608;
  assign n26055 = pi1153 & ~n26054;
  assign n26056 = ~n26053 & n26055;
  assign n26057 = pi608 & ~n25803;
  assign n26058 = ~n26056 & n26057;
  assign n26059 = ~n26052 & ~n26058;
  assign n26060 = pi778 & ~n26059;
  assign n26061 = ~pi778 & n26046;
  assign n26062 = ~n26060 & ~n26061;
  assign n26063 = ~pi609 & ~n26062;
  assign n26064 = pi609 & n25806;
  assign n26065 = ~pi1155 & ~n26064;
  assign n26066 = ~n26063 & n26065;
  assign n26067 = ~pi660 & ~n25616;
  assign n26068 = ~n26066 & n26067;
  assign n26069 = pi609 & ~n26062;
  assign n26070 = ~pi609 & n25806;
  assign n26071 = pi1155 & ~n26070;
  assign n26072 = ~n26069 & n26071;
  assign n26073 = pi660 & ~n25620;
  assign n26074 = ~n26072 & n26073;
  assign n26075 = ~n26068 & ~n26074;
  assign n26076 = pi785 & ~n26075;
  assign n26077 = ~pi785 & ~n26062;
  assign n26078 = ~n26076 & ~n26077;
  assign n26079 = ~pi618 & ~n26078;
  assign n26080 = pi618 & ~n59955;
  assign n26081 = ~pi1154 & ~n26080;
  assign n26082 = ~n26079 & n26081;
  assign n26083 = ~pi627 & ~n25628;
  assign n26084 = ~n26082 & n26083;
  assign n26085 = pi618 & ~n26078;
  assign n26086 = ~pi618 & ~n59955;
  assign n26087 = pi1154 & ~n26086;
  assign n26088 = ~n26085 & n26087;
  assign n26089 = pi627 & ~n25632;
  assign n26090 = ~n26088 & n26089;
  assign n26091 = ~n26084 & ~n26090;
  assign n26092 = pi781 & ~n26091;
  assign n26093 = ~pi781 & ~n26078;
  assign n26094 = ~n26092 & ~n26093;
  assign n26095 = pi619 & ~n26094;
  assign n26096 = ~pi619 & n59956;
  assign n26097 = pi1159 & ~n26096;
  assign n26098 = ~n26095 & n26097;
  assign n26099 = pi648 & ~n25644;
  assign n26100 = ~n26098 & n26099;
  assign n26101 = ~pi619 & ~n26094;
  assign n26102 = pi619 & n59956;
  assign n26103 = ~pi1159 & ~n26102;
  assign n26104 = ~n26101 & n26103;
  assign n26105 = ~pi648 & ~n25640;
  assign n26106 = ~n26104 & n26105;
  assign n26107 = pi789 & ~n26106;
  assign n26108 = pi789 & ~n26100;
  assign n26109 = ~n26106 & n26108;
  assign n26110 = ~n26100 & n26107;
  assign n26111 = ~pi789 & n26094;
  assign n26112 = n59242 & ~n26111;
  assign n26113 = ~n59966 & n26112;
  assign n26114 = ~n25870 & ~n26113;
  assign n26115 = ~n25854 & ~n26114;
  assign n26116 = n59357 & n25853;
  assign n26117 = ~n8108 & ~n26116;
  assign n26118 = ~n26115 & n26117;
  assign n26119 = ~n25847 & ~n26118;
  assign n26120 = ~n23537 & n26119;
  assign n26121 = pi1157 & ~n25838;
  assign n26122 = ~n25843 & ~n26121;
  assign n26123 = pi787 & ~n26122;
  assign n26124 = ~pi787 & ~n25835;
  assign n26125 = ~n23547 & ~n26124;
  assign n26126 = ~n26123 & n26125;
  assign n26127 = ~n23557 & ~n23562;
  assign n26128 = n12602 & n25406;
  assign n26129 = ~n26127 & ~n26128;
  assign n26130 = n25486 & n26129;
  assign n26131 = n25406 & ~n26127;
  assign n26132 = n12602 & n26131;
  assign n26133 = n25647 & n26132;
  assign n26134 = ~n26130 & ~n26133;
  assign n26135 = ~n26126 & n26134;
  assign n26136 = ~n26120 & n26135;
  assign n26137 = ~pi790 & ~n26119;
  assign n26138 = ~pi644 & n26119;
  assign n26139 = ~n26123 & ~n26124;
  assign n26140 = pi644 & n26139;
  assign n26141 = ~pi715 & ~n26140;
  assign n26142 = ~n26138 & n26141;
  assign n26143 = ~n7835 & n25655;
  assign n26144 = n7835 & n25486;
  assign n26145 = ~n26143 & ~n26144;
  assign n26146 = ~pi644 & ~n26145;
  assign n26147 = pi644 & n25486;
  assign n26148 = pi715 & ~n26147;
  assign n26149 = ~n26146 & n26148;
  assign n26150 = ~pi1160 & ~n26149;
  assign n26151 = ~n26142 & n26150;
  assign n26152 = pi644 & n26119;
  assign n26153 = ~pi644 & n26139;
  assign n26154 = pi715 & ~n26153;
  assign n26155 = ~n26152 & n26154;
  assign n26156 = pi644 & ~n26145;
  assign n26157 = ~pi644 & n25486;
  assign n26158 = ~pi715 & ~n26157;
  assign n26159 = ~n26156 & n26158;
  assign n26160 = pi1160 & ~n26159;
  assign n26161 = ~n26155 & n26160;
  assign n26162 = pi790 & ~n26161;
  assign n26163 = ~n26151 & n26162;
  assign n26164 = ~n26137 & ~n26163;
  assign n26165 = ~n26136 & ~n26137;
  assign n26166 = n58992 & ~n59967;
  assign n26167 = pi198 & ~n58992;
  assign n26168 = ~n26166 & ~n26167;
  assign n26169 = ~pi223 & ~n59154;
  assign n26170 = ~n6543 & ~n26169;
  assign n26171 = ~pi299 & ~n26170;
  assign n26172 = pi39 & ~n26171;
  assign n26173 = ~n6653 & n26172;
  assign n26174 = ~pi38 & ~n8180;
  assign n26175 = ~n26173 & n26174;
  assign n26176 = n9184 & ~n26175;
  assign n26177 = pi222 & ~n26176;
  assign n26178 = n7597 & ~n26177;
  assign n26179 = pi222 & ~n59132;
  assign n26180 = ~n2680 & n6593;
  assign n26181 = ~n6567 & ~n26180;
  assign n26182 = ~pi616 & ~n26181;
  assign n26183 = pi616 & n7014;
  assign n26184 = pi616 & ~n7014;
  assign n26185 = ~pi616 & n26181;
  assign n26186 = ~n26184 & ~n26185;
  assign n26187 = ~n26182 & ~n26183;
  assign n26188 = ~n6517 & ~n59968;
  assign n26189 = ~n2779 & n59968;
  assign n26190 = pi616 & n6701;
  assign n26191 = n6687 & ~n26190;
  assign n26192 = ~n6685 & ~n26191;
  assign n26193 = n2779 & ~n26192;
  assign n26194 = n6517 & ~n26193;
  assign n26195 = ~n26189 & n26194;
  assign n26196 = ~n26188 & ~n26195;
  assign n26197 = ~n58846 & n26196;
  assign n26198 = pi616 & ~n6702;
  assign n26199 = ~n6594 & ~n26198;
  assign n26200 = ~n6517 & ~n26199;
  assign n26201 = ~n2779 & n26199;
  assign n26202 = n2779 & ~n26190;
  assign n26203 = n6587 & n26202;
  assign n26204 = n6517 & ~n26203;
  assign n26205 = ~n26201 & n26204;
  assign n26206 = ~n26200 & ~n26205;
  assign n26207 = n58846 & n26206;
  assign n26208 = pi222 & ~n26207;
  assign n26209 = ~n26197 & n26208;
  assign n26210 = ~n2781 & ~n6803;
  assign n26211 = ~n2781 & n6803;
  assign n26212 = ~n6810 & ~n26211;
  assign n26213 = ~n6801 & ~n26210;
  assign n26214 = pi616 & ~n59969;
  assign n26215 = n58846 & ~n26214;
  assign n26216 = ~n6568 & n26190;
  assign n26217 = ~n6517 & ~n26216;
  assign n26218 = ~n2779 & n26216;
  assign n26219 = pi616 & n2779;
  assign n26220 = n6904 & n26219;
  assign n26221 = n6517 & ~n26220;
  assign n26222 = ~n26218 & n26221;
  assign n26223 = ~n26217 & ~n26222;
  assign n26224 = ~n58846 & ~n26223;
  assign n26225 = ~pi222 & ~n26224;
  assign n26226 = ~pi222 & ~n26215;
  assign n26227 = ~n26224 & n26226;
  assign n26228 = ~n26215 & n26225;
  assign n26229 = ~n6629 & ~n59970;
  assign n26230 = ~n26209 & n26229;
  assign n26231 = pi222 & ~n6464;
  assign n26232 = n6629 & ~n26231;
  assign n26233 = n6531 & n6701;
  assign n26234 = n26232 & ~n26233;
  assign n26235 = ~pi215 & ~n26234;
  assign n26236 = ~n26230 & n26235;
  assign n26237 = n6504 & n6517;
  assign n26238 = ~n2680 & n26237;
  assign n26239 = n2781 & n6489;
  assign n26240 = ~n6827 & ~n26211;
  assign n26241 = pi616 & ~n26240;
  assign n26242 = n26233 & ~n59971;
  assign n26243 = ~pi222 & n59972;
  assign n26244 = ~n6833 & n26243;
  assign n26245 = ~n6501 & ~n26198;
  assign n26246 = ~n6517 & ~n26245;
  assign n26247 = ~n2779 & n26245;
  assign n26248 = n6490 & n26202;
  assign n26249 = n6517 & ~n26248;
  assign n26250 = ~n26247 & n26249;
  assign n26251 = ~n26246 & ~n26250;
  assign n26252 = n58846 & n26251;
  assign n26253 = pi616 & ~n6731;
  assign n26254 = n6496 & ~n26253;
  assign n26255 = ~n6517 & ~n26254;
  assign n26256 = ~n2779 & ~n6496;
  assign n26257 = ~n6504 & ~n26253;
  assign n26258 = ~n26256 & n26257;
  assign n26259 = n6517 & ~n26258;
  assign n26260 = ~n26255 & ~n26259;
  assign n26261 = ~n58846 & n26260;
  assign n26262 = pi222 & ~n26261;
  assign n26263 = ~n26252 & n26262;
  assign n26264 = ~n26244 & ~n26263;
  assign n26265 = pi215 & ~n26264;
  assign n26266 = pi299 & ~n26265;
  assign n26267 = ~n26236 & n26266;
  assign n26268 = ~n2790 & n26196;
  assign n26269 = n2790 & n26206;
  assign n26270 = pi222 & ~n26269;
  assign n26271 = ~n26268 & n26270;
  assign n26272 = ~n2790 & n26223;
  assign n26273 = n2790 & n26214;
  assign n26274 = pi224 & ~n26273;
  assign n26275 = ~n26272 & n26274;
  assign n26276 = ~pi224 & ~n26233;
  assign n26277 = ~pi222 & ~n26276;
  assign n26278 = ~n26275 & n26277;
  assign n26279 = ~pi223 & ~n26278;
  assign n26280 = ~n26271 & n26279;
  assign n26281 = n2790 & n26251;
  assign n26282 = ~n2790 & n26260;
  assign n26283 = pi222 & ~n26282;
  assign n26284 = ~n26281 & n26283;
  assign n26285 = ~n6848 & n26243;
  assign n26286 = pi223 & ~n26285;
  assign n26287 = ~n26284 & n26286;
  assign n26288 = ~n26280 & ~n26287;
  assign n26289 = ~pi299 & ~n26288;
  assign n26290 = pi39 & ~n26289;
  assign n26291 = pi39 & ~n26267;
  assign n26292 = ~n26289 & n26291;
  assign n26293 = ~n26267 & n26290;
  assign n26294 = pi222 & n59157;
  assign n26295 = ~pi616 & n6798;
  assign n26296 = ~pi222 & ~n6798;
  assign n26297 = ~pi39 & ~n26296;
  assign n26298 = ~pi39 & ~n26295;
  assign n26299 = ~n26296 & n26298;
  assign n26300 = ~n26295 & n26297;
  assign n26301 = ~n26294 & n59974;
  assign n26302 = ~pi38 & ~n26301;
  assign n26303 = ~n59973 & n26302;
  assign n26304 = pi222 & ~n6863;
  assign n26305 = pi38 & ~n26304;
  assign n26306 = n6863 & n26190;
  assign n26307 = pi616 & n6865;
  assign n26308 = n26305 & ~n59975;
  assign n26309 = n59132 & ~n26308;
  assign n26310 = ~n26303 & n26309;
  assign n26311 = ~n26179 & ~n26310;
  assign n26312 = ~n7597 & n26311;
  assign n26313 = ~n7597 & ~n26311;
  assign n26314 = n7597 & n26177;
  assign n26315 = ~n26313 & ~n26314;
  assign n26316 = ~n26178 & ~n26312;
  assign n26317 = ~pi785 & ~n59976;
  assign n26318 = pi609 & n59976;
  assign n26319 = ~pi609 & ~n26177;
  assign n26320 = pi1155 & ~n26319;
  assign n26321 = ~n26318 & n26320;
  assign n26322 = ~pi609 & n59976;
  assign n26323 = pi609 & ~n26177;
  assign n26324 = ~pi1155 & ~n26323;
  assign n26325 = ~n26322 & n26324;
  assign n26326 = ~n26321 & ~n26325;
  assign n26327 = pi785 & ~n26326;
  assign n26328 = ~n26317 & ~n26327;
  assign n26329 = ~pi781 & ~n26328;
  assign n26330 = pi618 & n26328;
  assign n26331 = ~pi618 & ~n26177;
  assign n26332 = pi1154 & ~n26331;
  assign n26333 = ~n26330 & n26332;
  assign n26334 = ~pi618 & n26328;
  assign n26335 = pi618 & ~n26177;
  assign n26336 = ~pi1154 & ~n26335;
  assign n26337 = ~n26334 & n26336;
  assign n26338 = ~n26333 & ~n26337;
  assign n26339 = pi781 & ~n26338;
  assign n26340 = ~n26329 & ~n26339;
  assign n26341 = ~pi789 & ~n26340;
  assign n26342 = pi619 & n26340;
  assign n26343 = ~pi619 & ~n26177;
  assign n26344 = pi1159 & ~n26343;
  assign n26345 = ~n26342 & n26344;
  assign n26346 = ~pi619 & n26340;
  assign n26347 = pi619 & ~n26177;
  assign n26348 = ~pi1159 & ~n26347;
  assign n26349 = ~n26346 & n26348;
  assign n26350 = ~n26345 & ~n26349;
  assign n26351 = pi789 & ~n26350;
  assign n26352 = ~n26341 & ~n26351;
  assign n26353 = ~n8054 & ~n26352;
  assign n26354 = n8054 & n26177;
  assign n26355 = n8054 & ~n26177;
  assign n26356 = ~n8054 & n26352;
  assign n26357 = ~n26355 & ~n26356;
  assign n26358 = ~n26353 & ~n26354;
  assign n26359 = ~n11154 & n59977;
  assign n26360 = ~n9651 & ~n26177;
  assign n26361 = n59229 & ~n26177;
  assign n26362 = ~pi222 & ~n7327;
  assign n26363 = pi661 & pi680;
  assign n26364 = n7327 & ~n26363;
  assign n26365 = pi222 & n7304;
  assign n26366 = pi299 & ~n26365;
  assign n26367 = ~n26364 & n26366;
  assign n26368 = ~n26362 & n26366;
  assign n26369 = ~n26364 & n26368;
  assign n26370 = ~n26362 & n26367;
  assign n26371 = ~pi222 & ~n7318;
  assign n26372 = n7318 & ~n26363;
  assign n26373 = pi222 & n7298;
  assign n26374 = ~pi299 & ~n26373;
  assign n26375 = ~n26372 & n26374;
  assign n26376 = ~n26371 & n26374;
  assign n26377 = ~n26372 & n26376;
  assign n26378 = ~n26371 & n26375;
  assign n26379 = ~pi39 & ~n59979;
  assign n26380 = ~pi39 & ~n59978;
  assign n26381 = ~n59979 & n26380;
  assign n26382 = ~n59978 & n26379;
  assign n26383 = pi661 & ~n7418;
  assign n26384 = ~pi661 & n6596;
  assign n26385 = ~n2779 & ~n6595;
  assign n26386 = ~pi662 & n6606;
  assign n26387 = ~n26385 & ~n26386;
  assign n26388 = n6517 & ~n26387;
  assign n26389 = ~n26384 & ~n26388;
  assign n26390 = ~n26383 & n26389;
  assign n26391 = n2790 & n26390;
  assign n26392 = ~pi661 & ~n59152;
  assign n26393 = pi680 & n7209;
  assign n26394 = ~n6903 & ~n26393;
  assign n26395 = pi661 & ~n26394;
  assign n26396 = ~n26392 & ~n26395;
  assign n26397 = ~n2790 & n26396;
  assign n26398 = pi222 & ~n26397;
  assign n26399 = ~n26391 & n26398;
  assign n26400 = ~n7495 & n26363;
  assign n26401 = n2790 & n26400;
  assign n26402 = pi661 & n7490;
  assign n26403 = ~n2790 & n26402;
  assign n26404 = pi224 & ~n26403;
  assign n26405 = pi224 & ~n26401;
  assign n26406 = ~n26403 & n26405;
  assign n26407 = ~n26401 & n26404;
  assign n26408 = pi661 & n59222;
  assign n26409 = n7035 & n26363;
  assign n26410 = ~pi224 & ~n59982;
  assign n26411 = ~pi222 & ~n26410;
  assign n26412 = ~n59981 & n26411;
  assign n26413 = ~pi223 & ~n26412;
  assign n26414 = ~n26399 & n26413;
  assign n26415 = ~pi661 & ~n59149;
  assign n26416 = pi661 & ~n7440;
  assign n26417 = ~n26415 & ~n26416;
  assign n26418 = n2790 & n26417;
  assign n26419 = n6507 & n6517;
  assign n26420 = ~pi661 & n6497;
  assign n26421 = pi661 & ~n7445;
  assign n26422 = ~n26420 & ~n26421;
  assign n26423 = ~n26419 & n26422;
  assign n26424 = ~n2790 & n26423;
  assign n26425 = pi222 & ~n26424;
  assign n26426 = ~n26418 & n26425;
  assign n26427 = ~pi222 & pi661;
  assign n26428 = n7508 & n26427;
  assign n26429 = pi223 & ~n26428;
  assign n26430 = ~n26426 & n26429;
  assign n26431 = ~n26414 & ~n26430;
  assign n26432 = ~pi299 & ~n26431;
  assign n26433 = n58846 & n26390;
  assign n26434 = ~n58846 & n26396;
  assign n26435 = pi222 & ~n26434;
  assign n26436 = ~n26433 & n26435;
  assign n26437 = ~n58846 & ~n26402;
  assign n26438 = n58846 & ~n26400;
  assign n26439 = ~pi222 & ~n26438;
  assign n26440 = ~pi222 & ~n26437;
  assign n26441 = ~n26438 & n26440;
  assign n26442 = ~n26437 & n26439;
  assign n26443 = ~n6629 & ~n59983;
  assign n26444 = ~n26436 & n26443;
  assign n26445 = n26232 & ~n59982;
  assign n26446 = ~pi215 & ~n26445;
  assign n26447 = ~n26444 & n26446;
  assign n26448 = n7531 & n26427;
  assign n26449 = n58846 & n26417;
  assign n26450 = ~n58846 & n26423;
  assign n26451 = pi222 & ~n26450;
  assign n26452 = ~n26449 & n26451;
  assign n26453 = ~n26448 & ~n26452;
  assign n26454 = pi215 & ~n26453;
  assign n26455 = pi299 & ~n26454;
  assign n26456 = ~n26447 & n26455;
  assign n26457 = ~n26432 & ~n26456;
  assign n26458 = pi39 & ~n26457;
  assign n26459 = ~n59980 & ~n26458;
  assign n26460 = ~pi38 & ~n26459;
  assign n26461 = pi661 & n7546;
  assign n26462 = n26305 & ~n26461;
  assign n26463 = n59132 & ~n26462;
  assign n26464 = ~n26460 & n26463;
  assign n26465 = ~n26179 & ~n26464;
  assign n26466 = ~pi778 & ~n26465;
  assign n26467 = pi625 & n26465;
  assign n26468 = ~pi625 & ~n26177;
  assign n26469 = pi1153 & ~n26468;
  assign n26470 = ~n26467 & n26469;
  assign n26471 = ~pi625 & n26465;
  assign n26472 = pi625 & ~n26177;
  assign n26473 = ~pi1153 & ~n26472;
  assign n26474 = ~n26471 & n26473;
  assign n26475 = ~n26470 & ~n26474;
  assign n26476 = pi778 & ~n26475;
  assign n26477 = ~n26466 & ~n26476;
  assign n26478 = ~n59229 & n26477;
  assign n26479 = ~n59229 & ~n26477;
  assign n26480 = n59229 & n26177;
  assign n26481 = ~n26479 & ~n26480;
  assign n26482 = ~n26361 & ~n26478;
  assign n26483 = ~n59231 & n59984;
  assign n26484 = n59231 & ~n26177;
  assign n26485 = ~n59231 & ~n59984;
  assign n26486 = n59231 & n26177;
  assign n26487 = ~n26485 & ~n26486;
  assign n26488 = ~n26483 & ~n26484;
  assign n26489 = ~n7716 & n59985;
  assign n26490 = ~n7762 & n26489;
  assign n26491 = ~n26360 & ~n26490;
  assign n26492 = ~pi628 & ~n26491;
  assign n26493 = pi628 & ~n26177;
  assign n26494 = n7791 & ~n26493;
  assign n26495 = ~n26492 & n26494;
  assign n26496 = pi628 & ~n26491;
  assign n26497 = ~pi628 & ~n26177;
  assign n26498 = n7790 & ~n26497;
  assign n26499 = ~n26496 & n26498;
  assign n26500 = ~n26495 & ~n26499;
  assign n26501 = ~n26359 & n26500;
  assign n26502 = pi792 & ~n26501;
  assign n26503 = ~pi680 & n26199;
  assign n26504 = pi616 & ~n7192;
  assign n26505 = pi680 & ~n26504;
  assign n26506 = ~n6883 & n26505;
  assign n26507 = pi661 & ~n26506;
  assign n26508 = pi661 & ~n26503;
  assign n26509 = ~n26506 & n26508;
  assign n26510 = ~n26503 & n26507;
  assign n26511 = ~pi661 & pi681;
  assign n26512 = ~n26199 & n26511;
  assign n26513 = ~n26205 & ~n26512;
  assign n26514 = ~n59986 & n26513;
  assign n26515 = pi222 & ~n26514;
  assign n26516 = pi616 & ~n7132;
  assign n26517 = pi680 & ~n7047;
  assign n26518 = ~n26516 & n26517;
  assign n26519 = ~pi680 & n26233;
  assign n26520 = pi661 & ~n26519;
  assign n26521 = ~n26518 & n26520;
  assign n26522 = ~pi661 & ~n26233;
  assign n26523 = ~n2781 & ~n26522;
  assign n26524 = ~pi681 & n26219;
  assign n26525 = n6800 & n26524;
  assign n26526 = n6800 & n26219;
  assign n26527 = ~n2779 & n26233;
  assign n26528 = n6517 & ~n26527;
  assign n26529 = ~n26526 & n26528;
  assign n26530 = ~n26233 & n26511;
  assign n26531 = ~n26529 & ~n26530;
  assign n26532 = ~n26523 & ~n26525;
  assign n26533 = ~n26521 & n59987;
  assign n26534 = ~pi222 & n26533;
  assign n26535 = n58846 & ~n26534;
  assign n26536 = ~n26515 & n26535;
  assign n26537 = ~pi680 & n59968;
  assign n26538 = n2680 & n6889;
  assign n26539 = ~n6922 & ~n26538;
  assign n26540 = n6872 & ~n7010;
  assign n26541 = ~pi603 & n59988;
  assign n26542 = pi603 & n6566;
  assign n26543 = ~n6894 & ~n26542;
  assign n26544 = ~n26541 & n26543;
  assign n26545 = ~pi642 & n26544;
  assign n26546 = ~n7117 & n59988;
  assign n26547 = pi642 & ~n26546;
  assign n26548 = n2777 & ~n26547;
  assign n26549 = n2777 & ~n26545;
  assign n26550 = ~n26547 & n26549;
  assign n26551 = ~n26545 & n26548;
  assign n26552 = n7067 & n26546;
  assign n26553 = n7131 & ~n59988;
  assign n26554 = ~n7010 & n7131;
  assign n26555 = pi616 & ~n59990;
  assign n26556 = pi680 & ~n26555;
  assign n26557 = ~n26552 & n26556;
  assign n26558 = ~n59989 & n26557;
  assign n26559 = pi661 & ~n26558;
  assign n26560 = ~n26537 & n26559;
  assign n26561 = ~n59968 & n26511;
  assign n26562 = ~n26195 & ~n26561;
  assign n26563 = ~n26560 & n26562;
  assign n26564 = pi222 & ~n26563;
  assign n26565 = pi616 & n7118;
  assign n26566 = pi680 & ~n26565;
  assign n26567 = ~n59181 & n26566;
  assign n26568 = ~pi680 & n26216;
  assign n26569 = pi661 & ~n26568;
  assign n26570 = ~n26567 & n26569;
  assign n26571 = ~n26216 & n26511;
  assign n26572 = ~n26222 & ~n26571;
  assign n26573 = ~n26570 & n26572;
  assign n26574 = ~pi222 & n26573;
  assign n26575 = ~n58846 & ~n26574;
  assign n26576 = ~n26564 & n26575;
  assign n26577 = ~n58846 & ~n26563;
  assign n26578 = n58846 & ~n26514;
  assign n26579 = pi222 & ~n26578;
  assign n26580 = ~n26577 & n26579;
  assign n26581 = ~n58846 & n26573;
  assign n26582 = n58846 & n26533;
  assign n26583 = ~pi222 & ~n26582;
  assign n26584 = ~n26581 & n26583;
  assign n26585 = ~n26580 & ~n26584;
  assign n26586 = ~n26536 & ~n26576;
  assign n26587 = ~n6629 & ~n59991;
  assign n26588 = ~n26190 & ~n26363;
  assign n26589 = ~pi616 & ~n59182;
  assign n26590 = ~n26516 & ~n26589;
  assign n26591 = ~n26588 & n26590;
  assign n26592 = n26232 & ~n26591;
  assign n26593 = ~pi215 & ~n26592;
  assign n26594 = ~n26587 & n26593;
  assign n26595 = ~n6933 & n26505;
  assign n26596 = ~pi680 & n26245;
  assign n26597 = pi661 & ~n26596;
  assign n26598 = ~n26595 & n26597;
  assign n26599 = ~n26245 & n26511;
  assign n26600 = ~n26250 & ~n26599;
  assign n26601 = ~n26598 & n26600;
  assign n26602 = n58846 & ~n26601;
  assign n26603 = ~pi680 & n26254;
  assign n26604 = ~n6943 & n7131;
  assign n26605 = pi616 & ~n26604;
  assign n26606 = pi680 & ~n26605;
  assign n26607 = n6947 & n26606;
  assign n26608 = pi661 & ~n26607;
  assign n26609 = ~n26603 & n26608;
  assign n26610 = ~n26254 & n26511;
  assign n26611 = ~n26259 & ~n26610;
  assign n26612 = ~n26609 & n26611;
  assign n26613 = ~n58846 & ~n26612;
  assign n26614 = pi222 & ~n26613;
  assign n26615 = pi222 & ~n26602;
  assign n26616 = ~n26613 & n26615;
  assign n26617 = ~n26602 & n26614;
  assign n26618 = ~n6828 & ~n7169;
  assign n26619 = pi616 & n26618;
  assign n26620 = pi680 & ~n26619;
  assign n26621 = n59184 & n26620;
  assign n26622 = pi616 & n6828;
  assign n26623 = ~n6486 & n26233;
  assign n26624 = ~pi680 & n59993;
  assign n26625 = pi661 & ~n26624;
  assign n26626 = ~n26621 & n26625;
  assign n26627 = ~pi661 & ~n59993;
  assign n26628 = pi616 & n6920;
  assign n26629 = ~n6484 & n26233;
  assign n26630 = n2781 & ~n59994;
  assign n26631 = ~n26627 & ~n26630;
  assign n26632 = ~n26626 & n26631;
  assign n26633 = ~n58846 & n26632;
  assign n26634 = n7081 & n26363;
  assign n26635 = ~n59972 & ~n26634;
  assign n26636 = n58846 & ~n26635;
  assign n26637 = ~pi222 & ~n26636;
  assign n26638 = ~n26633 & n26637;
  assign n26639 = pi215 & ~n26638;
  assign n26640 = ~n59992 & n26639;
  assign n26641 = pi299 & ~n26640;
  assign n26642 = ~n26594 & n26641;
  assign n26643 = ~n2790 & n26573;
  assign n26644 = n2790 & n26533;
  assign n26645 = pi224 & ~n26644;
  assign n26646 = ~n26643 & n26645;
  assign n26647 = n26363 & n26590;
  assign n26648 = n26233 & ~n26363;
  assign n26649 = ~pi224 & ~n26648;
  assign n26650 = ~n26647 & n26649;
  assign n26651 = ~pi222 & pi224;
  assign n26652 = n26363 & ~n26590;
  assign n26653 = ~n26233 & ~n26363;
  assign n26654 = ~pi222 & ~n26653;
  assign n26655 = ~n26652 & n26654;
  assign n26656 = ~n26651 & ~n26655;
  assign n26657 = ~pi222 & ~n26650;
  assign n26658 = ~n26646 & ~n59995;
  assign n26659 = ~n2790 & n26563;
  assign n26660 = n2790 & n26514;
  assign n26661 = pi222 & ~n26660;
  assign n26662 = ~n26659 & n26661;
  assign n26663 = ~n26658 & ~n26662;
  assign n26664 = ~pi223 & ~n26663;
  assign n26665 = n2790 & ~n26601;
  assign n26666 = ~n2790 & ~n26612;
  assign n26667 = pi222 & ~n26666;
  assign n26668 = pi222 & ~n26665;
  assign n26669 = ~n26666 & n26668;
  assign n26670 = ~n26665 & n26667;
  assign n26671 = ~n2790 & n26632;
  assign n26672 = n2790 & ~n26635;
  assign n26673 = ~pi222 & ~n26672;
  assign n26674 = ~n26671 & n26673;
  assign n26675 = pi223 & ~n26674;
  assign n26676 = ~n59996 & n26675;
  assign n26677 = ~pi299 & ~n26676;
  assign n26678 = ~n26664 & n26677;
  assign n26679 = pi39 & ~n26678;
  assign n26680 = ~n26642 & n26679;
  assign n26681 = pi661 & n7323;
  assign n26682 = pi616 & n6791;
  assign n26683 = ~pi222 & ~n26682;
  assign n26684 = ~n26681 & n26683;
  assign n26685 = n7322 & ~n26363;
  assign n26686 = ~pi603 & ~n7298;
  assign n26687 = ~n6893 & ~n7320;
  assign n26688 = ~n26686 & n26687;
  assign n26689 = ~pi616 & n6791;
  assign n26690 = ~n26688 & ~n26689;
  assign n26691 = ~n26685 & n26690;
  assign n26692 = pi222 & ~n26691;
  assign n26693 = ~pi299 & ~n26692;
  assign n26694 = ~n26684 & n26693;
  assign n26695 = pi661 & n7331;
  assign n26696 = pi616 & n6796;
  assign n26697 = ~pi222 & ~n26696;
  assign n26698 = ~n26695 & n26697;
  assign n26699 = n7330 & ~n26363;
  assign n26700 = ~pi603 & ~n7304;
  assign n26701 = ~n6676 & ~n6893;
  assign n26702 = ~n26700 & n26701;
  assign n26703 = ~pi616 & n6796;
  assign n26704 = ~n26702 & ~n26703;
  assign n26705 = ~n26699 & n26704;
  assign n26706 = pi222 & ~n26705;
  assign n26707 = pi299 & ~n26706;
  assign n26708 = ~n26698 & n26707;
  assign n26709 = ~n26694 & ~n26708;
  assign n26710 = ~n26698 & ~n26706;
  assign n26711 = pi299 & ~n26710;
  assign n26712 = ~n26684 & ~n26692;
  assign n26713 = ~pi299 & ~n26712;
  assign n26714 = ~pi39 & ~n26713;
  assign n26715 = ~n26711 & n26714;
  assign n26716 = ~pi39 & ~n26709;
  assign n26717 = ~pi38 & ~n59997;
  assign n26718 = ~n26680 & n26717;
  assign n26719 = n6468 & n7131;
  assign n26720 = ~pi222 & ~pi616;
  assign n26721 = ~pi39 & pi616;
  assign n26722 = n26363 & n26721;
  assign n26723 = ~n26720 & ~n26722;
  assign n26724 = n26719 & ~n26723;
  assign n26725 = ~pi616 & ~n6914;
  assign n26726 = ~n26588 & ~n26725;
  assign n26727 = n6863 & n26726;
  assign n26728 = ~n26304 & ~n26727;
  assign n26729 = ~n26724 & ~n26728;
  assign n26730 = pi38 & ~n26729;
  assign n26731 = n59132 & ~n26730;
  assign n26732 = ~n26718 & n26731;
  assign n26733 = ~n26179 & ~n26732;
  assign n26734 = ~pi625 & n26733;
  assign n26735 = pi625 & n26311;
  assign n26736 = ~pi1153 & ~n26735;
  assign n26737 = ~n26734 & n26736;
  assign n26738 = ~pi608 & ~n26470;
  assign n26739 = ~n26737 & n26738;
  assign n26740 = pi625 & n26733;
  assign n26741 = ~pi625 & n26311;
  assign n26742 = pi1153 & ~n26741;
  assign n26743 = ~n26740 & n26742;
  assign n26744 = pi608 & ~n26474;
  assign n26745 = ~n26743 & n26744;
  assign n26746 = ~n26739 & ~n26745;
  assign n26747 = pi778 & ~n26746;
  assign n26748 = ~pi778 & n26733;
  assign n26749 = ~n26747 & ~n26748;
  assign n26750 = ~pi609 & ~n26749;
  assign n26751 = pi609 & n26477;
  assign n26752 = ~pi1155 & ~n26751;
  assign n26753 = ~n26750 & n26752;
  assign n26754 = ~pi660 & ~n26321;
  assign n26755 = ~n26753 & n26754;
  assign n26756 = pi609 & ~n26749;
  assign n26757 = ~pi609 & n26477;
  assign n26758 = pi1155 & ~n26757;
  assign n26759 = ~n26756 & n26758;
  assign n26760 = pi660 & ~n26325;
  assign n26761 = ~n26759 & n26760;
  assign n26762 = ~n26755 & ~n26761;
  assign n26763 = pi785 & ~n26762;
  assign n26764 = ~pi785 & ~n26749;
  assign n26765 = ~n26763 & ~n26764;
  assign n26766 = ~pi618 & ~n26765;
  assign n26767 = pi618 & n59984;
  assign n26768 = ~pi1154 & ~n26767;
  assign n26769 = ~n26766 & n26768;
  assign n26770 = ~pi627 & ~n26333;
  assign n26771 = ~n26769 & n26770;
  assign n26772 = pi618 & ~n26765;
  assign n26773 = ~pi618 & n59984;
  assign n26774 = pi1154 & ~n26773;
  assign n26775 = ~n26772 & n26774;
  assign n26776 = pi627 & ~n26337;
  assign n26777 = ~n26775 & n26776;
  assign n26778 = ~n26771 & ~n26777;
  assign n26779 = pi781 & ~n26778;
  assign n26780 = ~pi781 & ~n26765;
  assign n26781 = ~n26779 & ~n26780;
  assign n26782 = ~pi619 & ~n26781;
  assign n26783 = pi619 & n59985;
  assign n26784 = ~pi1159 & ~n26783;
  assign n26785 = ~n26782 & n26784;
  assign n26786 = ~pi648 & ~n26345;
  assign n26787 = ~n26785 & n26786;
  assign n26788 = pi619 & ~n26781;
  assign n26789 = ~pi619 & n59985;
  assign n26790 = pi1159 & ~n26789;
  assign n26791 = ~n26788 & n26790;
  assign n26792 = pi648 & ~n26349;
  assign n26793 = ~n26791 & n26792;
  assign n26794 = pi789 & ~n26793;
  assign n26795 = pi789 & ~n26787;
  assign n26796 = ~n26793 & n26795;
  assign n26797 = ~n26787 & n26794;
  assign n26798 = pi626 & n26352;
  assign n26799 = ~pi626 & ~n26177;
  assign n26800 = n7759 & ~n26799;
  assign n26801 = ~n26798 & n26800;
  assign n26802 = ~pi626 & n26352;
  assign n26803 = pi626 & ~n26177;
  assign n26804 = n7760 & ~n26803;
  assign n26805 = ~n26802 & n26804;
  assign n26806 = n7716 & ~n26177;
  assign n26807 = n7984 & ~n26806;
  assign n26808 = ~n26489 & n26807;
  assign n26809 = ~n26805 & ~n26808;
  assign n26810 = ~n26801 & ~n26808;
  assign n26811 = ~n26805 & n26810;
  assign n26812 = ~n26801 & n26809;
  assign n26813 = pi788 & ~n59999;
  assign n26814 = ~pi789 & n26781;
  assign n26815 = ~n26813 & ~n26814;
  assign n26816 = ~n59998 & n26815;
  assign n26817 = ~n59242 & n59999;
  assign n26818 = ~n59357 & ~n26817;
  assign n26819 = ~n26816 & n26818;
  assign n26820 = ~n26502 & ~n26819;
  assign n26821 = ~n8108 & ~n26820;
  assign n26822 = ~n7793 & ~n59977;
  assign n26823 = n7793 & ~n26177;
  assign n26824 = ~n7872 & ~n26823;
  assign n26825 = ~n7793 & n59977;
  assign n26826 = n7793 & n26177;
  assign n26827 = ~n26825 & ~n26826;
  assign n26828 = ~n7872 & ~n26827;
  assign n26829 = ~n26822 & n26824;
  assign n26830 = ~n59240 & n26491;
  assign n26831 = n59240 & n26177;
  assign n26832 = ~n59240 & ~n26491;
  assign n26833 = n59240 & ~n26177;
  assign n26834 = ~n26832 & ~n26833;
  assign n26835 = ~n26830 & ~n26831;
  assign n26836 = pi647 & ~n60001;
  assign n26837 = ~pi647 & ~n26177;
  assign n26838 = pi1157 & ~n26837;
  assign n26839 = ~n26836 & n26838;
  assign n26840 = ~pi630 & n26839;
  assign n26841 = ~pi647 & ~n60001;
  assign n26842 = pi647 & ~n26177;
  assign n26843 = ~pi1157 & ~n26842;
  assign n26844 = ~n26841 & n26843;
  assign n26845 = pi630 & n26844;
  assign n26846 = ~n26840 & ~n26845;
  assign n26847 = ~n60000 & n26846;
  assign n26848 = pi787 & ~n26847;
  assign n26849 = ~n26821 & ~n26848;
  assign n26850 = ~n23537 & ~n26849;
  assign n26851 = n12602 & ~n26352;
  assign n26852 = n23562 & n26851;
  assign n26853 = n23557 & n26177;
  assign n26854 = ~n26852 & ~n26853;
  assign n26855 = ~pi644 & ~n26854;
  assign n26856 = n23557 & n26851;
  assign n26857 = n23562 & n26177;
  assign n26858 = ~n26856 & ~n26857;
  assign n26859 = pi644 & ~n26858;
  assign n26860 = ~n12602 & ~n26127;
  assign n26861 = n26177 & n26860;
  assign n26862 = pi787 & ~n26839;
  assign n26863 = ~n26844 & n26862;
  assign n26864 = ~pi787 & ~n60001;
  assign n26865 = ~n23547 & ~n26864;
  assign n26866 = ~n26863 & n26865;
  assign n26867 = ~n26861 & ~n26866;
  assign n26868 = ~n26859 & n26867;
  assign n26869 = ~n26855 & n26868;
  assign n26870 = pi790 & ~n26869;
  assign n26871 = ~pi644 & n26849;
  assign n26872 = ~pi787 & n60001;
  assign n26873 = ~n26839 & ~n26844;
  assign n26874 = pi787 & ~n26873;
  assign n26875 = ~n26872 & ~n26874;
  assign n26876 = pi644 & n26875;
  assign n26877 = ~pi715 & ~n26876;
  assign n26878 = ~n26871 & n26877;
  assign n26879 = n7835 & ~n26177;
  assign n26880 = ~n7835 & n26827;
  assign n26881 = ~n26879 & ~n26880;
  assign n26882 = ~pi644 & ~n26881;
  assign n26883 = pi644 & ~n26177;
  assign n26884 = pi715 & ~n26883;
  assign n26885 = ~n26882 & n26884;
  assign n26886 = ~pi1160 & ~n26885;
  assign n26887 = ~n26878 & n26886;
  assign n26888 = pi644 & n26849;
  assign n26889 = ~pi644 & n26875;
  assign n26890 = pi715 & ~n26889;
  assign n26891 = ~n26888 & n26890;
  assign n26892 = pi644 & ~n26881;
  assign n26893 = ~pi644 & ~n26177;
  assign n26894 = ~pi715 & ~n26893;
  assign n26895 = ~n26892 & n26894;
  assign n26896 = pi1160 & ~n26895;
  assign n26897 = ~n26891 & n26896;
  assign n26898 = ~n26887 & ~n26897;
  assign n26899 = pi790 & ~n26898;
  assign n26900 = ~pi790 & n26849;
  assign n26901 = ~n26899 & ~n26900;
  assign n26902 = ~n26850 & ~n26870;
  assign n26903 = n58992 & n60002;
  assign n26904 = pi222 & ~n58992;
  assign n26905 = n58992 & ~n60002;
  assign n26906 = ~pi222 & ~n58992;
  assign n26907 = ~n26905 & ~n26906;
  assign n26908 = ~n26903 & ~n26904;
  assign n26909 = pi223 & ~n59132;
  assign n26910 = ~pi223 & pi642;
  assign n26911 = n6791 & n26910;
  assign n26912 = ~pi299 & ~n26911;
  assign n26913 = ~pi642 & n6791;
  assign n26914 = pi223 & ~n26913;
  assign n26915 = n6671 & n26914;
  assign n26916 = n26912 & ~n26915;
  assign n26917 = n6796 & n26910;
  assign n26918 = pi299 & ~n26917;
  assign n26919 = n2776 & n6795;
  assign n26920 = pi223 & ~n26919;
  assign n26921 = pi223 & ~n6677;
  assign n26922 = ~n26919 & n26921;
  assign n26923 = ~n6677 & n26920;
  assign n26924 = n26918 & ~n60004;
  assign n26925 = ~pi39 & ~n26924;
  assign n26926 = ~n26916 & n26925;
  assign n26927 = ~n2777 & n6464;
  assign n26928 = pi642 & n6701;
  assign n26929 = n26927 & ~n26928;
  assign n26930 = pi642 & ~n6702;
  assign n26931 = n2777 & ~n26930;
  assign n26932 = ~n6590 & n26931;
  assign n26933 = ~n26929 & ~n26932;
  assign n26934 = pi681 & n26933;
  assign n26935 = ~n2780 & ~n26933;
  assign n26936 = ~pi642 & n6587;
  assign n26937 = ~n6697 & ~n26936;
  assign n26938 = n2780 & ~n26937;
  assign n26939 = ~pi681 & ~n26938;
  assign n26940 = ~n26935 & n26939;
  assign n26941 = n58846 & ~n26940;
  assign n26942 = ~n26934 & n26941;
  assign n26943 = pi642 & ~n7014;
  assign n26944 = ~pi642 & n59151;
  assign n26945 = ~n26943 & ~n26944;
  assign n26946 = pi681 & ~n26945;
  assign n26947 = ~n2780 & n26945;
  assign n26948 = n6578 & ~n26928;
  assign n26949 = ~pi681 & ~n26948;
  assign n26950 = ~n26947 & n26949;
  assign n26951 = ~n58846 & ~n26950;
  assign n26952 = ~n26946 & n26951;
  assign n26953 = pi223 & ~n26952;
  assign n26954 = ~n26942 & n26953;
  assign n26955 = ~n6568 & n26928;
  assign n26956 = pi681 & ~n26955;
  assign n26957 = ~n2780 & n26955;
  assign n26958 = pi642 & n2780;
  assign n26959 = n6904 & n26958;
  assign n26960 = ~pi681 & ~n26959;
  assign n26961 = ~n26957 & n26960;
  assign n26962 = ~n26956 & ~n26961;
  assign n26963 = ~n2841 & n26962;
  assign n26964 = pi642 & n6803;
  assign n26965 = ~n2780 & n26964;
  assign n26966 = ~pi681 & ~n26965;
  assign n26967 = n6800 & n26958;
  assign n26968 = n26966 & ~n26967;
  assign n26969 = pi681 & ~n26964;
  assign n26970 = ~n26968 & ~n26969;
  assign n26971 = n2841 & n26970;
  assign n26972 = ~pi947 & ~n26971;
  assign n26973 = ~n26963 & n26972;
  assign n26974 = pi947 & ~n26962;
  assign n26975 = ~pi223 & ~n26974;
  assign n26976 = ~n26973 & n26975;
  assign n26977 = ~n6629 & ~n26976;
  assign n26978 = ~n26954 & n26977;
  assign n26979 = pi223 & ~n6464;
  assign n26980 = n6629 & ~n26979;
  assign n26981 = ~n26964 & n26980;
  assign n26982 = ~pi215 & ~n26981;
  assign n26983 = ~n26978 & n26982;
  assign n26984 = n6827 & n26958;
  assign n26985 = n26966 & ~n26984;
  assign n26986 = pi642 & ~n6731;
  assign n26987 = n2780 & ~n26986;
  assign n26988 = ~n6484 & n26987;
  assign n26989 = ~pi681 & ~n26988;
  assign n26990 = n6486 & n26989;
  assign n26991 = ~n26985 & ~n26990;
  assign n26992 = pi642 & n6828;
  assign n26993 = pi681 & ~n26992;
  assign n26994 = n26991 & ~n26993;
  assign n26995 = ~n2841 & n26994;
  assign n26996 = n58846 & ~n26985;
  assign n26997 = n26964 & n26996;
  assign n26998 = ~pi947 & ~n26997;
  assign n26999 = ~n26995 & n26998;
  assign n27000 = pi947 & ~n26994;
  assign n27001 = ~pi223 & ~n27000;
  assign n27002 = ~n26999 & n27001;
  assign n27003 = n26245 & ~n26930;
  assign n27004 = ~n26929 & ~n27003;
  assign n27005 = pi681 & n27004;
  assign n27006 = ~n2780 & ~n27004;
  assign n27007 = n6468 & ~n26928;
  assign n27008 = n2780 & n27007;
  assign n27009 = n6490 & n27008;
  assign n27010 = ~pi681 & ~n27009;
  assign n27011 = ~n27006 & n27010;
  assign n27012 = ~n27005 & ~n27011;
  assign n27013 = n58846 & n27012;
  assign n27014 = ~n6492 & n6700;
  assign n27015 = ~n6486 & ~n26986;
  assign n27016 = ~pi642 & ~n6496;
  assign n27017 = pi642 & ~n6732;
  assign n27018 = ~n27016 & ~n27017;
  assign n27019 = ~n27014 & n27015;
  assign n27020 = ~n2780 & n60005;
  assign n27021 = n26989 & ~n27020;
  assign n27022 = pi681 & ~n60005;
  assign n27023 = ~n27021 & ~n27022;
  assign n27024 = ~n58846 & n27023;
  assign n27025 = pi223 & ~n27024;
  assign n27026 = ~n27013 & n27025;
  assign n27027 = ~n27002 & ~n27026;
  assign n27028 = pi215 & ~n27027;
  assign n27029 = pi299 & ~n27028;
  assign n27030 = ~n26983 & n27029;
  assign n27031 = ~n2790 & n26962;
  assign n27032 = n2790 & n26970;
  assign n27033 = ~n6544 & ~n27032;
  assign n27034 = ~n27031 & n27033;
  assign n27035 = n6544 & ~n26964;
  assign n27036 = ~pi223 & ~n27035;
  assign n27037 = ~n27034 & n27036;
  assign n27038 = n2790 & n27012;
  assign n27039 = ~n2790 & n27023;
  assign n27040 = pi223 & ~n27039;
  assign n27041 = ~n27038 & n27040;
  assign n27042 = ~pi299 & ~n27041;
  assign n27043 = ~n27037 & n27042;
  assign n27044 = pi39 & ~n27043;
  assign n27045 = ~n27030 & n27044;
  assign n27046 = ~pi38 & ~n27045;
  assign n27047 = ~pi38 & ~n26926;
  assign n27048 = ~n27045 & n27047;
  assign n27049 = ~n26926 & n27046;
  assign n27050 = pi39 & pi223;
  assign n27051 = pi38 & ~n27050;
  assign n27052 = ~pi223 & ~n6468;
  assign n27053 = ~pi39 & ~n27052;
  assign n27054 = ~n27007 & n27053;
  assign n27055 = n27051 & ~n27054;
  assign n27056 = n59132 & ~n27055;
  assign n27057 = ~n60006 & n27056;
  assign n27058 = ~n26909 & ~n27057;
  assign n27059 = ~n7597 & ~n27058;
  assign n27060 = ~pi299 & ~n59150;
  assign n27061 = pi39 & ~n27060;
  assign n27062 = ~n6653 & n27061;
  assign n27063 = ~n8180 & n59292;
  assign n27064 = ~n27062 & n27063;
  assign n27065 = n9184 & ~n27064;
  assign n27066 = pi223 & ~n27065;
  assign n27067 = n7597 & n27066;
  assign n27068 = n7597 & ~n27066;
  assign n27069 = ~n7597 & n27058;
  assign n27070 = ~n27068 & ~n27069;
  assign n27071 = ~n27059 & ~n27067;
  assign n27072 = ~pi785 & n60007;
  assign n27073 = pi609 & ~n60007;
  assign n27074 = ~pi609 & ~n27066;
  assign n27075 = pi1155 & ~n27074;
  assign n27076 = ~n27073 & n27075;
  assign n27077 = ~pi609 & ~n60007;
  assign n27078 = pi609 & ~n27066;
  assign n27079 = ~pi1155 & ~n27078;
  assign n27080 = ~n27077 & n27079;
  assign n27081 = ~n27076 & ~n27080;
  assign n27082 = pi785 & ~n27081;
  assign n27083 = ~n27072 & ~n27082;
  assign n27084 = ~pi781 & ~n27083;
  assign n27085 = pi618 & n27083;
  assign n27086 = ~pi618 & ~n27066;
  assign n27087 = pi1154 & ~n27086;
  assign n27088 = ~n27085 & n27087;
  assign n27089 = ~pi618 & n27083;
  assign n27090 = pi618 & ~n27066;
  assign n27091 = ~pi1154 & ~n27090;
  assign n27092 = ~n27089 & n27091;
  assign n27093 = ~n27088 & ~n27092;
  assign n27094 = pi781 & ~n27093;
  assign n27095 = ~n27084 & ~n27094;
  assign n27096 = ~pi789 & ~n27095;
  assign n27097 = pi619 & n27095;
  assign n27098 = ~pi619 & ~n27066;
  assign n27099 = pi1159 & ~n27098;
  assign n27100 = ~n27097 & n27099;
  assign n27101 = ~pi619 & n27095;
  assign n27102 = pi619 & ~n27066;
  assign n27103 = ~pi1159 & ~n27102;
  assign n27104 = ~n27101 & n27103;
  assign n27105 = ~n27100 & ~n27104;
  assign n27106 = pi789 & ~n27105;
  assign n27107 = ~n27096 & ~n27106;
  assign n27108 = ~n8054 & ~n27107;
  assign n27109 = n8054 & n27066;
  assign n27110 = n8054 & ~n27066;
  assign n27111 = ~n8054 & n27107;
  assign n27112 = ~n27110 & ~n27111;
  assign n27113 = ~n27108 & ~n27109;
  assign n27114 = ~n7793 & ~n60008;
  assign n27115 = n7793 & ~n27066;
  assign n27116 = ~n7872 & ~n27115;
  assign n27117 = ~n7793 & n60008;
  assign n27118 = n7793 & n27066;
  assign n27119 = ~n27117 & ~n27118;
  assign n27120 = ~n7872 & ~n27119;
  assign n27121 = ~n27114 & n27116;
  assign n27122 = ~n9651 & ~n27066;
  assign n27123 = n59231 & ~n27066;
  assign n27124 = pi681 & n7490;
  assign n27125 = ~n2790 & n27124;
  assign n27126 = pi680 & pi681;
  assign n27127 = ~n7495 & n27126;
  assign n27128 = n2790 & n27127;
  assign n27129 = ~n27125 & ~n27128;
  assign n27130 = ~n6544 & ~n27129;
  assign n27131 = pi681 & n59222;
  assign n27132 = n7035 & n27126;
  assign n27133 = n6544 & n60010;
  assign n27134 = ~pi223 & ~n27133;
  assign n27135 = n6544 & ~n60010;
  assign n27136 = ~n6544 & ~n27125;
  assign n27137 = ~n6544 & ~n27128;
  assign n27138 = ~n27125 & n27137;
  assign n27139 = ~n27128 & n27136;
  assign n27140 = ~n27135 & ~n60011;
  assign n27141 = ~pi223 & ~n27140;
  assign n27142 = ~n27130 & n27134;
  assign n27143 = pi681 & ~n7445;
  assign n27144 = ~n6511 & ~n27143;
  assign n27145 = ~n2790 & ~n27144;
  assign n27146 = pi681 & ~n7440;
  assign n27147 = ~n6535 & ~n27146;
  assign n27148 = n2790 & ~n27147;
  assign n27149 = pi223 & ~n27148;
  assign n27150 = ~n27145 & n27149;
  assign n27151 = ~pi299 & ~n27150;
  assign n27152 = ~n60012 & n27151;
  assign n27153 = n26980 & ~n60010;
  assign n27154 = pi681 & ~n7418;
  assign n27155 = n58846 & ~n6614;
  assign n27156 = ~n27154 & n27155;
  assign n27157 = pi681 & ~n26394;
  assign n27158 = ~n58846 & ~n6580;
  assign n27159 = ~n27157 & n27158;
  assign n27160 = pi223 & ~n27159;
  assign n27161 = ~n27156 & n27160;
  assign n27162 = n58846 & ~n27127;
  assign n27163 = ~n58846 & ~n27124;
  assign n27164 = ~pi223 & ~n27163;
  assign n27165 = ~pi223 & ~n27162;
  assign n27166 = ~n27163 & n27165;
  assign n27167 = ~n27162 & n27164;
  assign n27168 = ~n6629 & ~n60013;
  assign n27169 = ~n27161 & n27168;
  assign n27170 = ~n27153 & ~n27169;
  assign n27171 = ~pi215 & ~n27170;
  assign n27172 = ~n58846 & n27144;
  assign n27173 = n58846 & n27147;
  assign n27174 = pi223 & ~n27173;
  assign n27175 = ~n27172 & n27174;
  assign n27176 = ~pi223 & pi681;
  assign n27177 = n7531 & n27176;
  assign n27178 = pi215 & ~n27177;
  assign n27179 = ~n27175 & n27178;
  assign n27180 = pi299 & ~n27179;
  assign n27181 = ~n27171 & n27180;
  assign n27182 = ~n27152 & ~n27181;
  assign n27183 = pi39 & ~n27182;
  assign n27184 = ~pi223 & ~n7318;
  assign n27185 = n7318 & ~n27126;
  assign n27186 = pi223 & n7298;
  assign n27187 = ~pi299 & ~n27186;
  assign n27188 = ~n27185 & n27187;
  assign n27189 = ~n27184 & n27187;
  assign n27190 = ~n27185 & n27189;
  assign n27191 = ~n27184 & n27188;
  assign n27192 = n7327 & ~n27126;
  assign n27193 = ~pi223 & ~n7327;
  assign n27194 = pi223 & n7304;
  assign n27195 = pi299 & ~n27194;
  assign n27196 = ~n27193 & n27195;
  assign n27197 = ~n27192 & n27195;
  assign n27198 = ~n27193 & n27197;
  assign n27199 = ~n27192 & n27196;
  assign n27200 = ~n60014 & ~n60015;
  assign n27201 = ~pi39 & ~n27200;
  assign n27202 = ~pi38 & ~n27201;
  assign n27203 = ~pi39 & ~n60015;
  assign n27204 = ~pi39 & ~n60014;
  assign n27205 = ~n60015 & n27204;
  assign n27206 = ~n60014 & n27203;
  assign n27207 = pi39 & ~n27152;
  assign n27208 = ~n27181 & n27207;
  assign n27209 = ~n60016 & ~n27208;
  assign n27210 = ~pi38 & ~n27209;
  assign n27211 = ~n27183 & n27202;
  assign n27212 = pi223 & ~n6863;
  assign n27213 = pi681 & n7546;
  assign n27214 = pi38 & ~n27213;
  assign n27215 = ~n27212 & n27214;
  assign n27216 = n59132 & ~n27215;
  assign n27217 = ~n60017 & n27216;
  assign n27218 = ~n26909 & ~n27217;
  assign n27219 = ~pi778 & ~n27218;
  assign n27220 = pi625 & n27218;
  assign n27221 = ~pi625 & ~n27066;
  assign n27222 = pi1153 & ~n27221;
  assign n27223 = ~n27220 & n27222;
  assign n27224 = ~pi625 & n27218;
  assign n27225 = pi625 & ~n27066;
  assign n27226 = ~pi1153 & ~n27225;
  assign n27227 = ~n27224 & n27226;
  assign n27228 = ~n27223 & ~n27227;
  assign n27229 = pi778 & ~n27228;
  assign n27230 = ~n27219 & ~n27229;
  assign n27231 = ~n59229 & ~n27230;
  assign n27232 = n59229 & n27066;
  assign n27233 = n59229 & ~n27066;
  assign n27234 = ~n59229 & n27230;
  assign n27235 = ~n27233 & ~n27234;
  assign n27236 = ~n27231 & ~n27232;
  assign n27237 = ~n59231 & ~n60018;
  assign n27238 = ~n59231 & n60018;
  assign n27239 = n59231 & n27066;
  assign n27240 = ~n27238 & ~n27239;
  assign n27241 = ~n27123 & ~n27237;
  assign n27242 = ~n7716 & n60019;
  assign n27243 = ~n7762 & n27242;
  assign n27244 = ~n27122 & ~n27243;
  assign n27245 = ~n59240 & n27244;
  assign n27246 = n59240 & n27066;
  assign n27247 = ~n59240 & ~n27244;
  assign n27248 = n59240 & ~n27066;
  assign n27249 = ~n27247 & ~n27248;
  assign n27250 = ~n27245 & ~n27246;
  assign n27251 = pi647 & ~n60020;
  assign n27252 = ~pi647 & ~n27066;
  assign n27253 = pi1157 & ~n27252;
  assign n27254 = ~n27251 & n27253;
  assign n27255 = ~pi630 & n27254;
  assign n27256 = ~pi647 & ~n60020;
  assign n27257 = pi647 & ~n27066;
  assign n27258 = ~pi1157 & ~n27257;
  assign n27259 = ~n27256 & n27258;
  assign n27260 = pi630 & n27259;
  assign n27261 = ~n27255 & ~n27260;
  assign n27262 = ~n60009 & n27261;
  assign n27263 = pi787 & ~n27262;
  assign n27264 = ~n11154 & n60008;
  assign n27265 = ~pi628 & ~n27244;
  assign n27266 = pi628 & ~n27066;
  assign n27267 = n7791 & ~n27266;
  assign n27268 = ~n27265 & n27267;
  assign n27269 = pi628 & ~n27244;
  assign n27270 = ~pi628 & ~n27066;
  assign n27271 = n7790 & ~n27270;
  assign n27272 = ~n27269 & n27271;
  assign n27273 = ~n27268 & ~n27272;
  assign n27274 = ~n27264 & n27273;
  assign n27275 = pi792 & ~n27274;
  assign n27276 = pi626 & ~n27107;
  assign n27277 = ~pi626 & n27066;
  assign n27278 = n7759 & ~n27277;
  assign n27279 = ~n27276 & n27278;
  assign n27280 = n7716 & ~n27066;
  assign n27281 = ~n27242 & ~n27280;
  assign n27282 = n7984 & ~n27281;
  assign n27283 = ~pi626 & ~n27107;
  assign n27284 = pi626 & n27066;
  assign n27285 = n7760 & ~n27284;
  assign n27286 = ~n27283 & n27285;
  assign n27287 = ~n27282 & ~n27286;
  assign n27288 = ~n27279 & ~n27282;
  assign n27289 = ~n27286 & n27288;
  assign n27290 = ~n27279 & n27287;
  assign n27291 = pi788 & ~n60021;
  assign n27292 = n7331 & n27176;
  assign n27293 = n7330 & ~n27126;
  assign n27294 = ~n26702 & n26920;
  assign n27295 = ~n27293 & n27294;
  assign n27296 = n26918 & ~n27295;
  assign n27297 = n26918 & ~n27292;
  assign n27298 = ~n27295 & n27297;
  assign n27299 = ~n27292 & n27296;
  assign n27300 = n7322 & ~n27126;
  assign n27301 = ~n26688 & n26914;
  assign n27302 = ~n27300 & n27301;
  assign n27303 = n7323 & n27176;
  assign n27304 = n26912 & ~n27303;
  assign n27305 = ~n27302 & n27304;
  assign n27306 = ~pi39 & ~n27305;
  assign n27307 = ~pi39 & ~n60022;
  assign n27308 = ~n27305 & n27307;
  assign n27309 = ~n60022 & n27306;
  assign n27310 = ~pi680 & ~n26964;
  assign n27311 = pi642 & ~n7192;
  assign n27312 = ~n6873 & ~n27311;
  assign n27313 = n26927 & ~n27312;
  assign n27314 = pi680 & ~n27313;
  assign n27315 = pi642 & ~n7132;
  assign n27316 = n2777 & ~n27315;
  assign n27317 = ~pi642 & ~n7043;
  assign n27318 = n27316 & ~n27317;
  assign n27319 = n27314 & ~n27318;
  assign n27320 = ~n27310 & ~n27319;
  assign n27321 = pi681 & ~n27320;
  assign n27322 = ~n26968 & ~n27321;
  assign n27323 = n58846 & ~n27322;
  assign n27324 = ~n26956 & ~n27126;
  assign n27325 = ~pi642 & ~n2777;
  assign n27326 = ~n7015 & n27325;
  assign n27327 = pi642 & n7118;
  assign n27328 = pi680 & ~n27327;
  assign n27329 = ~n7122 & n27328;
  assign n27330 = ~n27326 & n27329;
  assign n27331 = ~n27324 & ~n27330;
  assign n27332 = ~n26961 & ~n27331;
  assign n27333 = ~n58846 & ~n27332;
  assign n27334 = ~pi223 & ~n27333;
  assign n27335 = ~pi223 & ~n27323;
  assign n27336 = ~n27333 & n27335;
  assign n27337 = ~n27323 & n27334;
  assign n27338 = ~n26934 & ~n27126;
  assign n27339 = ~pi642 & ~n6873;
  assign n27340 = pi642 & n7131;
  assign n27341 = ~n27339 & ~n27340;
  assign n27342 = pi642 & ~n7131;
  assign n27343 = n13069 & ~n27342;
  assign n27344 = n6468 & ~n27341;
  assign n27345 = ~n6461 & n60025;
  assign n27346 = ~n2777 & ~n27345;
  assign n27347 = pi680 & ~n27346;
  assign n27348 = ~n6879 & ~n27311;
  assign n27349 = n2777 & ~n27348;
  assign n27350 = n27347 & ~n27349;
  assign n27351 = ~n27338 & ~n27350;
  assign n27352 = n26941 & ~n27351;
  assign n27353 = ~n26946 & ~n27126;
  assign n27354 = n6700 & ~n26544;
  assign n27355 = n26546 & n27325;
  assign n27356 = pi642 & ~n59990;
  assign n27357 = pi680 & ~n27356;
  assign n27358 = ~n27355 & n27357;
  assign n27359 = ~n27354 & n27357;
  assign n27360 = ~n27355 & n27359;
  assign n27361 = ~n27354 & n27358;
  assign n27362 = ~n27353 & ~n60026;
  assign n27363 = n26951 & ~n27362;
  assign n27364 = pi223 & ~n27363;
  assign n27365 = ~n27352 & n27364;
  assign n27366 = ~n6629 & ~n27365;
  assign n27367 = ~n27352 & ~n27363;
  assign n27368 = pi223 & ~n27367;
  assign n27369 = n58846 & n27322;
  assign n27370 = ~n58846 & n27332;
  assign n27371 = ~pi223 & ~n27370;
  assign n27372 = ~n27369 & n27371;
  assign n27373 = ~n27368 & ~n27372;
  assign n27374 = ~n6629 & ~n27373;
  assign n27375 = ~n60024 & n27366;
  assign n27376 = n26928 & ~n27126;
  assign n27377 = n27126 & ~n27339;
  assign n27378 = ~n26719 & n27377;
  assign n27379 = ~n27376 & ~n27378;
  assign n27380 = n6464 & ~n27379;
  assign n27381 = ~pi223 & n27380;
  assign n27382 = n27126 & n60025;
  assign n27383 = n27007 & ~n27126;
  assign n27384 = pi223 & ~n27383;
  assign n27385 = ~n27382 & n27384;
  assign n27386 = n26980 & ~n27385;
  assign n27387 = ~n27381 & n27386;
  assign n27388 = ~pi215 & ~n27387;
  assign n27389 = ~n60027 & n27388;
  assign n27390 = ~n27005 & ~n27126;
  assign n27391 = ~pi614 & n6929;
  assign n27392 = ~n27311 & ~n27391;
  assign n27393 = ~pi616 & ~n27392;
  assign n27394 = n27347 & ~n27393;
  assign n27395 = ~n27390 & ~n27394;
  assign n27396 = ~n27011 & ~n27395;
  assign n27397 = n58846 & ~n27396;
  assign n27398 = ~n2777 & n6944;
  assign n27399 = pi642 & ~n26604;
  assign n27400 = pi680 & ~n6946;
  assign n27401 = ~n27399 & n27400;
  assign n27402 = ~n27398 & n27401;
  assign n27403 = ~pi680 & n60005;
  assign n27404 = pi681 & ~n27403;
  assign n27405 = pi681 & ~n27402;
  assign n27406 = ~n27403 & n27405;
  assign n27407 = ~n27402 & n27404;
  assign n27408 = ~n27021 & ~n60028;
  assign n27409 = ~n58846 & ~n27408;
  assign n27410 = pi223 & ~n27409;
  assign n27411 = ~n27397 & n27410;
  assign n27412 = ~n26993 & ~n27126;
  assign n27413 = n7062 & n7169;
  assign n27414 = n6700 & ~n27413;
  assign n27415 = ~n7061 & n27325;
  assign n27416 = pi642 & n26618;
  assign n27417 = pi680 & ~n27416;
  assign n27418 = pi680 & ~n27415;
  assign n27419 = ~n27416 & n27418;
  assign n27420 = ~n27415 & n27417;
  assign n27421 = ~n27414 & n60029;
  assign n27422 = ~n27412 & ~n27421;
  assign n27423 = ~n58846 & n26991;
  assign n27424 = ~n27422 & n27423;
  assign n27425 = ~n7063 & n27316;
  assign n27426 = n27314 & ~n27425;
  assign n27427 = ~n27310 & ~n27426;
  assign n27428 = pi681 & ~n27427;
  assign n27429 = n26996 & ~n27428;
  assign n27430 = ~pi223 & ~n27429;
  assign n27431 = ~n27424 & n27430;
  assign n27432 = pi215 & ~n27431;
  assign n27433 = ~n27411 & n27432;
  assign n27434 = pi299 & ~n27433;
  assign n27435 = ~n27389 & n27434;
  assign n27436 = ~n2790 & n27332;
  assign n27437 = n2790 & n27322;
  assign n27438 = ~n6544 & ~n27437;
  assign n27439 = ~n6544 & ~n27436;
  assign n27440 = ~n27437 & n27439;
  assign n27441 = ~n27436 & n27438;
  assign n27442 = n6544 & ~n27380;
  assign n27443 = ~pi223 & ~n27442;
  assign n27444 = ~n60030 & n27443;
  assign n27445 = n2790 & n27396;
  assign n27446 = ~n2790 & n27408;
  assign n27447 = pi223 & ~n27446;
  assign n27448 = ~n27445 & n27447;
  assign n27449 = ~pi299 & ~n27448;
  assign n27450 = n2790 & ~n27396;
  assign n27451 = ~n2790 & ~n27408;
  assign n27452 = pi223 & ~n27451;
  assign n27453 = ~n27450 & n27452;
  assign n27454 = ~n27436 & ~n27437;
  assign n27455 = ~n6544 & ~n27454;
  assign n27456 = n6544 & n27380;
  assign n27457 = ~pi223 & ~n27456;
  assign n27458 = ~n27455 & n27457;
  assign n27459 = ~n27453 & ~n27458;
  assign n27460 = ~pi299 & ~n27459;
  assign n27461 = ~n27444 & n27449;
  assign n27462 = pi39 & ~n60031;
  assign n27463 = ~n27435 & n27462;
  assign n27464 = ~pi38 & ~n27463;
  assign n27465 = ~pi38 & ~n60023;
  assign n27466 = ~n27463 & n27465;
  assign n27467 = ~n60023 & n27464;
  assign n27468 = n27379 & ~n27385;
  assign n27469 = n27053 & ~n27468;
  assign n27470 = n27051 & ~n27469;
  assign n27471 = n59132 & ~n27470;
  assign n27472 = ~n60032 & n27471;
  assign n27473 = ~n26909 & ~n27472;
  assign n27474 = ~pi625 & n27473;
  assign n27475 = pi625 & n27058;
  assign n27476 = ~pi1153 & ~n27475;
  assign n27477 = ~n27474 & n27476;
  assign n27478 = ~pi608 & ~n27477;
  assign n27479 = ~n27223 & n27478;
  assign n27480 = pi625 & n27473;
  assign n27481 = ~pi625 & n27058;
  assign n27482 = pi1153 & ~n27481;
  assign n27483 = ~n27480 & n27482;
  assign n27484 = pi608 & ~n27483;
  assign n27485 = ~n27227 & n27484;
  assign n27486 = ~n27479 & ~n27485;
  assign n27487 = pi778 & ~n27486;
  assign n27488 = ~pi778 & n27473;
  assign n27489 = ~n27487 & ~n27488;
  assign n27490 = ~pi609 & ~n27489;
  assign n27491 = pi609 & n27230;
  assign n27492 = ~pi1155 & ~n27491;
  assign n27493 = ~n27490 & n27492;
  assign n27494 = ~pi660 & ~n27076;
  assign n27495 = ~n27493 & n27494;
  assign n27496 = pi609 & ~n27489;
  assign n27497 = ~pi609 & n27230;
  assign n27498 = pi1155 & ~n27497;
  assign n27499 = ~n27496 & n27498;
  assign n27500 = pi660 & ~n27080;
  assign n27501 = ~n27499 & n27500;
  assign n27502 = ~n27495 & ~n27501;
  assign n27503 = pi785 & ~n27502;
  assign n27504 = ~pi785 & ~n27489;
  assign n27505 = ~n27503 & ~n27504;
  assign n27506 = ~pi618 & ~n27505;
  assign n27507 = pi618 & ~n60018;
  assign n27508 = ~pi1154 & ~n27507;
  assign n27509 = ~n27506 & n27508;
  assign n27510 = ~pi627 & ~n27088;
  assign n27511 = ~n27509 & n27510;
  assign n27512 = pi618 & ~n27505;
  assign n27513 = ~pi618 & ~n60018;
  assign n27514 = pi1154 & ~n27513;
  assign n27515 = ~n27512 & n27514;
  assign n27516 = pi627 & ~n27092;
  assign n27517 = ~n27515 & n27516;
  assign n27518 = ~n27511 & ~n27517;
  assign n27519 = pi781 & ~n27518;
  assign n27520 = ~pi781 & ~n27505;
  assign n27521 = ~n27519 & ~n27520;
  assign n27522 = pi619 & ~n27521;
  assign n27523 = ~pi619 & n60019;
  assign n27524 = pi1159 & ~n27523;
  assign n27525 = ~n27522 & n27524;
  assign n27526 = pi648 & ~n27104;
  assign n27527 = ~n27525 & n27526;
  assign n27528 = ~pi619 & ~n27521;
  assign n27529 = pi619 & n60019;
  assign n27530 = ~pi1159 & ~n27529;
  assign n27531 = ~n27528 & n27530;
  assign n27532 = ~pi648 & ~n27100;
  assign n27533 = ~n27531 & n27532;
  assign n27534 = pi789 & ~n27533;
  assign n27535 = pi789 & ~n27527;
  assign n27536 = ~n27533 & n27535;
  assign n27537 = ~n27527 & n27534;
  assign n27538 = ~pi789 & n27521;
  assign n27539 = n59242 & ~n27538;
  assign n27540 = ~n60033 & n27539;
  assign n27541 = ~n27291 & ~n27540;
  assign n27542 = ~n27275 & ~n27541;
  assign n27543 = n59357 & n27274;
  assign n27544 = ~n8108 & ~n27543;
  assign n27545 = ~n27542 & n27544;
  assign n27546 = ~n27263 & ~n27545;
  assign n27547 = ~n23536 & n27546;
  assign n27548 = ~n27254 & ~n27259;
  assign n27549 = pi787 & ~n27548;
  assign n27550 = ~pi787 & n60020;
  assign n27551 = ~n23547 & ~n27550;
  assign n27552 = ~n27549 & n27551;
  assign n27553 = n26860 & ~n27066;
  assign n27554 = pi790 & ~n27553;
  assign n27555 = ~n27552 & n27554;
  assign n27556 = n12602 & n27107;
  assign n27557 = n23557 & n27556;
  assign n27558 = n23562 & ~n27066;
  assign n27559 = ~n27557 & ~n27558;
  assign n27560 = pi644 & ~n27559;
  assign n27561 = n23562 & n27556;
  assign n27562 = n23557 & ~n27066;
  assign n27563 = ~n27561 & ~n27562;
  assign n27564 = ~pi644 & ~n27563;
  assign n27565 = ~n27560 & ~n27564;
  assign n27566 = n27555 & n27565;
  assign n27567 = ~n27547 & n27566;
  assign n27568 = ~pi790 & ~n27546;
  assign n27569 = ~pi644 & n27546;
  assign n27570 = ~n27549 & ~n27550;
  assign n27571 = pi644 & n27570;
  assign n27572 = ~pi715 & ~n27571;
  assign n27573 = ~n27569 & n27572;
  assign n27574 = n7835 & ~n27066;
  assign n27575 = ~n7835 & n27119;
  assign n27576 = ~n27574 & ~n27575;
  assign n27577 = ~pi644 & ~n27576;
  assign n27578 = pi644 & ~n27066;
  assign n27579 = pi715 & ~n27578;
  assign n27580 = ~n27577 & n27579;
  assign n27581 = ~pi1160 & ~n27580;
  assign n27582 = ~n27573 & n27581;
  assign n27583 = pi644 & n27546;
  assign n27584 = ~pi644 & n27570;
  assign n27585 = pi715 & ~n27584;
  assign n27586 = ~n27583 & n27585;
  assign n27587 = pi644 & ~n27576;
  assign n27588 = ~pi644 & ~n27066;
  assign n27589 = ~pi715 & ~n27588;
  assign n27590 = ~n27587 & n27589;
  assign n27591 = pi1160 & ~n27590;
  assign n27592 = ~n27586 & n27591;
  assign n27593 = ~n27582 & ~n27592;
  assign n27594 = pi790 & ~n27593;
  assign n27595 = ~pi790 & n27546;
  assign n27596 = ~n27594 & ~n27595;
  assign n27597 = ~n27567 & ~n27568;
  assign n27598 = n58992 & n60034;
  assign n27599 = pi223 & ~n58992;
  assign n27600 = n58992 & ~n60034;
  assign n27601 = ~pi223 & ~n58992;
  assign n27602 = ~n27600 & ~n27601;
  assign n27603 = ~n27598 & ~n27599;
  assign n27604 = pi224 & ~n26176;
  assign n27605 = n7597 & ~n27604;
  assign n27606 = pi224 & ~n59132;
  assign n27607 = pi614 & n6701;
  assign n27608 = n6464 & ~n27607;
  assign n27609 = ~n2778 & ~n27608;
  assign n27610 = ~n6594 & ~n27609;
  assign n27611 = ~n6518 & ~n27610;
  assign n27612 = ~pi680 & ~n27610;
  assign n27613 = pi680 & n27607;
  assign n27614 = ~n6606 & ~n27613;
  assign n27615 = ~n27612 & n27614;
  assign n27616 = n6518 & ~n27615;
  assign n27617 = ~n27611 & ~n27616;
  assign n27618 = n58846 & n27617;
  assign n27619 = ~n2680 & n6591;
  assign n27620 = n2777 & ~n6567;
  assign n27621 = ~n27619 & n27620;
  assign n27622 = pi614 & ~n7014;
  assign n27623 = ~pi614 & pi616;
  assign n27624 = n6568 & n27623;
  assign n27625 = ~n27622 & ~n27624;
  assign n27626 = ~n2680 & n6600;
  assign n27627 = ~pi614 & ~n6567;
  assign n27628 = ~n27626 & n27627;
  assign n27629 = ~n27622 & ~n27628;
  assign n27630 = ~n27621 & n27625;
  assign n27631 = ~n6518 & ~n60036;
  assign n27632 = ~pi680 & ~n60036;
  assign n27633 = pi614 & n6904;
  assign n27634 = pi680 & ~n27633;
  assign n27635 = n6566 & n27634;
  assign n27636 = ~n27613 & ~n27635;
  assign n27637 = ~n27632 & n27636;
  assign n27638 = n6518 & ~n27637;
  assign n27639 = ~n27631 & ~n27638;
  assign n27640 = ~n58846 & n27639;
  assign n27641 = pi224 & ~n27640;
  assign n27642 = pi224 & ~n27618;
  assign n27643 = ~n27640 & n27642;
  assign n27644 = ~n27618 & n27641;
  assign n27645 = ~n6568 & n27607;
  assign n27646 = ~pi680 & ~n27645;
  assign n27647 = ~n27634 & ~n27646;
  assign n27648 = n6518 & ~n27647;
  assign n27649 = ~n6518 & ~n27645;
  assign n27650 = ~n27648 & ~n27649;
  assign n27651 = ~n58846 & ~n27650;
  assign n27652 = pi614 & ~n59969;
  assign n27653 = n58846 & ~n27652;
  assign n27654 = ~pi224 & ~n27653;
  assign n27655 = ~n27651 & n27654;
  assign n27656 = ~n6629 & ~n27655;
  assign n27657 = ~n60037 & n27656;
  assign n27658 = n6610 & n6701;
  assign n27659 = pi224 & ~n6464;
  assign n27660 = n6629 & ~n27659;
  assign n27661 = ~n27658 & n27660;
  assign n27662 = ~pi215 & ~n27661;
  assign n27663 = ~n27657 & n27662;
  assign n27664 = pi614 & ~n26240;
  assign n27665 = ~n59971 & n27658;
  assign n27666 = ~pi224 & n60038;
  assign n27667 = ~n6833 & n27666;
  assign n27668 = ~n6501 & ~n27609;
  assign n27669 = ~n6518 & ~n27668;
  assign n27670 = ~pi680 & ~n27668;
  assign n27671 = ~n6522 & ~n27613;
  assign n27672 = ~n27670 & n27671;
  assign n27673 = n6518 & ~n27672;
  assign n27674 = ~n27669 & ~n27673;
  assign n27675 = n58846 & n27674;
  assign n27676 = ~n7067 & ~n25459;
  assign n27677 = ~n25458 & n27676;
  assign n27678 = pi614 & ~n6732;
  assign n27679 = ~n27677 & ~n27678;
  assign n27680 = ~pi680 & ~n27679;
  assign n27681 = ~pi614 & ~n6484;
  assign n27682 = n6737 & ~n27681;
  assign n27683 = ~n27680 & ~n27682;
  assign n27684 = n6518 & ~n27683;
  assign n27685 = ~n6518 & ~n27679;
  assign n27686 = ~n27684 & ~n27685;
  assign n27687 = ~n58846 & n27686;
  assign n27688 = pi224 & ~n27687;
  assign n27689 = ~n27675 & n27688;
  assign n27690 = ~n27667 & ~n27689;
  assign n27691 = pi215 & ~n27690;
  assign n27692 = pi299 & ~n27691;
  assign n27693 = ~n27663 & n27692;
  assign n27694 = n2790 & n27674;
  assign n27695 = ~n2790 & n27686;
  assign n27696 = pi224 & ~n27695;
  assign n27697 = ~n27694 & n27696;
  assign n27698 = ~n6848 & n27666;
  assign n27699 = pi223 & ~n27698;
  assign n27700 = ~n27697 & n27699;
  assign n27701 = n2790 & n27617;
  assign n27702 = ~n2790 & n27639;
  assign n27703 = pi224 & ~n27702;
  assign n27704 = pi224 & ~n27701;
  assign n27705 = ~n27702 & n27704;
  assign n27706 = ~n27701 & n27703;
  assign n27707 = ~n2790 & ~n27650;
  assign n27708 = n2790 & ~n27652;
  assign n27709 = n2827 & ~n27708;
  assign n27710 = ~n27707 & n27709;
  assign n27711 = pi614 & n59169;
  assign n27712 = n59155 & n27607;
  assign n27713 = ~pi223 & ~n60040;
  assign n27714 = ~n27710 & n27713;
  assign n27715 = ~n60039 & n27714;
  assign n27716 = ~n27700 & ~n27715;
  assign n27717 = ~pi299 & ~n27716;
  assign n27718 = pi39 & ~n27717;
  assign n27719 = pi39 & ~n27693;
  assign n27720 = ~n27717 & n27719;
  assign n27721 = ~n27693 & n27718;
  assign n27722 = ~pi614 & n6791;
  assign n27723 = pi224 & ~n27722;
  assign n27724 = n6671 & n27723;
  assign n27725 = pi614 & n6791;
  assign n27726 = ~pi224 & n27725;
  assign n27727 = ~pi299 & ~n27726;
  assign n27728 = ~n27724 & n27727;
  assign n27729 = pi614 & n6796;
  assign n27730 = pi224 & ~n6453;
  assign n27731 = ~n27729 & ~n27730;
  assign n27732 = pi299 & n27731;
  assign n27733 = ~pi39 & ~n27732;
  assign n27734 = ~pi39 & ~n27728;
  assign n27735 = ~n27732 & n27734;
  assign n27736 = ~n27728 & n27733;
  assign n27737 = ~pi38 & ~n60042;
  assign n27738 = ~n60041 & n27737;
  assign n27739 = pi224 & ~n6863;
  assign n27740 = pi38 & ~n27739;
  assign n27741 = n6863 & n27607;
  assign n27742 = pi614 & n6865;
  assign n27743 = n27740 & ~n60043;
  assign n27744 = n59132 & ~n27743;
  assign n27745 = ~n27738 & n27744;
  assign n27746 = ~n27606 & ~n27745;
  assign n27747 = ~n7597 & n27746;
  assign n27748 = ~n7597 & ~n27746;
  assign n27749 = n7597 & n27604;
  assign n27750 = ~n27748 & ~n27749;
  assign n27751 = ~n27605 & ~n27747;
  assign n27752 = ~pi785 & ~n60044;
  assign n27753 = pi609 & n60044;
  assign n27754 = ~pi609 & ~n27604;
  assign n27755 = pi1155 & ~n27754;
  assign n27756 = ~n27753 & n27755;
  assign n27757 = ~pi609 & n60044;
  assign n27758 = pi609 & ~n27604;
  assign n27759 = ~pi1155 & ~n27758;
  assign n27760 = ~n27757 & n27759;
  assign n27761 = ~n27756 & ~n27760;
  assign n27762 = pi785 & ~n27761;
  assign n27763 = ~n27752 & ~n27762;
  assign n27764 = ~pi781 & ~n27763;
  assign n27765 = pi618 & n27763;
  assign n27766 = ~pi618 & ~n27604;
  assign n27767 = pi1154 & ~n27766;
  assign n27768 = ~n27765 & n27767;
  assign n27769 = ~pi618 & n27763;
  assign n27770 = pi618 & ~n27604;
  assign n27771 = ~pi1154 & ~n27770;
  assign n27772 = ~n27769 & n27771;
  assign n27773 = ~n27768 & ~n27772;
  assign n27774 = pi781 & ~n27773;
  assign n27775 = ~n27764 & ~n27774;
  assign n27776 = ~pi789 & ~n27775;
  assign n27777 = pi619 & n27775;
  assign n27778 = ~pi619 & ~n27604;
  assign n27779 = pi1159 & ~n27778;
  assign n27780 = ~n27777 & n27779;
  assign n27781 = ~pi619 & n27775;
  assign n27782 = pi619 & ~n27604;
  assign n27783 = ~pi1159 & ~n27782;
  assign n27784 = ~n27781 & n27783;
  assign n27785 = ~n27780 & ~n27784;
  assign n27786 = pi789 & ~n27785;
  assign n27787 = ~n27776 & ~n27786;
  assign n27788 = ~n8054 & n27787;
  assign n27789 = n8054 & ~n27604;
  assign n27790 = ~n27788 & ~n27789;
  assign n27791 = ~n7793 & ~n27790;
  assign n27792 = n7793 & ~n27604;
  assign n27793 = ~n7872 & ~n27792;
  assign n27794 = ~n7793 & n27790;
  assign n27795 = n7793 & n27604;
  assign n27796 = ~n27794 & ~n27795;
  assign n27797 = ~n7872 & ~n27796;
  assign n27798 = ~n27791 & n27793;
  assign n27799 = ~n9651 & ~n27604;
  assign n27800 = n59229 & ~n27604;
  assign n27801 = ~pi224 & ~n7327;
  assign n27802 = pi662 & pi680;
  assign n27803 = n7327 & ~n27802;
  assign n27804 = pi224 & n7304;
  assign n27805 = pi299 & ~n27804;
  assign n27806 = ~n27803 & n27805;
  assign n27807 = ~n27801 & n27805;
  assign n27808 = ~n27803 & n27807;
  assign n27809 = ~n27801 & n27806;
  assign n27810 = ~pi224 & ~n7318;
  assign n27811 = n7318 & ~n27802;
  assign n27812 = pi224 & n7298;
  assign n27813 = ~pi299 & ~n27812;
  assign n27814 = ~n27811 & n27813;
  assign n27815 = ~n27810 & n27813;
  assign n27816 = ~n27811 & n27815;
  assign n27817 = ~n27810 & n27814;
  assign n27818 = ~pi39 & ~n60047;
  assign n27819 = ~pi39 & ~n60046;
  assign n27820 = ~n60047 & n27819;
  assign n27821 = ~n60046 & n27818;
  assign n27822 = pi662 & n59222;
  assign n27823 = n7035 & n27802;
  assign n27824 = n27660 & ~n60049;
  assign n27825 = pi662 & ~n7418;
  assign n27826 = ~pi662 & ~n6615;
  assign n27827 = ~n27825 & ~n27826;
  assign n27828 = n58846 & n27827;
  assign n27829 = ~n2779 & ~n26394;
  assign n27830 = n59152 & ~n27829;
  assign n27831 = ~n58846 & n27830;
  assign n27832 = pi224 & ~n27831;
  assign n27833 = ~n27828 & n27832;
  assign n27834 = pi662 & n7490;
  assign n27835 = ~n58846 & ~n27834;
  assign n27836 = ~n7495 & n27802;
  assign n27837 = n58846 & ~n27836;
  assign n27838 = ~pi224 & ~n27837;
  assign n27839 = ~pi224 & ~n27835;
  assign n27840 = ~n27837 & n27839;
  assign n27841 = ~n27835 & n27838;
  assign n27842 = ~n6629 & ~n60050;
  assign n27843 = ~n27833 & n27842;
  assign n27844 = ~n27824 & ~n27843;
  assign n27845 = ~pi215 & ~n27844;
  assign n27846 = ~pi662 & ~n6512;
  assign n27847 = pi662 & ~n7445;
  assign n27848 = ~n27846 & ~n27847;
  assign n27849 = ~n58846 & n27848;
  assign n27850 = ~pi662 & ~n59149;
  assign n27851 = pi662 & ~n7440;
  assign n27852 = ~n27850 & ~n27851;
  assign n27853 = n58846 & n27852;
  assign n27854 = pi224 & ~n27853;
  assign n27855 = ~n27849 & n27854;
  assign n27856 = ~pi224 & pi662;
  assign n27857 = n7531 & n27856;
  assign n27858 = pi215 & ~n27857;
  assign n27859 = ~n27855 & n27858;
  assign n27860 = pi299 & ~n27859;
  assign n27861 = ~n27845 & n27860;
  assign n27862 = n2790 & n27827;
  assign n27863 = ~n2790 & n27830;
  assign n27864 = pi224 & ~n27863;
  assign n27865 = ~n27862 & n27864;
  assign n27866 = ~n2790 & ~n27834;
  assign n27867 = n2790 & ~n27836;
  assign n27868 = n2827 & ~n27867;
  assign n27869 = n2827 & ~n27866;
  assign n27870 = ~n27867 & n27869;
  assign n27871 = ~n27866 & n27868;
  assign n27872 = pi662 & n7489;
  assign n27873 = ~pi223 & ~n27872;
  assign n27874 = ~n60051 & n27873;
  assign n27875 = ~n27865 & n27874;
  assign n27876 = ~n2790 & n27848;
  assign n27877 = n2790 & n27852;
  assign n27878 = pi224 & ~n27877;
  assign n27879 = ~n27876 & n27878;
  assign n27880 = n7508 & n27856;
  assign n27881 = pi223 & ~n27880;
  assign n27882 = ~n27879 & n27881;
  assign n27883 = ~pi299 & ~n27882;
  assign n27884 = ~n27875 & n27883;
  assign n27885 = pi39 & ~n27884;
  assign n27886 = ~n27861 & n27885;
  assign n27887 = ~n60048 & ~n27886;
  assign n27888 = ~pi38 & ~n27887;
  assign n27889 = pi662 & n7546;
  assign n27890 = n27740 & ~n27889;
  assign n27891 = n59132 & ~n27890;
  assign n27892 = ~n27888 & n27891;
  assign n27893 = ~n27606 & ~n27892;
  assign n27894 = ~pi778 & ~n27893;
  assign n27895 = pi625 & n27893;
  assign n27896 = ~pi625 & ~n27604;
  assign n27897 = pi1153 & ~n27896;
  assign n27898 = ~n27895 & n27897;
  assign n27899 = ~pi625 & n27893;
  assign n27900 = pi625 & ~n27604;
  assign n27901 = ~pi1153 & ~n27900;
  assign n27902 = ~n27899 & n27901;
  assign n27903 = ~n27898 & ~n27902;
  assign n27904 = pi778 & ~n27903;
  assign n27905 = ~n27894 & ~n27904;
  assign n27906 = ~n59229 & n27905;
  assign n27907 = ~n59229 & ~n27905;
  assign n27908 = n59229 & n27604;
  assign n27909 = ~n27907 & ~n27908;
  assign n27910 = ~n27800 & ~n27906;
  assign n27911 = ~n59231 & n60052;
  assign n27912 = n59231 & ~n27604;
  assign n27913 = ~n59231 & ~n60052;
  assign n27914 = n59231 & n27604;
  assign n27915 = ~n27913 & ~n27914;
  assign n27916 = ~n27911 & ~n27912;
  assign n27917 = ~n7716 & n60053;
  assign n27918 = ~n7762 & n27917;
  assign n27919 = ~n27799 & ~n27918;
  assign n27920 = ~n59240 & n27919;
  assign n27921 = n59240 & n27604;
  assign n27922 = ~n59240 & ~n27919;
  assign n27923 = n59240 & ~n27604;
  assign n27924 = ~n27922 & ~n27923;
  assign n27925 = ~n27920 & ~n27921;
  assign n27926 = pi647 & ~n60054;
  assign n27927 = ~pi647 & ~n27604;
  assign n27928 = pi1157 & ~n27927;
  assign n27929 = ~n27926 & n27928;
  assign n27930 = ~pi630 & n27929;
  assign n27931 = ~pi647 & ~n60054;
  assign n27932 = pi647 & ~n27604;
  assign n27933 = ~pi1157 & ~n27932;
  assign n27934 = ~n27931 & n27933;
  assign n27935 = pi630 & n27934;
  assign n27936 = ~n27930 & ~n27935;
  assign n27937 = ~n60045 & n27936;
  assign n27938 = pi787 & ~n27937;
  assign n27939 = ~n11154 & n27790;
  assign n27940 = ~pi628 & ~n27919;
  assign n27941 = pi628 & ~n27604;
  assign n27942 = n7791 & ~n27941;
  assign n27943 = ~n27940 & n27942;
  assign n27944 = pi628 & ~n27919;
  assign n27945 = ~pi628 & ~n27604;
  assign n27946 = n7790 & ~n27945;
  assign n27947 = ~n27944 & n27946;
  assign n27948 = ~n27943 & ~n27947;
  assign n27949 = ~n27939 & n27948;
  assign n27950 = pi792 & ~n27949;
  assign n27951 = ~pi614 & ~n13069;
  assign n27952 = pi614 & ~n26719;
  assign n27953 = ~n27951 & ~n27952;
  assign n27954 = ~n6461 & n27953;
  assign n27955 = pi616 & ~n27954;
  assign n27956 = pi614 & ~n7192;
  assign n27957 = ~n6881 & ~n27956;
  assign n27958 = ~pi616 & ~n27957;
  assign n27959 = ~n27955 & ~n27958;
  assign n27960 = pi680 & ~n27959;
  assign n27961 = ~n27612 & ~n27960;
  assign n27962 = pi662 & ~n27961;
  assign n27963 = ~pi662 & ~n6517;
  assign n27964 = ~n27610 & n27963;
  assign n27965 = ~n27616 & ~n27964;
  assign n27966 = ~n27962 & n27965;
  assign n27967 = pi224 & ~n27966;
  assign n27968 = ~n59182 & n27623;
  assign n27969 = ~n26516 & ~n27968;
  assign n27970 = pi680 & ~n27969;
  assign n27971 = ~n26517 & ~n27658;
  assign n27972 = ~n27970 & ~n27971;
  assign n27973 = pi662 & ~n27972;
  assign n27974 = ~pi662 & ~n27652;
  assign n27975 = ~n27973 & ~n27974;
  assign n27976 = ~pi224 & n27975;
  assign n27977 = n58846 & ~n27976;
  assign n27978 = ~n27967 & n27977;
  assign n27979 = pi614 & ~n59990;
  assign n27980 = n26546 & n27623;
  assign n27981 = ~n27979 & ~n27980;
  assign n27982 = ~n59989 & n27981;
  assign n27983 = pi680 & ~n27982;
  assign n27984 = ~n27632 & ~n27983;
  assign n27985 = pi662 & ~n27984;
  assign n27986 = ~n60036 & n27963;
  assign n27987 = ~n27638 & ~n27986;
  assign n27988 = ~n27985 & n27987;
  assign n27989 = pi224 & ~n27988;
  assign n27990 = ~pi614 & n7028;
  assign n27991 = pi614 & ~n7118;
  assign n27992 = pi680 & ~n27991;
  assign n27993 = ~n27990 & n27992;
  assign n27994 = ~n27646 & ~n27993;
  assign n27995 = pi662 & ~n27994;
  assign n27996 = ~n27645 & n27963;
  assign n27997 = ~n27648 & ~n27996;
  assign n27998 = ~n27995 & n27997;
  assign n27999 = ~pi224 & n27998;
  assign n28000 = ~n58846 & ~n27999;
  assign n28001 = ~n27989 & n28000;
  assign n28002 = ~n27978 & ~n28001;
  assign n28003 = ~pi224 & ~n27998;
  assign n28004 = pi224 & n27988;
  assign n28005 = ~n58846 & ~n28004;
  assign n28006 = ~n58846 & ~n28003;
  assign n28007 = ~n28004 & n28006;
  assign n28008 = ~n28003 & n28005;
  assign n28009 = pi224 & n27966;
  assign n28010 = ~pi224 & ~n27975;
  assign n28011 = n58846 & ~n28010;
  assign n28012 = ~n28009 & n28011;
  assign n28013 = ~n6629 & ~n28012;
  assign n28014 = ~n60055 & n28013;
  assign n28015 = ~n6629 & ~n60055;
  assign n28016 = ~n28012 & n28015;
  assign n28017 = ~n6629 & ~n28002;
  assign n28018 = n59182 & n27802;
  assign n28019 = ~n27658 & ~n28018;
  assign n28020 = ~pi224 & ~n28019;
  assign n28021 = n27802 & n27953;
  assign n28022 = ~n27607 & ~n27802;
  assign n28023 = n6468 & n28022;
  assign n28024 = pi224 & ~n28023;
  assign n28025 = ~n28021 & n28024;
  assign n28026 = n27660 & ~n28025;
  assign n28027 = ~n28020 & n28026;
  assign n28028 = ~pi215 & ~n28027;
  assign n28029 = ~n60056 & n28028;
  assign n28030 = pi680 & ~n7082;
  assign n28031 = ~n27658 & ~n28030;
  assign n28032 = ~n27970 & ~n28031;
  assign n28033 = pi662 & ~n28032;
  assign n28034 = ~pi662 & ~n60038;
  assign n28035 = ~n28033 & ~n28034;
  assign n28036 = ~pi224 & ~n28035;
  assign n28037 = ~n6931 & ~n27956;
  assign n28038 = ~pi616 & ~n28037;
  assign n28039 = ~n27955 & ~n28038;
  assign n28040 = pi680 & ~n28039;
  assign n28041 = ~n27670 & ~n28040;
  assign n28042 = pi662 & ~n28041;
  assign n28043 = ~n27668 & n27963;
  assign n28044 = pi224 & ~n28043;
  assign n28045 = ~n27673 & n28044;
  assign n28046 = ~n27673 & ~n28043;
  assign n28047 = ~n28042 & n28046;
  assign n28048 = pi224 & n28047;
  assign n28049 = ~n28042 & n28045;
  assign n28050 = ~n28036 & ~n60057;
  assign n28051 = n58846 & ~n28050;
  assign n28052 = pi614 & ~n26604;
  assign n28053 = n6947 & ~n28052;
  assign n28054 = pi680 & ~n28053;
  assign n28055 = ~n27680 & ~n28054;
  assign n28056 = pi662 & ~n28055;
  assign n28057 = ~n27679 & n27963;
  assign n28058 = pi224 & ~n28057;
  assign n28059 = ~n27684 & n28058;
  assign n28060 = ~n27684 & ~n28057;
  assign n28061 = ~n28056 & n28060;
  assign n28062 = pi224 & n28061;
  assign n28063 = ~n28056 & n28059;
  assign n28064 = ~pi614 & n7073;
  assign n28065 = pi614 & n26618;
  assign n28066 = pi680 & ~n28065;
  assign n28067 = ~n28064 & n28066;
  assign n28068 = ~n7070 & n28067;
  assign n28069 = pi614 & ~pi680;
  assign n28070 = n6828 & n28069;
  assign n28071 = pi662 & ~n28070;
  assign n28072 = ~pi616 & n7063;
  assign n28073 = n7061 & ~n28072;
  assign n28074 = ~pi614 & ~n28073;
  assign n28075 = ~n6486 & n27658;
  assign n28076 = ~pi680 & ~n28075;
  assign n28077 = ~n28065 & ~n28076;
  assign n28078 = ~n28074 & n28077;
  assign n28079 = pi662 & ~n28078;
  assign n28080 = ~n28068 & n28071;
  assign n28081 = ~pi662 & n6486;
  assign n28082 = ~n6486 & n60038;
  assign n28083 = ~pi662 & ~n28082;
  assign n28084 = ~n28034 & ~n28081;
  assign n28085 = ~n60059 & ~n60060;
  assign n28086 = ~pi224 & ~n28085;
  assign n28087 = ~n60058 & ~n28086;
  assign n28088 = ~n58846 & ~n28087;
  assign n28089 = pi215 & ~n28088;
  assign n28090 = n58846 & ~n28047;
  assign n28091 = ~n58846 & ~n28061;
  assign n28092 = pi224 & ~n28091;
  assign n28093 = ~n28090 & n28092;
  assign n28094 = n58846 & n28035;
  assign n28095 = ~n58846 & n28085;
  assign n28096 = ~pi224 & ~n28095;
  assign n28097 = ~n28094 & n28096;
  assign n28098 = pi215 & ~n28097;
  assign n28099 = ~n28093 & n28098;
  assign n28100 = ~n28051 & n28089;
  assign n28101 = pi299 & ~n60061;
  assign n28102 = ~n28029 & n28101;
  assign n28103 = n2790 & ~n28036;
  assign n28104 = n2790 & n28050;
  assign n28105 = ~n60057 & n28103;
  assign n28106 = ~n2790 & ~n28086;
  assign n28107 = ~n60058 & n28106;
  assign n28108 = ~n2790 & n28087;
  assign n28109 = pi223 & ~n60063;
  assign n28110 = ~n60062 & n28109;
  assign n28111 = n2790 & n27966;
  assign n28112 = ~n2790 & n27988;
  assign n28113 = pi224 & ~n28112;
  assign n28114 = pi224 & ~n28111;
  assign n28115 = ~n28112 & n28114;
  assign n28116 = ~n28111 & n28113;
  assign n28117 = ~n2790 & ~n27998;
  assign n28118 = n2790 & ~n27975;
  assign n28119 = n2827 & ~n28118;
  assign n28120 = ~n28117 & n28119;
  assign n28121 = ~pi222 & n28020;
  assign n28122 = ~pi223 & ~n28121;
  assign n28123 = ~n28120 & n28122;
  assign n28124 = ~n60064 & n28123;
  assign n28125 = ~n28110 & ~n28124;
  assign n28126 = ~pi299 & ~n28125;
  assign n28127 = pi39 & ~n28126;
  assign n28128 = ~n28102 & n28127;
  assign n28129 = n7322 & n27802;
  assign n28130 = ~n27725 & ~n28129;
  assign n28131 = ~pi224 & ~n28130;
  assign n28132 = n7322 & ~n27802;
  assign n28133 = ~n26688 & n27723;
  assign n28134 = ~n28132 & n28133;
  assign n28135 = ~n28131 & ~n28134;
  assign n28136 = ~pi299 & ~n28135;
  assign n28137 = ~pi614 & n6796;
  assign n28138 = ~n26702 & ~n28137;
  assign n28139 = pi224 & ~n28138;
  assign n28140 = ~pi224 & ~n7330;
  assign n28141 = ~n27729 & n28140;
  assign n28142 = ~n28139 & ~n28141;
  assign n28143 = n27802 & ~n28142;
  assign n28144 = n27731 & ~n27802;
  assign n28145 = pi299 & ~n28144;
  assign n28146 = ~n28143 & n28145;
  assign n28147 = ~n28136 & ~n28146;
  assign n28148 = ~pi39 & ~n28147;
  assign n28149 = ~pi38 & ~n28148;
  assign n28150 = ~n28128 & n28149;
  assign n28151 = pi662 & n6914;
  assign n28152 = n6863 & n28151;
  assign n28153 = n27743 & ~n28152;
  assign n28154 = n59132 & ~n28153;
  assign n28155 = ~n28150 & n28154;
  assign n28156 = ~n27606 & ~n28155;
  assign n28157 = ~pi625 & n28156;
  assign n28158 = pi625 & n27746;
  assign n28159 = ~pi1153 & ~n28158;
  assign n28160 = ~n28157 & n28159;
  assign n28161 = ~pi608 & ~n27898;
  assign n28162 = ~n28160 & n28161;
  assign n28163 = pi625 & n28156;
  assign n28164 = ~pi625 & n27746;
  assign n28165 = pi1153 & ~n28164;
  assign n28166 = ~n28163 & n28165;
  assign n28167 = pi608 & ~n27902;
  assign n28168 = ~n28166 & n28167;
  assign n28169 = ~n28162 & ~n28168;
  assign n28170 = pi778 & ~n28169;
  assign n28171 = ~pi778 & n28156;
  assign n28172 = ~n28170 & ~n28171;
  assign n28173 = ~pi609 & ~n28172;
  assign n28174 = pi609 & n27905;
  assign n28175 = ~pi1155 & ~n28174;
  assign n28176 = ~n28173 & n28175;
  assign n28177 = ~pi660 & ~n27756;
  assign n28178 = ~n28176 & n28177;
  assign n28179 = pi609 & ~n28172;
  assign n28180 = ~pi609 & n27905;
  assign n28181 = pi1155 & ~n28180;
  assign n28182 = ~n28179 & n28181;
  assign n28183 = pi660 & ~n27760;
  assign n28184 = ~n28182 & n28183;
  assign n28185 = ~n28178 & ~n28184;
  assign n28186 = pi785 & ~n28185;
  assign n28187 = ~pi785 & ~n28172;
  assign n28188 = ~n28186 & ~n28187;
  assign n28189 = ~pi618 & ~n28188;
  assign n28190 = pi618 & n60052;
  assign n28191 = ~pi1154 & ~n28190;
  assign n28192 = ~n28189 & n28191;
  assign n28193 = ~pi627 & ~n27768;
  assign n28194 = ~n28192 & n28193;
  assign n28195 = pi618 & ~n28188;
  assign n28196 = ~pi618 & n60052;
  assign n28197 = pi1154 & ~n28196;
  assign n28198 = ~n28195 & n28197;
  assign n28199 = pi627 & ~n27772;
  assign n28200 = ~n28198 & n28199;
  assign n28201 = ~n28194 & ~n28200;
  assign n28202 = pi781 & ~n28201;
  assign n28203 = ~pi781 & ~n28188;
  assign n28204 = ~n28202 & ~n28203;
  assign n28205 = ~pi619 & ~n28204;
  assign n28206 = pi619 & n60053;
  assign n28207 = ~pi1159 & ~n28206;
  assign n28208 = ~n28205 & n28207;
  assign n28209 = ~pi648 & ~n27780;
  assign n28210 = ~n28208 & n28209;
  assign n28211 = pi619 & ~n28204;
  assign n28212 = ~pi619 & n60053;
  assign n28213 = pi1159 & ~n28212;
  assign n28214 = ~n28211 & n28213;
  assign n28215 = pi648 & ~n27784;
  assign n28216 = ~n28214 & n28215;
  assign n28217 = pi789 & ~n28216;
  assign n28218 = pi789 & ~n28210;
  assign n28219 = ~n28216 & n28218;
  assign n28220 = ~n28210 & n28217;
  assign n28221 = ~pi789 & n28204;
  assign n28222 = n59242 & ~n28221;
  assign n28223 = ~n60065 & n28222;
  assign n28224 = pi626 & ~n27787;
  assign n28225 = ~pi626 & n27604;
  assign n28226 = n7759 & ~n28225;
  assign n28227 = ~n28224 & n28226;
  assign n28228 = n7716 & ~n27604;
  assign n28229 = ~n27917 & ~n28228;
  assign n28230 = n7984 & ~n28229;
  assign n28231 = ~pi626 & ~n27787;
  assign n28232 = pi626 & n27604;
  assign n28233 = n7760 & ~n28232;
  assign n28234 = ~n28231 & n28233;
  assign n28235 = ~n28230 & ~n28234;
  assign n28236 = ~n28227 & ~n28230;
  assign n28237 = ~n28234 & n28236;
  assign n28238 = ~n28227 & n28235;
  assign n28239 = pi788 & ~n60066;
  assign n28240 = ~n59357 & ~n28239;
  assign n28241 = ~n28223 & n28240;
  assign n28242 = ~n27950 & ~n28241;
  assign n28243 = ~n8108 & ~n28242;
  assign n28244 = ~n27938 & ~n28243;
  assign n28245 = ~pi644 & n28244;
  assign n28246 = ~pi787 & n60054;
  assign n28247 = ~n27929 & ~n27934;
  assign n28248 = pi787 & ~n28247;
  assign n28249 = ~n28246 & ~n28248;
  assign n28250 = pi644 & n28249;
  assign n28251 = ~pi715 & ~n28250;
  assign n28252 = ~n28245 & n28251;
  assign n28253 = ~n12602 & ~n27604;
  assign n28254 = n11491 & n27788;
  assign n28255 = n7835 & ~n27604;
  assign n28256 = ~n7835 & n27796;
  assign n28257 = ~n28255 & ~n28256;
  assign n28258 = ~n28253 & ~n28254;
  assign n28259 = ~pi644 & ~n60067;
  assign n28260 = pi644 & ~n27604;
  assign n28261 = pi715 & ~n28260;
  assign n28262 = ~n28259 & n28261;
  assign n28263 = ~pi1160 & ~n28262;
  assign n28264 = ~n28252 & n28263;
  assign n28265 = pi644 & n28244;
  assign n28266 = ~pi644 & n28249;
  assign n28267 = pi715 & ~n28266;
  assign n28268 = ~n28265 & n28267;
  assign n28269 = pi644 & ~n60067;
  assign n28270 = ~pi644 & ~n27604;
  assign n28271 = ~pi715 & ~n28270;
  assign n28272 = ~n28269 & n28271;
  assign n28273 = pi1160 & ~n28272;
  assign n28274 = ~n28268 & n28273;
  assign n28275 = ~n28264 & ~n28274;
  assign n28276 = pi790 & ~n28275;
  assign n28277 = ~pi790 & n28244;
  assign n28278 = ~n28276 & ~n28277;
  assign n28279 = n58992 & ~n28278;
  assign n28280 = ~pi224 & ~n58992;
  assign po381 = ~n28279 & ~n28280;
  assign n28282 = pi57 & pi59;
  assign n28283 = ~pi55 & n6311;
  assign n28284 = n2634 & n59132;
  assign n28285 = ~pi39 & n59292;
  assign n28286 = n58815 & n6309;
  assign n28287 = ~pi87 & n58816;
  assign n28288 = n2439 & n60069;
  assign n28289 = n58815 & n6311;
  assign n28290 = ~pi55 & n28288;
  assign n28291 = n58815 & n28283;
  assign n28292 = n4437 & n60070;
  assign n28293 = n58822 & n28292;
  assign n28294 = ~n4438 & ~n28293;
  assign n28295 = ~n28282 & ~n28294;
  assign n28296 = ~pi95 & n58815;
  assign n28297 = n58815 & n58822;
  assign n28298 = n2661 & n28296;
  assign n28299 = ~pi54 & n6310;
  assign n28300 = n60071 & n28299;
  assign n28301 = pi74 & ~n28300;
  assign n28302 = n59171 & n59291;
  assign n28303 = pi75 & ~n28302;
  assign n28304 = n2635 & n9186;
  assign n28305 = n2636 & n6309;
  assign n28306 = n59171 & n60072;
  assign n28307 = pi92 & ~n28306;
  assign n28308 = ~n28303 & ~n28307;
  assign n28309 = pi38 & ~n59171;
  assign n28310 = pi145 & pi180;
  assign n28311 = pi181 & pi182;
  assign n28312 = n28310 & n28311;
  assign n28313 = pi95 & ~pi479;
  assign n28314 = n2661 & n28313;
  assign n28315 = ~pi51 & n59135;
  assign n28316 = n2579 & n59136;
  assign n28317 = n58801 & n60073;
  assign n28318 = pi72 & ~n28317;
  assign n28319 = n2621 & ~n28318;
  assign n28320 = pi70 & ~n2593;
  assign n28321 = n2653 & ~n28320;
  assign n28322 = pi841 & n2526;
  assign n28323 = pi93 & ~n28322;
  assign n28324 = ~pi35 & ~n28323;
  assign n28325 = pi90 & ~n58801;
  assign n28326 = ~pi91 & ~pi314;
  assign n28327 = pi46 & n2493;
  assign n28328 = pi46 & ~pi97;
  assign n28329 = n2746 & n28328;
  assign n28330 = n58833 & n28327;
  assign n28331 = n2446 & n2515;
  assign n28332 = ~pi60 & n58794;
  assign n28333 = pi53 & ~n60075;
  assign n28334 = pi60 & n58794;
  assign n28335 = ~pi53 & ~n28334;
  assign n28336 = pi50 & ~n58831;
  assign n28337 = ~pi60 & ~n28336;
  assign n28338 = pi77 & n2733;
  assign n28339 = ~pi50 & ~n28338;
  assign n28340 = pi69 & ~n2466;
  assign n28341 = pi83 & ~n58782;
  assign n28342 = ~pi103 & ~n28341;
  assign n28343 = ~n28340 & n28342;
  assign n28344 = n2455 & n2460;
  assign n28345 = ~pi84 & n28344;
  assign n28346 = ~pi68 & ~pi111;
  assign n28347 = pi82 & n28346;
  assign n28348 = ~pi68 & n28345;
  assign n28349 = pi82 & ~pi111;
  assign n28350 = n28348 & n28349;
  assign n28351 = n28345 & n28347;
  assign n28352 = pi66 & pi73;
  assign n28353 = ~n2455 & ~n2460;
  assign n28354 = ~n28352 & ~n28353;
  assign n28355 = pi85 & pi106;
  assign n28356 = n2448 & ~n28355;
  assign n28357 = pi61 & pi76;
  assign n28358 = n2449 & ~n28357;
  assign n28359 = ~n28356 & ~n28358;
  assign n28360 = ~pi48 & ~n28359;
  assign n28361 = ~n2450 & ~n28360;
  assign n28362 = pi89 & ~n2451;
  assign n28363 = ~pi49 & ~n28362;
  assign n28364 = ~n28361 & n28363;
  assign n28365 = ~n2452 & ~n28364;
  assign n28366 = pi104 & ~n2453;
  assign n28367 = ~pi45 & ~n28366;
  assign n28368 = ~n28365 & n28367;
  assign n28369 = ~n2454 & ~n28368;
  assign n28370 = ~n2455 & ~n28369;
  assign n28371 = pi85 & n28370;
  assign n28372 = n2460 & ~n28371;
  assign n28373 = n28354 & ~n28372;
  assign n28374 = n2456 & ~n28373;
  assign n28375 = pi84 & ~n28344;
  assign n28376 = pi68 & ~n28345;
  assign n28377 = ~n28375 & ~n28376;
  assign n28378 = ~n28374 & n28377;
  assign n28379 = n2457 & n28378;
  assign n28380 = ~n60076 & ~n28379;
  assign n28381 = n6320 & ~n28380;
  assign n28382 = pi67 & n58781;
  assign n28383 = n6324 & ~n28382;
  assign n28384 = ~n28381 & n28383;
  assign n28385 = n28343 & ~n28384;
  assign n28386 = ~pi71 & ~n28385;
  assign n28387 = pi71 & ~n2469;
  assign n28388 = ~pi65 & ~n28387;
  assign n28389 = ~pi64 & n2446;
  assign n28390 = n28388 & n28389;
  assign n28391 = ~n28386 & n28390;
  assign n28392 = ~pi81 & ~n28391;
  assign n28393 = ~pi83 & pi103;
  assign n28394 = pi103 & n6324;
  assign n28395 = n2466 & n28394;
  assign n28396 = n58782 & n28393;
  assign n28397 = n28390 & n60077;
  assign n28398 = n28392 & ~n28397;
  assign n28399 = pi81 & ~n2520;
  assign n28400 = ~pi102 & ~n28399;
  assign n28401 = n2470 & n28400;
  assign n28402 = ~pi77 & n28401;
  assign n28403 = n2472 & n28400;
  assign n28404 = ~n28398 & n60078;
  assign n28405 = n28339 & ~n28404;
  assign n28406 = n28337 & ~n28405;
  assign n28407 = n28335 & ~n28406;
  assign n28408 = ~n28333 & ~n28407;
  assign n28409 = ~pi86 & ~n28408;
  assign n28410 = pi86 & ~n58834;
  assign n28411 = ~pi94 & ~n28410;
  assign n28412 = n58787 & n28411;
  assign n28413 = ~n28409 & n28412;
  assign n28414 = ~n60074 & ~n28413;
  assign n28415 = n2533 & ~n28414;
  assign n28416 = n28326 & ~n28415;
  assign n28417 = pi91 & ~n58800;
  assign n28418 = ~pi58 & ~n28417;
  assign n28419 = ~pi91 & pi314;
  assign n28420 = ~n28392 & n60078;
  assign n28421 = n28339 & ~n28420;
  assign n28422 = n28337 & ~n28421;
  assign n28423 = n28335 & ~n28422;
  assign n28424 = ~n28333 & ~n28423;
  assign n28425 = ~pi86 & ~n28424;
  assign n28426 = n28412 & ~n28425;
  assign n28427 = ~n60074 & ~n28426;
  assign n28428 = n2533 & ~n28427;
  assign n28429 = n28419 & ~n28428;
  assign n28430 = n28418 & ~n28429;
  assign n28431 = ~n28416 & n28430;
  assign n28432 = ~pi90 & ~n28431;
  assign n28433 = ~n28325 & ~n28432;
  assign n28434 = ~pi93 & ~n28433;
  assign n28435 = n28324 & ~n28434;
  assign n28436 = ~pi70 & ~n28435;
  assign n28437 = n28321 & ~n28436;
  assign n28438 = ~pi72 & ~n28437;
  assign n28439 = n28319 & ~n28438;
  assign n28440 = ~n28314 & ~n28439;
  assign n28441 = pi32 & n6426;
  assign n28442 = ~pi95 & n28441;
  assign n28443 = ~pi198 & n28442;
  assign n28444 = n28440 & ~n28443;
  assign n28445 = n2680 & ~n28444;
  assign n28446 = n28312 & n28445;
  assign n28447 = pi109 & ~n2548;
  assign n28448 = n2540 & ~n28447;
  assign n28449 = ~pi109 & ~n60074;
  assign n28450 = ~n28413 & n28449;
  assign n28451 = n28448 & ~n28450;
  assign n28452 = n28326 & ~n28451;
  assign n28453 = ~n28426 & n28449;
  assign n28454 = n28448 & ~n28453;
  assign n28455 = n28419 & ~n28454;
  assign n28456 = n28418 & ~n28455;
  assign n28457 = ~n28452 & n28456;
  assign n28458 = ~pi90 & ~n28457;
  assign n28459 = ~n28325 & ~n28458;
  assign n28460 = ~pi93 & ~n28459;
  assign n28461 = n28324 & ~n28460;
  assign n28462 = ~pi70 & ~n28461;
  assign n28463 = n28321 & ~n28462;
  assign n28464 = ~pi72 & ~n28463;
  assign n28465 = n28319 & ~n28464;
  assign n28466 = ~n28314 & ~n28465;
  assign n28467 = ~n28443 & n28466;
  assign n28468 = ~n28312 & ~n28467;
  assign n28469 = ~n2680 & ~n28467;
  assign n28470 = ~pi299 & ~n28469;
  assign n28471 = ~n28468 & n28470;
  assign n28472 = ~n28446 & n28471;
  assign n28473 = pi160 & pi197;
  assign n28474 = ~pi210 & n28442;
  assign n28475 = n28440 & ~n28474;
  assign n28476 = n2680 & ~n28475;
  assign n28477 = n28473 & ~n28476;
  assign n28478 = n28466 & ~n28474;
  assign n28479 = ~n28473 & n28478;
  assign n28480 = ~n28477 & ~n28479;
  assign n28481 = ~n2680 & ~n28478;
  assign n28482 = pi158 & pi159;
  assign n28483 = pi299 & n28482;
  assign n28484 = ~n28481 & n28483;
  assign n28485 = ~n28480 & n28484;
  assign n28486 = pi299 & n28478;
  assign n28487 = ~n28482 & n28486;
  assign n28488 = pi232 & ~n28487;
  assign n28489 = ~n28485 & n28488;
  assign n28490 = ~n28472 & n28488;
  assign n28491 = ~n28485 & n28490;
  assign n28492 = ~n28472 & n28489;
  assign n28493 = ~pi299 & n28467;
  assign n28494 = ~pi232 & ~n28486;
  assign n28495 = ~n28493 & n28494;
  assign n28496 = ~pi39 & ~n28495;
  assign n28497 = ~n28472 & ~n28485;
  assign n28498 = pi232 & ~n28497;
  assign n28499 = ~n28486 & ~n28493;
  assign n28500 = ~n28488 & ~n28499;
  assign n28501 = ~n28498 & ~n28500;
  assign n28502 = ~pi39 & ~n28501;
  assign n28503 = ~n60079 & n28496;
  assign n28504 = ~pi829 & ~n2692;
  assign n28505 = pi1091 & ~n28504;
  assign n28506 = n2807 & n58849;
  assign n28507 = ~n28505 & n28506;
  assign n28508 = ~pi216 & ~n28507;
  assign n28509 = ~pi1091 & n28506;
  assign n28510 = pi1091 & n2692;
  assign n28511 = n2441 & ~n28510;
  assign n28512 = n2862 & n28511;
  assign n28513 = n58849 & ~n28510;
  assign n28514 = ~n58838 & ~n60081;
  assign n28515 = pi1091 & ~n28514;
  assign n28516 = n2807 & n28515;
  assign n28517 = ~n28509 & ~n28516;
  assign n28518 = pi216 & n28517;
  assign n28519 = pi216 & ~n28517;
  assign n28520 = ~pi216 & n28507;
  assign n28521 = ~n28519 & ~n28520;
  assign n28522 = ~n28508 & ~n28518;
  assign n28523 = n2852 & ~n60082;
  assign n28524 = pi299 & ~n2845;
  assign n28525 = n28523 & n28524;
  assign n28526 = pi224 & ~n28517;
  assign n28527 = ~pi224 & n28507;
  assign n28528 = ~pi224 & ~n28507;
  assign n28529 = pi224 & n28517;
  assign n28530 = ~n28528 & ~n28529;
  assign n28531 = ~n28526 & ~n28527;
  assign n28532 = ~pi299 & ~n2792;
  assign n28533 = n2829 & n28532;
  assign n28534 = pi222 & ~n2792;
  assign n28535 = n2828 & n28534;
  assign n28536 = ~n2792 & n58844;
  assign n28537 = n2829 & ~n28528;
  assign n28538 = n2829 & n60083;
  assign n28539 = ~n28529 & n28537;
  assign n28540 = n28532 & n60085;
  assign n28541 = n60083 & n60084;
  assign n28542 = pi39 & ~n60086;
  assign n28543 = ~n28525 & n28542;
  assign n28544 = ~n60080 & ~n28543;
  assign n28545 = ~pi38 & ~n28544;
  assign n28546 = ~n28309 & ~n28545;
  assign n28547 = ~pi100 & ~n28546;
  assign n28548 = ~pi38 & pi100;
  assign n28549 = n59171 & n28548;
  assign n28550 = ~pi252 & n58822;
  assign n28551 = ~pi142 & ~n2674;
  assign n28552 = ~pi299 & n28551;
  assign n28553 = ~pi146 & ~n2677;
  assign n28554 = pi299 & n28553;
  assign n28555 = pi146 & n2678;
  assign n28556 = pi142 & n2675;
  assign n28557 = ~n28555 & ~n28556;
  assign n28558 = ~n2679 & n28557;
  assign n28559 = ~n28552 & ~n28554;
  assign n28560 = n28550 & ~n60087;
  assign n28561 = ~pi683 & ~n2707;
  assign n28562 = ~pi250 & ~po740;
  assign n28563 = pi129 & pi250;
  assign n28564 = ~n28562 & ~n28563;
  assign n28565 = ~n28561 & ~n28564;
  assign n28566 = n60087 & ~n28565;
  assign n28567 = n2707 & n60087;
  assign n28568 = ~n28566 & ~n28567;
  assign n28569 = ~n28550 & ~n60087;
  assign n28570 = ~n2707 & n60087;
  assign n28571 = n28565 & n28570;
  assign n28572 = ~n28569 & ~n28571;
  assign n28573 = ~n28560 & n28568;
  assign n28574 = n28549 & n60088;
  assign n28575 = ~pi38 & n59171;
  assign n28576 = pi100 & ~n28575;
  assign n28577 = ~pi87 & ~n28576;
  assign n28578 = ~pi87 & ~n28574;
  assign n28579 = ~n28576 & n28578;
  assign n28580 = ~n28574 & n28577;
  assign n28581 = ~n28547 & n60089;
  assign n28582 = n6307 & ~n28581;
  assign n28583 = n28308 & ~n28582;
  assign n28584 = ~pi54 & ~n28583;
  assign n28585 = ~pi92 & n28306;
  assign n28586 = pi54 & ~n28585;
  assign n28587 = ~n28584 & ~n28586;
  assign n28588 = ~pi74 & ~n28587;
  assign n28589 = ~n28301 & ~n28588;
  assign n28590 = ~pi55 & ~n28589;
  assign n28591 = n6311 & n60071;
  assign n28592 = ~pi74 & n28300;
  assign n28593 = n58822 & n28288;
  assign n28594 = pi55 & ~n60090;
  assign n28595 = ~pi56 & ~n28594;
  assign n28596 = ~pi62 & n28595;
  assign n28597 = ~n28590 & n28596;
  assign n28598 = n4438 & ~n28597;
  assign po195 = n28295 & ~n28598;
  assign n28600 = ~pi954 & ~po195;
  assign n28601 = pi24 & pi954;
  assign po182 = ~n28600 & ~n28601;
  assign n28603 = ~pi31 & ~pi80;
  assign n28604 = pi818 & n28603;
  assign n28605 = ~n2439 & n3871;
  assign n28606 = ~n3213 & ~n28605;
  assign n28607 = ~pi120 & ~n2439;
  assign n28608 = ~pi1093 & n28607;
  assign n28609 = n28606 & ~n28608;
  assign n28610 = n58822 & n2710;
  assign n28611 = pi120 & ~n3871;
  assign n28612 = ~n2718 & n28611;
  assign n28613 = ~pi120 & pi1093;
  assign n28614 = pi120 & n2718;
  assign n28615 = n2718 & ~n28613;
  assign n28616 = ~pi120 & n28610;
  assign n28617 = ~n60091 & ~n28616;
  assign n28618 = n28610 & ~n28612;
  assign n28619 = n2720 & ~n60092;
  assign n28620 = ~pi1091 & n5304;
  assign n28621 = n28613 & ~n28620;
  assign n28622 = ~n28611 & ~n28621;
  assign n28623 = pi100 & ~n28622;
  assign n28624 = ~n28619 & n28623;
  assign n28625 = ~pi1093 & n2631;
  assign n28626 = pi120 & n28625;
  assign n28627 = ~pi39 & ~n28626;
  assign n28628 = pi97 & ~n58833;
  assign n28629 = ~pi108 & ~n28628;
  assign n28630 = ~pi110 & n28629;
  assign n28631 = ~pi46 & ~pi109;
  assign n28632 = n2492 & n28631;
  assign n28633 = ~n2582 & n28632;
  assign n28634 = n28630 & n28633;
  assign n28635 = ~n2732 & ~n28634;
  assign n28636 = n2445 & ~n28635;
  assign n28637 = n2556 & ~n28636;
  assign n28638 = n2529 & ~n28637;
  assign n28639 = ~pi51 & ~n28638;
  assign n28640 = ~n2596 & ~n28639;
  assign n28641 = ~pi96 & ~n28640;
  assign n28642 = n58837 & ~n28641;
  assign n28643 = n58811 & n2727;
  assign n28644 = ~pi829 & n28643;
  assign n28645 = ~pi122 & ~n28644;
  assign n28646 = ~n28642 & n28645;
  assign n28647 = pi122 & ~n2610;
  assign n28648 = ~n2692 & ~n28647;
  assign n28649 = ~n28646 & n28648;
  assign n28650 = n2797 & ~n28649;
  assign n28651 = n2878 & ~n28643;
  assign n28652 = ~n5304 & n28651;
  assign n28653 = ~n28650 & ~n28652;
  assign n28654 = n28627 & n28653;
  assign n28655 = ~n2783 & n28622;
  assign n28656 = ~n58842 & n28611;
  assign n28657 = pi1091 & pi1092;
  assign n28658 = n58840 & n28657;
  assign n28659 = n2793 & n58839;
  assign n28660 = n28621 & ~n60093;
  assign n28661 = ~n28656 & ~n28660;
  assign n28662 = n2783 & n28661;
  assign n28663 = ~n28655 & ~n28662;
  assign n28664 = n58846 & n28663;
  assign n28665 = n2822 & ~n28622;
  assign n28666 = ~n2822 & ~n28661;
  assign n28667 = ~n28665 & ~n28666;
  assign n28668 = ~n58846 & ~n28667;
  assign n28669 = n3906 & ~n28668;
  assign n28670 = n3906 & ~n28664;
  assign n28671 = ~n28668 & n28670;
  assign n28672 = ~n28664 & n28669;
  assign n28673 = ~n3906 & n28622;
  assign n28674 = pi299 & ~n28673;
  assign n28675 = ~n60094 & n28674;
  assign n28676 = n2790 & n28663;
  assign n28677 = ~n2790 & ~n28667;
  assign n28678 = n3890 & ~n28677;
  assign n28679 = n3890 & ~n28676;
  assign n28680 = ~n28677 & n28679;
  assign n28681 = ~n28676 & n28678;
  assign n28682 = ~n3890 & n28622;
  assign n28683 = ~pi299 & ~n28682;
  assign n28684 = ~n60095 & n28683;
  assign n28685 = pi39 & ~n28684;
  assign n28686 = pi39 & ~n28675;
  assign n28687 = ~n28684 & n28686;
  assign n28688 = ~n28675 & n28685;
  assign n28689 = ~n28654 & ~n60096;
  assign n28690 = ~pi38 & ~n28689;
  assign n28691 = ~pi120 & ~pi1093;
  assign n28692 = pi38 & n28691;
  assign n28693 = ~pi100 & ~n28692;
  assign n28694 = ~n3923 & n28693;
  assign n28695 = ~n28690 & n28694;
  assign n28696 = ~n28624 & ~n28695;
  assign n28697 = ~pi87 & ~n28696;
  assign n28698 = n2886 & ~n28691;
  assign n28699 = n2878 & ~n5304;
  assign n28700 = ~n3941 & n28699;
  assign n28701 = n2884 & ~n28700;
  assign n28702 = ~n58815 & n3871;
  assign n28703 = pi87 & ~n28702;
  assign n28704 = ~n28701 & n28703;
  assign n28705 = n28698 & n28704;
  assign n28706 = ~n28697 & ~n28705;
  assign n28707 = ~pi75 & ~n28706;
  assign n28708 = n2682 & n28622;
  assign n28709 = ~n2711 & n28621;
  assign n28710 = ~pi1091 & ~n3870;
  assign n28711 = ~n3863 & ~n28710;
  assign n28712 = pi120 & ~n28711;
  assign n28713 = ~n2682 & ~n28712;
  assign n28714 = ~n28709 & n28713;
  assign n28715 = ~n28708 & ~n28714;
  assign n28716 = n2672 & ~n28715;
  assign n28717 = ~n2672 & n28622;
  assign n28718 = pi75 & ~n28717;
  assign n28719 = ~n28716 & n28718;
  assign n28720 = n2439 & ~n28719;
  assign n28721 = ~n28707 & n28720;
  assign n28722 = n28609 & ~n28721;
  assign n28723 = ~n28650 & ~n28651;
  assign n28724 = n28627 & n28723;
  assign n28725 = pi299 & ~n28691;
  assign n28726 = ~n58975 & n28725;
  assign n28727 = ~pi299 & ~n28691;
  assign n28728 = ~n58982 & n28727;
  assign n28729 = pi39 & ~n28728;
  assign n28730 = pi39 & ~n28726;
  assign n28731 = ~n28728 & n28730;
  assign n28732 = ~n28726 & n28729;
  assign n28733 = ~n28724 & ~n60097;
  assign n28734 = ~pi38 & ~n28733;
  assign n28735 = n28693 & ~n28734;
  assign n28736 = pi100 & ~n28691;
  assign n28737 = ~n28619 & n28736;
  assign n28738 = ~n28735 & ~n28737;
  assign n28739 = ~pi87 & ~n28738;
  assign n28740 = ~n28698 & ~n28739;
  assign n28741 = ~pi75 & ~n28740;
  assign n28742 = n2714 & ~n28691;
  assign n28743 = n2439 & ~n28742;
  assign n28744 = ~n28741 & n28743;
  assign n28745 = n3213 & ~n28608;
  assign n28746 = ~n28744 & n28745;
  assign n28747 = ~n28722 & ~n28746;
  assign n28748 = n28604 & ~n28747;
  assign n28749 = n58992 & ~n28748;
  assign n28750 = ~n3213 & n28622;
  assign n28751 = pi120 & ~n28750;
  assign n28752 = n28604 & ~n28691;
  assign n28753 = ~n28750 & n28752;
  assign n28754 = ~n58992 & ~n28753;
  assign n28755 = ~n28751 & n28754;
  assign n28756 = ~n5138 & ~n28755;
  assign n28757 = pi951 & pi982;
  assign n28758 = pi1092 & n28757;
  assign n28759 = pi1093 & n28758;
  assign n28760 = ~pi120 & ~n28759;
  assign n28761 = ~n28750 & ~n28760;
  assign n28762 = n28754 & ~n28761;
  assign n28763 = n5138 & ~n28762;
  assign n28764 = ~n28756 & ~n28763;
  assign n28765 = ~n28749 & ~n28764;
  assign n28766 = pi120 & n2712;
  assign n28767 = ~pi1091 & n28759;
  assign n28768 = ~pi120 & ~n28767;
  assign n28769 = n2797 & n28758;
  assign n28770 = ~pi24 & ~pi90;
  assign n28771 = pi950 & n2440;
  assign n28772 = ~pi122 & n2795;
  assign n28773 = n28770 & n60098;
  assign n28774 = n2684 & n28773;
  assign n28775 = n6346 & n28770;
  assign n28776 = n60098 & n28775;
  assign n28777 = ~pi93 & ~pi122;
  assign n28778 = n2600 & n28777;
  assign n28779 = n2795 & n28770;
  assign n28780 = n28778 & n28779;
  assign n28781 = n2614 & n28780;
  assign n28782 = n59136 & n28776;
  assign n28783 = n2684 & n60099;
  assign n28784 = n59137 & n28774;
  assign n28785 = n2708 & n60100;
  assign n28786 = n58801 & n28785;
  assign n28787 = n28769 & ~n28786;
  assign n28788 = n28768 & ~n28787;
  assign n28789 = ~n28766 & ~n28788;
  assign n28790 = ~n2682 & ~n28789;
  assign n28791 = n2682 & n28760;
  assign n28792 = n2672 & ~n28791;
  assign n28793 = ~n28790 & n28792;
  assign n28794 = ~n2672 & ~n28760;
  assign n28795 = pi75 & ~n28794;
  assign n28796 = ~n28793 & n28795;
  assign n28797 = n2440 & n2708;
  assign n28798 = n2873 & n28797;
  assign n28799 = n28769 & ~n28798;
  assign n28800 = n28768 & ~n28799;
  assign n28801 = ~n60091 & ~n28800;
  assign n28802 = ~pi39 & n2719;
  assign n28803 = ~n28801 & n28802;
  assign n28804 = pi100 & ~n28803;
  assign n28805 = ~pi38 & ~n28804;
  assign n28806 = ~n2720 & n28760;
  assign n28807 = ~n28805 & ~n28806;
  assign n28808 = ~n28625 & n28723;
  assign n28809 = pi120 & n28808;
  assign n28810 = n58836 & ~n28641;
  assign n28811 = n2440 & n28758;
  assign n28812 = ~n28810 & n28811;
  assign n28813 = pi950 & n58810;
  assign n28814 = ~n2588 & n28813;
  assign n28815 = pi122 & n2761;
  assign n28816 = pi122 & n28757;
  assign n28817 = n2761 & n28816;
  assign n28818 = n28757 & n28815;
  assign n28819 = ~n28814 & n60101;
  assign n28820 = pi824 & n28814;
  assign n28821 = n28758 & ~n28820;
  assign n28822 = ~pi829 & n28821;
  assign n28823 = ~n28819 & ~n28822;
  assign n28824 = ~n28812 & n28823;
  assign n28825 = n2726 & ~n28824;
  assign n28826 = n2692 & n28759;
  assign n28827 = n2880 & n28758;
  assign n28828 = ~n28825 & ~n60102;
  assign n28829 = pi1091 & ~n28828;
  assign n28830 = n2878 & n28821;
  assign n28831 = n28767 & ~n28820;
  assign n28832 = ~pi120 & ~n60103;
  assign n28833 = ~n28829 & n28832;
  assign n28834 = ~pi39 & ~n28833;
  assign n28835 = ~pi39 & ~n28809;
  assign n28836 = ~n28833 & n28835;
  assign n28837 = ~n28809 & n28834;
  assign n28838 = pi39 & ~n28760;
  assign n28839 = ~n3890 & n28760;
  assign n28840 = ~pi299 & ~n28839;
  assign n28841 = ~n2819 & ~n28760;
  assign n28842 = n2790 & n28841;
  assign n28843 = ~n2823 & ~n28760;
  assign n28844 = ~n2790 & n28843;
  assign n28845 = n3890 & ~n28844;
  assign n28846 = ~n28842 & n28845;
  assign n28847 = n28840 & ~n28846;
  assign n28848 = n58846 & n28841;
  assign n28849 = ~n58846 & n28843;
  assign n28850 = n3906 & ~n28849;
  assign n28851 = ~n28848 & n28850;
  assign n28852 = ~n3906 & n28760;
  assign n28853 = pi299 & ~n28852;
  assign n28854 = ~n28851 & n28853;
  assign n28855 = ~n28847 & ~n28854;
  assign n28856 = pi39 & ~n28855;
  assign n28857 = n4293 & n28838;
  assign n28858 = ~n60104 & ~n60105;
  assign n28859 = n2636 & ~n28858;
  assign n28860 = ~n28807 & ~n28859;
  assign n28861 = ~pi87 & ~n28860;
  assign n28862 = ~n58815 & n28760;
  assign n28863 = pi87 & ~n28862;
  assign n28864 = n2873 & n6472;
  assign n28865 = n28769 & ~n28864;
  assign n28866 = ~n58851 & n28767;
  assign n28867 = ~n28865 & ~n28866;
  assign n28868 = ~pi120 & ~n28867;
  assign n28869 = ~n2879 & ~n2883;
  assign n28870 = pi120 & ~n28869;
  assign n28871 = n58815 & ~n28870;
  assign n28872 = ~n28868 & n28871;
  assign n28873 = n28863 & ~n28872;
  assign n28874 = ~pi75 & ~n28873;
  assign n28875 = ~n28861 & n28874;
  assign n28876 = ~n28796 & ~n28875;
  assign n28877 = n2439 & ~n28876;
  assign n28878 = n3213 & ~n28877;
  assign n28879 = ~n5304 & n28767;
  assign n28880 = ~n28799 & ~n28879;
  assign n28881 = ~pi120 & ~n28880;
  assign n28882 = ~n28612 & ~n28881;
  assign n28883 = n2719 & ~n28882;
  assign n28884 = ~n28622 & ~n28760;
  assign n28885 = ~n2719 & n28884;
  assign n28886 = n2634 & ~n28885;
  assign n28887 = ~n28883 & n28886;
  assign n28888 = ~n2634 & ~n28884;
  assign n28889 = pi100 & ~n28888;
  assign n28890 = ~n28887 & n28889;
  assign n28891 = ~n28625 & n28653;
  assign n28892 = pi120 & n28891;
  assign n28893 = n28699 & n28821;
  assign n28894 = ~pi120 & ~n28893;
  assign n28895 = ~n28829 & n28894;
  assign n28896 = ~n28892 & ~n28895;
  assign n28897 = ~pi39 & ~n28896;
  assign n28898 = ~n58840 & n28769;
  assign n28899 = ~n28879 & ~n28898;
  assign n28900 = ~pi120 & ~n28899;
  assign n28901 = ~n28656 & ~n28900;
  assign n28902 = n2783 & ~n28901;
  assign n28903 = ~n2783 & n28884;
  assign n28904 = ~n28902 & ~n28903;
  assign n28905 = n2790 & ~n28904;
  assign n28906 = ~n2822 & ~n28901;
  assign n28907 = n2822 & n28884;
  assign n28908 = ~n28906 & ~n28907;
  assign n28909 = ~n2790 & ~n28908;
  assign n28910 = n3890 & ~n28909;
  assign n28911 = n3890 & ~n28905;
  assign n28912 = ~n28909 & n28911;
  assign n28913 = ~n28905 & n28910;
  assign n28914 = ~n3890 & ~n28884;
  assign n28915 = ~pi299 & ~n28914;
  assign n28916 = ~n28682 & n28840;
  assign n28917 = ~n60106 & n60107;
  assign n28918 = n58846 & ~n28904;
  assign n28919 = ~n58846 & ~n28908;
  assign n28920 = n3906 & ~n28919;
  assign n28921 = n3906 & ~n28918;
  assign n28922 = ~n28919 & n28921;
  assign n28923 = ~n28918 & n28920;
  assign n28924 = pi299 & ~n3912;
  assign n28925 = ~n3912 & n28853;
  assign n28926 = ~n28852 & n28924;
  assign n28927 = ~n60108 & n60109;
  assign n28928 = pi39 & ~n28927;
  assign n28929 = pi39 & ~n28917;
  assign n28930 = ~n28927 & n28929;
  assign n28931 = ~n28917 & n28928;
  assign n28932 = ~n28897 & ~n60110;
  assign n28933 = ~pi38 & ~n28932;
  assign n28934 = pi38 & ~n28884;
  assign n28935 = ~pi100 & ~n28934;
  assign n28936 = ~n28933 & n28935;
  assign n28937 = ~n28890 & ~n28936;
  assign n28938 = ~pi87 & ~n28937;
  assign n28939 = ~n28701 & ~n28871;
  assign n28940 = ~n28865 & ~n28879;
  assign n28941 = n28868 & ~n28940;
  assign n28942 = ~n28939 & ~n28941;
  assign n28943 = ~n28702 & n28863;
  assign n28944 = ~n28942 & n28943;
  assign n28945 = ~n28938 & ~n28944;
  assign n28946 = ~pi75 & ~n28945;
  assign n28947 = n2682 & ~n28884;
  assign n28948 = ~n28787 & ~n28879;
  assign n28949 = ~pi120 & ~n28948;
  assign n28950 = n28713 & ~n28949;
  assign n28951 = ~n28947 & ~n28950;
  assign n28952 = n2672 & ~n28951;
  assign n28953 = ~n2672 & ~n28884;
  assign n28954 = pi75 & ~n28953;
  assign n28955 = ~n28952 & n28954;
  assign n28956 = n2439 & ~n28955;
  assign n28957 = ~n28946 & n28956;
  assign n28958 = n28609 & ~n28957;
  assign n28959 = ~n28878 & ~n28958;
  assign n28960 = n28607 & ~n28759;
  assign n28961 = n28763 & ~n28960;
  assign n28962 = ~n28959 & n28961;
  assign n28963 = ~pi39 & ~n28808;
  assign n28964 = n2859 & ~n28963;
  assign n28965 = ~pi100 & ~n28964;
  assign n28966 = ~n2725 & ~n28965;
  assign n28967 = ~pi87 & ~n28966;
  assign n28968 = ~n2886 & ~n28967;
  assign n28969 = ~pi75 & ~n28968;
  assign n28970 = ~n2714 & ~n28969;
  assign n28971 = n3213 & ~n28607;
  assign n28972 = ~n28970 & n28971;
  assign n28973 = n2725 & ~n3871;
  assign n28974 = ~pi39 & ~n28891;
  assign n28975 = pi1091 & n2822;
  assign n28976 = ~n28710 & ~n28975;
  assign n28977 = ~n3884 & ~n28710;
  assign n28978 = ~n28975 & n28977;
  assign n28979 = ~n2822 & ~n28977;
  assign n28980 = n2822 & ~n3871;
  assign n28981 = ~n28979 & ~n28980;
  assign n28982 = ~n3884 & n28976;
  assign n28983 = ~n58846 & ~n60111;
  assign n28984 = pi1091 & ~n2783;
  assign n28985 = ~n28710 & ~n28984;
  assign n28986 = n28977 & ~n28984;
  assign n28987 = n2783 & ~n28977;
  assign n28988 = ~n2783 & ~n3871;
  assign n28989 = ~n28987 & ~n28988;
  assign n28990 = ~n3884 & n28985;
  assign n28991 = n58846 & ~n60112;
  assign n28992 = n3906 & ~n28991;
  assign n28993 = ~n28983 & n28992;
  assign n28994 = n28924 & ~n28993;
  assign n28995 = n2790 & ~n60112;
  assign n28996 = ~n2790 & ~n60111;
  assign n28997 = n3890 & ~n28996;
  assign n28998 = n3890 & ~n28995;
  assign n28999 = ~n28996 & n28998;
  assign n29000 = ~n28995 & n28997;
  assign n29001 = ~pi299 & ~n3900;
  assign n29002 = ~n60113 & n29001;
  assign n29003 = ~n28994 & ~n29002;
  assign n29004 = pi39 & ~n29003;
  assign n29005 = ~pi38 & ~n29004;
  assign n29006 = ~n28974 & n29005;
  assign n29007 = ~pi100 & ~n3923;
  assign n29008 = ~n29006 & n29007;
  assign n29009 = ~n28973 & ~n29008;
  assign n29010 = ~pi87 & ~n29009;
  assign n29011 = ~n28704 & ~n29010;
  assign n29012 = ~pi75 & ~n29011;
  assign n29013 = n2683 & n28711;
  assign n29014 = ~n2683 & n3871;
  assign n29015 = pi75 & ~n29014;
  assign n29016 = ~n29013 & n29015;
  assign n29017 = ~n29012 & ~n29016;
  assign n29018 = n28606 & ~n29017;
  assign n29019 = ~n2439 & ~n28750;
  assign n29020 = ~n29018 & ~n29019;
  assign n29021 = ~n28972 & n29020;
  assign n29022 = pi120 & n28756;
  assign n29023 = ~n29021 & n29022;
  assign n29024 = ~n28962 & ~n29023;
  assign n29025 = ~n28604 & ~n29024;
  assign n29026 = ~n28765 & ~n29025;
  assign n29027 = ~pi149 & ~pi157;
  assign n29028 = pi197 & n29027;
  assign n29029 = ~pi197 & ~n29027;
  assign n29030 = ~n29028 & ~n29029;
  assign n29031 = pi162 & n2680;
  assign n29032 = n29030 & ~n29031;
  assign n29033 = n29028 & n29031;
  assign n29034 = n2680 & ~n29027;
  assign n29035 = ~pi162 & ~pi197;
  assign n29036 = n29034 & ~n29035;
  assign n29037 = n2680 & ~n29036;
  assign n29038 = ~n29033 & n29037;
  assign n29039 = ~n29030 & ~n29038;
  assign n29040 = ~n29032 & ~n29039;
  assign n29041 = pi232 & ~n2635;
  assign n29042 = pi232 & n29040;
  assign n29043 = ~n2635 & n29042;
  assign n29044 = n29040 & n29041;
  assign n29045 = n2635 & n2681;
  assign n29046 = pi167 & n2681;
  assign n29047 = n2635 & n29046;
  assign n29048 = pi167 & n29045;
  assign n29049 = ~n60114 & ~n60115;
  assign n29050 = ~pi74 & n29049;
  assign n29051 = pi148 & n29045;
  assign n29052 = pi74 & ~n29051;
  assign n29053 = ~n60114 & n29052;
  assign n29054 = ~n29050 & ~n29053;
  assign n29055 = ~n4438 & n29054;
  assign n29056 = ~pi54 & ~n60114;
  assign n29057 = pi38 & n29046;
  assign n29058 = pi38 & n60115;
  assign n29059 = n2635 & n29057;
  assign n29060 = n29056 & ~n60116;
  assign n29061 = ~pi74 & n29060;
  assign n29062 = n29054 & ~n29061;
  assign n29063 = ~n4437 & ~n29062;
  assign n29064 = n4438 & ~n29063;
  assign n29065 = ~pi40 & n2446;
  assign n29066 = ~pi38 & n29065;
  assign n29067 = n2635 & n29066;
  assign n29068 = n6306 & n29067;
  assign n29069 = ~n4437 & ~n29068;
  assign n29070 = n4438 & ~n29069;
  assign n29071 = ~n29064 & ~n29070;
  assign n29072 = pi299 & ~n29040;
  assign n29073 = ~pi178 & ~pi183;
  assign n29074 = n2680 & ~n29073;
  assign n29075 = pi140 & pi145;
  assign n29076 = ~pi140 & ~pi145;
  assign n29077 = ~n29075 & ~n29076;
  assign n29078 = n29074 & ~n29077;
  assign n29079 = n29073 & ~n29075;
  assign n29080 = n2680 & ~n29076;
  assign n29081 = n29079 & n29080;
  assign n29082 = ~pi299 & ~n29081;
  assign n29083 = ~n29078 & n29082;
  assign n29084 = pi232 & ~n29083;
  assign n29085 = ~n29072 & n29084;
  assign n29086 = pi100 & ~n29085;
  assign n29087 = pi75 & ~n29085;
  assign n29088 = ~n29086 & ~n29087;
  assign n29089 = pi141 & ~pi299;
  assign n29090 = pi148 & pi299;
  assign n29091 = ~n29089 & ~n29090;
  assign n29092 = n2681 & ~n29091;
  assign n29093 = n2635 & ~n29092;
  assign n29094 = n29088 & ~n29093;
  assign n29095 = pi74 & ~n29094;
  assign n29096 = ~pi55 & ~n29095;
  assign n29097 = ~pi167 & pi299;
  assign n29098 = ~pi188 & ~pi299;
  assign n29099 = pi188 & ~pi299;
  assign n29100 = pi167 & pi299;
  assign n29101 = ~n29099 & ~n29100;
  assign n29102 = ~n29097 & ~n29098;
  assign n29103 = n2681 & ~n60117;
  assign n29104 = ~pi100 & ~n29103;
  assign n29105 = ~pi75 & n29104;
  assign n29106 = n29088 & ~n29105;
  assign n29107 = pi54 & ~n29106;
  assign n29108 = pi95 & ~n29065;
  assign n29109 = ~n28313 & ~n29108;
  assign n29110 = ~pi40 & ~pi479;
  assign n29111 = ~pi58 & n58793;
  assign n29112 = n2580 & n29111;
  assign n29113 = ~pi32 & n58817;
  assign n29114 = n29112 & n29113;
  assign n29115 = n2446 & ~n29114;
  assign n29116 = n29110 & n29115;
  assign n29117 = ~n29109 & ~n29116;
  assign n29118 = pi32 & ~n29065;
  assign n29119 = n2446 & ~n2600;
  assign n29120 = n2446 & ~n29112;
  assign n29121 = pi70 & ~n29120;
  assign n29122 = n2446 & ~n58793;
  assign n29123 = pi58 & ~n29122;
  assign n29124 = pi53 & ~n2515;
  assign n29125 = pi50 & n58831;
  assign n29126 = ~pi60 & n29125;
  assign n29127 = n28335 & ~n29126;
  assign n29128 = ~n29124 & ~n29127;
  assign n29129 = ~pi68 & n2465;
  assign n29130 = ~pi111 & n2447;
  assign n29131 = ~pi36 & ~pi82;
  assign n29132 = ~pi82 & ~pi84;
  assign n29133 = ~pi36 & n29132;
  assign n29134 = ~pi84 & n29131;
  assign n29135 = n29130 & n60118;
  assign n29136 = n29129 & n60118;
  assign n29137 = n29130 & n29136;
  assign n29138 = n29129 & n29135;
  assign n29139 = ~pi66 & pi73;
  assign n29140 = ~pi36 & n29129;
  assign n29141 = n29130 & n29140;
  assign n29142 = pi73 & ~pi82;
  assign n29143 = n6318 & n29142;
  assign n29144 = n29141 & n29143;
  assign n29145 = n60119 & n29139;
  assign n29146 = n2478 & n29139;
  assign n29147 = n60119 & n29146;
  assign n29148 = n2483 & n29147;
  assign n29149 = n58785 & n60120;
  assign n29150 = n2455 & n60121;
  assign n29151 = n2489 & n29150;
  assign n29152 = n2446 & ~n29151;
  assign n29153 = ~n29128 & n29152;
  assign n29154 = n2501 & ~n29153;
  assign n29155 = ~n2446 & ~n2501;
  assign n29156 = n58788 & ~n29155;
  assign n29157 = ~n29154 & n29156;
  assign n29158 = n2446 & ~n58788;
  assign n29159 = ~pi58 & ~n29158;
  assign n29160 = ~n29157 & n29159;
  assign n29161 = ~n29123 & ~n29160;
  assign n29162 = ~pi90 & ~n29161;
  assign n29163 = ~pi841 & n29111;
  assign n29164 = n2446 & ~n29163;
  assign n29165 = pi90 & ~n29164;
  assign n29166 = n2592 & ~n29165;
  assign n29167 = ~n29162 & n29166;
  assign n29168 = n2446 & ~n2592;
  assign n29169 = ~pi70 & ~n29168;
  assign n29170 = ~n29167 & n29169;
  assign n29171 = ~n29121 & ~n29170;
  assign n29172 = ~pi51 & ~n29171;
  assign n29173 = pi51 & ~n2446;
  assign n29174 = n2600 & ~n29173;
  assign n29175 = ~n29172 & n29174;
  assign n29176 = ~n29119 & ~n29175;
  assign n29177 = ~pi40 & ~n29176;
  assign n29178 = ~pi32 & ~n29177;
  assign n29179 = ~n29118 & ~n29178;
  assign n29180 = ~pi95 & ~n29179;
  assign n29181 = ~n29117 & ~n29180;
  assign n29182 = pi210 & pi299;
  assign n29183 = pi198 & ~pi299;
  assign n29184 = ~pi198 & ~pi299;
  assign n29185 = ~pi210 & pi299;
  assign n29186 = ~n29184 & ~n29185;
  assign n29187 = ~n29182 & ~n29183;
  assign n29188 = n59138 & n29163;
  assign n29189 = n29065 & ~n29188;
  assign n29190 = pi32 & ~n29189;
  assign n29191 = ~n29178 & ~n29190;
  assign n29192 = ~pi95 & ~n29191;
  assign n29193 = ~n60122 & n29192;
  assign n29194 = n29181 & ~n29193;
  assign n29195 = ~pi232 & ~n29194;
  assign n29196 = ~pi198 & n29192;
  assign n29197 = n29181 & ~n29196;
  assign n29198 = ~n2680 & n29197;
  assign n29199 = ~pi40 & ~n2446;
  assign n29200 = pi32 & ~n29199;
  assign n29201 = n2445 & n2592;
  assign n29202 = ~n2446 & ~n29201;
  assign n29203 = n2580 & n29160;
  assign n29204 = ~n29202 & ~n29203;
  assign n29205 = ~pi70 & ~n29204;
  assign n29206 = ~n29121 & ~n29205;
  assign n29207 = ~pi51 & ~n29206;
  assign n29208 = n29174 & ~n29207;
  assign n29209 = ~pi40 & ~n29119;
  assign n29210 = ~n29208 & n29209;
  assign n29211 = ~pi32 & ~n29210;
  assign n29212 = ~n29200 & ~n29211;
  assign n29213 = ~n2601 & ~n29065;
  assign n29214 = ~n29212 & ~n29213;
  assign n29215 = ~pi95 & ~n29214;
  assign n29216 = ~n29117 & ~n29215;
  assign n29217 = n2680 & ~n29065;
  assign n29218 = ~n29108 & ~n29215;
  assign n29219 = pi95 & ~n29199;
  assign n29220 = ~pi40 & ~n29189;
  assign n29221 = pi32 & ~n29220;
  assign n29222 = ~n29211 & ~n29221;
  assign n29223 = ~pi95 & ~n29222;
  assign n29224 = ~n29219 & ~n29223;
  assign n29225 = n29218 & ~n29224;
  assign n29226 = ~pi198 & ~n29225;
  assign n29227 = n2680 & ~n29226;
  assign n29228 = ~n29217 & ~n29227;
  assign n29229 = n29216 & ~n29228;
  assign n29230 = ~n29198 & ~n29229;
  assign n29231 = ~pi142 & ~n29230;
  assign n29232 = pi142 & n29197;
  assign n29233 = ~pi140 & ~n29232;
  assign n29234 = ~n29231 & n29233;
  assign n29235 = ~pi32 & n6403;
  assign n29236 = ~pi32 & n29150;
  assign n29237 = n6403 & n29236;
  assign n29238 = n29150 & n29235;
  assign n29239 = n29065 & ~n60123;
  assign n29240 = ~pi95 & ~n29239;
  assign n29241 = n2680 & ~n29240;
  assign n29242 = ~n29117 & n29241;
  assign n29243 = ~n29198 & ~n29242;
  assign n29244 = ~pi142 & ~n29243;
  assign n29245 = ~n2680 & ~n29197;
  assign n29246 = ~pi40 & ~n29118;
  assign n29247 = n2446 & ~n58823;
  assign n29248 = ~pi32 & ~n29247;
  assign n29249 = pi93 & ~n2446;
  assign n29250 = n58823 & ~n29249;
  assign n29251 = n2446 & ~n29123;
  assign n29252 = ~pi90 & ~n29251;
  assign n29253 = ~n29165 & ~n29252;
  assign n29254 = n58797 & n29150;
  assign n29255 = ~pi90 & n29254;
  assign n29256 = n29253 & ~n29255;
  assign n29257 = ~pi93 & ~n29256;
  assign n29258 = n29250 & ~n29257;
  assign n29259 = n29248 & ~n29258;
  assign n29260 = n29246 & ~n29259;
  assign n29261 = ~pi95 & ~n29260;
  assign n29262 = ~n29117 & ~n29261;
  assign n29263 = n2680 & ~n29262;
  assign n29264 = pi142 & ~n29263;
  assign n29265 = ~n29245 & n29264;
  assign n29266 = pi140 & ~n29265;
  assign n29267 = ~n29244 & n29266;
  assign n29268 = ~n29234 & ~n29267;
  assign n29269 = ~pi181 & ~n29268;
  assign n29270 = n29218 & n29227;
  assign n29271 = ~n29198 & ~n29270;
  assign n29272 = ~pi142 & ~n29271;
  assign n29273 = ~pi40 & n2680;
  assign n29274 = ~n29108 & ~n29180;
  assign n29275 = ~n29196 & n29274;
  assign n29276 = n29273 & n29275;
  assign n29277 = ~n29198 & ~n29276;
  assign n29278 = pi142 & ~n29277;
  assign n29279 = ~pi140 & ~n29278;
  assign n29280 = ~n29272 & n29279;
  assign n29281 = n2680 & ~n29108;
  assign n29282 = ~n29108 & n29241;
  assign n29283 = ~n29240 & n29281;
  assign n29284 = ~n29198 & ~n60124;
  assign n29285 = ~pi142 & ~n29284;
  assign n29286 = ~n29261 & n29281;
  assign n29287 = ~n29198 & ~n29286;
  assign n29288 = pi142 & ~n29287;
  assign n29289 = pi140 & ~n29288;
  assign n29290 = pi140 & ~n29285;
  assign n29291 = ~n29288 & n29290;
  assign n29292 = ~n29285 & n29289;
  assign n29293 = ~n29280 & ~n60125;
  assign n29294 = pi181 & ~n29293;
  assign n29295 = pi144 & ~n29294;
  assign n29296 = ~n29269 & n29295;
  assign n29297 = ~pi93 & ~n29253;
  assign n29298 = n29250 & ~n29297;
  assign n29299 = n29248 & ~n29298;
  assign n29300 = n29246 & ~n29299;
  assign n29301 = ~pi95 & ~n29300;
  assign n29302 = n29281 & ~n29301;
  assign n29303 = ~n29198 & ~n29302;
  assign n29304 = pi142 & ~n29303;
  assign n29305 = ~n29217 & ~n29245;
  assign n29306 = ~pi142 & n29305;
  assign n29307 = pi140 & ~n29306;
  assign n29308 = pi140 & ~n29304;
  assign n29309 = ~n29306 & n29308;
  assign n29310 = ~n29304 & n29307;
  assign n29311 = n2502 & n29128;
  assign n29312 = n2446 & ~n29311;
  assign n29313 = ~pi58 & ~n29312;
  assign n29314 = n2580 & n29313;
  assign n29315 = ~n29202 & ~n29314;
  assign n29316 = ~pi70 & ~n29315;
  assign n29317 = ~n29121 & ~n29316;
  assign n29318 = ~pi51 & ~n29317;
  assign n29319 = n29174 & ~n29318;
  assign n29320 = ~n29119 & ~n29319;
  assign n29321 = ~pi40 & n29320;
  assign n29322 = ~pi32 & ~n29321;
  assign n29323 = ~n29200 & ~n29322;
  assign n29324 = ~pi95 & ~n29323;
  assign n29325 = pi198 & n29324;
  assign n29326 = ~n29221 & ~n29322;
  assign n29327 = ~pi95 & ~n29326;
  assign n29328 = ~pi198 & n29327;
  assign n29329 = ~n29219 & ~n29328;
  assign n29330 = ~n29219 & ~n29324;
  assign n29331 = pi198 & ~n29330;
  assign n29332 = ~n29219 & ~n29327;
  assign n29333 = ~pi198 & ~n29332;
  assign n29334 = ~n29331 & ~n29333;
  assign n29335 = ~n29325 & n29329;
  assign n29336 = n29273 & ~n60127;
  assign n29337 = ~n29198 & ~n29336;
  assign n29338 = ~pi142 & ~n29337;
  assign n29339 = ~n29123 & ~n29313;
  assign n29340 = ~pi90 & ~n29339;
  assign n29341 = n29166 & ~n29340;
  assign n29342 = n29169 & ~n29341;
  assign n29343 = ~n29121 & ~n29342;
  assign n29344 = ~pi51 & ~n29343;
  assign n29345 = n29174 & ~n29344;
  assign n29346 = ~n29119 & ~n29345;
  assign n29347 = ~pi40 & ~n29346;
  assign n29348 = ~pi32 & ~n29347;
  assign n29349 = ~n29118 & ~n29348;
  assign n29350 = ~pi95 & ~n29349;
  assign n29351 = n29281 & ~n29350;
  assign n29352 = ~n29190 & ~n29348;
  assign n29353 = ~pi95 & ~n29352;
  assign n29354 = ~pi198 & n29353;
  assign n29355 = n29351 & ~n29354;
  assign n29356 = ~n29198 & ~n29355;
  assign n29357 = pi142 & ~n29356;
  assign n29358 = ~pi140 & ~n29357;
  assign n29359 = ~pi140 & ~n29338;
  assign n29360 = ~n29357 & n29359;
  assign n29361 = ~n29338 & n29358;
  assign n29362 = ~n60126 & ~n60128;
  assign n29363 = pi181 & ~n29362;
  assign n29364 = ~pi40 & ~n29320;
  assign n29365 = ~pi32 & ~n29364;
  assign n29366 = ~n29118 & ~n29365;
  assign n29367 = ~pi95 & ~n29366;
  assign n29368 = ~n29117 & ~n29367;
  assign n29369 = ~n29190 & ~n29365;
  assign n29370 = ~pi95 & ~n29369;
  assign n29371 = ~pi198 & n29370;
  assign n29372 = n29368 & ~n29371;
  assign n29373 = n2680 & ~n29372;
  assign n29374 = ~n29245 & ~n29373;
  assign n29375 = ~pi142 & n29374;
  assign n29376 = ~n29117 & ~n29350;
  assign n29377 = ~n29354 & n29376;
  assign n29378 = n2680 & ~n29377;
  assign n29379 = pi142 & ~n29378;
  assign n29380 = ~n29245 & n29379;
  assign n29381 = ~pi140 & ~n29380;
  assign n29382 = ~n29375 & n29381;
  assign n29383 = ~pi95 & ~n29065;
  assign n29384 = ~n29117 & ~n29383;
  assign n29385 = n2680 & n29384;
  assign n29386 = ~n29198 & ~n29385;
  assign n29387 = ~pi142 & ~n29386;
  assign n29388 = ~n29117 & ~n29301;
  assign n29389 = n2680 & ~n29388;
  assign n29390 = pi142 & ~n29389;
  assign n29391 = ~n29245 & n29390;
  assign n29392 = pi140 & ~n29391;
  assign n29393 = ~n29387 & n29392;
  assign n29394 = ~n29382 & ~n29393;
  assign n29395 = ~pi181 & ~n29394;
  assign n29396 = ~pi144 & ~n29395;
  assign n29397 = ~n29363 & n29396;
  assign n29398 = ~pi299 & ~n29397;
  assign n29399 = pi181 & ~n60128;
  assign n29400 = ~n60126 & n29399;
  assign n29401 = ~pi140 & n29377;
  assign n29402 = pi140 & n29388;
  assign n29403 = pi142 & ~n29402;
  assign n29404 = ~n29401 & n29403;
  assign n29405 = ~pi140 & n29372;
  assign n29406 = pi140 & n29384;
  assign n29407 = ~pi142 & ~n29406;
  assign n29408 = ~n29405 & n29407;
  assign n29409 = ~n29404 & ~n29408;
  assign n29410 = n2680 & ~n29409;
  assign n29411 = ~pi181 & ~n29245;
  assign n29412 = ~n29410 & n29411;
  assign n29413 = ~pi144 & ~n29412;
  assign n29414 = ~n29400 & n29413;
  assign n29415 = ~pi181 & ~n29267;
  assign n29416 = ~n29234 & n29415;
  assign n29417 = pi181 & ~n60125;
  assign n29418 = ~n29280 & n29417;
  assign n29419 = pi144 & ~n29418;
  assign n29420 = ~n29416 & n29419;
  assign n29421 = ~n29414 & ~n29420;
  assign n29422 = ~pi299 & ~n29421;
  assign n29423 = ~n29296 & n29398;
  assign n29424 = ~pi159 & pi299;
  assign n29425 = ~pi210 & n29192;
  assign n29426 = n29181 & ~n29425;
  assign n29427 = ~n2680 & n29426;
  assign n29428 = ~n29242 & ~n29427;
  assign n29429 = ~pi146 & ~n29428;
  assign n29430 = ~n2680 & ~n29426;
  assign n29431 = ~n29263 & ~n29430;
  assign n29432 = pi146 & n29431;
  assign n29433 = pi161 & ~n29432;
  assign n29434 = pi161 & ~n29429;
  assign n29435 = ~n29432 & n29434;
  assign n29436 = ~n29429 & n29433;
  assign n29437 = ~n29385 & ~n29427;
  assign n29438 = ~pi146 & ~n29437;
  assign n29439 = ~n29389 & ~n29430;
  assign n29440 = pi146 & n29439;
  assign n29441 = ~pi161 & ~n29440;
  assign n29442 = ~pi161 & ~n29438;
  assign n29443 = ~n29440 & n29442;
  assign n29444 = ~n29438 & n29441;
  assign n29445 = ~n60130 & ~n60131;
  assign n29446 = pi162 & ~n29445;
  assign n29447 = ~pi210 & ~n29225;
  assign n29448 = n2680 & ~n29447;
  assign n29449 = ~n29217 & ~n29448;
  assign n29450 = n29216 & ~n29449;
  assign n29451 = pi161 & ~n29450;
  assign n29452 = ~n29108 & ~n29370;
  assign n29453 = ~pi210 & ~n29452;
  assign n29454 = n2680 & ~n29453;
  assign n29455 = ~n29217 & ~n29454;
  assign n29456 = n29368 & ~n29455;
  assign n29457 = ~pi161 & ~n29456;
  assign n29458 = ~pi146 & ~n29457;
  assign n29459 = ~n29451 & n29458;
  assign n29460 = ~pi162 & ~n29427;
  assign n29461 = ~pi210 & n29353;
  assign n29462 = n29376 & ~n29461;
  assign n29463 = n2680 & n29462;
  assign n29464 = ~pi161 & ~n29463;
  assign n29465 = pi161 & ~n29426;
  assign n29466 = pi146 & ~n29465;
  assign n29467 = pi146 & ~n29464;
  assign n29468 = ~n29465 & n29467;
  assign n29469 = ~n29464 & n29466;
  assign n29470 = n29460 & ~n60132;
  assign n29471 = pi161 & n29426;
  assign n29472 = ~pi161 & n29463;
  assign n29473 = pi146 & ~n29472;
  assign n29474 = ~n29471 & n29473;
  assign n29475 = pi161 & n29450;
  assign n29476 = ~pi161 & n29456;
  assign n29477 = ~pi146 & ~n29476;
  assign n29478 = ~n29475 & n29477;
  assign n29479 = ~n29474 & ~n29478;
  assign n29480 = n29460 & ~n29479;
  assign n29481 = ~n29459 & n29470;
  assign n29482 = ~n29446 & ~n60133;
  assign n29483 = n29424 & ~n29482;
  assign n29484 = ~n29302 & ~n29427;
  assign n29485 = pi146 & ~n29484;
  assign n29486 = ~n29217 & ~n29430;
  assign n29487 = ~pi146 & n29486;
  assign n29488 = ~pi161 & ~n29487;
  assign n29489 = ~n29485 & n29488;
  assign n29490 = ~n29286 & ~n29427;
  assign n29491 = pi146 & ~n29490;
  assign n29492 = ~n60124 & ~n29427;
  assign n29493 = ~pi146 & ~n29492;
  assign n29494 = pi161 & ~n29493;
  assign n29495 = pi161 & ~n29491;
  assign n29496 = ~n29493 & n29495;
  assign n29497 = ~n29491 & n29494;
  assign n29498 = pi162 & ~n60134;
  assign n29499 = pi162 & ~n29489;
  assign n29500 = ~n60134 & n29499;
  assign n29501 = ~n29489 & n29498;
  assign n29502 = pi159 & pi299;
  assign n29503 = ~n29108 & ~n29367;
  assign n29504 = n29454 & n29503;
  assign n29505 = ~n29427 & ~n29504;
  assign n29506 = ~pi146 & ~n29505;
  assign n29507 = n29351 & ~n29461;
  assign n29508 = ~n29427 & ~n29507;
  assign n29509 = pi146 & ~n29508;
  assign n29510 = ~pi161 & ~n29509;
  assign n29511 = ~n29506 & n29510;
  assign n29512 = n29218 & n29448;
  assign n29513 = ~n29427 & ~n29512;
  assign n29514 = ~pi146 & ~n29513;
  assign n29515 = n29274 & ~n29425;
  assign n29516 = n2680 & ~n29515;
  assign n29517 = ~n29430 & ~n29516;
  assign n29518 = pi146 & n29517;
  assign n29519 = pi161 & ~n29518;
  assign n29520 = ~n29514 & n29519;
  assign n29521 = ~pi162 & ~n29520;
  assign n29522 = ~n29511 & n29521;
  assign n29523 = n29502 & ~n29522;
  assign n29524 = ~n60135 & n29502;
  assign n29525 = ~n29522 & n29524;
  assign n29526 = ~n60135 & n29523;
  assign n29527 = ~n29483 & ~n60136;
  assign n29528 = ~n60129 & n29527;
  assign n29529 = pi232 & ~n29528;
  assign n29530 = ~n29195 & ~n29529;
  assign n29531 = n2634 & ~n29530;
  assign n29532 = pi216 & n2852;
  assign n29533 = ~pi95 & n29114;
  assign n29534 = n58838 & n6471;
  assign n29535 = pi1092 & n6471;
  assign n29536 = n2862 & ~n28505;
  assign n29537 = n29535 & n29536;
  assign n29538 = ~n29534 & ~n29537;
  assign n29539 = n29533 & ~n29538;
  assign n29540 = n2783 & n29539;
  assign n29541 = n29065 & ~n29540;
  assign n29542 = n2680 & n29539;
  assign n29543 = n29065 & ~n29542;
  assign n29544 = ~n58846 & ~n29543;
  assign n29545 = n29541 & ~n29544;
  assign n29546 = n29533 & n29534;
  assign n29547 = ~n2822 & n29546;
  assign n29548 = n29065 & ~n29547;
  assign n29549 = n2680 & n29548;
  assign n29550 = ~pi161 & n29549;
  assign n29551 = ~n29545 & ~n29550;
  assign n29552 = n29532 & ~n29551;
  assign n29553 = n29065 & ~n29532;
  assign n29554 = pi299 & ~n29553;
  assign n29555 = ~pi38 & ~pi155;
  assign n29556 = n29554 & n29555;
  assign n29557 = ~n29552 & n29556;
  assign n29558 = n29533 & n29537;
  assign n29559 = n29065 & ~n29558;
  assign n29560 = n2844 & ~n29559;
  assign n29561 = pi161 & n29560;
  assign n29562 = n29532 & n29541;
  assign n29563 = ~n29561 & n29562;
  assign n29564 = ~pi38 & pi155;
  assign n29565 = n29554 & n29564;
  assign n29566 = ~n29563 & n29565;
  assign n29567 = ~n29552 & n29555;
  assign n29568 = ~n29563 & n29564;
  assign n29569 = ~n29567 & ~n29568;
  assign n29570 = n29554 & ~n29569;
  assign n29571 = ~n29557 & ~n29566;
  assign n29572 = pi224 & n2829;
  assign n29573 = n29065 & ~n29572;
  assign n29574 = ~n2790 & ~n29543;
  assign n29575 = n29541 & ~n29574;
  assign n29576 = ~n29541 & ~n29573;
  assign n29577 = ~n29573 & n29574;
  assign n29578 = ~n29576 & ~n29577;
  assign n29579 = ~n29573 & ~n29575;
  assign n29580 = pi144 & n60138;
  assign n29581 = ~pi177 & ~pi299;
  assign n29582 = n2791 & n29546;
  assign n29583 = n29065 & n29572;
  assign n29584 = ~n29582 & n29583;
  assign n29585 = ~n29573 & ~n29584;
  assign n29586 = ~pi144 & ~n29576;
  assign n29587 = ~n29585 & n29586;
  assign n29588 = n29581 & ~n29587;
  assign n29589 = ~n29580 & n29588;
  assign n29590 = n2680 & n29572;
  assign n29591 = n29558 & n29590;
  assign n29592 = n29065 & ~n29591;
  assign n29593 = n2680 & n29558;
  assign n29594 = n29065 & ~n29593;
  assign n29595 = ~n2790 & ~n29594;
  assign n29596 = ~n29573 & n29595;
  assign n29597 = ~n2790 & ~n29592;
  assign n29598 = ~n29576 & ~n60139;
  assign n29599 = ~pi299 & ~n29598;
  assign n29600 = pi177 & ~n29586;
  assign n29601 = pi177 & ~pi299;
  assign n29602 = ~n29586 & n29601;
  assign n29603 = ~n29598 & n29602;
  assign n29604 = n29599 & n29600;
  assign n29605 = ~n29589 & ~n60140;
  assign n29606 = ~pi38 & ~n29605;
  assign n29607 = ~n60137 & ~n29606;
  assign n29608 = pi232 & ~n29607;
  assign n29609 = ~n29545 & n29554;
  assign n29610 = ~pi299 & ~n60138;
  assign n29611 = ~n29609 & ~n29610;
  assign n29612 = ~pi232 & ~n29611;
  assign n29613 = ~pi38 & n29612;
  assign n29614 = pi232 & ~n29605;
  assign n29615 = ~n29612 & ~n29614;
  assign n29616 = ~pi38 & ~n29615;
  assign n29617 = pi232 & n29554;
  assign n29618 = pi232 & n60137;
  assign n29619 = ~n29569 & n29617;
  assign n29620 = ~n29616 & ~n60141;
  assign n29621 = ~n29608 & ~n29613;
  assign n29622 = pi39 & ~n60142;
  assign n29623 = ~pi299 & n2681;
  assign n29624 = ~n59171 & n29623;
  assign n29625 = ~pi167 & ~n29624;
  assign n29626 = n2681 & ~n59171;
  assign n29627 = pi167 & ~n29626;
  assign n29628 = pi188 & ~n29627;
  assign n29629 = ~n29625 & n29628;
  assign n29630 = pi299 & ~n59171;
  assign n29631 = ~pi188 & n29046;
  assign n29632 = n29630 & n29631;
  assign n29633 = pi38 & ~n29632;
  assign n29634 = pi188 & n29624;
  assign n29635 = ~pi167 & ~n29634;
  assign n29636 = pi167 & pi188;
  assign n29637 = ~n29626 & n29636;
  assign n29638 = pi299 & n2681;
  assign n29639 = n2681 & n29630;
  assign n29640 = ~n59171 & n29638;
  assign n29641 = ~pi188 & ~n60143;
  assign n29642 = ~n29637 & ~n29641;
  assign n29643 = pi188 & ~n29625;
  assign n29644 = pi167 & n60143;
  assign n29645 = ~n29643 & ~n29644;
  assign n29646 = ~n29637 & ~n29645;
  assign n29647 = ~n29635 & n29642;
  assign n29648 = pi38 & ~n60144;
  assign n29649 = ~n29629 & n29633;
  assign n29650 = ~pi87 & ~n60145;
  assign n29651 = ~n29622 & n29650;
  assign n29652 = ~n29531 & n29651;
  assign n29653 = ~pi38 & ~n29065;
  assign n29654 = pi38 & ~n29103;
  assign n29655 = ~n29653 & ~n29654;
  assign n29656 = pi87 & n29655;
  assign n29657 = ~pi100 & ~n29656;
  assign n29658 = ~n29652 & n29657;
  assign n29659 = ~n29086 & ~n29658;
  assign n29660 = n6307 & ~n29659;
  assign n29661 = ~pi75 & pi92;
  assign n29662 = ~pi87 & n6860;
  assign n29663 = n2671 & n29533;
  assign n29664 = n29114 & n29662;
  assign n29665 = ~pi155 & pi299;
  assign n29666 = pi155 & pi299;
  assign n29667 = ~n29601 & ~n29666;
  assign n29668 = ~n29581 & ~n29665;
  assign n29669 = ~pi38 & n60147;
  assign n29670 = n2681 & ~n29669;
  assign n29671 = n60146 & ~n29670;
  assign n29672 = n29655 & ~n29671;
  assign n29673 = ~pi100 & ~n29672;
  assign n29674 = ~n29086 & ~n29673;
  assign n29675 = n29661 & ~n29674;
  assign n29676 = ~n29087 & ~n29675;
  assign n29677 = ~n29660 & n29676;
  assign n29678 = ~pi54 & ~n29677;
  assign n29679 = ~n29107 & ~n29678;
  assign n29680 = ~pi74 & ~n29679;
  assign n29681 = n29096 & ~n29680;
  assign n29682 = pi55 & ~n29053;
  assign n29683 = pi54 & n29049;
  assign n29684 = n29060 & ~n29067;
  assign n29685 = ~n2438 & ~n29684;
  assign n29686 = ~n2635 & n29040;
  assign n29687 = n29031 & n29067;
  assign n29688 = ~n29686 & ~n29687;
  assign n29689 = pi232 & ~n29688;
  assign n29690 = n29066 & ~n60146;
  assign n29691 = ~n29057 & ~n29690;
  assign n29692 = n2635 & ~n29691;
  assign n29693 = ~n29689 & ~n29692;
  assign n29694 = pi100 & ~n29042;
  assign n29695 = ~n29031 & n60146;
  assign n29696 = n29066 & ~n29695;
  assign n29697 = ~pi100 & ~n29696;
  assign n29698 = ~pi232 & n60146;
  assign n29699 = ~n29697 & ~n29698;
  assign n29700 = ~n29057 & ~n29699;
  assign n29701 = ~n29694 & ~n29700;
  assign n29702 = ~pi75 & ~n29701;
  assign n29703 = pi75 & ~n29042;
  assign n29704 = ~pi92 & ~n29703;
  assign n29705 = ~n29702 & n29704;
  assign n29706 = ~pi92 & ~n29693;
  assign n29707 = ~n29685 & ~n60148;
  assign n29708 = ~n29683 & ~n29707;
  assign n29709 = ~pi74 & ~n29708;
  assign n29710 = n29682 & ~n29709;
  assign n29711 = n4437 & ~n29710;
  assign n29712 = ~n29681 & n29711;
  assign n29713 = ~n29071 & ~n29712;
  assign n29714 = ~n29055 & ~n29713;
  assign n29715 = ~pi34 & n29714;
  assign n29716 = pi159 & n28314;
  assign n29717 = n2599 & n28321;
  assign n29718 = pi90 & ~n2554;
  assign n29719 = pi58 & n58795;
  assign n29720 = ~pi90 & ~n29719;
  assign n29721 = n2592 & ~n29720;
  assign n29722 = ~n29718 & ~n29720;
  assign n29723 = n2592 & n29722;
  assign n29724 = ~n29718 & n29721;
  assign n29725 = n2501 & ~n28333;
  assign n29726 = n2577 & n2592;
  assign n29727 = n29725 & n29726;
  assign n29728 = n2446 & n29727;
  assign n29729 = n29154 & n29728;
  assign n29730 = ~pi70 & ~n29729;
  assign n29731 = ~n60149 & n29730;
  assign n29732 = n29717 & ~n29731;
  assign n29733 = ~pi146 & n29732;
  assign n29734 = n29717 & ~n29730;
  assign n29735 = ~n28474 & ~n29734;
  assign n29736 = ~pi161 & n29735;
  assign n29737 = ~n29733 & n29736;
  assign n29738 = ~n29127 & n29727;
  assign n29739 = ~pi70 & ~n29738;
  assign n29740 = ~n60149 & n29739;
  assign n29741 = n29717 & ~n29740;
  assign n29742 = ~pi146 & n29741;
  assign n29743 = n29717 & ~n29739;
  assign n29744 = ~n28474 & ~n29743;
  assign n29745 = pi161 & n29744;
  assign n29746 = ~n29742 & n29745;
  assign n29747 = pi162 & ~n29746;
  assign n29748 = ~n29737 & n29747;
  assign n29749 = ~n29716 & ~n29748;
  assign n29750 = n2680 & ~n29749;
  assign n29751 = n2446 & n29254;
  assign n29752 = n29720 & ~n29751;
  assign n29753 = n59137 & ~n29718;
  assign n29754 = ~n29752 & n29753;
  assign n29755 = n2598 & n2680;
  assign n29756 = ~pi40 & n29755;
  assign n29757 = n29754 & n29756;
  assign n29758 = ~pi146 & ~n29757;
  assign n29759 = n59138 & n29751;
  assign n29760 = n2598 & n29759;
  assign n29761 = n29273 & n29760;
  assign n29762 = pi146 & ~n29761;
  assign n29763 = ~pi161 & ~n29762;
  assign n29764 = ~n29758 & n29763;
  assign n29765 = n59137 & n29722;
  assign n29766 = ~n29720 & n29753;
  assign n29767 = n29756 & n60150;
  assign n29768 = ~pi146 & pi161;
  assign n29769 = n29767 & n29768;
  assign n29770 = ~n29764 & ~n29769;
  assign n29771 = ~pi162 & ~n29770;
  assign n29772 = pi299 & ~n29771;
  assign n29773 = ~n29733 & n29735;
  assign n29774 = ~pi161 & ~n29773;
  assign n29775 = ~n29742 & n29744;
  assign n29776 = pi161 & ~n29775;
  assign n29777 = pi299 & ~n29716;
  assign n29778 = ~n29776 & n29777;
  assign n29779 = ~n29774 & n29778;
  assign n29780 = ~pi162 & ~n29716;
  assign n29781 = n2680 & ~n29780;
  assign n29782 = n2680 & n28314;
  assign n29783 = ~pi162 & n29782;
  assign n29784 = n29502 & ~n29783;
  assign n29785 = ~n29424 & ~n29784;
  assign n29786 = ~n29031 & ~n29785;
  assign n29787 = pi299 & ~n29781;
  assign n29788 = ~n29779 & ~n60151;
  assign n29789 = ~n29771 & ~n29788;
  assign n29790 = ~n29750 & n29772;
  assign n29791 = ~pi142 & n29732;
  assign n29792 = ~n28443 & ~n29734;
  assign n29793 = ~pi144 & n29792;
  assign n29794 = ~n29791 & n29793;
  assign n29795 = ~pi142 & n29741;
  assign n29796 = ~n28443 & ~n29743;
  assign n29797 = pi144 & n29796;
  assign n29798 = ~n29795 & n29797;
  assign n29799 = pi140 & n2680;
  assign n29800 = ~n29798 & n29799;
  assign n29801 = ~n29794 & n29800;
  assign n29802 = ~pi142 & ~n29757;
  assign n29803 = pi142 & ~n29761;
  assign n29804 = ~pi144 & ~n29803;
  assign n29805 = ~n29802 & n29804;
  assign n29806 = ~pi142 & pi144;
  assign n29807 = n29767 & n29806;
  assign n29808 = ~n29805 & ~n29807;
  assign n29809 = ~pi140 & ~n29808;
  assign n29810 = pi181 & n29782;
  assign n29811 = ~pi299 & ~n29810;
  assign n29812 = ~n29809 & n29811;
  assign n29813 = ~pi142 & n29757;
  assign n29814 = pi142 & n29761;
  assign n29815 = ~pi140 & ~n29814;
  assign n29816 = ~n29813 & n29815;
  assign n29817 = pi140 & n29792;
  assign n29818 = ~n29791 & n29817;
  assign n29819 = ~n29816 & ~n29818;
  assign n29820 = ~pi144 & ~n29819;
  assign n29821 = ~n29795 & n29796;
  assign n29822 = pi140 & ~n29821;
  assign n29823 = pi144 & ~n29822;
  assign n29824 = ~pi142 & n29767;
  assign n29825 = ~pi140 & ~n29824;
  assign n29826 = pi140 & ~n29795;
  assign n29827 = n29796 & n29826;
  assign n29828 = ~n29825 & ~n29827;
  assign n29829 = pi144 & ~n29828;
  assign n29830 = n29823 & ~n29824;
  assign n29831 = pi140 & ~n2680;
  assign n29832 = n2680 & ~n29823;
  assign n29833 = pi140 & ~n29832;
  assign n29834 = ~n60153 & ~n29833;
  assign n29835 = ~n60153 & ~n29831;
  assign n29836 = ~n29820 & n60154;
  assign n29837 = n29811 & ~n29836;
  assign n29838 = ~n29801 & n29812;
  assign n29839 = pi232 & ~n60155;
  assign n29840 = pi232 & ~n60152;
  assign n29841 = ~n60155 & n29840;
  assign n29842 = ~n60152 & n29839;
  assign n29843 = n2634 & ~n60156;
  assign n29844 = n2844 & ~n28517;
  assign n29845 = ~pi161 & ~n29844;
  assign n29846 = n2680 & n58842;
  assign n29847 = ~n58846 & n29846;
  assign n29848 = n58842 & n2844;
  assign n29849 = pi161 & ~n60157;
  assign n29850 = n29532 & ~n29849;
  assign n29851 = n29532 & ~n29845;
  assign n29852 = ~n29849 & n29851;
  assign n29853 = ~n29845 & n29850;
  assign n29854 = n29564 & ~n60158;
  assign n29855 = n2844 & n28507;
  assign n29856 = ~pi161 & n29532;
  assign n29857 = n29855 & n29856;
  assign n29858 = n29555 & ~n29857;
  assign n29859 = ~n29854 & ~n29858;
  assign n29860 = pi299 & ~n29859;
  assign n29861 = ~n2790 & n29572;
  assign n29862 = n2680 & n29861;
  assign n29863 = n2791 & n29572;
  assign n29864 = ~n28517 & n29572;
  assign n29865 = n2791 & n29864;
  assign n29866 = ~n28517 & n60159;
  assign n29867 = ~pi144 & n60160;
  assign n29868 = n58842 & n60159;
  assign n29869 = pi144 & n29868;
  assign n29870 = n29601 & ~n29869;
  assign n29871 = n29601 & ~n29867;
  assign n29872 = ~n29869 & n29871;
  assign n29873 = ~n29867 & n29870;
  assign n29874 = n2791 & n28507;
  assign n29875 = n29572 & n29874;
  assign n29876 = n28507 & n60159;
  assign n29877 = ~pi144 & n60162;
  assign n29878 = n29581 & ~n29877;
  assign n29879 = pi232 & ~n29878;
  assign n29880 = ~n60161 & n29879;
  assign n29881 = ~pi38 & ~n29880;
  assign n29882 = ~n29860 & ~n29881;
  assign n29883 = pi39 & ~n29882;
  assign n29884 = ~n60145 & ~n29883;
  assign n29885 = ~n29843 & n29884;
  assign n29886 = ~pi100 & ~n29885;
  assign n29887 = ~n29086 & ~n29886;
  assign n29888 = ~pi87 & ~n29887;
  assign n29889 = ~n2636 & ~n29104;
  assign n29890 = ~n29086 & n29889;
  assign n29891 = pi87 & ~n29890;
  assign n29892 = ~n29888 & ~n29891;
  assign n29893 = n6307 & ~n29892;
  assign n29894 = pi38 & ~n60117;
  assign n29895 = n2634 & ~n60147;
  assign n29896 = n28575 & ~n60147;
  assign n29897 = n58822 & n29895;
  assign n29898 = ~n29894 & ~n60163;
  assign n29899 = n2681 & ~n29898;
  assign n29900 = ~pi100 & ~n29899;
  assign n29901 = ~n29086 & ~n29900;
  assign n29902 = ~pi87 & ~n29901;
  assign n29903 = ~n29891 & ~n29902;
  assign n29904 = n29661 & ~n29903;
  assign n29905 = ~n29087 & ~n29904;
  assign n29906 = ~n29893 & n29905;
  assign n29907 = ~pi54 & ~n29906;
  assign n29908 = ~n29107 & ~n29907;
  assign n29909 = ~pi74 & ~n29908;
  assign n29910 = n29096 & ~n29909;
  assign n29911 = n58822 & n2680;
  assign n29912 = ~pi39 & pi232;
  assign n29913 = ~pi92 & pi162;
  assign n29914 = n29912 & n29913;
  assign n29915 = n9186 & n29913;
  assign n29916 = n29912 & n29915;
  assign n29917 = n9186 & n29914;
  assign n29918 = n29911 & n60164;
  assign n29919 = ~n29057 & ~n29918;
  assign n29920 = n2635 & ~n29919;
  assign n29921 = n29056 & ~n29920;
  assign n29922 = ~n29683 & ~n29921;
  assign n29923 = ~pi74 & ~n29922;
  assign n29924 = n29682 & ~n29923;
  assign n29925 = n4437 & ~n29924;
  assign n29926 = ~n29910 & n29925;
  assign n29927 = n29064 & ~n29926;
  assign n29928 = ~n29055 & ~n29927;
  assign n29929 = pi34 & n29928;
  assign n29930 = ~pi33 & ~pi954;
  assign n29931 = ~n29929 & ~n29930;
  assign n29932 = ~n29715 & n29931;
  assign n29933 = ~pi195 & ~pi196;
  assign n29934 = ~pi138 & n29933;
  assign n29935 = ~pi139 & n29934;
  assign n29936 = ~pi118 & n29935;
  assign n29937 = ~pi79 & n29936;
  assign n29938 = ~pi34 & ~n29937;
  assign n29939 = n29714 & ~n29938;
  assign n29940 = n29928 & n29938;
  assign n29941 = n29930 & ~n29940;
  assign n29942 = ~n29939 & n29941;
  assign po192 = ~n29932 & ~n29942;
  assign n29944 = pi163 & ~n29038;
  assign n29945 = ~pi163 & ~n29033;
  assign n29946 = ~n29036 & n29945;
  assign n29947 = ~n29944 & ~n29946;
  assign n29948 = pi232 & n29947;
  assign n29949 = pi75 & ~n29948;
  assign n29950 = pi100 & ~n29948;
  assign n29951 = ~n29949 & ~n29950;
  assign n29952 = pi147 & n2681;
  assign n29953 = n2635 & n29952;
  assign n29954 = n29951 & ~n29953;
  assign n29955 = ~n2635 & n29948;
  assign n29956 = pi74 & ~n29955;
  assign n29957 = ~n4438 & ~n29956;
  assign n29958 = n29954 & n29957;
  assign n29959 = pi299 & ~n29947;
  assign n29960 = ~n29079 & n29080;
  assign n29961 = pi184 & n2680;
  assign n29962 = ~n29960 & n29961;
  assign n29963 = ~pi184 & n29960;
  assign n29964 = ~pi299 & ~n29963;
  assign n29965 = ~n29962 & n29964;
  assign n29966 = pi232 & ~n29965;
  assign n29967 = ~n29959 & n29966;
  assign n29968 = ~n2635 & n29967;
  assign n29969 = pi74 & ~n29968;
  assign n29970 = ~pi55 & ~n29969;
  assign n29971 = ~pi187 & ~pi299;
  assign n29972 = ~pi147 & pi299;
  assign n29973 = ~n29971 & ~n29972;
  assign n29974 = n2681 & n29973;
  assign n29975 = n2635 & ~n29974;
  assign n29976 = pi54 & ~n29975;
  assign n29977 = ~n29968 & n29976;
  assign n29978 = ~pi187 & ~n60143;
  assign n29979 = pi187 & ~n29626;
  assign n29980 = pi147 & ~n29979;
  assign n29981 = ~n29978 & n29980;
  assign n29982 = ~pi147 & pi187;
  assign n29983 = n29624 & n29982;
  assign n29984 = ~n29981 & ~n29983;
  assign n29985 = pi38 & ~n29984;
  assign n29986 = ~pi40 & ~n29300;
  assign n29987 = ~pi95 & ~n29986;
  assign n29988 = ~pi40 & ~n29260;
  assign n29989 = pi166 & n29988;
  assign n29990 = n29987 & ~n29989;
  assign n29991 = n2680 & ~n29219;
  assign n29992 = ~n29990 & n29991;
  assign n29993 = ~pi153 & ~n29992;
  assign n29994 = ~pi40 & ~n29239;
  assign n29995 = ~pi95 & ~n29994;
  assign n29996 = pi166 & ~n29995;
  assign n29997 = n29991 & n29996;
  assign n29998 = ~pi166 & n2680;
  assign n29999 = n29199 & n29998;
  assign n30000 = pi153 & ~n29999;
  assign n30001 = ~n29997 & n30000;
  assign n30002 = pi160 & ~n30001;
  assign n30003 = ~n29993 & n30002;
  assign n30004 = ~pi153 & n29990;
  assign n30005 = ~n28313 & ~n29219;
  assign n30006 = n29110 & ~n29115;
  assign n30007 = ~n30005 & ~n30006;
  assign n30008 = n2579 & n2621;
  assign n30009 = n58823 & n30008;
  assign n30010 = n2621 & n59138;
  assign n30011 = n2599 & n60073;
  assign n30012 = n2621 & n29759;
  assign n30013 = n29751 & n60165;
  assign n30014 = ~n29995 & ~n60166;
  assign n30015 = pi153 & ~n29996;
  assign n30016 = ~n30014 & n30015;
  assign n30017 = ~pi160 & n2680;
  assign n30018 = ~n30016 & n30017;
  assign n30019 = ~n30007 & n30018;
  assign n30020 = ~n30004 & n30019;
  assign n30021 = pi163 & ~n30020;
  assign n30022 = ~n30003 & n30021;
  assign n30023 = ~pi40 & ~n29515;
  assign n30024 = ~pi95 & ~n30023;
  assign n30025 = ~n30007 & ~n30024;
  assign n30026 = pi166 & n30025;
  assign n30027 = ~pi40 & n29346;
  assign n30028 = ~pi32 & ~n30027;
  assign n30029 = ~n29200 & ~n30028;
  assign n30030 = ~pi95 & ~n30029;
  assign n30031 = ~n30007 & ~n30030;
  assign n30032 = pi210 & ~n30031;
  assign n30033 = ~n29221 & ~n30028;
  assign n30034 = ~pi95 & ~n30033;
  assign n30035 = ~n30007 & ~n30034;
  assign n30036 = ~pi210 & ~n30035;
  assign n30037 = n29998 & ~n30036;
  assign n30038 = n29998 & ~n30032;
  assign n30039 = ~n30036 & n30038;
  assign n30040 = ~n30032 & n30037;
  assign n30041 = ~pi153 & ~n60167;
  assign n30042 = ~n30026 & n30041;
  assign n30043 = pi210 & n29324;
  assign n30044 = ~pi210 & n29327;
  assign n30045 = n29998 & ~n30044;
  assign n30046 = ~n30043 & n30045;
  assign n30047 = ~pi95 & ~n29212;
  assign n30048 = pi210 & n30047;
  assign n30049 = pi166 & n2680;
  assign n30050 = ~pi210 & n29223;
  assign n30051 = n30049 & ~n30050;
  assign n30052 = ~n30048 & n30051;
  assign n30053 = ~n30046 & ~n30052;
  assign n30054 = ~n30007 & ~n30053;
  assign n30055 = ~n29324 & ~n30007;
  assign n30056 = pi210 & ~n30055;
  assign n30057 = ~n29327 & ~n30007;
  assign n30058 = ~pi210 & ~n30057;
  assign n30059 = n29998 & ~n30058;
  assign n30060 = ~n30056 & n30059;
  assign n30061 = ~n29223 & ~n30007;
  assign n30062 = ~pi210 & ~n30061;
  assign n30063 = ~n30007 & ~n30047;
  assign n30064 = pi210 & ~n30063;
  assign n30065 = n30049 & ~n30064;
  assign n30066 = ~n30062 & n30065;
  assign n30067 = pi153 & ~n30066;
  assign n30068 = ~n30060 & n30067;
  assign n30069 = pi153 & ~n30060;
  assign n30070 = ~n30066 & n30069;
  assign n30071 = pi153 & ~n30054;
  assign n30072 = ~pi160 & ~n60168;
  assign n30073 = ~n30042 & n30072;
  assign n30074 = n30023 & n30049;
  assign n30075 = ~n29219 & ~n30034;
  assign n30076 = ~pi210 & ~n30075;
  assign n30077 = ~n29219 & ~n30030;
  assign n30078 = pi210 & ~n30077;
  assign n30079 = n29998 & ~n30078;
  assign n30080 = n29998 & ~n30076;
  assign n30081 = ~n30078 & n30080;
  assign n30082 = ~n30076 & n30079;
  assign n30083 = ~pi153 & ~n60169;
  assign n30084 = ~n30074 & n30083;
  assign n30085 = ~n29219 & ~n30053;
  assign n30086 = ~n29219 & ~n30047;
  assign n30087 = pi210 & ~n30086;
  assign n30088 = ~pi210 & ~n29224;
  assign n30089 = n30049 & ~n30088;
  assign n30090 = ~n30087 & n30089;
  assign n30091 = pi210 & ~n29330;
  assign n30092 = ~pi210 & ~n29332;
  assign n30093 = n29998 & ~n30092;
  assign n30094 = n29998 & ~n30091;
  assign n30095 = ~n30092 & n30094;
  assign n30096 = ~n30091 & n30093;
  assign n30097 = pi153 & ~n60170;
  assign n30098 = ~n30090 & n30097;
  assign n30099 = pi153 & ~n30090;
  assign n30100 = ~n60170 & n30099;
  assign n30101 = pi153 & ~n30085;
  assign n30102 = pi160 & ~n60171;
  assign n30103 = ~n30084 & n30102;
  assign n30104 = ~pi163 & ~n30103;
  assign n30105 = ~n30073 & n30104;
  assign n30106 = ~n30022 & ~n30105;
  assign n30107 = ~n2680 & n30025;
  assign n30108 = pi299 & ~n30107;
  assign n30109 = ~n30106 & n30108;
  assign n30110 = ~pi40 & ~n29275;
  assign n30111 = ~pi95 & ~n30110;
  assign n30112 = ~n30007 & ~n30111;
  assign n30113 = ~n2680 & n30112;
  assign n30114 = ~pi175 & ~pi299;
  assign n30115 = pi189 & n29988;
  assign n30116 = n29987 & ~n30115;
  assign n30117 = ~pi182 & n30007;
  assign n30118 = pi182 & n29219;
  assign n30119 = n2680 & ~n30118;
  assign n30120 = n2680 & ~n30117;
  assign n30121 = ~n30118 & n30120;
  assign n30122 = ~n30117 & n30119;
  assign n30123 = ~n30116 & n60172;
  assign n30124 = pi184 & ~n30123;
  assign n30125 = pi189 & n2680;
  assign n30126 = n30110 & n30125;
  assign n30127 = pi198 & ~n30077;
  assign n30128 = ~pi189 & n2680;
  assign n30129 = ~pi198 & ~n30075;
  assign n30130 = n30128 & ~n30129;
  assign n30131 = ~n30127 & n30128;
  assign n30132 = ~n30129 & n30131;
  assign n30133 = ~n30127 & n30130;
  assign n30134 = pi182 & ~pi184;
  assign n30135 = ~n60173 & n30134;
  assign n30136 = ~n30126 & n30135;
  assign n30137 = ~n30124 & ~n30136;
  assign n30138 = n30114 & ~n30137;
  assign n30139 = pi198 & ~n30047;
  assign n30140 = ~pi198 & ~n29223;
  assign n30141 = ~n30139 & ~n30140;
  assign n30142 = pi189 & n60172;
  assign n30143 = ~n30141 & n30142;
  assign n30144 = pi95 & ~pi182;
  assign n30145 = ~n60127 & ~n30144;
  assign n30146 = ~pi189 & n30120;
  assign n30147 = ~n30007 & n30128;
  assign n30148 = ~n30145 & n30147;
  assign n30149 = ~n30145 & n30146;
  assign n30150 = n60127 & n30128;
  assign n30151 = pi198 & ~n30086;
  assign n30152 = ~pi198 & ~n29224;
  assign n30153 = n30125 & ~n30152;
  assign n30154 = ~n30151 & n30153;
  assign n30155 = pi182 & ~n30154;
  assign n30156 = pi182 & ~n30150;
  assign n30157 = ~n30154 & n30156;
  assign n30158 = ~n30150 & n30155;
  assign n30159 = pi198 & ~n30063;
  assign n30160 = ~pi198 & ~n30061;
  assign n30161 = n30125 & ~n30160;
  assign n30162 = ~n30159 & n30161;
  assign n30163 = ~pi182 & ~n30162;
  assign n30164 = ~n60175 & ~n30163;
  assign n30165 = ~n60174 & ~n30164;
  assign n30166 = ~n30143 & ~n60174;
  assign n30167 = ~pi184 & ~n60176;
  assign n30168 = pi175 & ~pi299;
  assign n30169 = ~pi95 & pi189;
  assign n30170 = n2446 & ~n30169;
  assign n30171 = n29994 & ~n30170;
  assign n30172 = ~n30144 & ~n30171;
  assign n30173 = n29961 & ~n30172;
  assign n30174 = ~n30117 & n30173;
  assign n30175 = n30168 & ~n30174;
  assign n30176 = ~n30167 & n30175;
  assign n30177 = ~n30138 & ~n30176;
  assign n30178 = ~n30113 & ~n30177;
  assign n30179 = n30112 & ~n30128;
  assign n30180 = pi198 & ~n30031;
  assign n30181 = ~pi198 & ~n30035;
  assign n30182 = n30128 & ~n30181;
  assign n30183 = n30128 & ~n30180;
  assign n30184 = ~n30181 & n30183;
  assign n30185 = ~n30180 & n30182;
  assign n30186 = ~pi182 & ~pi184;
  assign n30187 = n30114 & n30186;
  assign n30188 = ~n60177 & n30187;
  assign n30189 = ~n30179 & n30188;
  assign n30190 = ~n30178 & ~n30189;
  assign n30191 = ~n30109 & n30190;
  assign n30192 = pi232 & ~n30191;
  assign n30193 = pi299 & n30025;
  assign n30194 = ~pi299 & n30112;
  assign n30195 = ~pi232 & ~n30194;
  assign n30196 = ~n30193 & n30195;
  assign n30197 = ~pi39 & ~n30196;
  assign n30198 = ~n30192 & n30197;
  assign n30199 = ~n29199 & ~n29572;
  assign n30200 = ~pi40 & ~n29541;
  assign n30201 = ~pi189 & ~n30200;
  assign n30202 = n2446 & ~n29558;
  assign n30203 = n29273 & ~n30202;
  assign n30204 = n2822 & n29199;
  assign n30205 = n2446 & ~n29539;
  assign n30206 = ~pi40 & ~n30205;
  assign n30207 = n2783 & n30206;
  assign n30208 = ~n30204 & ~n30207;
  assign n30209 = ~n30203 & n30208;
  assign n30210 = pi189 & ~n2790;
  assign n30211 = n30209 & n30210;
  assign n30212 = ~n30201 & ~n30211;
  assign n30213 = pi179 & ~n30212;
  assign n30214 = n2790 & ~n30200;
  assign n30215 = n2446 & ~n29546;
  assign n30216 = n29273 & n29546;
  assign n30217 = ~n2446 & n29273;
  assign n30218 = ~n30216 & ~n30217;
  assign n30219 = n29273 & ~n30215;
  assign n30220 = n30208 & n60178;
  assign n30221 = ~pi189 & ~n30220;
  assign n30222 = ~n2822 & n30206;
  assign n30223 = ~n30204 & ~n30222;
  assign n30224 = pi189 & ~n30223;
  assign n30225 = ~pi179 & ~n2790;
  assign n30226 = ~n30224 & n30225;
  assign n30227 = ~n30221 & n30226;
  assign n30228 = ~n30214 & ~n30227;
  assign n30229 = ~n30213 & n30228;
  assign n30230 = n29572 & ~n30229;
  assign n30231 = ~n30199 & ~n30230;
  assign n30232 = ~pi299 & ~n30231;
  assign n30233 = n29199 & ~n29532;
  assign n30234 = pi299 & ~n30233;
  assign n30235 = ~n58846 & ~n30223;
  assign n30236 = n58846 & n30200;
  assign n30237 = n58846 & ~n30200;
  assign n30238 = ~n58846 & n30223;
  assign n30239 = ~n30237 & ~n30238;
  assign n30240 = ~n30235 & ~n30236;
  assign n30241 = ~pi166 & ~n58846;
  assign n30242 = ~n60179 & ~n30241;
  assign n30243 = n30220 & n30241;
  assign n30244 = n29532 & ~n30243;
  assign n30245 = ~n30242 & n30244;
  assign n30246 = n30234 & ~n30245;
  assign n30247 = ~n30232 & ~n30246;
  assign n30248 = ~pi156 & pi232;
  assign n30249 = ~n30247 & n30248;
  assign n30250 = pi166 & ~n58846;
  assign n30251 = n30209 & n30250;
  assign n30252 = ~n30200 & ~n30250;
  assign n30253 = n29532 & ~n30252;
  assign n30254 = ~n30251 & n30253;
  assign n30255 = n30234 & ~n30254;
  assign n30256 = ~n30232 & ~n30255;
  assign n30257 = pi156 & pi232;
  assign n30258 = ~n30256 & n30257;
  assign n30259 = ~n2790 & n30223;
  assign n30260 = ~n30214 & ~n30259;
  assign n30261 = n29572 & ~n30260;
  assign n30262 = ~pi299 & ~n30199;
  assign n30263 = ~n30261 & n30262;
  assign n30264 = n29554 & n60179;
  assign n30265 = ~pi232 & ~n30264;
  assign n30266 = ~n30263 & n30265;
  assign n30267 = pi39 & ~n30266;
  assign n30268 = ~n30258 & n30267;
  assign n30269 = ~n30249 & n30267;
  assign n30270 = ~n30258 & n30269;
  assign n30271 = ~n30249 & n30268;
  assign n30272 = ~pi38 & ~n60180;
  assign n30273 = ~n30198 & n30272;
  assign n30274 = ~n29985 & ~n30273;
  assign n30275 = n6305 & ~n30274;
  assign n30276 = pi100 & ~n29967;
  assign n30277 = pi38 & ~n29974;
  assign n30278 = ~pi100 & ~n30277;
  assign n30279 = ~pi38 & ~pi40;
  assign n30280 = pi87 & ~n2446;
  assign n30281 = n30279 & n30280;
  assign n30282 = n30278 & ~n30281;
  assign n30283 = pi87 & n30282;
  assign n30284 = ~n30276 & ~n30283;
  assign n30285 = ~n30275 & n30284;
  assign n30286 = n6307 & ~n30285;
  assign n30287 = pi75 & ~n29967;
  assign n30288 = pi39 & ~n29199;
  assign n30289 = n9186 & ~n30288;
  assign n30290 = n2446 & ~n29533;
  assign n30291 = ~pi40 & ~n30290;
  assign n30292 = ~pi179 & ~pi299;
  assign n30293 = ~pi156 & pi299;
  assign n30294 = ~n30292 & ~n30293;
  assign n30295 = n2681 & n30294;
  assign n30296 = n2446 & n30295;
  assign n30297 = n30291 & ~n30296;
  assign n30298 = ~pi39 & ~n30297;
  assign n30299 = n30289 & ~n30298;
  assign n30300 = n30282 & ~n30299;
  assign n30301 = ~n30276 & ~n30300;
  assign n30302 = n29661 & ~n30301;
  assign n30303 = ~n30287 & ~n30302;
  assign n30304 = ~n30286 & n30303;
  assign n30305 = ~pi54 & ~n30304;
  assign n30306 = ~n29977 & ~n30305;
  assign n30307 = ~pi74 & ~n30306;
  assign n30308 = n29970 & ~n30307;
  assign n30309 = pi55 & ~n29956;
  assign n30310 = pi54 & ~n29954;
  assign n30311 = pi163 & pi232;
  assign n30312 = ~n2680 & n29533;
  assign n30313 = n29065 & ~n30312;
  assign n30314 = n30311 & n30313;
  assign n30315 = n30291 & ~n30314;
  assign n30316 = ~pi39 & ~n30315;
  assign n30317 = n30289 & ~n30316;
  assign n30318 = pi38 & ~n29952;
  assign n30319 = ~pi100 & ~n30318;
  assign n30320 = ~n30281 & n30319;
  assign n30321 = ~n30317 & n30320;
  assign n30322 = ~n29950 & ~n30321;
  assign n30323 = n6307 & ~n30322;
  assign n30324 = n2636 & n29065;
  assign n30325 = ~n30279 & n30319;
  assign n30326 = ~n29950 & ~n30325;
  assign n30327 = ~n30324 & n30326;
  assign n30328 = n29661 & ~n30327;
  assign n30329 = ~n29949 & ~n30328;
  assign n30330 = ~n30323 & n30329;
  assign n30331 = ~pi54 & ~n30330;
  assign n30332 = ~n30310 & ~n30331;
  assign n30333 = ~pi74 & ~n30332;
  assign n30334 = n30309 & ~n30333;
  assign n30335 = n4437 & ~n30334;
  assign n30336 = ~n30308 & n30335;
  assign n30337 = ~n4437 & n29068;
  assign n30338 = ~pi75 & ~n30326;
  assign n30339 = ~n29949 & ~n30338;
  assign n30340 = ~pi54 & ~n30339;
  assign n30341 = ~n30310 & ~n30340;
  assign n30342 = ~pi74 & ~n30341;
  assign n30343 = ~n29956 & ~n30342;
  assign n30344 = ~n4437 & ~n30343;
  assign n30345 = n4438 & ~n30344;
  assign n30346 = ~n30337 & n30345;
  assign n30347 = ~n30336 & n30346;
  assign n30348 = ~n29958 & ~n30347;
  assign n30349 = ~pi79 & n30348;
  assign n30350 = ~n28442 & ~n29734;
  assign n30351 = ~pi198 & ~n30350;
  assign n30352 = ~n29732 & ~n30351;
  assign n30353 = ~pi189 & ~n30352;
  assign n30354 = ~n28443 & ~n29741;
  assign n30355 = pi189 & ~n30354;
  assign n30356 = ~pi32 & pi95;
  assign n30357 = ~pi479 & n30356;
  assign n30358 = n58824 & n30357;
  assign n30359 = pi184 & ~n30358;
  assign n30360 = ~n30355 & n30359;
  assign n30361 = ~n30353 & n30360;
  assign n30362 = ~pi189 & ~n29754;
  assign n30363 = pi189 & ~n60150;
  assign n30364 = n2598 & ~n30363;
  assign n30365 = ~n30362 & n30364;
  assign n30366 = pi182 & n30358;
  assign n30367 = ~pi184 & ~n30366;
  assign n30368 = ~n30365 & n30367;
  assign n30369 = ~pi182 & pi184;
  assign n30370 = n2680 & ~n30369;
  assign n30371 = ~n30368 & n30370;
  assign n30372 = ~n30361 & n30371;
  assign n30373 = ~n30353 & ~n30355;
  assign n30374 = n2680 & n30369;
  assign n30375 = ~n30373 & n30374;
  assign n30376 = ~n30372 & ~n30375;
  assign n30377 = n30168 & ~n30376;
  assign n30378 = n2680 & n30358;
  assign n30379 = pi160 & n30378;
  assign n30380 = ~pi153 & n29735;
  assign n30381 = n29998 & ~n30380;
  assign n30382 = ~n30379 & ~n30381;
  assign n30383 = ~pi160 & n29735;
  assign n30384 = ~pi210 & ~n30350;
  assign n30385 = pi153 & pi160;
  assign n30386 = ~n30378 & n30385;
  assign n30387 = ~n30384 & n30386;
  assign n30388 = ~n30383 & ~n30387;
  assign n30389 = ~n29732 & ~n30388;
  assign n30390 = ~n30382 & ~n30389;
  assign n30391 = pi153 & n29741;
  assign n30392 = n29744 & ~n30391;
  assign n30393 = n30049 & ~n30392;
  assign n30394 = ~pi40 & pi163;
  assign n30395 = ~n30393 & n30394;
  assign n30396 = ~n30390 & n30395;
  assign n30397 = pi153 & n29755;
  assign n30398 = n60150 & n30397;
  assign n30399 = n29760 & n29998;
  assign n30400 = ~pi40 & ~pi163;
  assign n30401 = ~n30399 & n30400;
  assign n30402 = ~n30379 & n30401;
  assign n30403 = ~n30398 & n30402;
  assign n30404 = pi299 & ~n30403;
  assign n30405 = ~pi40 & ~n30358;
  assign n30406 = n29735 & n30405;
  assign n30407 = n29998 & ~n30406;
  assign n30408 = n29744 & n30405;
  assign n30409 = n30049 & ~n30408;
  assign n30410 = ~pi153 & ~n30409;
  assign n30411 = ~n30407 & n30410;
  assign n30412 = ~n29732 & n30405;
  assign n30413 = ~n30384 & n30412;
  assign n30414 = n29998 & ~n30413;
  assign n30415 = ~n29741 & n30408;
  assign n30416 = n30049 & ~n30415;
  assign n30417 = pi153 & ~n30416;
  assign n30418 = ~n30414 & n30417;
  assign n30419 = ~n30411 & ~n30418;
  assign n30420 = pi40 & ~n2680;
  assign n30421 = pi163 & ~n30420;
  assign n30422 = ~n30419 & n30421;
  assign n30423 = pi160 & ~n30422;
  assign n30424 = pi153 & n29732;
  assign n30425 = n29735 & ~n30424;
  assign n30426 = n29998 & ~n30425;
  assign n30427 = n30395 & ~n30426;
  assign n30428 = ~n30398 & n30401;
  assign n30429 = ~pi160 & ~n30428;
  assign n30430 = ~n30427 & n30429;
  assign n30431 = ~n30423 & ~n30430;
  assign n30432 = ~n30378 & n30428;
  assign n30433 = pi299 & ~n30432;
  assign n30434 = ~n30431 & n30433;
  assign n30435 = ~n30396 & n30404;
  assign n30436 = pi40 & ~pi299;
  assign n30437 = pi184 & n29792;
  assign n30438 = ~pi184 & ~n29760;
  assign n30439 = ~pi189 & ~n30438;
  assign n30440 = ~n30437 & n30439;
  assign n30441 = pi184 & pi189;
  assign n30442 = ~n29796 & n30441;
  assign n30443 = ~n30366 & ~n30442;
  assign n30444 = ~n30440 & n30443;
  assign n30445 = n2680 & n30114;
  assign n30446 = ~n30444 & n30445;
  assign n30447 = ~n30436 & ~n30446;
  assign n30448 = ~n60181 & n30447;
  assign n30449 = n2680 & ~n30444;
  assign n30450 = ~pi40 & ~n30449;
  assign n30451 = n30114 & ~n30450;
  assign n30452 = ~n30365 & ~n30366;
  assign n30453 = n2680 & ~n30452;
  assign n30454 = ~pi184 & ~n30453;
  assign n30455 = n30128 & ~n30352;
  assign n30456 = n2680 & ~n30354;
  assign n30457 = pi189 & n30456;
  assign n30458 = n30369 & ~n30457;
  assign n30459 = ~n30455 & n30458;
  assign n30460 = ~n30454 & ~n30459;
  assign n30461 = ~pi40 & ~n30460;
  assign n30462 = ~n30351 & n30412;
  assign n30463 = n30128 & ~n30462;
  assign n30464 = n30354 & n30405;
  assign n30465 = n30125 & ~n30464;
  assign n30466 = pi182 & pi184;
  assign n30467 = ~n30420 & n30466;
  assign n30468 = ~n30465 & n30467;
  assign n30469 = ~n30463 & n30468;
  assign n30470 = n30168 & ~n30469;
  assign n30471 = ~n30461 & n30470;
  assign n30472 = ~n30451 & ~n30471;
  assign n30473 = ~n60181 & n30472;
  assign n30474 = ~n30377 & n30448;
  assign n30475 = ~pi39 & ~n60182;
  assign n30476 = n58824 & n29755;
  assign n30477 = pi156 & n29534;
  assign n30478 = ~pi166 & n29537;
  assign n30479 = ~n30477 & ~n30478;
  assign n30480 = ~n58846 & n29532;
  assign n30481 = ~n30479 & n30480;
  assign n30482 = n30476 & n30481;
  assign n30483 = ~pi40 & pi299;
  assign n30484 = ~n30482 & n30483;
  assign n30485 = ~pi189 & n29537;
  assign n30486 = pi179 & n29534;
  assign n30487 = ~n30485 & ~n30486;
  assign n30488 = n29861 & ~n30487;
  assign n30489 = n30476 & n30488;
  assign n30490 = ~pi40 & ~pi299;
  assign n30491 = ~n30489 & n30490;
  assign n30492 = pi39 & ~n30491;
  assign n30493 = pi39 & ~n30484;
  assign n30494 = ~n30491 & n30493;
  assign n30495 = ~n30484 & n30492;
  assign n30496 = pi232 & ~n60183;
  assign n30497 = ~n30475 & n30496;
  assign n30498 = ~pi40 & ~pi232;
  assign n30499 = ~pi38 & ~n30498;
  assign n30500 = ~n30497 & n30499;
  assign n30501 = ~n29985 & ~n30500;
  assign n30502 = n6305 & ~n30501;
  assign n30503 = pi87 & ~n30279;
  assign n30504 = n30278 & n30503;
  assign n30505 = ~n30276 & ~n30504;
  assign n30506 = ~n30502 & n30505;
  assign n30507 = n6307 & ~n30506;
  assign n30508 = n2598 & n2671;
  assign n30509 = n30295 & n30508;
  assign n30510 = n58824 & n30509;
  assign n30511 = n30279 & ~n30510;
  assign n30512 = n30278 & ~n30511;
  assign n30513 = ~n30276 & ~n30512;
  assign n30514 = n29661 & ~n30513;
  assign n30515 = ~n30287 & ~n30514;
  assign n30516 = ~n30507 & n30515;
  assign n30517 = ~pi54 & ~n30516;
  assign n30518 = ~n29977 & ~n30517;
  assign n30519 = ~pi74 & ~n30518;
  assign n30520 = n29970 & ~n30519;
  assign n30521 = ~pi92 & n2671;
  assign n30522 = n30311 & n30521;
  assign n30523 = n30476 & n30522;
  assign n30524 = n30279 & ~n30523;
  assign n30525 = ~pi75 & n30319;
  assign n30526 = ~n30524 & n30525;
  assign n30527 = n29951 & ~n30526;
  assign n30528 = ~pi54 & ~n30527;
  assign n30529 = ~n30310 & ~n30528;
  assign n30530 = ~pi74 & ~n30529;
  assign n30531 = n30309 & ~n30530;
  assign n30532 = n4437 & ~n30531;
  assign n30533 = ~n30520 & n30532;
  assign n30534 = n30345 & ~n30533;
  assign n30535 = ~n29958 & ~n30534;
  assign n30536 = pi79 & n30535;
  assign n30537 = ~pi34 & n29930;
  assign n30538 = ~n30536 & ~n30537;
  assign n30539 = ~n30349 & n30538;
  assign n30540 = ~pi79 & ~n29936;
  assign n30541 = n30348 & ~n30540;
  assign n30542 = n30535 & n30540;
  assign n30543 = n30537 & ~n30542;
  assign n30544 = ~n30541 & n30543;
  assign n30545 = ~n30539 & ~n30544;
  assign n30546 = pi163 & n2680;
  assign n30547 = ~n29947 & ~n30546;
  assign n30548 = ~pi150 & ~n30547;
  assign n30549 = pi150 & n29037;
  assign n30550 = n29945 & n30549;
  assign n30551 = ~n30548 & ~n30550;
  assign n30552 = pi232 & ~n30551;
  assign n30553 = ~n2635 & n30552;
  assign n30554 = n29041 & ~n30551;
  assign n30555 = pi74 & ~n60184;
  assign n30556 = ~pi74 & ~n60184;
  assign n30557 = pi165 & n2681;
  assign n30558 = ~pi38 & ~pi54;
  assign n30559 = ~n30557 & ~n30558;
  assign n30560 = n2635 & n30559;
  assign n30561 = n30556 & ~n30560;
  assign n30562 = ~n30555 & ~n30561;
  assign n30563 = ~n4437 & ~n30562;
  assign n30564 = n4438 & ~n30563;
  assign n30565 = ~n29070 & ~n30564;
  assign n30566 = pi299 & n30551;
  assign n30567 = ~pi184 & ~n29960;
  assign n30568 = ~pi185 & n30567;
  assign n30569 = pi185 & ~n30567;
  assign n30570 = n2680 & ~n30569;
  assign n30571 = ~n30568 & n30570;
  assign n30572 = ~pi299 & ~n30571;
  assign n30573 = pi232 & ~n30572;
  assign n30574 = ~n30566 & n30573;
  assign n30575 = ~n2635 & n30574;
  assign n30576 = pi74 & ~n30575;
  assign n30577 = ~pi55 & ~n30576;
  assign n30578 = ~pi143 & ~pi299;
  assign n30579 = ~pi165 & pi299;
  assign n30580 = ~n30578 & ~n30579;
  assign n30581 = n2681 & n30580;
  assign n30582 = n2635 & ~n30581;
  assign n30583 = pi54 & ~n30582;
  assign n30584 = ~n30575 & n30583;
  assign n30585 = ~pi143 & ~n60143;
  assign n30586 = pi143 & ~n29626;
  assign n30587 = pi165 & ~n30586;
  assign n30588 = ~n30585 & n30587;
  assign n30589 = pi143 & ~pi165;
  assign n30590 = n29624 & n30589;
  assign n30591 = pi38 & ~n30590;
  assign n30592 = ~n30588 & n30591;
  assign n30593 = n6305 & ~n30592;
  assign n30594 = ~n2680 & n29384;
  assign n30595 = pi151 & ~pi168;
  assign n30596 = ~n29463 & n30595;
  assign n30597 = pi168 & n29450;
  assign n30598 = ~pi168 & n29456;
  assign n30599 = ~pi151 & ~n30598;
  assign n30600 = ~n30597 & n30599;
  assign n30601 = ~n30596 & ~n30600;
  assign n30602 = ~n30594 & ~n30601;
  assign n30603 = ~n2680 & ~n29384;
  assign n30604 = n2680 & ~n29426;
  assign n30605 = ~n30603 & ~n30604;
  assign n30606 = pi151 & pi168;
  assign n30607 = ~n30605 & n30606;
  assign n30608 = pi150 & ~n30607;
  assign n30609 = ~n30602 & n30608;
  assign n30610 = ~n29263 & ~n30603;
  assign n30611 = pi168 & n30610;
  assign n30612 = ~n29389 & ~n30603;
  assign n30613 = ~pi168 & n30612;
  assign n30614 = pi151 & ~n30613;
  assign n30615 = ~n30611 & n30614;
  assign n30616 = pi168 & n29242;
  assign n30617 = pi168 & n2680;
  assign n30618 = n29384 & ~n30617;
  assign n30619 = ~pi151 & ~n30618;
  assign n30620 = ~n30616 & n30619;
  assign n30621 = ~pi150 & ~n30620;
  assign n30622 = ~n30615 & n30621;
  assign n30623 = pi299 & ~n30622;
  assign n30624 = ~n30609 & n30623;
  assign n30625 = ~n29229 & ~n30594;
  assign n30626 = ~pi173 & ~n30625;
  assign n30627 = n2680 & ~n29197;
  assign n30628 = pi173 & ~n30603;
  assign n30629 = ~n30627 & n30628;
  assign n30630 = pi185 & ~n30629;
  assign n30631 = ~n30626 & n30630;
  assign n30632 = pi173 & n30610;
  assign n30633 = ~n29242 & ~n30594;
  assign n30634 = ~pi173 & ~n30633;
  assign n30635 = ~pi185 & ~n30634;
  assign n30636 = pi173 & ~n30610;
  assign n30637 = ~pi173 & ~n29242;
  assign n30638 = ~n30594 & n30637;
  assign n30639 = ~n30636 & ~n30638;
  assign n30640 = ~pi185 & ~n30639;
  assign n30641 = ~n30632 & n30635;
  assign n30642 = pi190 & ~n60185;
  assign n30643 = ~n30631 & n30642;
  assign n30644 = pi173 & ~n29377;
  assign n30645 = ~pi173 & ~n29372;
  assign n30646 = n2680 & ~n30645;
  assign n30647 = ~pi173 & n29372;
  assign n30648 = pi173 & n29377;
  assign n30649 = ~n30647 & ~n30648;
  assign n30650 = n2680 & ~n30649;
  assign n30651 = ~n30644 & n30646;
  assign n30652 = pi185 & ~n30594;
  assign n30653 = ~n60186 & n30652;
  assign n30654 = pi173 & n30612;
  assign n30655 = ~pi173 & n29384;
  assign n30656 = ~pi185 & ~n30655;
  assign n30657 = ~n30654 & n30656;
  assign n30658 = ~pi190 & ~n30657;
  assign n30659 = ~n30653 & n30658;
  assign n30660 = ~pi299 & ~n30659;
  assign n30661 = ~n30643 & n30660;
  assign n30662 = pi232 & ~n30661;
  assign n30663 = ~n30624 & n30662;
  assign n30664 = ~pi232 & n29384;
  assign n30665 = ~pi39 & ~n30664;
  assign n30666 = ~n30663 & n30665;
  assign n30667 = pi178 & ~n29539;
  assign n30668 = ~pi178 & ~n29558;
  assign n30669 = pi190 & ~n30668;
  assign n30670 = ~n30667 & n30669;
  assign n30671 = pi178 & ~pi190;
  assign n30672 = n29546 & n30671;
  assign n30673 = ~n30670 & ~n30672;
  assign n30674 = pi222 & pi224;
  assign n30675 = pi224 & n58844;
  assign n30676 = n2828 & n30674;
  assign n30677 = n2791 & n60187;
  assign n30678 = ~n30673 & n30677;
  assign n30679 = pi168 & n29558;
  assign n30680 = pi157 & n29546;
  assign n30681 = ~n30679 & ~n30680;
  assign n30682 = pi216 & pi221;
  assign n30683 = pi299 & n29532;
  assign n30684 = n2851 & n30682;
  assign n30685 = n2844 & n60188;
  assign n30686 = ~n30681 & n30685;
  assign n30687 = pi232 & n29065;
  assign n30688 = ~n30686 & n30687;
  assign n30689 = ~pi178 & ~pi299;
  assign n30690 = n2680 & n30480;
  assign n30691 = n2844 & n29532;
  assign n30692 = ~n30681 & n60189;
  assign n30693 = pi299 & ~n30692;
  assign n30694 = ~n30689 & ~n30693;
  assign n30695 = n29065 & ~n30694;
  assign n30696 = pi178 & ~n29585;
  assign n30697 = ~pi190 & ~n30696;
  assign n30698 = ~pi299 & ~n30697;
  assign n30699 = ~n30695 & ~n30698;
  assign n30700 = n2790 & ~n29065;
  assign n30701 = n29572 & ~n30700;
  assign n30702 = pi178 & n30701;
  assign n30703 = ~n29574 & n30702;
  assign n30704 = ~pi178 & n30701;
  assign n30705 = ~n29595 & n30704;
  assign n30706 = ~pi299 & ~n29573;
  assign n30707 = pi190 & n30706;
  assign n30708 = ~n30705 & n30707;
  assign n30709 = ~n30703 & n30708;
  assign n30710 = pi232 & ~n30709;
  assign n30711 = ~n30699 & n30710;
  assign n30712 = ~n30678 & n30688;
  assign n30713 = ~pi232 & n29065;
  assign n30714 = pi39 & ~n30713;
  assign n30715 = ~n60190 & n30714;
  assign n30716 = ~pi38 & ~n30715;
  assign n30717 = ~n30666 & n30716;
  assign n30718 = n30593 & ~n30717;
  assign n30719 = pi100 & ~n30574;
  assign n30720 = pi38 & ~n30581;
  assign n30721 = ~pi100 & ~n30720;
  assign n30722 = pi87 & n30721;
  assign n30723 = n2903 & ~n30720;
  assign n30724 = ~n29066 & n60191;
  assign n30725 = ~n30719 & ~n30724;
  assign n30726 = ~n30718 & n30725;
  assign n30727 = n6307 & ~n30726;
  assign n30728 = pi75 & ~n30574;
  assign n30729 = ~pi157 & pi299;
  assign n30730 = ~n30689 & ~n30729;
  assign n30731 = n2681 & n30730;
  assign n30732 = n60146 & n30731;
  assign n30733 = n29066 & ~n30732;
  assign n30734 = n30721 & ~n30733;
  assign n30735 = ~n30719 & ~n30734;
  assign n30736 = n29661 & ~n30735;
  assign n30737 = ~n30728 & ~n30736;
  assign n30738 = ~n30727 & n30737;
  assign n30739 = ~pi54 & ~n30738;
  assign n30740 = ~n30584 & ~n30739;
  assign n30741 = ~pi74 & ~n30740;
  assign n30742 = n30577 & ~n30741;
  assign n30743 = pi55 & ~n30555;
  assign n30744 = pi150 & n2681;
  assign n30745 = ~pi92 & n60146;
  assign n30746 = n30744 & n30745;
  assign n30747 = n29065 & n30558;
  assign n30748 = ~n30746 & n30747;
  assign n30749 = ~n30559 & ~n30748;
  assign n30750 = n2635 & ~n30749;
  assign n30751 = n30556 & ~n30750;
  assign n30752 = n30743 & ~n30751;
  assign n30753 = n4437 & ~n30752;
  assign n30754 = ~n30742 & n30753;
  assign n30755 = ~n30565 & ~n30754;
  assign n30756 = ~pi74 & n2635;
  assign n30757 = ~n30557 & n30756;
  assign n30758 = ~n60184 & ~n30757;
  assign n30759 = n2635 & ~n30557;
  assign n30760 = ~n60184 & ~n30759;
  assign n30761 = ~n2635 & ~n30552;
  assign n30762 = n2635 & n30557;
  assign n30763 = ~n4438 & ~n30762;
  assign n30764 = ~n30761 & n30763;
  assign n30765 = ~n4438 & ~n30760;
  assign n30766 = ~n30555 & n60192;
  assign n30767 = ~n4438 & ~n30758;
  assign n30768 = ~n30755 & ~n60193;
  assign n30769 = pi118 & n30768;
  assign n30770 = ~pi79 & n30537;
  assign n30771 = n2783 & ~n28517;
  assign n30772 = ~pi178 & n28517;
  assign n30773 = pi178 & ~n28507;
  assign n30774 = ~pi190 & ~n30773;
  assign n30775 = ~n30772 & n30774;
  assign n30776 = ~pi178 & pi190;
  assign n30777 = n58842 & n30776;
  assign n30778 = ~n30775 & ~n30777;
  assign n30779 = n2791 & ~n30778;
  assign n30780 = ~pi178 & ~n2790;
  assign n30781 = n29846 & n30780;
  assign n30782 = ~n30771 & ~n30781;
  assign n30783 = pi190 & ~n30782;
  assign n30784 = pi178 & ~n29874;
  assign n30785 = ~n30771 & n30784;
  assign n30786 = ~n2792 & ~n28517;
  assign n30787 = ~pi178 & ~n30786;
  assign n30788 = ~pi190 & ~n30787;
  assign n30789 = ~pi190 & ~n30785;
  assign n30790 = ~n30787 & n30789;
  assign n30791 = ~n30785 & n30788;
  assign n30792 = ~n30783 & ~n60194;
  assign n30793 = ~n30771 & ~n30779;
  assign n30794 = n60187 & ~n60195;
  assign n30795 = ~pi168 & ~n29844;
  assign n30796 = pi168 & ~n60157;
  assign n30797 = ~pi157 & ~n30796;
  assign n30798 = ~n30795 & n30797;
  assign n30799 = pi157 & ~pi168;
  assign n30800 = n29855 & n30799;
  assign n30801 = ~n30771 & ~n30800;
  assign n30802 = ~pi157 & n60157;
  assign n30803 = pi168 & ~n30802;
  assign n30804 = pi157 & ~n29855;
  assign n30805 = ~pi157 & ~pi168;
  assign n30806 = ~n29844 & n30805;
  assign n30807 = ~n30804 & ~n30806;
  assign n30808 = ~n30803 & n30807;
  assign n30809 = ~n30771 & ~n30808;
  assign n30810 = ~n30798 & n30801;
  assign n30811 = n60188 & ~n60196;
  assign n30812 = pi232 & ~n30811;
  assign n30813 = pi232 & ~n30794;
  assign n30814 = ~n30811 & n30813;
  assign n30815 = ~n30794 & n30812;
  assign n30816 = pi224 & n60084;
  assign n30817 = ~n2792 & n60187;
  assign n30818 = pi216 & ~n2845;
  assign n30819 = n2853 & n30818;
  assign n30820 = ~n2845 & n60188;
  assign n30821 = ~n60198 & ~n60199;
  assign n30822 = ~n28517 & ~n30821;
  assign n30823 = n28532 & n29864;
  assign n30824 = ~n28517 & n60199;
  assign n30825 = ~pi232 & ~n30824;
  assign n30826 = ~n30823 & n30825;
  assign n30827 = ~pi232 & ~n30822;
  assign n30828 = pi39 & ~n60200;
  assign n30829 = ~n60197 & n30828;
  assign n30830 = pi173 & n60166;
  assign n30831 = ~pi173 & n2621;
  assign n30832 = n29754 & n30831;
  assign n30833 = ~n30830 & ~n30832;
  assign n30834 = ~pi190 & n2680;
  assign n30835 = ~n30833 & n30834;
  assign n30836 = ~pi173 & pi190;
  assign n30837 = n29767 & n30836;
  assign n30838 = pi185 & ~n30837;
  assign n30839 = ~n30835 & n30838;
  assign n30840 = ~pi173 & n29732;
  assign n30841 = n29792 & ~n30840;
  assign n30842 = ~pi190 & ~n30841;
  assign n30843 = pi173 & n29796;
  assign n30844 = pi190 & ~n30843;
  assign n30845 = pi190 & n30456;
  assign n30846 = ~n30843 & n30845;
  assign n30847 = n30456 & n30844;
  assign n30848 = ~pi185 & ~n60201;
  assign n30849 = ~n30842 & n30848;
  assign n30850 = ~n30839 & ~n30849;
  assign n30851 = ~n2680 & ~n30352;
  assign n30852 = ~pi299 & ~n30851;
  assign n30853 = ~n30850 & n30852;
  assign n30854 = n29759 & n30595;
  assign n30855 = pi168 & ~n60150;
  assign n30856 = ~pi168 & ~n29754;
  assign n30857 = ~pi151 & ~n30856;
  assign n30858 = ~pi151 & ~n30855;
  assign n30859 = ~n30856 & n30858;
  assign n30860 = ~n30855 & n30857;
  assign n30861 = ~n30854 & ~n60202;
  assign n30862 = n29756 & ~n30861;
  assign n30863 = pi150 & ~n30862;
  assign n30864 = ~pi151 & n29732;
  assign n30865 = n29735 & ~n30864;
  assign n30866 = ~pi168 & ~n30865;
  assign n30867 = ~pi151 & n29741;
  assign n30868 = n29744 & ~n30867;
  assign n30869 = n30617 & ~n30868;
  assign n30870 = ~pi150 & ~n30869;
  assign n30871 = ~n30866 & n30870;
  assign n30872 = ~n30863 & ~n30871;
  assign n30873 = ~n29732 & ~n30384;
  assign n30874 = ~n2680 & ~n30873;
  assign n30875 = pi299 & ~n30874;
  assign n30876 = ~n30872 & n30875;
  assign n30877 = ~n30853 & ~n30876;
  assign n30878 = pi232 & ~n30877;
  assign n30879 = ~n60122 & ~n30350;
  assign n30880 = ~pi232 & ~n29732;
  assign n30881 = ~n30879 & n30880;
  assign n30882 = ~pi39 & ~n30881;
  assign n30883 = ~n30878 & n30882;
  assign n30884 = ~n30829 & ~n30883;
  assign n30885 = ~pi38 & ~n30884;
  assign n30886 = n30593 & ~n30885;
  assign n30887 = ~n30719 & ~n60191;
  assign n30888 = ~n30886 & n30887;
  assign n30889 = n6307 & ~n30888;
  assign n30890 = ~pi87 & n2634;
  assign n30891 = ~n30731 & n30890;
  assign n30892 = n58822 & n30891;
  assign n30893 = n30721 & ~n30892;
  assign n30894 = ~n30719 & ~n30893;
  assign n30895 = n29661 & ~n30894;
  assign n30896 = ~n30728 & ~n30895;
  assign n30897 = ~n30889 & n30896;
  assign n30898 = ~pi54 & ~n30897;
  assign n30899 = ~n30584 & ~n30898;
  assign n30900 = ~pi74 & ~n30899;
  assign n30901 = n30577 & ~n30900;
  assign n30902 = pi54 & n30557;
  assign n30903 = ~pi92 & n2635;
  assign n30904 = n30890 & n30903;
  assign n30905 = n2672 & n6307;
  assign n30906 = n58815 & n6310;
  assign n30907 = ~n30744 & n60203;
  assign n30908 = ~n30902 & n30907;
  assign n30909 = n58822 & n30908;
  assign n30910 = n30561 & ~n30909;
  assign n30911 = n30743 & ~n30910;
  assign n30912 = n4437 & ~n30911;
  assign n30913 = ~n30901 & n30912;
  assign n30914 = n30564 & ~n30913;
  assign n30915 = ~n60193 & ~n30914;
  assign n30916 = ~pi118 & n30915;
  assign n30917 = ~n30770 & ~n30916;
  assign n30918 = ~n30769 & n30917;
  assign n30919 = ~pi118 & ~n29935;
  assign n30920 = n30768 & n30919;
  assign n30921 = n30915 & ~n30919;
  assign n30922 = n30770 & ~n30921;
  assign n30923 = ~n30920 & n30922;
  assign n30924 = ~n30918 & ~n30923;
  assign n30925 = ~pi34 & n29937;
  assign n30926 = ~pi33 & ~n30925;
  assign n30927 = pi149 & pi157;
  assign n30928 = n29034 & ~n30927;
  assign n30929 = pi232 & n30928;
  assign n30930 = pi75 & ~n30929;
  assign n30931 = pi100 & ~n30929;
  assign n30932 = ~n30930 & ~n30931;
  assign n30933 = pi164 & n2681;
  assign n30934 = pi164 & n29045;
  assign n30935 = n2635 & n30933;
  assign n30936 = n30932 & ~n60204;
  assign n30937 = ~pi74 & ~n30936;
  assign n30938 = pi169 & n2681;
  assign n30939 = n2635 & n30938;
  assign n30940 = pi169 & n29045;
  assign n30941 = n30932 & ~n60205;
  assign n30942 = pi74 & ~n30941;
  assign n30943 = ~n4438 & ~n30942;
  assign n30944 = ~n4438 & ~n30937;
  assign n30945 = ~n30942 & n30944;
  assign n30946 = ~n30937 & n30943;
  assign n30947 = pi299 & ~n30928;
  assign n30948 = pi178 & pi183;
  assign n30949 = n29074 & ~n30948;
  assign n30950 = ~pi299 & ~n30949;
  assign n30951 = pi232 & ~n30950;
  assign n30952 = pi232 & ~n30947;
  assign n30953 = ~n30950 & n30952;
  assign n30954 = ~n30947 & n30951;
  assign n30955 = pi100 & ~n60207;
  assign n30956 = pi75 & ~n60207;
  assign n30957 = ~n30955 & ~n30956;
  assign n30958 = pi191 & ~pi299;
  assign n30959 = pi169 & pi299;
  assign n30960 = ~n30958 & ~n30959;
  assign n30961 = n29045 & ~n30960;
  assign n30962 = n30957 & ~n30961;
  assign n30963 = pi74 & ~n30962;
  assign n30964 = ~pi55 & ~n30963;
  assign n30965 = ~pi186 & ~pi299;
  assign n30966 = ~pi164 & pi299;
  assign n30967 = ~n30965 & ~n30966;
  assign n30968 = n2681 & n30967;
  assign n30969 = n2635 & n30968;
  assign n30970 = n30957 & ~n30969;
  assign n30971 = pi54 & ~n30970;
  assign n30972 = ~pi186 & ~n60143;
  assign n30973 = pi186 & ~n29626;
  assign n30974 = pi164 & ~n30973;
  assign n30975 = ~n30972 & n30974;
  assign n30976 = ~pi164 & pi186;
  assign n30977 = n29624 & n30976;
  assign n30978 = ~n30975 & ~n30977;
  assign n30979 = pi38 & ~n30978;
  assign n30980 = ~pi152 & n29549;
  assign n30981 = ~pi154 & ~n29545;
  assign n30982 = ~n30980 & n30981;
  assign n30983 = pi152 & n29560;
  assign n30984 = n29541 & ~n30983;
  assign n30985 = pi154 & ~n30984;
  assign n30986 = n29532 & ~n30985;
  assign n30987 = ~n30982 & n30986;
  assign n30988 = n29554 & ~n30987;
  assign n30989 = ~pi176 & ~pi299;
  assign n30990 = n29585 & n30989;
  assign n30991 = ~pi174 & ~n29576;
  assign n30992 = pi174 & n60139;
  assign n30993 = ~n29576 & ~n30992;
  assign n30994 = ~pi299 & ~n30993;
  assign n30995 = ~pi299 & ~n30991;
  assign n30996 = ~n29598 & n30995;
  assign n30997 = n29599 & ~n30991;
  assign n30998 = ~n30990 & ~n60208;
  assign n30999 = ~n30988 & n30998;
  assign n31000 = pi232 & ~n30999;
  assign n31001 = pi39 & ~n29612;
  assign n31002 = ~pi176 & pi232;
  assign n31003 = ~n30988 & ~n60208;
  assign n31004 = ~pi299 & n29585;
  assign n31005 = n31003 & ~n31004;
  assign n31006 = n31002 & ~n31005;
  assign n31007 = pi176 & pi232;
  assign n31008 = ~n31003 & n31007;
  assign n31009 = n31001 & ~n31008;
  assign n31010 = ~n31006 & n31009;
  assign n31011 = ~n31000 & n31001;
  assign n31012 = ~pi183 & ~n29356;
  assign n31013 = pi183 & ~n29303;
  assign n31014 = ~n31012 & ~n31013;
  assign n31015 = ~pi174 & ~n31014;
  assign n31016 = pi183 & n29287;
  assign n31017 = ~pi183 & n29277;
  assign n31018 = pi174 & ~n31017;
  assign n31019 = pi183 & ~n29287;
  assign n31020 = ~pi183 & ~n29277;
  assign n31021 = ~n31019 & ~n31020;
  assign n31022 = pi174 & ~n31021;
  assign n31023 = ~n31016 & n31018;
  assign n31024 = pi180 & ~n60210;
  assign n31025 = pi180 & ~n31015;
  assign n31026 = ~n60210 & n31025;
  assign n31027 = ~n31015 & n31024;
  assign n31028 = ~pi95 & n31014;
  assign n31029 = ~pi174 & ~n29117;
  assign n31030 = ~n31028 & n31029;
  assign n31031 = pi183 & n2680;
  assign n31032 = ~n29197 & ~n31031;
  assign n31033 = pi183 & n29263;
  assign n31034 = pi174 & ~n31033;
  assign n31035 = ~n31032 & n31034;
  assign n31036 = ~pi180 & ~n31035;
  assign n31037 = ~n31030 & n31036;
  assign n31038 = ~pi193 & ~n31037;
  assign n31039 = ~n60211 & n31038;
  assign n31040 = ~pi183 & ~n29230;
  assign n31041 = pi183 & ~n29243;
  assign n31042 = pi174 & ~n31041;
  assign n31043 = ~n31040 & n31042;
  assign n31044 = ~pi183 & n29372;
  assign n31045 = pi183 & n29384;
  assign n31046 = ~n31044 & ~n31045;
  assign n31047 = n2680 & ~n31046;
  assign n31048 = ~pi174 & ~n29198;
  assign n31049 = pi183 & ~n29386;
  assign n31050 = ~pi183 & n29374;
  assign n31051 = ~pi174 & ~n31050;
  assign n31052 = ~n31049 & n31051;
  assign n31053 = ~pi174 & ~n31049;
  assign n31054 = ~n31050 & n31053;
  assign n31055 = ~n31047 & n31048;
  assign n31056 = ~pi180 & ~n60212;
  assign n31057 = ~n31043 & n31056;
  assign n31058 = pi183 & n29305;
  assign n31059 = ~pi183 & ~n29337;
  assign n31060 = ~pi174 & ~n31059;
  assign n31061 = ~pi174 & ~n31058;
  assign n31062 = ~n31059 & n31061;
  assign n31063 = ~n31058 & n31060;
  assign n31064 = ~pi183 & ~n29271;
  assign n31065 = pi183 & ~n29284;
  assign n31066 = pi174 & ~n31065;
  assign n31067 = ~n31064 & n31066;
  assign n31068 = pi180 & ~n31067;
  assign n31069 = pi180 & ~n60213;
  assign n31070 = ~n31067 & n31069;
  assign n31071 = ~n60213 & n31068;
  assign n31072 = ~n31057 & ~n60214;
  assign n31073 = pi193 & ~n31072;
  assign n31074 = ~pi299 & ~n31073;
  assign n31075 = ~n60211 & ~n31037;
  assign n31076 = ~pi193 & ~n31075;
  assign n31077 = pi193 & ~n60214;
  assign n31078 = pi193 & ~n31057;
  assign n31079 = ~n60214 & n31078;
  assign n31080 = ~n31057 & n31077;
  assign n31081 = ~n31076 & ~n60215;
  assign n31082 = ~pi299 & ~n31081;
  assign n31083 = ~n31039 & n31074;
  assign n31084 = ~pi158 & pi299;
  assign n31085 = pi152 & ~n29428;
  assign n31086 = ~pi152 & ~n29437;
  assign n31087 = pi172 & ~n31086;
  assign n31088 = pi172 & ~n31085;
  assign n31089 = ~n31086 & n31088;
  assign n31090 = ~n31085 & n31087;
  assign n31091 = ~pi152 & n29439;
  assign n31092 = pi152 & n29431;
  assign n31093 = ~pi172 & ~n31092;
  assign n31094 = ~pi172 & ~n31091;
  assign n31095 = ~n31092 & n31094;
  assign n31096 = ~n31091 & n31093;
  assign n31097 = ~n60217 & ~n60218;
  assign n31098 = n31084 & ~n31097;
  assign n31099 = pi158 & pi299;
  assign n31100 = pi152 & ~n29490;
  assign n31101 = ~pi152 & ~n29484;
  assign n31102 = ~pi172 & ~n31101;
  assign n31103 = ~pi172 & ~n31100;
  assign n31104 = ~n31101 & n31103;
  assign n31105 = ~n31100 & n31102;
  assign n31106 = pi152 & ~n29492;
  assign n31107 = ~pi152 & n29486;
  assign n31108 = pi172 & ~n31107;
  assign n31109 = pi172 & ~n31106;
  assign n31110 = ~n31107 & n31109;
  assign n31111 = ~n31106 & n31108;
  assign n31112 = ~n60219 & ~n60220;
  assign n31113 = n31099 & ~n31112;
  assign n31114 = ~n31098 & ~n31113;
  assign n31115 = pi149 & ~n31114;
  assign n31116 = pi152 & ~n29513;
  assign n31117 = ~pi152 & ~n29505;
  assign n31118 = pi172 & ~n31117;
  assign n31119 = ~n31116 & n31118;
  assign n31120 = pi152 & n29517;
  assign n31121 = ~pi152 & ~n29508;
  assign n31122 = ~pi172 & ~n31121;
  assign n31123 = ~pi172 & ~n31120;
  assign n31124 = ~n31121 & n31123;
  assign n31125 = ~n31120 & n31122;
  assign n31126 = ~n31119 & ~n60221;
  assign n31127 = n31099 & ~n31126;
  assign n31128 = pi152 & ~n29450;
  assign n31129 = ~pi152 & ~n29456;
  assign n31130 = pi172 & ~n31129;
  assign n31131 = ~n31128 & n31130;
  assign n31132 = pi152 & ~n29426;
  assign n31133 = ~pi152 & ~n29463;
  assign n31134 = ~pi172 & ~n31133;
  assign n31135 = ~pi172 & ~n31132;
  assign n31136 = ~n31133 & n31135;
  assign n31137 = ~n31132 & n31134;
  assign n31138 = ~n29427 & n31084;
  assign n31139 = ~n60222 & n31138;
  assign n31140 = ~n31131 & n31139;
  assign n31141 = ~n31127 & ~n31140;
  assign n31142 = ~pi149 & ~n31141;
  assign n31143 = ~pi149 & ~n31140;
  assign n31144 = ~n31127 & n31143;
  assign n31145 = pi149 & ~n31098;
  assign n31146 = pi149 & ~n31113;
  assign n31147 = ~n31098 & n31146;
  assign n31148 = ~n31113 & n31145;
  assign n31149 = ~n31144 & ~n60223;
  assign n31150 = ~n31115 & ~n31142;
  assign n31151 = ~n60216 & ~n60224;
  assign n31152 = pi232 & ~n31151;
  assign n31153 = ~pi39 & ~n29195;
  assign n31154 = ~n31152 & n31153;
  assign n31155 = ~n60209 & ~n31154;
  assign n31156 = ~pi38 & ~n31155;
  assign n31157 = ~n30979 & ~n31156;
  assign n31158 = ~pi100 & ~n31157;
  assign n31159 = ~pi87 & ~n30955;
  assign n31160 = ~n31158 & n31159;
  assign n31161 = pi38 & n30968;
  assign n31162 = ~pi100 & n31161;
  assign n31163 = ~n30955 & ~n31162;
  assign n31164 = pi87 & ~n30324;
  assign n31165 = n31163 & n31164;
  assign n31166 = n6307 & ~n31165;
  assign n31167 = ~n31160 & n31166;
  assign n31168 = ~pi154 & pi299;
  assign n31169 = pi232 & ~n31168;
  assign n31170 = n2680 & ~n30989;
  assign n31171 = n31169 & n31170;
  assign n31172 = n60146 & ~n31171;
  assign n31173 = n30324 & ~n31172;
  assign n31174 = n31163 & ~n31173;
  assign n31175 = n29661 & ~n31174;
  assign n31176 = ~n30956 & ~n31175;
  assign n31177 = ~n31167 & n31176;
  assign n31178 = ~pi54 & ~n31177;
  assign n31179 = ~n30971 & ~n31178;
  assign n31180 = ~pi74 & ~n31179;
  assign n31181 = n30964 & ~n31180;
  assign n31182 = pi55 & ~n30942;
  assign n31183 = pi54 & ~n30936;
  assign n31184 = ~pi92 & n30932;
  assign n31185 = pi149 & n2681;
  assign n31186 = ~pi38 & ~n31185;
  assign n31187 = n60146 & n31186;
  assign n31188 = pi38 & ~n30933;
  assign n31189 = n2635 & ~n29653;
  assign n31190 = ~pi100 & ~n29653;
  assign n31191 = ~n31188 & n31190;
  assign n31192 = ~pi75 & n31191;
  assign n31193 = ~n31188 & n31189;
  assign n31194 = ~n31187 & n60225;
  assign n31195 = ~pi92 & ~n30930;
  assign n31196 = n6305 & ~n31188;
  assign n31197 = ~pi39 & ~n31185;
  assign n31198 = n29533 & n31197;
  assign n31199 = n29065 & ~n31198;
  assign n31200 = ~pi38 & ~n31199;
  assign n31201 = n31196 & ~n31200;
  assign n31202 = pi87 & n31191;
  assign n31203 = ~n30931 & ~n31202;
  assign n31204 = ~n31201 & n31203;
  assign n31205 = ~pi75 & ~n31204;
  assign n31206 = n31195 & ~n31205;
  assign n31207 = n31184 & ~n31194;
  assign n31208 = pi92 & n30932;
  assign n31209 = ~n60225 & n31208;
  assign n31210 = ~pi54 & ~n31209;
  assign n31211 = ~n60226 & n31210;
  assign n31212 = ~n31183 & ~n31211;
  assign n31213 = ~pi74 & ~n31212;
  assign n31214 = n31182 & ~n31213;
  assign n31215 = n4437 & ~n31214;
  assign n31216 = ~n31181 & n31215;
  assign n31217 = pi38 & n30933;
  assign n31218 = pi38 & n60204;
  assign n31219 = n2635 & n31217;
  assign n31220 = n30932 & ~n60227;
  assign n31221 = ~n31183 & n31220;
  assign n31222 = ~pi74 & ~n31221;
  assign n31223 = ~n30942 & ~n31222;
  assign n31224 = ~n4437 & ~n31223;
  assign n31225 = n4438 & ~n31224;
  assign n31226 = ~n30337 & n31225;
  assign n31227 = ~n31216 & n31226;
  assign n31228 = ~n60206 & ~n31227;
  assign n31229 = ~n30926 & ~n31228;
  assign n31230 = pi154 & ~n29844;
  assign n31231 = ~pi154 & ~n29855;
  assign n31232 = ~pi152 & ~n31231;
  assign n31233 = ~n31230 & n31232;
  assign n31234 = pi152 & pi154;
  assign n31235 = n60157 & n31234;
  assign n31236 = ~n31233 & ~n31235;
  assign n31237 = n29532 & ~n31236;
  assign n31238 = pi299 & ~n31237;
  assign n31239 = pi39 & pi232;
  assign n31240 = ~pi174 & n60160;
  assign n31241 = pi174 & n29868;
  assign n31242 = ~pi299 & ~n31241;
  assign n31243 = ~n31240 & n31242;
  assign n31244 = pi176 & ~n31243;
  assign n31245 = ~pi174 & n60162;
  assign n31246 = ~pi299 & ~n31245;
  assign n31247 = ~pi176 & ~n31246;
  assign n31248 = ~n31244 & ~n31247;
  assign n31249 = n31002 & ~n31246;
  assign n31250 = n31007 & ~n31243;
  assign n31251 = ~n31249 & ~n31250;
  assign n31252 = pi39 & ~n31251;
  assign n31253 = n31239 & ~n31248;
  assign n31254 = pi39 & ~n31238;
  assign n31255 = ~n31251 & n31254;
  assign n31256 = ~n31238 & n60228;
  assign n31257 = ~n30352 & n31031;
  assign n31258 = ~pi183 & n29757;
  assign n31259 = pi193 & ~n31258;
  assign n31260 = ~n31257 & n31259;
  assign n31261 = ~n29792 & n31031;
  assign n31262 = ~pi183 & n29761;
  assign n31263 = ~pi193 & ~n31262;
  assign n31264 = ~n31261 & n31263;
  assign n31265 = ~pi174 & ~n31264;
  assign n31266 = ~n31260 & n31265;
  assign n31267 = pi183 & ~n30456;
  assign n31268 = ~pi183 & ~n29767;
  assign n31269 = pi193 & ~n31268;
  assign n31270 = ~n31267 & n31269;
  assign n31271 = ~pi193 & n31031;
  assign n31272 = ~n29796 & n31271;
  assign n31273 = ~n31270 & ~n31272;
  assign n31274 = pi174 & ~n31273;
  assign n31275 = pi180 & n29782;
  assign n31276 = ~pi299 & ~n31275;
  assign n31277 = ~n31274 & n31276;
  assign n31278 = ~pi174 & ~n31258;
  assign n31279 = ~n31257 & n31278;
  assign n31280 = pi183 & n30456;
  assign n31281 = ~pi183 & n29767;
  assign n31282 = pi174 & ~n31281;
  assign n31283 = ~n31280 & n31282;
  assign n31284 = ~n31279 & ~n31283;
  assign n31285 = pi193 & ~n31284;
  assign n31286 = ~pi174 & n29792;
  assign n31287 = pi174 & n29796;
  assign n31288 = n31031 & ~n31287;
  assign n31289 = ~n31286 & n31288;
  assign n31290 = ~pi174 & ~pi183;
  assign n31291 = n29761 & n31290;
  assign n31292 = ~pi193 & ~n31291;
  assign n31293 = ~n31289 & n31292;
  assign n31294 = ~n31285 & ~n31293;
  assign n31295 = n31276 & ~n31294;
  assign n31296 = ~n31266 & n31277;
  assign n31297 = pi172 & n29732;
  assign n31298 = ~pi152 & n29735;
  assign n31299 = ~n31297 & n31298;
  assign n31300 = pi149 & n2680;
  assign n31301 = pi172 & n29741;
  assign n31302 = pi152 & n29744;
  assign n31303 = pi152 & ~n31301;
  assign n31304 = n29744 & n31303;
  assign n31305 = ~n31301 & n31302;
  assign n31306 = n31300 & ~n60231;
  assign n31307 = n29744 & ~n31301;
  assign n31308 = pi152 & ~n31307;
  assign n31309 = n29735 & ~n31297;
  assign n31310 = ~pi152 & ~n31309;
  assign n31311 = ~n31308 & ~n31310;
  assign n31312 = n31300 & ~n31311;
  assign n31313 = ~n31299 & n31306;
  assign n31314 = ~pi152 & n29757;
  assign n31315 = pi172 & ~n29767;
  assign n31316 = ~n31314 & n31315;
  assign n31317 = ~pi152 & n29761;
  assign n31318 = ~pi172 & ~n31317;
  assign n31319 = ~pi149 & ~n31318;
  assign n31320 = ~n29767 & ~n31314;
  assign n31321 = pi172 & ~n31320;
  assign n31322 = ~pi152 & ~pi172;
  assign n31323 = n29761 & n31322;
  assign n31324 = ~n31321 & ~n31323;
  assign n31325 = ~pi149 & ~n31324;
  assign n31326 = ~n31316 & n31319;
  assign n31327 = pi158 & n29782;
  assign n31328 = pi299 & ~n31327;
  assign n31329 = ~n60233 & n31328;
  assign n31330 = ~n60232 & n31329;
  assign n31331 = n29912 & ~n31330;
  assign n31332 = n29912 & ~n60230;
  assign n31333 = ~n31330 & n31332;
  assign n31334 = ~n60230 & n31331;
  assign n31335 = ~n60229 & ~n60234;
  assign n31336 = ~pi38 & ~n31335;
  assign n31337 = ~pi87 & ~n30979;
  assign n31338 = ~n31336 & n31337;
  assign n31339 = pi87 & ~n31161;
  assign n31340 = ~pi100 & ~n31339;
  assign n31341 = ~n31338 & n31340;
  assign n31342 = ~n30955 & ~n31341;
  assign n31343 = n6307 & ~n31342;
  assign n31344 = n59291 & n31171;
  assign n31345 = n59171 & n31344;
  assign n31346 = n31163 & ~n31345;
  assign n31347 = n29661 & ~n31346;
  assign n31348 = ~n30956 & ~n31347;
  assign n31349 = ~n31343 & n31348;
  assign n31350 = ~pi54 & ~n31349;
  assign n31351 = ~n30971 & ~n31350;
  assign n31352 = ~pi74 & ~n31351;
  assign n31353 = n30964 & ~n31352;
  assign n31354 = n9186 & n31185;
  assign n31355 = n59171 & n31354;
  assign n31356 = ~n31217 & ~n31355;
  assign n31357 = n2635 & ~n31356;
  assign n31358 = n59171 & n31185;
  assign n31359 = ~pi38 & ~n31358;
  assign n31360 = n31196 & ~n31359;
  assign n31361 = pi38 & pi87;
  assign n31362 = ~pi100 & n31361;
  assign n31363 = n2903 & n31217;
  assign n31364 = n30933 & n31362;
  assign n31365 = ~n30931 & ~n60235;
  assign n31366 = ~n31360 & n31365;
  assign n31367 = ~pi75 & ~n31366;
  assign n31368 = n31195 & ~n31367;
  assign n31369 = n31184 & ~n31357;
  assign n31370 = pi92 & n31220;
  assign n31371 = n31208 & ~n60227;
  assign n31372 = ~pi54 & ~n60237;
  assign n31373 = ~n60236 & n31372;
  assign n31374 = ~n31183 & ~n31373;
  assign n31375 = ~pi74 & ~n31374;
  assign n31376 = n31182 & ~n31375;
  assign n31377 = n4437 & ~n31376;
  assign n31378 = ~n31353 & n31377;
  assign n31379 = n31225 & ~n31378;
  assign n31380 = ~n60206 & ~n31379;
  assign n31381 = n30926 & ~n31380;
  assign n31382 = ~pi954 & ~n31381;
  assign n31383 = ~n31229 & n31382;
  assign n31384 = ~pi33 & ~n31228;
  assign n31385 = pi33 & ~n31380;
  assign n31386 = pi954 & ~n31385;
  assign n31387 = ~n31384 & n31386;
  assign po191 = ~n31383 & ~n31387;
  assign n31389 = n3871 & n5053;
  assign n31390 = n2439 & n28970;
  assign n31391 = n3213 & ~n31390;
  assign n31392 = n2439 & n29017;
  assign n31393 = n28606 & ~n31392;
  assign n31394 = n58992 & ~n31393;
  assign n31395 = ~n31391 & n31394;
  assign n31396 = ~n31389 & ~n31395;
  assign n31397 = pi57 & ~n28295;
  assign n31398 = ~pi55 & ~n28301;
  assign n31399 = ~pi100 & ~n28309;
  assign n31400 = pi95 & ~n2661;
  assign n31401 = ~pi32 & ~n6380;
  assign n31402 = ~pi40 & ~n28318;
  assign n31403 = ~pi91 & n2589;
  assign n31404 = n2530 & n2579;
  assign n31405 = n2614 & n60238;
  assign n31406 = n58800 & n31405;
  assign n31407 = pi96 & n31406;
  assign n31408 = ~pi72 & ~n31407;
  assign n31409 = pi108 & ~n6365;
  assign n31410 = ~pi46 & ~n31409;
  assign n31411 = ~pi86 & pi94;
  assign n31412 = n58834 & n31411;
  assign n31413 = ~pi97 & ~n31412;
  assign n31414 = ~n6335 & ~n28399;
  assign n31415 = pi64 & ~n2519;
  assign n31416 = n2460 & ~n28370;
  assign n31417 = n28354 & ~n31416;
  assign n31418 = ~pi84 & ~n31417;
  assign n31419 = ~n28375 & ~n31418;
  assign n31420 = n28346 & ~n31419;
  assign n31421 = pi111 & ~n28348;
  assign n31422 = ~pi82 & ~n31421;
  assign n31423 = ~n28376 & n31422;
  assign n31424 = ~n31420 & n31423;
  assign n31425 = n6320 & ~n60076;
  assign n31426 = ~n31424 & n31425;
  assign n31427 = pi67 & ~n58781;
  assign n31428 = n2457 & n28348;
  assign n31429 = pi36 & ~n31428;
  assign n31430 = ~n31427 & ~n31429;
  assign n31431 = ~n31426 & n31430;
  assign n31432 = n6324 & ~n31431;
  assign n31433 = n28343 & ~n31432;
  assign n31434 = ~pi71 & ~n60077;
  assign n31435 = ~n31433 & n31434;
  assign n31436 = n28388 & ~n31435;
  assign n31437 = ~pi107 & ~n31436;
  assign n31438 = pi65 & ~pi71;
  assign n31439 = n2469 & n31438;
  assign n31440 = n31437 & ~n31439;
  assign n31441 = pi107 & ~n2486;
  assign n31442 = ~pi63 & ~n31441;
  assign n31443 = ~n31440 & n31442;
  assign n31444 = ~pi64 & ~n31443;
  assign n31445 = ~n31415 & ~n31444;
  assign n31446 = ~pi81 & ~pi102;
  assign n31447 = ~n31445 & n31446;
  assign n31448 = ~n31437 & n31442;
  assign n31449 = pi63 & ~pi107;
  assign n31450 = n2486 & n31449;
  assign n31451 = ~pi64 & ~n31450;
  assign n31452 = ~n31448 & n31451;
  assign n31453 = ~n31415 & ~n31452;
  assign n31454 = n31447 & ~n31453;
  assign n31455 = n31414 & ~n31454;
  assign n31456 = n2470 & ~n31455;
  assign n31457 = pi98 & ~n2559;
  assign n31458 = ~pi77 & ~n31457;
  assign n31459 = ~n6390 & n31458;
  assign n31460 = ~n31456 & n31459;
  assign n31461 = n58832 & n31460;
  assign n31462 = n31413 & ~n31461;
  assign n31463 = ~n28628 & ~n31462;
  assign n31464 = ~pi108 & ~n31463;
  assign n31465 = n31410 & ~n31464;
  assign n31466 = ~pi110 & n28449;
  assign n31467 = ~n31465 & n31466;
  assign n31468 = ~pi109 & n2548;
  assign n31469 = pi110 & ~n31468;
  assign n31470 = ~n28447 & ~n31469;
  assign n31471 = ~n31467 & n31470;
  assign n31472 = ~pi47 & ~n31471;
  assign n31473 = n6362 & ~n31472;
  assign n31474 = n29720 & ~n31473;
  assign n31475 = ~n28325 & ~n31474;
  assign n31476 = ~pi93 & ~n31475;
  assign n31477 = ~n2528 & ~n31476;
  assign n31478 = ~pi35 & ~n31477;
  assign n31479 = pi35 & ~n58807;
  assign n31480 = ~pi70 & ~n31479;
  assign n31481 = ~n31478 & n31480;
  assign n31482 = ~pi51 & ~n31481;
  assign n31483 = n2604 & ~n31482;
  assign n31484 = n31408 & ~n31483;
  assign n31485 = n31402 & ~n31484;
  assign n31486 = n31401 & ~n31485;
  assign n31487 = n2597 & n28317;
  assign n31488 = pi32 & ~n31487;
  assign n31489 = n60122 & ~n31488;
  assign n31490 = ~pi93 & n28322;
  assign n31491 = ~pi35 & ~pi40;
  assign n31492 = ~pi40 & n58823;
  assign n31493 = ~pi35 & n58820;
  assign n31494 = n58817 & n31491;
  assign n31495 = n31490 & n60239;
  assign n31496 = pi32 & ~n31495;
  assign n31497 = ~n60122 & ~n31496;
  assign n31498 = ~n31489 & ~n31497;
  assign n31499 = ~n31486 & ~n31498;
  assign n31500 = ~pi95 & ~n31499;
  assign n31501 = ~n31400 & ~n31500;
  assign n31502 = ~pi39 & ~n31501;
  assign n31503 = pi1093 & ~n2793;
  assign n31504 = pi824 & ~pi1091;
  assign n31505 = n31503 & ~n31504;
  assign n31506 = pi829 & ~n31503;
  assign n31507 = ~pi824 & ~n31506;
  assign n31508 = ~n6416 & ~n31507;
  assign n31509 = ~n2442 & ~n31505;
  assign n31510 = n29535 & n60240;
  assign n31511 = n2783 & n31510;
  assign n31512 = ~n2680 & ~n31510;
  assign n31513 = ~n2782 & ~n31512;
  assign n31514 = n58822 & ~n31513;
  assign n31515 = ~n2782 & n29911;
  assign n31516 = ~n31514 & ~n31515;
  assign n31517 = n58822 & ~n31511;
  assign n31518 = n58846 & ~n60241;
  assign n31519 = ~n2822 & n31510;
  assign n31520 = n58822 & ~n31519;
  assign n31521 = ~n58846 & n31520;
  assign n31522 = pi215 & ~n31521;
  assign n31523 = ~n31518 & n31522;
  assign n31524 = n29534 & n30682;
  assign n31525 = pi221 & n29534;
  assign n31526 = n30818 & n31525;
  assign n31527 = ~n2845 & n31524;
  assign n31528 = n58822 & ~n60242;
  assign n31529 = ~pi215 & ~n31528;
  assign n31530 = pi299 & ~n31529;
  assign n31531 = n58846 & n60241;
  assign n31532 = ~n58846 & ~n31520;
  assign n31533 = pi215 & ~n31532;
  assign n31534 = ~n31531 & n31533;
  assign n31535 = ~pi215 & ~n60242;
  assign n31536 = n58822 & n31535;
  assign n31537 = ~n31534 & ~n31536;
  assign n31538 = pi299 & ~n31537;
  assign n31539 = ~n31523 & n31530;
  assign n31540 = n2790 & ~n60241;
  assign n31541 = ~n2790 & n31520;
  assign n31542 = pi223 & ~n31541;
  assign n31543 = ~n31540 & n31542;
  assign n31544 = n29534 & n30674;
  assign n31545 = pi224 & n29534;
  assign n31546 = n28534 & n31545;
  assign n31547 = ~n2792 & n31544;
  assign n31548 = n58822 & ~n60244;
  assign n31549 = ~pi223 & ~n31548;
  assign n31550 = ~pi299 & ~n31549;
  assign n31551 = ~n31543 & n31550;
  assign n31552 = pi39 & ~n31551;
  assign n31553 = pi39 & ~n60243;
  assign n31554 = ~n31551 & n31553;
  assign n31555 = ~n60243 & n31552;
  assign n31556 = ~n31502 & ~n60245;
  assign n31557 = ~pi38 & ~n31556;
  assign n31558 = n31399 & ~n31557;
  assign n31559 = n28578 & ~n31558;
  assign n31560 = pi87 & ~n60071;
  assign n31561 = ~pi75 & ~n31560;
  assign n31562 = n2438 & n31561;
  assign n31563 = ~n31559 & n31562;
  assign n31564 = ~pi74 & ~n31563;
  assign n31565 = n31398 & ~n31564;
  assign n31566 = ~pi56 & ~n31565;
  assign n31567 = ~pi55 & ~pi74;
  assign n31568 = n28300 & n31567;
  assign n31569 = n28283 & n60071;
  assign n31570 = pi56 & ~n60246;
  assign n31571 = ~n31566 & ~n31570;
  assign n31572 = ~pi62 & ~n31571;
  assign n31573 = ~pi56 & n28283;
  assign n31574 = n60071 & n31573;
  assign n31575 = pi62 & ~n31574;
  assign n31576 = ~pi59 & ~n31575;
  assign n31577 = ~n31572 & n31576;
  assign n31578 = ~pi57 & ~n31577;
  assign po167 = ~n31397 & ~n31578;
  assign n31580 = ~pi228 & ~n4441;
  assign n31581 = pi57 & ~n31580;
  assign n31582 = ~n2680 & ~n2781;
  assign n31583 = ~pi907 & n2680;
  assign n31584 = ~n31582 & ~n31583;
  assign n31585 = pi30 & pi228;
  assign n31586 = ~pi228 & n58822;
  assign n31587 = n2634 & n31586;
  assign n31588 = ~pi100 & n31586;
  assign n31589 = n30890 & n31588;
  assign n31590 = n6305 & n31587;
  assign n31591 = n6308 & n60247;
  assign n31592 = n58815 & n28299;
  assign n31593 = ~pi54 & n6307;
  assign n31594 = n60247 & n31593;
  assign n31595 = n31586 & n31592;
  assign n31596 = ~pi74 & n60249;
  assign n31597 = ~pi228 & n60090;
  assign n31598 = ~n31585 & ~n31586;
  assign n31599 = ~pi228 & ~n28288;
  assign n31600 = ~n31598 & ~n31599;
  assign n31601 = ~n31585 & ~n60248;
  assign n31602 = n31584 & n60250;
  assign n31603 = n31581 & n31602;
  assign n31604 = ~pi602 & n2680;
  assign n31605 = ~n31582 & ~n31604;
  assign n31606 = ~pi228 & ~n28467;
  assign n31607 = ~n31585 & ~n31606;
  assign n31608 = n31605 & ~n31607;
  assign n31609 = ~pi299 & ~n31608;
  assign n31610 = ~pi299 & n28312;
  assign n31611 = ~n31609 & ~n31610;
  assign n31612 = n31585 & n31605;
  assign n31613 = ~n28445 & ~n28469;
  assign n31614 = ~pi228 & n31605;
  assign n31615 = ~n31613 & n31614;
  assign n31616 = ~n31612 & ~n31615;
  assign n31617 = n28312 & ~n31616;
  assign n31618 = ~n31611 & ~n31617;
  assign n31619 = n31584 & n31585;
  assign n31620 = pi299 & ~n31619;
  assign n31621 = n28473 & n28482;
  assign n31622 = ~n28476 & ~n28481;
  assign n31623 = n31584 & ~n31622;
  assign n31624 = n31621 & ~n31623;
  assign n31625 = ~n28478 & n31584;
  assign n31626 = ~n31621 & ~n31625;
  assign n31627 = ~pi228 & ~n31626;
  assign n31628 = ~n31624 & n31627;
  assign n31629 = n31620 & ~n31628;
  assign n31630 = pi232 & ~n31629;
  assign n31631 = pi232 & ~n31618;
  assign n31632 = ~n31629 & n31631;
  assign n31633 = ~n31618 & n31630;
  assign n31634 = ~pi228 & n31625;
  assign n31635 = n31620 & ~n31634;
  assign n31636 = ~pi232 & ~n31635;
  assign n31637 = ~n31609 & n31636;
  assign n31638 = ~n60251 & ~n31637;
  assign n31639 = ~pi39 & ~n31638;
  assign n31640 = ~pi228 & ~n60082;
  assign n31641 = ~n31585 & ~n31640;
  assign n31642 = n2852 & ~n31641;
  assign n31643 = ~n31585 & ~n31642;
  assign n31644 = n31584 & ~n31643;
  assign n31645 = pi299 & ~n31644;
  assign n31646 = ~pi228 & n60085;
  assign n31647 = ~n31585 & ~n31646;
  assign n31648 = n31605 & ~n31647;
  assign n31649 = ~pi299 & ~n31648;
  assign n31650 = pi39 & ~n31649;
  assign n31651 = ~n31645 & n31650;
  assign n31652 = ~pi38 & ~n31651;
  assign n31653 = ~n31639 & n31652;
  assign n31654 = pi299 & n31584;
  assign n31655 = ~pi299 & n31605;
  assign n31656 = ~n31654 & ~n31655;
  assign n31657 = ~pi39 & ~n31598;
  assign n31658 = ~n31656 & n31657;
  assign n31659 = n31585 & ~n31656;
  assign n31660 = pi38 & ~n31659;
  assign n31661 = ~n31658 & n31660;
  assign n31662 = ~n31653 & ~n31661;
  assign n31663 = ~pi100 & ~n31662;
  assign n31664 = n58822 & ~n28564;
  assign n31665 = pi683 & ~n2707;
  assign n31666 = n31664 & n31665;
  assign n31667 = ~n31582 & n31666;
  assign n31668 = n28551 & n31667;
  assign n31669 = pi252 & n29911;
  assign n31670 = ~n2781 & ~n31669;
  assign n31671 = ~n58825 & n2781;
  assign n31672 = ~n2781 & n31669;
  assign n31673 = n58825 & n2781;
  assign n31674 = ~n31672 & ~n31673;
  assign n31675 = ~n31670 & ~n31671;
  assign n31676 = pi252 & ~n28551;
  assign n31677 = ~n60252 & n31676;
  assign n31678 = ~n31668 & ~n31677;
  assign n31679 = ~pi228 & ~n31604;
  assign n31680 = ~n31678 & n31679;
  assign n31681 = ~pi299 & ~n31612;
  assign n31682 = ~n31680 & n31681;
  assign n31683 = ~n28553 & n60252;
  assign n31684 = n28553 & ~n31667;
  assign n31685 = ~pi228 & ~n31583;
  assign n31686 = ~n31684 & n31685;
  assign n31687 = ~n31683 & n31686;
  assign n31688 = n31620 & ~n31687;
  assign n31689 = n2634 & ~n31688;
  assign n31690 = ~n31682 & n31689;
  assign n31691 = ~n2634 & n31659;
  assign n31692 = pi100 & ~n31691;
  assign n31693 = ~n31690 & n31692;
  assign n31694 = ~pi87 & ~n31693;
  assign n31695 = ~n31663 & n31694;
  assign n31696 = pi87 & n31659;
  assign n31697 = ~pi75 & ~n31696;
  assign n31698 = ~n31695 & n31697;
  assign n31699 = ~n2672 & n31659;
  assign n31700 = n59291 & n31658;
  assign n31701 = ~n31699 & ~n31700;
  assign n31702 = pi75 & n31701;
  assign n31703 = ~pi92 & ~n31702;
  assign n31704 = ~n31698 & n31703;
  assign n31705 = ~pi75 & n31701;
  assign n31706 = pi75 & ~n31659;
  assign n31707 = pi92 & ~n31706;
  assign n31708 = ~n31705 & n31707;
  assign n31709 = ~pi54 & ~n31708;
  assign n31710 = ~n31704 & n31709;
  assign n31711 = n6307 & n31701;
  assign n31712 = ~n6307 & ~n31659;
  assign n31713 = ~n31711 & ~n31712;
  assign n31714 = pi54 & ~n31713;
  assign n31715 = ~pi74 & ~n31714;
  assign n31716 = ~n31710 & n31715;
  assign n31717 = ~pi54 & n31711;
  assign n31718 = ~n31593 & ~n31659;
  assign n31719 = pi74 & ~n31718;
  assign n31720 = ~n31717 & n31719;
  assign n31721 = ~pi55 & ~n31720;
  assign n31722 = ~n31716 & n31721;
  assign n31723 = pi55 & ~n31602;
  assign n31724 = n4437 & ~n31723;
  assign n31725 = ~n31722 & n31724;
  assign n31726 = ~n4437 & n31619;
  assign n31727 = ~pi59 & ~n31726;
  assign n31728 = ~n31725 & n31727;
  assign n31729 = ~pi228 & ~n4440;
  assign n31730 = n31602 & ~n31729;
  assign n31731 = pi59 & ~n31730;
  assign n31732 = ~pi57 & ~n31731;
  assign n31733 = ~n31728 & n31732;
  assign po171 = ~n31603 & ~n31733;
  assign n31735 = ~pi947 & n2680;
  assign n31736 = ~n2821 & ~n31735;
  assign n31737 = n60250 & n31736;
  assign n31738 = n31581 & n31737;
  assign n31739 = ~pi587 & n2680;
  assign n31740 = ~n2821 & ~n31739;
  assign n31741 = n31585 & n31740;
  assign n31742 = ~pi228 & n31740;
  assign n31743 = ~n31613 & n31742;
  assign n31744 = ~n31741 & ~n31743;
  assign n31745 = n28312 & ~n31744;
  assign n31746 = ~n31607 & n31740;
  assign n31747 = ~n28312 & n31746;
  assign n31748 = ~pi299 & ~n31747;
  assign n31749 = ~n31745 & n31748;
  assign n31750 = n31585 & n31736;
  assign n31751 = pi299 & ~n31750;
  assign n31752 = ~n31622 & n31736;
  assign n31753 = n31621 & ~n31752;
  assign n31754 = ~n28478 & n31736;
  assign n31755 = ~n31621 & ~n31754;
  assign n31756 = ~pi228 & ~n31755;
  assign n31757 = ~n31753 & n31756;
  assign n31758 = n31751 & ~n31757;
  assign n31759 = pi232 & ~n31758;
  assign n31760 = pi232 & ~n31749;
  assign n31761 = ~n31758 & n31760;
  assign n31762 = ~n31749 & n31759;
  assign n31763 = ~pi299 & ~n31746;
  assign n31764 = ~pi228 & n31754;
  assign n31765 = n31751 & ~n31764;
  assign n31766 = ~pi232 & ~n31765;
  assign n31767 = ~n31763 & n31766;
  assign n31768 = ~n60253 & ~n31767;
  assign n31769 = ~pi39 & ~n31768;
  assign n31770 = ~n2853 & ~n31751;
  assign n31771 = n31642 & n31736;
  assign n31772 = ~n31770 & ~n31771;
  assign n31773 = ~n31647 & n31740;
  assign n31774 = ~pi299 & ~n31773;
  assign n31775 = pi39 & ~n31774;
  assign n31776 = pi39 & ~n31772;
  assign n31777 = ~n31774 & n31776;
  assign n31778 = ~n31772 & n31775;
  assign n31779 = ~pi38 & ~n60254;
  assign n31780 = ~n31769 & n31779;
  assign n31781 = pi299 & ~n31736;
  assign n31782 = ~pi299 & ~n31740;
  assign n31783 = ~n31781 & ~n31782;
  assign n31784 = n31657 & n31783;
  assign n31785 = n31585 & n31783;
  assign n31786 = pi38 & ~n31785;
  assign n31787 = ~n31784 & n31786;
  assign n31788 = ~n31780 & ~n31787;
  assign n31789 = ~pi100 & ~n31788;
  assign n31790 = ~pi228 & n2674;
  assign n31791 = ~n2778 & n31669;
  assign n31792 = n58825 & n2778;
  assign n31793 = ~n58825 & n2778;
  assign n31794 = ~n2778 & ~n31669;
  assign n31795 = ~n31793 & ~n31794;
  assign n31796 = ~n31791 & ~n31792;
  assign n31797 = ~n31739 & n60255;
  assign n31798 = n31790 & ~n31797;
  assign n31799 = pi142 & ~n60255;
  assign n31800 = ~n2821 & n31666;
  assign n31801 = ~pi142 & ~n31800;
  assign n31802 = ~n2680 & n2778;
  assign n31803 = ~pi587 & ~n31802;
  assign n31804 = ~pi228 & ~n31803;
  assign n31805 = ~n31801 & n31804;
  assign n31806 = ~n31799 & n31805;
  assign n31807 = ~n31741 & ~n31790;
  assign n31808 = ~n31806 & n31807;
  assign n31809 = ~n31798 & ~n31808;
  assign n31810 = ~pi299 & ~n31809;
  assign n31811 = n28553 & ~n31735;
  assign n31812 = n31800 & n31811;
  assign n31813 = ~pi947 & ~n31802;
  assign n31814 = ~n28553 & ~n31813;
  assign n31815 = n60255 & n31814;
  assign n31816 = ~n31812 & ~n31815;
  assign n31817 = ~pi228 & ~n31816;
  assign n31818 = n31751 & ~n31817;
  assign n31819 = n2634 & ~n31818;
  assign n31820 = ~n31810 & n31819;
  assign n31821 = ~n2634 & n31785;
  assign n31822 = pi100 & ~n31821;
  assign n31823 = ~n31820 & n31822;
  assign n31824 = ~pi87 & ~n31823;
  assign n31825 = ~n31789 & n31824;
  assign n31826 = pi87 & n31785;
  assign n31827 = ~pi75 & ~n31826;
  assign n31828 = ~n31825 & n31827;
  assign n31829 = ~n2672 & n31785;
  assign n31830 = n59291 & n31784;
  assign n31831 = ~n31829 & ~n31830;
  assign n31832 = pi75 & n31831;
  assign n31833 = ~pi92 & ~n31832;
  assign n31834 = ~n31828 & n31833;
  assign n31835 = ~pi75 & n31831;
  assign n31836 = pi75 & ~n31785;
  assign n31837 = pi92 & ~n31836;
  assign n31838 = ~n31835 & n31837;
  assign n31839 = ~pi54 & ~n31838;
  assign n31840 = ~n31834 & n31839;
  assign n31841 = n6307 & n31831;
  assign n31842 = ~n6307 & ~n31785;
  assign n31843 = ~n31841 & ~n31842;
  assign n31844 = pi54 & ~n31843;
  assign n31845 = ~pi74 & ~n31844;
  assign n31846 = ~n31840 & n31845;
  assign n31847 = ~pi54 & n31841;
  assign n31848 = ~n31593 & ~n31785;
  assign n31849 = pi74 & ~n31848;
  assign n31850 = ~n31847 & n31849;
  assign n31851 = ~pi55 & ~n31850;
  assign n31852 = ~n31846 & n31851;
  assign n31853 = pi55 & ~n31737;
  assign n31854 = n4437 & ~n31853;
  assign n31855 = ~n31852 & n31854;
  assign n31856 = ~n4437 & n31750;
  assign n31857 = ~pi59 & ~n31856;
  assign n31858 = ~n31855 & n31857;
  assign n31859 = ~n31729 & n31737;
  assign n31860 = pi59 & ~n31859;
  assign n31861 = ~pi57 & ~n31860;
  assign n31862 = ~n31858 & n31861;
  assign po172 = ~n31738 & ~n31862;
  assign n31864 = pi30 & n2680;
  assign n31865 = pi228 & n31864;
  assign n31866 = pi970 & n31865;
  assign n31867 = ~pi228 & pi970;
  assign n31868 = n29911 & n31867;
  assign n31869 = n28288 & n31868;
  assign n31870 = n4441 & n31869;
  assign n31871 = ~n31866 & ~n31870;
  assign n31872 = pi57 & ~n31871;
  assign n31873 = pi299 & ~n31866;
  assign n31874 = n2680 & ~n28478;
  assign n31875 = n31867 & n31874;
  assign n31876 = n31873 & ~n31875;
  assign n31877 = ~n28483 & ~n31876;
  assign n31878 = n2680 & n28480;
  assign n31879 = n31867 & n31878;
  assign n31880 = ~n31866 & ~n31879;
  assign n31881 = n28482 & ~n31880;
  assign n31882 = ~n31877 & ~n31881;
  assign n31883 = n2680 & ~n31607;
  assign n31884 = ~n28312 & ~n31883;
  assign n31885 = ~pi228 & n28445;
  assign n31886 = ~n28468 & ~n31865;
  assign n31887 = ~n31885 & n31886;
  assign n31888 = ~n31884 & ~n31887;
  assign n31889 = pi967 & n31888;
  assign n31890 = ~pi299 & ~n31889;
  assign n31891 = pi232 & ~n31890;
  assign n31892 = ~n31882 & n31891;
  assign n31893 = pi967 & n31883;
  assign n31894 = ~pi299 & ~n31893;
  assign n31895 = ~pi232 & ~n31876;
  assign n31896 = ~n31894 & n31895;
  assign n31897 = ~n31892 & ~n31896;
  assign n31898 = ~pi39 & ~n31897;
  assign n31899 = pi299 & pi970;
  assign n31900 = n2680 & n28523;
  assign n31901 = ~pi228 & ~n31900;
  assign n31902 = n31899 & ~n31901;
  assign n31903 = ~pi299 & pi967;
  assign n31904 = n2680 & n60085;
  assign n31905 = ~pi228 & ~n31904;
  assign n31906 = n31903 & ~n31905;
  assign n31907 = ~n31902 & ~n31906;
  assign n31908 = pi228 & ~n31864;
  assign n31909 = pi39 & ~n31908;
  assign n31910 = ~n31907 & n31909;
  assign n31911 = ~pi38 & ~n31910;
  assign n31912 = ~n31898 & n31911;
  assign n31913 = ~pi228 & ~n29911;
  assign n31914 = ~n31908 & ~n31913;
  assign n31915 = n2680 & ~n31598;
  assign n31916 = pi967 & n60256;
  assign n31917 = ~pi299 & ~n31916;
  assign n31918 = ~n31868 & n31873;
  assign n31919 = ~pi39 & ~n31918;
  assign n31920 = ~n31917 & n31919;
  assign n31921 = ~n31899 & ~n31903;
  assign n31922 = n31865 & ~n31921;
  assign n31923 = pi39 & n31922;
  assign n31924 = pi38 & ~n31923;
  assign n31925 = ~n31920 & n31924;
  assign n31926 = ~n31912 & ~n31925;
  assign n31927 = ~pi100 & ~n31926;
  assign n31928 = n2680 & n31666;
  assign n31929 = n28551 & n31928;
  assign n31930 = ~n28551 & n31669;
  assign n31931 = ~pi228 & ~n31930;
  assign n31932 = ~pi228 & ~n31929;
  assign n31933 = ~n31930 & n31932;
  assign n31934 = ~n31929 & n31931;
  assign n31935 = ~n31908 & ~n60257;
  assign n31936 = pi967 & n31935;
  assign n31937 = ~pi299 & ~n31936;
  assign n31938 = n28553 & ~n31928;
  assign n31939 = ~n28553 & ~n31669;
  assign n31940 = ~pi228 & ~n31939;
  assign n31941 = ~n31938 & n31940;
  assign n31942 = pi970 & n31941;
  assign n31943 = n31873 & ~n31942;
  assign n31944 = n2634 & ~n31943;
  assign n31945 = ~n31937 & n31944;
  assign n31946 = ~n2634 & n31922;
  assign n31947 = pi100 & ~n31946;
  assign n31948 = ~n31945 & n31947;
  assign n31949 = ~pi87 & ~n31948;
  assign n31950 = ~n31927 & n31949;
  assign n31951 = pi87 & n31922;
  assign n31952 = ~pi75 & ~n31951;
  assign n31953 = ~n31950 & n31952;
  assign n31954 = ~n2672 & n31922;
  assign n31955 = n59291 & n31920;
  assign n31956 = ~n31954 & ~n31955;
  assign n31957 = pi75 & n31956;
  assign n31958 = ~pi92 & ~n31957;
  assign n31959 = ~n31953 & n31958;
  assign n31960 = ~pi75 & n31956;
  assign n31961 = pi75 & ~n31922;
  assign n31962 = pi92 & ~n31961;
  assign n31963 = ~n31960 & n31962;
  assign n31964 = ~pi54 & ~n31963;
  assign n31965 = ~n31959 & n31964;
  assign n31966 = n6307 & n31956;
  assign n31967 = ~n6307 & ~n31922;
  assign n31968 = ~n31966 & ~n31967;
  assign n31969 = pi54 & ~n31968;
  assign n31970 = ~pi74 & ~n31969;
  assign n31971 = ~n31965 & n31970;
  assign n31972 = ~pi54 & n31966;
  assign n31973 = ~n31593 & ~n31922;
  assign n31974 = pi74 & ~n31973;
  assign n31975 = ~n31972 & n31974;
  assign n31976 = ~pi55 & ~n31975;
  assign n31977 = ~n31971 & n31976;
  assign n31978 = pi55 & ~n31866;
  assign n31979 = ~n31869 & n31978;
  assign n31980 = n4437 & ~n31979;
  assign n31981 = ~n31977 & n31980;
  assign n31982 = ~n4437 & n31866;
  assign n31983 = ~pi59 & ~n31982;
  assign n31984 = ~n31981 & n31983;
  assign n31985 = n4440 & n31869;
  assign n31986 = pi59 & ~n31866;
  assign n31987 = ~n31985 & n31986;
  assign n31988 = ~pi57 & ~n31987;
  assign n31989 = ~n31984 & n31988;
  assign po173 = ~n31872 & ~n31989;
  assign n31991 = pi972 & n31865;
  assign n31992 = ~pi228 & pi972;
  assign n31993 = n29911 & n31992;
  assign n31994 = n28288 & n31993;
  assign n31995 = n4441 & n31994;
  assign n31996 = ~n31991 & ~n31995;
  assign n31997 = pi57 & ~n31996;
  assign n31998 = pi299 & ~n31991;
  assign n31999 = n31874 & n31992;
  assign n32000 = n31998 & ~n31999;
  assign n32001 = ~n28483 & ~n32000;
  assign n32002 = n31878 & n31992;
  assign n32003 = ~n31991 & ~n32002;
  assign n32004 = n28482 & ~n32003;
  assign n32005 = ~n32001 & ~n32004;
  assign n32006 = pi961 & n31888;
  assign n32007 = ~pi299 & ~n32006;
  assign n32008 = pi232 & ~n32007;
  assign n32009 = ~n32005 & n32008;
  assign n32010 = pi961 & n31883;
  assign n32011 = ~pi299 & ~n32010;
  assign n32012 = ~pi232 & ~n32000;
  assign n32013 = ~n32011 & n32012;
  assign n32014 = ~n32009 & ~n32013;
  assign n32015 = ~pi39 & ~n32014;
  assign n32016 = ~pi299 & pi961;
  assign n32017 = ~n31905 & n32016;
  assign n32018 = pi299 & pi972;
  assign n32019 = ~n31901 & n32018;
  assign n32020 = ~n32017 & ~n32019;
  assign n32021 = n31909 & ~n32020;
  assign n32022 = ~pi38 & ~n32021;
  assign n32023 = ~n32015 & n32022;
  assign n32024 = pi961 & n60256;
  assign n32025 = ~pi299 & ~n32024;
  assign n32026 = ~n31993 & n31998;
  assign n32027 = ~pi39 & ~n32026;
  assign n32028 = ~n32025 & n32027;
  assign n32029 = ~n32016 & ~n32018;
  assign n32030 = n31865 & ~n32029;
  assign n32031 = pi39 & n32030;
  assign n32032 = pi38 & ~n32031;
  assign n32033 = ~n32028 & n32032;
  assign n32034 = ~n32023 & ~n32033;
  assign n32035 = ~pi100 & ~n32034;
  assign n32036 = pi961 & n31935;
  assign n32037 = ~pi299 & ~n32036;
  assign n32038 = pi972 & n31941;
  assign n32039 = n31998 & ~n32038;
  assign n32040 = n2634 & ~n32039;
  assign n32041 = ~n32037 & n32040;
  assign n32042 = ~n2634 & n32030;
  assign n32043 = pi100 & ~n32042;
  assign n32044 = ~n32041 & n32043;
  assign n32045 = ~pi87 & ~n32044;
  assign n32046 = ~n32035 & n32045;
  assign n32047 = pi87 & n32030;
  assign n32048 = ~pi75 & ~n32047;
  assign n32049 = ~n32046 & n32048;
  assign n32050 = ~n2672 & n32030;
  assign n32051 = n59291 & n32028;
  assign n32052 = ~n32050 & ~n32051;
  assign n32053 = pi75 & n32052;
  assign n32054 = ~pi92 & ~n32053;
  assign n32055 = ~n32049 & n32054;
  assign n32056 = ~pi75 & n32052;
  assign n32057 = pi75 & ~n32030;
  assign n32058 = pi92 & ~n32057;
  assign n32059 = ~n32056 & n32058;
  assign n32060 = ~pi54 & ~n32059;
  assign n32061 = ~n32055 & n32060;
  assign n32062 = n6307 & n32052;
  assign n32063 = ~n6307 & ~n32030;
  assign n32064 = ~n32062 & ~n32063;
  assign n32065 = pi54 & ~n32064;
  assign n32066 = ~pi74 & ~n32065;
  assign n32067 = ~n32061 & n32066;
  assign n32068 = ~pi54 & n32062;
  assign n32069 = ~n31593 & ~n32030;
  assign n32070 = pi74 & ~n32069;
  assign n32071 = ~n32068 & n32070;
  assign n32072 = ~pi55 & ~n32071;
  assign n32073 = ~n32067 & n32072;
  assign n32074 = pi55 & ~n31991;
  assign n32075 = ~n31994 & n32074;
  assign n32076 = n4437 & ~n32075;
  assign n32077 = ~n32073 & n32076;
  assign n32078 = ~n4437 & n31991;
  assign n32079 = ~pi59 & ~n32078;
  assign n32080 = ~n32077 & n32079;
  assign n32081 = n4440 & n31994;
  assign n32082 = pi59 & ~n31991;
  assign n32083 = ~n32081 & n32082;
  assign n32084 = ~pi57 & ~n32083;
  assign n32085 = ~n32080 & n32084;
  assign po174 = ~n31997 & ~n32085;
  assign n32087 = pi960 & n31865;
  assign n32088 = ~pi228 & pi960;
  assign n32089 = n29911 & n32088;
  assign n32090 = n28288 & n32089;
  assign n32091 = n4441 & n32090;
  assign n32092 = ~n32087 & ~n32091;
  assign n32093 = pi57 & ~n32092;
  assign n32094 = pi299 & ~n32087;
  assign n32095 = n31874 & n32088;
  assign n32096 = n32094 & ~n32095;
  assign n32097 = ~n28483 & ~n32096;
  assign n32098 = n31878 & n32088;
  assign n32099 = ~n32087 & ~n32098;
  assign n32100 = n28482 & ~n32099;
  assign n32101 = ~n32097 & ~n32100;
  assign n32102 = pi977 & n31888;
  assign n32103 = ~pi299 & ~n32102;
  assign n32104 = pi232 & ~n32103;
  assign n32105 = ~n32101 & n32104;
  assign n32106 = pi977 & n31883;
  assign n32107 = ~pi299 & ~n32106;
  assign n32108 = ~pi232 & ~n32096;
  assign n32109 = ~n32107 & n32108;
  assign n32110 = ~n32105 & ~n32109;
  assign n32111 = ~pi39 & ~n32110;
  assign n32112 = ~pi299 & pi977;
  assign n32113 = ~n31905 & n32112;
  assign n32114 = pi299 & pi960;
  assign n32115 = ~n31901 & n32114;
  assign n32116 = ~n32113 & ~n32115;
  assign n32117 = n31909 & ~n32116;
  assign n32118 = ~pi38 & ~n32117;
  assign n32119 = ~n32111 & n32118;
  assign n32120 = pi977 & n60256;
  assign n32121 = ~pi299 & ~n32120;
  assign n32122 = ~n32089 & n32094;
  assign n32123 = ~pi39 & ~n32122;
  assign n32124 = ~n32121 & n32123;
  assign n32125 = ~n32112 & ~n32114;
  assign n32126 = n31865 & ~n32125;
  assign n32127 = pi39 & n32126;
  assign n32128 = pi38 & ~n32127;
  assign n32129 = ~n32124 & n32128;
  assign n32130 = ~n32119 & ~n32129;
  assign n32131 = ~pi100 & ~n32130;
  assign n32132 = pi977 & n31935;
  assign n32133 = ~pi299 & ~n32132;
  assign n32134 = pi960 & n31941;
  assign n32135 = n32094 & ~n32134;
  assign n32136 = n2634 & ~n32135;
  assign n32137 = ~n32133 & n32136;
  assign n32138 = ~n2634 & n32126;
  assign n32139 = pi100 & ~n32138;
  assign n32140 = ~n32137 & n32139;
  assign n32141 = ~pi87 & ~n32140;
  assign n32142 = ~n32131 & n32141;
  assign n32143 = pi87 & n32126;
  assign n32144 = ~pi75 & ~n32143;
  assign n32145 = ~n32142 & n32144;
  assign n32146 = ~n2672 & n32126;
  assign n32147 = n59291 & n32124;
  assign n32148 = ~n32146 & ~n32147;
  assign n32149 = pi75 & n32148;
  assign n32150 = ~pi92 & ~n32149;
  assign n32151 = ~n32145 & n32150;
  assign n32152 = ~pi75 & n32148;
  assign n32153 = pi75 & ~n32126;
  assign n32154 = pi92 & ~n32153;
  assign n32155 = ~n32152 & n32154;
  assign n32156 = ~pi54 & ~n32155;
  assign n32157 = ~n32151 & n32156;
  assign n32158 = n6307 & n32148;
  assign n32159 = ~n6307 & ~n32126;
  assign n32160 = ~n32158 & ~n32159;
  assign n32161 = pi54 & ~n32160;
  assign n32162 = ~pi74 & ~n32161;
  assign n32163 = ~n32157 & n32162;
  assign n32164 = ~pi54 & n32158;
  assign n32165 = ~n31593 & ~n32126;
  assign n32166 = pi74 & ~n32165;
  assign n32167 = ~n32164 & n32166;
  assign n32168 = ~pi55 & ~n32167;
  assign n32169 = ~n32163 & n32168;
  assign n32170 = pi55 & ~n32087;
  assign n32171 = ~n32090 & n32170;
  assign n32172 = n4437 & ~n32171;
  assign n32173 = ~n32169 & n32172;
  assign n32174 = ~n4437 & n32087;
  assign n32175 = ~pi59 & ~n32174;
  assign n32176 = ~n32173 & n32175;
  assign n32177 = n4440 & n32090;
  assign n32178 = pi59 & ~n32087;
  assign n32179 = ~n32177 & n32178;
  assign n32180 = ~pi57 & ~n32179;
  assign n32181 = ~n32176 & n32180;
  assign po175 = ~n32093 & ~n32181;
  assign n32183 = pi963 & n31865;
  assign n32184 = ~pi228 & pi963;
  assign n32185 = n29911 & n32184;
  assign n32186 = n28288 & n32185;
  assign n32187 = n4441 & n32186;
  assign n32188 = ~n32183 & ~n32187;
  assign n32189 = pi57 & ~n32188;
  assign n32190 = pi299 & ~n32183;
  assign n32191 = n31874 & n32184;
  assign n32192 = n32190 & ~n32191;
  assign n32193 = ~n28483 & ~n32192;
  assign n32194 = n31878 & n32184;
  assign n32195 = ~n32183 & ~n32194;
  assign n32196 = n28482 & ~n32195;
  assign n32197 = ~n32193 & ~n32196;
  assign n32198 = pi969 & n31888;
  assign n32199 = ~pi299 & ~n32198;
  assign n32200 = pi232 & ~n32199;
  assign n32201 = ~n32197 & n32200;
  assign n32202 = pi969 & n31883;
  assign n32203 = ~pi299 & ~n32202;
  assign n32204 = ~pi232 & ~n32192;
  assign n32205 = ~n32203 & n32204;
  assign n32206 = ~n32201 & ~n32205;
  assign n32207 = ~pi39 & ~n32206;
  assign n32208 = ~pi299 & pi969;
  assign n32209 = ~n31905 & n32208;
  assign n32210 = pi299 & pi963;
  assign n32211 = ~n31901 & n32210;
  assign n32212 = ~n32209 & ~n32211;
  assign n32213 = n31909 & ~n32212;
  assign n32214 = ~pi38 & ~n32213;
  assign n32215 = ~n32207 & n32214;
  assign n32216 = pi969 & n60256;
  assign n32217 = ~pi299 & ~n32216;
  assign n32218 = ~n32185 & n32190;
  assign n32219 = ~pi39 & ~n32218;
  assign n32220 = ~n32217 & n32219;
  assign n32221 = ~n32208 & ~n32210;
  assign n32222 = n31865 & ~n32221;
  assign n32223 = pi39 & n32222;
  assign n32224 = pi38 & ~n32223;
  assign n32225 = ~n32220 & n32224;
  assign n32226 = ~n32215 & ~n32225;
  assign n32227 = ~pi100 & ~n32226;
  assign n32228 = pi969 & n31935;
  assign n32229 = ~pi299 & ~n32228;
  assign n32230 = pi963 & n31941;
  assign n32231 = n32190 & ~n32230;
  assign n32232 = n2634 & ~n32231;
  assign n32233 = ~n32229 & n32232;
  assign n32234 = ~n2634 & n32222;
  assign n32235 = pi100 & ~n32234;
  assign n32236 = ~n32233 & n32235;
  assign n32237 = ~pi87 & ~n32236;
  assign n32238 = ~n32227 & n32237;
  assign n32239 = pi87 & n32222;
  assign n32240 = ~pi75 & ~n32239;
  assign n32241 = ~n32238 & n32240;
  assign n32242 = ~n2672 & n32222;
  assign n32243 = n59291 & n32220;
  assign n32244 = ~n32242 & ~n32243;
  assign n32245 = pi75 & n32244;
  assign n32246 = ~pi92 & ~n32245;
  assign n32247 = ~n32241 & n32246;
  assign n32248 = ~pi75 & n32244;
  assign n32249 = pi75 & ~n32222;
  assign n32250 = pi92 & ~n32249;
  assign n32251 = ~n32248 & n32250;
  assign n32252 = ~pi54 & ~n32251;
  assign n32253 = ~n32247 & n32252;
  assign n32254 = n6307 & n32244;
  assign n32255 = ~n6307 & ~n32222;
  assign n32256 = ~n32254 & ~n32255;
  assign n32257 = pi54 & ~n32256;
  assign n32258 = ~pi74 & ~n32257;
  assign n32259 = ~n32253 & n32258;
  assign n32260 = ~pi54 & n32254;
  assign n32261 = ~n31593 & ~n32222;
  assign n32262 = pi74 & ~n32261;
  assign n32263 = ~n32260 & n32262;
  assign n32264 = ~pi55 & ~n32263;
  assign n32265 = ~n32259 & n32264;
  assign n32266 = pi55 & ~n32183;
  assign n32267 = ~n32186 & n32266;
  assign n32268 = n4437 & ~n32267;
  assign n32269 = ~n32265 & n32268;
  assign n32270 = ~n4437 & n32183;
  assign n32271 = ~pi59 & ~n32270;
  assign n32272 = ~n32269 & n32271;
  assign n32273 = n4440 & n32186;
  assign n32274 = pi59 & ~n32183;
  assign n32275 = ~n32273 & n32274;
  assign n32276 = ~pi57 & ~n32275;
  assign n32277 = ~n32272 & n32276;
  assign po176 = ~n32189 & ~n32277;
  assign n32279 = pi975 & n31865;
  assign n32280 = ~pi228 & pi975;
  assign n32281 = n29911 & n32280;
  assign n32282 = n28288 & n32281;
  assign n32283 = n4441 & n32282;
  assign n32284 = ~n32279 & ~n32283;
  assign n32285 = pi57 & ~n32284;
  assign n32286 = pi299 & ~n32279;
  assign n32287 = n31874 & n32280;
  assign n32288 = n32286 & ~n32287;
  assign n32289 = ~n28483 & ~n32288;
  assign n32290 = n31878 & n32280;
  assign n32291 = ~n32279 & ~n32290;
  assign n32292 = n28482 & ~n32291;
  assign n32293 = ~n32289 & ~n32292;
  assign n32294 = pi971 & n31888;
  assign n32295 = ~pi299 & ~n32294;
  assign n32296 = pi232 & ~n32295;
  assign n32297 = ~n32293 & n32296;
  assign n32298 = pi971 & n31883;
  assign n32299 = ~pi299 & ~n32298;
  assign n32300 = ~pi232 & ~n32288;
  assign n32301 = ~n32299 & n32300;
  assign n32302 = ~n32297 & ~n32301;
  assign n32303 = ~pi39 & ~n32302;
  assign n32304 = ~pi299 & pi971;
  assign n32305 = ~n31905 & n32304;
  assign n32306 = pi299 & pi975;
  assign n32307 = ~n31901 & n32306;
  assign n32308 = ~n32305 & ~n32307;
  assign n32309 = n31909 & ~n32308;
  assign n32310 = ~pi38 & ~n32309;
  assign n32311 = ~n32303 & n32310;
  assign n32312 = pi971 & n60256;
  assign n32313 = ~pi299 & ~n32312;
  assign n32314 = ~n32281 & n32286;
  assign n32315 = ~pi39 & ~n32314;
  assign n32316 = ~n32313 & n32315;
  assign n32317 = ~n32304 & ~n32306;
  assign n32318 = n31865 & ~n32317;
  assign n32319 = pi39 & n32318;
  assign n32320 = pi38 & ~n32319;
  assign n32321 = ~n32316 & n32320;
  assign n32322 = ~n32311 & ~n32321;
  assign n32323 = ~pi100 & ~n32322;
  assign n32324 = pi971 & n31935;
  assign n32325 = ~pi299 & ~n32324;
  assign n32326 = pi975 & n31941;
  assign n32327 = n32286 & ~n32326;
  assign n32328 = n2634 & ~n32327;
  assign n32329 = ~n32325 & n32328;
  assign n32330 = ~n2634 & n32318;
  assign n32331 = pi100 & ~n32330;
  assign n32332 = ~n32329 & n32331;
  assign n32333 = ~pi87 & ~n32332;
  assign n32334 = ~n32323 & n32333;
  assign n32335 = pi87 & n32318;
  assign n32336 = ~pi75 & ~n32335;
  assign n32337 = ~n32334 & n32336;
  assign n32338 = ~n2672 & n32318;
  assign n32339 = n59291 & n32316;
  assign n32340 = ~n32338 & ~n32339;
  assign n32341 = pi75 & n32340;
  assign n32342 = ~pi92 & ~n32341;
  assign n32343 = ~n32337 & n32342;
  assign n32344 = ~pi75 & n32340;
  assign n32345 = pi75 & ~n32318;
  assign n32346 = pi92 & ~n32345;
  assign n32347 = ~n32344 & n32346;
  assign n32348 = ~pi54 & ~n32347;
  assign n32349 = ~n32343 & n32348;
  assign n32350 = n6307 & n32340;
  assign n32351 = ~n6307 & ~n32318;
  assign n32352 = ~n32350 & ~n32351;
  assign n32353 = pi54 & ~n32352;
  assign n32354 = ~pi74 & ~n32353;
  assign n32355 = ~n32349 & n32354;
  assign n32356 = ~pi54 & n32350;
  assign n32357 = ~n31593 & ~n32318;
  assign n32358 = pi74 & ~n32357;
  assign n32359 = ~n32356 & n32358;
  assign n32360 = ~pi55 & ~n32359;
  assign n32361 = ~n32355 & n32360;
  assign n32362 = pi55 & ~n32279;
  assign n32363 = ~n32282 & n32362;
  assign n32364 = n4437 & ~n32363;
  assign n32365 = ~n32361 & n32364;
  assign n32366 = ~n4437 & n32279;
  assign n32367 = ~pi59 & ~n32366;
  assign n32368 = ~n32365 & n32367;
  assign n32369 = n4440 & n32282;
  assign n32370 = pi59 & ~n32279;
  assign n32371 = ~n32369 & n32370;
  assign n32372 = ~pi57 & ~n32371;
  assign n32373 = ~n32368 & n32372;
  assign po177 = ~n32285 & ~n32373;
  assign n32375 = pi978 & n31865;
  assign n32376 = ~pi228 & pi978;
  assign n32377 = n2680 & n32376;
  assign n32378 = n28288 & n32376;
  assign n32379 = n29911 & n32378;
  assign n32380 = n60090 & n32377;
  assign n32381 = n4441 & n60258;
  assign n32382 = ~n32375 & ~n32381;
  assign n32383 = pi57 & ~n32382;
  assign n32384 = ~pi299 & pi974;
  assign n32385 = pi299 & pi978;
  assign n32386 = ~n32384 & ~n32385;
  assign n32387 = n60256 & ~n32386;
  assign n32388 = ~pi39 & n32387;
  assign n32389 = n31865 & ~n32386;
  assign n32390 = pi39 & n32389;
  assign n32391 = pi38 & ~n32390;
  assign n32392 = ~n32388 & n32391;
  assign n32393 = pi299 & ~n32375;
  assign n32394 = n31874 & n32376;
  assign n32395 = n32393 & ~n32394;
  assign n32396 = ~n28483 & ~n32395;
  assign n32397 = n31878 & n32376;
  assign n32398 = ~n32375 & ~n32397;
  assign n32399 = n28482 & ~n32398;
  assign n32400 = ~n32396 & ~n32399;
  assign n32401 = pi974 & n31888;
  assign n32402 = ~pi299 & ~n32401;
  assign n32403 = pi232 & ~n32402;
  assign n32404 = ~n32400 & n32403;
  assign n32405 = pi974 & n31883;
  assign n32406 = ~pi299 & ~n32405;
  assign n32407 = ~pi232 & ~n32395;
  assign n32408 = ~n32406 & n32407;
  assign n32409 = ~n32404 & ~n32408;
  assign n32410 = ~pi39 & ~n32409;
  assign n32411 = ~n31905 & n32384;
  assign n32412 = ~n31901 & n32385;
  assign n32413 = ~n32411 & ~n32412;
  assign n32414 = n31909 & ~n32413;
  assign n32415 = ~pi38 & ~n32414;
  assign n32416 = ~n32410 & n32415;
  assign n32417 = ~n32392 & ~n32416;
  assign n32418 = ~pi100 & ~n32417;
  assign n32419 = pi974 & n31935;
  assign n32420 = ~pi299 & ~n32419;
  assign n32421 = pi978 & n31941;
  assign n32422 = n32393 & ~n32421;
  assign n32423 = n2634 & ~n32422;
  assign n32424 = ~n32420 & n32423;
  assign n32425 = ~n2634 & n32389;
  assign n32426 = pi100 & ~n32425;
  assign n32427 = ~n32424 & n32426;
  assign n32428 = ~pi87 & ~n32427;
  assign n32429 = ~n32418 & n32428;
  assign n32430 = pi87 & n32389;
  assign n32431 = ~pi75 & ~n32430;
  assign n32432 = ~n32429 & n32431;
  assign n32433 = ~pi228 & ~n2672;
  assign n32434 = n32387 & ~n32433;
  assign n32435 = pi75 & ~n32434;
  assign n32436 = ~pi92 & ~n32435;
  assign n32437 = ~n32432 & n32436;
  assign n32438 = ~pi75 & ~n32434;
  assign n32439 = pi75 & ~n32389;
  assign n32440 = pi92 & ~n32439;
  assign n32441 = ~n32438 & n32440;
  assign n32442 = ~pi54 & ~n32441;
  assign n32443 = ~n32437 & n32442;
  assign n32444 = n6307 & ~n32434;
  assign n32445 = ~n6307 & ~n32389;
  assign n32446 = ~n32444 & ~n32445;
  assign n32447 = pi54 & ~n32446;
  assign n32448 = ~pi74 & ~n32447;
  assign n32449 = ~n32443 & n32448;
  assign n32450 = ~pi54 & n32444;
  assign n32451 = ~n31593 & ~n32389;
  assign n32452 = pi74 & ~n32451;
  assign n32453 = ~n32450 & n32452;
  assign n32454 = ~pi55 & ~n32453;
  assign n32455 = ~n32449 & n32454;
  assign n32456 = pi55 & ~n32375;
  assign n32457 = ~n60258 & n32456;
  assign n32458 = n4437 & ~n32457;
  assign n32459 = ~n32455 & n32458;
  assign n32460 = ~n4437 & n32375;
  assign n32461 = ~pi59 & ~n32460;
  assign n32462 = ~n32459 & n32461;
  assign n32463 = n4440 & n60258;
  assign n32464 = pi59 & ~n32375;
  assign n32465 = ~n32463 & n32464;
  assign n32466 = ~pi57 & ~n32465;
  assign n32467 = ~n32462 & n32466;
  assign po178 = ~n32383 & ~n32467;
  assign n32469 = ~pi110 & n29537;
  assign n32470 = ~n2845 & n2852;
  assign n32471 = ~n2845 & n32469;
  assign n32472 = n2852 & n32471;
  assign n32473 = n32469 & n32470;
  assign n32474 = pi39 & ~n60259;
  assign n32475 = n2677 & n2681;
  assign n32476 = n2727 & ~n6416;
  assign n32477 = pi110 & n32476;
  assign n32478 = ~n32475 & n32477;
  assign n32479 = ~n2707 & n32478;
  assign n32480 = ~pi39 & ~n32479;
  assign n32481 = ~n58992 & ~n32480;
  assign n32482 = ~pi39 & pi110;
  assign n32483 = n32476 & n32482;
  assign n32484 = ~n32475 & n32483;
  assign n32485 = ~n2707 & n32484;
  assign n32486 = pi39 & n2852;
  assign n32487 = n32471 & n32486;
  assign n32488 = ~n32485 & ~n32487;
  assign n32489 = ~n58992 & ~n32488;
  assign n32490 = ~n32474 & n32481;
  assign n32491 = pi299 & n60259;
  assign n32492 = n2853 & n32471;
  assign n32493 = n60084 & n32469;
  assign n32494 = pi39 & ~n32493;
  assign n32495 = ~n60261 & n32494;
  assign n32496 = ~n2682 & ~n2707;
  assign n32497 = n32476 & n32496;
  assign n32498 = n2531 & n31468;
  assign n32499 = pi72 & n60073;
  assign n32500 = n32498 & n32499;
  assign n32501 = n58798 & n2565;
  assign n32502 = n2471 & n58797;
  assign n32503 = ~pi50 & n58797;
  assign n32504 = n60078 & n32503;
  assign n32505 = n28401 & n60262;
  assign n32506 = ~pi111 & ~n28378;
  assign n32507 = ~pi36 & n31422;
  assign n32508 = ~n32506 & n32507;
  assign n32509 = n2465 & ~n32508;
  assign n32510 = ~n28340 & ~n31427;
  assign n32511 = ~n32509 & n32510;
  assign n32512 = ~pi83 & ~n32511;
  assign n32513 = n28342 & ~n32512;
  assign n32514 = ~pi71 & ~n32513;
  assign n32515 = n28390 & ~n32514;
  assign n32516 = ~pi81 & ~n32515;
  assign n32517 = n60263 & ~n32516;
  assign n32518 = ~pi90 & ~n32517;
  assign n32519 = n59136 & ~n32518;
  assign n32520 = pi90 & ~n32498;
  assign n32521 = n6346 & ~n32520;
  assign n32522 = n32519 & n32521;
  assign n32523 = ~n32500 & ~n32522;
  assign n32524 = n2621 & ~n32523;
  assign n32525 = ~pi110 & ~n32524;
  assign n32526 = n32497 & ~n32525;
  assign n32527 = ~pi93 & ~n28325;
  assign n32528 = n32519 & n32527;
  assign n32529 = ~pi72 & ~n32528;
  assign n32530 = n28319 & ~n32497;
  assign n32531 = ~n32529 & n32530;
  assign n32532 = ~pi39 & ~n32531;
  assign n32533 = ~n32526 & n32532;
  assign n32534 = ~n32495 & ~n32533;
  assign n32535 = n59292 & ~n32534;
  assign n32536 = pi110 & n32497;
  assign n32537 = ~pi39 & ~n32536;
  assign n32538 = ~n32495 & ~n32537;
  assign n32539 = ~n59292 & ~n32538;
  assign n32540 = n58992 & ~n32539;
  assign n32541 = ~n32535 & n32540;
  assign po281 = ~n60260 & ~n32541;
  assign n32543 = n2635 & n29690;
  assign n32544 = n29067 & ~n60146;
  assign n32545 = pi92 & ~n60264;
  assign n32546 = n6306 & ~n32545;
  assign n32547 = ~pi75 & ~n31164;
  assign n32548 = ~pi299 & ~n29377;
  assign n32549 = pi299 & ~n29462;
  assign n32550 = ~pi232 & ~n32549;
  assign n32551 = ~n32548 & n32550;
  assign n32552 = ~pi39 & ~n32551;
  assign n32553 = pi148 & n2680;
  assign n32554 = ~n29462 & ~n32553;
  assign n32555 = pi148 & n30604;
  assign n32556 = ~n32554 & ~n32555;
  assign n32557 = pi299 & ~n32556;
  assign n32558 = ~n2680 & ~n29377;
  assign n32559 = ~n30627 & ~n32558;
  assign n32560 = ~pi299 & ~n32559;
  assign n32561 = pi141 & n32560;
  assign n32562 = n29089 & ~n32559;
  assign n32563 = ~pi141 & n32548;
  assign n32564 = pi232 & ~n32563;
  assign n32565 = ~n60265 & n32564;
  assign n32566 = ~n32557 & n32564;
  assign n32567 = ~n60265 & n32566;
  assign n32568 = ~n32557 & n32565;
  assign n32569 = n32552 & ~n60266;
  assign n32570 = ~n29548 & ~n30313;
  assign n32571 = n29584 & ~n32570;
  assign n32572 = n30706 & ~n32571;
  assign n32573 = ~n58846 & ~n29548;
  assign n32574 = n29532 & ~n32570;
  assign n32575 = ~n32573 & n32574;
  assign n32576 = n29554 & ~n32575;
  assign n32577 = ~n32572 & ~n32576;
  assign n32578 = ~pi232 & ~n32577;
  assign n32579 = ~n29544 & ~n32570;
  assign n32580 = ~n29553 & ~n32579;
  assign n32581 = pi148 & ~n32580;
  assign n32582 = ~n29090 & ~n32576;
  assign n32583 = ~n32581 & ~n32582;
  assign n32584 = pi141 & n29574;
  assign n32585 = n32571 & ~n32584;
  assign n32586 = ~pi141 & n32572;
  assign n32587 = ~n29574 & n32571;
  assign n32588 = n30706 & ~n32587;
  assign n32589 = pi141 & n32588;
  assign n32590 = ~n32586 & ~n32589;
  assign n32591 = n30706 & ~n32585;
  assign n32592 = ~n32583 & n60267;
  assign n32593 = pi232 & ~n32592;
  assign n32594 = ~n32578 & ~n32593;
  assign n32595 = pi39 & ~n32594;
  assign n32596 = n2636 & ~n32595;
  assign n32597 = ~n32569 & n32596;
  assign n32598 = ~pi87 & ~n32597;
  assign n32599 = n32547 & ~n32598;
  assign n32600 = ~pi92 & ~n32599;
  assign n32601 = n32546 & ~n32600;
  assign n32602 = ~pi55 & ~n32601;
  assign n32603 = n29068 & ~n30745;
  assign n32604 = pi55 & ~n32603;
  assign n32605 = ~n32602 & ~n32604;
  assign n32606 = n4437 & ~n32605;
  assign n32607 = n29070 & ~n32606;
  assign n32608 = pi138 & n32607;
  assign n32609 = ~n2783 & n29090;
  assign n32610 = n2783 & n28507;
  assign n32611 = n29572 & n32610;
  assign n32612 = n29089 & ~n32611;
  assign n32613 = ~n32609 & ~n32612;
  assign n32614 = pi232 & ~n32613;
  assign n32615 = ~n2792 & n28507;
  assign n32616 = n29572 & n32615;
  assign n32617 = ~pi299 & ~n32616;
  assign n32618 = ~n2845 & n28507;
  assign n32619 = n29532 & n32618;
  assign n32620 = pi299 & ~n32619;
  assign n32621 = ~n32617 & ~n32620;
  assign n32622 = pi232 & ~pi299;
  assign n32623 = pi141 & n32622;
  assign n32624 = ~n32621 & ~n32623;
  assign n32625 = ~pi232 & ~n32621;
  assign n32626 = ~n29089 & ~n32621;
  assign n32627 = n32613 & ~n32626;
  assign n32628 = pi232 & ~n32627;
  assign n32629 = ~n32625 & ~n32628;
  assign n32630 = ~n32614 & ~n32624;
  assign n32631 = pi39 & ~n60268;
  assign n32632 = ~pi38 & n59928;
  assign n32633 = ~n29092 & n60166;
  assign n32634 = ~pi39 & ~n32633;
  assign n32635 = n32632 & ~n32634;
  assign n32636 = ~n32631 & n32635;
  assign n32637 = ~pi138 & n32636;
  assign n32638 = ~pi118 & n30770;
  assign n32639 = ~pi139 & n32638;
  assign n32640 = ~n32637 & ~n32639;
  assign n32641 = ~n32608 & n32640;
  assign n32642 = ~pi138 & ~n29933;
  assign n32643 = n32607 & n32642;
  assign n32644 = n32636 & ~n32642;
  assign n32645 = n32639 & ~n32644;
  assign n32646 = ~n32643 & n32645;
  assign po295 = ~n32641 & ~n32646;
  assign n32648 = pi169 & n2680;
  assign n32649 = ~n29462 & ~n32648;
  assign n32650 = pi169 & n30604;
  assign n32651 = ~n32649 & ~n32650;
  assign n32652 = pi299 & ~n32651;
  assign n32653 = pi191 & n32560;
  assign n32654 = n30958 & ~n32559;
  assign n32655 = ~pi191 & n32548;
  assign n32656 = pi232 & ~n32655;
  assign n32657 = ~n60269 & n32656;
  assign n32658 = ~n32652 & n32656;
  assign n32659 = ~n60269 & n32658;
  assign n32660 = ~n32652 & n32657;
  assign n32661 = n32552 & ~n60270;
  assign n32662 = ~pi169 & n29548;
  assign n32663 = ~n32579 & ~n32662;
  assign n32664 = n29532 & ~n32663;
  assign n32665 = n29554 & ~n32664;
  assign n32666 = pi191 & n32588;
  assign n32667 = ~n32665 & ~n32666;
  assign n32668 = pi232 & ~n32667;
  assign n32669 = ~pi191 & n32572;
  assign n32670 = ~n32578 & ~n32669;
  assign n32671 = ~n32665 & ~n32669;
  assign n32672 = ~n32666 & n32671;
  assign n32673 = pi232 & ~n32672;
  assign n32674 = ~n32578 & ~n32673;
  assign n32675 = ~n32668 & n32670;
  assign n32676 = pi39 & ~n60271;
  assign n32677 = n2636 & ~n32676;
  assign n32678 = ~n32661 & n32677;
  assign n32679 = ~pi87 & ~n32678;
  assign n32680 = n32547 & ~n32679;
  assign n32681 = ~pi92 & ~n32680;
  assign n32682 = n32546 & ~n32681;
  assign n32683 = ~pi55 & ~n32682;
  assign n32684 = ~n32604 & ~n32683;
  assign n32685 = n4437 & ~n32684;
  assign n32686 = n29070 & ~n32685;
  assign n32687 = pi139 & n32686;
  assign n32688 = ~n2783 & n30959;
  assign n32689 = ~n32620 & ~n32688;
  assign n32690 = ~pi191 & ~pi299;
  assign n32691 = ~n32616 & n32690;
  assign n32692 = n30958 & ~n32611;
  assign n32693 = ~n32691 & ~n32692;
  assign n32694 = n32689 & n32693;
  assign n32695 = pi232 & ~n32694;
  assign n32696 = ~n32625 & ~n32695;
  assign n32697 = pi39 & ~n32696;
  assign n32698 = n2681 & ~n30960;
  assign n32699 = n60166 & ~n32698;
  assign n32700 = ~pi39 & ~n32699;
  assign n32701 = n32632 & ~n32700;
  assign n32702 = ~n32697 & n32701;
  assign n32703 = ~pi139 & n32702;
  assign n32704 = ~n32638 & ~n32703;
  assign n32705 = ~n32687 & n32704;
  assign n32706 = ~pi139 & ~n29934;
  assign n32707 = n32686 & n32706;
  assign n32708 = n32702 & ~n32706;
  assign n32709 = n32638 & ~n32708;
  assign n32710 = ~n32707 & n32709;
  assign po296 = ~n32705 & ~n32710;
  assign n32712 = pi171 & pi299;
  assign n32713 = ~n2783 & n32712;
  assign n32714 = ~n32620 & ~n32713;
  assign n32715 = ~pi192 & ~pi299;
  assign n32716 = ~n32616 & n32715;
  assign n32717 = pi192 & ~pi299;
  assign n32718 = ~n32611 & n32717;
  assign n32719 = ~n32716 & ~n32718;
  assign n32720 = n32714 & n32719;
  assign n32721 = pi232 & ~n32720;
  assign n32722 = ~n32625 & ~n32721;
  assign n32723 = pi39 & ~n32722;
  assign n32724 = ~n32712 & ~n32717;
  assign n32725 = n2681 & ~n32724;
  assign n32726 = n60166 & ~n32725;
  assign n32727 = ~pi39 & ~n32726;
  assign n32728 = ~pi138 & n32639;
  assign n32729 = ~pi196 & n32728;
  assign n32730 = pi195 & ~n32729;
  assign n32731 = n32632 & ~n32730;
  assign n32732 = ~n32727 & n32731;
  assign n32733 = ~n32723 & n32732;
  assign n32734 = pi171 & n2680;
  assign n32735 = ~n29462 & ~n32734;
  assign n32736 = pi171 & n30604;
  assign n32737 = ~n32735 & ~n32736;
  assign n32738 = pi299 & ~n32737;
  assign n32739 = pi192 & n32560;
  assign n32740 = ~n32559 & n32717;
  assign n32741 = ~pi192 & n32548;
  assign n32742 = pi232 & ~n32741;
  assign n32743 = ~n60272 & n32742;
  assign n32744 = ~n32738 & n32742;
  assign n32745 = ~n60272 & n32744;
  assign n32746 = ~n32738 & n32743;
  assign n32747 = n32552 & ~n60273;
  assign n32748 = ~pi171 & n29548;
  assign n32749 = ~n32579 & ~n32748;
  assign n32750 = n29532 & ~n32749;
  assign n32751 = n29554 & ~n32750;
  assign n32752 = pi192 & n32588;
  assign n32753 = ~n32751 & ~n32752;
  assign n32754 = pi232 & ~n32753;
  assign n32755 = ~pi192 & n32572;
  assign n32756 = ~n32578 & ~n32755;
  assign n32757 = ~n32751 & ~n32755;
  assign n32758 = ~n32752 & n32757;
  assign n32759 = pi232 & ~n32758;
  assign n32760 = ~n32578 & ~n32759;
  assign n32761 = ~n32754 & n32756;
  assign n32762 = pi39 & ~n60274;
  assign n32763 = n2636 & ~n32762;
  assign n32764 = ~n32747 & n32763;
  assign n32765 = ~pi87 & ~n32764;
  assign n32766 = n32547 & ~n32765;
  assign n32767 = ~pi92 & ~n32766;
  assign n32768 = n32546 & ~n32767;
  assign n32769 = ~pi55 & ~n32768;
  assign n32770 = ~n32604 & ~n32769;
  assign n32771 = n4437 & ~n32770;
  assign n32772 = n29070 & n32730;
  assign n32773 = ~n32771 & n32772;
  assign n32774 = ~n32733 & ~n32773;
  assign n32775 = ~pi170 & n29548;
  assign n32776 = ~n32579 & ~n32775;
  assign n32777 = n29532 & ~n32776;
  assign n32778 = n29554 & ~n32777;
  assign n32779 = ~n32572 & ~n32778;
  assign n32780 = pi232 & ~n32779;
  assign n32781 = ~n32578 & ~n32780;
  assign n32782 = pi232 & n32588;
  assign n32783 = n32781 & ~n32782;
  assign n32784 = pi39 & ~n32783;
  assign n32785 = ~pi38 & pi194;
  assign n32786 = ~n32784 & n32785;
  assign n32787 = pi39 & ~n32781;
  assign n32788 = ~pi38 & ~pi194;
  assign n32789 = ~n32787 & n32788;
  assign n32790 = ~n32786 & ~n32789;
  assign n32791 = pi170 & n30604;
  assign n32792 = pi232 & pi299;
  assign n32793 = pi170 & n2680;
  assign n32794 = ~n29462 & ~n32793;
  assign n32795 = n32792 & ~n32794;
  assign n32796 = ~n32791 & n32795;
  assign n32797 = n32552 & ~n32796;
  assign n32798 = ~n32790 & ~n32797;
  assign n32799 = n29377 & n32789;
  assign n32800 = n32559 & n32786;
  assign n32801 = ~n32799 & ~n32800;
  assign n32802 = n32622 & ~n32801;
  assign n32803 = ~n32552 & ~n32790;
  assign n32804 = ~n32560 & n32786;
  assign n32805 = ~n32548 & n32789;
  assign n32806 = ~n32804 & ~n32805;
  assign n32807 = ~n32791 & ~n32794;
  assign n32808 = pi299 & ~n32807;
  assign n32809 = pi232 & ~n32808;
  assign n32810 = ~n32806 & n32809;
  assign n32811 = ~n32803 & ~n32810;
  assign n32812 = ~n32798 & ~n32802;
  assign n32813 = ~pi100 & ~n60275;
  assign n32814 = ~pi87 & ~n32813;
  assign n32815 = n32547 & ~n32814;
  assign n32816 = ~pi92 & ~n32815;
  assign n32817 = n32546 & ~n32816;
  assign n32818 = ~pi55 & ~n32817;
  assign n32819 = ~n32604 & ~n32818;
  assign n32820 = n4437 & ~n32819;
  assign n32821 = n29070 & ~n32820;
  assign n32822 = pi196 & ~n32821;
  assign n32823 = ~pi170 & n29855;
  assign n32824 = ~n32610 & ~n32823;
  assign n32825 = n60188 & ~n32824;
  assign n32826 = ~pi299 & n32611;
  assign n32827 = n60187 & n32610;
  assign n32828 = pi232 & ~n60276;
  assign n32829 = ~n32825 & n32828;
  assign n32830 = ~n32625 & ~n32829;
  assign n32831 = pi299 & ~n32830;
  assign n32832 = ~n32617 & ~n32831;
  assign n32833 = pi39 & ~n32832;
  assign n32834 = n32792 & n32793;
  assign n32835 = n60166 & ~n32834;
  assign n32836 = ~pi39 & ~n32835;
  assign n32837 = ~pi38 & ~n32836;
  assign n32838 = ~n32833 & n32837;
  assign n32839 = ~pi194 & ~n32838;
  assign n32840 = pi39 & ~n32830;
  assign n32841 = pi170 & n2681;
  assign n32842 = ~n29623 & ~n32841;
  assign n32843 = n60166 & n32842;
  assign n32844 = ~pi39 & ~n32843;
  assign n32845 = ~pi38 & ~n32844;
  assign n32846 = ~n32840 & n32845;
  assign n32847 = pi194 & ~n32846;
  assign n32848 = n59928 & ~n32847;
  assign n32849 = ~n32839 & n32848;
  assign n32850 = ~pi196 & ~n32849;
  assign n32851 = ~n32728 & ~n32850;
  assign n32852 = ~n32822 & n32851;
  assign n32853 = pi195 & ~pi196;
  assign n32854 = ~n32821 & n32853;
  assign n32855 = ~n32849 & ~n32853;
  assign n32856 = n32728 & ~n32855;
  assign n32857 = ~n32854 & n32856;
  assign n32858 = ~n32852 & ~n32857;
  assign n32859 = n58992 & n6306;
  assign n32860 = pi128 & pi228;
  assign n32861 = ~n32859 & n32860;
  assign n32862 = n2828 & ~n6544;
  assign n32863 = n58843 & n32862;
  assign n32864 = n2851 & ~n6629;
  assign n32865 = n58847 & n32864;
  assign n32866 = ~n32863 & ~n32865;
  assign n32867 = pi39 & ~n32866;
  assign n32868 = pi93 & n2526;
  assign n32869 = n2562 & n28338;
  assign n32870 = ~pi86 & ~n32869;
  assign n32871 = ~pi83 & n31428;
  assign n32872 = n2446 & n2470;
  assign n32873 = ~pi65 & n2446;
  assign n32874 = ~pi65 & n2470;
  assign n32875 = n2446 & n32874;
  assign n32876 = n2470 & n32873;
  assign n32877 = n2479 & n60277;
  assign n32878 = n2477 & n32872;
  assign n32879 = ~pi69 & n60278;
  assign n32880 = ~pi67 & ~pi71;
  assign n32881 = pi36 & ~pi103;
  assign n32882 = n32880 & n32881;
  assign n32883 = n32879 & n32882;
  assign n32884 = n32871 & n32883;
  assign n32885 = n58802 & n32884;
  assign n32886 = n32870 & ~n32885;
  assign n32887 = n28411 & ~n32886;
  assign n32888 = ~pi97 & ~n32887;
  assign n32889 = ~pi46 & n58838;
  assign n32890 = n28629 & n32889;
  assign n32891 = ~n32888 & n32890;
  assign n32892 = pi299 & n31621;
  assign n32893 = ~n31610 & ~n32892;
  assign n32894 = n2681 & ~n32893;
  assign n32895 = pi109 & ~n32894;
  assign n32896 = n28412 & ~n32870;
  assign n32897 = ~n58838 & n32896;
  assign n32898 = ~n32895 & ~n32897;
  assign n32899 = ~n32891 & n32898;
  assign n32900 = ~n2533 & n32894;
  assign n32901 = ~n28448 & ~n32894;
  assign n32902 = ~n32900 & ~n32901;
  assign n32903 = ~n32899 & n32902;
  assign n32904 = ~pi91 & ~n32903;
  assign n32905 = n2589 & ~n28417;
  assign n32906 = ~n32904 & n32905;
  assign n32907 = ~n32868 & ~n32906;
  assign n32908 = ~pi32 & n6860;
  assign n32909 = ~pi39 & n58809;
  assign n32910 = ~pi39 & n2599;
  assign n32911 = n2597 & n32908;
  assign n32912 = ~pi96 & n60280;
  assign n32913 = n2601 & n32908;
  assign n32914 = n58809 & n2614;
  assign n32915 = ~pi39 & n32914;
  assign n32916 = n2614 & n60279;
  assign n32917 = ~n32907 & n60281;
  assign n32918 = ~n32867 & ~n32917;
  assign n32919 = ~pi38 & ~n32918;
  assign n32920 = ~pi228 & n32919;
  assign n32921 = ~n32860 & ~n32920;
  assign n32922 = ~pi100 & ~n32921;
  assign n32923 = ~n31587 & ~n32860;
  assign n32924 = pi100 & ~n32923;
  assign n32925 = ~pi87 & ~n32924;
  assign n32926 = ~n32922 & n32925;
  assign n32927 = pi87 & ~n32860;
  assign n32928 = ~pi75 & ~n32927;
  assign n32929 = ~n32926 & n32928;
  assign n32930 = ~n60247 & ~n32860;
  assign n32931 = pi75 & ~n32930;
  assign n32932 = ~pi92 & ~n32931;
  assign n32933 = ~n32929 & n32932;
  assign n32934 = n58815 & n31586;
  assign n32935 = n6309 & n32934;
  assign n32936 = ~pi75 & n60247;
  assign n32937 = n60069 & n31586;
  assign n32938 = pi92 & ~n32860;
  assign n32939 = ~n60282 & n32938;
  assign n32940 = n32859 & ~n32939;
  assign n32941 = ~n32933 & n32940;
  assign n32942 = ~n32861 & ~n32941;
  assign n32943 = pi743 & pi947;
  assign n32944 = pi907 & ~pi947;
  assign n32945 = pi735 & n32944;
  assign n32946 = ~n32943 & ~n32945;
  assign n32947 = n59152 & ~n32946;
  assign n32948 = pi146 & n59293;
  assign n32949 = pi146 & ~n59152;
  assign n32950 = ~n2841 & n32949;
  assign n32951 = pi146 & ~n6615;
  assign n32952 = n2841 & n32951;
  assign n32953 = pi735 & pi907;
  assign n32954 = n59152 & n32953;
  assign n32955 = ~pi947 & ~n32954;
  assign n32956 = ~n32952 & n32955;
  assign n32957 = pi743 & n59152;
  assign n32958 = pi947 & ~n32949;
  assign n32959 = ~n32957 & n32958;
  assign n32960 = ~n32956 & ~n32959;
  assign n32961 = ~n32950 & ~n32960;
  assign n32962 = ~n32947 & ~n32948;
  assign n32963 = ~n6629 & ~n60283;
  assign n32964 = ~pi146 & ~n6464;
  assign n32965 = n6464 & n32946;
  assign n32966 = n6464 & ~n32946;
  assign n32967 = pi146 & ~n6464;
  assign n32968 = ~n32966 & ~n32967;
  assign n32969 = ~n32964 & ~n32965;
  assign n32970 = n6629 & ~n60284;
  assign n32971 = ~pi215 & ~n32970;
  assign n32972 = ~n32963 & n32971;
  assign n32973 = pi146 & n6650;
  assign n32974 = n6512 & ~n32946;
  assign n32975 = pi215 & ~n32974;
  assign n32976 = ~n32973 & n32975;
  assign n32977 = pi299 & ~n32976;
  assign n32978 = ~n32972 & n32977;
  assign n32979 = n6615 & ~n32946;
  assign n32980 = n2790 & ~n32951;
  assign n32981 = ~n32979 & n32980;
  assign n32982 = ~n2790 & ~n32947;
  assign n32983 = ~n2790 & ~n32949;
  assign n32984 = ~n32947 & n32983;
  assign n32985 = ~n32949 & n32982;
  assign n32986 = ~n6544 & ~n60285;
  assign n32987 = ~n32981 & n32986;
  assign n32988 = n6544 & ~n60284;
  assign n32989 = ~pi223 & ~n32988;
  assign n32990 = ~n32987 & n32989;
  assign n32991 = pi146 & ~n6512;
  assign n32992 = ~n32974 & ~n32991;
  assign n32993 = ~n2790 & ~n32992;
  assign n32994 = n59149 & n32946;
  assign n32995 = ~pi146 & ~n59149;
  assign n32996 = n2790 & ~n32995;
  assign n32997 = n2790 & ~n32994;
  assign n32998 = ~n32995 & n32997;
  assign n32999 = ~n32994 & n32996;
  assign n33000 = pi223 & ~n60286;
  assign n33001 = ~n32993 & n33000;
  assign n33002 = ~pi299 & ~n33001;
  assign n33003 = ~n32990 & n33002;
  assign n33004 = pi39 & ~n33003;
  assign n33005 = ~n32972 & ~n32976;
  assign n33006 = pi299 & ~n33005;
  assign n33007 = ~n32981 & ~n60285;
  assign n33008 = ~n6544 & ~n33007;
  assign n33009 = n6544 & n60284;
  assign n33010 = ~pi223 & ~n33009;
  assign n33011 = ~n33008 & n33010;
  assign n33012 = ~n32993 & ~n60286;
  assign n33013 = pi223 & ~n33012;
  assign n33014 = ~pi299 & ~n33013;
  assign n33015 = ~n33011 & n33014;
  assign n33016 = ~n33006 & ~n33015;
  assign n33017 = pi39 & ~n33016;
  assign n33018 = ~n32978 & n33004;
  assign n33019 = n6453 & ~n32946;
  assign n33020 = pi146 & ~n6453;
  assign n33021 = pi299 & ~n33020;
  assign n33022 = ~n33019 & n33021;
  assign n33023 = n6449 & ~n32946;
  assign n33024 = pi146 & ~n6449;
  assign n33025 = ~pi299 & ~n33024;
  assign n33026 = ~n33023 & n33025;
  assign n33027 = ~n33022 & ~n33026;
  assign n33028 = n6449 & n32946;
  assign n33029 = ~pi146 & ~n6449;
  assign n33030 = ~pi299 & ~n33029;
  assign n33031 = ~n33028 & n33030;
  assign n33032 = ~pi146 & ~n6453;
  assign n33033 = n6453 & n32946;
  assign n33034 = pi299 & ~n33033;
  assign n33035 = pi299 & ~n33032;
  assign n33036 = ~n33033 & n33035;
  assign n33037 = ~n33032 & n33034;
  assign n33038 = ~pi39 & ~n60288;
  assign n33039 = ~n33031 & n33038;
  assign n33040 = ~pi39 & ~n33031;
  assign n33041 = ~n60288 & n33040;
  assign n33042 = ~pi39 & ~n33027;
  assign n33043 = ~pi38 & ~n60289;
  assign n33044 = ~n60287 & n33043;
  assign n33045 = ~pi146 & ~n6863;
  assign n33046 = n2794 & n32946;
  assign n33047 = n6863 & n32946;
  assign n33048 = n59171 & n33046;
  assign n33049 = pi38 & ~n60290;
  assign n33050 = pi38 & ~n33045;
  assign n33051 = ~n60290 & n33050;
  assign n33052 = ~n33045 & n33049;
  assign n33053 = n59928 & ~n60291;
  assign n33054 = ~n33044 & n33053;
  assign n33055 = ~pi146 & ~n59928;
  assign n33056 = ~pi832 & ~n33055;
  assign n33057 = ~n33054 & n33056;
  assign n33058 = ~pi146 & ~n2794;
  assign n33059 = pi832 & ~n33058;
  assign n33060 = ~n33046 & n33059;
  assign n33061 = ~n33057 & ~n33060;
  assign n33062 = ~pi770 & pi947;
  assign n33063 = pi726 & n32944;
  assign n33064 = ~n33062 & ~n33063;
  assign n33065 = n2794 & ~n33064;
  assign n33066 = ~pi147 & ~n2794;
  assign n33067 = pi832 & ~n33066;
  assign n33068 = ~n33065 & n33067;
  assign n33069 = pi215 & pi947;
  assign n33070 = n6512 & n33069;
  assign n33071 = pi215 & ~n6649;
  assign n33072 = n6637 & ~n32944;
  assign n33073 = pi947 & n59152;
  assign n33074 = ~n6633 & ~n33073;
  assign n33075 = ~n6629 & ~n33074;
  assign n33076 = ~pi215 & ~n33075;
  assign n33077 = ~n33072 & n33076;
  assign n33078 = ~n33071 & ~n33077;
  assign n33079 = ~n33070 & ~n33078;
  assign n33080 = pi299 & ~n33079;
  assign n33081 = ~pi299 & ~n32944;
  assign n33082 = ~pi299 & n6627;
  assign n33083 = ~n32944 & n33082;
  assign n33084 = n6627 & n33081;
  assign n33085 = ~n33080 & ~n60292;
  assign n33086 = pi39 & ~n33085;
  assign n33087 = n59147 & ~n32944;
  assign n33088 = ~pi39 & n33087;
  assign n33089 = ~n33086 & ~n33088;
  assign n33090 = ~pi147 & n33089;
  assign n33091 = n6512 & n32944;
  assign n33092 = pi215 & ~n33091;
  assign n33093 = n59152 & n32944;
  assign n33094 = ~n6629 & ~n33093;
  assign n33095 = pi907 & n6464;
  assign n33096 = ~pi947 & n33095;
  assign n33097 = n6629 & ~n33096;
  assign n33098 = ~n33094 & ~n33097;
  assign n33099 = ~pi215 & ~n33098;
  assign n33100 = ~n33092 & ~n33099;
  assign n33101 = pi299 & ~n33100;
  assign n33102 = n6627 & n32944;
  assign n33103 = ~pi299 & ~n33102;
  assign n33104 = ~n33101 & ~n33103;
  assign n33105 = pi39 & ~n33104;
  assign n33106 = n59147 & n32944;
  assign n33107 = ~pi39 & ~n33106;
  assign n33108 = ~n33105 & ~n33107;
  assign n33109 = pi147 & n33108;
  assign n33110 = ~pi38 & ~n33109;
  assign n33111 = ~n33090 & n33110;
  assign n33112 = ~pi147 & ~n6863;
  assign n33113 = n6863 & n32944;
  assign n33114 = pi38 & ~n33113;
  assign n33115 = ~n33112 & n33114;
  assign n33116 = pi770 & ~n33115;
  assign n33117 = ~n33111 & n33116;
  assign n33118 = pi299 & ~n33078;
  assign n33119 = ~n6621 & ~n59155;
  assign n33120 = n2840 & ~n33119;
  assign n33121 = ~pi223 & ~n33120;
  assign n33122 = ~pi947 & n59150;
  assign n33123 = pi223 & ~n33122;
  assign n33124 = n59150 & ~n32944;
  assign n33125 = pi223 & ~n33124;
  assign n33126 = ~n33123 & ~n33125;
  assign n33127 = ~n33121 & n33126;
  assign n33128 = ~pi299 & ~n33127;
  assign n33129 = pi299 & pi947;
  assign n33130 = ~n33128 & ~n33129;
  assign n33131 = ~n33118 & ~n33129;
  assign n33132 = ~n33128 & n33131;
  assign n33133 = ~n33118 & n33130;
  assign n33134 = pi39 & n60293;
  assign n33135 = ~n2840 & n59147;
  assign n33136 = ~pi39 & ~n33135;
  assign n33137 = n59147 & n33136;
  assign n33138 = ~n33134 & ~n33137;
  assign n33139 = ~pi147 & n33138;
  assign n33140 = pi215 & ~n6645;
  assign n33141 = ~n2840 & n6464;
  assign n33142 = n6629 & n33141;
  assign n33143 = ~n2840 & n6637;
  assign n33144 = ~pi215 & ~n60294;
  assign n33145 = n6629 & ~n33141;
  assign n33146 = ~n6640 & ~n33145;
  assign n33147 = ~pi215 & ~n33146;
  assign n33148 = ~n6636 & n33144;
  assign n33149 = ~n33140 & ~n60295;
  assign n33150 = pi299 & ~n33149;
  assign n33151 = ~n2840 & n6627;
  assign n33152 = ~pi299 & ~n33151;
  assign n33153 = ~pi299 & n33151;
  assign n33154 = pi299 & ~n60295;
  assign n33155 = pi299 & ~n33140;
  assign n33156 = ~n60295 & n33155;
  assign n33157 = ~n33140 & n33154;
  assign n33158 = ~n33153 & ~n60296;
  assign n33159 = ~n33150 & ~n33152;
  assign n33160 = pi39 & n60297;
  assign n33161 = ~n33136 & ~n33160;
  assign n33162 = pi147 & n33161;
  assign n33163 = ~pi38 & ~n33162;
  assign n33164 = ~n33139 & n33163;
  assign n33165 = n2840 & n6863;
  assign n33166 = ~pi147 & ~n33165;
  assign n33167 = ~n2840 & n6863;
  assign n33168 = pi38 & ~n33167;
  assign n33169 = ~n33166 & n33168;
  assign n33170 = ~pi770 & ~n33169;
  assign n33171 = ~n33164 & n33170;
  assign n33172 = pi726 & ~n33171;
  assign n33173 = pi726 & ~n33117;
  assign n33174 = ~n33171 & n33173;
  assign n33175 = ~n33117 & n33172;
  assign n33176 = ~pi947 & n59147;
  assign n33177 = ~pi39 & ~n33176;
  assign n33178 = ~pi947 & n6637;
  assign n33179 = ~n6633 & ~n33093;
  assign n33180 = ~n6629 & ~n33179;
  assign n33181 = ~pi215 & ~n33180;
  assign n33182 = ~n33178 & n33181;
  assign n33183 = n33071 & ~n33091;
  assign n33184 = ~n33182 & ~n33183;
  assign n33185 = pi299 & ~n33184;
  assign n33186 = ~n6628 & ~n33185;
  assign n33187 = pi947 & n6627;
  assign n33188 = pi947 & n33082;
  assign n33189 = ~pi299 & n33187;
  assign n33190 = n33186 & ~n60299;
  assign n33191 = pi39 & ~n33190;
  assign n33192 = ~n33177 & ~n33191;
  assign n33193 = ~pi38 & n33192;
  assign n33194 = pi38 & ~pi947;
  assign n33195 = n6863 & n33194;
  assign n33196 = ~n33193 & ~n33195;
  assign n33197 = ~pi770 & ~n33196;
  assign n33198 = ~pi147 & ~n19469;
  assign n33199 = ~pi770 & n33196;
  assign n33200 = ~n19475 & ~n33199;
  assign n33201 = ~pi147 & ~n33200;
  assign n33202 = ~n33197 & n33198;
  assign n33203 = ~n7552 & ~n33195;
  assign n33204 = pi947 & n59147;
  assign n33205 = ~pi39 & ~n33204;
  assign n33206 = ~pi299 & ~n33187;
  assign n33207 = pi299 & ~n33070;
  assign n33208 = ~n6629 & ~n33073;
  assign n33209 = pi947 & n6464;
  assign n33210 = n6629 & ~n33209;
  assign n33211 = ~pi215 & ~n33210;
  assign n33212 = ~n33208 & n33211;
  assign n33213 = n33207 & ~n33212;
  assign n33214 = ~n33206 & ~n33213;
  assign n33215 = pi39 & ~n33214;
  assign n33216 = ~n33205 & ~n33215;
  assign n33217 = ~pi38 & ~n33216;
  assign n33218 = n33203 & ~n33217;
  assign n33219 = pi147 & ~pi770;
  assign n33220 = n33218 & n33219;
  assign n33221 = ~pi726 & ~n33220;
  assign n33222 = ~n60300 & n33221;
  assign n33223 = n59928 & ~n33222;
  assign n33224 = n59928 & ~n60298;
  assign n33225 = ~n33222 & n33224;
  assign n33226 = ~n60298 & n33223;
  assign n33227 = ~pi147 & ~n59928;
  assign n33228 = ~pi832 & ~n33227;
  assign n33229 = ~n60301 & n33228;
  assign po304 = ~n33068 & ~n33229;
  assign n33231 = ~pi148 & n60293;
  assign n33232 = pi148 & n60297;
  assign n33233 = pi749 & ~n33232;
  assign n33234 = ~n33231 & n33233;
  assign n33235 = ~n29090 & ~n33085;
  assign n33236 = ~n6628 & ~n33101;
  assign n33237 = pi148 & ~n33236;
  assign n33238 = ~pi749 & ~n33237;
  assign n33239 = ~n33235 & n33238;
  assign n33240 = pi39 & ~n33239;
  assign n33241 = ~n33235 & ~n33237;
  assign n33242 = ~pi749 & ~n33241;
  assign n33243 = ~pi148 & ~n60293;
  assign n33244 = pi148 & ~n60297;
  assign n33245 = pi749 & ~n33244;
  assign n33246 = ~n33243 & n33245;
  assign n33247 = ~n33242 & ~n33246;
  assign n33248 = pi39 & ~n33247;
  assign n33249 = pi39 & ~n33234;
  assign n33250 = ~n33239 & n33249;
  assign n33251 = ~n33234 & n33240;
  assign n33252 = ~pi148 & ~n59147;
  assign n33253 = ~pi39 & ~n33252;
  assign n33254 = ~pi749 & pi947;
  assign n33255 = n33135 & ~n33254;
  assign n33256 = n33253 & ~n33255;
  assign n33257 = ~pi38 & ~n33256;
  assign n33258 = ~n60302 & n33257;
  assign n33259 = n33167 & ~n33254;
  assign n33260 = ~pi148 & ~n6863;
  assign n33261 = ~n33259 & ~n33260;
  assign n33262 = pi38 & ~n33261;
  assign n33263 = pi706 & ~n33262;
  assign n33264 = ~n33258 & n33263;
  assign n33265 = ~pi148 & ~n33184;
  assign n33266 = ~n33070 & ~n33212;
  assign n33267 = pi148 & ~n33266;
  assign n33268 = pi299 & ~n33267;
  assign n33269 = ~n33265 & n33268;
  assign n33270 = ~pi148 & ~n6627;
  assign n33271 = n33206 & ~n33270;
  assign n33272 = pi749 & ~n33271;
  assign n33273 = ~n33269 & n33272;
  assign n33274 = ~pi148 & ~pi749;
  assign n33275 = ~n6654 & n33274;
  assign n33276 = pi39 & ~n33275;
  assign n33277 = ~n33273 & n33276;
  assign n33278 = pi749 & pi947;
  assign n33279 = n59147 & n33278;
  assign n33280 = n33253 & ~n33279;
  assign n33281 = ~pi38 & ~n33280;
  assign n33282 = ~n33277 & n33281;
  assign n33283 = pi148 & ~n6863;
  assign n33284 = n2794 & ~n33278;
  assign n33285 = n6863 & ~n33278;
  assign n33286 = n59171 & n33284;
  assign n33287 = pi38 & ~n60303;
  assign n33288 = ~n33283 & n33287;
  assign n33289 = ~pi706 & ~n33288;
  assign n33290 = ~n33282 & n33289;
  assign n33291 = n25257 & ~n33290;
  assign n33292 = ~n33264 & n33291;
  assign n33293 = ~pi148 & ~n25257;
  assign n33294 = ~pi57 & ~n33293;
  assign n33295 = ~n33292 & n33294;
  assign n33296 = pi57 & pi148;
  assign n33297 = ~pi832 & ~n33296;
  assign n33298 = ~n33295 & n33297;
  assign n33299 = pi706 & n32944;
  assign n33300 = n33284 & ~n33299;
  assign n33301 = pi148 & ~n2794;
  assign n33302 = pi832 & ~n33301;
  assign n33303 = ~n33300 & n33302;
  assign n33304 = ~n33298 & ~n33303;
  assign n33305 = ~pi755 & pi947;
  assign n33306 = ~pi725 & n32944;
  assign n33307 = ~n33305 & ~n33306;
  assign n33308 = n2794 & ~n33307;
  assign n33309 = ~pi149 & ~n2794;
  assign n33310 = pi832 & ~n33309;
  assign n33311 = ~n33308 & n33310;
  assign n33312 = ~pi149 & n60293;
  assign n33313 = pi149 & n60297;
  assign n33314 = ~pi755 & ~n33313;
  assign n33315 = ~n33312 & n33314;
  assign n33316 = ~pi149 & n33080;
  assign n33317 = pi149 & ~n33236;
  assign n33318 = pi755 & ~n60292;
  assign n33319 = ~n33317 & n33318;
  assign n33320 = ~n33316 & n33319;
  assign n33321 = pi39 & ~n33320;
  assign n33322 = ~n60292 & ~n33317;
  assign n33323 = ~n33316 & n33322;
  assign n33324 = pi755 & ~n33323;
  assign n33325 = ~pi149 & ~n60293;
  assign n33326 = pi149 & ~n60297;
  assign n33327 = ~pi755 & ~n33326;
  assign n33328 = ~n33325 & n33327;
  assign n33329 = ~n33324 & ~n33328;
  assign n33330 = pi39 & ~n33329;
  assign n33331 = ~n33315 & n33321;
  assign n33332 = n59147 & n33305;
  assign n33333 = ~pi149 & ~n59147;
  assign n33334 = ~pi39 & ~n33333;
  assign n33335 = ~pi39 & ~n33332;
  assign n33336 = ~n33333 & n33335;
  assign n33337 = ~n33332 & n33334;
  assign n33338 = ~n33106 & n60305;
  assign n33339 = ~pi38 & ~n33338;
  assign n33340 = ~n60304 & n33339;
  assign n33341 = n6863 & ~n33305;
  assign n33342 = ~n32944 & n33341;
  assign n33343 = pi149 & ~n6863;
  assign n33344 = pi38 & ~n33343;
  assign n33345 = ~n33342 & n33344;
  assign n33346 = ~pi725 & ~n33345;
  assign n33347 = ~n33340 & n33346;
  assign n33348 = ~pi149 & ~n33184;
  assign n33349 = ~pi149 & pi299;
  assign n33350 = ~n33213 & ~n33349;
  assign n33351 = ~n33348 & ~n33350;
  assign n33352 = ~pi149 & ~n6627;
  assign n33353 = n33206 & ~n33352;
  assign n33354 = ~pi755 & ~n33353;
  assign n33355 = ~n33351 & n33354;
  assign n33356 = ~pi149 & pi755;
  assign n33357 = ~n6654 & n33356;
  assign n33358 = pi39 & ~n33357;
  assign n33359 = ~n33355 & n33358;
  assign n33360 = ~pi38 & ~n60305;
  assign n33361 = ~n33359 & n33360;
  assign n33362 = pi38 & ~n33341;
  assign n33363 = ~n33343 & n33362;
  assign n33364 = pi725 & ~n33363;
  assign n33365 = ~n33361 & n33364;
  assign n33366 = n59928 & ~n33365;
  assign n33367 = ~n33361 & ~n33363;
  assign n33368 = pi725 & ~n33367;
  assign n33369 = ~n60304 & ~n33338;
  assign n33370 = ~pi38 & ~n33369;
  assign n33371 = ~n32944 & ~n33305;
  assign n33372 = ~n2840 & n6468;
  assign n33373 = pi755 & pi947;
  assign n33374 = ~pi39 & ~n33373;
  assign n33375 = n33372 & n33374;
  assign n33376 = n6863 & ~n33371;
  assign n33377 = ~pi149 & ~n6863;
  assign n33378 = pi38 & ~n33377;
  assign n33379 = ~n60306 & n33378;
  assign n33380 = ~pi725 & ~n33379;
  assign n33381 = ~n33370 & n33380;
  assign n33382 = ~n33368 & ~n33381;
  assign n33383 = n59928 & ~n33382;
  assign n33384 = ~n33347 & n33366;
  assign n33385 = ~pi149 & ~n59928;
  assign n33386 = ~pi832 & ~n33385;
  assign n33387 = ~n60307 & n33386;
  assign po306 = ~n33311 & ~n33387;
  assign n33389 = ~pi751 & pi947;
  assign n33390 = ~n32944 & ~n33389;
  assign n33391 = n2794 & ~n33390;
  assign n33392 = pi701 & ~n33389;
  assign n33393 = ~pi701 & n32944;
  assign n33394 = ~n33389 & ~n33393;
  assign n33395 = n2794 & ~n33394;
  assign n33396 = n33391 & ~n33392;
  assign n33397 = ~pi150 & ~n2794;
  assign n33398 = pi832 & ~n33397;
  assign n33399 = ~n60308 & n33398;
  assign n33400 = ~pi150 & ~n60293;
  assign n33401 = pi150 & ~n60297;
  assign n33402 = ~pi751 & ~n33401;
  assign n33403 = ~n33400 & n33402;
  assign n33404 = ~pi150 & n33085;
  assign n33405 = pi150 & n33104;
  assign n33406 = pi751 & ~n33405;
  assign n33407 = ~n33404 & n33406;
  assign n33408 = pi39 & ~n33407;
  assign n33409 = ~pi150 & ~n33085;
  assign n33410 = pi150 & ~n33104;
  assign n33411 = pi751 & ~n33410;
  assign n33412 = ~n33409 & n33411;
  assign n33413 = ~pi150 & n60293;
  assign n33414 = pi150 & n60297;
  assign n33415 = ~pi751 & ~n33414;
  assign n33416 = ~n33413 & n33415;
  assign n33417 = ~n33412 & ~n33416;
  assign n33418 = pi39 & ~n33417;
  assign n33419 = ~n33403 & n33408;
  assign n33420 = n33087 & ~n33389;
  assign n33421 = pi150 & ~n59147;
  assign n33422 = ~pi39 & ~n33421;
  assign n33423 = ~n33420 & n33422;
  assign n33424 = ~pi38 & ~n33423;
  assign n33425 = ~n60309 & n33424;
  assign n33426 = ~pi150 & ~n6863;
  assign n33427 = pi751 & pi947;
  assign n33428 = ~pi39 & ~n33427;
  assign n33429 = n33372 & n33428;
  assign n33430 = n6863 & ~n33390;
  assign n33431 = n59171 & n33391;
  assign n33432 = pi38 & ~n60310;
  assign n33433 = pi38 & ~n33426;
  assign n33434 = ~n60310 & n33433;
  assign n33435 = ~n33426 & n33432;
  assign n33436 = ~pi701 & ~n60311;
  assign n33437 = ~n33425 & n33436;
  assign n33438 = ~pi150 & n33190;
  assign n33439 = pi150 & ~n33214;
  assign n33440 = ~pi751 & ~n33439;
  assign n33441 = ~n33438 & n33440;
  assign n33442 = ~pi150 & pi751;
  assign n33443 = ~n6654 & n33442;
  assign n33444 = ~n33441 & ~n33443;
  assign n33445 = pi39 & ~n33444;
  assign n33446 = ~n18433 & ~n33421;
  assign n33447 = n33177 & n33446;
  assign n33448 = ~pi38 & ~n33447;
  assign n33449 = ~n33445 & n33448;
  assign n33450 = pi150 & ~n6863;
  assign n33451 = n6863 & ~n33389;
  assign n33452 = ~n33450 & ~n33451;
  assign n33453 = pi38 & ~n33452;
  assign n33454 = pi701 & ~n33453;
  assign n33455 = ~n33449 & n33454;
  assign n33456 = ~n33437 & ~n33455;
  assign n33457 = n59928 & ~n33456;
  assign n33458 = ~pi150 & ~n59928;
  assign n33459 = ~pi832 & ~n33458;
  assign n33460 = ~n33457 & n33459;
  assign po307 = ~n33399 & ~n33460;
  assign n33462 = ~pi745 & pi947;
  assign n33463 = ~pi723 & n32944;
  assign n33464 = ~n33462 & ~n33463;
  assign n33465 = n2794 & ~n33464;
  assign n33466 = ~pi151 & ~n2794;
  assign n33467 = pi832 & ~n33466;
  assign n33468 = ~n33465 & n33467;
  assign n33469 = ~pi151 & ~n59147;
  assign n33470 = ~pi745 & n33204;
  assign n33471 = ~n33469 & ~n33470;
  assign n33472 = n33107 & n33471;
  assign n33473 = pi151 & ~n33151;
  assign n33474 = n33128 & ~n33473;
  assign n33475 = ~n6649 & ~n33091;
  assign n33476 = ~pi151 & n33475;
  assign n33477 = ~n6645 & ~n33476;
  assign n33478 = pi215 & ~n33477;
  assign n33479 = pi151 & ~n6629;
  assign n33480 = pi151 & n6640;
  assign n33481 = ~n6635 & n33479;
  assign n33482 = ~n6634 & ~n60312;
  assign n33483 = ~pi151 & ~n6464;
  assign n33484 = n33097 & ~n33483;
  assign n33485 = ~n33141 & n33484;
  assign n33486 = ~pi215 & ~n33485;
  assign n33487 = n33482 & n33486;
  assign n33488 = ~n33478 & ~n33487;
  assign n33489 = pi299 & ~n33488;
  assign n33490 = ~n33474 & ~n33489;
  assign n33491 = ~pi745 & ~n33490;
  assign n33492 = n33482 & ~n33484;
  assign n33493 = n33076 & n33492;
  assign n33494 = ~n33478 & ~n33493;
  assign n33495 = ~n33070 & ~n33494;
  assign n33496 = pi299 & ~n33495;
  assign n33497 = ~pi151 & ~n6627;
  assign n33498 = n33103 & ~n33497;
  assign n33499 = pi745 & ~n33498;
  assign n33500 = ~n33496 & n33499;
  assign n33501 = pi39 & ~n33500;
  assign n33502 = ~n33496 & ~n33498;
  assign n33503 = pi745 & ~n33502;
  assign n33504 = ~pi745 & ~n33489;
  assign n33505 = ~n33474 & n33504;
  assign n33506 = ~n33503 & ~n33505;
  assign n33507 = pi39 & ~n33506;
  assign n33508 = ~n33491 & n33501;
  assign n33509 = ~n33472 & ~n60313;
  assign n33510 = ~pi38 & ~n33509;
  assign n33511 = ~n32944 & ~n33462;
  assign n33512 = pi745 & pi947;
  assign n33513 = ~pi39 & ~n33512;
  assign n33514 = n33372 & n33513;
  assign n33515 = n6863 & ~n33511;
  assign n33516 = ~pi151 & ~n6863;
  assign n33517 = pi38 & ~n33516;
  assign n33518 = pi151 & ~n6863;
  assign n33519 = n6863 & ~n33462;
  assign n33520 = ~n32944 & n33519;
  assign n33521 = ~n33518 & ~n33520;
  assign n33522 = pi38 & ~n33521;
  assign n33523 = ~n60314 & n33517;
  assign n33524 = ~pi723 & ~n60315;
  assign n33525 = ~n33510 & n33524;
  assign n33526 = ~pi745 & ~n6628;
  assign n33527 = ~pi151 & ~n6654;
  assign n33528 = ~n33526 & n33527;
  assign n33529 = n33210 & ~n33483;
  assign n33530 = n33482 & ~n33529;
  assign n33531 = n33181 & n33530;
  assign n33532 = ~n33091 & n33478;
  assign n33533 = n33092 & ~n33477;
  assign n33534 = pi299 & ~n60316;
  assign n33535 = ~n33531 & n33534;
  assign n33536 = ~pi745 & ~n33206;
  assign n33537 = ~n33535 & n33536;
  assign n33538 = ~n33528 & ~n33537;
  assign n33539 = pi39 & ~n33538;
  assign n33540 = ~pi39 & ~n33471;
  assign n33541 = ~pi38 & ~n33540;
  assign n33542 = ~n33539 & n33541;
  assign n33543 = ~n33518 & ~n33519;
  assign n33544 = pi38 & ~n33543;
  assign n33545 = pi723 & ~n33544;
  assign n33546 = ~n33542 & n33545;
  assign n33547 = ~n33525 & ~n33546;
  assign n33548 = n59928 & ~n33547;
  assign n33549 = ~pi151 & ~n59928;
  assign n33550 = ~pi832 & ~n33549;
  assign n33551 = ~n33548 & n33550;
  assign po308 = ~n33468 & ~n33551;
  assign n33553 = pi152 & ~n6464;
  assign n33554 = ~n33141 & ~n33553;
  assign n33555 = n6629 & n33554;
  assign n33556 = ~pi215 & ~n33555;
  assign n33557 = pi152 & n33074;
  assign n33558 = n33094 & ~n33557;
  assign n33559 = ~n6635 & n33558;
  assign n33560 = n33556 & ~n33559;
  assign n33561 = ~pi152 & ~n6645;
  assign n33562 = n33071 & ~n33561;
  assign n33563 = pi299 & ~n33562;
  assign n33564 = ~n33560 & n33563;
  assign n33565 = ~pi152 & ~n59154;
  assign n33566 = ~pi947 & n59154;
  assign n33567 = ~n6544 & ~n33566;
  assign n33568 = ~n33565 & n33567;
  assign n33569 = ~n2840 & n59154;
  assign n33570 = ~n6544 & ~n33569;
  assign n33571 = ~n33568 & n33570;
  assign n33572 = n6544 & n33554;
  assign n33573 = ~pi223 & ~n33572;
  assign n33574 = ~n33571 & n33573;
  assign n33575 = ~pi152 & ~n59150;
  assign n33576 = n33125 & ~n33575;
  assign n33577 = n33123 & ~n33575;
  assign n33578 = ~pi299 & ~n33577;
  assign n33579 = ~n33576 & n33578;
  assign n33580 = ~n33574 & n33579;
  assign n33581 = pi759 & ~n33580;
  assign n33582 = pi759 & ~n33564;
  assign n33583 = ~n33580 & n33582;
  assign n33584 = ~n33564 & n33581;
  assign n33585 = ~n33096 & ~n33553;
  assign n33586 = n6544 & ~n33585;
  assign n33587 = n59154 & ~n32944;
  assign n33588 = ~n6544 & ~n33587;
  assign n33589 = ~n33565 & n33588;
  assign n33590 = ~n33586 & ~n33589;
  assign n33591 = ~pi223 & ~n33590;
  assign n33592 = ~pi299 & ~n33576;
  assign n33593 = ~n33591 & n33592;
  assign n33594 = ~n33072 & n33556;
  assign n33595 = ~n33558 & n33594;
  assign n33596 = ~n32944 & ~n33140;
  assign n33597 = n33562 & ~n33596;
  assign n33598 = pi299 & ~n33597;
  assign n33599 = ~n33595 & n33598;
  assign n33600 = ~pi759 & ~n33599;
  assign n33601 = ~n33593 & n33600;
  assign n33602 = pi39 & ~n33601;
  assign n33603 = ~n60317 & n33602;
  assign n33604 = pi759 & n33204;
  assign n33605 = pi152 & ~n59147;
  assign n33606 = ~pi39 & ~n33605;
  assign n33607 = pi759 & pi947;
  assign n33608 = ~pi39 & ~n33607;
  assign n33609 = ~n6459 & ~n33608;
  assign n33610 = ~n33605 & ~n33609;
  assign n33611 = ~n33604 & n33606;
  assign n33612 = ~n33106 & n60318;
  assign n33613 = ~pi38 & ~n33612;
  assign n33614 = ~n33603 & n33613;
  assign n33615 = n6468 & ~n32944;
  assign n33616 = n6863 & ~n33607;
  assign n33617 = ~n32944 & n33616;
  assign n33618 = n33608 & n33615;
  assign n33619 = ~pi152 & ~n6863;
  assign n33620 = pi38 & ~n33619;
  assign n33621 = ~n60319 & n33620;
  assign n33622 = pi696 & ~n33621;
  assign n33623 = ~n33614 & n33622;
  assign n33624 = ~n33180 & ~n33558;
  assign n33625 = ~n33073 & ~n33624;
  assign n33626 = ~n33209 & ~n33553;
  assign n33627 = n6629 & n33626;
  assign n33628 = ~pi215 & ~n33627;
  assign n33629 = ~n33625 & n33628;
  assign n33630 = pi152 & n33183;
  assign n33631 = n33207 & ~n33630;
  assign n33632 = ~n33629 & n33631;
  assign n33633 = n6544 & ~n33626;
  assign n33634 = ~n33568 & ~n33633;
  assign n33635 = ~pi223 & ~n33634;
  assign n33636 = n33578 & ~n33635;
  assign n33637 = pi759 & ~n33636;
  assign n33638 = ~n33632 & n33637;
  assign n33639 = pi152 & n12074;
  assign n33640 = pi39 & ~n33639;
  assign n33641 = ~n33638 & n33640;
  assign n33642 = ~pi38 & ~n60318;
  assign n33643 = ~n33641 & n33642;
  assign n33644 = pi38 & ~n33616;
  assign n33645 = ~n33619 & n33644;
  assign n33646 = ~pi696 & ~n33645;
  assign n33647 = ~n33643 & n33646;
  assign n33648 = ~n33623 & ~n33647;
  assign n33649 = n59928 & ~n33648;
  assign n33650 = ~pi152 & ~n59928;
  assign n33651 = ~pi832 & ~n33650;
  assign n33652 = ~n33649 & n33651;
  assign n33653 = pi696 & n32944;
  assign n33654 = n2794 & ~n33607;
  assign n33655 = ~n33653 & n33654;
  assign n33656 = ~pi152 & ~n2794;
  assign n33657 = pi832 & ~n33656;
  assign n33658 = ~n33655 & n33657;
  assign n33659 = ~n33652 & ~n33658;
  assign n33660 = pi153 & ~n6863;
  assign n33661 = pi766 & pi947;
  assign n33662 = n2794 & ~n33661;
  assign n33663 = n6863 & ~n33661;
  assign n33664 = n59171 & n33662;
  assign n33665 = pi38 & ~n60320;
  assign n33666 = ~n33660 & n33665;
  assign n33667 = ~pi153 & ~n6627;
  assign n33668 = n33206 & ~n33667;
  assign n33669 = ~pi153 & ~n6464;
  assign n33670 = n33210 & ~n33669;
  assign n33671 = pi153 & ~n6629;
  assign n33672 = pi153 & n6640;
  assign n33673 = ~n6635 & n33671;
  assign n33674 = ~n6634 & ~n60321;
  assign n33675 = ~n33670 & n33674;
  assign n33676 = n33181 & n33675;
  assign n33677 = pi153 & ~n6645;
  assign n33678 = n33071 & ~n33677;
  assign n33679 = ~n33091 & n33678;
  assign n33680 = n33183 & ~n33677;
  assign n33681 = pi299 & ~n60322;
  assign n33682 = ~n33676 & n33681;
  assign n33683 = pi766 & ~n33682;
  assign n33684 = ~n33668 & n33683;
  assign n33685 = ~pi153 & ~pi766;
  assign n33686 = ~n6654 & n33685;
  assign n33687 = pi39 & ~n33686;
  assign n33688 = ~n33684 & n33687;
  assign n33689 = ~pi153 & ~n59147;
  assign n33690 = ~n12925 & ~n33205;
  assign n33691 = ~n33689 & ~n33690;
  assign n33692 = ~pi38 & ~n33691;
  assign n33693 = ~n33688 & n33692;
  assign n33694 = ~n33666 & ~n33693;
  assign n33695 = ~pi700 & ~n33694;
  assign n33696 = ~n33106 & n33691;
  assign n33697 = pi153 & ~n33151;
  assign n33698 = n33128 & ~n33697;
  assign n33699 = ~n33095 & n33670;
  assign n33700 = ~pi215 & ~n33699;
  assign n33701 = n33674 & n33700;
  assign n33702 = ~n33678 & ~n33701;
  assign n33703 = pi299 & ~n33702;
  assign n33704 = ~n33698 & ~n33703;
  assign n33705 = pi766 & ~n33704;
  assign n33706 = n33097 & ~n33669;
  assign n33707 = ~n33075 & ~n33706;
  assign n33708 = n33674 & n33707;
  assign n33709 = ~pi215 & ~n33708;
  assign n33710 = n33140 & ~n33678;
  assign n33711 = ~n33070 & ~n33710;
  assign n33712 = ~n33709 & n33711;
  assign n33713 = pi299 & ~n33712;
  assign n33714 = n33103 & ~n33667;
  assign n33715 = ~pi766 & ~n33714;
  assign n33716 = ~n33713 & n33715;
  assign n33717 = pi39 & ~n33716;
  assign n33718 = ~n33713 & ~n33714;
  assign n33719 = ~pi766 & ~n33718;
  assign n33720 = pi766 & ~n33703;
  assign n33721 = ~n33698 & n33720;
  assign n33722 = ~n33719 & ~n33721;
  assign n33723 = pi39 & ~n33722;
  assign n33724 = ~n33705 & n33717;
  assign n33725 = ~n33696 & ~n60323;
  assign n33726 = ~pi38 & ~n33725;
  assign n33727 = ~n32944 & ~n33661;
  assign n33728 = ~pi766 & pi947;
  assign n33729 = ~pi39 & ~n33728;
  assign n33730 = n33372 & n33729;
  assign n33731 = n6863 & ~n33727;
  assign n33732 = ~pi153 & ~n6863;
  assign n33733 = pi38 & ~n33732;
  assign n33734 = pi38 & ~n60324;
  assign n33735 = ~n33732 & n33734;
  assign n33736 = ~n60324 & n33733;
  assign n33737 = pi700 & ~n60325;
  assign n33738 = ~n33726 & n33737;
  assign n33739 = ~n33695 & ~n33738;
  assign n33740 = ~n33726 & ~n60325;
  assign n33741 = pi700 & ~n33740;
  assign n33742 = ~pi700 & ~n33666;
  assign n33743 = ~n33693 & n33742;
  assign n33744 = n25257 & ~n33743;
  assign n33745 = ~n33741 & n33744;
  assign n33746 = n25257 & ~n33739;
  assign n33747 = ~pi153 & ~n25257;
  assign n33748 = ~pi57 & ~n33747;
  assign n33749 = ~n60326 & n33748;
  assign n33750 = pi57 & pi153;
  assign n33751 = ~pi832 & ~n33750;
  assign n33752 = ~n33749 & n33751;
  assign n33753 = pi700 & n32944;
  assign n33754 = ~pi700 & ~n33661;
  assign n33755 = ~n33727 & ~n33754;
  assign n33756 = n2794 & ~n33755;
  assign n33757 = n33662 & ~n33753;
  assign n33758 = pi153 & ~n2794;
  assign n33759 = pi832 & ~n33758;
  assign n33760 = ~n60327 & n33759;
  assign n33761 = ~n33752 & ~n33760;
  assign n33762 = ~pi742 & pi947;
  assign n33763 = ~pi704 & n32944;
  assign n33764 = ~n33762 & ~n33763;
  assign n33765 = n2794 & ~n33764;
  assign n33766 = ~pi154 & ~n2794;
  assign n33767 = pi832 & ~n33766;
  assign n33768 = ~n33765 & n33767;
  assign n33769 = ~pi154 & ~n59147;
  assign n33770 = n33107 & ~n33769;
  assign n33771 = ~n33135 & n33770;
  assign n33772 = ~pi154 & ~n60293;
  assign n33773 = pi154 & ~n60297;
  assign n33774 = pi39 & ~n33773;
  assign n33775 = ~n33772 & n33774;
  assign n33776 = ~n33771 & ~n33775;
  assign n33777 = ~pi38 & ~n33776;
  assign n33778 = ~pi154 & ~n6863;
  assign n33779 = n33168 & ~n33778;
  assign n33780 = ~pi742 & ~n33779;
  assign n33781 = ~n33777 & n33780;
  assign n33782 = ~pi154 & n33085;
  assign n33783 = pi154 & n33104;
  assign n33784 = pi39 & ~n33783;
  assign n33785 = ~n33782 & n33784;
  assign n33786 = ~n33770 & ~n33785;
  assign n33787 = ~pi38 & ~n33786;
  assign n33788 = n33114 & ~n33778;
  assign n33789 = pi742 & ~n33788;
  assign n33790 = ~n33787 & n33789;
  assign n33791 = ~pi704 & ~n33790;
  assign n33792 = ~n33781 & n33791;
  assign n33793 = n33205 & ~n33769;
  assign n33794 = ~pi154 & ~n33190;
  assign n33795 = pi154 & n33214;
  assign n33796 = pi39 & ~n33795;
  assign n33797 = ~n33794 & n33796;
  assign n33798 = ~n33793 & ~n33797;
  assign n33799 = ~pi38 & ~n33798;
  assign n33800 = ~n33203 & ~n33778;
  assign n33801 = ~pi742 & ~n33800;
  assign n33802 = ~n33799 & n33801;
  assign n33803 = ~pi154 & pi742;
  assign n33804 = ~n7553 & n33803;
  assign n33805 = pi704 & ~n33804;
  assign n33806 = ~n33802 & n33805;
  assign n33807 = n59928 & ~n33806;
  assign n33808 = ~n33792 & n33807;
  assign n33809 = ~pi154 & ~n59928;
  assign n33810 = ~pi832 & ~n33809;
  assign n33811 = ~n33808 & n33810;
  assign po311 = ~n33768 & ~n33811;
  assign n33813 = ~pi38 & ~n33108;
  assign n33814 = ~n33114 & ~n33813;
  assign n33815 = pi757 & n33814;
  assign n33816 = ~pi38 & ~n33161;
  assign n33817 = ~n33168 & ~n33816;
  assign n33818 = ~pi757 & n33817;
  assign n33819 = ~pi686 & ~n33818;
  assign n33820 = ~pi686 & ~n33815;
  assign n33821 = ~n33818 & n33820;
  assign n33822 = ~n33815 & n33819;
  assign n33823 = ~pi757 & n33218;
  assign n33824 = pi686 & ~n33823;
  assign n33825 = n59928 & ~n33824;
  assign n33826 = ~n60328 & n33825;
  assign n33827 = pi155 & ~n33826;
  assign n33828 = ~pi38 & ~n33089;
  assign n33829 = n24385 & ~n32944;
  assign n33830 = n6863 & n33114;
  assign n33831 = n24385 & n33615;
  assign n33832 = n6468 & n33829;
  assign n33833 = ~n33828 & ~n60329;
  assign n33834 = pi757 & n33833;
  assign n33835 = ~pi38 & ~n33138;
  assign n33836 = pi38 & n33165;
  assign n33837 = ~n33835 & ~n33836;
  assign n33838 = ~pi757 & n33837;
  assign n33839 = ~pi686 & ~n33838;
  assign n33840 = ~pi686 & ~n33834;
  assign n33841 = ~n33838 & n33840;
  assign n33842 = ~n33834 & n33839;
  assign n33843 = ~pi757 & n33196;
  assign n33844 = pi686 & ~n13914;
  assign n33845 = ~n33843 & n33844;
  assign n33846 = ~n60330 & ~n33845;
  assign n33847 = ~pi155 & n59928;
  assign n33848 = ~n33846 & n33847;
  assign n33849 = ~n33827 & ~n33848;
  assign n33850 = ~pi832 & ~n33849;
  assign n33851 = ~pi757 & pi947;
  assign n33852 = ~pi686 & n32944;
  assign n33853 = ~n33851 & ~n33852;
  assign n33854 = n2794 & ~n33853;
  assign n33855 = ~pi155 & ~n2794;
  assign n33856 = pi832 & ~n33855;
  assign n33857 = ~n33854 & n33856;
  assign po312 = ~n33850 & ~n33857;
  assign n33859 = ~pi741 & pi947;
  assign n33860 = ~pi724 & n32944;
  assign n33861 = ~n33859 & ~n33860;
  assign n33862 = n2794 & ~n33861;
  assign n33863 = ~pi156 & ~n2794;
  assign n33864 = pi832 & ~n33863;
  assign n33865 = ~n33862 & n33864;
  assign n33866 = ~pi741 & ~n33837;
  assign n33867 = pi741 & ~n33833;
  assign n33868 = ~pi724 & ~n33867;
  assign n33869 = ~pi724 & ~n33866;
  assign n33870 = ~n33867 & n33869;
  assign n33871 = ~n33866 & n33868;
  assign n33872 = ~pi741 & ~n33196;
  assign n33873 = pi724 & ~n15124;
  assign n33874 = ~n33872 & n33873;
  assign n33875 = n59928 & ~n33874;
  assign n33876 = ~n60331 & n33875;
  assign n33877 = ~pi156 & ~n33876;
  assign n33878 = ~pi741 & ~n33817;
  assign n33879 = pi741 & ~n33814;
  assign n33880 = ~pi724 & ~n33879;
  assign n33881 = ~pi724 & ~n33878;
  assign n33882 = ~n33879 & n33881;
  assign n33883 = ~n33878 & n33880;
  assign n33884 = pi724 & ~pi741;
  assign n33885 = n33218 & n33884;
  assign n33886 = ~n60332 & ~n33885;
  assign n33887 = pi156 & n59928;
  assign n33888 = ~n33886 & n33887;
  assign n33889 = ~pi832 & ~n33888;
  assign n33890 = ~n33877 & n33889;
  assign po313 = ~n33865 & ~n33890;
  assign n33892 = ~pi760 & pi947;
  assign n33893 = ~pi688 & n32944;
  assign n33894 = ~n33892 & ~n33893;
  assign n33895 = n2794 & ~n33894;
  assign n33896 = ~pi157 & ~n2794;
  assign n33897 = pi832 & ~n33896;
  assign n33898 = ~n33895 & n33897;
  assign n33899 = pi760 & ~n33085;
  assign n33900 = ~pi760 & n60293;
  assign n33901 = ~pi157 & ~n33900;
  assign n33902 = ~pi157 & ~n33899;
  assign n33903 = ~n33900 & n33902;
  assign n33904 = ~n33899 & n33901;
  assign n33905 = pi760 & ~n33104;
  assign n33906 = ~pi760 & n60297;
  assign n33907 = pi157 & ~n33906;
  assign n33908 = ~n33905 & n33907;
  assign n33909 = pi39 & ~n33908;
  assign n33910 = pi760 & n33104;
  assign n33911 = ~pi760 & ~n60297;
  assign n33912 = pi157 & ~n33911;
  assign n33913 = ~n33910 & n33912;
  assign n33914 = ~pi760 & ~n60293;
  assign n33915 = pi760 & n33085;
  assign n33916 = ~pi157 & ~n33915;
  assign n33917 = ~n33914 & n33916;
  assign n33918 = ~n33913 & ~n33917;
  assign n33919 = pi39 & ~n33918;
  assign n33920 = ~n60333 & n33909;
  assign n33921 = n59147 & n33892;
  assign n33922 = ~pi157 & ~n59147;
  assign n33923 = ~pi39 & ~n33922;
  assign n33924 = ~pi39 & ~n33921;
  assign n33925 = ~n33922 & n33924;
  assign n33926 = ~n33921 & n33923;
  assign n33927 = ~n33106 & n60335;
  assign n33928 = ~pi38 & ~n33927;
  assign n33929 = ~n60334 & n33928;
  assign n33930 = n6863 & ~n33892;
  assign n33931 = ~n32944 & n33930;
  assign n33932 = pi157 & ~n6863;
  assign n33933 = pi38 & ~n33932;
  assign n33934 = ~n33931 & n33933;
  assign n33935 = ~pi688 & ~n33934;
  assign n33936 = ~n33929 & n33935;
  assign n33937 = ~pi157 & ~n33184;
  assign n33938 = ~n30729 & ~n33213;
  assign n33939 = ~n33937 & ~n33938;
  assign n33940 = ~pi157 & ~n6627;
  assign n33941 = n33206 & ~n33940;
  assign n33942 = ~pi760 & ~n33941;
  assign n33943 = ~n33939 & n33942;
  assign n33944 = ~pi157 & pi760;
  assign n33945 = ~n6654 & n33944;
  assign n33946 = pi39 & ~n33945;
  assign n33947 = ~n33943 & n33946;
  assign n33948 = ~pi38 & ~n60335;
  assign n33949 = ~n33947 & n33948;
  assign n33950 = pi38 & ~n33930;
  assign n33951 = ~n33932 & n33950;
  assign n33952 = pi688 & ~n33951;
  assign n33953 = ~n33949 & n33952;
  assign n33954 = n59928 & ~n33953;
  assign n33955 = ~n33949 & ~n33951;
  assign n33956 = pi688 & ~n33955;
  assign n33957 = ~n60334 & ~n33927;
  assign n33958 = ~pi38 & ~n33957;
  assign n33959 = ~n32944 & ~n33892;
  assign n33960 = pi760 & pi947;
  assign n33961 = ~pi39 & ~n33960;
  assign n33962 = n33372 & n33961;
  assign n33963 = n6863 & ~n33959;
  assign n33964 = ~pi157 & ~n6863;
  assign n33965 = pi38 & ~n33964;
  assign n33966 = ~n60336 & n33965;
  assign n33967 = ~pi688 & ~n33966;
  assign n33968 = ~n33958 & n33967;
  assign n33969 = ~n33956 & ~n33968;
  assign n33970 = n59928 & ~n33969;
  assign n33971 = ~n33936 & n33954;
  assign n33972 = ~pi157 & ~n59928;
  assign n33973 = ~pi832 & ~n33972;
  assign n33974 = ~n60337 & n33973;
  assign po314 = ~n33898 & ~n33974;
  assign n33976 = ~pi753 & pi947;
  assign n33977 = ~n32944 & ~n33976;
  assign n33978 = n2794 & ~n33977;
  assign n33979 = pi702 & ~n33976;
  assign n33980 = ~pi702 & n32944;
  assign n33981 = ~n33976 & ~n33980;
  assign n33982 = n2794 & ~n33981;
  assign n33983 = n33978 & ~n33979;
  assign n33984 = ~pi158 & ~n2794;
  assign n33985 = pi832 & ~n33984;
  assign n33986 = ~n60338 & n33985;
  assign n33987 = ~pi158 & ~n60293;
  assign n33988 = pi158 & ~n60297;
  assign n33989 = ~pi753 & ~n33988;
  assign n33990 = ~n33987 & n33989;
  assign n33991 = ~pi158 & n33085;
  assign n33992 = pi158 & n33104;
  assign n33993 = pi753 & ~n33992;
  assign n33994 = ~n33991 & n33993;
  assign n33995 = pi39 & ~n33994;
  assign n33996 = ~pi158 & ~n33085;
  assign n33997 = pi158 & ~n33104;
  assign n33998 = pi753 & ~n33997;
  assign n33999 = ~n33996 & n33998;
  assign n34000 = ~pi158 & n60293;
  assign n34001 = pi158 & n60297;
  assign n34002 = ~pi753 & ~n34001;
  assign n34003 = ~n34000 & n34002;
  assign n34004 = ~n33999 & ~n34003;
  assign n34005 = pi39 & ~n34004;
  assign n34006 = ~n33990 & n33995;
  assign n34007 = n33087 & ~n33976;
  assign n34008 = pi158 & ~n59147;
  assign n34009 = ~pi39 & ~n34008;
  assign n34010 = ~n34007 & n34009;
  assign n34011 = ~pi38 & ~n34010;
  assign n34012 = ~n60339 & n34011;
  assign n34013 = ~pi158 & ~n6863;
  assign n34014 = pi753 & pi947;
  assign n34015 = ~pi39 & ~n34014;
  assign n34016 = n33372 & n34015;
  assign n34017 = n6863 & ~n33977;
  assign n34018 = n59171 & n33978;
  assign n34019 = pi38 & ~n60340;
  assign n34020 = pi38 & ~n34013;
  assign n34021 = ~n60340 & n34020;
  assign n34022 = ~n34013 & n34019;
  assign n34023 = ~pi702 & ~n60341;
  assign n34024 = ~n34012 & n34023;
  assign n34025 = ~pi158 & n33190;
  assign n34026 = pi158 & ~n33214;
  assign n34027 = ~pi753 & ~n34026;
  assign n34028 = ~n34025 & n34027;
  assign n34029 = ~pi158 & pi753;
  assign n34030 = ~n6654 & n34029;
  assign n34031 = ~n34028 & ~n34030;
  assign n34032 = pi39 & ~n34031;
  assign n34033 = ~n15731 & ~n34008;
  assign n34034 = n33177 & n34033;
  assign n34035 = ~pi38 & ~n34034;
  assign n34036 = ~n34032 & n34035;
  assign n34037 = pi158 & ~n6863;
  assign n34038 = n6863 & ~n33976;
  assign n34039 = ~n34037 & ~n34038;
  assign n34040 = pi38 & ~n34039;
  assign n34041 = pi702 & ~n34040;
  assign n34042 = ~n34036 & n34041;
  assign n34043 = ~n34024 & ~n34042;
  assign n34044 = n59928 & ~n34043;
  assign n34045 = ~pi158 & ~n59928;
  assign n34046 = ~pi832 & ~n34045;
  assign n34047 = ~n34044 & n34046;
  assign po315 = ~n33986 & ~n34047;
  assign n34049 = ~pi754 & pi947;
  assign n34050 = ~n32944 & ~n34049;
  assign n34051 = n2794 & ~n34050;
  assign n34052 = pi709 & ~n34049;
  assign n34053 = ~pi709 & n32944;
  assign n34054 = ~n34049 & ~n34053;
  assign n34055 = n2794 & ~n34054;
  assign n34056 = n34051 & ~n34052;
  assign n34057 = ~pi159 & ~n2794;
  assign n34058 = pi832 & ~n34057;
  assign n34059 = ~n60342 & n34058;
  assign n34060 = ~pi159 & ~n60293;
  assign n34061 = pi159 & ~n60297;
  assign n34062 = ~pi754 & ~n34061;
  assign n34063 = ~n34060 & n34062;
  assign n34064 = ~pi159 & n33085;
  assign n34065 = pi159 & n33104;
  assign n34066 = pi754 & ~n34065;
  assign n34067 = ~n34064 & n34066;
  assign n34068 = pi39 & ~n34067;
  assign n34069 = ~pi159 & ~n33085;
  assign n34070 = pi159 & ~n33104;
  assign n34071 = pi754 & ~n34070;
  assign n34072 = ~n34069 & n34071;
  assign n34073 = ~pi159 & n60293;
  assign n34074 = pi159 & n60297;
  assign n34075 = ~pi754 & ~n34074;
  assign n34076 = ~n34073 & n34075;
  assign n34077 = ~n34072 & ~n34076;
  assign n34078 = pi39 & ~n34077;
  assign n34079 = ~n34063 & n34068;
  assign n34080 = n33087 & ~n34049;
  assign n34081 = pi159 & ~n59147;
  assign n34082 = ~pi39 & ~n34081;
  assign n34083 = ~n34080 & n34082;
  assign n34084 = ~pi38 & ~n34083;
  assign n34085 = ~n60343 & n34084;
  assign n34086 = ~pi159 & ~n6863;
  assign n34087 = pi754 & pi947;
  assign n34088 = ~pi39 & ~n34087;
  assign n34089 = n33372 & n34088;
  assign n34090 = n6863 & ~n34050;
  assign n34091 = n59171 & n34051;
  assign n34092 = pi38 & ~n60344;
  assign n34093 = pi38 & ~n34086;
  assign n34094 = ~n60344 & n34093;
  assign n34095 = ~n34086 & n34092;
  assign n34096 = ~pi709 & ~n60345;
  assign n34097 = ~n34085 & n34096;
  assign n34098 = ~pi159 & n33190;
  assign n34099 = pi159 & ~n33214;
  assign n34100 = ~pi754 & ~n34099;
  assign n34101 = ~n34098 & n34100;
  assign n34102 = ~pi159 & pi754;
  assign n34103 = ~n6654 & n34102;
  assign n34104 = ~n34101 & ~n34103;
  assign n34105 = pi39 & ~n34104;
  assign n34106 = ~n16272 & ~n34081;
  assign n34107 = n33177 & n34106;
  assign n34108 = ~pi38 & ~n34107;
  assign n34109 = ~n34105 & n34108;
  assign n34110 = pi159 & ~n6863;
  assign n34111 = n6863 & ~n34049;
  assign n34112 = ~n34110 & ~n34111;
  assign n34113 = pi38 & ~n34112;
  assign n34114 = pi709 & ~n34113;
  assign n34115 = ~n34109 & n34114;
  assign n34116 = ~n34097 & ~n34115;
  assign n34117 = n59928 & ~n34116;
  assign n34118 = ~pi159 & ~n59928;
  assign n34119 = ~pi832 & ~n34118;
  assign n34120 = ~n34117 & n34119;
  assign po316 = ~n34059 & ~n34120;
  assign n34122 = ~pi756 & pi947;
  assign n34123 = ~pi734 & n32944;
  assign n34124 = ~n34122 & ~n34123;
  assign n34125 = n2794 & ~n34124;
  assign n34126 = ~pi160 & ~n2794;
  assign n34127 = pi832 & ~n34126;
  assign n34128 = ~n34125 & n34127;
  assign n34129 = ~pi160 & n60293;
  assign n34130 = pi160 & n60297;
  assign n34131 = ~pi756 & ~n34130;
  assign n34132 = ~n34129 & n34131;
  assign n34133 = ~pi160 & n33080;
  assign n34134 = pi160 & ~n33236;
  assign n34135 = pi756 & ~n60292;
  assign n34136 = ~n34134 & n34135;
  assign n34137 = ~n34133 & n34136;
  assign n34138 = pi39 & ~n34137;
  assign n34139 = ~n60292 & ~n34134;
  assign n34140 = ~n34133 & n34139;
  assign n34141 = pi756 & ~n34140;
  assign n34142 = ~pi160 & ~n60293;
  assign n34143 = pi160 & ~n60297;
  assign n34144 = ~pi756 & ~n34143;
  assign n34145 = ~n34142 & n34144;
  assign n34146 = ~n34141 & ~n34145;
  assign n34147 = pi39 & ~n34146;
  assign n34148 = ~n34132 & n34138;
  assign n34149 = n59147 & n34122;
  assign n34150 = ~pi160 & ~n59147;
  assign n34151 = ~pi39 & ~n34150;
  assign n34152 = ~pi39 & ~n34149;
  assign n34153 = ~n34150 & n34152;
  assign n34154 = ~n34149 & n34151;
  assign n34155 = ~n33106 & n60347;
  assign n34156 = ~pi38 & ~n34155;
  assign n34157 = ~n60346 & n34156;
  assign n34158 = n6863 & ~n34122;
  assign n34159 = ~n32944 & n34158;
  assign n34160 = pi160 & ~n6863;
  assign n34161 = pi38 & ~n34160;
  assign n34162 = ~n34159 & n34161;
  assign n34163 = ~pi734 & ~n34162;
  assign n34164 = ~n34157 & n34163;
  assign n34165 = ~pi160 & ~n33184;
  assign n34166 = pi160 & ~n33266;
  assign n34167 = pi299 & ~n34166;
  assign n34168 = ~n34165 & n34167;
  assign n34169 = ~pi160 & ~n6627;
  assign n34170 = n33206 & ~n34169;
  assign n34171 = ~pi756 & ~n34170;
  assign n34172 = ~n34168 & n34171;
  assign n34173 = ~pi160 & pi756;
  assign n34174 = ~n6654 & n34173;
  assign n34175 = pi39 & ~n34174;
  assign n34176 = ~n34172 & n34175;
  assign n34177 = ~pi38 & ~n60347;
  assign n34178 = ~n34176 & n34177;
  assign n34179 = pi38 & ~n34158;
  assign n34180 = ~n34160 & n34179;
  assign n34181 = pi734 & ~n34180;
  assign n34182 = ~n34178 & n34181;
  assign n34183 = n59928 & ~n34182;
  assign n34184 = ~n34178 & ~n34180;
  assign n34185 = pi734 & ~n34184;
  assign n34186 = ~n60346 & ~n34155;
  assign n34187 = ~pi38 & ~n34186;
  assign n34188 = ~n32944 & ~n34122;
  assign n34189 = pi756 & pi947;
  assign n34190 = ~pi39 & ~n34189;
  assign n34191 = n33372 & n34190;
  assign n34192 = n6863 & ~n34188;
  assign n34193 = ~pi160 & ~n6863;
  assign n34194 = pi38 & ~n34193;
  assign n34195 = ~n60348 & n34194;
  assign n34196 = ~pi734 & ~n34195;
  assign n34197 = ~n34187 & n34196;
  assign n34198 = ~n34185 & ~n34197;
  assign n34199 = n59928 & ~n34198;
  assign n34200 = ~n34164 & n34183;
  assign n34201 = ~pi160 & ~n59928;
  assign n34202 = ~pi832 & ~n34201;
  assign n34203 = ~n60349 & n34202;
  assign po317 = ~n34128 & ~n34203;
  assign n34205 = pi161 & ~n6464;
  assign n34206 = ~n33141 & ~n34205;
  assign n34207 = n6629 & n34206;
  assign n34208 = ~pi215 & ~n34207;
  assign n34209 = pi161 & n33074;
  assign n34210 = n33094 & ~n34209;
  assign n34211 = ~n6635 & n34210;
  assign n34212 = n34208 & ~n34211;
  assign n34213 = ~pi161 & ~n6645;
  assign n34214 = n33071 & ~n34213;
  assign n34215 = pi299 & ~n34214;
  assign n34216 = ~n34212 & n34215;
  assign n34217 = ~pi161 & ~n59154;
  assign n34218 = n33567 & ~n34217;
  assign n34219 = n33570 & ~n34218;
  assign n34220 = n6544 & n34206;
  assign n34221 = ~pi223 & ~n34220;
  assign n34222 = ~n34219 & n34221;
  assign n34223 = ~pi161 & ~n59150;
  assign n34224 = n33125 & ~n34223;
  assign n34225 = n33123 & ~n34223;
  assign n34226 = ~pi299 & ~n34225;
  assign n34227 = ~n34224 & n34226;
  assign n34228 = ~n34222 & n34227;
  assign n34229 = pi758 & ~n34228;
  assign n34230 = pi758 & ~n34216;
  assign n34231 = ~n34228 & n34230;
  assign n34232 = ~n34216 & n34229;
  assign n34233 = ~n33096 & ~n34205;
  assign n34234 = n6544 & ~n34233;
  assign n34235 = n33588 & ~n34217;
  assign n34236 = ~n34234 & ~n34235;
  assign n34237 = ~pi223 & ~n34236;
  assign n34238 = ~pi299 & ~n34224;
  assign n34239 = ~n34237 & n34238;
  assign n34240 = ~n33072 & n34208;
  assign n34241 = ~n34210 & n34240;
  assign n34242 = ~n33596 & n34214;
  assign n34243 = pi299 & ~n34242;
  assign n34244 = ~n34241 & n34243;
  assign n34245 = ~pi758 & ~n34244;
  assign n34246 = ~n34239 & n34245;
  assign n34247 = pi39 & ~n34246;
  assign n34248 = ~n60350 & n34247;
  assign n34249 = pi758 & pi947;
  assign n34250 = n59147 & n34249;
  assign n34251 = pi161 & ~n59147;
  assign n34252 = ~pi39 & ~n34251;
  assign n34253 = ~pi39 & ~n34250;
  assign n34254 = ~n34251 & n34253;
  assign n34255 = ~n34250 & n34252;
  assign n34256 = ~n33106 & n60351;
  assign n34257 = ~pi38 & ~n34256;
  assign n34258 = ~n34248 & n34257;
  assign n34259 = ~pi39 & ~n34249;
  assign n34260 = n6863 & ~n34249;
  assign n34261 = ~n32944 & n34260;
  assign n34262 = n33615 & n34259;
  assign n34263 = ~pi161 & ~n6863;
  assign n34264 = pi38 & ~n34263;
  assign n34265 = ~n60352 & n34264;
  assign n34266 = pi736 & ~n34265;
  assign n34267 = ~n34258 & n34266;
  assign n34268 = ~n33180 & ~n34210;
  assign n34269 = ~n33073 & ~n34268;
  assign n34270 = ~n33209 & ~n34205;
  assign n34271 = n6629 & n34270;
  assign n34272 = ~pi215 & ~n34271;
  assign n34273 = ~n34269 & n34272;
  assign n34274 = pi161 & n33183;
  assign n34275 = n33207 & ~n34274;
  assign n34276 = ~n34273 & n34275;
  assign n34277 = n6544 & ~n34270;
  assign n34278 = ~n34218 & ~n34277;
  assign n34279 = ~pi223 & ~n34278;
  assign n34280 = n34226 & ~n34279;
  assign n34281 = pi758 & ~n34280;
  assign n34282 = ~n34276 & n34281;
  assign n34283 = pi161 & n10364;
  assign n34284 = pi39 & ~n34283;
  assign n34285 = ~n34282 & n34284;
  assign n34286 = ~pi38 & ~n60351;
  assign n34287 = ~n34285 & n34286;
  assign n34288 = pi38 & ~n34260;
  assign n34289 = ~n34263 & n34288;
  assign n34290 = ~pi736 & ~n34289;
  assign n34291 = ~n34287 & n34290;
  assign n34292 = ~n34267 & ~n34291;
  assign n34293 = n59928 & ~n34292;
  assign n34294 = ~pi161 & ~n59928;
  assign n34295 = ~pi832 & ~n34294;
  assign n34296 = ~n34293 & n34295;
  assign n34297 = pi736 & n32944;
  assign n34298 = n2794 & ~n34249;
  assign n34299 = ~n34297 & n34298;
  assign n34300 = ~pi161 & ~n2794;
  assign n34301 = pi832 & ~n34300;
  assign n34302 = ~n34299 & n34301;
  assign n34303 = ~n34296 & ~n34302;
  assign n34304 = ~pi761 & pi947;
  assign n34305 = ~n32944 & ~n34304;
  assign n34306 = n2794 & ~n34305;
  assign n34307 = pi738 & ~n34304;
  assign n34308 = ~pi738 & n32944;
  assign n34309 = ~n34304 & ~n34308;
  assign n34310 = n2794 & ~n34309;
  assign n34311 = n34306 & ~n34307;
  assign n34312 = ~pi162 & ~n2794;
  assign n34313 = pi832 & ~n34312;
  assign n34314 = ~n60353 & n34313;
  assign n34315 = pi162 & ~n6863;
  assign n34316 = n6863 & ~n34304;
  assign n34317 = pi38 & ~n34316;
  assign n34318 = ~n34315 & n34317;
  assign n34319 = ~pi761 & n33186;
  assign n34320 = pi761 & n6654;
  assign n34321 = ~pi162 & ~n34320;
  assign n34322 = ~n34319 & n34321;
  assign n34323 = pi162 & pi299;
  assign n34324 = ~n33266 & n34323;
  assign n34325 = ~n60299 & ~n34324;
  assign n34326 = ~pi761 & ~n34325;
  assign n34327 = pi39 & ~n34326;
  assign n34328 = ~pi162 & ~n6654;
  assign n34329 = pi761 & ~n34328;
  assign n34330 = ~pi162 & ~n34319;
  assign n34331 = n34325 & ~n34330;
  assign n34332 = ~n34329 & ~n34331;
  assign n34333 = pi39 & ~n34332;
  assign n34334 = ~n34322 & n34327;
  assign n34335 = n59147 & n34304;
  assign n34336 = ~pi162 & ~n59147;
  assign n34337 = ~pi39 & ~n34336;
  assign n34338 = ~pi39 & ~n34335;
  assign n34339 = ~n34336 & n34338;
  assign n34340 = ~n34335 & n34337;
  assign n34341 = ~pi38 & ~n60355;
  assign n34342 = ~n60354 & n34341;
  assign n34343 = ~n34318 & ~n34342;
  assign n34344 = pi738 & ~n34343;
  assign n34345 = ~n33106 & n60355;
  assign n34346 = ~pi162 & n60293;
  assign n34347 = pi162 & n60297;
  assign n34348 = ~pi761 & ~n34347;
  assign n34349 = ~n34346 & n34348;
  assign n34350 = ~n33085 & ~n34323;
  assign n34351 = pi162 & ~n33236;
  assign n34352 = pi761 & ~n34351;
  assign n34353 = ~n34350 & n34352;
  assign n34354 = pi39 & ~n34353;
  assign n34355 = ~n34350 & ~n34351;
  assign n34356 = pi761 & ~n34355;
  assign n34357 = ~pi162 & ~n60293;
  assign n34358 = pi162 & ~n60297;
  assign n34359 = ~pi761 & ~n34358;
  assign n34360 = ~n34357 & n34359;
  assign n34361 = ~n34356 & ~n34360;
  assign n34362 = pi39 & ~n34361;
  assign n34363 = ~n34349 & n34354;
  assign n34364 = ~n34345 & ~n60356;
  assign n34365 = ~pi38 & ~n34364;
  assign n34366 = ~pi162 & ~n6863;
  assign n34367 = pi761 & pi947;
  assign n34368 = ~pi39 & ~n34367;
  assign n34369 = n33372 & n34368;
  assign n34370 = n6863 & ~n34305;
  assign n34371 = n59171 & n34306;
  assign n34372 = pi38 & ~n60357;
  assign n34373 = pi38 & ~n34366;
  assign n34374 = ~n60357 & n34373;
  assign n34375 = ~n34366 & n34372;
  assign n34376 = ~pi738 & ~n60358;
  assign n34377 = ~n34365 & n34376;
  assign n34378 = ~n34344 & ~n34377;
  assign n34379 = n59928 & ~n34378;
  assign n34380 = ~pi162 & ~n59928;
  assign n34381 = ~pi832 & ~n34380;
  assign n34382 = ~n34379 & n34381;
  assign po319 = ~n34314 & ~n34382;
  assign n34384 = ~pi777 & pi947;
  assign n34385 = ~pi737 & n32944;
  assign n34386 = ~n34384 & ~n34385;
  assign n34387 = n2794 & ~n34386;
  assign n34388 = ~pi163 & ~n2794;
  assign n34389 = pi832 & ~n34388;
  assign n34390 = ~n34387 & n34389;
  assign n34391 = ~pi163 & n60293;
  assign n34392 = pi163 & n60297;
  assign n34393 = ~pi777 & ~n34392;
  assign n34394 = ~n34391 & n34393;
  assign n34395 = ~pi163 & n33080;
  assign n34396 = pi163 & ~n33236;
  assign n34397 = pi777 & ~n60292;
  assign n34398 = ~n34396 & n34397;
  assign n34399 = ~n34395 & n34398;
  assign n34400 = pi39 & ~n34399;
  assign n34401 = ~n60292 & ~n34396;
  assign n34402 = ~n34395 & n34401;
  assign n34403 = pi777 & ~n34402;
  assign n34404 = ~pi163 & ~n60293;
  assign n34405 = pi163 & ~n60297;
  assign n34406 = ~pi777 & ~n34405;
  assign n34407 = ~n34404 & n34406;
  assign n34408 = ~n34403 & ~n34407;
  assign n34409 = pi39 & ~n34408;
  assign n34410 = ~n34394 & n34400;
  assign n34411 = n59147 & n34384;
  assign n34412 = ~pi163 & ~n59147;
  assign n34413 = ~pi39 & ~n34412;
  assign n34414 = ~pi39 & ~n34411;
  assign n34415 = ~n34412 & n34414;
  assign n34416 = ~n34411 & n34413;
  assign n34417 = ~n33106 & n60360;
  assign n34418 = ~pi38 & ~n34417;
  assign n34419 = ~n60359 & n34418;
  assign n34420 = n6863 & ~n34384;
  assign n34421 = ~n32944 & n34420;
  assign n34422 = pi163 & ~n6863;
  assign n34423 = pi38 & ~n34422;
  assign n34424 = ~n34421 & n34423;
  assign n34425 = ~pi737 & ~n34424;
  assign n34426 = ~n34419 & n34425;
  assign n34427 = ~pi163 & ~n33184;
  assign n34428 = ~pi163 & pi299;
  assign n34429 = ~n33213 & ~n34428;
  assign n34430 = ~n34427 & ~n34429;
  assign n34431 = ~pi163 & ~n6627;
  assign n34432 = n33206 & ~n34431;
  assign n34433 = ~pi777 & ~n34432;
  assign n34434 = ~n34430 & n34433;
  assign n34435 = ~pi163 & pi777;
  assign n34436 = ~n6654 & n34435;
  assign n34437 = pi39 & ~n34436;
  assign n34438 = ~n34434 & n34437;
  assign n34439 = ~pi38 & ~n60360;
  assign n34440 = ~n34438 & n34439;
  assign n34441 = pi38 & ~n34420;
  assign n34442 = ~n34422 & n34441;
  assign n34443 = pi737 & ~n34442;
  assign n34444 = ~n34440 & n34443;
  assign n34445 = n59928 & ~n34444;
  assign n34446 = ~n34440 & ~n34442;
  assign n34447 = pi737 & ~n34446;
  assign n34448 = ~n60359 & ~n34417;
  assign n34449 = ~pi38 & ~n34448;
  assign n34450 = ~n32944 & ~n34384;
  assign n34451 = pi777 & pi947;
  assign n34452 = ~pi39 & ~n34451;
  assign n34453 = n33372 & n34452;
  assign n34454 = n6863 & ~n34450;
  assign n34455 = ~pi163 & ~n6863;
  assign n34456 = pi38 & ~n34455;
  assign n34457 = ~n60361 & n34456;
  assign n34458 = ~pi737 & ~n34457;
  assign n34459 = ~n34449 & n34458;
  assign n34460 = ~n34447 & ~n34459;
  assign n34461 = n59928 & ~n34460;
  assign n34462 = ~n34426 & n34445;
  assign n34463 = ~pi163 & ~n59928;
  assign n34464 = ~pi832 & ~n34463;
  assign n34465 = ~n60362 & n34464;
  assign po320 = ~n34390 & ~n34465;
  assign n34467 = ~pi752 & pi947;
  assign n34468 = pi703 & n32944;
  assign n34469 = ~n34467 & ~n34468;
  assign n34470 = n2794 & ~n34469;
  assign n34471 = ~pi164 & ~n2794;
  assign n34472 = pi832 & ~n34471;
  assign n34473 = ~n34470 & n34472;
  assign n34474 = ~pi164 & n33138;
  assign n34475 = pi164 & n33161;
  assign n34476 = ~pi38 & ~n34475;
  assign n34477 = ~n34474 & n34476;
  assign n34478 = ~pi164 & ~n33165;
  assign n34479 = n33168 & ~n34478;
  assign n34480 = ~pi752 & ~n34479;
  assign n34481 = ~n34477 & n34480;
  assign n34482 = ~pi164 & n33089;
  assign n34483 = pi164 & n33108;
  assign n34484 = ~pi38 & ~n34483;
  assign n34485 = ~n34482 & n34484;
  assign n34486 = ~pi164 & ~n6863;
  assign n34487 = n33114 & ~n34486;
  assign n34488 = pi752 & ~n34487;
  assign n34489 = ~n34485 & n34488;
  assign n34490 = ~n34481 & ~n34489;
  assign n34491 = pi703 & ~n34490;
  assign n34492 = pi164 & ~n33195;
  assign n34493 = ~pi752 & ~n34492;
  assign n34494 = ~n33196 & n34493;
  assign n34495 = ~pi164 & ~n7553;
  assign n34496 = pi752 & ~n34495;
  assign n34497 = pi164 & ~n33218;
  assign n34498 = ~pi703 & ~n34497;
  assign n34499 = ~pi752 & n33218;
  assign n34500 = pi164 & ~n34499;
  assign n34501 = pi752 & n7553;
  assign n34502 = ~pi703 & ~n34501;
  assign n34503 = ~n34500 & n34502;
  assign n34504 = ~n34496 & n34498;
  assign n34505 = ~n34494 & n60363;
  assign n34506 = ~n34491 & ~n34505;
  assign n34507 = n59928 & ~n34506;
  assign n34508 = ~pi164 & ~n59928;
  assign n34509 = ~pi832 & ~n34508;
  assign n34510 = ~n34507 & n34509;
  assign po321 = ~n34473 & ~n34510;
  assign n34512 = ~pi774 & pi947;
  assign n34513 = pi687 & n32944;
  assign n34514 = ~n34512 & ~n34513;
  assign n34515 = n2794 & ~n34514;
  assign n34516 = ~pi165 & ~n2794;
  assign n34517 = pi832 & ~n34516;
  assign n34518 = ~n34515 & n34517;
  assign n34519 = ~pi165 & n33138;
  assign n34520 = pi165 & n33161;
  assign n34521 = ~pi38 & ~n34520;
  assign n34522 = ~n34519 & n34521;
  assign n34523 = ~pi165 & ~n33165;
  assign n34524 = n33168 & ~n34523;
  assign n34525 = ~pi774 & ~n34524;
  assign n34526 = ~n34522 & n34525;
  assign n34527 = ~pi165 & n33089;
  assign n34528 = pi165 & n33108;
  assign n34529 = ~pi38 & ~n34528;
  assign n34530 = ~n34527 & n34529;
  assign n34531 = ~pi165 & ~n6863;
  assign n34532 = n33114 & ~n34531;
  assign n34533 = pi774 & ~n34532;
  assign n34534 = ~n34530 & n34533;
  assign n34535 = ~n34526 & ~n34534;
  assign n34536 = pi687 & ~n34535;
  assign n34537 = pi165 & ~n33195;
  assign n34538 = ~pi774 & ~n34537;
  assign n34539 = ~n33196 & n34538;
  assign n34540 = ~pi165 & ~n7553;
  assign n34541 = pi774 & ~n34540;
  assign n34542 = pi165 & ~n33218;
  assign n34543 = ~pi687 & ~n34542;
  assign n34544 = ~pi774 & n33218;
  assign n34545 = pi165 & ~n34544;
  assign n34546 = pi774 & n7553;
  assign n34547 = ~pi687 & ~n34546;
  assign n34548 = ~n34545 & n34547;
  assign n34549 = ~n34541 & n34543;
  assign n34550 = ~n34539 & n60364;
  assign n34551 = ~n34536 & ~n34550;
  assign n34552 = n59928 & ~n34551;
  assign n34553 = ~pi165 & ~n59928;
  assign n34554 = ~pi832 & ~n34553;
  assign n34555 = ~n34552 & n34554;
  assign po322 = ~n34518 & ~n34555;
  assign n34557 = pi166 & ~n6464;
  assign n34558 = ~n33141 & ~n34557;
  assign n34559 = n6629 & n34558;
  assign n34560 = ~pi215 & ~n34559;
  assign n34561 = pi166 & n33074;
  assign n34562 = n33094 & ~n34561;
  assign n34563 = ~n6635 & n34562;
  assign n34564 = n34560 & ~n34563;
  assign n34565 = ~pi166 & ~n6645;
  assign n34566 = n33071 & ~n34565;
  assign n34567 = pi299 & ~n34566;
  assign n34568 = ~n34564 & n34567;
  assign n34569 = n6544 & n34558;
  assign n34570 = ~pi223 & ~n34569;
  assign n34571 = ~pi166 & ~n59154;
  assign n34572 = ~n33587 & ~n34571;
  assign n34573 = n33570 & ~n34572;
  assign n34574 = n34570 & ~n34573;
  assign n34575 = ~n2840 & n59150;
  assign n34576 = ~pi166 & ~n34575;
  assign n34577 = n33125 & ~n34576;
  assign n34578 = ~pi299 & ~n34577;
  assign n34579 = ~pi166 & ~n59150;
  assign n34580 = n33123 & ~n34579;
  assign n34581 = ~pi299 & ~n34580;
  assign n34582 = ~n34577 & n34581;
  assign n34583 = n34578 & ~n34580;
  assign n34584 = ~n34574 & n60365;
  assign n34585 = pi772 & ~n34584;
  assign n34586 = ~n34568 & n34585;
  assign n34587 = ~n33072 & n34560;
  assign n34588 = ~n34562 & n34587;
  assign n34589 = ~n33596 & n34566;
  assign n34590 = pi299 & ~n34589;
  assign n34591 = ~n34588 & n34590;
  assign n34592 = ~n6544 & ~n34572;
  assign n34593 = pi947 & n59155;
  assign n34594 = n6544 & n33209;
  assign n34595 = n34570 & ~n60366;
  assign n34596 = ~n34592 & n34595;
  assign n34597 = n34578 & ~n34596;
  assign n34598 = ~pi772 & ~n34597;
  assign n34599 = ~n34591 & n34598;
  assign n34600 = pi39 & ~n34599;
  assign n34601 = pi39 & ~n34586;
  assign n34602 = ~n34599 & n34601;
  assign n34603 = ~n34586 & n34600;
  assign n34604 = pi772 & pi947;
  assign n34605 = n59147 & n34604;
  assign n34606 = pi166 & ~n59147;
  assign n34607 = ~pi39 & ~n34606;
  assign n34608 = ~pi39 & ~n34604;
  assign n34609 = ~n6459 & ~n34608;
  assign n34610 = ~n34606 & ~n34609;
  assign n34611 = ~n34605 & n34607;
  assign n34612 = ~n33106 & n60368;
  assign n34613 = ~pi38 & ~n34612;
  assign n34614 = ~n60367 & n34613;
  assign n34615 = n2794 & ~n34604;
  assign n34616 = n6863 & ~n34604;
  assign n34617 = n59171 & n34615;
  assign n34618 = n33615 & n34608;
  assign n34619 = ~n32944 & n60369;
  assign n34620 = ~pi166 & ~n6863;
  assign n34621 = pi38 & ~n34620;
  assign n34622 = pi38 & ~n60370;
  assign n34623 = ~n34620 & n34622;
  assign n34624 = ~n60370 & n34621;
  assign n34625 = pi727 & ~n60371;
  assign n34626 = ~n34614 & n34625;
  assign n34627 = ~n33180 & ~n34562;
  assign n34628 = ~n33073 & ~n34627;
  assign n34629 = ~n33209 & ~n34557;
  assign n34630 = n6629 & n34629;
  assign n34631 = ~pi215 & ~n34630;
  assign n34632 = ~n34628 & n34631;
  assign n34633 = pi166 & n33183;
  assign n34634 = n33207 & ~n34633;
  assign n34635 = ~n34632 & n34634;
  assign n34636 = n6544 & ~n34629;
  assign n34637 = n33567 & ~n34571;
  assign n34638 = ~n34636 & ~n34637;
  assign n34639 = ~pi223 & ~n34638;
  assign n34640 = n34581 & ~n34639;
  assign n34641 = pi772 & ~n34640;
  assign n34642 = ~n34635 & n34641;
  assign n34643 = pi166 & n20623;
  assign n34644 = pi39 & ~n34643;
  assign n34645 = ~n34642 & n34644;
  assign n34646 = ~pi38 & ~n60368;
  assign n34647 = ~n34645 & n34646;
  assign n34648 = pi38 & ~n60369;
  assign n34649 = ~n34620 & n34648;
  assign n34650 = ~pi727 & ~n34649;
  assign n34651 = ~n34647 & n34650;
  assign n34652 = ~n34626 & ~n34651;
  assign n34653 = n59928 & ~n34652;
  assign n34654 = ~pi166 & ~n59928;
  assign n34655 = ~pi832 & ~n34654;
  assign n34656 = ~n34653 & n34655;
  assign n34657 = pi727 & n32944;
  assign n34658 = n34615 & ~n34657;
  assign n34659 = ~pi166 & ~n2794;
  assign n34660 = pi832 & ~n34659;
  assign n34661 = ~n34658 & n34660;
  assign n34662 = ~n34656 & ~n34661;
  assign n34663 = ~pi768 & pi947;
  assign n34664 = pi705 & n32944;
  assign n34665 = ~n34663 & ~n34664;
  assign n34666 = n2794 & ~n34665;
  assign n34667 = ~pi167 & ~n2794;
  assign n34668 = pi832 & ~n34667;
  assign n34669 = ~n34666 & n34668;
  assign n34670 = ~pi167 & n33138;
  assign n34671 = pi167 & n33161;
  assign n34672 = ~pi38 & ~n34671;
  assign n34673 = ~n34670 & n34672;
  assign n34674 = ~pi167 & ~n33165;
  assign n34675 = n33168 & ~n34674;
  assign n34676 = ~pi768 & ~n34675;
  assign n34677 = ~n34673 & n34676;
  assign n34678 = ~pi167 & n33089;
  assign n34679 = pi167 & n33108;
  assign n34680 = ~pi38 & ~n34679;
  assign n34681 = ~n34678 & n34680;
  assign n34682 = ~pi167 & ~n6863;
  assign n34683 = n33114 & ~n34682;
  assign n34684 = pi768 & ~n34683;
  assign n34685 = ~n34681 & n34684;
  assign n34686 = pi705 & ~n34685;
  assign n34687 = pi705 & ~n34677;
  assign n34688 = ~n34685 & n34687;
  assign n34689 = ~n34677 & n34686;
  assign n34690 = ~pi167 & ~n33192;
  assign n34691 = pi167 & n33216;
  assign n34692 = ~pi38 & ~n34691;
  assign n34693 = ~n34690 & n34692;
  assign n34694 = ~n33203 & ~n34682;
  assign n34695 = ~pi768 & ~n34694;
  assign n34696 = ~n34693 & n34695;
  assign n34697 = ~pi167 & pi768;
  assign n34698 = ~pi167 & n20066;
  assign n34699 = ~n7553 & n34697;
  assign n34700 = ~pi705 & ~n60373;
  assign n34701 = ~n34696 & n34700;
  assign n34702 = n59928 & ~n34701;
  assign n34703 = ~n60372 & n34702;
  assign n34704 = ~pi167 & ~n59928;
  assign n34705 = ~pi832 & ~n34704;
  assign n34706 = ~n34703 & n34705;
  assign po324 = ~n34669 & ~n34706;
  assign n34708 = pi168 & ~n6863;
  assign n34709 = pi763 & pi947;
  assign n34710 = n2794 & ~n34709;
  assign n34711 = n6863 & ~n34709;
  assign n34712 = n59171 & n34710;
  assign n34713 = pi38 & ~n60374;
  assign n34714 = ~n34708 & n34713;
  assign n34715 = ~pi168 & ~n6627;
  assign n34716 = n33206 & ~n34715;
  assign n34717 = ~pi168 & ~n6464;
  assign n34718 = n33210 & ~n34717;
  assign n34719 = pi168 & ~n6629;
  assign n34720 = pi168 & n6640;
  assign n34721 = ~n6635 & n34719;
  assign n34722 = ~n6634 & ~n60375;
  assign n34723 = ~n34718 & n34722;
  assign n34724 = n33181 & n34723;
  assign n34725 = pi168 & ~n6645;
  assign n34726 = n33071 & ~n34725;
  assign n34727 = ~n33091 & n34726;
  assign n34728 = n33183 & ~n34725;
  assign n34729 = pi299 & ~n60376;
  assign n34730 = ~n34724 & n34729;
  assign n34731 = pi763 & ~n34730;
  assign n34732 = ~n34716 & n34731;
  assign n34733 = ~pi168 & ~pi763;
  assign n34734 = ~n6654 & n34733;
  assign n34735 = pi39 & ~n34734;
  assign n34736 = ~n34732 & n34735;
  assign n34737 = ~pi168 & ~n59147;
  assign n34738 = ~n21316 & ~n33205;
  assign n34739 = ~n34737 & ~n34738;
  assign n34740 = ~pi38 & ~n34739;
  assign n34741 = ~n34736 & n34740;
  assign n34742 = ~n34714 & ~n34741;
  assign n34743 = ~pi699 & ~n34742;
  assign n34744 = ~n33106 & n34739;
  assign n34745 = pi168 & ~n33151;
  assign n34746 = n33128 & ~n34745;
  assign n34747 = ~n33095 & n34718;
  assign n34748 = ~pi215 & ~n34747;
  assign n34749 = n34722 & n34748;
  assign n34750 = ~n34726 & ~n34749;
  assign n34751 = pi299 & ~n34750;
  assign n34752 = ~n34746 & ~n34751;
  assign n34753 = pi763 & ~n34752;
  assign n34754 = n33097 & ~n34717;
  assign n34755 = ~n33075 & ~n34754;
  assign n34756 = n34722 & n34755;
  assign n34757 = ~pi215 & ~n34756;
  assign n34758 = n33140 & ~n34726;
  assign n34759 = ~n33070 & ~n34758;
  assign n34760 = ~n34757 & n34759;
  assign n34761 = pi299 & ~n34760;
  assign n34762 = n33103 & ~n34715;
  assign n34763 = ~pi763 & ~n34762;
  assign n34764 = ~n34761 & n34763;
  assign n34765 = pi39 & ~n34764;
  assign n34766 = ~n34761 & ~n34762;
  assign n34767 = ~pi763 & ~n34766;
  assign n34768 = pi763 & ~n34751;
  assign n34769 = ~n34746 & n34768;
  assign n34770 = ~n34767 & ~n34769;
  assign n34771 = pi39 & ~n34770;
  assign n34772 = ~n34753 & n34765;
  assign n34773 = ~n34744 & ~n60377;
  assign n34774 = ~pi38 & ~n34773;
  assign n34775 = ~n32944 & ~n34709;
  assign n34776 = ~pi763 & pi947;
  assign n34777 = ~pi39 & ~n34776;
  assign n34778 = n33372 & n34777;
  assign n34779 = n6863 & ~n34775;
  assign n34780 = ~pi168 & ~n6863;
  assign n34781 = pi38 & ~n34780;
  assign n34782 = pi38 & ~n60378;
  assign n34783 = ~n34780 & n34782;
  assign n34784 = ~n60378 & n34781;
  assign n34785 = pi699 & ~n60379;
  assign n34786 = ~n34774 & n34785;
  assign n34787 = ~n34743 & ~n34786;
  assign n34788 = ~n34774 & ~n60379;
  assign n34789 = pi699 & ~n34788;
  assign n34790 = ~pi699 & ~n34714;
  assign n34791 = ~n34741 & n34790;
  assign n34792 = n25257 & ~n34791;
  assign n34793 = ~n34789 & n34792;
  assign n34794 = n25257 & ~n34787;
  assign n34795 = ~pi168 & ~n25257;
  assign n34796 = ~pi57 & ~n34795;
  assign n34797 = ~n60380 & n34796;
  assign n34798 = pi57 & pi168;
  assign n34799 = ~pi832 & ~n34798;
  assign n34800 = ~n34797 & n34799;
  assign n34801 = pi699 & n32944;
  assign n34802 = ~pi699 & ~n34709;
  assign n34803 = ~n34775 & ~n34802;
  assign n34804 = n2794 & ~n34803;
  assign n34805 = n34710 & ~n34801;
  assign n34806 = pi168 & ~n2794;
  assign n34807 = pi832 & ~n34806;
  assign n34808 = ~n60381 & n34807;
  assign n34809 = ~n34800 & ~n34808;
  assign n34810 = pi169 & ~n6863;
  assign n34811 = pi746 & pi947;
  assign n34812 = n2794 & ~n34811;
  assign n34813 = n6863 & ~n34811;
  assign n34814 = n59171 & n34812;
  assign n34815 = pi38 & ~n60382;
  assign n34816 = ~n34810 & n34815;
  assign n34817 = ~pi169 & ~n6627;
  assign n34818 = n33206 & ~n34817;
  assign n34819 = ~pi169 & ~n6464;
  assign n34820 = n33210 & ~n34819;
  assign n34821 = pi169 & ~n6629;
  assign n34822 = pi169 & n6640;
  assign n34823 = ~n6635 & n34821;
  assign n34824 = ~n6634 & ~n60383;
  assign n34825 = ~n34820 & n34824;
  assign n34826 = n33181 & n34825;
  assign n34827 = pi169 & ~n6645;
  assign n34828 = n33071 & ~n34827;
  assign n34829 = ~n33091 & n34828;
  assign n34830 = n33183 & ~n34827;
  assign n34831 = pi299 & ~n60384;
  assign n34832 = ~n34826 & n34831;
  assign n34833 = pi746 & ~n34832;
  assign n34834 = ~n34818 & n34833;
  assign n34835 = ~pi169 & ~pi746;
  assign n34836 = ~n6654 & n34835;
  assign n34837 = pi39 & ~n34836;
  assign n34838 = ~n34834 & n34837;
  assign n34839 = ~pi169 & ~n59147;
  assign n34840 = ~n21865 & ~n33205;
  assign n34841 = ~n34839 & ~n34840;
  assign n34842 = ~pi38 & ~n34841;
  assign n34843 = ~n34838 & n34842;
  assign n34844 = ~n34816 & ~n34843;
  assign n34845 = ~pi729 & ~n34844;
  assign n34846 = ~n33106 & n34841;
  assign n34847 = pi169 & ~n33151;
  assign n34848 = n33128 & ~n34847;
  assign n34849 = ~n33095 & n34820;
  assign n34850 = ~pi215 & ~n34849;
  assign n34851 = n34824 & n34850;
  assign n34852 = ~n34828 & ~n34851;
  assign n34853 = pi299 & ~n34852;
  assign n34854 = ~n34848 & ~n34853;
  assign n34855 = pi746 & ~n34854;
  assign n34856 = n33097 & ~n34819;
  assign n34857 = ~n33075 & ~n34856;
  assign n34858 = n34824 & n34857;
  assign n34859 = ~pi215 & ~n34858;
  assign n34860 = n33140 & ~n34828;
  assign n34861 = ~n33070 & ~n34860;
  assign n34862 = ~n34859 & n34861;
  assign n34863 = pi299 & ~n34862;
  assign n34864 = n33103 & ~n34817;
  assign n34865 = ~pi746 & ~n34864;
  assign n34866 = ~n34863 & n34865;
  assign n34867 = pi39 & ~n34866;
  assign n34868 = ~n34863 & ~n34864;
  assign n34869 = ~pi746 & ~n34868;
  assign n34870 = pi746 & ~n34853;
  assign n34871 = ~n34848 & n34870;
  assign n34872 = ~n34869 & ~n34871;
  assign n34873 = pi39 & ~n34872;
  assign n34874 = ~n34855 & n34867;
  assign n34875 = ~n34846 & ~n60385;
  assign n34876 = ~pi38 & ~n34875;
  assign n34877 = ~n32944 & ~n34811;
  assign n34878 = ~pi746 & pi947;
  assign n34879 = ~pi39 & ~n34878;
  assign n34880 = n33372 & n34879;
  assign n34881 = n6863 & ~n34877;
  assign n34882 = ~pi169 & ~n6863;
  assign n34883 = pi38 & ~n34882;
  assign n34884 = pi38 & ~n60386;
  assign n34885 = ~n34882 & n34884;
  assign n34886 = ~n60386 & n34883;
  assign n34887 = pi729 & ~n60387;
  assign n34888 = ~n34876 & n34887;
  assign n34889 = ~n34845 & ~n34888;
  assign n34890 = ~n34876 & ~n60387;
  assign n34891 = pi729 & ~n34890;
  assign n34892 = ~pi729 & ~n34816;
  assign n34893 = ~n34843 & n34892;
  assign n34894 = n25257 & ~n34893;
  assign n34895 = ~n34891 & n34894;
  assign n34896 = n25257 & ~n34889;
  assign n34897 = ~pi169 & ~n25257;
  assign n34898 = ~pi57 & ~n34897;
  assign n34899 = ~n60388 & n34898;
  assign n34900 = pi57 & pi169;
  assign n34901 = ~pi832 & ~n34900;
  assign n34902 = ~n34899 & n34901;
  assign n34903 = pi729 & n32944;
  assign n34904 = ~pi729 & ~n34811;
  assign n34905 = ~n34877 & ~n34904;
  assign n34906 = n2794 & ~n34905;
  assign n34907 = n34812 & ~n34903;
  assign n34908 = pi169 & ~n2794;
  assign n34909 = pi832 & ~n34908;
  assign n34910 = ~n60389 & n34909;
  assign n34911 = ~n34902 & ~n34910;
  assign n34912 = pi730 & n32944;
  assign n34913 = pi748 & pi947;
  assign n34914 = n2794 & ~n34913;
  assign n34915 = ~n34912 & n34914;
  assign n34916 = pi170 & ~n2794;
  assign n34917 = pi832 & ~n34916;
  assign n34918 = ~n34915 & n34917;
  assign n34919 = pi170 & ~n6629;
  assign n34920 = pi170 & n6640;
  assign n34921 = ~n6635 & n34919;
  assign n34922 = ~n6634 & ~n60390;
  assign n34923 = ~pi170 & ~n6464;
  assign n34924 = n33097 & ~n34923;
  assign n34925 = ~n33075 & ~n34924;
  assign n34926 = n34922 & n34925;
  assign n34927 = ~pi215 & ~n34926;
  assign n34928 = pi170 & ~n6645;
  assign n34929 = n33071 & ~n34928;
  assign n34930 = n33140 & ~n34929;
  assign n34931 = ~n33070 & ~n34930;
  assign n34932 = ~n34927 & n34931;
  assign n34933 = pi299 & ~n34932;
  assign n34934 = ~pi170 & ~n6627;
  assign n34935 = ~pi299 & ~n34934;
  assign n34936 = ~n33102 & n34935;
  assign n34937 = ~n34933 & ~n34936;
  assign n34938 = pi39 & ~n34937;
  assign n34939 = ~pi170 & ~n59147;
  assign n34940 = n33107 & ~n34939;
  assign n34941 = ~n34938 & ~n34940;
  assign n34942 = ~pi38 & ~n34941;
  assign n34943 = ~pi170 & ~n6863;
  assign n34944 = n33114 & ~n34943;
  assign n34945 = ~pi748 & ~n34944;
  assign n34946 = ~n34942 & n34945;
  assign n34947 = n33136 & ~n34939;
  assign n34948 = pi170 & ~n33151;
  assign n34949 = n33128 & ~n34948;
  assign n34950 = n33210 & ~n34923;
  assign n34951 = ~n33095 & n34950;
  assign n34952 = ~pi215 & ~n34951;
  assign n34953 = n34922 & n34952;
  assign n34954 = ~n34929 & ~n34953;
  assign n34955 = pi299 & ~n34954;
  assign n34956 = pi39 & ~n34955;
  assign n34957 = ~n34949 & n34956;
  assign n34958 = ~n34947 & ~n34957;
  assign n34959 = ~pi38 & ~n34958;
  assign n34960 = n33168 & ~n34943;
  assign n34961 = pi748 & ~n34960;
  assign n34962 = ~n34959 & n34961;
  assign n34963 = pi730 & ~n34962;
  assign n34964 = ~n34946 & n34963;
  assign n34965 = n33205 & ~n34939;
  assign n34966 = n34922 & ~n34950;
  assign n34967 = n33181 & n34966;
  assign n34968 = n33183 & ~n34928;
  assign n34969 = ~n33091 & n34929;
  assign n34970 = pi299 & ~n60391;
  assign n34971 = ~n34967 & n34970;
  assign n34972 = ~n33187 & n34935;
  assign n34973 = ~n34971 & ~n34972;
  assign n34974 = pi39 & ~n34973;
  assign n34975 = ~n34965 & ~n34974;
  assign n34976 = ~pi38 & ~n34975;
  assign n34977 = ~n33203 & ~n34943;
  assign n34978 = pi748 & ~n34977;
  assign n34979 = ~n34976 & n34978;
  assign n34980 = ~pi170 & ~pi748;
  assign n34981 = ~n7553 & n34980;
  assign n34982 = ~pi730 & ~n34981;
  assign n34983 = ~n34979 & n34982;
  assign n34984 = n25257 & ~n34983;
  assign n34985 = ~n34964 & n34984;
  assign n34986 = ~pi170 & ~n25257;
  assign n34987 = ~pi57 & ~n34986;
  assign n34988 = ~n34985 & n34987;
  assign n34989 = pi57 & pi170;
  assign n34990 = ~pi832 & ~n34989;
  assign n34991 = ~n34988 & n34990;
  assign n34992 = ~n34918 & ~n34991;
  assign n34993 = pi171 & ~n6863;
  assign n34994 = pi764 & pi947;
  assign n34995 = n2794 & ~n34994;
  assign n34996 = n6863 & ~n34994;
  assign n34997 = n59171 & n34995;
  assign n34998 = pi38 & ~n60392;
  assign n34999 = ~n34993 & n34998;
  assign n35000 = ~pi171 & ~n6627;
  assign n35001 = n33206 & ~n35000;
  assign n35002 = ~pi171 & ~n6464;
  assign n35003 = n33210 & ~n35002;
  assign n35004 = pi171 & ~n6629;
  assign n35005 = pi171 & n6640;
  assign n35006 = ~n6635 & n35004;
  assign n35007 = ~n6634 & ~n60393;
  assign n35008 = ~n35003 & n35007;
  assign n35009 = n33181 & n35008;
  assign n35010 = pi171 & ~n6645;
  assign n35011 = n33071 & ~n35010;
  assign n35012 = ~n33091 & n35011;
  assign n35013 = n33183 & ~n35010;
  assign n35014 = pi299 & ~n60394;
  assign n35015 = ~n35009 & n35014;
  assign n35016 = pi764 & ~n35015;
  assign n35017 = ~n35001 & n35016;
  assign n35018 = ~pi171 & ~pi764;
  assign n35019 = ~n6654 & n35018;
  assign n35020 = pi39 & ~n35019;
  assign n35021 = ~n35017 & n35020;
  assign n35022 = ~pi171 & ~n59147;
  assign n35023 = ~n22414 & ~n33205;
  assign n35024 = ~n35022 & ~n35023;
  assign n35025 = ~pi38 & ~n35024;
  assign n35026 = ~n35021 & n35025;
  assign n35027 = ~n34999 & ~n35026;
  assign n35028 = ~pi691 & ~n35027;
  assign n35029 = ~n33106 & n35024;
  assign n35030 = pi171 & ~n33151;
  assign n35031 = n33128 & ~n35030;
  assign n35032 = ~n33095 & n35003;
  assign n35033 = ~pi215 & ~n35032;
  assign n35034 = n35007 & n35033;
  assign n35035 = ~n35011 & ~n35034;
  assign n35036 = pi299 & ~n35035;
  assign n35037 = ~n35031 & ~n35036;
  assign n35038 = pi764 & ~n35037;
  assign n35039 = n33097 & ~n35002;
  assign n35040 = ~n33075 & ~n35039;
  assign n35041 = n35007 & n35040;
  assign n35042 = ~pi215 & ~n35041;
  assign n35043 = n33140 & ~n35011;
  assign n35044 = ~n33070 & ~n35043;
  assign n35045 = ~n35042 & n35044;
  assign n35046 = pi299 & ~n35045;
  assign n35047 = n33103 & ~n35000;
  assign n35048 = ~pi764 & ~n35047;
  assign n35049 = ~n35046 & n35048;
  assign n35050 = pi39 & ~n35049;
  assign n35051 = ~n35046 & ~n35047;
  assign n35052 = ~pi764 & ~n35051;
  assign n35053 = pi764 & ~n35036;
  assign n35054 = ~n35031 & n35053;
  assign n35055 = ~n35052 & ~n35054;
  assign n35056 = pi39 & ~n35055;
  assign n35057 = ~n35038 & n35050;
  assign n35058 = ~n35029 & ~n60395;
  assign n35059 = ~pi38 & ~n35058;
  assign n35060 = ~n32944 & ~n34994;
  assign n35061 = ~pi764 & pi947;
  assign n35062 = ~pi39 & ~n35061;
  assign n35063 = n33372 & n35062;
  assign n35064 = n6863 & ~n35060;
  assign n35065 = ~pi171 & ~n6863;
  assign n35066 = pi38 & ~n35065;
  assign n35067 = pi38 & ~n60396;
  assign n35068 = ~n35065 & n35067;
  assign n35069 = ~n60396 & n35066;
  assign n35070 = pi691 & ~n60397;
  assign n35071 = ~n35059 & n35070;
  assign n35072 = ~n35028 & ~n35071;
  assign n35073 = ~n35059 & ~n60397;
  assign n35074 = pi691 & ~n35073;
  assign n35075 = ~pi691 & ~n34999;
  assign n35076 = ~n35026 & n35075;
  assign n35077 = n25257 & ~n35076;
  assign n35078 = ~n35074 & n35077;
  assign n35079 = n25257 & ~n35072;
  assign n35080 = ~pi171 & ~n25257;
  assign n35081 = ~pi57 & ~n35080;
  assign n35082 = ~n60398 & n35081;
  assign n35083 = pi57 & pi171;
  assign n35084 = ~pi832 & ~n35083;
  assign n35085 = ~n35082 & n35084;
  assign n35086 = pi691 & n32944;
  assign n35087 = ~pi691 & ~n34994;
  assign n35088 = ~n35060 & ~n35087;
  assign n35089 = n2794 & ~n35088;
  assign n35090 = n34995 & ~n35086;
  assign n35091 = pi171 & ~n2794;
  assign n35092 = pi832 & ~n35091;
  assign n35093 = ~n60399 & n35092;
  assign n35094 = ~n35085 & ~n35093;
  assign n35095 = pi690 & n32944;
  assign n35096 = pi739 & pi947;
  assign n35097 = n2794 & ~n35096;
  assign n35098 = ~n35095 & n35097;
  assign n35099 = pi172 & ~n2794;
  assign n35100 = pi832 & ~n35099;
  assign n35101 = ~n35098 & n35100;
  assign n35102 = pi172 & ~n6863;
  assign n35103 = n6863 & ~n35096;
  assign n35104 = n59171 & n35097;
  assign n35105 = pi38 & ~n60400;
  assign n35106 = ~n35102 & n35105;
  assign n35107 = ~pi172 & ~n6627;
  assign n35108 = n33206 & ~n35107;
  assign n35109 = ~pi172 & ~n6464;
  assign n35110 = n33210 & ~n35109;
  assign n35111 = pi172 & ~n6629;
  assign n35112 = pi172 & n6640;
  assign n35113 = ~n6635 & n35111;
  assign n35114 = ~n6634 & ~n60401;
  assign n35115 = ~n35110 & n35114;
  assign n35116 = n33181 & n35115;
  assign n35117 = pi172 & ~n6645;
  assign n35118 = n33071 & ~n35117;
  assign n35119 = ~n33091 & n35118;
  assign n35120 = n33183 & ~n35117;
  assign n35121 = pi299 & ~n60402;
  assign n35122 = ~n35116 & n35121;
  assign n35123 = pi739 & ~n35122;
  assign n35124 = ~n35108 & n35123;
  assign n35125 = ~pi172 & ~pi739;
  assign n35126 = ~n6654 & n35125;
  assign n35127 = pi39 & ~n35126;
  assign n35128 = ~n35124 & n35127;
  assign n35129 = n59147 & n35096;
  assign n35130 = ~pi172 & ~n59147;
  assign n35131 = ~pi39 & ~n35130;
  assign n35132 = ~pi39 & ~n35129;
  assign n35133 = ~n35130 & n35132;
  assign n35134 = ~n35129 & n35131;
  assign n35135 = ~pi38 & ~n60403;
  assign n35136 = ~n35128 & n35135;
  assign n35137 = ~n35106 & ~n35136;
  assign n35138 = ~pi690 & ~n35137;
  assign n35139 = ~n33106 & n60403;
  assign n35140 = pi172 & ~n33151;
  assign n35141 = n33128 & ~n35140;
  assign n35142 = ~n33095 & n35110;
  assign n35143 = ~pi215 & ~n35142;
  assign n35144 = n35114 & n35143;
  assign n35145 = ~n35118 & ~n35144;
  assign n35146 = pi299 & ~n35145;
  assign n35147 = ~n35141 & ~n35146;
  assign n35148 = pi739 & ~n35147;
  assign n35149 = n33097 & ~n35109;
  assign n35150 = ~n33075 & ~n35149;
  assign n35151 = n35114 & n35150;
  assign n35152 = ~pi215 & ~n35151;
  assign n35153 = n33140 & ~n35118;
  assign n35154 = ~n33070 & ~n35153;
  assign n35155 = ~n35152 & n35154;
  assign n35156 = pi299 & ~n35155;
  assign n35157 = n33103 & ~n35107;
  assign n35158 = ~pi739 & ~n35157;
  assign n35159 = ~n35156 & n35158;
  assign n35160 = pi39 & ~n35159;
  assign n35161 = ~n35156 & ~n35157;
  assign n35162 = ~pi739 & ~n35161;
  assign n35163 = pi739 & ~n35146;
  assign n35164 = ~n35141 & n35163;
  assign n35165 = ~n35162 & ~n35164;
  assign n35166 = pi39 & ~n35165;
  assign n35167 = ~n35148 & n35160;
  assign n35168 = ~n35139 & ~n60404;
  assign n35169 = ~pi38 & ~n35168;
  assign n35170 = ~n32944 & ~n35096;
  assign n35171 = ~pi739 & pi947;
  assign n35172 = ~pi39 & ~n35171;
  assign n35173 = n33372 & n35172;
  assign n35174 = n6863 & ~n35170;
  assign n35175 = ~pi172 & ~n6863;
  assign n35176 = pi38 & ~n35175;
  assign n35177 = pi38 & ~n60405;
  assign n35178 = ~n35175 & n35177;
  assign n35179 = ~n60405 & n35176;
  assign n35180 = pi690 & ~n60406;
  assign n35181 = ~n35169 & n35180;
  assign n35182 = ~n35138 & ~n35181;
  assign n35183 = ~n35169 & ~n60406;
  assign n35184 = pi690 & ~n35183;
  assign n35185 = ~pi690 & ~n35106;
  assign n35186 = ~n35136 & n35185;
  assign n35187 = n25257 & ~n35186;
  assign n35188 = ~n35184 & n35187;
  assign n35189 = n25257 & ~n35182;
  assign n35190 = ~pi172 & ~n25257;
  assign n35191 = ~pi57 & ~n35190;
  assign n35192 = ~n60407 & n35191;
  assign n35193 = pi57 & pi172;
  assign n35194 = ~pi832 & ~n35193;
  assign n35195 = ~n35192 & n35194;
  assign n35196 = ~n35101 & ~n35195;
  assign n35197 = ~pi767 & pi947;
  assign n35198 = ~pi698 & n32944;
  assign n35199 = ~n35197 & ~n35198;
  assign n35200 = n2794 & ~n35199;
  assign n35201 = ~pi197 & ~n2794;
  assign n35202 = pi832 & ~n35201;
  assign n35203 = ~n35200 & n35202;
  assign n35204 = ~pi197 & n60293;
  assign n35205 = pi197 & n60297;
  assign n35206 = ~pi767 & ~n35205;
  assign n35207 = ~n35204 & n35206;
  assign n35208 = ~pi197 & n33079;
  assign n35209 = pi197 & n33100;
  assign n35210 = pi299 & ~n35209;
  assign n35211 = ~n35208 & n35210;
  assign n35212 = ~pi197 & ~n6627;
  assign n35213 = n33103 & ~n35212;
  assign n35214 = pi767 & ~n35213;
  assign n35215 = ~n35211 & n35214;
  assign n35216 = pi39 & ~n35215;
  assign n35217 = ~n35207 & n35216;
  assign n35218 = n59147 & n35197;
  assign n35219 = ~pi197 & ~n59147;
  assign n35220 = ~pi39 & ~n35219;
  assign n35221 = ~pi39 & ~n35218;
  assign n35222 = ~n35219 & n35221;
  assign n35223 = ~n35218 & n35220;
  assign n35224 = ~n33106 & n60408;
  assign n35225 = ~pi38 & ~n35224;
  assign n35226 = ~n35217 & n35225;
  assign n35227 = n6863 & ~n35197;
  assign n35228 = ~n32944 & n35227;
  assign n35229 = pi197 & ~n6863;
  assign n35230 = pi38 & ~n35229;
  assign n35231 = ~n35228 & n35230;
  assign n35232 = ~pi698 & ~n35231;
  assign n35233 = ~n35226 & n35232;
  assign n35234 = ~pi197 & ~n33184;
  assign n35235 = pi197 & ~n33266;
  assign n35236 = pi299 & ~n35235;
  assign n35237 = ~n35234 & n35236;
  assign n35238 = n33206 & ~n35212;
  assign n35239 = ~pi767 & ~n35238;
  assign n35240 = ~n35237 & n35239;
  assign n35241 = ~pi197 & pi767;
  assign n35242 = ~n6654 & n35241;
  assign n35243 = pi39 & ~n35242;
  assign n35244 = ~n35240 & n35243;
  assign n35245 = ~pi38 & ~n60408;
  assign n35246 = ~n35244 & n35245;
  assign n35247 = pi38 & ~n35227;
  assign n35248 = ~n35229 & n35247;
  assign n35249 = pi698 & ~n35248;
  assign n35250 = ~n35246 & n35249;
  assign n35251 = n59928 & ~n35250;
  assign n35252 = ~n35246 & ~n35248;
  assign n35253 = pi698 & ~n35252;
  assign n35254 = ~n35217 & ~n35224;
  assign n35255 = ~pi38 & ~n35254;
  assign n35256 = ~n32944 & ~n35197;
  assign n35257 = pi767 & pi947;
  assign n35258 = ~pi39 & ~n35257;
  assign n35259 = n33372 & n35258;
  assign n35260 = n6863 & ~n35256;
  assign n35261 = ~pi197 & ~n6863;
  assign n35262 = pi38 & ~n35261;
  assign n35263 = ~n60409 & n35262;
  assign n35264 = ~pi698 & ~n35263;
  assign n35265 = ~n35255 & n35264;
  assign n35266 = ~n35253 & ~n35265;
  assign n35267 = n59928 & ~n35266;
  assign n35268 = ~n35233 & n35251;
  assign n35269 = ~pi197 & ~n59928;
  assign n35270 = ~pi832 & ~n35269;
  assign n35271 = ~n60410 & n35270;
  assign po354 = ~n35203 & ~n35271;
  assign n35273 = ~pi100 & ~n32919;
  assign n35274 = n28577 & ~n35273;
  assign n35275 = ~pi75 & ~n35274;
  assign n35276 = ~n28303 & ~n35275;
  assign n35277 = ~pi92 & ~n35276;
  assign n35278 = ~pi74 & n4440;
  assign n35279 = n4437 & n31567;
  assign n35280 = n4439 & n31567;
  assign n35281 = ~pi74 & n58992;
  assign n35282 = n4438 & n60411;
  assign n35283 = ~pi54 & ~n28307;
  assign n35284 = n60412 & n35283;
  assign n35285 = ~n28307 & n32859;
  assign po288 = ~n35277 & n60413;
  assign n35287 = n59132 & ~n33837;
  assign n35288 = pi606 & n35287;
  assign n35289 = n59132 & ~n33833;
  assign n35290 = ~pi606 & n35289;
  assign n35291 = pi643 & ~n35290;
  assign n35292 = pi643 & ~n35288;
  assign n35293 = ~n35290 & n35292;
  assign n35294 = ~n35288 & n35291;
  assign n35295 = n59132 & ~n33196;
  assign n35296 = pi606 & n35295;
  assign n35297 = ~pi606 & n7560;
  assign n35298 = n7553 & n24377;
  assign n35299 = ~pi643 & ~n60415;
  assign n35300 = ~n35296 & n35299;
  assign n35301 = n58992 & ~n35300;
  assign n35302 = ~n60414 & n35301;
  assign n35303 = pi211 & ~n35302;
  assign n35304 = n59132 & n33817;
  assign n35305 = pi606 & ~n35304;
  assign n35306 = n59132 & n33814;
  assign n35307 = ~pi606 & ~n35306;
  assign n35308 = pi643 & ~n35307;
  assign n35309 = pi643 & ~n35305;
  assign n35310 = ~n35307 & n35309;
  assign n35311 = ~n35305 & n35308;
  assign n35312 = n59132 & n33218;
  assign n35313 = pi606 & ~pi643;
  assign n35314 = n35312 & n35313;
  assign n35315 = ~n60416 & ~n35314;
  assign n35316 = ~pi211 & n58992;
  assign n35317 = ~n35315 & n35316;
  assign n35318 = ~n35303 & ~n35317;
  assign n35319 = pi607 & n35287;
  assign n35320 = ~pi607 & n35289;
  assign n35321 = pi638 & ~n35320;
  assign n35322 = pi638 & ~n35319;
  assign n35323 = ~n35320 & n35322;
  assign n35324 = ~n35319 & n35321;
  assign n35325 = pi607 & n35295;
  assign n35326 = ~pi607 & n7560;
  assign n35327 = ~pi638 & ~n35326;
  assign n35328 = ~n35325 & n35327;
  assign n35329 = n58992 & ~n35328;
  assign n35330 = ~n60417 & n35329;
  assign n35331 = ~pi212 & ~n35330;
  assign n35332 = pi607 & ~n35304;
  assign n35333 = ~pi607 & ~n35306;
  assign n35334 = pi638 & ~n35333;
  assign n35335 = pi638 & ~n35332;
  assign n35336 = ~n35333 & n35335;
  assign n35337 = ~n35332 & n35334;
  assign n35338 = pi607 & ~pi638;
  assign n35339 = n35312 & n35338;
  assign n35340 = ~n60418 & ~n35339;
  assign n35341 = pi212 & n58992;
  assign n35342 = ~n35340 & n35341;
  assign n35343 = ~n35331 & ~n35342;
  assign n35344 = pi213 & n58992;
  assign n35345 = pi622 & ~n35304;
  assign n35346 = ~pi622 & ~n35306;
  assign n35347 = pi639 & ~n35346;
  assign n35348 = pi639 & ~n35345;
  assign n35349 = ~n35346 & n35348;
  assign n35350 = ~n35345 & n35347;
  assign n35351 = pi622 & ~pi639;
  assign n35352 = n35312 & n35351;
  assign n35353 = ~n60419 & ~n35352;
  assign n35354 = n35344 & ~n35353;
  assign n35355 = ~pi639 & n35295;
  assign n35356 = pi639 & n35287;
  assign n35357 = pi622 & ~n35356;
  assign n35358 = pi622 & ~n35355;
  assign n35359 = ~n35356 & n35358;
  assign n35360 = ~n35355 & n35357;
  assign n35361 = pi639 & n35289;
  assign n35362 = ~pi639 & n7560;
  assign n35363 = ~pi622 & ~n35362;
  assign n35364 = ~n35361 & n35363;
  assign n35365 = n58992 & ~n35364;
  assign n35366 = pi639 & ~n35287;
  assign n35367 = ~pi639 & ~n35295;
  assign n35368 = pi622 & ~n35367;
  assign n35369 = ~n35366 & n35368;
  assign n35370 = pi639 & ~n35289;
  assign n35371 = ~pi639 & ~n7560;
  assign n35372 = ~pi622 & ~n35371;
  assign n35373 = ~n35370 & n35372;
  assign n35374 = ~n35369 & ~n35373;
  assign n35375 = n58992 & ~n35374;
  assign n35376 = ~n60420 & n35365;
  assign n35377 = ~pi213 & ~n60421;
  assign n35378 = ~n35354 & ~n35377;
  assign n35379 = pi623 & n35287;
  assign n35380 = ~pi623 & n35289;
  assign n35381 = pi710 & ~n35380;
  assign n35382 = pi710 & ~n35379;
  assign n35383 = ~n35380 & n35382;
  assign n35384 = ~n35379 & n35381;
  assign n35385 = pi623 & n35295;
  assign n35386 = ~pi623 & n7560;
  assign n35387 = ~pi710 & ~n35386;
  assign n35388 = ~n35385 & n35387;
  assign n35389 = n58992 & ~n35388;
  assign n35390 = ~n60422 & n35389;
  assign n35391 = ~pi214 & ~n35390;
  assign n35392 = pi623 & ~n35304;
  assign n35393 = ~pi623 & ~n35306;
  assign n35394 = pi710 & ~n35393;
  assign n35395 = pi710 & ~n35392;
  assign n35396 = ~n35393 & n35395;
  assign n35397 = ~n35392 & n35394;
  assign n35398 = pi623 & ~pi710;
  assign n35399 = n35312 & n35398;
  assign n35400 = ~n60423 & ~n35399;
  assign n35401 = pi214 & n58992;
  assign n35402 = ~n35400 & n35401;
  assign n35403 = ~n35391 & ~n35402;
  assign n35404 = ~pi219 & n58992;
  assign n35405 = pi617 & ~n35304;
  assign n35406 = ~pi617 & ~n35306;
  assign n35407 = pi637 & ~n35406;
  assign n35408 = pi637 & ~n35405;
  assign n35409 = ~n35406 & n35408;
  assign n35410 = ~n35405 & n35407;
  assign n35411 = pi617 & ~pi637;
  assign n35412 = n35312 & n35411;
  assign n35413 = ~n60424 & ~n35412;
  assign n35414 = n35404 & ~n35413;
  assign n35415 = ~pi617 & n35289;
  assign n35416 = pi617 & n35287;
  assign n35417 = pi637 & ~n35416;
  assign n35418 = pi637 & ~n35415;
  assign n35419 = ~n35416 & n35418;
  assign n35420 = ~n35415 & n35417;
  assign n35421 = pi617 & n35295;
  assign n35422 = ~pi617 & n7560;
  assign n35423 = ~pi637 & ~n35422;
  assign n35424 = ~n35421 & n35423;
  assign n35425 = n58992 & ~n35424;
  assign n35426 = pi617 & ~n35287;
  assign n35427 = ~pi617 & ~n35289;
  assign n35428 = pi637 & ~n35427;
  assign n35429 = ~n35426 & n35428;
  assign n35430 = pi617 & ~n35295;
  assign n35431 = ~pi617 & ~n7560;
  assign n35432 = ~pi637 & ~n35431;
  assign n35433 = ~n35430 & n35432;
  assign n35434 = ~n35429 & ~n35433;
  assign n35435 = n58992 & ~n35434;
  assign n35436 = ~n60425 & n35425;
  assign n35437 = pi219 & ~n60426;
  assign n35438 = ~n35414 & ~n35437;
  assign n35439 = pi634 & n32944;
  assign n35440 = pi633 & pi947;
  assign n35441 = ~n35439 & ~n35440;
  assign n35442 = n6863 & ~n35441;
  assign n35443 = pi210 & ~n6863;
  assign n35444 = pi38 & ~n35443;
  assign n35445 = pi38 & ~n35442;
  assign n35446 = ~n35443 & n35445;
  assign n35447 = ~n35442 & n35444;
  assign n35448 = pi210 & ~n6464;
  assign n35449 = n2782 & n35448;
  assign n35450 = pi210 & ~n2782;
  assign n35451 = ~n6587 & n35450;
  assign n35452 = ~n35449 & ~n35451;
  assign n35453 = ~pi907 & n35452;
  assign n35454 = ~n25722 & ~n35448;
  assign n35455 = ~n2783 & ~n35454;
  assign n35456 = pi907 & ~n35455;
  assign n35457 = pi210 & n6566;
  assign n35458 = pi634 & ~n6566;
  assign n35459 = ~n35457 & ~n35458;
  assign n35460 = n2783 & ~n35459;
  assign n35461 = n35456 & ~n35460;
  assign n35462 = ~pi947 & ~n35461;
  assign n35463 = ~n35453 & n35462;
  assign n35464 = ~n25489 & ~n35448;
  assign n35465 = n2782 & n35464;
  assign n35466 = pi947 & ~n35465;
  assign n35467 = ~n2782 & n35464;
  assign n35468 = ~n2783 & ~n35467;
  assign n35469 = pi633 & ~n6566;
  assign n35470 = ~n35457 & ~n35469;
  assign n35471 = ~n2680 & ~n35470;
  assign n35472 = ~n35468 & ~n35471;
  assign n35473 = n35466 & ~n35472;
  assign n35474 = n2790 & ~n35473;
  assign n35475 = ~n35463 & n35474;
  assign n35476 = n2822 & n35454;
  assign n35477 = pi907 & ~n35476;
  assign n35478 = ~n2822 & n35459;
  assign n35479 = n35477 & ~n35478;
  assign n35480 = pi210 & ~n59152;
  assign n35481 = ~pi907 & n35480;
  assign n35482 = ~n35479 & ~n35481;
  assign n35483 = ~pi947 & ~n35482;
  assign n35484 = n2822 & n35464;
  assign n35485 = pi947 & ~n35484;
  assign n35486 = ~n2822 & n35470;
  assign n35487 = n35485 & ~n35486;
  assign n35488 = ~n2790 & ~n35487;
  assign n35489 = ~n35483 & n35488;
  assign n35490 = ~n35475 & ~n35489;
  assign n35491 = ~n6544 & ~n35490;
  assign n35492 = n6464 & ~n35441;
  assign n35493 = ~n35448 & ~n35492;
  assign n35494 = n6544 & n35493;
  assign n35495 = ~pi223 & ~n35494;
  assign n35496 = ~n35491 & n35495;
  assign n35497 = ~n6490 & n35450;
  assign n35498 = ~n35449 & ~n35497;
  assign n35499 = ~pi907 & n35498;
  assign n35500 = pi210 & n6484;
  assign n35501 = ~n25663 & ~n35500;
  assign n35502 = n2783 & ~n35501;
  assign n35503 = n35456 & ~n35502;
  assign n35504 = ~pi947 & ~n35503;
  assign n35505 = ~n35499 & n35504;
  assign n35506 = pi633 & ~n6484;
  assign n35507 = ~n35500 & ~n35506;
  assign n35508 = ~n2680 & ~n35507;
  assign n35509 = ~n35468 & ~n35508;
  assign n35510 = n35466 & ~n35509;
  assign n35511 = n2790 & ~n35510;
  assign n35512 = ~n35505 & n35511;
  assign n35513 = ~n2822 & n35501;
  assign n35514 = n35477 & ~n35513;
  assign n35515 = n2822 & n6463;
  assign n35516 = n2794 & n35515;
  assign n35517 = n35500 & ~n35516;
  assign n35518 = ~n35514 & ~n35517;
  assign n35519 = ~pi947 & ~n35518;
  assign n35520 = ~n2822 & n35507;
  assign n35521 = n35485 & ~n35520;
  assign n35522 = ~n2790 & ~n35521;
  assign n35523 = ~n35519 & n35522;
  assign n35524 = pi223 & ~n35523;
  assign n35525 = pi223 & ~n35512;
  assign n35526 = ~n35523 & n35525;
  assign n35527 = ~n35512 & n35524;
  assign n35528 = ~pi299 & ~n60428;
  assign n35529 = ~n35496 & n35528;
  assign n35530 = ~n2839 & ~n35480;
  assign n35531 = n2839 & n35452;
  assign n35532 = ~pi907 & ~n35531;
  assign n35533 = ~n35530 & n35532;
  assign n35534 = ~n35479 & ~n35533;
  assign n35535 = ~pi947 & ~n35534;
  assign n35536 = ~n6629 & ~n35487;
  assign n35537 = ~n35535 & n35536;
  assign n35538 = n6629 & n35493;
  assign n35539 = ~pi215 & ~n35538;
  assign n35540 = ~n35537 & n35539;
  assign n35541 = n2839 & n35498;
  assign n35542 = ~n2839 & ~n35517;
  assign n35543 = ~pi907 & ~n35542;
  assign n35544 = ~n35541 & n35543;
  assign n35545 = ~n35514 & ~n35544;
  assign n35546 = ~pi947 & ~n35545;
  assign n35547 = ~n35521 & ~n35546;
  assign n35548 = pi215 & ~n35547;
  assign n35549 = pi299 & ~n35548;
  assign n35550 = ~n35540 & n35549;
  assign n35551 = pi39 & ~n35550;
  assign n35552 = ~n35529 & n35551;
  assign n35553 = n6449 & ~n35441;
  assign n35554 = pi210 & ~n6449;
  assign n35555 = ~pi299 & ~n35554;
  assign n35556 = ~pi299 & ~n35553;
  assign n35557 = ~n35554 & n35556;
  assign n35558 = ~n35553 & n35555;
  assign n35559 = ~n6451 & ~n35441;
  assign n35560 = pi299 & ~n35559;
  assign n35561 = pi299 & ~n6452;
  assign n35562 = ~n35559 & n35561;
  assign n35563 = ~n6452 & n35560;
  assign n35564 = ~pi39 & ~n60430;
  assign n35565 = ~n60429 & n35564;
  assign n35566 = ~pi38 & ~n35565;
  assign n35567 = ~n35552 & n35566;
  assign n35568 = ~n60427 & ~n35567;
  assign n35569 = n59928 & ~n35568;
  assign n35570 = ~pi210 & ~n59928;
  assign po367 = ~n35569 & ~n35570;
  assign n35572 = ~pi51 & pi70;
  assign n35573 = n2593 & n35572;
  assign n35574 = ~pi96 & n35573;
  assign n35575 = pi24 & n60280;
  assign n35576 = pi24 & n32908;
  assign n35577 = n2618 & n35573;
  assign n35578 = n2597 & n35574;
  assign n35579 = n35576 & n60431;
  assign n35580 = n35574 & n35575;
  assign n35581 = pi198 & pi589;
  assign n35582 = n2828 & n6544;
  assign n35583 = ~pi223 & n6544;
  assign n35584 = n28532 & n35583;
  assign n35585 = ~n2792 & n35582;
  assign n35586 = n35581 & n60433;
  assign n35587 = pi210 & pi589;
  assign n35588 = ~pi221 & n2851;
  assign n35589 = ~pi216 & n60434;
  assign n35590 = n2851 & n6629;
  assign n35591 = ~pi215 & n6629;
  assign n35592 = n28524 & n35591;
  assign n35593 = ~n2845 & n60435;
  assign n35594 = n35587 & n60436;
  assign n35595 = ~n35586 & ~n35594;
  assign n35596 = ~pi593 & n2806;
  assign n35597 = ~n28514 & n35596;
  assign n35598 = ~n35595 & n35597;
  assign n35599 = ~pi287 & ~n35598;
  assign n35600 = pi39 & ~n35599;
  assign n35601 = n58822 & n35600;
  assign n35602 = ~n60432 & ~n35601;
  assign po228 = n32632 & ~n35602;
  assign n35604 = ~n35587 & n60436;
  assign n35605 = ~n2792 & n2828;
  assign n35606 = n6544 & ~n35581;
  assign n35607 = n35605 & n35606;
  assign n35608 = ~n35604 & ~n35607;
  assign n35609 = ~n28517 & ~n35608;
  assign n35610 = ~n35581 & n35582;
  assign n35611 = n30786 & n35610;
  assign n35612 = ~n28517 & n35604;
  assign n35613 = pi39 & ~n35612;
  assign n35614 = ~n35611 & n35613;
  assign n35615 = pi39 & ~n35609;
  assign n35616 = pi24 & n28317;
  assign n35617 = n2597 & n30356;
  assign n35618 = n35616 & n35617;
  assign n35619 = ~pi71 & n2446;
  assign n35620 = ~pi104 & n2450;
  assign n35621 = n35619 & n35620;
  assign n35622 = ~pi49 & ~pi66;
  assign n35623 = ~pi45 & ~pi73;
  assign n35624 = n35622 & n35623;
  assign n35625 = ~pi48 & ~pi65;
  assign n35626 = pi89 & n35625;
  assign n35627 = n35624 & n35626;
  assign n35628 = pi89 & n29132;
  assign n35629 = n35625 & n35628;
  assign n35630 = n35624 & n35629;
  assign n35631 = n29141 & n35630;
  assign n35632 = n60119 & n35627;
  assign n35633 = n35621 & n60438;
  assign n35634 = n2547 & n35633;
  assign n35635 = ~pi841 & n2579;
  assign n35636 = ~pi332 & n60165;
  assign n35637 = n35635 & n35636;
  assign n35638 = n35634 & n35637;
  assign n35639 = ~pi39 & ~n35638;
  assign n35640 = ~n35618 & n35639;
  assign n35641 = n32632 & ~n35640;
  assign po253 = ~n60437 & n35641;
  assign n35643 = pi39 & pi593;
  assign n35644 = ~n35595 & n35643;
  assign n35645 = ~n28517 & n35644;
  assign n35646 = n58835 & n31405;
  assign n35647 = pi829 & ~pi1093;
  assign n35648 = n2441 & n35647;
  assign n35649 = ~n58838 & ~n35648;
  assign n35650 = pi479 & n35649;
  assign n35651 = n60122 & n35650;
  assign n35652 = ~po740 & ~n35651;
  assign n35653 = n60279 & ~n35652;
  assign n35654 = n35646 & n35653;
  assign n35655 = ~n35645 & ~n35654;
  assign po255 = n32632 & ~n35655;
  assign n35657 = pi215 & ~n59928;
  assign n35658 = pi681 & pi907;
  assign n35659 = n33566 & ~n35658;
  assign n35660 = n6589 & n6700;
  assign n35661 = ~pi642 & n26927;
  assign n35662 = ~n2781 & ~n35661;
  assign n35663 = ~n35660 & n35662;
  assign n35664 = n2781 & ~n26936;
  assign n35665 = n2790 & ~n35664;
  assign n35666 = ~n35663 & n35665;
  assign n35667 = ~pi642 & n59152;
  assign n35668 = ~n2790 & n35667;
  assign n35669 = ~n35666 & ~n35668;
  assign n35670 = ~n35660 & ~n35661;
  assign n35671 = ~n2781 & ~n35670;
  assign n35672 = n2781 & n26936;
  assign n35673 = n2790 & ~n35672;
  assign n35674 = ~n35663 & ~n35664;
  assign n35675 = n2790 & ~n35674;
  assign n35676 = ~n35671 & n35673;
  assign n35677 = ~n2790 & ~n35667;
  assign n35678 = pi947 & ~n35677;
  assign n35679 = ~n60439 & n35678;
  assign n35680 = pi947 & ~n35669;
  assign n35681 = ~n6544 & ~n60440;
  assign n35682 = ~n35659 & n35681;
  assign n35683 = ~n6464 & n6544;
  assign n35684 = ~pi947 & n35658;
  assign n35685 = pi642 & pi947;
  assign n35686 = ~n35684 & ~n35685;
  assign n35687 = n6544 & ~n35686;
  assign n35688 = ~pi223 & ~n35687;
  assign n35689 = ~n35683 & n35688;
  assign n35690 = ~n35682 & n35689;
  assign n35691 = ~n2781 & ~n6502;
  assign n35692 = n6518 & n6522;
  assign n35693 = n2781 & ~n6490;
  assign n35694 = ~pi642 & ~n60441;
  assign n35695 = ~pi642 & n59149;
  assign n35696 = ~n35691 & n35694;
  assign n35697 = n2790 & ~n60442;
  assign n35698 = ~n2781 & ~n6496;
  assign n35699 = ~pi642 & ~n26237;
  assign n35700 = ~n35698 & n35699;
  assign n35701 = ~n2790 & ~n35700;
  assign n35702 = pi947 & ~n35701;
  assign n35703 = ~n35697 & n35702;
  assign n35704 = ~n33122 & ~n35703;
  assign n35705 = pi223 & ~n35684;
  assign n35706 = ~n35704 & n35705;
  assign n35707 = ~pi299 & ~n35706;
  assign n35708 = ~n35690 & n35707;
  assign n35709 = ~pi947 & n33475;
  assign n35710 = pi947 & ~n35700;
  assign n35711 = ~n35684 & ~n35710;
  assign n35712 = ~n35709 & n35711;
  assign n35713 = pi299 & ~n35712;
  assign n35714 = ~n35708 & ~n35713;
  assign n35715 = pi215 & ~n35714;
  assign n35716 = n6595 & n35684;
  assign n35717 = pi642 & ~n6518;
  assign n35718 = n6464 & n35717;
  assign n35719 = pi642 & n6518;
  assign n35720 = ~n6527 & n35719;
  assign n35721 = ~n6606 & n35720;
  assign n35722 = ~n35718 & ~n35721;
  assign n35723 = pi947 & ~n35722;
  assign n35724 = n2790 & ~n35723;
  assign n35725 = ~n35716 & n35724;
  assign n35726 = ~n59151 & n35658;
  assign n35727 = ~pi947 & ~n35726;
  assign n35728 = ~n2781 & n6568;
  assign n35729 = ~n6576 & ~n35728;
  assign n35730 = n35719 & n35729;
  assign n35731 = ~n6568 & n35717;
  assign n35732 = pi947 & ~n35731;
  assign n35733 = ~n35730 & n35732;
  assign n35734 = ~n35727 & ~n35733;
  assign n35735 = ~n2790 & ~n35734;
  assign n35736 = ~n6544 & ~n35735;
  assign n35737 = ~n35725 & n35736;
  assign n35738 = n59155 & ~n35686;
  assign n35739 = n6464 & n35687;
  assign n35740 = ~pi223 & ~n60443;
  assign n35741 = ~n35737 & n35740;
  assign n35742 = n2790 & ~n6502;
  assign n35743 = n35658 & ~n35742;
  assign n35744 = ~pi947 & ~n35743;
  assign n35745 = pi947 & ~n6486;
  assign n35746 = ~n6496 & ~n35745;
  assign n35747 = ~n2790 & n35746;
  assign n35748 = ~n6522 & n35720;
  assign n35749 = pi947 & ~n35718;
  assign n35750 = ~n35748 & n35749;
  assign n35751 = ~n35747 & ~n35750;
  assign n35752 = ~n35744 & n35751;
  assign n35753 = pi223 & ~n35752;
  assign n35754 = ~n35741 & ~n35753;
  assign n35755 = ~pi299 & ~n35754;
  assign n35756 = ~n6629 & n35734;
  assign n35757 = n6637 & ~n35686;
  assign n35758 = pi299 & ~n35757;
  assign n35759 = ~n35756 & n35758;
  assign n35760 = ~pi215 & ~n35759;
  assign n35761 = ~n35755 & n35760;
  assign n35762 = ~n35715 & ~n35761;
  assign n35763 = pi39 & ~n35762;
  assign n35764 = n6453 & n35686;
  assign n35765 = ~pi215 & ~n6453;
  assign n35766 = pi299 & ~n35765;
  assign n35767 = ~n35764 & n35766;
  assign n35768 = n6449 & n35686;
  assign n35769 = ~pi215 & ~n6449;
  assign n35770 = ~pi299 & ~n35769;
  assign n35771 = ~n35768 & n35770;
  assign n35772 = ~n35767 & ~n35771;
  assign n35773 = pi215 & ~n6449;
  assign n35774 = n6449 & ~n35686;
  assign n35775 = ~pi299 & ~n35774;
  assign n35776 = ~n35773 & n35775;
  assign n35777 = pi215 & ~n6453;
  assign n35778 = n6453 & ~n35686;
  assign n35779 = pi299 & ~n35778;
  assign n35780 = pi299 & ~n35777;
  assign n35781 = ~n35778 & n35780;
  assign n35782 = ~n35777 & n35779;
  assign n35783 = ~pi39 & ~n60444;
  assign n35784 = ~n35776 & n35783;
  assign n35785 = ~pi39 & ~n35776;
  assign n35786 = ~n60444 & n35785;
  assign n35787 = ~pi39 & ~n35772;
  assign n35788 = ~pi38 & ~n60445;
  assign n35789 = ~n35763 & n35788;
  assign n35790 = n6863 & ~n35686;
  assign n35791 = pi215 & ~n6863;
  assign n35792 = pi38 & ~n35791;
  assign n35793 = pi38 & ~n35790;
  assign n35794 = ~n35791 & n35793;
  assign n35795 = ~n35790 & n35792;
  assign n35796 = n59928 & ~n60446;
  assign n35797 = ~n35789 & n35796;
  assign n35798 = ~n35657 & ~n35797;
  assign n35799 = pi216 & ~n6863;
  assign n35800 = pi662 & pi907;
  assign n35801 = ~pi947 & n35800;
  assign n35802 = pi614 & pi947;
  assign n35803 = ~n35801 & ~n35802;
  assign n35804 = n6863 & ~n35803;
  assign n35805 = pi38 & ~n35804;
  assign n35806 = pi38 & ~n35799;
  assign n35807 = ~n35804 & n35806;
  assign n35808 = ~n35799 & n35805;
  assign n35809 = ~n6522 & n6608;
  assign n35810 = pi947 & ~n6611;
  assign n35811 = ~n35809 & n35810;
  assign n35812 = ~n35745 & ~n35801;
  assign n35813 = ~n35811 & ~n35812;
  assign n35814 = n6496 & n35800;
  assign n35815 = ~pi947 & ~n35814;
  assign n35816 = pi947 & n6486;
  assign n35817 = ~n35811 & ~n35816;
  assign n35818 = ~n35815 & n35817;
  assign n35819 = ~n35746 & n35813;
  assign n35820 = ~pi216 & ~n60448;
  assign n35821 = n6598 & ~n27677;
  assign n35822 = n2781 & n27681;
  assign n35823 = ~n35821 & ~n35822;
  assign n35824 = pi947 & n35823;
  assign n35825 = pi216 & ~n35801;
  assign n35826 = ~n35824 & n35825;
  assign n35827 = ~n35709 & n35826;
  assign n35828 = ~n35820 & ~n35827;
  assign n35829 = pi215 & ~n35828;
  assign n35830 = pi947 & ~n59152;
  assign n35831 = ~pi614 & n59152;
  assign n35832 = pi947 & ~n35831;
  assign n35833 = ~n35801 & ~n35832;
  assign n35834 = n35803 & ~n35830;
  assign n35835 = ~pi947 & n33179;
  assign n35836 = n60449 & ~n35835;
  assign n35837 = ~n59293 & n35803;
  assign n35838 = pi216 & ~n60450;
  assign n35839 = n35729 & n35802;
  assign n35840 = ~n59151 & n35801;
  assign n35841 = ~n35839 & ~n35840;
  assign n35842 = n2850 & ~n35841;
  assign n35843 = n6637 & ~n35803;
  assign n35844 = ~pi215 & ~n35843;
  assign n35845 = ~n35842 & n35844;
  assign n35846 = ~n35838 & n35845;
  assign n35847 = ~n35829 & ~n35846;
  assign n35848 = ~n35842 & ~n35843;
  assign n35849 = ~n35838 & n35848;
  assign n35850 = ~pi215 & ~n35849;
  assign n35851 = pi215 & ~n35820;
  assign n35852 = ~n35827 & n35851;
  assign n35853 = pi299 & ~n35852;
  assign n35854 = ~n35850 & n35853;
  assign n35855 = pi299 & ~n35847;
  assign n35856 = pi947 & ~n6605;
  assign n35857 = ~pi947 & ~n35800;
  assign n35858 = ~pi947 & n6615;
  assign n35859 = ~n35800 & n35858;
  assign n35860 = n6615 & n35857;
  assign n35861 = ~n35856 & ~n60452;
  assign n35862 = n2790 & ~n35861;
  assign n35863 = ~pi947 & ~n59152;
  assign n35864 = ~n2790 & ~n35801;
  assign n35865 = ~n35832 & n35864;
  assign n35866 = ~n35863 & n35865;
  assign n35867 = ~n2790 & ~n35863;
  assign n35868 = n60449 & n35867;
  assign n35869 = n6584 & n35803;
  assign n35870 = ~n6544 & ~n60453;
  assign n35871 = ~n35862 & n35870;
  assign n35872 = n6544 & ~n35803;
  assign n35873 = ~pi223 & ~n35872;
  assign n35874 = ~n35683 & n35873;
  assign n35875 = ~n35871 & n35874;
  assign n35876 = ~pi616 & n6492;
  assign n35877 = ~n2781 & ~n6531;
  assign n35878 = ~n35876 & n35877;
  assign n35879 = ~pi614 & ~n60441;
  assign n35880 = ~pi616 & ~n6492;
  assign n35881 = ~n2781 & ~n6498;
  assign n35882 = ~n35880 & n35881;
  assign n35883 = ~n6514 & ~n35882;
  assign n35884 = ~pi614 & ~n35883;
  assign n35885 = ~n35878 & n35879;
  assign n35886 = n2790 & ~n60454;
  assign n35887 = ~n2790 & n35823;
  assign n35888 = pi947 & ~n35887;
  assign n35889 = ~n35886 & n35888;
  assign n35890 = ~n33122 & ~n35889;
  assign n35891 = pi223 & ~n35801;
  assign n35892 = ~n35890 & n35891;
  assign n35893 = pi216 & ~n35892;
  assign n35894 = ~n35875 & n35893;
  assign n35895 = n6595 & n35801;
  assign n35896 = pi947 & ~n6612;
  assign n35897 = n2790 & ~n35896;
  assign n35898 = ~n35895 & n35897;
  assign n35899 = ~n2790 & n35841;
  assign n35900 = ~n6544 & ~n35899;
  assign n35901 = ~n35898 & n35900;
  assign n35902 = n59155 & ~n35803;
  assign n35903 = n6464 & n35872;
  assign n35904 = ~pi223 & ~n60455;
  assign n35905 = ~n35901 & n35904;
  assign n35906 = ~n35742 & n35800;
  assign n35907 = ~pi947 & ~n35906;
  assign n35908 = ~n35747 & ~n35811;
  assign n35909 = ~n35907 & n35908;
  assign n35910 = pi223 & ~n35909;
  assign n35911 = ~pi216 & ~n35910;
  assign n35912 = ~n35905 & n35911;
  assign n35913 = ~pi299 & ~n35912;
  assign n35914 = ~n35894 & n35913;
  assign n35915 = pi39 & ~n35914;
  assign n35916 = ~n60451 & n35915;
  assign n35917 = n6453 & n35803;
  assign n35918 = ~pi216 & ~n6453;
  assign n35919 = pi299 & ~n35918;
  assign n35920 = ~n35917 & n35919;
  assign n35921 = n6449 & n35803;
  assign n35922 = ~pi216 & ~n6449;
  assign n35923 = ~pi299 & ~n35922;
  assign n35924 = ~n35921 & n35923;
  assign n35925 = ~n35920 & ~n35924;
  assign n35926 = pi216 & ~n6449;
  assign n35927 = n6449 & ~n35803;
  assign n35928 = ~pi299 & ~n35927;
  assign n35929 = ~n35926 & n35928;
  assign n35930 = pi216 & ~n6453;
  assign n35931 = n6453 & ~n35803;
  assign n35932 = pi299 & ~n35931;
  assign n35933 = pi299 & ~n35930;
  assign n35934 = ~n35931 & n35933;
  assign n35935 = ~n35930 & n35932;
  assign n35936 = ~pi39 & ~n60456;
  assign n35937 = ~n35929 & n35936;
  assign n35938 = ~pi39 & ~n35929;
  assign n35939 = ~n60456 & n35938;
  assign n35940 = ~pi39 & ~n35925;
  assign n35941 = ~pi38 & ~n60457;
  assign n35942 = ~n35916 & n35941;
  assign n35943 = ~n60447 & ~n35942;
  assign n35944 = n59928 & ~n35943;
  assign n35945 = ~pi216 & ~n59928;
  assign po373 = ~n35944 & ~n35945;
  assign n35947 = n6605 & ~n6609;
  assign n35948 = n6523 & ~n35947;
  assign n35949 = n6519 & n6593;
  assign n35950 = ~n35948 & ~n35949;
  assign n35951 = pi947 & ~n35950;
  assign n35952 = n2790 & ~n35858;
  assign n35953 = ~n35951 & n35952;
  assign n35954 = pi661 & pi907;
  assign n35955 = ~pi947 & n35954;
  assign n35956 = ~n6518 & n26182;
  assign n35957 = n6519 & ~n26181;
  assign n35958 = ~n35667 & ~n35730;
  assign n35959 = n6523 & ~n35958;
  assign n35960 = pi947 & ~n35959;
  assign n35961 = ~n60458 & ~n35959;
  assign n35962 = pi947 & n35961;
  assign n35963 = ~n60458 & n35960;
  assign n35964 = ~n35863 & ~n60459;
  assign n35965 = ~n2790 & ~n35964;
  assign n35966 = ~n35955 & ~n35965;
  assign n35967 = n2790 & ~n35949;
  assign n35968 = ~n35948 & n35967;
  assign n35969 = ~n2790 & n35961;
  assign n35970 = ~n35968 & ~n35969;
  assign n35971 = pi947 & ~n35970;
  assign n35972 = ~pi947 & ~n59154;
  assign n35973 = ~n35955 & ~n35972;
  assign n35974 = ~n35971 & n35973;
  assign n35975 = ~n35953 & n35966;
  assign n35976 = ~n6544 & ~n60460;
  assign n35977 = pi616 & pi947;
  assign n35978 = ~n35955 & ~n35977;
  assign n35979 = n6464 & ~n35978;
  assign n35980 = n6544 & n35979;
  assign n35981 = n59155 & ~n35978;
  assign n35982 = ~pi223 & ~n60461;
  assign n35983 = ~n35683 & n35982;
  assign n35984 = ~n35976 & n35983;
  assign n35985 = ~pi947 & ~n6512;
  assign n35986 = ~n6486 & ~n6493;
  assign n35987 = ~n2781 & ~n35986;
  assign n35988 = ~pi616 & ~n26237;
  assign n35989 = ~n35987 & n35988;
  assign n35990 = pi947 & ~n35989;
  assign n35991 = ~n35985 & ~n35990;
  assign n35992 = ~n2790 & ~n35991;
  assign n35993 = ~pi947 & n59149;
  assign n35994 = pi947 & ~n6526;
  assign n35995 = n2790 & ~n35994;
  assign n35996 = ~n35993 & n35995;
  assign n35997 = pi223 & ~n35955;
  assign n35998 = ~n35996 & n35997;
  assign n35999 = ~n35992 & n35998;
  assign n36000 = pi221 & ~n35999;
  assign n36001 = ~n35984 & n36000;
  assign n36002 = n6595 & n35955;
  assign n36003 = n6529 & ~n6606;
  assign n36004 = ~n6532 & ~n36003;
  assign n36005 = pi947 & ~n36004;
  assign n36006 = n2790 & ~n36005;
  assign n36007 = ~n36002 & n36006;
  assign n36008 = n35729 & n35977;
  assign n36009 = ~n59151 & n35955;
  assign n36010 = ~n36008 & ~n36009;
  assign n36011 = ~n2790 & n36010;
  assign n36012 = ~n6544 & ~n36011;
  assign n36013 = ~n36007 & n36012;
  assign n36014 = n35982 & ~n36013;
  assign n36015 = pi947 & ~n6533;
  assign n36016 = ~n35955 & ~n36015;
  assign n36017 = ~n35747 & ~n36016;
  assign n36018 = ~n35742 & n36017;
  assign n36019 = pi223 & ~n36018;
  assign n36020 = ~pi221 & ~n36019;
  assign n36021 = ~n36014 & n36020;
  assign n36022 = ~pi299 & ~n36021;
  assign n36023 = ~n36001 & n36022;
  assign n36024 = ~n33179 & ~n35954;
  assign n36025 = ~pi947 & ~n36024;
  assign n36026 = pi221 & ~n60459;
  assign n36027 = ~n36025 & n36026;
  assign n36028 = pi216 & ~n36010;
  assign n36029 = ~pi216 & ~n35978;
  assign n36030 = ~pi216 & n35979;
  assign n36031 = n6464 & n36029;
  assign n36032 = ~pi221 & ~n60462;
  assign n36033 = ~n36028 & n36032;
  assign n36034 = ~pi215 & ~n36033;
  assign n36035 = ~n36027 & n36034;
  assign n36036 = pi221 & ~n35955;
  assign n36037 = ~n35990 & n36036;
  assign n36038 = ~n35709 & n36037;
  assign n36039 = ~n35746 & ~n36016;
  assign n36040 = ~pi221 & ~n36039;
  assign n36041 = pi215 & ~n36040;
  assign n36042 = ~n36038 & n36041;
  assign n36043 = pi299 & ~n36042;
  assign n36044 = ~n36035 & n36043;
  assign n36045 = pi39 & ~n36044;
  assign n36046 = pi39 & ~n36023;
  assign n36047 = ~n36044 & n36046;
  assign n36048 = ~n36023 & n36045;
  assign n36049 = n6453 & n35978;
  assign n36050 = ~pi221 & ~n6453;
  assign n36051 = pi299 & ~n36050;
  assign n36052 = ~n36049 & n36051;
  assign n36053 = n6449 & n35978;
  assign n36054 = ~pi221 & ~n6449;
  assign n36055 = ~pi299 & ~n36054;
  assign n36056 = ~n36053 & n36055;
  assign n36057 = ~n36052 & ~n36056;
  assign n36058 = pi221 & ~n6449;
  assign n36059 = n6449 & ~n35978;
  assign n36060 = ~pi299 & ~n36059;
  assign n36061 = ~n36058 & n36060;
  assign n36062 = pi221 & ~n6453;
  assign n36063 = n6453 & ~n35978;
  assign n36064 = pi299 & ~n36063;
  assign n36065 = pi299 & ~n36062;
  assign n36066 = ~n36063 & n36065;
  assign n36067 = ~n36062 & n36064;
  assign n36068 = ~pi39 & ~n60464;
  assign n36069 = ~n36061 & n36068;
  assign n36070 = ~pi39 & ~n36061;
  assign n36071 = ~n60464 & n36070;
  assign n36072 = ~pi39 & ~n36057;
  assign n36073 = ~pi38 & ~n60465;
  assign n36074 = ~n60463 & n36073;
  assign n36075 = pi221 & ~n6863;
  assign n36076 = n6863 & ~n35978;
  assign n36077 = pi38 & ~n36076;
  assign n36078 = pi38 & ~n36075;
  assign n36079 = ~n36076 & n36078;
  assign n36080 = ~n36075 & n36077;
  assign n36081 = ~n36074 & ~n60466;
  assign n36082 = n59928 & ~n36081;
  assign n36083 = ~pi221 & ~n59928;
  assign po378 = ~n36082 & ~n36083;
  assign n36085 = n59928 & ~n28309;
  assign n36086 = pi829 & pi1091;
  assign n36087 = ~pi824 & ~n36086;
  assign n36088 = n2441 & ~n36087;
  assign n36089 = n6384 & ~n36088;
  assign n36090 = n6438 & n36086;
  assign n36091 = ~n59145 & ~n36090;
  assign n36092 = pi824 & ~n6431;
  assign n36093 = n6439 & n36086;
  assign n36094 = ~pi824 & ~n36093;
  assign n36095 = ~n28510 & ~n36094;
  assign n36096 = ~n36092 & n36095;
  assign n36097 = ~n28510 & ~n36092;
  assign n36098 = ~n36094 & n36097;
  assign n36099 = ~n28510 & ~n36091;
  assign n36100 = ~n36089 & ~n60467;
  assign n36101 = n60122 & ~n36100;
  assign n36102 = ~n2727 & n6384;
  assign n36103 = ~n6409 & ~n36102;
  assign n36104 = ~n28510 & ~n60122;
  assign n36105 = ~n36103 & n36104;
  assign n36106 = n6384 & n28510;
  assign n36107 = pi1093 & ~n36106;
  assign n36108 = ~n36105 & n36107;
  assign n36109 = ~n6384 & ~n60467;
  assign n36110 = ~n36104 & ~n36109;
  assign n36111 = pi1093 & ~n36105;
  assign n36112 = ~n36110 & n36111;
  assign n36113 = ~n36101 & n36108;
  assign n36114 = ~n2443 & n6384;
  assign n36115 = n58823 & n59139;
  assign n36116 = n59138 & n6362;
  assign n36117 = ~n6372 & n60469;
  assign n36118 = ~pi40 & ~n36117;
  assign n36119 = n6316 & ~n36118;
  assign n36120 = pi252 & ~n36119;
  assign n36121 = n2443 & ~n6357;
  assign n36122 = ~n36120 & n36121;
  assign n36123 = ~pi1093 & ~n36122;
  assign n36124 = ~n36114 & n36123;
  assign n36125 = ~pi39 & ~n36124;
  assign n36126 = ~n60468 & n36125;
  assign n36127 = ~n2442 & n2726;
  assign n36128 = n6551 & n36127;
  assign n36129 = n6460 & ~n36127;
  assign n36130 = pi1091 & ~n36129;
  assign n36131 = pi1091 & ~n36128;
  assign n36132 = ~n36129 & n36131;
  assign n36133 = ~n36128 & n36130;
  assign n36134 = ~n2862 & n6460;
  assign n36135 = n2862 & n6551;
  assign n36136 = ~pi1091 & ~n36135;
  assign n36137 = ~pi1091 & ~n36134;
  assign n36138 = ~n36135 & n36137;
  assign n36139 = ~n36134 & n36136;
  assign n36140 = ~n60470 & ~n60471;
  assign n36141 = ~pi120 & ~n36140;
  assign n36142 = ~n6462 & ~n36141;
  assign n36143 = ~n2822 & n36142;
  assign n36144 = ~n35515 & ~n36143;
  assign n36145 = ~n2790 & n36144;
  assign n36146 = ~n2783 & n6463;
  assign n36147 = n2783 & n36142;
  assign n36148 = ~n36146 & ~n36147;
  assign n36149 = n2790 & n36148;
  assign n36150 = ~n6544 & ~n36149;
  assign n36151 = ~n6544 & ~n36145;
  assign n36152 = ~n36149 & n36151;
  assign n36153 = ~n36145 & n36150;
  assign n36154 = ~pi223 & ~n6622;
  assign n36155 = ~n60472 & n36154;
  assign n36156 = pi120 & n31510;
  assign n36157 = n6463 & ~n36156;
  assign n36158 = ~n36146 & ~n36157;
  assign n36159 = n2790 & ~n36158;
  assign n36160 = ~n35515 & ~n36157;
  assign n36161 = ~n2790 & ~n36160;
  assign n36162 = pi223 & ~n36161;
  assign n36163 = ~n36159 & n36162;
  assign n36164 = ~pi299 & ~n36163;
  assign n36165 = ~n36155 & n36164;
  assign n36166 = ~n58846 & n36144;
  assign n36167 = n58846 & n36148;
  assign n36168 = ~n6629 & ~n36167;
  assign n36169 = ~n6629 & ~n36166;
  assign n36170 = ~n36167 & n36169;
  assign n36171 = ~n36166 & n36168;
  assign n36172 = ~pi215 & ~n6821;
  assign n36173 = ~n60473 & n36172;
  assign n36174 = n58846 & ~n36158;
  assign n36175 = ~n58846 & ~n36160;
  assign n36176 = pi215 & ~n36175;
  assign n36177 = ~n36174 & n36176;
  assign n36178 = pi299 & ~n36177;
  assign n36179 = ~n36173 & n36178;
  assign n36180 = ~n36165 & ~n36179;
  assign n36181 = pi39 & ~n36180;
  assign n36182 = ~pi38 & ~n36181;
  assign n36183 = ~n36126 & n36182;
  assign po387 = n36085 & ~n36183;
  assign n36185 = ~n6550 & n60240;
  assign n36186 = pi1093 & n36185;
  assign n36187 = n2801 & n2805;
  assign n36188 = ~n36186 & n36187;
  assign n36189 = ~pi223 & n36188;
  assign n36190 = n2783 & n36185;
  assign n36191 = n36187 & ~n36190;
  assign n36192 = n2790 & n36191;
  assign n36193 = ~n2822 & n36185;
  assign n36194 = n36187 & ~n36193;
  assign n36195 = ~n2790 & n36194;
  assign n36196 = ~pi299 & ~n36195;
  assign n36197 = ~pi299 & ~n36192;
  assign n36198 = ~n36195 & n36197;
  assign n36199 = ~n36192 & n36196;
  assign n36200 = ~n36189 & n60474;
  assign n36201 = ~pi215 & n36188;
  assign n36202 = n58846 & n36191;
  assign n36203 = ~n58846 & n36194;
  assign n36204 = pi299 & ~n36203;
  assign n36205 = pi299 & ~n36202;
  assign n36206 = ~n36203 & n36205;
  assign n36207 = ~n36202 & n36204;
  assign n36208 = ~n36201 & n60475;
  assign n36209 = pi786 & ~pi1082;
  assign n36210 = ~n36208 & ~n36209;
  assign n36211 = ~n36200 & ~n36209;
  assign n36212 = ~n36208 & n36211;
  assign n36213 = ~n36200 & n36210;
  assign n36214 = ~n2845 & n2851;
  assign n36215 = ~n35605 & ~n36214;
  assign n36216 = po740 & n36209;
  assign n36217 = ~n36215 & n36216;
  assign n36218 = n2807 & n36217;
  assign n36219 = ~n60476 & ~n36218;
  assign n36220 = pi39 & ~n36219;
  assign n36221 = n28441 & n60122;
  assign n36222 = n2490 & n31410;
  assign n36223 = n2491 & ~n31409;
  assign n36224 = ~pi89 & ~pi102;
  assign n36225 = n2471 & n36224;
  assign n36226 = n2470 & n6320;
  assign n36227 = n36225 & n36226;
  assign n36228 = n29130 & n36227;
  assign n36229 = ~pi65 & ~pi69;
  assign n36230 = n6319 & n36229;
  assign n36231 = pi48 & ~pi49;
  assign n36232 = ~pi68 & ~pi82;
  assign n36233 = n36231 & n36232;
  assign n36234 = n35623 & n36233;
  assign n36235 = n36230 & n36234;
  assign n36236 = n36228 & n36235;
  assign n36237 = n35621 & n36236;
  assign n36238 = ~pi841 & n2489;
  assign n36239 = n2501 & n36238;
  assign n36240 = ~pi841 & n2507;
  assign n36241 = ~pi97 & n60478;
  assign n36242 = n36237 & n36241;
  assign n36243 = n60477 & n36242;
  assign n36244 = ~pi47 & ~n6369;
  assign n36245 = ~n36243 & n36244;
  assign n36246 = ~pi986 & ~po740;
  assign n36247 = pi252 & ~n36246;
  assign n36248 = pi314 & ~n36247;
  assign n36249 = n6362 & n36248;
  assign n36250 = ~n36245 & n36249;
  assign n36251 = ~pi47 & ~pi841;
  assign n36252 = n36237 & n36251;
  assign n36253 = ~n6358 & ~n36252;
  assign n36254 = n58791 & n2530;
  assign n36255 = ~n36248 & n36254;
  assign n36256 = ~n36253 & n36255;
  assign n36257 = ~n36250 & ~n36256;
  assign n36258 = n2579 & ~n36257;
  assign n36259 = ~pi35 & ~n36258;
  assign n36260 = n2620 & n6377;
  assign n36261 = ~n36259 & n36260;
  assign n36262 = ~n36221 & ~n36261;
  assign n36263 = n6860 & ~n36262;
  assign n36264 = ~n36220 & ~n36263;
  assign po197 = n32632 & ~n36264;
  assign n36266 = pi39 & ~n32621;
  assign n36267 = ~pi314 & pi1050;
  assign n36268 = n60166 & n36267;
  assign n36269 = ~pi39 & ~n36268;
  assign n36270 = n32632 & ~n36269;
  assign n36271 = pi39 & n32621;
  assign n36272 = ~pi39 & n36267;
  assign n36273 = n60166 & n36272;
  assign n36274 = ~n36271 & ~n36273;
  assign n36275 = n32632 & ~n36274;
  assign n36276 = ~n36266 & n36270;
  assign n36277 = pi72 & n35616;
  assign n36278 = pi88 & n60262;
  assign n36279 = n59138 & n60081;
  assign n36280 = n36278 & n36279;
  assign n36281 = n6389 & n36278;
  assign n36282 = n36279 & n36281;
  assign n36283 = n6389 & n36280;
  assign n36284 = ~n36277 & ~n60480;
  assign n36285 = n2621 & ~n36284;
  assign n36286 = ~pi39 & ~n36285;
  assign n36287 = n58845 & n32615;
  assign n36288 = n58848 & n32618;
  assign n36289 = pi39 & ~n36288;
  assign n36290 = ~n36287 & n36289;
  assign n36291 = n32632 & ~n36290;
  assign po230 = ~n36286 & n36291;
  assign n36293 = ~pi100 & n25479;
  assign n36294 = n6310 & n36293;
  assign n36295 = ~n30821 & n36294;
  assign n36296 = n58847 & n60188;
  assign n36297 = n58843 & n60187;
  assign n36298 = ~n36296 & ~n36297;
  assign n36299 = n36294 & ~n36298;
  assign n36300 = n58842 & n36295;
  assign n36301 = pi92 & n58822;
  assign n36302 = n60069 & n36267;
  assign n36303 = n36301 & n36302;
  assign n36304 = ~n60481 & ~n36303;
  assign po250 = n32859 & ~n36304;
  assign n36306 = ~pi39 & pi228;
  assign n36307 = ~n60433 & ~n60436;
  assign n36308 = pi39 & ~n36307;
  assign n36309 = n28516 & n36308;
  assign n36310 = ~pi96 & ~n35646;
  assign n36311 = pi96 & ~n31406;
  assign n36312 = n2597 & ~n36311;
  assign n36313 = ~n2797 & ~n35648;
  assign n36314 = n32908 & ~n36313;
  assign n36315 = n36312 & n36314;
  assign n36316 = ~n36310 & n36315;
  assign n36317 = ~n36309 & ~n36316;
  assign n36318 = n32632 & ~n36317;
  assign n36319 = ~n36306 & ~n36318;
  assign n36320 = pi207 & pi208;
  assign n36321 = ~pi115 & n2793;
  assign n36322 = pi42 & ~pi114;
  assign n36323 = pi72 & pi116;
  assign n36324 = pi72 & pi113;
  assign n36325 = pi72 & ~n2693;
  assign n36326 = ~pi72 & pi101;
  assign n36327 = ~pi41 & ~n36326;
  assign n36328 = pi44 & pi72;
  assign n36329 = n2625 & ~n2628;
  assign n36330 = ~pi72 & ~n58811;
  assign n36331 = ~n2613 & n36330;
  assign n36332 = ~pi1093 & ~n36331;
  assign n36333 = ~n36329 & n36332;
  assign n36334 = n58811 & ~n2613;
  assign n36335 = ~pi122 & n28642;
  assign n36336 = n58813 & ~n28641;
  assign n36337 = ~n36334 & ~n60482;
  assign n36338 = ~pi72 & n36337;
  assign n36339 = pi1093 & ~n36338;
  assign n36340 = ~n36333 & ~n36339;
  assign n36341 = ~pi44 & ~n36340;
  assign n36342 = ~n36328 & ~n36341;
  assign n36343 = ~pi101 & n36342;
  assign n36344 = n36327 & ~n36343;
  assign n36345 = ~pi99 & n36344;
  assign n36346 = ~n36325 & ~n36345;
  assign n36347 = ~pi113 & ~n36346;
  assign n36348 = ~n36324 & ~n36347;
  assign n36349 = ~pi116 & ~n36348;
  assign n36350 = ~n36323 & ~n36349;
  assign n36351 = n36322 & ~n36350;
  assign n36352 = pi42 & ~pi72;
  assign n36353 = pi114 & ~n36352;
  assign n36354 = ~pi1093 & ~n36334;
  assign n36355 = ~pi1093 & ~n58814;
  assign n36356 = ~n36334 & n36355;
  assign n36357 = ~n58814 & n36354;
  assign n36358 = ~pi44 & ~n60483;
  assign n36359 = pi1093 & n36337;
  assign n36360 = n36358 & ~n36359;
  assign n36361 = ~pi101 & n36360;
  assign n36362 = n2693 & n36361;
  assign n36363 = n2695 & n36362;
  assign n36364 = ~pi42 & ~n36363;
  assign n36365 = ~n36353 & ~n36364;
  assign n36366 = ~n36351 & n36365;
  assign n36367 = n36321 & ~n36366;
  assign n36368 = n36330 & ~n36333;
  assign n36369 = ~pi44 & ~n36368;
  assign n36370 = ~n36328 & ~n36369;
  assign n36371 = ~pi101 & n36370;
  assign n36372 = n36327 & ~n36371;
  assign n36373 = ~pi99 & n36372;
  assign n36374 = ~n36325 & ~n36373;
  assign n36375 = ~pi113 & ~n36374;
  assign n36376 = ~n36324 & ~n36375;
  assign n36377 = ~pi116 & ~n36376;
  assign n36378 = ~n36323 & ~n36377;
  assign n36379 = pi42 & n36378;
  assign n36380 = pi1093 & ~n58811;
  assign n36381 = n36358 & ~n36380;
  assign n36382 = ~pi101 & n36381;
  assign n36383 = n2693 & n36382;
  assign n36384 = n2695 & n36383;
  assign n36385 = ~pi42 & n36384;
  assign n36386 = ~pi114 & ~n36385;
  assign n36387 = ~n36379 & n36386;
  assign n36388 = ~n36353 & ~n36387;
  assign n36389 = ~pi115 & ~n2793;
  assign n36390 = ~n36388 & n36389;
  assign n36391 = pi115 & ~n36352;
  assign n36392 = pi228 & ~n36391;
  assign n36393 = ~n36390 & n36392;
  assign n36394 = ~n36367 & n36393;
  assign n36395 = n2539 & n31412;
  assign n36396 = ~pi110 & ~n36395;
  assign n36397 = n2530 & ~n31469;
  assign n36398 = ~pi480 & pi949;
  assign n36399 = n60073 & n36398;
  assign n36400 = ~pi47 & n36399;
  assign n36401 = n36397 & n36400;
  assign n36402 = ~n36396 & n36401;
  assign n36403 = pi901 & ~pi959;
  assign n36404 = n58798 & n31412;
  assign n36405 = n60073 & ~n36398;
  assign n36406 = n60073 & n36404;
  assign n36407 = ~n36398 & n36406;
  assign n36408 = n36404 & n36405;
  assign n36409 = n36403 & ~n60484;
  assign n36410 = ~n36402 & n36403;
  assign n36411 = ~n60484 & n36410;
  assign n36412 = ~n36402 & n36409;
  assign n36413 = pi110 & n32498;
  assign n36414 = n36399 & n36413;
  assign n36415 = ~n36403 & ~n36414;
  assign n36416 = ~pi250 & pi252;
  assign n36417 = n2621 & n36416;
  assign n36418 = ~n36415 & n36417;
  assign n36419 = ~n60485 & n36418;
  assign n36420 = n2621 & ~n36416;
  assign n36421 = n36414 & n36420;
  assign n36422 = ~pi72 & ~n36421;
  assign n36423 = ~n36419 & n36422;
  assign n36424 = ~pi44 & ~n36423;
  assign n36425 = ~n36328 & ~n36424;
  assign n36426 = ~pi101 & n36425;
  assign n36427 = n36327 & ~n36426;
  assign n36428 = ~pi99 & n36427;
  assign n36429 = ~n36325 & ~n36428;
  assign n36430 = ~pi113 & ~n36429;
  assign n36431 = ~n36324 & ~n36430;
  assign n36432 = ~pi116 & ~n36431;
  assign n36433 = ~n36323 & ~n36432;
  assign n36434 = n36322 & ~n36433;
  assign n36435 = ~pi72 & n36419;
  assign n36436 = n60165 & n36413;
  assign n36437 = n36398 & ~n36416;
  assign n36438 = n36436 & n36437;
  assign n36439 = ~n36435 & ~n36438;
  assign n36440 = ~pi44 & ~n36439;
  assign n36441 = ~pi101 & n36440;
  assign n36442 = n2693 & n36441;
  assign n36443 = ~pi113 & n36442;
  assign n36444 = ~pi116 & n36443;
  assign n36445 = n2695 & n36442;
  assign n36446 = ~pi42 & ~n60486;
  assign n36447 = ~n36353 & ~n36446;
  assign n36448 = ~n36434 & n36447;
  assign n36449 = ~pi115 & ~n36448;
  assign n36450 = ~pi228 & ~n36391;
  assign n36451 = ~n36449 & n36450;
  assign n36452 = ~pi39 & ~n36451;
  assign n36453 = ~n36394 & n36452;
  assign n36454 = ~pi72 & ~n30128;
  assign n36455 = pi287 & n58822;
  assign n36456 = n2680 & n36455;
  assign n36457 = pi287 & n29911;
  assign n36458 = ~pi189 & n60487;
  assign n36459 = n30128 & n36455;
  assign n36460 = ~n36454 & ~n60488;
  assign n36461 = pi199 & ~n36460;
  assign n36462 = pi232 & ~n36461;
  assign n36463 = ~pi299 & n36462;
  assign n36464 = n32622 & ~n36461;
  assign n36465 = ~pi166 & n60487;
  assign n36466 = n29998 & n36455;
  assign n36467 = pi232 & n29998;
  assign n36468 = ~pi166 & n2681;
  assign n36469 = ~pi72 & ~n60491;
  assign n36470 = n32792 & ~n36469;
  assign n36471 = ~n60490 & n36470;
  assign n36472 = ~pi72 & pi199;
  assign n36473 = ~pi232 & ~n36472;
  assign n36474 = pi72 & ~pi232;
  assign n36475 = pi299 & ~n36474;
  assign n36476 = n36473 & ~n36475;
  assign n36477 = ~n36471 & ~n36476;
  assign n36478 = ~n60489 & n36477;
  assign n36479 = pi39 & ~n36478;
  assign n36480 = ~n36453 & ~n36479;
  assign n36481 = n2636 & ~n36480;
  assign n36482 = ~n2719 & ~n36352;
  assign n36483 = ~n36321 & n36352;
  assign n36484 = n2719 & ~n36483;
  assign n36485 = n36321 & ~n36353;
  assign n36486 = ~pi44 & n58822;
  assign n36487 = ~pi101 & n36486;
  assign n36488 = n2693 & n36487;
  assign n36489 = n2695 & n36488;
  assign n36490 = n2715 & n36489;
  assign n36491 = ~pi114 & ~n2702;
  assign n36492 = n36490 & n36491;
  assign n36493 = ~pi42 & n36492;
  assign n36494 = ~pi72 & ~n2715;
  assign n36495 = n2621 & n28317;
  assign n36496 = ~pi44 & n36495;
  assign n36497 = n2694 & n36496;
  assign n36498 = n2695 & n36497;
  assign n36499 = ~pi72 & ~n36498;
  assign n36500 = ~n36494 & ~n36499;
  assign n36501 = pi42 & ~n36500;
  assign n36502 = ~pi114 & ~n36501;
  assign n36503 = ~pi114 & ~n36493;
  assign n36504 = ~n36501 & n36503;
  assign n36505 = ~n36493 & n36502;
  assign n36506 = n36485 & ~n60492;
  assign n36507 = n36484 & ~n36506;
  assign n36508 = ~n36482 & ~n36507;
  assign n36509 = ~pi39 & ~n36508;
  assign n36510 = ~pi299 & ~n36473;
  assign n36511 = pi199 & n36454;
  assign n36512 = pi232 & ~n36511;
  assign n36513 = n36510 & ~n36512;
  assign n36514 = pi299 & n36469;
  assign n36515 = pi39 & ~n36514;
  assign n36516 = ~n36513 & n36515;
  assign n36517 = ~n36509 & ~n36516;
  assign n36518 = n28548 & ~n36517;
  assign n36519 = ~pi39 & ~n36352;
  assign n36520 = ~n36516 & ~n36519;
  assign n36521 = pi38 & ~n36520;
  assign n36522 = ~pi87 & ~n36521;
  assign n36523 = ~n36518 & n36522;
  assign n36524 = ~n36481 & n36523;
  assign n36525 = ~pi42 & n2698;
  assign n36526 = pi228 & n36525;
  assign n36527 = pi228 & n36489;
  assign n36528 = ~pi115 & n36527;
  assign n36529 = ~pi114 & n36528;
  assign n36530 = n2698 & n36527;
  assign n36531 = ~pi42 & n60493;
  assign n36532 = n36489 & n36526;
  assign n36533 = pi228 & n36497;
  assign n36534 = pi228 & n36498;
  assign n36535 = ~pi115 & n36534;
  assign n36536 = ~pi114 & n36535;
  assign n36537 = n2703 & n36533;
  assign n36538 = n36352 & ~n60495;
  assign n36539 = n58815 & ~n36538;
  assign n36540 = n58815 & ~n60494;
  assign n36541 = ~n36538 & n36540;
  assign n36542 = ~n60494 & n36539;
  assign n36543 = ~n2636 & n36519;
  assign n36544 = pi87 & ~n36543;
  assign n36545 = ~n60496 & n36544;
  assign n36546 = ~n36516 & n36545;
  assign n36547 = ~pi75 & ~n36546;
  assign n36548 = ~n36524 & n36547;
  assign n36549 = n58827 & n36492;
  assign n36550 = ~pi42 & n36549;
  assign n36551 = n58827 & n36493;
  assign n36552 = ~pi24 & n28317;
  assign n36553 = n2684 & n2715;
  assign n36554 = n36552 & n36553;
  assign n36555 = ~pi44 & n36554;
  assign n36556 = n2694 & n36555;
  assign n36557 = ~pi113 & n36556;
  assign n36558 = ~pi116 & n36557;
  assign n36559 = n36352 & ~n36558;
  assign n36560 = ~pi114 & ~n36559;
  assign n36561 = ~pi114 & ~n60497;
  assign n36562 = ~n36559 & n36561;
  assign n36563 = ~n60497 & n36560;
  assign n36564 = n36485 & ~n60498;
  assign n36565 = n36484 & ~n36564;
  assign n36566 = n59291 & ~n36482;
  assign n36567 = ~n36565 & n36566;
  assign n36568 = ~n59291 & n36352;
  assign n36569 = ~pi39 & ~n36568;
  assign n36570 = ~n36567 & n36569;
  assign n36571 = ~n36516 & ~n36570;
  assign n36572 = pi75 & ~n36571;
  assign n36573 = n2439 & ~n36572;
  assign n36574 = ~n36548 & n36573;
  assign n36575 = ~n36320 & ~n36574;
  assign n36576 = ~pi72 & pi200;
  assign n36577 = ~pi232 & ~n36576;
  assign n36578 = ~pi299 & ~n36577;
  assign n36579 = pi200 & n36454;
  assign n36580 = pi232 & ~n36579;
  assign n36581 = n36578 & ~n36580;
  assign n36582 = pi39 & ~n36581;
  assign n36583 = ~n36513 & n36582;
  assign n36584 = ~n36519 & ~n36583;
  assign n36585 = ~n2439 & n36584;
  assign n36586 = n36320 & ~n36585;
  assign n36587 = pi200 & ~n36460;
  assign n36588 = pi232 & ~n36587;
  assign n36589 = ~pi299 & n36588;
  assign n36590 = n32622 & ~n36587;
  assign n36591 = n36462 & ~n36587;
  assign n36592 = ~n36461 & n36588;
  assign n36593 = ~pi299 & n60500;
  assign n36594 = ~n36461 & n60499;
  assign n36595 = n36476 & ~n36576;
  assign n36596 = ~n36471 & ~n36595;
  assign n36597 = ~n60501 & n36596;
  assign n36598 = pi39 & ~n36597;
  assign n36599 = ~n36453 & ~n36598;
  assign n36600 = n2636 & ~n36599;
  assign n36601 = pi38 & ~n36584;
  assign n36602 = ~pi87 & ~n36601;
  assign n36603 = ~n36522 & ~n36602;
  assign n36604 = n36516 & n36582;
  assign n36605 = ~n36509 & ~n36604;
  assign n36606 = n28548 & ~n36605;
  assign n36607 = ~n36603 & ~n36606;
  assign n36608 = ~n36600 & n36607;
  assign n36609 = n36544 & ~n36604;
  assign n36610 = n36545 & ~n36604;
  assign n36611 = ~n60496 & n36609;
  assign n36612 = ~pi75 & ~n60502;
  assign n36613 = ~n36608 & n36612;
  assign n36614 = ~n36570 & ~n36604;
  assign n36615 = pi75 & ~n36614;
  assign n36616 = n2439 & ~n36615;
  assign n36617 = ~n36613 & n36616;
  assign n36618 = n36586 & ~n36617;
  assign n36619 = ~n36575 & ~n36618;
  assign n36620 = pi211 & pi214;
  assign n36621 = pi212 & pi214;
  assign n36622 = pi211 & n36621;
  assign n36623 = pi212 & n36620;
  assign n36624 = ~pi219 & ~n60503;
  assign n36625 = ~n2439 & n36520;
  assign n36626 = ~n36624 & ~n36625;
  assign n36627 = ~n36619 & n36626;
  assign n36628 = ~n36462 & n36510;
  assign n36629 = pi39 & ~n36628;
  assign n36630 = ~n36453 & ~n36629;
  assign n36631 = n2636 & ~n36630;
  assign n36632 = pi39 & ~n36513;
  assign n36633 = ~n36509 & ~n36632;
  assign n36634 = n28548 & ~n36633;
  assign n36635 = ~n36519 & ~n36632;
  assign n36636 = pi38 & ~n36635;
  assign n36637 = ~pi87 & ~n36636;
  assign n36638 = ~n36634 & n36637;
  assign n36639 = ~n36631 & n36638;
  assign n36640 = n36545 & ~n36632;
  assign n36641 = ~pi75 & ~n36640;
  assign n36642 = ~n36639 & n36641;
  assign n36643 = ~n36570 & ~n36632;
  assign n36644 = pi75 & ~n36643;
  assign n36645 = n2439 & ~n36644;
  assign n36646 = ~n36642 & n36645;
  assign n36647 = ~n2439 & n36635;
  assign n36648 = ~n36320 & ~n36647;
  assign n36649 = ~n36646 & n36648;
  assign n36650 = ~n36510 & ~n36578;
  assign n36651 = ~n60500 & ~n36650;
  assign n36652 = pi39 & ~n36651;
  assign n36653 = ~n36453 & ~n36652;
  assign n36654 = n2636 & ~n36653;
  assign n36655 = ~n36509 & ~n36583;
  assign n36656 = n28548 & ~n36655;
  assign n36657 = n36602 & ~n36656;
  assign n36658 = ~n36654 & n36657;
  assign n36659 = n36545 & ~n36583;
  assign n36660 = ~pi75 & ~n36659;
  assign n36661 = ~n36658 & n36660;
  assign n36662 = ~n36570 & ~n36583;
  assign n36663 = pi75 & ~n36662;
  assign n36664 = n2439 & ~n36663;
  assign n36665 = ~n36661 & n36664;
  assign n36666 = n36586 & ~n36665;
  assign n36667 = ~n36649 & ~n36666;
  assign n36668 = n36624 & ~n36667;
  assign n36669 = n58992 & ~n36668;
  assign n36670 = n58992 & ~n36627;
  assign n36671 = ~n36668 & n36670;
  assign n36672 = ~n36627 & n36669;
  assign n36673 = n36469 & ~n36624;
  assign n36674 = pi39 & ~n36673;
  assign n36675 = ~n58992 & ~n36519;
  assign n36676 = ~n36674 & n36675;
  assign n36677 = ~n60504 & ~n36676;
  assign n36678 = ~pi211 & ~n36621;
  assign n36679 = ~pi211 & ~pi219;
  assign n36680 = n36621 & ~n36679;
  assign n36681 = ~pi211 & pi219;
  assign n36682 = ~n60503 & ~n36678;
  assign n36683 = ~n36681 & n36682;
  assign n36684 = pi211 & ~n36621;
  assign n36685 = n36621 & n36679;
  assign n36686 = ~n36684 & ~n36685;
  assign n36687 = ~n36678 & ~n36680;
  assign n36688 = ~n2793 & ~n36383;
  assign n36689 = n2793 & ~n36362;
  assign n36690 = ~n36688 & ~n36689;
  assign n36691 = pi228 & ~n36690;
  assign n36692 = ~pi228 & ~n36442;
  assign n36693 = n2695 & ~n36692;
  assign n36694 = n2793 & n36363;
  assign n36695 = ~n2793 & n36384;
  assign n36696 = pi228 & ~n36695;
  assign n36697 = n2695 & n36690;
  assign n36698 = pi228 & ~n36697;
  assign n36699 = ~n36694 & n36696;
  assign n36700 = ~pi228 & ~n60486;
  assign n36701 = ~n60506 & ~n36700;
  assign n36702 = ~n36691 & n36693;
  assign n36703 = ~pi43 & ~n60507;
  assign n36704 = pi43 & ~pi72;
  assign n36705 = ~n36525 & ~n36704;
  assign n36706 = n36525 & ~n36703;
  assign n36707 = ~n36704 & ~n36706;
  assign n36708 = ~n36703 & ~n36705;
  assign n36709 = ~pi228 & ~n36433;
  assign n36710 = n2793 & ~n36350;
  assign n36711 = ~n2793 & ~n36378;
  assign n36712 = ~n36710 & ~n36711;
  assign n36713 = pi228 & ~n36712;
  assign n36714 = ~n36709 & ~n36713;
  assign n36715 = pi43 & n36525;
  assign n36716 = ~n36714 & n36715;
  assign n36717 = ~n60508 & ~n36716;
  assign n36718 = ~pi39 & ~n36717;
  assign n36719 = ~pi199 & ~pi200;
  assign n36720 = ~pi299 & ~n36719;
  assign n36721 = ~pi72 & ~n36720;
  assign n36722 = ~pi232 & ~n36721;
  assign n36723 = ~pi299 & ~n36722;
  assign n36724 = ~n36460 & n36719;
  assign n36725 = pi232 & ~n36724;
  assign n36726 = n36723 & ~n36725;
  assign n36727 = pi39 & ~n36726;
  assign n36728 = ~n36718 & ~n36727;
  assign n36729 = n2636 & ~n36728;
  assign n36730 = ~n2719 & ~n36704;
  assign n36731 = n2793 & n36525;
  assign n36732 = n36704 & ~n36731;
  assign n36733 = n2719 & ~n36732;
  assign n36734 = ~pi43 & pi52;
  assign n36735 = n36490 & n36734;
  assign n36736 = pi43 & ~n36500;
  assign n36737 = ~n36735 & ~n36736;
  assign n36738 = n36731 & ~n36737;
  assign n36739 = n36733 & ~n36738;
  assign n36740 = ~n36730 & ~n36739;
  assign n36741 = ~pi39 & ~n36740;
  assign n36742 = n36454 & n36719;
  assign n36743 = pi232 & ~n36742;
  assign n36744 = n36723 & ~n36743;
  assign n36745 = pi39 & ~n36744;
  assign n36746 = ~n36741 & ~n36745;
  assign n36747 = n28548 & ~n36746;
  assign n36748 = ~pi39 & ~n36704;
  assign n36749 = ~n36745 & ~n36748;
  assign n36750 = pi38 & ~n36749;
  assign n36751 = ~pi87 & ~n36750;
  assign n36752 = ~n36747 & n36751;
  assign n36753 = ~n36729 & n36752;
  assign n36754 = ~pi43 & ~n36489;
  assign n36755 = pi43 & ~n36499;
  assign n36756 = n36526 & ~n36755;
  assign n36757 = ~n36754 & n36756;
  assign n36758 = ~n36526 & n36704;
  assign n36759 = n58815 & ~n36758;
  assign n36760 = ~pi42 & n60495;
  assign n36761 = n36704 & ~n36760;
  assign n36762 = n2699 & n36528;
  assign n36763 = n58815 & ~n36762;
  assign n36764 = ~n36761 & n36763;
  assign n36765 = ~n36757 & n36759;
  assign n36766 = ~n2636 & n36748;
  assign n36767 = pi87 & ~n36766;
  assign n36768 = ~n60509 & n36767;
  assign n36769 = ~n58815 & ~n36749;
  assign n36770 = n36768 & ~n36769;
  assign n36771 = ~pi75 & ~n36770;
  assign n36772 = ~n36753 & n36771;
  assign n36773 = ~pi72 & ~n36558;
  assign n36774 = pi43 & n36773;
  assign n36775 = n58827 & n36490;
  assign n36776 = n36734 & n36775;
  assign n36777 = ~n36774 & ~n36776;
  assign n36778 = n36731 & ~n36777;
  assign n36779 = n36733 & ~n36778;
  assign n36780 = n59291 & ~n36730;
  assign n36781 = ~n36779 & n36780;
  assign n36782 = ~n59291 & n36704;
  assign n36783 = ~pi39 & ~n36782;
  assign n36784 = ~n36730 & ~n36779;
  assign n36785 = ~pi39 & ~n36784;
  assign n36786 = n59291 & ~n36785;
  assign n36787 = ~n59291 & ~n36748;
  assign n36788 = ~n36786 & ~n36787;
  assign n36789 = ~n36781 & n36783;
  assign n36790 = ~n36745 & ~n60510;
  assign n36791 = pi75 & ~n36790;
  assign n36792 = n2439 & ~n36791;
  assign n36793 = ~n36772 & n36792;
  assign n36794 = ~n2439 & n36749;
  assign n36795 = n36320 & ~n36794;
  assign n36796 = ~n36793 & n36795;
  assign n36797 = n36578 & ~n36588;
  assign n36798 = pi39 & ~n36797;
  assign n36799 = ~n36718 & ~n36798;
  assign n36800 = n2636 & ~n36799;
  assign n36801 = ~n36582 & ~n36741;
  assign n36802 = n28548 & ~n36801;
  assign n36803 = ~n36582 & ~n36748;
  assign n36804 = pi38 & ~n36803;
  assign n36805 = ~pi87 & ~n36804;
  assign n36806 = ~n36802 & n36805;
  assign n36807 = ~n36800 & n36806;
  assign n36808 = ~n36582 & n36768;
  assign n36809 = ~pi75 & ~n36808;
  assign n36810 = ~n36807 & n36809;
  assign n36811 = ~n36582 & ~n60510;
  assign n36812 = pi75 & ~n36811;
  assign n36813 = n2439 & ~n36812;
  assign n36814 = ~n36810 & n36813;
  assign n36815 = ~n2439 & n36803;
  assign n36816 = ~n36320 & ~n36815;
  assign n36817 = ~n36814 & n36816;
  assign n36818 = ~n36796 & ~n36817;
  assign n36819 = ~n60505 & ~n36818;
  assign n36820 = ~n36475 & n36577;
  assign n36821 = ~n36471 & ~n36820;
  assign n36822 = ~n60499 & n36821;
  assign n36823 = pi39 & ~n36822;
  assign n36824 = ~n36718 & ~n36823;
  assign n36825 = n2636 & ~n36824;
  assign n36826 = n36515 & ~n36581;
  assign n36827 = ~n36741 & ~n36826;
  assign n36828 = n28548 & ~n36827;
  assign n36829 = ~n36748 & ~n36826;
  assign n36830 = pi38 & ~n36829;
  assign n36831 = ~pi87 & ~n36830;
  assign n36832 = ~n36828 & n36831;
  assign n36833 = ~n36825 & n36832;
  assign n36834 = n36768 & ~n36826;
  assign n36835 = ~pi75 & ~n36834;
  assign n36836 = ~n36833 & n36835;
  assign n36837 = ~n60510 & ~n36826;
  assign n36838 = pi75 & ~n36837;
  assign n36839 = n2439 & ~n36838;
  assign n36840 = ~n36836 & n36839;
  assign n36841 = ~n2439 & n36829;
  assign n36842 = ~n36320 & ~n36841;
  assign n36843 = ~n36840 & n36842;
  assign n36844 = n32622 & ~n36724;
  assign n36845 = ~n36471 & ~n36722;
  assign n36846 = ~n36844 & n36845;
  assign n36847 = pi39 & ~n36846;
  assign n36848 = ~n36718 & ~n36847;
  assign n36849 = n2636 & ~n36848;
  assign n36850 = ~n36514 & n36745;
  assign n36851 = ~n36741 & ~n36850;
  assign n36852 = n28548 & ~n36851;
  assign n36853 = ~n36748 & ~n36850;
  assign n36854 = pi38 & ~n36853;
  assign n36855 = ~pi87 & ~n36854;
  assign n36856 = ~n36852 & n36855;
  assign n36857 = ~n36849 & n36856;
  assign n36858 = n36768 & ~n36850;
  assign n36859 = ~pi75 & ~n36858;
  assign n36860 = ~n36857 & n36859;
  assign n36861 = ~n60510 & ~n36850;
  assign n36862 = pi75 & ~n36861;
  assign n36863 = n2439 & ~n36862;
  assign n36864 = ~n36860 & n36863;
  assign n36865 = ~n2439 & n36853;
  assign n36866 = n36320 & ~n36865;
  assign n36867 = ~n36864 & n36866;
  assign n36868 = ~n36843 & ~n36867;
  assign n36869 = n60505 & ~n36868;
  assign n36870 = n58992 & ~n36869;
  assign n36871 = n58992 & ~n36819;
  assign n36872 = ~n36869 & n36871;
  assign n36873 = ~n36819 & n36870;
  assign n36874 = n36469 & n60505;
  assign n36875 = pi39 & ~n36874;
  assign n36876 = ~n58992 & ~n36748;
  assign n36877 = ~n36875 & n36876;
  assign n36878 = ~n60511 & ~n36877;
  assign n36879 = ~pi219 & n36678;
  assign n36880 = ~n36621 & n36679;
  assign n36881 = pi52 & ~pi72;
  assign n36882 = ~pi39 & n36881;
  assign n36883 = pi38 & ~n36882;
  assign n36884 = ~pi43 & n36526;
  assign n36885 = pi228 & n58828;
  assign n36886 = ~pi52 & n36489;
  assign n36887 = pi52 & n36499;
  assign n36888 = ~n36886 & ~n36887;
  assign n36889 = n60513 & ~n36888;
  assign n36890 = n36881 & ~n60513;
  assign n36891 = ~n36889 & ~n36890;
  assign n36892 = ~pi38 & n36891;
  assign n36893 = ~n36883 & ~n36892;
  assign n36894 = ~pi100 & ~n36893;
  assign n36895 = pi100 & ~n36882;
  assign n36896 = pi87 & ~n36293;
  assign n36897 = ~n36895 & n36896;
  assign n36898 = ~n36894 & n36897;
  assign n36899 = pi52 & n36712;
  assign n36900 = n2696 & n36690;
  assign n36901 = n58828 & ~n36900;
  assign n36902 = pi52 & n36350;
  assign n36903 = ~pi52 & n36363;
  assign n36904 = n36321 & ~n36903;
  assign n36905 = ~n36902 & n36904;
  assign n36906 = pi52 & n36378;
  assign n36907 = ~pi52 & n36384;
  assign n36908 = n36389 & ~n36907;
  assign n36909 = ~n36906 & n36908;
  assign n36910 = ~n36905 & ~n36909;
  assign n36911 = n2699 & ~n36910;
  assign n36912 = ~n36899 & n36901;
  assign n36913 = ~n58828 & ~n36881;
  assign n36914 = pi228 & ~n36913;
  assign n36915 = ~n60514 & n36914;
  assign n36916 = pi52 & n36433;
  assign n36917 = ~pi52 & n60486;
  assign n36918 = n58828 & ~n36917;
  assign n36919 = ~n36916 & n36918;
  assign n36920 = ~pi228 & ~n36913;
  assign n36921 = ~n36919 & n36920;
  assign n36922 = ~pi39 & ~n36921;
  assign n36923 = ~n36915 & n36922;
  assign n36924 = ~pi100 & n36923;
  assign n36925 = n2719 & n36321;
  assign n36926 = n2699 & n36925;
  assign n36927 = n2715 & n36926;
  assign n36928 = n36498 & n36927;
  assign n36929 = n36881 & ~n36928;
  assign n36930 = pi100 & ~n36929;
  assign n36931 = ~pi39 & ~n36930;
  assign n36932 = ~n36924 & n36931;
  assign n36933 = ~pi38 & ~n36932;
  assign n36934 = ~pi87 & ~n36883;
  assign n36935 = ~n36933 & n36934;
  assign n36936 = ~n36898 & ~n36935;
  assign n36937 = ~pi75 & ~n36936;
  assign n36938 = n59291 & n36926;
  assign n36939 = n36558 & n36926;
  assign n36940 = n59291 & n36939;
  assign n36941 = n36558 & n36938;
  assign n36942 = n36881 & ~n60515;
  assign n36943 = ~pi39 & pi75;
  assign n36944 = n36882 & ~n60515;
  assign n36945 = pi75 & n36944;
  assign n36946 = n36942 & n36943;
  assign n36947 = n2439 & ~n60516;
  assign n36948 = ~n36937 & n36947;
  assign n36949 = ~n2439 & ~n36882;
  assign n36950 = n36320 & ~n36949;
  assign n36951 = ~n36948 & n36950;
  assign n36952 = ~n36727 & ~n36923;
  assign n36953 = n2636 & ~n36952;
  assign n36954 = ~pi39 & ~n36929;
  assign n36955 = ~n36745 & ~n36954;
  assign n36956 = n28548 & ~n36955;
  assign n36957 = ~pi39 & ~n36881;
  assign n36958 = ~n36745 & ~n36957;
  assign n36959 = pi38 & ~n36958;
  assign n36960 = ~pi87 & ~n36959;
  assign n36961 = ~n36956 & n36960;
  assign n36962 = ~n36953 & n36961;
  assign n36963 = ~n2636 & n36958;
  assign n36964 = ~pi39 & n36891;
  assign n36965 = n2636 & ~n36745;
  assign n36966 = ~n36964 & n36965;
  assign n36967 = ~n36963 & ~n36966;
  assign n36968 = pi87 & ~n36967;
  assign n36969 = ~pi75 & ~n36968;
  assign n36970 = ~n36962 & n36969;
  assign n36971 = n2439 & ~n36320;
  assign n36972 = n36881 & ~n36939;
  assign n36973 = ~pi39 & ~n36972;
  assign n36974 = ~pi87 & n36965;
  assign n36975 = n59291 & ~n36745;
  assign n36976 = ~n36973 & n60517;
  assign n36977 = ~n59291 & n36958;
  assign n36978 = pi75 & ~n36977;
  assign n36979 = ~n36976 & n36978;
  assign n36980 = n36971 & ~n36979;
  assign n36981 = ~n36962 & ~n36968;
  assign n36982 = ~pi75 & ~n36981;
  assign n36983 = ~pi39 & ~n36944;
  assign n36984 = ~pi39 & ~n36942;
  assign n36985 = pi75 & ~n36745;
  assign n36986 = ~n60518 & n36985;
  assign n36987 = ~n36982 & ~n36986;
  assign n36988 = n36971 & ~n36987;
  assign n36989 = ~n36970 & n36980;
  assign n36990 = ~n36951 & ~n60519;
  assign n36991 = ~n60512 & ~n36990;
  assign n36992 = ~n36471 & n36475;
  assign n36993 = pi39 & ~n36992;
  assign n36994 = ~n36923 & ~n36993;
  assign n36995 = n2636 & ~n36994;
  assign n36996 = ~n36515 & ~n36957;
  assign n36997 = pi38 & ~n36996;
  assign n36998 = ~n36515 & ~n36954;
  assign n36999 = n28548 & ~n36998;
  assign n37000 = ~n36997 & ~n36999;
  assign n37001 = ~n36995 & n37000;
  assign n37002 = ~pi87 & ~n37001;
  assign n37003 = ~n2636 & n36996;
  assign n37004 = pi87 & ~n37003;
  assign n37005 = n2636 & ~n36515;
  assign n37006 = ~n36964 & n37005;
  assign n37007 = n37004 & ~n37006;
  assign n37008 = n36320 & ~n37007;
  assign n37009 = ~n37002 & n37008;
  assign n37010 = ~n36847 & ~n36923;
  assign n37011 = n2636 & ~n37010;
  assign n37012 = n36959 & ~n36996;
  assign n37013 = ~n36850 & ~n36954;
  assign n37014 = n28548 & ~n37013;
  assign n37015 = ~n37012 & ~n37014;
  assign n37016 = ~n37011 & n37015;
  assign n37017 = ~pi87 & ~n37016;
  assign n37018 = n2636 & ~n36850;
  assign n37019 = ~n36964 & n37018;
  assign n37020 = ~n36963 & n37004;
  assign n37021 = ~n37019 & n37020;
  assign n37022 = ~n36320 & ~n37021;
  assign n37023 = ~n37017 & n37022;
  assign n37024 = ~n37009 & ~n37023;
  assign n37025 = ~pi75 & ~n37024;
  assign n37026 = ~n36320 & n36744;
  assign n37027 = n36515 & ~n37026;
  assign n37028 = ~n36320 & n36850;
  assign n37029 = n36320 & n36515;
  assign n37030 = pi75 & ~n37029;
  assign n37031 = ~n37028 & n37030;
  assign n37032 = pi75 & ~n37027;
  assign n37033 = ~n60518 & n60520;
  assign n37034 = n2439 & ~n37033;
  assign n37035 = ~n37025 & n37034;
  assign n37036 = ~n2439 & ~n36996;
  assign n37037 = n60512 & ~n37036;
  assign n37038 = ~n37035 & n37037;
  assign n37039 = ~n2439 & ~n36320;
  assign n37040 = n36958 & n37039;
  assign n37041 = n58992 & ~n37040;
  assign n37042 = ~n37038 & n37041;
  assign n37043 = ~n36991 & n37042;
  assign n37044 = pi39 & n60512;
  assign n37045 = n36469 & n37044;
  assign n37046 = ~n58992 & ~n36882;
  assign n37047 = ~n37045 & n37046;
  assign po210 = ~n37043 & ~n37047;
  assign n37049 = n59928 & n25479;
  assign n37050 = pi216 & ~pi221;
  assign n37051 = n2851 & n37050;
  assign n37052 = n32618 & n37051;
  assign n37053 = n2828 & n26651;
  assign n37054 = n32615 & n37053;
  assign n37055 = ~n37052 & ~n37054;
  assign po226 = n37049 & ~n37055;
  assign n37057 = n60262 & n32884;
  assign n37058 = ~pi58 & n2731;
  assign n37059 = ~n37057 & ~n37058;
  assign n37060 = n58838 & n60165;
  assign n37061 = ~n37059 & n37060;
  assign n37062 = pi24 & n2589;
  assign n37063 = ~n58838 & n37062;
  assign n37064 = n32914 & n37063;
  assign n37065 = n2731 & n37064;
  assign n37066 = ~pi39 & ~n37065;
  assign n37067 = ~n37061 & n37066;
  assign n37068 = n59928 & ~n37067;
  assign po249 = n2859 & n37068;
  assign n37070 = n60073 & n28418;
  assign n37071 = ~pi82 & n2452;
  assign n37072 = ~pi84 & pi104;
  assign n37073 = n28346 & n37072;
  assign n37074 = n35624 & n37073;
  assign n37075 = n37071 & n37074;
  assign n37076 = ~pi36 & ~n37075;
  assign n37077 = n58784 & n6324;
  assign n37078 = n2479 & n6325;
  assign n37079 = ~pi67 & ~pi103;
  assign n37080 = n2446 & n37079;
  assign n37081 = ~pi98 & n37080;
  assign n37082 = n60521 & n37081;
  assign n37083 = ~n37076 & n37082;
  assign n37084 = ~pi36 & n37083;
  assign n37085 = ~pi88 & ~n37084;
  assign n37086 = n6391 & ~n37085;
  assign n37087 = n58796 & n6547;
  assign n37088 = n37086 & n37087;
  assign n37089 = ~pi91 & ~n6359;
  assign n37090 = ~n31429 & n37083;
  assign n37091 = ~pi88 & ~n37090;
  assign n37092 = n58796 & ~n37091;
  assign n37093 = n6391 & n37092;
  assign n37094 = ~n2441 & n37093;
  assign n37095 = n37089 & ~n37094;
  assign n37096 = ~n37088 & n37095;
  assign n37097 = n37070 & ~n37096;
  assign n37098 = ~pi72 & ~n37097;
  assign n37099 = n28319 & ~n37098;
  assign n37100 = n31506 & ~n37099;
  assign n37101 = n2727 & n60073;
  assign n37102 = ~n37059 & n37101;
  assign n37103 = n28319 & n37101;
  assign n37104 = ~n37059 & n37103;
  assign n37105 = n28319 & n37102;
  assign n37106 = ~n28505 & ~n60522;
  assign n37107 = pi1093 & ~n37106;
  assign n37108 = n37070 & n37093;
  assign n37109 = ~n2727 & n37108;
  assign n37110 = n37070 & ~n37089;
  assign n37111 = ~pi72 & ~n37110;
  assign n37112 = ~n35647 & n37111;
  assign n37113 = ~n37109 & n37112;
  assign n37114 = n28319 & ~n37113;
  assign n37115 = ~n37107 & ~n37114;
  assign n37116 = ~n37108 & n37111;
  assign n37117 = n28319 & ~n37116;
  assign n37118 = n6416 & ~n37117;
  assign n37119 = ~n37115 & ~n37118;
  assign n37120 = ~n37100 & n37119;
  assign n37121 = ~pi39 & ~n37120;
  assign n37122 = n36291 & ~n37121;
  assign n37123 = pi100 & n2634;
  assign n37124 = n28567 & n31664;
  assign n37125 = pi137 & n37124;
  assign n37126 = pi129 & n58822;
  assign n37127 = ~pi137 & pi252;
  assign n37128 = pi683 & n32476;
  assign n37129 = pi252 & ~n37128;
  assign n37130 = pi252 & ~n2707;
  assign n37131 = ~n37128 & n37130;
  assign n37132 = ~n2707 & n37129;
  assign n37133 = ~n60087 & ~n60523;
  assign n37134 = ~n2682 & ~n37133;
  assign n37135 = ~n37127 & ~n37134;
  assign n37136 = ~n60087 & ~n32496;
  assign n37137 = ~n60087 & ~n37136;
  assign n37138 = ~n60087 & n32496;
  assign n37139 = ~n60523 & n60524;
  assign n37140 = ~n37135 & ~n37139;
  assign n37141 = n37126 & ~n37140;
  assign n37142 = ~n37125 & ~n37141;
  assign n37143 = n37123 & ~n37142;
  assign n37144 = ~pi90 & n29719;
  assign n37145 = ~pi93 & ~n37144;
  assign n37146 = ~n2528 & ~n37145;
  assign n37147 = ~pi35 & ~n37146;
  assign n37148 = pi35 & ~n31490;
  assign n37149 = n58820 & ~n37148;
  assign n37150 = ~n37147 & n37149;
  assign n37151 = ~pi32 & n37150;
  assign n37152 = n28770 & n60239;
  assign n37153 = pi32 & ~pi93;
  assign n37154 = n37152 & n37153;
  assign n37155 = n2554 & n37154;
  assign n37156 = ~n37151 & ~n37155;
  assign n37157 = ~pi95 & ~n60122;
  assign n37158 = ~n37156 & n37157;
  assign n37159 = ~n6380 & ~n37150;
  assign n37160 = pi1082 & n2598;
  assign n37161 = ~n37159 & n37160;
  assign n37162 = n60122 & ~n37147;
  assign n37163 = n2715 & n2793;
  assign n37164 = ~pi122 & n58838;
  assign n37165 = ~n3213 & n60525;
  assign n37166 = ~pi122 & ~po740;
  assign n37167 = n3213 & n37166;
  assign n37168 = ~n3213 & ~n60525;
  assign n37169 = n3213 & ~n37166;
  assign n37170 = ~n37168 & ~n37169;
  assign n37171 = ~n37165 & ~n37167;
  assign n37172 = ~n37162 & ~n60526;
  assign n37173 = pi76 & ~pi84;
  assign n37174 = n2457 & n37173;
  assign n37175 = n6323 & n35622;
  assign n37176 = ~pi73 & pi76;
  assign n37177 = n28346 & n37176;
  assign n37178 = n29132 & n35622;
  assign n37179 = n37177 & n37178;
  assign n37180 = n37174 & n37175;
  assign n37181 = n2446 & n2475;
  assign n37182 = n36225 & n37181;
  assign n37183 = n60527 & n37182;
  assign n37184 = ~pi103 & n2449;
  assign n37185 = n36226 & n37184;
  assign n37186 = ~pi45 & ~pi48;
  assign n37187 = ~pi61 & ~pi104;
  assign n37188 = n37186 & n37187;
  assign n37189 = n6325 & n37188;
  assign n37190 = n37185 & n37189;
  assign n37191 = n37183 & n37190;
  assign n37192 = n2503 & n37191;
  assign n37193 = n59134 & n37192;
  assign n37194 = n2579 & n37193;
  assign n37195 = n37147 & ~n37194;
  assign n37196 = ~pi137 & ~n60122;
  assign n37197 = n2598 & ~n37196;
  assign n37198 = n37149 & n37197;
  assign n37199 = ~n37195 & n37198;
  assign n37200 = ~n3213 & ~n37196;
  assign n37201 = n60525 & n37200;
  assign n37202 = n3213 & ~n37196;
  assign n37203 = n37166 & n37202;
  assign n37204 = ~n37201 & ~n37203;
  assign n37205 = n37147 & ~n60526;
  assign n37206 = n60122 & ~n37205;
  assign n37207 = pi137 & n60526;
  assign n37208 = ~n37206 & ~n37207;
  assign n37209 = ~n37162 & n37204;
  assign n37210 = n2598 & n37149;
  assign n37211 = ~n37195 & n37210;
  assign n37212 = ~n60528 & n37211;
  assign n37213 = ~n37172 & n37199;
  assign n37214 = ~pi38 & ~n60529;
  assign n37215 = ~pi38 & ~n37161;
  assign n37216 = ~n60529 & n37215;
  assign n37217 = ~n37161 & n37214;
  assign n37218 = ~n37158 & n60530;
  assign n37219 = pi38 & ~n58826;
  assign n37220 = ~pi39 & ~pi100;
  assign n37221 = ~n37219 & n37220;
  assign n37222 = ~n37218 & n37221;
  assign n37223 = ~n37143 & ~n37222;
  assign n37224 = n6309 & ~n37223;
  assign n37225 = pi75 & ~pi100;
  assign n37226 = n30890 & n37225;
  assign n37227 = ~pi24 & n37226;
  assign n37228 = pi252 & ~n32496;
  assign n37229 = pi137 & n35649;
  assign n37230 = ~n28570 & n37229;
  assign n37231 = ~n37228 & ~n37230;
  assign n37232 = n37227 & ~n37231;
  assign n37233 = n37226 & ~n37231;
  assign n37234 = n58826 & n37233;
  assign n37235 = n58822 & n37232;
  assign n37236 = ~n37224 & ~n60531;
  assign n37237 = n2438 & ~n37236;
  assign n37238 = ~pi24 & pi54;
  assign n37239 = n28585 & n37238;
  assign n37240 = ~n37237 & ~n37239;
  assign n37241 = ~pi92 & ~n37236;
  assign n37242 = ~pi54 & ~n37241;
  assign n37243 = ~pi24 & n28585;
  assign n37244 = pi54 & ~n37243;
  assign n37245 = n60411 & ~n37244;
  assign n37246 = ~n37242 & n37245;
  assign n37247 = n60411 & ~n37240;
  assign n37248 = ~pi59 & ~n60532;
  assign n37249 = n4437 & n28288;
  assign n37250 = n58826 & n37249;
  assign n37251 = ~pi55 & n37250;
  assign n37252 = pi59 & ~n37251;
  assign n37253 = ~pi57 & ~n37252;
  assign po193 = ~n37248 & n37253;
  assign n37255 = n58847 & n37051;
  assign n37256 = n58843 & n37053;
  assign n37257 = ~n37255 & ~n37256;
  assign po244 = n37049 & ~n37257;
  assign n37259 = ~pi979 & ~pi984;
  assign n37260 = pi1001 & n37259;
  assign n37261 = n6470 & n37260;
  assign n37262 = ~n2442 & n37261;
  assign n37263 = n2801 & n37262;
  assign n37264 = ~pi252 & ~n37263;
  assign n37265 = pi1092 & ~pi1093;
  assign n37266 = ~n37264 & n37265;
  assign n37267 = n28517 & ~n37266;
  assign n37268 = ~n2822 & ~n37267;
  assign n37269 = pi252 & pi1092;
  assign n37270 = ~pi1093 & n37269;
  assign n37271 = n2822 & n37270;
  assign n37272 = ~n37268 & ~n37271;
  assign n37273 = ~n2790 & ~n37272;
  assign n37274 = ~n2783 & n37270;
  assign n37275 = n2783 & ~n37267;
  assign n37276 = ~n37274 & ~n37275;
  assign n37277 = n2790 & ~n37276;
  assign n37278 = ~pi299 & ~n37277;
  assign n37279 = ~n37273 & n37278;
  assign n37280 = n58846 & ~n37276;
  assign n37281 = ~n58846 & ~n37272;
  assign n37282 = pi299 & ~n37281;
  assign n37283 = pi299 & ~n37280;
  assign n37284 = ~n37281 & n37283;
  assign n37285 = ~n37280 & n37282;
  assign n37286 = n37049 & ~n60533;
  assign n37287 = ~n37279 & n37286;
  assign n37288 = ~n37049 & n37270;
  assign n37289 = ~n5138 & ~n37288;
  assign n37290 = ~n37287 & n37289;
  assign n37291 = ~n28524 & ~n28532;
  assign n37292 = n25479 & n37261;
  assign n37293 = n25257 & n37292;
  assign n37294 = n60240 & n37293;
  assign n37295 = ~n37291 & n37294;
  assign n37296 = n2801 & n37295;
  assign n37297 = ~pi252 & ~n37296;
  assign n37298 = ~pi57 & pi1092;
  assign n37299 = ~n37297 & n37298;
  assign n37300 = pi57 & n37269;
  assign n37301 = n5138 & ~n37300;
  assign n37302 = ~n37299 & n37301;
  assign po409 = ~n37290 & ~n37302;
  assign n37304 = n2438 & n60412;
  assign n37305 = ~n3213 & n35649;
  assign n37306 = ~pi137 & ~n37305;
  assign n37307 = ~n29125 & ~n37191;
  assign n37308 = n58797 & ~n37307;
  assign n37309 = ~pi24 & ~n37308;
  assign n37310 = pi24 & ~n37193;
  assign n37311 = ~pi40 & n59138;
  assign n37312 = n2580 & n58820;
  assign n37313 = ~n37310 & n60534;
  assign n37314 = ~n37309 & n37313;
  assign n37315 = n37306 & ~n37314;
  assign n37316 = n2503 & n29125;
  assign n37317 = ~pi93 & n59134;
  assign n37318 = n37316 & n37317;
  assign n37319 = n37152 & n37318;
  assign n37320 = ~n37306 & ~n37319;
  assign n37321 = ~pi32 & ~n37320;
  assign n37322 = ~n37306 & n37319;
  assign n37323 = ~pi137 & n2580;
  assign n37324 = n58820 & n37323;
  assign n37325 = ~n37305 & n37324;
  assign n37326 = ~n37310 & n37325;
  assign n37327 = ~n37309 & n37326;
  assign n37328 = ~n37322 & ~n37327;
  assign n37329 = ~pi32 & ~n37328;
  assign n37330 = ~n37315 & n37321;
  assign n37331 = ~pi24 & ~pi841;
  assign n37332 = pi32 & ~n37331;
  assign n37333 = n31487 & n37332;
  assign n37334 = ~n60122 & ~n37333;
  assign n37335 = ~n60535 & n37334;
  assign n37336 = ~pi32 & ~n37319;
  assign n37337 = ~n31496 & ~n37336;
  assign n37338 = n60122 & ~n37337;
  assign n37339 = n28296 & ~n37338;
  assign n37340 = ~n60535 & ~n37333;
  assign n37341 = ~n60122 & ~n37340;
  assign n37342 = n60122 & ~n31496;
  assign n37343 = ~n37336 & n37342;
  assign n37344 = ~n37341 & ~n37343;
  assign n37345 = n28296 & ~n37344;
  assign n37346 = ~n37335 & n37339;
  assign n37347 = ~n60087 & n37228;
  assign n37348 = n37126 & n37347;
  assign n37349 = ~n37124 & ~n37348;
  assign n37350 = ~pi137 & n37123;
  assign n37351 = ~pi137 & n37124;
  assign n37352 = ~n60087 & n37127;
  assign n37353 = n37127 & n37136;
  assign n37354 = ~n32496 & n37352;
  assign n37355 = n37126 & n60537;
  assign n37356 = ~n37351 & ~n37355;
  assign n37357 = n37123 & ~n37356;
  assign n37358 = ~n37349 & n37350;
  assign n37359 = ~n60536 & ~n60538;
  assign n37360 = n6309 & ~n37359;
  assign n37361 = n58826 & n35649;
  assign n37362 = ~pi137 & n37226;
  assign n37363 = ~n28570 & n37362;
  assign n37364 = ~n37228 & n37363;
  assign n37365 = n37361 & n37364;
  assign n37366 = ~n37360 & ~n37365;
  assign po190 = n37304 & ~n37366;
  assign n37368 = pi39 & n36209;
  assign n37369 = n32632 & n37368;
  assign n37370 = n36209 & n37049;
  assign n37371 = ~n60475 & n60539;
  assign n37372 = ~n60474 & n60539;
  assign n37373 = ~n60475 & n37372;
  assign n37374 = ~n60474 & n37371;
  assign n37375 = ~n28301 & ~n28594;
  assign n37376 = pi93 & ~n2526;
  assign n37377 = ~n31479 & ~n37376;
  assign n37378 = pi58 & ~n58795;
  assign n37379 = ~n28325 & ~n37378;
  assign n37380 = n2445 & ~n2731;
  assign n37381 = ~pi91 & ~n31469;
  assign n37382 = ~n6360 & n37381;
  assign n37383 = n6361 & ~n31469;
  assign n37384 = ~pi81 & ~n31453;
  assign n37385 = n28400 & ~n37384;
  assign n37386 = n2470 & ~n37385;
  assign n37387 = n31459 & ~n37386;
  assign n37388 = n28339 & ~n37387;
  assign n37389 = n28337 & ~n37388;
  assign n37390 = n28335 & ~n37389;
  assign n37391 = ~n28333 & ~n37390;
  assign n37392 = ~pi86 & ~n37391;
  assign n37393 = n28411 & ~n37392;
  assign n37394 = n31413 & ~n37393;
  assign n37395 = ~n28628 & ~n37394;
  assign n37396 = ~pi108 & ~n37395;
  assign n37397 = n31410 & ~n37396;
  assign n37398 = n28449 & ~n37397;
  assign n37399 = ~n28447 & ~n37398;
  assign n37400 = n2540 & ~n37399;
  assign n37401 = n60541 & ~n37400;
  assign n37402 = n37380 & ~n37401;
  assign n37403 = n37379 & ~n37402;
  assign n37404 = n2592 & ~n37403;
  assign n37405 = n37377 & ~n37404;
  assign n37406 = ~pi70 & ~n37405;
  assign n37407 = ~n28320 & ~n37406;
  assign n37408 = ~pi51 & ~n37407;
  assign n37409 = n2604 & ~n37408;
  assign n37410 = n31408 & ~n37409;
  assign n37411 = n31402 & ~n37410;
  assign n37412 = ~pi1082 & n6380;
  assign n37413 = ~pi32 & ~n37412;
  assign n37414 = ~n37411 & n37413;
  assign n37415 = ~n31488 & ~n37414;
  assign n37416 = ~pi95 & ~n37415;
  assign n37417 = ~n31400 & ~n37416;
  assign n37418 = ~pi39 & ~n37417;
  assign n37419 = pi39 & ~n58822;
  assign n37420 = n2441 & n60240;
  assign n37421 = n2806 & n37420;
  assign n37422 = ~n37291 & n37421;
  assign n37423 = n6469 & n37368;
  assign n37424 = ~n37422 & n37423;
  assign n37425 = ~n37419 & ~n37424;
  assign n37426 = ~n37418 & n37425;
  assign n37427 = ~pi38 & ~n37426;
  assign n37428 = n31399 & ~n37427;
  assign n37429 = ~pi87 & ~n28549;
  assign n37430 = ~n37428 & n37429;
  assign n37431 = ~n31560 & ~n37430;
  assign n37432 = n6307 & ~n37431;
  assign n37433 = n28308 & ~n37432;
  assign n37434 = ~pi54 & ~n37433;
  assign n37435 = ~n28586 & ~n37434;
  assign n37436 = n31567 & ~n37435;
  assign n37437 = n37375 & ~n37436;
  assign n37438 = ~pi56 & ~n37437;
  assign n37439 = ~n31570 & ~n37438;
  assign n37440 = ~pi62 & ~n37439;
  assign n37441 = ~n31575 & ~n37440;
  assign n37442 = n4438 & ~n37441;
  assign po389 = n28295 & ~n37442;
  assign n37444 = pi41 & ~n36361;
  assign n37445 = n2793 & ~n36344;
  assign n37446 = ~n37444 & n37445;
  assign n37447 = pi41 & ~n36382;
  assign n37448 = ~n2793 & ~n37447;
  assign n37449 = ~n2793 & ~n36372;
  assign n37450 = ~n37447 & n37449;
  assign n37451 = ~n36372 & n37448;
  assign n37452 = pi228 & ~n60542;
  assign n37453 = ~n37446 & n37452;
  assign n37454 = pi41 & ~n36441;
  assign n37455 = ~n36427 & ~n37454;
  assign n37456 = ~pi228 & ~n37455;
  assign n37457 = ~pi39 & ~n37456;
  assign n37458 = ~n37453 & n37457;
  assign n37459 = pi144 & n30128;
  assign n37460 = ~pi174 & n37459;
  assign n37461 = ~pi299 & ~n37460;
  assign n37462 = pi161 & n29998;
  assign n37463 = ~pi152 & n37462;
  assign n37464 = ~n2675 & ~n37463;
  assign n37465 = pi232 & ~n37464;
  assign n37466 = pi232 & ~n37461;
  assign n37467 = ~n37464 & n37466;
  assign n37468 = ~n37461 & n37465;
  assign n37469 = ~pi72 & ~n60543;
  assign n37470 = n36455 & n60543;
  assign n37471 = ~n37469 & ~n37470;
  assign n37472 = pi39 & ~n37471;
  assign n37473 = n2636 & ~n37472;
  assign n37474 = ~n37458 & n37473;
  assign n37475 = pi39 & ~n37469;
  assign n37476 = ~pi41 & ~pi72;
  assign n37477 = ~n2719 & ~n37476;
  assign n37478 = ~n2793 & n37476;
  assign n37479 = n2719 & ~n37478;
  assign n37480 = ~pi99 & n58829;
  assign n37481 = ~pi41 & pi72;
  assign n37482 = n36327 & n36496;
  assign n37483 = ~n37481 & ~n37482;
  assign n37484 = ~n36494 & ~n37483;
  assign n37485 = ~n37480 & n37484;
  assign n37486 = n2715 & n36487;
  assign n37487 = pi41 & ~n37486;
  assign n37488 = n2793 & ~n37481;
  assign n37489 = n2793 & ~n37480;
  assign n37490 = ~n37488 & ~n37489;
  assign n37491 = ~n37487 & ~n37490;
  assign n37492 = ~n37485 & ~n37490;
  assign n37493 = ~n37487 & n37492;
  assign n37494 = ~n37485 & n37491;
  assign n37495 = n37479 & ~n60544;
  assign n37496 = ~n37477 & ~n37495;
  assign n37497 = ~pi39 & ~n37496;
  assign n37498 = ~n37475 & ~n37497;
  assign n37499 = n28548 & ~n37498;
  assign n37500 = ~pi39 & ~n37476;
  assign n37501 = ~n37475 & ~n37500;
  assign n37502 = pi38 & ~n37501;
  assign n37503 = ~pi87 & ~n37502;
  assign n37504 = ~n37499 & n37503;
  assign n37505 = ~n37474 & n37504;
  assign n37506 = pi41 & ~n36487;
  assign n37507 = pi228 & n37483;
  assign n37508 = pi228 & ~n37506;
  assign n37509 = n37483 & n37508;
  assign n37510 = ~n37506 & n37507;
  assign n37511 = ~pi228 & n37476;
  assign n37512 = n58815 & ~n37511;
  assign n37513 = ~n60545 & n37512;
  assign n37514 = ~n2636 & n37500;
  assign n37515 = pi87 & ~n37514;
  assign n37516 = ~n37475 & n37515;
  assign n37517 = ~n37513 & n37516;
  assign n37518 = ~pi75 & ~n37517;
  assign n37519 = ~n37505 & n37518;
  assign n37520 = n58827 & n37486;
  assign n37521 = pi41 & ~n37520;
  assign n37522 = n36327 & n36555;
  assign n37523 = ~n37480 & n37522;
  assign n37524 = n37488 & ~n37523;
  assign n37525 = n37488 & ~n37521;
  assign n37526 = ~n37523 & n37525;
  assign n37527 = ~n37521 & n37524;
  assign n37528 = n37479 & ~n60546;
  assign n37529 = ~n37477 & ~n37528;
  assign n37530 = ~pi39 & ~n37529;
  assign n37531 = n59291 & ~n37475;
  assign n37532 = ~n37530 & n37531;
  assign n37533 = ~n59291 & n37501;
  assign n37534 = pi75 & ~n37533;
  assign n37535 = ~n37532 & n37534;
  assign n37536 = ~n37519 & ~n37535;
  assign n37537 = n2439 & ~n37536;
  assign n37538 = ~n2439 & ~n37501;
  assign n37539 = n58992 & ~n37538;
  assign n37540 = ~n37537 & n37539;
  assign n37541 = n31239 & n37463;
  assign n37542 = ~pi72 & ~n37500;
  assign n37543 = ~n58992 & n37542;
  assign n37544 = ~n37541 & n37543;
  assign po199 = ~n37540 & ~n37544;
  assign n37546 = pi44 & ~pi72;
  assign n37547 = ~n2719 & ~n37546;
  assign n37548 = ~pi39 & ~n37547;
  assign n37549 = ~n2793 & n37546;
  assign n37550 = n2719 & ~n37549;
  assign n37551 = n2709 & ~n36328;
  assign n37552 = n2715 & n36486;
  assign n37553 = n58827 & n37552;
  assign n37554 = pi44 & ~n36554;
  assign n37555 = ~n37553 & ~n37554;
  assign n37556 = n37551 & ~n37555;
  assign n37557 = n37550 & ~n37556;
  assign n37558 = n37548 & ~n37557;
  assign n37559 = ~pi72 & n2682;
  assign n37560 = pi39 & n2682;
  assign n37561 = ~pi72 & n37560;
  assign n37562 = pi39 & n37559;
  assign n37563 = ~n37558 & ~n60547;
  assign n37564 = n59291 & ~n37563;
  assign n37565 = pi39 & ~n37559;
  assign n37566 = ~pi39 & ~n37546;
  assign n37567 = ~n37565 & ~n37566;
  assign n37568 = ~n59291 & n37567;
  assign n37569 = pi75 & ~n37568;
  assign n37570 = ~n37564 & n37569;
  assign n37571 = pi44 & n36368;
  assign n37572 = ~n2793 & ~n36381;
  assign n37573 = ~n37571 & n37572;
  assign n37574 = pi44 & n36340;
  assign n37575 = n2793 & ~n36360;
  assign n37576 = ~n37574 & n37575;
  assign n37577 = ~n37573 & ~n37576;
  assign n37578 = pi228 & ~n37577;
  assign n37579 = pi44 & n36423;
  assign n37580 = ~pi228 & ~n37579;
  assign n37581 = ~n36440 & n37580;
  assign n37582 = ~pi39 & ~n37581;
  assign n37583 = ~n37578 & n37582;
  assign n37584 = pi287 & n36495;
  assign n37585 = ~pi72 & ~n37584;
  assign n37586 = n37560 & n37585;
  assign n37587 = n60547 & ~n37584;
  assign n37588 = n2636 & ~n60548;
  assign n37589 = ~n37583 & n37588;
  assign n37590 = n2715 & n36495;
  assign n37591 = pi44 & ~n37590;
  assign n37592 = ~n37552 & ~n37591;
  assign n37593 = n37551 & ~n37592;
  assign n37594 = n37550 & ~n37593;
  assign n37595 = n37548 & ~n37594;
  assign n37596 = n28548 & ~n60547;
  assign n37597 = ~n37595 & n37596;
  assign n37598 = pi38 & ~n37567;
  assign n37599 = ~pi87 & ~n37598;
  assign n37600 = ~n37597 & n37599;
  assign n37601 = ~n37589 & n37600;
  assign n37602 = pi228 & n2636;
  assign n37603 = n36486 & n37602;
  assign n37604 = n36495 & n37602;
  assign n37605 = n37546 & ~n37604;
  assign n37606 = ~pi39 & ~n37605;
  assign n37607 = ~pi39 & ~n37603;
  assign n37608 = ~n37605 & n37607;
  assign n37609 = ~n37603 & n37606;
  assign n37610 = pi87 & ~n37565;
  assign n37611 = ~n60549 & n37610;
  assign n37612 = ~pi75 & ~n37611;
  assign n37613 = ~n37601 & n37612;
  assign n37614 = ~n37570 & ~n37613;
  assign n37615 = n2439 & ~n37614;
  assign n37616 = ~n2439 & ~n37567;
  assign n37617 = n58992 & ~n37616;
  assign n37618 = ~n37615 & n37617;
  assign n37619 = ~pi72 & n32475;
  assign n37620 = pi39 & ~n37619;
  assign n37621 = ~n58992 & ~n37566;
  assign n37622 = ~n37620 & n37621;
  assign n37623 = ~n37618 & ~n37622;
  assign n37624 = ~pi72 & pi99;
  assign n37625 = ~n2719 & ~n37624;
  assign n37626 = ~n2793 & n37624;
  assign n37627 = n2719 & ~n37626;
  assign n37628 = ~n37522 & n37624;
  assign n37629 = n2694 & n37553;
  assign n37630 = ~n37628 & ~n37629;
  assign n37631 = n37489 & ~n37630;
  assign n37632 = n37627 & ~n37631;
  assign n37633 = ~n37625 & ~n37632;
  assign n37634 = ~pi39 & ~n37633;
  assign n37635 = ~pi72 & pi152;
  assign n37636 = n37462 & n37635;
  assign n37637 = pi299 & n37636;
  assign n37638 = ~pi72 & pi174;
  assign n37639 = ~pi299 & n37638;
  assign n37640 = n37459 & n37639;
  assign n37641 = ~n37637 & ~n37640;
  assign n37642 = pi232 & ~n37641;
  assign n37643 = pi39 & ~n37642;
  assign n37644 = n59291 & ~n37643;
  assign n37645 = ~n37634 & n37644;
  assign n37646 = ~pi39 & ~n37624;
  assign n37647 = ~n37643 & ~n37646;
  assign n37648 = ~n59291 & n37647;
  assign n37649 = pi75 & ~n37648;
  assign n37650 = ~n37645 & n37649;
  assign n37651 = pi41 & pi72;
  assign n37652 = pi99 & ~n37651;
  assign n37653 = ~n36344 & n37652;
  assign n37654 = n36689 & ~n37653;
  assign n37655 = ~n36372 & n37652;
  assign n37656 = n36688 & ~n37655;
  assign n37657 = ~n37654 & ~n37656;
  assign n37658 = pi228 & ~n37657;
  assign n37659 = ~n36427 & n37652;
  assign n37660 = n36692 & ~n37659;
  assign n37661 = ~pi39 & ~n37660;
  assign n37662 = ~n37658 & n37661;
  assign n37663 = n31239 & ~n37641;
  assign n37664 = ~n37584 & n37663;
  assign n37665 = n2636 & ~n37664;
  assign n37666 = ~n37662 & n37665;
  assign n37667 = ~n37484 & n37624;
  assign n37668 = n2693 & n37486;
  assign n37669 = ~n37667 & ~n37668;
  assign n37670 = n37489 & ~n37669;
  assign n37671 = n37627 & ~n37670;
  assign n37672 = ~n37625 & ~n37671;
  assign n37673 = ~pi39 & ~n37672;
  assign n37674 = ~n37643 & ~n37673;
  assign n37675 = n28548 & ~n37674;
  assign n37676 = pi38 & ~n37647;
  assign n37677 = ~pi87 & ~n37676;
  assign n37678 = ~n37675 & n37677;
  assign n37679 = ~n37666 & n37678;
  assign n37680 = pi228 & n36488;
  assign n37681 = pi228 & n37482;
  assign n37682 = n37624 & ~n37681;
  assign n37683 = n58815 & ~n37682;
  assign n37684 = n58815 & ~n37680;
  assign n37685 = ~n37682 & n37684;
  assign n37686 = ~n37680 & n37683;
  assign n37687 = ~n58815 & ~n37647;
  assign n37688 = pi87 & ~n37687;
  assign n37689 = ~n60550 & n37688;
  assign n37690 = ~pi75 & ~n37689;
  assign n37691 = ~n37679 & n37690;
  assign n37692 = ~n37650 & ~n37691;
  assign n37693 = n2439 & ~n37692;
  assign n37694 = ~n2439 & ~n37647;
  assign n37695 = n58992 & ~n37694;
  assign n37696 = ~n37693 & n37695;
  assign n37697 = pi232 & n37636;
  assign n37698 = pi39 & ~n37697;
  assign n37699 = ~n58992 & ~n37646;
  assign n37700 = ~n37698 & n37699;
  assign n37701 = ~n37696 & ~n37700;
  assign n37702 = ~n2719 & ~n36326;
  assign n37703 = ~n2793 & n36326;
  assign n37704 = n2719 & ~n37703;
  assign n37705 = ~n2706 & n2793;
  assign n37706 = n36326 & ~n36555;
  assign n37707 = ~n37520 & ~n37706;
  assign n37708 = n37705 & ~n37707;
  assign n37709 = n37704 & ~n37708;
  assign n37710 = ~n37702 & ~n37709;
  assign n37711 = ~pi39 & ~n37710;
  assign n37712 = ~pi144 & pi174;
  assign n37713 = n30128 & n37712;
  assign n37714 = ~pi72 & n37713;
  assign n37715 = ~pi299 & ~n37714;
  assign n37716 = pi152 & ~pi161;
  assign n37717 = ~pi72 & n37716;
  assign n37718 = ~pi161 & ~pi166;
  assign n37719 = pi152 & n37718;
  assign n37720 = n2680 & n37719;
  assign n37721 = ~pi72 & n37720;
  assign n37722 = n29998 & n37717;
  assign n37723 = pi299 & ~n60551;
  assign n37724 = pi232 & ~n37723;
  assign n37725 = ~n37715 & n37724;
  assign n37726 = pi39 & ~n37725;
  assign n37727 = n59291 & ~n37726;
  assign n37728 = ~n37711 & n37727;
  assign n37729 = ~pi39 & ~n36326;
  assign n37730 = ~n37726 & ~n37729;
  assign n37731 = ~n59291 & n37730;
  assign n37732 = pi75 & ~n37731;
  assign n37733 = ~n37728 & n37732;
  assign n37734 = pi101 & n36370;
  assign n37735 = ~n2793 & ~n36382;
  assign n37736 = ~n37734 & n37735;
  assign n37737 = pi101 & n36342;
  assign n37738 = n2793 & ~n36361;
  assign n37739 = ~n37737 & n37738;
  assign n37740 = ~n37736 & ~n37739;
  assign n37741 = pi228 & ~n37740;
  assign n37742 = pi101 & n36425;
  assign n37743 = ~pi228 & ~n36441;
  assign n37744 = ~n37742 & n37743;
  assign n37745 = ~pi39 & ~n37744;
  assign n37746 = ~n37741 & n37745;
  assign n37747 = ~pi299 & n37713;
  assign n37748 = pi299 & n37716;
  assign n37749 = n29998 & n37748;
  assign n37750 = ~n37747 & ~n37749;
  assign n37751 = ~pi72 & n31239;
  assign n37752 = ~n37750 & n37751;
  assign n37753 = n37585 & n37713;
  assign n37754 = ~pi299 & ~n37753;
  assign n37755 = n37585 & n37720;
  assign n37756 = pi299 & ~n37755;
  assign n37757 = n31239 & ~n37756;
  assign n37758 = ~n37754 & n37757;
  assign n37759 = ~n37584 & n37752;
  assign n37760 = n2636 & ~n60552;
  assign n37761 = ~n37746 & n37760;
  assign n37762 = n2715 & n36496;
  assign n37763 = ~pi44 & n37590;
  assign n37764 = n36326 & ~n60553;
  assign n37765 = ~n37486 & ~n37764;
  assign n37766 = n37705 & ~n37765;
  assign n37767 = n37704 & ~n37766;
  assign n37768 = ~n37702 & ~n37767;
  assign n37769 = ~pi39 & ~n37768;
  assign n37770 = ~n37726 & ~n37769;
  assign n37771 = n28548 & ~n37770;
  assign n37772 = pi38 & ~n37730;
  assign n37773 = ~pi87 & ~n37772;
  assign n37774 = ~n37771 & n37773;
  assign n37775 = ~n37761 & n37774;
  assign n37776 = ~pi101 & n37603;
  assign n37777 = n36496 & n37602;
  assign n37778 = n36326 & ~n37777;
  assign n37779 = ~pi39 & ~n37778;
  assign n37780 = ~pi39 & ~n37776;
  assign n37781 = ~n37778 & n37780;
  assign n37782 = ~n37776 & n37779;
  assign n37783 = pi87 & ~n37726;
  assign n37784 = ~n60554 & n37783;
  assign n37785 = ~pi75 & ~n37784;
  assign n37786 = ~n37775 & n37785;
  assign n37787 = ~n37733 & ~n37786;
  assign n37788 = n2439 & ~n37787;
  assign n37789 = ~n2439 & ~n37730;
  assign n37790 = n58992 & ~n37789;
  assign n37791 = ~n37788 & n37790;
  assign n37792 = pi232 & n60551;
  assign n37793 = pi39 & ~n37792;
  assign n37794 = ~n58992 & ~n37729;
  assign n37795 = ~n37793 & n37794;
  assign n37796 = ~n37791 & ~n37795;
  assign n37797 = pi252 & n2757;
  assign n37798 = n58798 & n60165;
  assign n37799 = n2599 & n36406;
  assign n37800 = n31412 & n37798;
  assign n37801 = ~n37797 & n60555;
  assign n37802 = ~pi137 & n37801;
  assign n37803 = ~pi137 & n2793;
  assign n37804 = pi94 & ~n31412;
  assign n37805 = ~pi94 & ~n37192;
  assign n37806 = n37798 & ~n37805;
  assign n37807 = ~n59134 & ~n36404;
  assign n37808 = n60165 & ~n37805;
  assign n37809 = ~n37807 & n37808;
  assign n37810 = ~n37804 & n37806;
  assign n37811 = ~n2757 & ~n60556;
  assign n37812 = ~pi252 & n60556;
  assign n37813 = n58819 & n29201;
  assign n37814 = n2621 & n29201;
  assign n37815 = n58792 & n37814;
  assign n37816 = n58817 & n37815;
  assign n37817 = n2621 & n6403;
  assign n37818 = n58792 & n37813;
  assign n37819 = n37191 & n60557;
  assign n37820 = pi252 & n37819;
  assign n37821 = n2757 & ~n37820;
  assign n37822 = ~n37812 & n37821;
  assign n37823 = ~n37811 & ~n37822;
  assign n37824 = pi122 & ~n37823;
  assign n37825 = n2727 & n37811;
  assign n37826 = ~n2443 & ~n60555;
  assign n37827 = ~n37822 & ~n37826;
  assign n37828 = ~n37825 & n37827;
  assign n37829 = ~pi122 & ~n37828;
  assign n37830 = ~n37824 & ~n37829;
  assign n37831 = ~pi1093 & ~n37830;
  assign n37832 = ~pi122 & ~n37801;
  assign n37833 = ~n37824 & ~n37832;
  assign n37834 = pi1093 & ~n37833;
  assign n37835 = ~n37831 & ~n37834;
  assign n37836 = n2793 & ~n37835;
  assign n37837 = ~n37803 & ~n37836;
  assign n37838 = ~n37802 & ~n37837;
  assign n37839 = ~pi122 & n60555;
  assign n37840 = pi1093 & ~n60556;
  assign n37841 = ~n3865 & ~n37840;
  assign n37842 = ~n37839 & ~n37841;
  assign n37843 = ~n37831 & ~n37842;
  assign n37844 = ~n2793 & ~n37843;
  assign n37845 = ~pi137 & ~n2793;
  assign n37846 = ~n37844 & ~n37845;
  assign n37847 = n2795 & n37270;
  assign n37848 = ~pi137 & ~n37847;
  assign n37849 = n60555 & n37848;
  assign n37850 = ~n37846 & ~n37849;
  assign n37851 = ~n37838 & ~n37850;
  assign n37852 = n2707 & ~n37851;
  assign n37853 = ~n37166 & n37819;
  assign n37854 = ~n2707 & ~n37853;
  assign n37855 = ~pi137 & ~n2707;
  assign n37856 = ~n37854 & ~n37855;
  assign n37857 = ~n37852 & n37856;
  assign n37858 = ~pi210 & ~n37857;
  assign n37859 = ~n37836 & ~n37844;
  assign n37860 = n2707 & ~n37859;
  assign n37861 = ~n37854 & ~n37860;
  assign n37862 = pi210 & ~n37861;
  assign n37863 = ~n37858 & ~n37862;
  assign n37864 = n2676 & n29998;
  assign n37865 = ~n37863 & ~n37864;
  assign n37866 = ~pi210 & n37851;
  assign n37867 = pi210 & n37859;
  assign n37868 = n37864 & ~n37867;
  assign n37869 = pi210 & ~n37859;
  assign n37870 = ~pi210 & ~n37851;
  assign n37871 = ~n37869 & ~n37870;
  assign n37872 = n37864 & ~n37871;
  assign n37873 = ~n37866 & n37868;
  assign n37874 = pi299 & ~n60558;
  assign n37875 = ~n37865 & n37874;
  assign n37876 = ~pi198 & ~n37857;
  assign n37877 = pi198 & ~n37861;
  assign n37878 = ~n37876 & ~n37877;
  assign n37879 = n2674 & n2680;
  assign n37880 = ~n37878 & ~n37879;
  assign n37881 = ~pi198 & n37851;
  assign n37882 = pi198 & n37859;
  assign n37883 = n37879 & ~n37882;
  assign n37884 = pi198 & ~n37859;
  assign n37885 = ~pi198 & ~n37851;
  assign n37886 = ~n37884 & ~n37885;
  assign n37887 = n37879 & ~n37886;
  assign n37888 = ~n37881 & n37883;
  assign n37889 = ~pi299 & ~n60559;
  assign n37890 = ~n37880 & n37889;
  assign n37891 = ~n37875 & ~n37890;
  assign n37892 = pi232 & ~n37891;
  assign n37893 = pi299 & ~n37863;
  assign n37894 = ~pi299 & ~n37878;
  assign n37895 = ~pi232 & ~n37894;
  assign n37896 = ~pi232 & ~n37893;
  assign n37897 = ~n37894 & n37896;
  assign n37898 = ~n37893 & n37895;
  assign n37899 = n3213 & ~n60560;
  assign n37900 = ~n37892 & n37899;
  assign n37901 = n31593 & n60412;
  assign n37902 = n6307 & n32859;
  assign n37903 = n58992 & n6308;
  assign n37904 = n2672 & n60561;
  assign n37905 = n60069 & n32859;
  assign n37906 = ~pi92 & n37905;
  assign n37907 = n58992 & n31592;
  assign n37908 = ~pi74 & n37907;
  assign n37909 = n60203 & n32859;
  assign n37910 = n58992 & n28288;
  assign n37911 = n2757 & ~n60555;
  assign n37912 = ~n37797 & ~n37911;
  assign n37913 = ~n37797 & ~n37811;
  assign n37914 = ~n37911 & n37913;
  assign n37915 = ~n37811 & n37912;
  assign n37916 = n3865 & ~n60564;
  assign n37917 = ~n37824 & ~n37916;
  assign n37918 = n2793 & ~n37917;
  assign n37919 = ~n2793 & n37840;
  assign n37920 = ~pi1093 & ~n37823;
  assign n37921 = ~n37919 & ~n37920;
  assign n37922 = ~n37918 & n37921;
  assign n37923 = n2707 & n37922;
  assign n37924 = ~n2707 & n37819;
  assign n37925 = ~n60525 & n37924;
  assign n37926 = ~n37923 & ~n37925;
  assign n37927 = pi210 & ~n37926;
  assign n37928 = pi137 & n37920;
  assign n37929 = ~pi137 & ~n60564;
  assign n37930 = ~pi1093 & n37929;
  assign n37931 = ~n37840 & ~n37930;
  assign n37932 = ~n37840 & ~n37928;
  assign n37933 = ~n37930 & n37932;
  assign n37934 = ~n37928 & n37931;
  assign n37935 = n2707 & n60565;
  assign n37936 = ~n37924 & ~n37935;
  assign n37937 = n35648 & n37855;
  assign n37938 = ~n2793 & ~n37937;
  assign n37939 = ~n37936 & n37938;
  assign n37940 = pi137 & ~n37917;
  assign n37941 = ~n37928 & ~n37929;
  assign n37942 = ~n37940 & n37941;
  assign n37943 = n2707 & ~n37942;
  assign n37944 = pi137 & ~n3865;
  assign n37945 = n2757 & ~n37944;
  assign n37946 = n37819 & ~n37945;
  assign n37947 = ~n2707 & ~n37946;
  assign n37948 = n2793 & ~n37947;
  assign n37949 = ~n37943 & n37948;
  assign n37950 = ~n37939 & ~n37949;
  assign n37951 = ~pi210 & ~n37950;
  assign n37952 = ~n37927 & ~n37951;
  assign n37953 = ~n37864 & ~n37952;
  assign n37954 = ~n2793 & n60565;
  assign n37955 = n2793 & n37942;
  assign n37956 = ~n37954 & ~n37955;
  assign n37957 = ~pi210 & n37956;
  assign n37958 = pi210 & ~n37922;
  assign n37959 = n37864 & ~n37958;
  assign n37960 = ~pi210 & ~n37956;
  assign n37961 = pi210 & n37922;
  assign n37962 = ~n37960 & ~n37961;
  assign n37963 = n37864 & ~n37962;
  assign n37964 = ~n37957 & n37959;
  assign n37965 = pi299 & ~n60566;
  assign n37966 = ~n37953 & n37965;
  assign n37967 = pi198 & ~n37926;
  assign n37968 = ~pi198 & ~n37950;
  assign n37969 = ~n37967 & ~n37968;
  assign n37970 = ~n37879 & ~n37969;
  assign n37971 = ~pi198 & n37956;
  assign n37972 = pi198 & ~n37922;
  assign n37973 = n37879 & ~n37972;
  assign n37974 = ~pi198 & ~n37956;
  assign n37975 = pi198 & n37922;
  assign n37976 = ~n37974 & ~n37975;
  assign n37977 = n37879 & ~n37976;
  assign n37978 = ~n37971 & n37973;
  assign n37979 = ~pi299 & ~n60567;
  assign n37980 = ~n37970 & n37979;
  assign n37981 = ~n37966 & ~n37980;
  assign n37982 = pi232 & ~n37981;
  assign n37983 = pi299 & ~n37952;
  assign n37984 = ~pi299 & ~n37969;
  assign n37985 = ~pi232 & ~n37984;
  assign n37986 = ~n37983 & n37985;
  assign n37987 = ~n37982 & ~n37986;
  assign n37988 = ~n3213 & ~n37987;
  assign n37989 = n60562 & ~n37988;
  assign n37990 = ~n37892 & ~n60560;
  assign n37991 = n3213 & ~n37990;
  assign n37992 = ~n3213 & ~n37986;
  assign n37993 = ~n37982 & n37992;
  assign n37994 = ~n37991 & ~n37993;
  assign n37995 = n60562 & ~n37994;
  assign n37996 = ~n37900 & n37989;
  assign n37997 = ~pi99 & ~n37449;
  assign n37998 = ~n37445 & n37997;
  assign n37999 = pi113 & ~n36325;
  assign n38000 = ~n37998 & n37999;
  assign n38001 = ~pi113 & n36690;
  assign n38002 = pi228 & ~n38001;
  assign n38003 = ~n38000 & n38002;
  assign n38004 = pi113 & n36429;
  assign n38005 = ~pi228 & ~n36443;
  assign n38006 = ~n38004 & n38005;
  assign n38007 = ~pi39 & ~n38006;
  assign n38008 = ~n38003 & n38007;
  assign n38009 = n2636 & ~n38008;
  assign n38010 = ~pi72 & pi113;
  assign n38011 = ~pi39 & n38010;
  assign n38012 = pi38 & ~n38011;
  assign n38013 = n2719 & n2793;
  assign n38014 = n2715 & n36497;
  assign n38015 = ~n58829 & ~n38014;
  assign n38016 = n38013 & ~n38015;
  assign n38017 = n38010 & ~n38016;
  assign n38018 = ~n58829 & n38013;
  assign n38019 = ~pi113 & n38018;
  assign n38020 = n37668 & n38019;
  assign n38021 = ~n38017 & ~n38020;
  assign n38022 = ~pi39 & ~n38021;
  assign n38023 = n28548 & ~n38022;
  assign n38024 = ~n38012 & ~n38023;
  assign n38025 = ~n38009 & n38024;
  assign n38026 = ~pi87 & ~n38025;
  assign n38027 = ~n36533 & n38010;
  assign n38028 = ~pi113 & n37680;
  assign n38029 = ~n38027 & ~n38028;
  assign n38030 = n58815 & ~n38029;
  assign n38031 = ~n2636 & n38011;
  assign n38032 = pi87 & ~n38031;
  assign n38033 = ~n38030 & n38032;
  assign n38034 = ~n38026 & ~n38033;
  assign n38035 = ~pi75 & ~n38034;
  assign n38036 = n58827 & n38020;
  assign n38037 = ~n58829 & ~n36556;
  assign n38038 = n38013 & ~n38037;
  assign n38039 = n38010 & ~n38038;
  assign n38040 = ~n38036 & ~n38039;
  assign n38041 = n2672 & ~n38040;
  assign n38042 = ~n59291 & n38011;
  assign n38043 = pi75 & ~n38042;
  assign n38044 = ~n38041 & n38043;
  assign n38045 = ~n38035 & ~n38044;
  assign n38046 = n37304 & ~n38045;
  assign n38047 = ~n37304 & ~n38011;
  assign po271 = ~n38046 & ~n38047;
  assign n38049 = ~pi72 & pi114;
  assign n38050 = pi114 & n36773;
  assign n38051 = ~n36558 & n38049;
  assign n38052 = n36925 & ~n60569;
  assign n38053 = ~n36549 & n36925;
  assign n38054 = ~n60569 & n38053;
  assign n38055 = ~n36549 & n38052;
  assign n38056 = ~n36925 & ~n38049;
  assign n38057 = n2672 & ~n38056;
  assign n38058 = ~n60570 & n38057;
  assign n38059 = ~pi39 & n38049;
  assign n38060 = ~n59291 & n38059;
  assign n38061 = pi75 & ~n38060;
  assign n38062 = ~n38058 & n38061;
  assign n38063 = pi114 & n36714;
  assign n38064 = ~pi114 & n60507;
  assign n38065 = ~pi115 & ~n38064;
  assign n38066 = pi114 & ~n36714;
  assign n38067 = ~pi114 & ~n60507;
  assign n38068 = ~n38066 & ~n38067;
  assign n38069 = ~pi115 & ~n38068;
  assign n38070 = ~n38063 & n38065;
  assign n38071 = pi115 & ~n38049;
  assign n38072 = ~pi39 & ~n38071;
  assign n38073 = ~n60571 & n38072;
  assign n38074 = n2636 & ~n38073;
  assign n38075 = pi114 & ~n36500;
  assign n38076 = n36925 & ~n38075;
  assign n38077 = ~n36492 & n36925;
  assign n38078 = ~n38075 & n38077;
  assign n38079 = ~n36492 & n38076;
  assign n38080 = ~pi39 & ~n38056;
  assign n38081 = ~n60572 & n38080;
  assign n38082 = n28548 & ~n38081;
  assign n38083 = pi38 & ~n38059;
  assign n38084 = ~pi87 & ~n38083;
  assign n38085 = ~n38082 & n38084;
  assign n38086 = ~n38074 & n38085;
  assign n38087 = ~n36535 & n38049;
  assign n38088 = n2636 & ~n38087;
  assign n38089 = n2636 & ~n60493;
  assign n38090 = ~n38087 & n38089;
  assign n38091 = ~n60493 & n38088;
  assign n38092 = ~n2636 & ~n38059;
  assign n38093 = n36896 & ~n38092;
  assign n38094 = ~n60573 & n38093;
  assign n38095 = ~pi75 & ~n38094;
  assign n38096 = ~n38086 & n38095;
  assign n38097 = ~n38062 & ~n38096;
  assign n38098 = n37304 & ~n38097;
  assign n38099 = ~n37304 & ~n38059;
  assign po272 = ~n38098 & ~n38099;
  assign n38101 = ~pi52 & n2699;
  assign n38102 = ~pi115 & ~n38101;
  assign n38103 = n36490 & n38102;
  assign n38104 = n58827 & n38103;
  assign n38105 = pi115 & n36773;
  assign n38106 = n38013 & ~n38105;
  assign n38107 = n38013 & ~n38104;
  assign n38108 = ~n38105 & n38107;
  assign n38109 = ~n38104 & n38106;
  assign n38110 = ~pi72 & pi115;
  assign n38111 = ~n38013 & ~n38110;
  assign n38112 = n2672 & ~n38111;
  assign n38113 = ~n60574 & n38112;
  assign n38114 = ~pi39 & n38110;
  assign n38115 = ~n59291 & n38114;
  assign n38116 = pi75 & ~n38115;
  assign n38117 = ~n38113 & n38116;
  assign n38118 = pi115 & ~n36714;
  assign n38119 = ~pi115 & ~n60507;
  assign n38120 = ~pi39 & ~n38119;
  assign n38121 = ~n38118 & n38120;
  assign n38122 = n2636 & ~n38121;
  assign n38123 = pi115 & ~n36500;
  assign n38124 = n38013 & ~n38123;
  assign n38125 = n38013 & ~n38103;
  assign n38126 = ~n38123 & n38125;
  assign n38127 = ~n38103 & n38124;
  assign n38128 = ~pi39 & ~n38111;
  assign n38129 = ~n60575 & n38128;
  assign n38130 = n28548 & ~n38129;
  assign n38131 = pi38 & ~n38114;
  assign n38132 = ~pi87 & ~n38131;
  assign n38133 = ~n38130 & n38132;
  assign n38134 = ~n38122 & n38133;
  assign n38135 = ~n36534 & n38110;
  assign n38136 = n2636 & ~n38135;
  assign n38137 = n2636 & ~n36528;
  assign n38138 = ~n38135 & n38137;
  assign n38139 = ~n36528 & n38136;
  assign n38140 = ~n2636 & ~n38114;
  assign n38141 = n36896 & ~n38140;
  assign n38142 = ~n60576 & n38141;
  assign n38143 = ~pi75 & ~n38142;
  assign n38144 = ~n38134 & n38143;
  assign n38145 = ~n38117 & ~n38144;
  assign n38146 = n37304 & ~n38145;
  assign n38147 = ~n37304 & ~n38114;
  assign po273 = ~n38146 & ~n38147;
  assign n38149 = ~pi72 & pi116;
  assign n38150 = ~n38013 & n38149;
  assign n38151 = ~n36557 & n38149;
  assign n38152 = ~n36775 & ~n38151;
  assign n38153 = n38018 & ~n38152;
  assign n38154 = ~n38150 & ~n38153;
  assign n38155 = n2672 & ~n38154;
  assign n38156 = ~pi39 & n38149;
  assign n38157 = ~n59291 & n38156;
  assign n38158 = pi75 & ~n38157;
  assign n38159 = ~n38155 & n38158;
  assign n38160 = n2793 & ~n36348;
  assign n38161 = ~n2793 & ~n36376;
  assign n38162 = pi116 & ~n38161;
  assign n38163 = ~n38160 & n38162;
  assign n38164 = pi116 & n36376;
  assign n38165 = ~n2793 & ~n38164;
  assign n38166 = pi116 & ~n38160;
  assign n38167 = ~n36363 & ~n38166;
  assign n38168 = ~n38165 & ~n38167;
  assign n38169 = n36696 & ~n38168;
  assign n38170 = n60506 & ~n38163;
  assign n38171 = pi116 & n36431;
  assign n38172 = n36700 & ~n38171;
  assign n38173 = ~pi39 & ~n38172;
  assign n38174 = ~n60577 & n38173;
  assign n38175 = n2636 & ~n38174;
  assign n38176 = ~pi113 & n38014;
  assign n38177 = n38149 & ~n38176;
  assign n38178 = ~n36490 & ~n38177;
  assign n38179 = n38018 & ~n38178;
  assign n38180 = ~n38150 & ~n38179;
  assign n38181 = ~pi39 & ~n38180;
  assign n38182 = n28548 & ~n38181;
  assign n38183 = pi38 & ~n38156;
  assign n38184 = ~pi87 & ~n38183;
  assign n38185 = ~n38182 & n38184;
  assign n38186 = ~n38175 & n38185;
  assign n38187 = ~pi38 & ~pi113;
  assign n38188 = n36533 & n38187;
  assign n38189 = n38149 & ~n38188;
  assign n38190 = ~n36527 & ~n38189;
  assign n38191 = ~pi113 & n36533;
  assign n38192 = n38149 & ~n38191;
  assign n38193 = ~pi38 & ~n38192;
  assign n38194 = ~n36527 & n38193;
  assign n38195 = ~n38183 & ~n38194;
  assign n38196 = ~n38183 & ~n38190;
  assign n38197 = ~pi100 & ~n60578;
  assign n38198 = pi100 & ~n38156;
  assign n38199 = n36896 & ~n38198;
  assign n38200 = ~n38197 & n38199;
  assign n38201 = ~pi75 & ~n38200;
  assign n38202 = ~n38186 & n38201;
  assign n38203 = ~n38159 & ~n38202;
  assign n38204 = n37304 & ~n38203;
  assign n38205 = ~n37304 & ~n38156;
  assign po274 = ~n38204 & ~n38205;
  assign n38207 = ~pi332 & ~pi1144;
  assign n38208 = pi215 & ~n38207;
  assign n38209 = pi265 & ~pi332;
  assign n38210 = pi216 & ~n38209;
  assign n38211 = pi105 & pi228;
  assign n38212 = pi234 & n28313;
  assign n38213 = ~pi332 & ~n38212;
  assign n38214 = n38211 & n38213;
  assign n38215 = pi153 & ~pi332;
  assign n38216 = ~n38211 & n38215;
  assign n38217 = ~pi216 & ~n38216;
  assign n38218 = ~n38214 & n38217;
  assign n38219 = ~n38210 & ~n38218;
  assign n38220 = ~pi221 & ~n38219;
  assign n38221 = ~pi216 & pi833;
  assign n38222 = pi929 & n38221;
  assign n38223 = pi1144 & ~n38221;
  assign n38224 = ~pi332 & ~n38223;
  assign n38225 = ~n38222 & n38224;
  assign n38226 = pi221 & ~n38225;
  assign n38227 = ~n38220 & ~n38226;
  assign n38228 = ~pi215 & ~n38227;
  assign n38229 = ~n38208 & ~n38228;
  assign n38230 = pi137 & n58822;
  assign n38231 = ~n58822 & ~n28313;
  assign n38232 = pi234 & ~n38231;
  assign n38233 = ~pi234 & n58822;
  assign n38234 = ~n38232 & ~n38233;
  assign n38235 = ~n58822 & ~n38212;
  assign n38236 = pi137 & ~n60579;
  assign n38237 = n38213 & ~n38236;
  assign n38238 = n38213 & ~n38230;
  assign n38239 = ~pi215 & ~pi221;
  assign n38240 = n38217 & n38239;
  assign n38241 = ~n60580 & n38240;
  assign n38242 = n28292 & n38241;
  assign n38243 = ~pi59 & n38242;
  assign n38244 = n38229 & ~n38243;
  assign n38245 = pi57 & ~n38244;
  assign n38246 = ~pi105 & ~n38215;
  assign n38247 = pi479 & n31400;
  assign n38248 = n2642 & n31491;
  assign n38249 = ~pi40 & n2642;
  assign n38250 = ~pi51 & n2597;
  assign n38251 = n2593 & n60581;
  assign n38252 = n58807 & n38248;
  assign n38253 = n31407 & n60582;
  assign n38254 = n2604 & ~n35572;
  assign n38255 = pi35 & n58807;
  assign n38256 = ~pi225 & n38255;
  assign n38257 = ~n31479 & ~n38256;
  assign n38258 = ~pi35 & ~n32868;
  assign n38259 = n28339 & ~n31460;
  assign n38260 = n28337 & ~n38259;
  assign n38261 = n28335 & ~n38260;
  assign n38262 = ~n28333 & ~n38261;
  assign n38263 = ~pi86 & ~n38262;
  assign n38264 = n28411 & ~n38263;
  assign n38265 = n31413 & ~n38264;
  assign n38266 = ~n28628 & ~n38265;
  assign n38267 = ~pi108 & ~n38266;
  assign n38268 = n31410 & ~n38267;
  assign n38269 = n28449 & ~n38268;
  assign n38270 = ~n28447 & ~n38269;
  assign n38271 = n2540 & ~n38270;
  assign n38272 = n60541 & ~n38271;
  assign n38273 = n37380 & ~n38272;
  assign n38274 = n32527 & ~n37378;
  assign n38275 = ~n38273 & n38274;
  assign n38276 = n38258 & ~n38275;
  assign n38277 = n38257 & ~n38276;
  assign n38278 = ~pi51 & ~n38277;
  assign n38279 = n38254 & ~n38278;
  assign n38280 = ~pi72 & ~n38279;
  assign n38281 = n31402 & ~n38280;
  assign n38282 = n31401 & ~n38281;
  assign n38283 = ~n38253 & n38282;
  assign n38284 = n2642 & n31490;
  assign n38285 = pi225 & n2641;
  assign n38286 = pi225 & n31491;
  assign n38287 = n2641 & n38286;
  assign n38288 = n31491 & n38285;
  assign n38289 = n38284 & n60583;
  assign n38290 = pi32 & ~n38289;
  assign n38291 = ~n38283 & ~n38290;
  assign n38292 = ~pi95 & ~n38291;
  assign n38293 = ~n38247 & ~n38292;
  assign n38294 = pi137 & ~n38293;
  assign n38295 = pi95 & pi479;
  assign n38296 = ~n28335 & n29725;
  assign n38297 = n58798 & n2579;
  assign n38298 = n38296 & n38297;
  assign n38299 = ~pi35 & ~n38298;
  assign n38300 = ~pi70 & ~n38256;
  assign n38301 = ~pi51 & n38300;
  assign n38302 = ~n31479 & n38301;
  assign n38303 = ~n38299 & n38302;
  assign n38304 = ~pi96 & ~n38303;
  assign n38305 = n36312 & ~n38304;
  assign n38306 = ~pi32 & ~n38305;
  assign n38307 = ~n38290 & ~n38306;
  assign n38308 = ~pi95 & ~n38307;
  assign n38309 = ~n38295 & ~n38308;
  assign n38310 = ~pi137 & ~n38309;
  assign n38311 = ~n38294 & ~n38310;
  assign n38312 = ~pi210 & ~n38311;
  assign n38313 = pi225 & n31487;
  assign n38314 = pi32 & ~n38313;
  assign n38315 = ~pi95 & ~n38314;
  assign n38316 = ~n38306 & n38315;
  assign n38317 = ~n28313 & ~n38316;
  assign n38318 = ~pi137 & n38317;
  assign n38319 = ~n38283 & ~n38314;
  assign n38320 = ~pi95 & ~n38319;
  assign n38321 = ~n38247 & ~n38320;
  assign n38322 = pi137 & ~n38321;
  assign n38323 = ~n38318 & ~n38322;
  assign n38324 = pi210 & ~n38323;
  assign n38325 = ~pi146 & ~n38324;
  assign n38326 = ~n38312 & n38325;
  assign n38327 = pi234 & ~pi332;
  assign n38328 = ~pi97 & ~n38296;
  assign n38329 = n2589 & n28632;
  assign n38330 = ~n38328 & n38329;
  assign n38331 = n28630 & n38329;
  assign n38332 = ~n38328 & n38331;
  assign n38333 = n28630 & n38330;
  assign n38334 = ~pi35 & ~n60584;
  assign n38335 = n38302 & ~n38334;
  assign n38336 = ~pi96 & ~n38335;
  assign n38337 = n36312 & ~n38336;
  assign n38338 = ~pi32 & ~n38337;
  assign n38339 = ~n38290 & ~n38338;
  assign n38340 = ~pi95 & ~n38339;
  assign n38341 = ~n38295 & ~n38340;
  assign n38342 = n58838 & n38341;
  assign n38343 = ~n58838 & n38309;
  assign n38344 = ~pi137 & ~n38343;
  assign n38345 = ~n38342 & n38344;
  assign n38346 = ~n2793 & n38311;
  assign n38347 = n2796 & ~n38295;
  assign n38348 = ~n38340 & n38347;
  assign n38349 = ~n2796 & n38309;
  assign n38350 = ~pi137 & ~n38349;
  assign n38351 = ~pi137 & ~n38348;
  assign n38352 = ~n38349 & n38351;
  assign n38353 = ~n38348 & n38350;
  assign n38354 = n2793 & ~n60585;
  assign n38355 = ~n38294 & n38354;
  assign n38356 = ~n38346 & ~n38355;
  assign n38357 = ~n38294 & ~n38345;
  assign n38358 = ~pi210 & n60586;
  assign n38359 = ~n38324 & ~n38358;
  assign n38360 = pi146 & n38359;
  assign n38361 = n38327 & ~n38360;
  assign n38362 = ~n38326 & n38327;
  assign n38363 = ~n38360 & n38362;
  assign n38364 = ~n38326 & n38361;
  assign n38365 = ~n28313 & ~n31400;
  assign n38366 = ~n38282 & ~n38290;
  assign n38367 = ~pi95 & ~n38366;
  assign n38368 = n38365 & ~n38367;
  assign n38369 = pi137 & ~n38368;
  assign n38370 = n2601 & n38303;
  assign n38371 = ~pi32 & ~n38370;
  assign n38372 = ~pi95 & ~n38290;
  assign n38373 = ~n38371 & n38372;
  assign n38374 = ~pi137 & ~n38373;
  assign n38375 = ~n38369 & ~n38374;
  assign n38376 = ~pi210 & ~n38375;
  assign n38377 = n38315 & ~n38371;
  assign n38378 = ~pi137 & ~n38377;
  assign n38379 = ~n38282 & ~n38314;
  assign n38380 = ~pi95 & ~n38379;
  assign n38381 = n38365 & ~n38380;
  assign n38382 = pi137 & ~n38381;
  assign n38383 = ~n38378 & ~n38382;
  assign n38384 = pi210 & ~n38383;
  assign n38385 = ~pi146 & ~n38384;
  assign n38386 = ~n38376 & n38385;
  assign n38387 = ~pi234 & ~pi332;
  assign n38388 = n58838 & n38334;
  assign n38389 = ~n58838 & n38299;
  assign n38390 = n2601 & n38302;
  assign n38391 = n58820 & n38257;
  assign n38392 = ~n38389 & n60588;
  assign n38393 = ~n58838 & ~n38299;
  assign n38394 = n58838 & ~n38334;
  assign n38395 = ~n38393 & ~n38394;
  assign n38396 = n60588 & ~n38395;
  assign n38397 = ~n38388 & n38392;
  assign n38398 = ~pi32 & ~n60589;
  assign n38399 = n38372 & ~n38398;
  assign n38400 = ~pi137 & ~n38399;
  assign n38401 = ~n38369 & ~n38400;
  assign n38402 = ~pi210 & ~n38401;
  assign n38403 = ~n38384 & ~n38402;
  assign n38404 = pi146 & n38403;
  assign n38405 = n38387 & ~n38404;
  assign n38406 = ~n38386 & n38405;
  assign n38407 = ~n60587 & ~n38406;
  assign n38408 = ~n2677 & ~n38407;
  assign n38409 = pi234 & n38359;
  assign n38410 = ~pi234 & n38403;
  assign n38411 = ~pi332 & n2677;
  assign n38412 = ~n38410 & n38411;
  assign n38413 = ~n38409 & n38412;
  assign n38414 = pi105 & ~n38413;
  assign n38415 = ~pi332 & ~n38410;
  assign n38416 = ~n38409 & n38415;
  assign n38417 = n2677 & ~n38416;
  assign n38418 = ~n2677 & ~n38406;
  assign n38419 = ~n60587 & n38418;
  assign n38420 = ~n38417 & ~n38419;
  assign n38421 = pi105 & ~n38420;
  assign n38422 = ~n38408 & n38414;
  assign n38423 = ~n38246 & ~n60590;
  assign n38424 = pi228 & ~n38423;
  assign n38425 = ~pi35 & ~n37376;
  assign n38426 = ~pi53 & n38260;
  assign n38427 = ~pi86 & ~n38426;
  assign n38428 = n28411 & ~n38427;
  assign n38429 = n31413 & ~n38428;
  assign n38430 = ~n28628 & ~n38429;
  assign n38431 = ~pi108 & ~n38430;
  assign n38432 = n31410 & ~n38431;
  assign n38433 = ~pi109 & ~n38432;
  assign n38434 = ~n28447 & ~n38433;
  assign n38435 = n2540 & ~n38434;
  assign n38436 = n60541 & ~n38435;
  assign n38437 = n37380 & ~n38436;
  assign n38438 = n37379 & ~n38437;
  assign n38439 = ~pi93 & ~n38438;
  assign n38440 = n38425 & ~n38439;
  assign n38441 = n38301 & ~n38440;
  assign n38442 = n2604 & ~n28320;
  assign n38443 = ~n38441 & n38442;
  assign n38444 = n31408 & ~n38443;
  assign n38445 = n31402 & ~n38444;
  assign n38446 = n31401 & ~n38445;
  assign n38447 = ~n58838 & n38446;
  assign n38448 = pi225 & pi841;
  assign n38449 = n31487 & ~n38448;
  assign n38450 = pi32 & ~n38449;
  assign n38451 = n58838 & n31401;
  assign n38452 = ~pi97 & ~n38429;
  assign n38453 = ~pi108 & ~n38452;
  assign n38454 = n31410 & ~n38453;
  assign n38455 = ~pi109 & ~n38454;
  assign n38456 = ~n28447 & ~n38455;
  assign n38457 = n2540 & ~n38456;
  assign n38458 = n60541 & ~n38457;
  assign n38459 = n37380 & ~n38458;
  assign n38460 = n37379 & ~n38459;
  assign n38461 = ~pi93 & ~n38460;
  assign n38462 = n38425 & ~n38461;
  assign n38463 = n38301 & ~n38462;
  assign n38464 = n38442 & ~n38463;
  assign n38465 = n31408 & ~n38464;
  assign n38466 = n31402 & ~n38465;
  assign n38467 = n38451 & ~n38466;
  assign n38468 = ~n38450 & ~n38467;
  assign n38469 = ~n38447 & n38468;
  assign n38470 = ~pi95 & ~n38469;
  assign n38471 = ~n31400 & ~n38470;
  assign n38472 = ~pi137 & ~n38471;
  assign n38473 = ~pi95 & ~n38450;
  assign n38474 = n2597 & ~n38300;
  assign n38475 = n2597 & n28321;
  assign n38476 = ~n38300 & n38475;
  assign n38477 = n28321 & n38474;
  assign n38478 = ~pi32 & ~n60591;
  assign n38479 = ~pi72 & n2620;
  assign n38480 = n31407 & n38479;
  assign n38481 = n38478 & ~n38480;
  assign n38482 = n38473 & ~n38481;
  assign n38483 = pi137 & ~n28314;
  assign n38484 = ~n38482 & n38483;
  assign n38485 = ~n38472 & ~n38484;
  assign n38486 = ~pi210 & ~n38485;
  assign n38487 = pi146 & n38486;
  assign n38488 = ~pi137 & ~n31400;
  assign n38489 = ~pi225 & n31487;
  assign n38490 = pi32 & ~n38489;
  assign n38491 = ~n38446 & ~n38490;
  assign n38492 = ~pi95 & ~n38491;
  assign n38493 = n38488 & ~n38492;
  assign n38494 = ~pi95 & ~n38490;
  assign n38495 = ~n38481 & n38494;
  assign n38496 = ~n28314 & ~n38495;
  assign n38497 = pi137 & ~n38496;
  assign n38498 = pi210 & ~n38497;
  assign n38499 = ~n38493 & n38498;
  assign n38500 = n38387 & ~n38499;
  assign n38501 = ~pi146 & ~pi210;
  assign n38502 = ~n38446 & ~n38450;
  assign n38503 = ~pi95 & ~n38502;
  assign n38504 = ~n31400 & ~n38503;
  assign n38505 = ~pi137 & ~n38504;
  assign n38506 = ~n38484 & ~n38505;
  assign n38507 = n38501 & ~n38506;
  assign n38508 = n38500 & ~n38507;
  assign n38509 = ~n38487 & n38508;
  assign n38510 = n38473 & ~n38478;
  assign n38511 = pi137 & ~n38510;
  assign n38512 = ~pi72 & ~n38443;
  assign n38513 = n31402 & ~n38512;
  assign n38514 = n31401 & ~n38513;
  assign n38515 = ~n58838 & n38514;
  assign n38516 = ~pi72 & ~n38464;
  assign n38517 = n31402 & ~n38516;
  assign n38518 = n38451 & ~n38517;
  assign n38519 = ~n38450 & ~n38518;
  assign n38520 = ~n38515 & n38519;
  assign n38521 = ~pi95 & ~n38520;
  assign n38522 = n38365 & ~n38521;
  assign n38523 = ~pi137 & ~n38522;
  assign n38524 = ~n38511 & ~n38523;
  assign n38525 = ~pi210 & ~n38524;
  assign n38526 = pi146 & n38525;
  assign n38527 = ~n38490 & ~n38514;
  assign n38528 = ~pi95 & ~n38527;
  assign n38529 = ~pi137 & n38365;
  assign n38530 = ~n38528 & n38529;
  assign n38531 = pi137 & n38494;
  assign n38532 = pi137 & ~n38478;
  assign n38533 = n38494 & n38532;
  assign n38534 = ~n38478 & n38531;
  assign n38535 = pi210 & ~n60592;
  assign n38536 = ~n38530 & n38535;
  assign n38537 = n38327 & ~n38536;
  assign n38538 = ~n38450 & ~n38514;
  assign n38539 = ~pi95 & ~n38538;
  assign n38540 = n38365 & ~n38539;
  assign n38541 = ~pi137 & ~n38540;
  assign n38542 = ~n38511 & ~n38541;
  assign n38543 = n38501 & ~n38542;
  assign n38544 = n38537 & ~n38543;
  assign n38545 = ~n38526 & n38544;
  assign n38546 = ~n2677 & ~n38545;
  assign n38547 = ~n2677 & ~n38509;
  assign n38548 = ~n38545 & n38547;
  assign n38549 = ~n38509 & n38546;
  assign n38550 = ~n38486 & n38500;
  assign n38551 = ~n38525 & n38537;
  assign n38552 = n2677 & ~n38551;
  assign n38553 = ~n38550 & n38552;
  assign n38554 = ~pi153 & ~n38553;
  assign n38555 = ~n60593 & n38554;
  assign n38556 = ~pi109 & ~n38268;
  assign n38557 = ~n28447 & ~n38556;
  assign n38558 = n2540 & ~n38557;
  assign n38559 = n60541 & ~n38558;
  assign n38560 = n37380 & ~n38559;
  assign n38561 = n38274 & ~n38560;
  assign n38562 = n38258 & ~n38561;
  assign n38563 = n38257 & ~n38562;
  assign n38564 = ~pi51 & ~n38563;
  assign n38565 = n38254 & ~n38564;
  assign n38566 = ~pi72 & ~n38565;
  assign n38567 = n31402 & ~n38566;
  assign n38568 = n31401 & ~n38567;
  assign n38569 = ~n38253 & n38568;
  assign n38570 = ~n38290 & ~n38569;
  assign n38571 = ~pi95 & pi137;
  assign n38572 = ~n38570 & n38571;
  assign n38573 = n2793 & ~n28553;
  assign n38574 = n2796 & n38573;
  assign n38575 = n38341 & n38574;
  assign n38576 = n38309 & ~n38574;
  assign n38577 = ~pi137 & ~n38576;
  assign n38578 = ~n38575 & n38577;
  assign n38579 = ~n31400 & ~n38578;
  assign n38580 = ~pi95 & ~n38570;
  assign n38581 = ~n31400 & ~n38580;
  assign n38582 = pi137 & ~n38581;
  assign n38583 = ~n31400 & n38573;
  assign n38584 = n38348 & n38583;
  assign n38585 = ~n38349 & n38573;
  assign n38586 = ~n31400 & n38309;
  assign n38587 = ~n38585 & n38586;
  assign n38588 = ~pi137 & ~n38587;
  assign n38589 = ~pi137 & ~n38584;
  assign n38590 = ~n38587 & n38589;
  assign n38591 = ~n38584 & n38588;
  assign n38592 = ~n38582 & ~n60594;
  assign n38593 = ~n38572 & n38579;
  assign n38594 = ~pi210 & ~n60595;
  assign n38595 = pi234 & ~n38594;
  assign n38596 = ~n38290 & ~n38568;
  assign n38597 = ~pi95 & ~n38596;
  assign n38598 = n38365 & ~n38597;
  assign n38599 = pi137 & ~n38598;
  assign n38600 = ~n28553 & n38400;
  assign n38601 = n28553 & n38374;
  assign n38602 = ~pi210 & ~pi234;
  assign n38603 = ~n38601 & n38602;
  assign n38604 = ~n38600 & n38603;
  assign n38605 = ~n38599 & n38604;
  assign n38606 = ~n38314 & ~n38568;
  assign n38607 = ~pi95 & ~n38606;
  assign n38608 = n38365 & ~n38607;
  assign n38609 = pi137 & ~n38608;
  assign n38610 = pi210 & ~n38378;
  assign n38611 = ~n38609 & n38610;
  assign n38612 = ~n38605 & ~n38611;
  assign n38613 = ~n38595 & n38612;
  assign n38614 = ~n38314 & ~n38569;
  assign n38615 = ~pi95 & ~n38614;
  assign n38616 = pi137 & ~n31400;
  assign n38617 = ~n38615 & n38616;
  assign n38618 = ~n38317 & n38488;
  assign n38619 = pi210 & pi234;
  assign n38620 = ~n38618 & n38619;
  assign n38621 = ~n38617 & n38620;
  assign n38622 = ~n38613 & ~n38621;
  assign n38623 = n38215 & ~n38622;
  assign n38624 = ~pi228 & ~n38623;
  assign n38625 = ~pi228 & ~n38555;
  assign n38626 = ~n38623 & n38625;
  assign n38627 = ~n38555 & n38624;
  assign n38628 = ~n38424 & ~n60596;
  assign n38629 = ~pi216 & ~n38628;
  assign n38630 = ~n38210 & ~n38629;
  assign n38631 = ~pi221 & ~n38630;
  assign n38632 = ~n38226 & ~n38631;
  assign n38633 = ~pi215 & ~n38632;
  assign n38634 = pi299 & ~n38208;
  assign n38635 = ~n38633 & n38634;
  assign n38636 = ~pi224 & pi833;
  assign n38637 = pi222 & ~n38636;
  assign n38638 = ~pi223 & ~n38637;
  assign n38639 = n38207 & ~n38638;
  assign n38640 = pi224 & ~n38209;
  assign n38641 = ~pi222 & ~n38640;
  assign n38642 = ~pi332 & ~pi929;
  assign n38643 = n38636 & n38642;
  assign n38644 = ~n38641 & ~n38643;
  assign n38645 = ~pi223 & ~n38644;
  assign n38646 = ~n38639 & ~n38645;
  assign n38647 = ~pi299 & ~n38646;
  assign n38648 = ~pi223 & n2674;
  assign n38649 = pi198 & ~n38323;
  assign n38650 = ~pi198 & n60586;
  assign n38651 = ~n38649 & ~n38650;
  assign n38652 = pi234 & n38651;
  assign n38653 = pi198 & ~n38383;
  assign n38654 = ~pi198 & ~n38401;
  assign n38655 = ~n38653 & ~n38654;
  assign n38656 = ~pi234 & n38655;
  assign n38657 = ~pi332 & ~n38656;
  assign n38658 = ~n38652 & n38657;
  assign n38659 = n38648 & ~n38658;
  assign n38660 = ~pi198 & ~n38311;
  assign n38661 = ~pi142 & ~n38649;
  assign n38662 = ~n38660 & n38661;
  assign n38663 = pi142 & n38651;
  assign n38664 = n38327 & ~n38663;
  assign n38665 = n38327 & ~n38662;
  assign n38666 = ~n38663 & n38665;
  assign n38667 = ~n38662 & n38664;
  assign n38668 = ~pi223 & ~n2674;
  assign n38669 = ~pi198 & ~n38375;
  assign n38670 = ~pi142 & ~n38653;
  assign n38671 = ~n38669 & n38670;
  assign n38672 = pi142 & n38655;
  assign n38673 = n38387 & ~n38672;
  assign n38674 = ~n38671 & n38673;
  assign n38675 = n38668 & ~n38674;
  assign n38676 = ~n60597 & n38675;
  assign n38677 = ~n38659 & ~n38676;
  assign n38678 = n6544 & ~n38677;
  assign n38679 = n38647 & ~n38678;
  assign n38680 = ~pi39 & ~n38679;
  assign n38681 = ~n38635 & n38680;
  assign n38682 = n35583 & ~n60580;
  assign n38683 = ~n38646 & ~n38682;
  assign n38684 = ~pi299 & ~n38683;
  assign n38685 = pi105 & ~n60580;
  assign n38686 = ~n38246 & ~n38685;
  assign n38687 = pi228 & ~n38686;
  assign n38688 = n38215 & ~n38230;
  assign n38689 = ~pi137 & ~pi153;
  assign n38690 = ~pi332 & n38689;
  assign n38691 = ~pi332 & n58822;
  assign n38692 = n38689 & n38691;
  assign n38693 = n58822 & n38690;
  assign n38694 = ~pi228 & ~n60598;
  assign n38695 = ~pi228 & ~n38688;
  assign n38696 = ~n60598 & n38695;
  assign n38697 = ~n38688 & n38694;
  assign n38698 = ~n38687 & ~n60599;
  assign n38699 = ~pi216 & ~n38698;
  assign n38700 = ~n38210 & ~n38699;
  assign n38701 = ~pi221 & ~n38700;
  assign n38702 = ~n38226 & ~n38701;
  assign n38703 = ~pi215 & ~n38702;
  assign n38704 = ~n38208 & ~n38703;
  assign n38705 = pi299 & ~n38704;
  assign n38706 = ~n38684 & ~n38705;
  assign n38707 = pi39 & ~n38706;
  assign n38708 = ~pi38 & ~n38707;
  assign n38709 = ~n38681 & n38708;
  assign n38710 = n38229 & ~n38241;
  assign n38711 = pi299 & ~n38710;
  assign n38712 = ~n38684 & ~n38711;
  assign n38713 = ~pi39 & ~n38712;
  assign n38714 = n35583 & ~n38213;
  assign n38715 = n38647 & ~n38714;
  assign n38716 = pi299 & n38229;
  assign n38717 = ~n38715 & ~n38716;
  assign n38718 = pi39 & n38717;
  assign n38719 = pi38 & ~n38718;
  assign n38720 = ~n38713 & n38719;
  assign n38721 = ~pi100 & ~n38720;
  assign n38722 = ~n38709 & n38721;
  assign n38723 = n28550 & ~n28553;
  assign n38724 = n28553 & n38230;
  assign n38725 = pi153 & ~n38724;
  assign n38726 = ~n38723 & n38725;
  assign n38727 = ~pi210 & ~n28553;
  assign n38728 = ~pi137 & ~n38727;
  assign n38729 = pi252 & ~n28553;
  assign n38730 = n38728 & ~n38729;
  assign n38731 = n58822 & n38730;
  assign n38732 = ~n38726 & ~n38731;
  assign n38733 = ~pi228 & ~pi332;
  assign n38734 = ~pi137 & pi210;
  assign n38735 = ~pi252 & ~n38734;
  assign n38736 = ~n28553 & n38735;
  assign n38737 = n38691 & n38736;
  assign n38738 = n38215 & ~n38724;
  assign n38739 = ~n38737 & n38738;
  assign n38740 = ~n38727 & ~n38729;
  assign n38741 = n60598 & n38740;
  assign n38742 = ~n38739 & ~n38741;
  assign n38743 = ~pi228 & ~n38742;
  assign n38744 = ~n38732 & n38733;
  assign n38745 = pi228 & ~n38246;
  assign n38746 = pi95 & pi234;
  assign n38747 = ~pi137 & ~n38746;
  assign n38748 = n38728 & ~n38746;
  assign n38749 = ~n38727 & n38747;
  assign n38750 = ~n60579 & ~n60601;
  assign n38751 = ~pi332 & ~n38750;
  assign n38752 = pi105 & ~n38751;
  assign n38753 = n38745 & ~n38752;
  assign n38754 = ~pi216 & ~n38753;
  assign n38755 = ~pi216 & ~n60600;
  assign n38756 = ~n38753 & n38755;
  assign n38757 = ~n60600 & n38754;
  assign n38758 = ~n38210 & ~n60602;
  assign n38759 = ~pi221 & ~n38758;
  assign n38760 = ~n38226 & ~n38759;
  assign n38761 = ~pi215 & ~n38760;
  assign n38762 = ~n38208 & ~n38761;
  assign n38763 = pi299 & ~n38762;
  assign n38764 = pi142 & ~pi198;
  assign n38765 = ~pi137 & ~n38764;
  assign n38766 = n58822 & ~n38765;
  assign n38767 = ~n60579 & ~n38765;
  assign n38768 = n38213 & ~n38767;
  assign n38769 = n38213 & ~n38766;
  assign n38770 = n38668 & ~n60603;
  assign n38771 = ~pi137 & pi198;
  assign n38772 = ~pi95 & n38771;
  assign n38773 = n58822 & ~n38772;
  assign n38774 = n58822 & ~n38771;
  assign n38775 = n38387 & ~n60604;
  assign n38776 = ~n28313 & n38327;
  assign n38777 = ~n38231 & ~n38772;
  assign n38778 = n38327 & ~n38777;
  assign n38779 = ~n60604 & n38776;
  assign n38780 = n38648 & ~n60605;
  assign n38781 = n38648 & ~n38775;
  assign n38782 = ~n60605 & n38781;
  assign n38783 = ~n38775 & n38780;
  assign n38784 = ~n38770 & ~n60606;
  assign n38785 = n6544 & ~n38784;
  assign n38786 = ~n38646 & ~n38785;
  assign n38787 = ~pi299 & ~n38786;
  assign n38788 = n2634 & ~n38787;
  assign n38789 = ~n38763 & n38788;
  assign n38790 = ~n2634 & ~n38717;
  assign n38791 = pi100 & ~n38790;
  assign n38792 = ~n38789 & n38791;
  assign n38793 = ~pi87 & ~n38792;
  assign n38794 = ~n38722 & n38793;
  assign n38795 = ~n58815 & ~n38717;
  assign n38796 = n58815 & n38706;
  assign n38797 = ~n38795 & ~n38796;
  assign n38798 = pi87 & ~n38797;
  assign n38799 = ~pi75 & ~n38798;
  assign n38800 = ~n38794 & n38799;
  assign n38801 = n38217 & ~n38753;
  assign n38802 = ~n38210 & ~n38801;
  assign n38803 = ~pi221 & ~n38802;
  assign n38804 = ~n38226 & ~n38803;
  assign n38805 = ~pi215 & ~n38804;
  assign n38806 = ~n38208 & ~n38805;
  assign n38807 = pi299 & ~n38806;
  assign n38808 = n2672 & ~n38787;
  assign n38809 = ~n38807 & n38808;
  assign n38810 = ~n2672 & ~n38717;
  assign n38811 = pi75 & ~n38810;
  assign n38812 = ~n38809 & n38811;
  assign n38813 = ~n38800 & ~n38812;
  assign n38814 = ~pi92 & ~n38813;
  assign n38815 = n6309 & ~n38797;
  assign n38816 = ~n6309 & ~n38717;
  assign n38817 = pi92 & ~n38816;
  assign n38818 = ~n38815 & n38817;
  assign n38819 = ~pi54 & ~n38818;
  assign n38820 = ~n38814 & n38819;
  assign n38821 = ~n60203 & n38717;
  assign n38822 = n9189 & n38713;
  assign n38823 = ~n38821 & ~n38822;
  assign n38824 = pi54 & n38823;
  assign n38825 = ~pi74 & ~n38824;
  assign n38826 = ~n38820 & n38825;
  assign n38827 = ~pi54 & n38823;
  assign n38828 = pi54 & ~n38717;
  assign n38829 = pi74 & ~n38828;
  assign n38830 = ~n38827 & n38829;
  assign n38831 = ~n38826 & ~n38830;
  assign n38832 = ~pi55 & ~n38831;
  assign n38833 = ~pi332 & n60579;
  assign n38834 = pi105 & ~n38833;
  assign n38835 = n38745 & ~n38834;
  assign n38836 = ~pi228 & n38215;
  assign n38837 = ~n58822 & n38836;
  assign n38838 = ~pi216 & ~n38837;
  assign n38839 = ~n38835 & n38838;
  assign n38840 = ~n38210 & ~n38839;
  assign n38841 = ~pi221 & ~n38840;
  assign n38842 = ~n38226 & ~n38841;
  assign n38843 = ~pi215 & ~n38842;
  assign n38844 = n28288 & ~n38208;
  assign n38845 = ~n38843 & n38844;
  assign n38846 = ~n28288 & n38229;
  assign n38847 = pi55 & ~n38846;
  assign n38848 = ~n38845 & n38847;
  assign n38849 = ~pi56 & ~n38848;
  assign n38850 = ~n38832 & n38849;
  assign n38851 = ~n60070 & n38229;
  assign n38852 = n60070 & n38704;
  assign n38853 = ~n38851 & ~n38852;
  assign n38854 = pi56 & ~n38853;
  assign n38855 = ~pi62 & ~n38854;
  assign n38856 = ~n38850 & n38855;
  assign n38857 = ~pi56 & ~n38853;
  assign n38858 = pi56 & n38229;
  assign n38859 = pi62 & ~n38858;
  assign n38860 = ~n38857 & n38859;
  assign n38861 = ~pi59 & ~n38860;
  assign n38862 = ~n38856 & n38861;
  assign n38863 = pi59 & n38229;
  assign n38864 = ~n38242 & n38863;
  assign n38865 = ~pi57 & ~n38864;
  assign n38866 = ~n38862 & n38865;
  assign n38867 = ~n38245 & ~n38866;
  assign n38868 = n28570 & n37226;
  assign n38869 = n37361 & n38868;
  assign n38870 = pi24 & ~pi94;
  assign n38871 = n58798 & n38870;
  assign n38872 = pi24 & n59134;
  assign n38873 = ~n36404 & ~n60607;
  assign n38874 = ~n37316 & n38870;
  assign n38875 = pi252 & n35649;
  assign n38876 = ~pi252 & ~n32496;
  assign n38877 = pi252 & ~n35649;
  assign n38878 = ~pi252 & n32496;
  assign n38879 = ~n38877 & ~n38878;
  assign n38880 = ~n38875 & ~n38876;
  assign n38881 = n60165 & ~n60608;
  assign n38882 = ~n38874 & n38881;
  assign n38883 = ~n38873 & n38882;
  assign n38884 = pi24 & ~pi90;
  assign n38885 = n32914 & n38884;
  assign n38886 = n60608 & n38885;
  assign n38887 = n37318 & n38886;
  assign n38888 = ~n38883 & ~n38887;
  assign n38889 = ~pi100 & ~n38888;
  assign n38890 = pi100 & n60087;
  assign n38891 = n31666 & n38890;
  assign n38892 = ~n38889 & ~n38891;
  assign n38893 = ~pi75 & n30890;
  assign n38894 = n2634 & n6309;
  assign n38895 = ~n38892 & n60609;
  assign n38896 = ~n38869 & ~n38895;
  assign po208 = n37304 & ~n38896;
  assign n38898 = n2681 & n28557;
  assign n38899 = n60523 & ~n38898;
  assign n38900 = pi129 & ~n38899;
  assign n38901 = ~n60087 & ~n38900;
  assign n38902 = ~n2681 & n60523;
  assign n38903 = pi129 & ~n38902;
  assign n38904 = n2679 & ~n38903;
  assign n38905 = pi129 & ~n60523;
  assign n38906 = ~n28557 & ~n38905;
  assign n38907 = ~n28566 & ~n38906;
  assign n38908 = ~n38904 & n38907;
  assign n38909 = ~n28566 & ~n38901;
  assign n38910 = ~pi75 & n2671;
  assign n38911 = n28548 & n38910;
  assign n38912 = ~n60610 & n38911;
  assign n38913 = ~n35649 & n37227;
  assign n38914 = ~n37228 & n38913;
  assign n38915 = ~n38912 & ~n38914;
  assign n38916 = n37304 & ~n38915;
  assign po258 = n58822 & n38916;
  assign n38918 = pi51 & n2680;
  assign n38919 = ~pi146 & n38918;
  assign n38920 = pi161 & ~n38919;
  assign n38921 = n2456 & n32880;
  assign n38922 = ~pi51 & n38921;
  assign n38923 = n2680 & ~n38922;
  assign n38924 = pi51 & pi146;
  assign n38925 = n38923 & ~n38924;
  assign n38926 = ~n38920 & ~n38924;
  assign n38927 = n38923 & n38926;
  assign n38928 = ~n38920 & n38925;
  assign n38929 = ~pi87 & ~n60611;
  assign n38930 = pi87 & ~n30546;
  assign n38931 = pi232 & ~n38930;
  assign n38932 = ~n38929 & n38931;
  assign n38933 = ~pi134 & ~pi135;
  assign n38934 = ~pi136 & n38933;
  assign n38935 = ~pi130 & n38934;
  assign n38936 = ~pi132 & n38935;
  assign n38937 = ~pi126 & n38936;
  assign n38938 = ~pi121 & n38937;
  assign n38939 = ~pi125 & ~pi133;
  assign n38940 = pi121 & ~n38939;
  assign n38941 = ~pi121 & n38939;
  assign n38942 = ~n38940 & ~n38941;
  assign n38943 = ~n38938 & ~n38942;
  assign n38944 = ~pi87 & n38922;
  assign n38945 = ~n38943 & n38944;
  assign n38946 = ~n58992 & ~n38945;
  assign n38947 = ~n58992 & ~n38932;
  assign n38948 = ~n38945 & n38947;
  assign n38949 = ~n38932 & n38946;
  assign n38950 = ~pi142 & n38918;
  assign n38951 = pi144 & ~n38950;
  assign n38952 = pi51 & pi142;
  assign n38953 = n38923 & ~n38952;
  assign n38954 = ~n38951 & n38953;
  assign n38955 = ~pi299 & ~n38954;
  assign n38956 = pi299 & ~n60611;
  assign n38957 = pi232 & ~n38956;
  assign n38958 = pi232 & ~n38955;
  assign n38959 = ~n38956 & n38958;
  assign n38960 = ~n38955 & n38957;
  assign n38961 = pi38 & ~n60613;
  assign n38962 = ~pi100 & ~n38961;
  assign n38963 = pi38 & ~n38922;
  assign n38964 = ~pi100 & ~n38963;
  assign n38965 = ~n38962 & ~n38964;
  assign n38966 = n2458 & n28344;
  assign n38967 = n2447 & n2562;
  assign n38968 = n32879 & n38967;
  assign n38969 = n38966 & n38968;
  assign n38970 = pi77 & ~pi86;
  assign n38971 = n2447 & n32879;
  assign n38972 = n38966 & n38971;
  assign n38973 = ~pi50 & pi77;
  assign n38974 = n2503 & n38973;
  assign n38975 = n38972 & n38974;
  assign n38976 = n38969 & n38970;
  assign n38977 = ~pi24 & pi314;
  assign n38978 = n59135 & n38977;
  assign n38979 = ~pi24 & n58798;
  assign n38980 = ~pi94 & n38979;
  assign n38981 = ~pi24 & n59134;
  assign n38982 = pi314 & n59135;
  assign n38983 = n60615 & n38982;
  assign n38984 = n59134 & n38978;
  assign n38985 = n60614 & n60616;
  assign n38986 = n2599 & n38985;
  assign n38987 = ~n59135 & n38921;
  assign n38988 = ~pi51 & ~n38987;
  assign n38989 = n58802 & n38972;
  assign n38990 = ~pi77 & n38969;
  assign n38991 = pi86 & n60617;
  assign n38992 = ~n60614 & ~n38991;
  assign n38993 = n60607 & ~n38992;
  assign n38994 = pi86 & n59134;
  assign n38995 = ~pi24 & n38994;
  assign n38996 = n60615 & n38991;
  assign n38997 = n60617 & n38995;
  assign n38998 = n38921 & ~n60618;
  assign n38999 = ~n38993 & n38998;
  assign n39000 = n38988 & ~n38999;
  assign n39001 = n2599 & n39000;
  assign n39002 = n38922 & ~n39001;
  assign n39003 = ~pi58 & n59135;
  assign n39004 = n2502 & n39003;
  assign n39005 = n60617 & n39004;
  assign n39006 = pi72 & n2621;
  assign n39007 = n39005 & n39006;
  assign n39008 = n39002 & ~n39007;
  assign n39009 = ~n38986 & n39008;
  assign n39010 = ~n2680 & n39009;
  assign n39011 = n58834 & n38994;
  assign n39012 = ~pi24 & ~n39011;
  assign n39013 = n2532 & n32896;
  assign n39014 = pi24 & ~n39013;
  assign n39015 = ~n39012 & ~n39014;
  assign n39016 = ~pi314 & ~n39015;
  assign n39017 = pi314 & ~n39013;
  assign n39018 = ~n39016 & ~n39017;
  assign n39019 = n60073 & n39018;
  assign n39020 = ~pi72 & ~n39019;
  assign n39021 = n28319 & ~n39020;
  assign n39022 = n2680 & ~n39021;
  assign n39023 = ~n39010 & ~n39022;
  assign n39024 = ~pi142 & ~n39023;
  assign n39025 = ~n2680 & ~n39009;
  assign n39026 = n2580 & n58818;
  assign n39027 = n2581 & n58809;
  assign n39028 = n39018 & n60619;
  assign n39029 = ~pi51 & ~n39028;
  assign n39030 = pi72 & n36495;
  assign n39031 = n39029 & ~n39030;
  assign n39032 = n2680 & ~n39031;
  assign n39033 = ~n39025 & ~n39032;
  assign n39034 = pi142 & n39033;
  assign n39035 = ~pi144 & ~n39034;
  assign n39036 = ~pi144 & ~n39024;
  assign n39037 = ~n39034 & n39036;
  assign n39038 = ~n39024 & n39035;
  assign n39039 = n38951 & ~n39009;
  assign n39040 = ~pi180 & ~n39039;
  assign n39041 = ~n60620 & n39040;
  assign n39042 = n60073 & n39015;
  assign n39043 = ~pi72 & ~n39042;
  assign n39044 = n28319 & ~n39043;
  assign n39045 = n2680 & ~n39044;
  assign n39046 = ~n39010 & ~n39045;
  assign n39047 = ~pi142 & ~n39046;
  assign n39048 = n2599 & n2680;
  assign n39049 = n2597 & n29755;
  assign n39050 = n39042 & n60621;
  assign n39051 = ~n38918 & ~n39030;
  assign n39052 = n2680 & ~n39051;
  assign n39053 = ~n39050 & ~n39052;
  assign n39054 = ~n39025 & n39053;
  assign n39055 = pi142 & n39054;
  assign n39056 = ~pi144 & ~n39055;
  assign n39057 = ~n39047 & n39056;
  assign n39058 = ~pi51 & ~n38921;
  assign n39059 = n2680 & n39058;
  assign n39060 = ~n60621 & ~n39059;
  assign n39061 = n2599 & ~n39000;
  assign n39062 = ~n39060 & ~n39061;
  assign n39063 = pi142 & ~n39062;
  assign n39064 = n2680 & ~n39002;
  assign n39065 = ~pi142 & ~n39064;
  assign n39066 = ~n39063 & ~n39065;
  assign n39067 = n38922 & ~n38986;
  assign n39068 = ~n39001 & n39067;
  assign n39069 = ~n2680 & ~n39068;
  assign n39070 = ~n38923 & ~n39069;
  assign n39071 = ~n39066 & ~n39070;
  assign n39072 = ~pi51 & n2680;
  assign n39073 = ~n39008 & n39072;
  assign n39074 = ~n39025 & ~n39073;
  assign n39075 = ~n39071 & n39074;
  assign n39076 = pi144 & ~n39075;
  assign n39077 = pi180 & ~n39076;
  assign n39078 = ~n39057 & n39077;
  assign n39079 = ~pi179 & ~n39078;
  assign n39080 = ~n60620 & ~n39039;
  assign n39081 = ~pi180 & ~n39080;
  assign n39082 = ~pi142 & n39046;
  assign n39083 = pi142 & ~n39054;
  assign n39084 = ~pi144 & ~n39083;
  assign n39085 = ~n39082 & n39084;
  assign n39086 = pi144 & n39074;
  assign n39087 = ~n39071 & n39086;
  assign n39088 = pi180 & ~n39087;
  assign n39089 = ~n39085 & n39088;
  assign n39090 = ~n39081 & ~n39089;
  assign n39091 = ~pi179 & ~n39090;
  assign n39092 = ~n39041 & n39079;
  assign n39093 = n2501 & n58798;
  assign n39094 = ~pi86 & n59134;
  assign n39095 = n32869 & n60623;
  assign n39096 = n28338 & n32503;
  assign n39097 = ~pi24 & ~pi51;
  assign n39098 = ~pi51 & n38978;
  assign n39099 = n38982 & n39097;
  assign n39100 = pi314 & n60623;
  assign n39101 = n32869 & n39100;
  assign n39102 = ~pi24 & n60073;
  assign n39103 = n39101 & n39102;
  assign n39104 = n60624 & n60625;
  assign n39105 = ~pi72 & ~n60626;
  assign n39106 = n28319 & ~n39105;
  assign n39107 = n2680 & ~n39106;
  assign n39108 = ~n39010 & ~n39107;
  assign n39109 = ~pi142 & ~n39108;
  assign n39110 = n60621 & n60626;
  assign n39111 = ~n39025 & ~n39052;
  assign n39112 = ~n39110 & n39111;
  assign n39113 = pi142 & n39112;
  assign n39114 = ~pi144 & ~n39113;
  assign n39115 = ~pi144 & ~n39109;
  assign n39116 = ~n39113 & n39115;
  assign n39117 = ~n39109 & n39114;
  assign n39118 = ~n39007 & n39070;
  assign n39119 = ~n38986 & n39118;
  assign n39120 = n38951 & ~n39119;
  assign n39121 = ~pi180 & ~n39120;
  assign n39122 = ~n60627 & n39121;
  assign n39123 = ~pi144 & n39111;
  assign n39124 = pi144 & n39118;
  assign n39125 = ~n38950 & ~n39124;
  assign n39126 = pi144 & ~n39118;
  assign n39127 = ~pi144 & ~n39111;
  assign n39128 = ~n39126 & ~n39127;
  assign n39129 = ~n38950 & ~n39128;
  assign n39130 = ~n39123 & n39125;
  assign n39131 = pi180 & ~n60628;
  assign n39132 = pi179 & ~n39131;
  assign n39133 = ~n39122 & n39132;
  assign n39134 = ~n60622 & ~n39133;
  assign n39135 = ~pi299 & ~n39134;
  assign n39136 = ~pi161 & ~n38919;
  assign n39137 = ~n39111 & n39136;
  assign n39138 = pi146 & n39118;
  assign n39139 = n38921 & ~n39007;
  assign n39140 = n39072 & ~n39139;
  assign n39141 = ~pi146 & ~n39140;
  assign n39142 = ~n39025 & n39141;
  assign n39143 = pi161 & ~n39142;
  assign n39144 = pi161 & ~n39138;
  assign n39145 = ~n39142 & n39144;
  assign n39146 = ~n39138 & n39143;
  assign n39147 = ~n39137 & ~n60629;
  assign n39148 = n31099 & ~n39147;
  assign n39149 = ~pi146 & ~n39108;
  assign n39150 = pi146 & n39112;
  assign n39151 = ~pi161 & ~n39150;
  assign n39152 = ~pi161 & ~n39149;
  assign n39153 = ~n39150 & n39152;
  assign n39154 = ~n39149 & n39151;
  assign n39155 = n39072 & n39139;
  assign n39156 = ~n38986 & n39155;
  assign n39157 = ~n38918 & ~n39156;
  assign n39158 = pi146 & ~n38922;
  assign n39159 = ~n39157 & ~n39158;
  assign n39160 = pi161 & ~n39159;
  assign n39161 = ~n39010 & n39160;
  assign n39162 = ~n60630 & ~n39161;
  assign n39163 = n31084 & ~n39162;
  assign n39164 = ~n39148 & ~n39163;
  assign n39165 = pi156 & ~n39164;
  assign n39166 = ~pi146 & ~n39023;
  assign n39167 = pi146 & n39033;
  assign n39168 = n31084 & ~n39167;
  assign n39169 = n31084 & ~n39166;
  assign n39170 = ~n39167 & n39169;
  assign n39171 = ~n39166 & n39168;
  assign n39172 = ~pi146 & ~n39046;
  assign n39173 = pi146 & n39054;
  assign n39174 = n31099 & ~n39173;
  assign n39175 = ~n39172 & n39174;
  assign n39176 = ~pi161 & ~n39175;
  assign n39177 = ~n60631 & n39176;
  assign n39178 = pi146 & ~n39062;
  assign n39179 = ~pi146 & ~n39064;
  assign n39180 = ~n39178 & ~n39179;
  assign n39181 = ~n39070 & ~n39180;
  assign n39182 = n39074 & ~n39181;
  assign n39183 = n31099 & ~n39182;
  assign n39184 = n31084 & ~n38919;
  assign n39185 = ~n39009 & n39184;
  assign n39186 = pi161 & ~n39185;
  assign n39187 = ~n39183 & n39186;
  assign n39188 = ~pi156 & ~n39187;
  assign n39189 = ~n39177 & n39188;
  assign n39190 = ~n39165 & ~n39189;
  assign n39191 = ~n39135 & n39190;
  assign n39192 = n29912 & ~n39191;
  assign n39193 = n2599 & n39005;
  assign n39194 = n38922 & ~n39193;
  assign n39195 = ~n38919 & ~n39194;
  assign n39196 = pi161 & ~n39195;
  assign n39197 = ~n2680 & ~n39194;
  assign n39198 = n2593 & n58818;
  assign n39199 = n58808 & n58809;
  assign n39200 = ~pi51 & ~n60632;
  assign n39201 = n2680 & ~n39200;
  assign n39202 = ~n39197 & ~n39201;
  assign n39203 = pi146 & ~n39202;
  assign n39204 = ~n29911 & ~n39197;
  assign n39205 = ~pi146 & ~n39204;
  assign n39206 = ~pi161 & ~n39205;
  assign n39207 = ~pi161 & ~n39203;
  assign n39208 = ~n39205 & n39207;
  assign n39209 = ~n39203 & n39206;
  assign n39210 = ~n39196 & ~n60633;
  assign n39211 = n2852 & ~n39210;
  assign n39212 = ~n29532 & ~n39211;
  assign n39213 = ~pi287 & n2680;
  assign n39214 = ~pi51 & n39213;
  assign n39215 = ~n39202 & ~n39214;
  assign n39216 = n39136 & n39215;
  assign n39217 = n39193 & ~n39213;
  assign n39218 = n38922 & ~n39217;
  assign n39219 = n38920 & ~n39218;
  assign n39220 = ~n39216 & ~n39219;
  assign n39221 = pi216 & ~n39220;
  assign n39222 = ~n39212 & ~n39221;
  assign n39223 = ~n38922 & ~n60611;
  assign n39224 = ~n2852 & ~n39223;
  assign n39225 = n29502 & ~n39224;
  assign n39226 = ~n39222 & n39225;
  assign n39227 = pi142 & ~n39202;
  assign n39228 = ~pi142 & ~n39204;
  assign n39229 = n2829 & ~n39228;
  assign n39230 = n2829 & ~n39227;
  assign n39231 = ~n39228 & n39230;
  assign n39232 = ~n39227 & n39229;
  assign n39233 = ~n29572 & ~n60634;
  assign n39234 = pi224 & ~n38950;
  assign n39235 = n39215 & n39234;
  assign n39236 = ~n39233 & ~n39235;
  assign n39237 = ~n38922 & ~n38950;
  assign n39238 = ~n2829 & ~n39237;
  assign n39239 = pi144 & ~n39238;
  assign n39240 = ~n2829 & n39059;
  assign n39241 = ~n39238 & ~n39240;
  assign n39242 = ~n39239 & n39241;
  assign n39243 = ~n39236 & n39242;
  assign n39244 = ~pi51 & ~n39194;
  assign n39245 = ~pi287 & ~n39244;
  assign n39246 = ~n39059 & ~n39213;
  assign n39247 = ~n39245 & ~n39246;
  assign n39248 = ~n38953 & ~n39247;
  assign n39249 = n29572 & ~n39248;
  assign n39250 = n38921 & n39249;
  assign n39251 = pi51 & ~n2680;
  assign n39252 = ~n39244 & ~n39251;
  assign n39253 = n2829 & ~n38952;
  assign n39254 = n39252 & n39253;
  assign n39255 = n39239 & ~n39254;
  assign n39256 = ~n39250 & n39255;
  assign n39257 = pi181 & ~n39256;
  assign n39258 = ~n39243 & n39257;
  assign n39259 = ~n60634 & n39242;
  assign n39260 = ~pi181 & ~n39255;
  assign n39261 = ~n39259 & n39260;
  assign n39262 = ~pi299 & ~n39261;
  assign n39263 = ~n39258 & n39262;
  assign n39264 = n29424 & ~n39224;
  assign n39265 = ~n39211 & n39264;
  assign n39266 = pi232 & ~n39265;
  assign n39267 = ~n39263 & n39266;
  assign n39268 = ~n39226 & n39267;
  assign n39269 = ~n58844 & ~n2853;
  assign n39270 = n39193 & ~n39269;
  assign n39271 = ~pi232 & n38922;
  assign n39272 = ~n39270 & n39271;
  assign n39273 = pi39 & ~n39272;
  assign n39274 = ~n39268 & n39273;
  assign n39275 = ~pi39 & ~pi232;
  assign n39276 = ~n39009 & n39275;
  assign n39277 = ~n39274 & ~n39276;
  assign n39278 = ~n39192 & n39277;
  assign n39279 = ~pi38 & ~n39278;
  assign n39280 = ~n38965 & ~n39279;
  assign n39281 = pi100 & n60613;
  assign n39282 = pi100 & n38922;
  assign n39283 = n6311 & ~n39282;
  assign n39284 = ~n39281 & n39283;
  assign n39285 = ~n39280 & n39284;
  assign n39286 = ~pi87 & ~n6308;
  assign n39287 = ~n38922 & n39286;
  assign n39288 = ~n60613 & n39287;
  assign n39289 = ~pi184 & ~pi299;
  assign n39290 = ~n34428 & ~n39289;
  assign n39291 = n2681 & n39290;
  assign n39292 = pi87 & ~n39291;
  assign n39293 = ~n38943 & ~n39292;
  assign n39294 = ~n39288 & n39293;
  assign n39295 = ~n39285 & n39294;
  assign n39296 = n2680 & ~n39029;
  assign n39297 = ~n38952 & n39296;
  assign n39298 = pi144 & ~n39297;
  assign n39299 = n38921 & ~n38985;
  assign n39300 = n59135 & n39299;
  assign n39301 = n38999 & n39300;
  assign n39302 = n38988 & ~n39301;
  assign n39303 = n2599 & ~n39302;
  assign n39304 = ~n39060 & ~n39303;
  assign n39305 = pi142 & n39304;
  assign n39306 = n2680 & ~n39068;
  assign n39307 = ~pi142 & n39306;
  assign n39308 = ~pi144 & ~n39307;
  assign n39309 = ~n39305 & n39308;
  assign n39310 = pi180 & ~n39309;
  assign n39311 = ~n39298 & n39310;
  assign n39312 = n38951 & ~n39050;
  assign n39313 = ~pi144 & ~n39066;
  assign n39314 = ~pi180 & ~n39313;
  assign n39315 = ~n39312 & n39314;
  assign n39316 = pi179 & ~n39315;
  assign n39317 = ~n39311 & n39316;
  assign n39318 = n38951 & ~n39110;
  assign n39319 = ~pi51 & ~n39299;
  assign n39320 = n2599 & ~n39319;
  assign n39321 = ~n39060 & ~n39320;
  assign n39322 = pi142 & n39321;
  assign n39323 = n2680 & ~n39067;
  assign n39324 = ~pi142 & n39323;
  assign n39325 = ~pi144 & ~n39324;
  assign n39326 = ~n39322 & n39325;
  assign n39327 = pi180 & ~n39326;
  assign n39328 = ~n39318 & n39327;
  assign n39329 = ~pi180 & n38954;
  assign n39330 = ~pi179 & ~n39329;
  assign n39331 = ~n39328 & n39330;
  assign n39332 = ~n39317 & ~n39331;
  assign n39333 = ~pi299 & ~n39332;
  assign n39334 = ~n38924 & n39296;
  assign n39335 = pi161 & ~n39334;
  assign n39336 = ~pi146 & n39306;
  assign n39337 = pi146 & n39304;
  assign n39338 = ~pi161 & ~n39337;
  assign n39339 = ~pi161 & ~n39336;
  assign n39340 = ~n39337 & n39339;
  assign n39341 = ~n39336 & n39338;
  assign n39342 = ~n39335 & ~n60635;
  assign n39343 = n31099 & ~n39342;
  assign n39344 = n38920 & ~n39050;
  assign n39345 = ~pi161 & ~n39180;
  assign n39346 = ~n39344 & ~n39345;
  assign n39347 = n31084 & ~n39346;
  assign n39348 = pi232 & ~n39347;
  assign n39349 = ~n39343 & n39348;
  assign n39350 = pi156 & ~n39349;
  assign n39351 = ~pi39 & ~n39350;
  assign n39352 = ~pi39 & ~n39333;
  assign n39353 = ~n39350 & n39352;
  assign n39354 = ~n39333 & n39351;
  assign n39355 = ~pi144 & ~n38953;
  assign n39356 = ~n39249 & n39355;
  assign n39357 = n29572 & n39213;
  assign n39358 = ~n38952 & n39357;
  assign n39359 = ~pi142 & ~n60632;
  assign n39360 = pi142 & ~n58822;
  assign n39361 = n39357 & ~n39360;
  assign n39362 = ~n39359 & n39361;
  assign n39363 = n60632 & n39358;
  assign n39364 = n38951 & ~n60637;
  assign n39365 = pi181 & ~n39364;
  assign n39366 = pi181 & ~n39356;
  assign n39367 = ~n39364 & n39366;
  assign n39368 = ~n39356 & n39365;
  assign n39369 = ~pi181 & n38954;
  assign n39370 = ~pi299 & ~n39369;
  assign n39371 = ~n60638 & n39370;
  assign n39372 = n2680 & n2801;
  assign n39373 = n38920 & ~n39372;
  assign n39374 = n39136 & ~n39247;
  assign n39375 = n29532 & ~n39374;
  assign n39376 = ~n39373 & n39375;
  assign n39377 = ~n29532 & n60611;
  assign n39378 = n29502 & ~n39377;
  assign n39379 = ~n39376 & n39378;
  assign n39380 = ~pi159 & n38956;
  assign n39381 = n31239 & ~n39380;
  assign n39382 = ~n39379 & n39381;
  assign n39383 = ~n39371 & n39382;
  assign n39384 = ~pi38 & ~n39383;
  assign n39385 = ~n60636 & n39384;
  assign n39386 = n38920 & ~n39110;
  assign n39387 = pi146 & n39321;
  assign n39388 = ~pi146 & n39323;
  assign n39389 = ~pi161 & ~n39388;
  assign n39390 = ~n39387 & n39389;
  assign n39391 = ~n39386 & ~n39390;
  assign n39392 = n31099 & ~n39391;
  assign n39393 = ~pi158 & n38956;
  assign n39394 = pi232 & ~n39393;
  assign n39395 = ~n39392 & n39394;
  assign n39396 = ~pi156 & n2634;
  assign n39397 = ~n39395 & n39396;
  assign n39398 = n38962 & ~n39397;
  assign n39399 = ~n39385 & n39398;
  assign n39400 = n6311 & ~n39281;
  assign n39401 = ~n39399 & n39400;
  assign n39402 = ~n60613 & n39286;
  assign n39403 = n38943 & ~n39292;
  assign n39404 = ~n39402 & n39403;
  assign n39405 = ~n39401 & n39404;
  assign n39406 = n58992 & ~n39405;
  assign n39407 = ~n39295 & n39406;
  assign n39408 = ~n60612 & ~n39407;
  assign n39409 = ~pi125 & n38938;
  assign n39410 = pi125 & pi133;
  assign n39411 = ~n38939 & ~n39410;
  assign n39412 = ~n39409 & ~n39411;
  assign n39413 = n38922 & ~n39412;
  assign n39414 = pi172 & n38918;
  assign n39415 = ~pi152 & n39059;
  assign n39416 = ~n39414 & ~n39415;
  assign n39417 = pi232 & ~n39416;
  assign n39418 = ~n39413 & ~n39417;
  assign n39419 = ~pi87 & ~n39418;
  assign n39420 = pi87 & n2681;
  assign n39421 = pi162 & n39420;
  assign n39422 = ~n58992 & ~n39421;
  assign n39423 = ~n39419 & n39422;
  assign n39424 = ~pi152 & n2680;
  assign n39425 = n39030 & ~n39424;
  assign n39426 = ~pi152 & n39140;
  assign n39427 = ~pi197 & ~n39426;
  assign n39428 = ~n39425 & n39427;
  assign n39429 = ~n2680 & n39030;
  assign n39430 = ~n39072 & ~n39429;
  assign n39431 = ~n39156 & ~n39430;
  assign n39432 = ~pi152 & pi197;
  assign n39433 = ~n39431 & n39432;
  assign n39434 = ~n39428 & ~n39433;
  assign n39435 = ~n39414 & ~n39434;
  assign n39436 = ~n2680 & ~n39030;
  assign n39437 = ~n39107 & ~n39436;
  assign n39438 = ~pi172 & n39437;
  assign n39439 = ~n38918 & ~n39110;
  assign n39440 = ~n39030 & n39439;
  assign n39441 = n39051 & ~n39110;
  assign n39442 = pi172 & ~n60639;
  assign n39443 = pi152 & pi197;
  assign n39444 = ~n39442 & n39443;
  assign n39445 = ~n39438 & n39444;
  assign n39446 = ~n39435 & ~n39445;
  assign n39447 = n29555 & ~n39446;
  assign n39448 = ~n39022 & ~n39436;
  assign n39449 = ~pi172 & n39448;
  assign n39450 = ~n39031 & ~n39436;
  assign n39451 = pi172 & n39450;
  assign n39452 = pi152 & ~n39451;
  assign n39453 = ~n39449 & n39452;
  assign n39454 = n2680 & n39009;
  assign n39455 = ~n39430 & ~n39454;
  assign n39456 = ~pi152 & ~n39414;
  assign n39457 = ~n39455 & n39456;
  assign n39458 = pi197 & ~n39457;
  assign n39459 = ~n39414 & ~n39455;
  assign n39460 = ~pi152 & ~n39459;
  assign n39461 = ~pi172 & ~n39448;
  assign n39462 = pi172 & ~n39450;
  assign n39463 = pi152 & ~n39462;
  assign n39464 = ~n39461 & n39463;
  assign n39465 = ~n39460 & ~n39464;
  assign n39466 = pi197 & ~n39465;
  assign n39467 = ~n39453 & n39458;
  assign n39468 = ~n39045 & ~n39436;
  assign n39469 = pi152 & n39468;
  assign n39470 = ~n39073 & ~n39429;
  assign n39471 = ~pi152 & ~n39470;
  assign n39472 = ~pi172 & ~n39471;
  assign n39473 = ~n39469 & n39472;
  assign n39474 = ~n39050 & n39051;
  assign n39475 = pi152 & ~n39474;
  assign n39476 = n39008 & n39155;
  assign n39477 = n39002 & n39155;
  assign n39478 = ~n39436 & ~n60641;
  assign n39479 = ~pi152 & n39478;
  assign n39480 = pi172 & ~n39479;
  assign n39481 = ~n39475 & n39480;
  assign n39482 = ~pi197 & ~n39481;
  assign n39483 = ~n39473 & n39482;
  assign n39484 = n29564 & ~n39483;
  assign n39485 = ~n60640 & n39484;
  assign n39486 = ~n39447 & ~n39485;
  assign n39487 = pi299 & ~n39486;
  assign n39488 = pi145 & n39437;
  assign n39489 = ~pi145 & n39030;
  assign n39490 = pi174 & ~n39489;
  assign n39491 = ~n39488 & n39490;
  assign n39492 = pi145 & n39431;
  assign n39493 = ~n39140 & ~n39429;
  assign n39494 = ~pi145 & ~n39493;
  assign n39495 = ~pi174 & ~n39494;
  assign n39496 = ~n39492 & n39495;
  assign n39497 = ~n39491 & ~n39496;
  assign n39498 = ~pi193 & ~n39497;
  assign n39499 = ~pi145 & n39110;
  assign n39500 = pi174 & ~n60639;
  assign n39501 = ~n39439 & ~n39499;
  assign n39502 = ~n39030 & ~n39501;
  assign n39503 = pi174 & ~n39502;
  assign n39504 = ~n39499 & n39500;
  assign n39505 = ~n38918 & ~n38986;
  assign n39506 = pi145 & ~n39505;
  assign n39507 = n39155 & ~n39506;
  assign n39508 = ~pi174 & ~n39507;
  assign n39509 = ~n39436 & n39508;
  assign n39510 = pi193 & ~n39509;
  assign n39511 = ~n60642 & n39510;
  assign n39512 = ~n39498 & ~n39511;
  assign n39513 = n29581 & ~n39512;
  assign n39514 = pi145 & n39448;
  assign n39515 = ~pi145 & n39468;
  assign n39516 = ~pi193 & ~n39515;
  assign n39517 = ~n39514 & n39516;
  assign n39518 = pi145 & n39450;
  assign n39519 = ~pi145 & ~n39474;
  assign n39520 = pi193 & ~n39519;
  assign n39521 = ~n39518 & n39520;
  assign n39522 = pi174 & ~n39521;
  assign n39523 = pi145 & ~n39450;
  assign n39524 = ~pi145 & n39474;
  assign n39525 = pi193 & ~n39524;
  assign n39526 = ~n39523 & n39525;
  assign n39527 = pi145 & ~n39448;
  assign n39528 = ~pi145 & ~n39468;
  assign n39529 = ~pi193 & ~n39528;
  assign n39530 = ~n39527 & n39529;
  assign n39531 = ~n39526 & ~n39530;
  assign n39532 = pi174 & ~n39531;
  assign n39533 = ~n39517 & n39522;
  assign n39534 = ~pi193 & ~n39470;
  assign n39535 = pi193 & n39478;
  assign n39536 = ~pi145 & ~n39535;
  assign n39537 = ~pi145 & ~n39534;
  assign n39538 = ~n39535 & n39537;
  assign n39539 = ~n39534 & n39536;
  assign n39540 = pi193 & n38918;
  assign n39541 = pi145 & ~n39540;
  assign n39542 = ~n39455 & n39541;
  assign n39543 = ~pi174 & ~n39542;
  assign n39544 = ~n60644 & n39543;
  assign n39545 = n29601 & ~n39544;
  assign n39546 = ~n60643 & n39545;
  assign n39547 = ~n39513 & ~n39546;
  assign n39548 = ~pi38 & ~n39547;
  assign n39549 = ~n39487 & ~n39548;
  assign n39550 = n29912 & ~n39549;
  assign n39551 = ~pi299 & ~n3890;
  assign n39552 = pi299 & ~n3906;
  assign n39553 = ~n39551 & ~n39552;
  assign n39554 = ~n58845 & ~n58848;
  assign n39555 = n58822 & n60645;
  assign n39556 = ~pi232 & ~n39555;
  assign n39557 = pi39 & ~n39556;
  assign n39558 = n60632 & n39213;
  assign n39559 = ~n38918 & ~n39558;
  assign n39560 = pi224 & n39559;
  assign n39561 = n2829 & ~n39560;
  assign n39562 = n58822 & ~n2680;
  assign n39563 = ~n39201 & ~n39562;
  assign n39564 = ~n39200 & ~n39251;
  assign n39565 = n3890 & n60646;
  assign n39566 = n39561 & ~n39565;
  assign n39567 = ~n38918 & ~n39566;
  assign n39568 = pi174 & ~n39567;
  assign n39569 = n2680 & ~n39194;
  assign n39570 = ~n39562 & ~n39569;
  assign n39571 = n3890 & n39570;
  assign n39572 = n39193 & n39213;
  assign n39573 = pi224 & ~n39572;
  assign n39574 = n2829 & ~n39573;
  assign n39575 = ~n38923 & ~n39574;
  assign n39576 = ~n39571 & ~n39575;
  assign n39577 = ~pi174 & n39576;
  assign n39578 = pi193 & ~n39577;
  assign n39579 = ~n39568 & n39578;
  assign n39580 = n2680 & n39244;
  assign n39581 = ~n39562 & ~n39580;
  assign n39582 = ~pi224 & n39581;
  assign n39583 = pi224 & ~n39247;
  assign n39584 = n2829 & ~n39583;
  assign n39585 = ~n39582 & n39584;
  assign n39586 = ~n39240 & ~n39585;
  assign n39587 = ~pi174 & ~n39586;
  assign n39588 = ~n3890 & ~n39357;
  assign n39589 = n58822 & ~n39588;
  assign n39590 = pi174 & n39589;
  assign n39591 = ~pi193 & ~n39590;
  assign n39592 = ~n39587 & n39591;
  assign n39593 = pi180 & ~n39592;
  assign n39594 = ~n39579 & n39593;
  assign n39595 = ~n3890 & ~n38923;
  assign n39596 = ~n39581 & ~n39595;
  assign n39597 = ~pi174 & n39596;
  assign n39598 = n3890 & n60632;
  assign n39599 = ~pi51 & n39598;
  assign n39600 = n58822 & n3890;
  assign n39601 = pi174 & n60647;
  assign n39602 = ~n39540 & ~n39601;
  assign n39603 = ~n39597 & n39602;
  assign n39604 = ~pi180 & ~n39603;
  assign n39605 = ~pi299 & ~n39604;
  assign n39606 = ~n39594 & n39605;
  assign n39607 = ~n3906 & n39416;
  assign n39608 = pi152 & n60646;
  assign n39609 = ~pi152 & n39570;
  assign n39610 = pi51 & ~pi172;
  assign n39611 = ~n39609 & ~n39610;
  assign n39612 = ~pi152 & ~n39570;
  assign n39613 = pi152 & ~n60646;
  assign n39614 = ~n39612 & ~n39613;
  assign n39615 = ~n39610 & ~n39614;
  assign n39616 = ~n39608 & ~n39610;
  assign n39617 = ~n39609 & n39616;
  assign n39618 = ~n39608 & n39611;
  assign n39619 = ~pi216 & ~n60648;
  assign n39620 = n2852 & n39619;
  assign n39621 = ~n39607 & ~n39620;
  assign n39622 = n31084 & ~n39621;
  assign n39623 = pi152 & ~n39559;
  assign n39624 = ~n38923 & ~n39572;
  assign n39625 = ~pi152 & ~n39624;
  assign n39626 = pi172 & ~n39625;
  assign n39627 = ~n39623 & n39626;
  assign n39628 = pi152 & n39372;
  assign n39629 = ~pi152 & n39247;
  assign n39630 = ~pi172 & ~n39629;
  assign n39631 = ~n39628 & n39630;
  assign n39632 = ~n39627 & ~n39631;
  assign n39633 = pi152 & ~n39372;
  assign n39634 = ~pi152 & ~n39247;
  assign n39635 = ~pi172 & ~n39634;
  assign n39636 = ~n39633 & n39635;
  assign n39637 = pi152 & n39559;
  assign n39638 = ~pi152 & n39624;
  assign n39639 = pi172 & ~n39638;
  assign n39640 = ~n39637 & n39639;
  assign n39641 = pi216 & ~n39640;
  assign n39642 = ~n39636 & n39641;
  assign n39643 = pi216 & ~n39632;
  assign n39644 = n2852 & ~n39619;
  assign n39645 = n2852 & ~n60649;
  assign n39646 = ~n39619 & n39645;
  assign n39647 = ~n60649 & n39644;
  assign n39648 = ~n2852 & ~n39416;
  assign n39649 = n31099 & ~n39648;
  assign n39650 = ~n60650 & n39649;
  assign n39651 = ~n39622 & ~n39650;
  assign n39652 = ~n39606 & n39651;
  assign n39653 = pi232 & ~n39652;
  assign n39654 = n39557 & ~n39653;
  assign n39655 = ~pi232 & ~n39030;
  assign n39656 = ~pi39 & ~n39655;
  assign n39657 = ~pi38 & ~n39656;
  assign n39658 = ~n39654 & n39657;
  assign n39659 = pi299 & n39416;
  assign n39660 = ~pi174 & n39059;
  assign n39661 = ~pi299 & ~n39540;
  assign n39662 = ~n39660 & n39661;
  assign n39663 = pi232 & ~n39662;
  assign n39664 = ~n39659 & n39663;
  assign n39665 = pi38 & ~n39664;
  assign n39666 = ~pi100 & ~n39665;
  assign n39667 = ~n39658 & n39666;
  assign n39668 = ~n39550 & n39667;
  assign n39669 = pi100 & n39664;
  assign n39670 = n6311 & ~n39669;
  assign n39671 = ~n39668 & n39670;
  assign n39672 = n39286 & ~n39664;
  assign n39673 = pi140 & ~pi299;
  assign n39674 = ~n34323 & ~n39673;
  assign n39675 = n2681 & ~n39674;
  assign n39676 = pi87 & ~n39675;
  assign n39677 = n39412 & ~n39676;
  assign n39678 = ~n39672 & n39677;
  assign n39679 = ~n39671 & n39678;
  assign n39680 = ~pi232 & ~n39068;
  assign n39681 = ~pi39 & ~n39680;
  assign n39682 = n29572 & n39193;
  assign n39683 = n38922 & ~n39682;
  assign n39684 = ~pi299 & ~n39683;
  assign n39685 = n29532 & n39193;
  assign n39686 = n38922 & ~n39685;
  assign n39687 = pi299 & ~n39686;
  assign n39688 = ~n39684 & ~n39687;
  assign n39689 = ~pi232 & ~n39688;
  assign n39690 = pi39 & ~n39689;
  assign n39691 = ~n38922 & n39416;
  assign n39692 = ~n29532 & ~n39691;
  assign n39693 = n39215 & n39456;
  assign n39694 = pi152 & ~n39414;
  assign n39695 = ~n39218 & n39694;
  assign n39696 = n29532 & ~n39695;
  assign n39697 = ~pi152 & ~n39215;
  assign n39698 = pi152 & n39218;
  assign n39699 = ~n39414 & ~n39698;
  assign n39700 = ~n39697 & n39699;
  assign n39701 = n29532 & ~n39700;
  assign n39702 = ~n39693 & n39696;
  assign n39703 = n31099 & ~n60651;
  assign n39704 = ~n39194 & ~n39424;
  assign n39705 = ~pi152 & n39201;
  assign n39706 = ~n39704 & ~n39705;
  assign n39707 = ~pi172 & ~n39706;
  assign n39708 = ~pi152 & n39204;
  assign n39709 = pi152 & n39252;
  assign n39710 = pi172 & ~n39709;
  assign n39711 = ~n39708 & n39710;
  assign n39712 = n29532 & ~n39711;
  assign n39713 = n29532 & ~n39707;
  assign n39714 = ~n39711 & n39713;
  assign n39715 = ~n39707 & n39712;
  assign n39716 = n31084 & ~n60652;
  assign n39717 = ~n39703 & ~n39716;
  assign n39718 = ~n39692 & ~n39717;
  assign n39719 = ~n2680 & ~n38921;
  assign n39720 = ~n29572 & ~n39719;
  assign n39721 = ~n39251 & n39720;
  assign n39722 = n29572 & n39204;
  assign n39723 = ~n39721 & ~n39722;
  assign n39724 = ~pi174 & n39723;
  assign n39725 = ~n38918 & ~n39683;
  assign n39726 = pi174 & n39725;
  assign n39727 = ~pi180 & ~n39726;
  assign n39728 = ~n39724 & n39727;
  assign n39729 = n29572 & ~n39197;
  assign n39730 = ~n60487 & n39729;
  assign n39731 = ~n39721 & ~n39730;
  assign n39732 = ~pi174 & n39731;
  assign n39733 = ~pi51 & ~n39218;
  assign n39734 = n2680 & ~n39733;
  assign n39735 = ~n39683 & ~n39734;
  assign n39736 = pi174 & n39735;
  assign n39737 = pi180 & ~n39736;
  assign n39738 = ~n39732 & n39737;
  assign n39739 = ~n39728 & ~n39738;
  assign n39740 = ~pi174 & ~n39723;
  assign n39741 = pi174 & ~n39725;
  assign n39742 = ~pi180 & ~n39741;
  assign n39743 = ~n39740 & n39742;
  assign n39744 = ~pi174 & ~n39731;
  assign n39745 = pi174 & ~n39735;
  assign n39746 = pi180 & ~n39745;
  assign n39747 = ~n39744 & n39746;
  assign n39748 = pi193 & ~n39747;
  assign n39749 = ~n39743 & n39748;
  assign n39750 = pi193 & ~n39739;
  assign n39751 = ~pi51 & n39720;
  assign n39752 = n29572 & n39202;
  assign n39753 = ~n39751 & ~n39752;
  assign n39754 = pi180 & n39214;
  assign n39755 = ~pi174 & ~n39754;
  assign n39756 = n39753 & n39755;
  assign n39757 = pi180 & n39218;
  assign n39758 = pi174 & ~n39683;
  assign n39759 = ~n39757 & n39758;
  assign n39760 = ~pi193 & ~n39759;
  assign n39761 = ~n39756 & n39760;
  assign n39762 = ~pi299 & ~n39761;
  assign n39763 = ~n60653 & n39762;
  assign n39764 = ~n39718 & ~n39763;
  assign n39765 = pi232 & ~n39764;
  assign n39766 = n39690 & ~n39765;
  assign n39767 = ~n39681 & ~n39766;
  assign n39768 = ~pi145 & ~n39069;
  assign n39769 = ~n39296 & n39768;
  assign n39770 = ~n39050 & ~n39069;
  assign n39771 = pi145 & n39770;
  assign n39772 = ~pi51 & n39771;
  assign n39773 = ~pi174 & ~n39772;
  assign n39774 = ~n39769 & n39773;
  assign n39775 = ~pi145 & ~n39067;
  assign n39776 = ~n2680 & ~n39067;
  assign n39777 = ~n38923 & ~n39776;
  assign n39778 = ~n39001 & n39777;
  assign n39779 = ~n39775 & n39778;
  assign n39780 = pi174 & ~n39779;
  assign n39781 = ~pi193 & ~n39780;
  assign n39782 = ~n39774 & n39781;
  assign n39783 = n39019 & n60621;
  assign n39784 = ~n39069 & ~n39783;
  assign n39785 = ~pi145 & n39784;
  assign n39786 = ~pi174 & ~n39771;
  assign n39787 = ~n39785 & n39786;
  assign n39788 = n2599 & n39779;
  assign n39789 = ~n39069 & ~n39304;
  assign n39790 = pi174 & ~n39789;
  assign n39791 = ~n39788 & n39790;
  assign n39792 = pi193 & ~n39791;
  assign n39793 = ~n39787 & n39792;
  assign n39794 = n29581 & ~n39793;
  assign n39795 = ~n39782 & n39794;
  assign n39796 = ~n38918 & ~n39069;
  assign n39797 = ~pi174 & ~n39499;
  assign n39798 = pi145 & n38921;
  assign n39799 = ~n39797 & ~n39798;
  assign n39800 = n39796 & ~n39799;
  assign n39801 = ~n39069 & ~n39323;
  assign n39802 = pi174 & n39801;
  assign n39803 = ~n39800 & ~n39802;
  assign n39804 = ~pi193 & ~n39803;
  assign n39805 = pi145 & ~n39059;
  assign n39806 = ~pi145 & pi174;
  assign n39807 = ~n39321 & n39806;
  assign n39808 = ~n39805 & ~n39807;
  assign n39809 = ~n39797 & n39808;
  assign n39810 = pi193 & ~n39069;
  assign n39811 = ~n39809 & n39810;
  assign n39812 = n29601 & ~n39811;
  assign n39813 = ~n39804 & n39812;
  assign n39814 = ~n39795 & ~n39813;
  assign n39815 = n29912 & ~n39814;
  assign n39816 = ~n39767 & ~n39815;
  assign n39817 = ~pi38 & ~n39816;
  assign n39818 = ~n38964 & ~n39666;
  assign n39819 = ~pi152 & ~n39784;
  assign n39820 = pi152 & ~n39789;
  assign n39821 = pi172 & ~n39820;
  assign n39822 = ~n39819 & n39821;
  assign n39823 = ~pi152 & n39296;
  assign n39824 = ~n39068 & ~n39424;
  assign n39825 = ~pi172 & ~n39824;
  assign n39826 = ~n39823 & n39825;
  assign n39827 = ~n39822 & ~n39826;
  assign n39828 = ~pi197 & ~n39827;
  assign n39829 = ~pi152 & ~n39770;
  assign n39830 = ~n39062 & ~n39069;
  assign n39831 = pi172 & n39830;
  assign n39832 = ~pi172 & n39778;
  assign n39833 = pi152 & ~n39832;
  assign n39834 = pi172 & ~n39830;
  assign n39835 = ~pi172 & ~n39778;
  assign n39836 = ~n39834 & ~n39835;
  assign n39837 = pi152 & ~n39836;
  assign n39838 = ~n39831 & n39833;
  assign n39839 = ~pi172 & n38918;
  assign n39840 = pi197 & ~n39839;
  assign n39841 = ~n60654 & n39840;
  assign n39842 = ~n39829 & n39841;
  assign n39843 = pi299 & n29555;
  assign n39844 = ~n39842 & n39843;
  assign n39845 = ~n39828 & n39844;
  assign n39846 = ~n39069 & ~n39110;
  assign n39847 = ~pi152 & n39846;
  assign n39848 = ~n38918 & n39847;
  assign n39849 = pi152 & n39801;
  assign n39850 = ~pi172 & ~n39849;
  assign n39851 = ~n39848 & n39850;
  assign n39852 = ~n39069 & ~n39321;
  assign n39853 = pi152 & n39852;
  assign n39854 = pi172 & ~n39853;
  assign n39855 = ~n39847 & n39854;
  assign n39856 = ~pi197 & ~n39855;
  assign n39857 = ~n39851 & n39856;
  assign n39858 = pi299 & n29564;
  assign n39859 = pi152 & n39059;
  assign n39860 = ~n39069 & ~n39859;
  assign n39861 = pi172 & ~n39860;
  assign n39862 = ~pi172 & ~n39415;
  assign n39863 = ~n39070 & n39862;
  assign n39864 = pi197 & ~n39863;
  assign n39865 = pi197 & ~n39861;
  assign n39866 = ~n39863 & n39865;
  assign n39867 = ~n39861 & n39864;
  assign n39868 = n39858 & ~n60655;
  assign n39869 = ~n39861 & ~n39863;
  assign n39870 = pi197 & ~n39869;
  assign n39871 = ~n39839 & n39846;
  assign n39872 = ~pi152 & ~n39871;
  assign n39873 = pi172 & n39852;
  assign n39874 = ~pi172 & n39801;
  assign n39875 = pi152 & ~n39874;
  assign n39876 = ~n39873 & n39875;
  assign n39877 = ~n39872 & ~n39876;
  assign n39878 = ~pi197 & ~n39877;
  assign n39879 = ~n39870 & ~n39878;
  assign n39880 = n39858 & ~n39879;
  assign n39881 = ~n39857 & n39868;
  assign n39882 = ~n39845 & ~n60656;
  assign n39883 = n29912 & ~n39882;
  assign n39884 = ~n39818 & ~n39883;
  assign n39885 = ~pi38 & ~n39814;
  assign n39886 = n39882 & ~n39885;
  assign n39887 = n29912 & ~n39886;
  assign n39888 = ~pi38 & ~n39681;
  assign n39889 = ~n39766 & n39888;
  assign n39890 = ~n39818 & ~n39889;
  assign n39891 = ~n39887 & n39890;
  assign n39892 = ~n39817 & n39884;
  assign n39893 = ~n39282 & n39670;
  assign n39894 = n39283 & ~n39669;
  assign n39895 = ~n60657 & n60658;
  assign n39896 = n39287 & ~n39664;
  assign n39897 = ~n39412 & ~n39676;
  assign n39898 = ~n39896 & n39897;
  assign n39899 = ~n39895 & n39898;
  assign n39900 = n58992 & ~n39899;
  assign n39901 = ~n39679 & n39900;
  assign n39902 = ~n39423 & ~n39901;
  assign n39903 = ~pi189 & n39455;
  assign n39904 = pi189 & n39448;
  assign n39905 = ~n39903 & ~n39904;
  assign n39906 = pi178 & ~n39905;
  assign n39907 = pi189 & ~n39437;
  assign n39908 = ~pi189 & ~n39431;
  assign n39909 = ~pi178 & ~n39908;
  assign n39910 = ~n39907 & n39909;
  assign n39911 = ~n39906 & ~n39910;
  assign n39912 = pi181 & ~n39911;
  assign n39913 = pi189 & n39468;
  assign n39914 = ~pi189 & ~n39470;
  assign n39915 = pi178 & ~n39914;
  assign n39916 = ~n39913 & n39915;
  assign n39917 = ~pi189 & ~n39493;
  assign n39918 = pi189 & n39030;
  assign n39919 = ~pi178 & ~n39918;
  assign n39920 = ~n38918 & n39919;
  assign n39921 = ~n39917 & n39920;
  assign n39922 = ~pi181 & ~n39921;
  assign n39923 = n39493 & n39919;
  assign n39924 = n39922 & ~n39923;
  assign n39925 = ~n39916 & n39924;
  assign n39926 = n30114 & ~n39925;
  assign n39927 = ~n39912 & n39926;
  assign n39928 = ~pi153 & n39448;
  assign n39929 = pi153 & n39450;
  assign n39930 = pi157 & ~n39929;
  assign n39931 = ~n39928 & n39930;
  assign n39932 = ~pi153 & n39437;
  assign n39933 = pi153 & ~n60639;
  assign n39934 = ~pi157 & ~n39933;
  assign n39935 = ~n39932 & n39934;
  assign n39936 = ~n39931 & ~n39935;
  assign n39937 = pi166 & ~n39936;
  assign n39938 = pi157 & n39455;
  assign n39939 = ~pi157 & n39431;
  assign n39940 = pi153 & n38918;
  assign n39941 = ~pi166 & ~n39940;
  assign n39942 = ~n39939 & n39941;
  assign n39943 = ~n39938 & n39941;
  assign n39944 = ~n39939 & n39943;
  assign n39945 = ~n39938 & n39942;
  assign n39946 = ~n39937 & ~n60659;
  assign n39947 = n29502 & ~n39946;
  assign n39948 = pi166 & ~n39474;
  assign n39949 = ~pi166 & n39478;
  assign n39950 = pi153 & ~n39949;
  assign n39951 = ~n39948 & n39950;
  assign n39952 = pi166 & n39468;
  assign n39953 = ~pi166 & ~n39470;
  assign n39954 = ~pi153 & ~n39953;
  assign n39955 = ~n39952 & n39954;
  assign n39956 = ~n39951 & ~n39955;
  assign n39957 = pi157 & ~n39956;
  assign n39958 = ~pi166 & ~n39493;
  assign n39959 = pi166 & n39030;
  assign n39960 = ~pi157 & ~n39940;
  assign n39961 = ~n39959 & n39960;
  assign n39962 = ~n39958 & n39961;
  assign n39963 = ~n39957 & ~n39962;
  assign n39964 = n29424 & ~n39963;
  assign n39965 = ~pi189 & n39796;
  assign n39966 = n39450 & ~n39965;
  assign n39967 = pi178 & ~n39903;
  assign n39968 = ~n39966 & n39967;
  assign n39969 = pi189 & n60639;
  assign n39970 = ~n38918 & n39908;
  assign n39971 = ~n39969 & ~n39970;
  assign n39972 = ~pi178 & ~n39971;
  assign n39973 = pi181 & ~n39972;
  assign n39974 = ~n39968 & n39973;
  assign n39975 = pi189 & ~n39474;
  assign n39976 = ~pi189 & n39478;
  assign n39977 = pi178 & ~n39976;
  assign n39978 = ~n39975 & n39977;
  assign n39979 = n39922 & ~n39978;
  assign n39980 = n30168 & ~n39979;
  assign n39981 = ~n39974 & n39980;
  assign n39982 = ~n39964 & ~n39981;
  assign n39983 = ~n39947 & n39982;
  assign n39984 = ~n39927 & n39983;
  assign n39985 = pi232 & ~n39984;
  assign n39986 = n39656 & ~n39985;
  assign n39987 = ~pi126 & n38941;
  assign n39988 = pi126 & ~n38941;
  assign n39989 = ~n39987 & ~n39988;
  assign n39990 = ~n38937 & ~n39989;
  assign n39991 = ~pi189 & n39596;
  assign n39992 = pi189 & n60647;
  assign n39993 = ~pi182 & ~n39992;
  assign n39994 = ~n39991 & n39993;
  assign n39995 = ~n38918 & n39994;
  assign n39996 = pi189 & ~n39567;
  assign n39997 = ~pi189 & n39576;
  assign n39998 = pi182 & ~n39997;
  assign n39999 = ~n39996 & n39998;
  assign n40000 = ~n39995 & ~n39999;
  assign n40001 = n30168 & ~n40000;
  assign n40002 = ~pi189 & ~n39586;
  assign n40003 = pi189 & n39589;
  assign n40004 = pi182 & ~n40003;
  assign n40005 = ~n40002 & n40004;
  assign n40006 = ~n39994 & ~n40005;
  assign n40007 = n30114 & ~n40006;
  assign n40008 = pi166 & n39559;
  assign n40009 = ~pi166 & n39624;
  assign n40010 = pi153 & ~n40009;
  assign n40011 = ~n40008 & n40010;
  assign n40012 = pi166 & ~n39372;
  assign n40013 = ~pi166 & ~n39247;
  assign n40014 = ~pi153 & ~n40013;
  assign n40015 = ~n40012 & n40014;
  assign n40016 = ~n40011 & ~n40015;
  assign n40017 = pi166 & ~n39559;
  assign n40018 = ~pi166 & ~n39624;
  assign n40019 = pi153 & ~n40018;
  assign n40020 = ~n40017 & n40019;
  assign n40021 = pi166 & n39372;
  assign n40022 = n2801 & n30049;
  assign n40023 = ~pi166 & n39247;
  assign n40024 = ~pi153 & ~n40023;
  assign n40025 = ~n60660 & n40024;
  assign n40026 = pi160 & ~n40025;
  assign n40027 = ~n40020 & n40026;
  assign n40028 = pi160 & ~n40016;
  assign n40029 = pi216 & ~n60661;
  assign n40030 = ~pi166 & n39570;
  assign n40031 = pi166 & n60646;
  assign n40032 = pi51 & ~pi153;
  assign n40033 = ~n40031 & ~n40032;
  assign n40034 = ~pi166 & ~n39570;
  assign n40035 = pi166 & ~n60646;
  assign n40036 = ~n40034 & ~n40035;
  assign n40037 = ~n40032 & ~n40036;
  assign n40038 = ~n40030 & n40033;
  assign n40039 = ~pi216 & ~n60662;
  assign n40040 = n2852 & ~n40039;
  assign n40041 = n2852 & ~n40029;
  assign n40042 = ~n40039 & n40041;
  assign n40043 = ~n40029 & n40040;
  assign n40044 = ~pi51 & ~n39059;
  assign n40045 = ~n29998 & ~n38921;
  assign n40046 = ~pi51 & ~n40045;
  assign n40047 = ~n39940 & ~n40046;
  assign n40048 = ~n40044 & ~n40047;
  assign n40049 = ~pi160 & pi216;
  assign n40050 = n2852 & ~n40049;
  assign n40051 = n40048 & ~n40050;
  assign n40052 = pi299 & ~n40051;
  assign n40053 = ~n60663 & n40052;
  assign n40054 = ~n40007 & ~n40053;
  assign n40055 = ~n40001 & ~n40007;
  assign n40056 = ~n40053 & n40055;
  assign n40057 = ~n40001 & n40054;
  assign n40058 = pi232 & ~n60664;
  assign n40059 = n39557 & ~n40058;
  assign n40060 = n39990 & ~n40059;
  assign n40061 = ~n39986 & n40060;
  assign n40062 = ~n29998 & ~n39068;
  assign n40063 = ~pi166 & n39296;
  assign n40064 = ~n40062 & ~n40063;
  assign n40065 = ~pi153 & ~n40064;
  assign n40066 = ~pi166 & n39784;
  assign n40067 = pi166 & n39789;
  assign n40068 = pi153 & ~n40067;
  assign n40069 = ~n40066 & n40068;
  assign n40070 = ~pi157 & ~n40069;
  assign n40071 = ~pi166 & ~n39784;
  assign n40072 = pi166 & ~n39789;
  assign n40073 = pi153 & ~n40072;
  assign n40074 = ~n40071 & n40073;
  assign n40075 = ~pi153 & ~n40062;
  assign n40076 = ~n40063 & n40075;
  assign n40077 = ~n40074 & ~n40076;
  assign n40078 = ~pi157 & ~n40077;
  assign n40079 = ~n40065 & n40070;
  assign n40080 = pi166 & ~n39801;
  assign n40081 = pi51 & n29998;
  assign n40082 = ~n40080 & ~n40081;
  assign n40083 = ~pi153 & ~n40082;
  assign n40084 = ~pi166 & ~n39846;
  assign n40085 = pi153 & pi166;
  assign n40086 = ~n39852 & n40085;
  assign n40087 = pi157 & ~n40086;
  assign n40088 = ~n40084 & n40087;
  assign n40089 = ~n40083 & n40087;
  assign n40090 = ~n40084 & n40089;
  assign n40091 = ~n40083 & n40088;
  assign n40092 = n29424 & ~n60666;
  assign n40093 = ~n60665 & n40092;
  assign n40094 = ~n30128 & ~n39068;
  assign n40095 = ~pi189 & n39296;
  assign n40096 = ~n40094 & ~n40095;
  assign n40097 = ~pi178 & ~n40096;
  assign n40098 = pi189 & n39801;
  assign n40099 = pi178 & ~n39965;
  assign n40100 = ~pi189 & n39846;
  assign n40101 = pi178 & ~n40100;
  assign n40102 = ~n40099 & ~n40101;
  assign n40103 = ~n40098 & ~n40102;
  assign n40104 = ~pi181 & ~n40103;
  assign n40105 = ~n40097 & n40104;
  assign n40106 = ~n39050 & n39965;
  assign n40107 = pi189 & n39778;
  assign n40108 = ~pi178 & ~n40107;
  assign n40109 = ~n40106 & n40108;
  assign n40110 = pi189 & n39070;
  assign n40111 = n40099 & ~n40110;
  assign n40112 = pi181 & ~n40111;
  assign n40113 = ~n40109 & n40112;
  assign n40114 = n30114 & ~n40113;
  assign n40115 = ~n40105 & n40114;
  assign n40116 = ~pi189 & n39784;
  assign n40117 = pi189 & n39789;
  assign n40118 = ~pi178 & ~n40117;
  assign n40119 = ~n40116 & n40118;
  assign n40120 = pi189 & n39852;
  assign n40121 = n40101 & ~n40120;
  assign n40122 = ~pi181 & ~n40121;
  assign n40123 = ~n40119 & n40122;
  assign n40124 = ~pi189 & ~n39050;
  assign n40125 = pi189 & ~n39062;
  assign n40126 = ~pi178 & ~n40125;
  assign n40127 = ~n40124 & n40126;
  assign n40128 = pi178 & n30125;
  assign n40129 = n39058 & n40128;
  assign n40130 = pi181 & ~n40129;
  assign n40131 = ~n39069 & n40130;
  assign n40132 = ~n40127 & n40131;
  assign n40133 = n30168 & ~n40132;
  assign n40134 = ~n40123 & n40133;
  assign n40135 = ~pi166 & ~n39770;
  assign n40136 = ~n39830 & n40085;
  assign n40137 = pi166 & ~n39778;
  assign n40138 = ~n40081 & ~n40137;
  assign n40139 = ~pi153 & ~n40138;
  assign n40140 = ~pi157 & ~n40139;
  assign n40141 = ~pi157 & ~n40136;
  assign n40142 = ~n40139 & n40141;
  assign n40143 = ~n40136 & n40140;
  assign n40144 = ~n40135 & n60667;
  assign n40145 = ~pi153 & ~n40048;
  assign n40146 = ~n39070 & n40145;
  assign n40147 = pi166 & n39059;
  assign n40148 = n30049 & n39058;
  assign n40149 = ~n39069 & ~n60668;
  assign n40150 = pi153 & ~n40149;
  assign n40151 = pi157 & ~n40150;
  assign n40152 = ~n40146 & n40151;
  assign n40153 = n29502 & ~n40152;
  assign n40154 = ~n40144 & n40153;
  assign n40155 = ~n40134 & ~n40154;
  assign n40156 = ~n40115 & n40155;
  assign n40157 = ~n40093 & n40155;
  assign n40158 = ~n40115 & n40157;
  assign n40159 = ~n40093 & n40156;
  assign n40160 = pi232 & ~n60669;
  assign n40161 = n39681 & ~n40160;
  assign n40162 = ~pi166 & ~n39215;
  assign n40163 = pi166 & n39218;
  assign n40164 = pi160 & ~n39940;
  assign n40165 = ~n40163 & n40164;
  assign n40166 = ~pi166 & n39215;
  assign n40167 = pi166 & ~n39218;
  assign n40168 = ~n40166 & ~n40167;
  assign n40169 = n40164 & ~n40168;
  assign n40170 = ~n40162 & n40165;
  assign n40171 = ~pi166 & n39201;
  assign n40172 = ~n29998 & ~n39194;
  assign n40173 = ~pi153 & ~n40172;
  assign n40174 = ~n40171 & n40173;
  assign n40175 = ~pi166 & ~n39204;
  assign n40176 = pi166 & ~n39252;
  assign n40177 = pi153 & ~n40176;
  assign n40178 = ~n40175 & n40177;
  assign n40179 = ~pi160 & ~n40178;
  assign n40180 = ~n40171 & ~n40172;
  assign n40181 = ~pi153 & ~n40180;
  assign n40182 = ~pi166 & n39204;
  assign n40183 = pi166 & n39252;
  assign n40184 = pi153 & ~n40183;
  assign n40185 = ~n40182 & n40184;
  assign n40186 = ~n40181 & ~n40185;
  assign n40187 = ~pi160 & ~n40186;
  assign n40188 = ~n40174 & n40179;
  assign n40189 = n29532 & ~n60671;
  assign n40190 = n29532 & ~n60670;
  assign n40191 = ~n60671 & n40190;
  assign n40192 = ~n60670 & n40189;
  assign n40193 = ~n29532 & ~n40047;
  assign n40194 = pi299 & ~n40193;
  assign n40195 = ~n60672 & n40194;
  assign n40196 = ~pi189 & ~n39723;
  assign n40197 = pi189 & ~n39725;
  assign n40198 = ~pi182 & ~n40197;
  assign n40199 = ~n40196 & n40198;
  assign n40200 = ~pi189 & ~n39731;
  assign n40201 = pi189 & ~n39735;
  assign n40202 = pi182 & ~n40201;
  assign n40203 = ~n40200 & n40202;
  assign n40204 = ~n40199 & ~n40203;
  assign n40205 = n30168 & ~n40204;
  assign n40206 = pi182 & n39218;
  assign n40207 = pi189 & ~n39683;
  assign n40208 = ~n40206 & n40207;
  assign n40209 = pi182 & n39214;
  assign n40210 = ~pi189 & ~n40209;
  assign n40211 = n39753 & n40210;
  assign n40212 = ~n40208 & ~n40211;
  assign n40213 = n30114 & ~n40212;
  assign n40214 = ~n40205 & ~n40213;
  assign n40215 = ~n40195 & n40214;
  assign n40216 = pi232 & ~n40215;
  assign n40217 = n39690 & ~n40216;
  assign n40218 = ~n39990 & ~n40217;
  assign n40219 = ~n40161 & n40218;
  assign n40220 = n2636 & ~n40219;
  assign n40221 = ~n40061 & n40220;
  assign n40222 = pi299 & ~n40048;
  assign n40223 = ~pi189 & n39059;
  assign n40224 = n30128 & n39058;
  assign n40225 = pi175 & n38918;
  assign n40226 = ~pi299 & ~n40225;
  assign n40227 = ~n60673 & n40226;
  assign n40228 = pi232 & ~n40227;
  assign n40229 = ~n40222 & n40228;
  assign n40230 = ~n2636 & n40229;
  assign n40231 = ~n2636 & n38922;
  assign n40232 = ~n39990 & n40231;
  assign n40233 = n6311 & ~n40232;
  assign n40234 = n38922 & ~n39990;
  assign n40235 = ~n40229 & ~n40234;
  assign n40236 = ~n2636 & ~n40235;
  assign n40237 = n6311 & ~n40236;
  assign n40238 = ~n40230 & n40233;
  assign n40239 = ~n40221 & n60674;
  assign n40240 = n39286 & ~n40229;
  assign n40241 = ~pi150 & pi299;
  assign n40242 = ~pi185 & ~pi299;
  assign n40243 = ~n40241 & ~n40242;
  assign n40244 = n2681 & n40243;
  assign n40245 = pi87 & ~n40244;
  assign n40246 = ~n40240 & ~n40245;
  assign n40247 = n38944 & ~n39990;
  assign n40248 = ~n40246 & ~n40247;
  assign n40249 = n58992 & ~n40248;
  assign n40250 = ~n40239 & n40249;
  assign n40251 = pi232 & ~n40044;
  assign n40252 = n39990 & ~n40251;
  assign n40253 = ~pi232 & ~n38922;
  assign n40254 = ~n40047 & ~n40253;
  assign n40255 = ~n40252 & n40254;
  assign n40256 = ~pi87 & ~n40255;
  assign n40257 = pi87 & ~n30744;
  assign n40258 = ~n58992 & ~n40257;
  assign n40259 = ~n40256 & n40258;
  assign n40260 = n39990 & n40044;
  assign n40261 = pi232 & ~n40260;
  assign n40262 = ~n40234 & ~n40261;
  assign n40263 = ~pi87 & ~n40047;
  assign n40264 = ~n40262 & n40263;
  assign n40265 = pi87 & n30744;
  assign n40266 = ~n58992 & ~n40265;
  assign n40267 = ~n40264 & n40266;
  assign n40268 = ~n40239 & ~n40248;
  assign n40269 = n58992 & ~n40268;
  assign n40270 = ~n40267 & ~n40269;
  assign n40271 = ~n40250 & ~n40259;
  assign n40272 = n3213 & ~n32496;
  assign n40273 = n32476 & ~n40272;
  assign n40274 = n36436 & ~n40273;
  assign n40275 = ~pi94 & n6317;
  assign n40276 = n2539 & n40275;
  assign n40277 = n2568 & n5152;
  assign n40278 = n37084 & n60676;
  assign n40279 = n2727 & n60165;
  assign n40280 = n58799 & n40279;
  assign n40281 = n40278 & n40280;
  assign n40282 = n32496 & n40281;
  assign n40283 = ~pi110 & ~n40278;
  assign n40284 = ~pi47 & ~n32496;
  assign n40285 = n40279 & n40284;
  assign n40286 = ~n40283 & n40285;
  assign n40287 = n36397 & n40286;
  assign n40288 = ~n40282 & ~n40287;
  assign n40289 = ~n3213 & ~n6416;
  assign n40290 = ~pi47 & n40279;
  assign n40291 = ~n40283 & n40290;
  assign n40292 = n36397 & n40291;
  assign n40293 = n2707 & ~n40292;
  assign n40294 = ~n2707 & ~n40281;
  assign n40295 = ~n2682 & ~n6416;
  assign n40296 = ~n40294 & n40295;
  assign n40297 = ~n40293 & n40296;
  assign n40298 = n2682 & ~n6416;
  assign n40299 = n40292 & n40298;
  assign n40300 = ~n40297 & ~n40299;
  assign n40301 = ~n3213 & ~n40300;
  assign n40302 = ~n32496 & ~n40292;
  assign n40303 = n32496 & ~n40281;
  assign n40304 = n40289 & ~n40303;
  assign n40305 = ~n40302 & n40304;
  assign n40306 = ~n40288 & n40289;
  assign n40307 = ~n40274 & ~n60677;
  assign po262 = n60562 & ~n40307;
  assign n40309 = pi51 & ~pi151;
  assign n40310 = ~n30617 & ~n38918;
  assign n40311 = ~n40309 & ~n40310;
  assign n40312 = n38923 & n40311;
  assign n40313 = pi232 & n40312;
  assign n40314 = ~pi132 & n39987;
  assign n40315 = pi132 & ~n39987;
  assign n40316 = ~n40314 & ~n40315;
  assign n40317 = ~n38936 & ~n40316;
  assign n40318 = n38922 & ~n40317;
  assign n40319 = ~n40313 & ~n40318;
  assign n40320 = ~pi87 & ~n40319;
  assign n40321 = pi164 & n39420;
  assign n40322 = ~n58992 & ~n40321;
  assign n40323 = ~n40320 & n40322;
  assign n40324 = pi299 & ~n40312;
  assign n40325 = pi190 & n39059;
  assign n40326 = pi173 & n38918;
  assign n40327 = ~pi299 & ~n40326;
  assign n40328 = ~n40325 & n40327;
  assign n40329 = pi232 & ~n40328;
  assign n40330 = ~n40324 & n40329;
  assign n40331 = ~n2636 & n40330;
  assign n40332 = n6311 & ~n40331;
  assign n40333 = ~pi168 & ~n39559;
  assign n40334 = pi168 & ~n39624;
  assign n40335 = pi151 & ~n40334;
  assign n40336 = ~n40333 & n40335;
  assign n40337 = ~pi168 & n39372;
  assign n40338 = pi168 & n39247;
  assign n40339 = ~pi151 & ~n40338;
  assign n40340 = ~n40337 & n40339;
  assign n40341 = pi149 & ~n40340;
  assign n40342 = pi149 & ~n40336;
  assign n40343 = ~n40340 & n40342;
  assign n40344 = ~n40336 & n40341;
  assign n40345 = pi216 & ~n60678;
  assign n40346 = pi168 & n39570;
  assign n40347 = ~pi168 & n60646;
  assign n40348 = ~n40309 & ~n40347;
  assign n40349 = pi168 & ~n39570;
  assign n40350 = ~pi168 & ~n60646;
  assign n40351 = ~n40349 & ~n40350;
  assign n40352 = ~n40309 & ~n40351;
  assign n40353 = ~n40346 & n40348;
  assign n40354 = ~pi216 & ~n60679;
  assign n40355 = n2852 & ~n40354;
  assign n40356 = n2852 & ~n40345;
  assign n40357 = ~n40354 & n40356;
  assign n40358 = ~n40345 & n40355;
  assign n40359 = ~pi149 & pi216;
  assign n40360 = n2852 & ~n40359;
  assign n40361 = n40312 & ~n40360;
  assign n40362 = pi299 & ~n40361;
  assign n40363 = ~n60680 & n40362;
  assign n40364 = pi190 & ~pi299;
  assign n40365 = pi183 & ~n39586;
  assign n40366 = ~pi183 & ~n39581;
  assign n40367 = ~pi173 & ~n40366;
  assign n40368 = ~n40365 & n40367;
  assign n40369 = ~pi183 & n39595;
  assign n40370 = ~pi183 & ~n39571;
  assign n40371 = pi173 & ~n39576;
  assign n40372 = ~n40370 & n40371;
  assign n40373 = ~n40369 & ~n40372;
  assign n40374 = ~n40368 & n40373;
  assign n40375 = n40364 & ~n40374;
  assign n40376 = pi183 & n39566;
  assign n40377 = ~pi183 & n60647;
  assign n40378 = ~n38918 & ~n40377;
  assign n40379 = ~n40376 & n40378;
  assign n40380 = pi183 & n39567;
  assign n40381 = ~pi183 & ~n38918;
  assign n40382 = ~n60647 & n40381;
  assign n40383 = pi173 & ~n40382;
  assign n40384 = ~n40380 & n40383;
  assign n40385 = pi173 & ~n40379;
  assign n40386 = ~pi183 & ~n3890;
  assign n40387 = ~pi173 & ~n40386;
  assign n40388 = n39589 & n40387;
  assign n40389 = ~pi190 & ~pi299;
  assign n40390 = ~n40388 & n40389;
  assign n40391 = ~n60681 & n40390;
  assign n40392 = ~n40375 & ~n40391;
  assign n40393 = ~n40363 & n40392;
  assign n40394 = pi232 & ~n40393;
  assign n40395 = n39557 & ~n40394;
  assign n40396 = ~pi232 & n39044;
  assign n40397 = ~pi151 & ~n39021;
  assign n40398 = pi151 & n39031;
  assign n40399 = ~pi168 & ~n40398;
  assign n40400 = ~pi168 & ~n40397;
  assign n40401 = ~n40398 & n40400;
  assign n40402 = ~n40397 & n40399;
  assign n40403 = pi168 & ~n40309;
  assign n40404 = ~n39009 & n40403;
  assign n40405 = n2680 & ~n40404;
  assign n40406 = ~n60682 & n40405;
  assign n40407 = ~n2680 & ~n39044;
  assign n40408 = pi160 & ~n40407;
  assign n40409 = ~n40406 & n40408;
  assign n40410 = ~n2680 & n39044;
  assign n40411 = n39053 & ~n40410;
  assign n40412 = ~pi168 & ~n40411;
  assign n40413 = pi168 & ~n60641;
  assign n40414 = ~n40407 & n40413;
  assign n40415 = pi151 & ~n40414;
  assign n40416 = ~n40412 & n40415;
  assign n40417 = ~n30617 & n39044;
  assign n40418 = pi168 & n39073;
  assign n40419 = ~pi151 & ~n40418;
  assign n40420 = ~n40417 & n40419;
  assign n40421 = ~pi160 & ~n40420;
  assign n40422 = ~n40416 & n40421;
  assign n40423 = pi299 & ~n40422;
  assign n40424 = ~pi168 & n40411;
  assign n40425 = ~n60641 & ~n40407;
  assign n40426 = pi168 & ~n40425;
  assign n40427 = pi151 & ~n40426;
  assign n40428 = ~n40424 & n40427;
  assign n40429 = ~n40417 & ~n40418;
  assign n40430 = ~pi151 & ~n40429;
  assign n40431 = ~pi160 & ~n40430;
  assign n40432 = ~n40428 & n40431;
  assign n40433 = ~n60682 & ~n40404;
  assign n40434 = n2680 & ~n40433;
  assign n40435 = pi160 & ~n40410;
  assign n40436 = ~n40434 & n40435;
  assign n40437 = ~n40432 & ~n40436;
  assign n40438 = pi299 & ~n40437;
  assign n40439 = ~n40409 & n40423;
  assign n40440 = pi182 & ~n40407;
  assign n40441 = ~n39022 & n40440;
  assign n40442 = ~pi182 & n39044;
  assign n40443 = ~pi173 & ~n40442;
  assign n40444 = ~n40441 & n40443;
  assign n40445 = ~n39032 & ~n40410;
  assign n40446 = pi182 & ~n40445;
  assign n40447 = ~pi182 & ~n40411;
  assign n40448 = pi173 & ~n40447;
  assign n40449 = ~n40446 & n40448;
  assign n40450 = ~n40444 & ~n40449;
  assign n40451 = n40389 & ~n40450;
  assign n40452 = pi182 & n38986;
  assign n40453 = n39008 & ~n40452;
  assign n40454 = pi51 & ~pi173;
  assign n40455 = n2680 & ~n40454;
  assign n40456 = ~n40453 & n40455;
  assign n40457 = n40364 & ~n40456;
  assign n40458 = ~n40410 & n40457;
  assign n40459 = pi232 & ~n40458;
  assign n40460 = ~n40451 & n40459;
  assign n40461 = ~n60683 & n40459;
  assign n40462 = ~n40451 & n40461;
  assign n40463 = ~n60683 & n40460;
  assign n40464 = ~n40396 & ~n60684;
  assign n40465 = ~pi39 & ~n40464;
  assign n40466 = ~n40395 & ~n40465;
  assign n40467 = n2636 & ~n40466;
  assign n40468 = n40332 & ~n40467;
  assign n40469 = n39286 & ~n40330;
  assign n40470 = pi87 & ~n30968;
  assign n40471 = n40317 & ~n40470;
  assign n40472 = ~n40469 & n40471;
  assign n40473 = ~n40468 & n40472;
  assign n40474 = ~pi183 & ~n39723;
  assign n40475 = pi183 & ~n39731;
  assign n40476 = pi173 & ~n40475;
  assign n40477 = ~n40474 & n40476;
  assign n40478 = pi183 & n39214;
  assign n40479 = ~pi173 & ~n40478;
  assign n40480 = n39753 & n40479;
  assign n40481 = ~n40477 & ~n40480;
  assign n40482 = n40364 & ~n40481;
  assign n40483 = ~n38922 & n40324;
  assign n40484 = ~n60188 & ~n40483;
  assign n40485 = pi168 & ~n39204;
  assign n40486 = ~pi168 & ~n39252;
  assign n40487 = pi151 & ~n40486;
  assign n40488 = ~n40485 & n40487;
  assign n40489 = pi168 & n39201;
  assign n40490 = ~n30617 & ~n39194;
  assign n40491 = ~pi151 & ~n40490;
  assign n40492 = ~n40489 & n40491;
  assign n40493 = ~pi149 & ~n40492;
  assign n40494 = ~n40488 & n40493;
  assign n40495 = ~n39559 & ~n40309;
  assign n40496 = ~n39202 & ~n40495;
  assign n40497 = pi168 & ~n40496;
  assign n40498 = ~n39218 & ~n40311;
  assign n40499 = ~pi168 & ~n40498;
  assign n40500 = pi149 & ~n40499;
  assign n40501 = ~n40497 & n40500;
  assign n40502 = n29532 & ~n40501;
  assign n40503 = n29532 & ~n40494;
  assign n40504 = ~n40501 & n40503;
  assign n40505 = ~n40494 & n40502;
  assign n40506 = ~n40484 & ~n60685;
  assign n40507 = pi183 & n39218;
  assign n40508 = ~n40326 & n40389;
  assign n40509 = ~n39683 & n40508;
  assign n40510 = ~n40507 & n40509;
  assign n40511 = ~n40506 & ~n40510;
  assign n40512 = ~n40482 & ~n40510;
  assign n40513 = ~n40506 & n40512;
  assign n40514 = ~n40482 & n40511;
  assign n40515 = pi232 & ~n60686;
  assign n40516 = ~n39689 & ~n40515;
  assign n40517 = pi39 & ~n40516;
  assign n40518 = pi151 & n39321;
  assign n40519 = ~pi151 & ~n39067;
  assign n40520 = ~pi168 & ~n40519;
  assign n40521 = ~n40518 & n40520;
  assign n40522 = ~pi151 & n38918;
  assign n40523 = pi168 & ~n40522;
  assign n40524 = ~n39110 & n40523;
  assign n40525 = ~n40521 & ~n40524;
  assign n40526 = ~pi160 & ~n39776;
  assign n40527 = ~n40525 & n40526;
  assign n40528 = ~pi151 & ~n40312;
  assign n40529 = ~n39777 & n40528;
  assign n40530 = ~pi168 & n39059;
  assign n40531 = ~n39776 & ~n40530;
  assign n40532 = pi151 & ~n40531;
  assign n40533 = pi160 & ~n40532;
  assign n40534 = ~n40529 & n40533;
  assign n40535 = pi299 & ~n40534;
  assign n40536 = ~n40527 & n40535;
  assign n40537 = ~pi182 & n39110;
  assign n40538 = ~n39776 & ~n40454;
  assign n40539 = ~n40537 & n40538;
  assign n40540 = n40364 & ~n40539;
  assign n40541 = pi182 & n39777;
  assign n40542 = ~n39067 & n40508;
  assign n40543 = ~n40541 & n40542;
  assign n40544 = pi232 & ~n40543;
  assign n40545 = ~n40540 & n40544;
  assign n40546 = ~n40536 & n40545;
  assign n40547 = ~pi232 & n39067;
  assign n40548 = ~pi39 & ~n40547;
  assign n40549 = ~n40546 & n40548;
  assign n40550 = n2636 & ~n40549;
  assign n40551 = ~n40517 & n40550;
  assign n40552 = n6311 & ~n40231;
  assign n40553 = ~n40231 & n40332;
  assign n40554 = ~n40331 & n40552;
  assign n40555 = ~n40551 & n60687;
  assign n40556 = n39287 & ~n40330;
  assign n40557 = ~n40317 & ~n40470;
  assign n40558 = ~n40556 & n40557;
  assign n40559 = ~n40555 & n40558;
  assign n40560 = n58992 & ~n40559;
  assign n40561 = ~n40473 & n40560;
  assign n40562 = ~n40323 & ~n40561;
  assign n40563 = n2446 & n58783;
  assign n40564 = ~pi102 & ~pi104;
  assign n40565 = ~pi111 & n40564;
  assign n40566 = ~pi45 & pi49;
  assign n40567 = n40565 & n40566;
  assign n40568 = n40563 & n40567;
  assign n40569 = n6327 & n40568;
  assign n40570 = n37071 & n40569;
  assign n40571 = n60478 & n40570;
  assign n40572 = ~n31412 & ~n40571;
  assign n40573 = n58797 & n6343;
  assign n40574 = n6343 & n40570;
  assign n40575 = n58797 & n40574;
  assign n40576 = n40570 & n40573;
  assign n40577 = n58818 & n35635;
  assign n40578 = n60688 & n40577;
  assign n40579 = n32496 & n38875;
  assign n40580 = ~n40578 & ~n40579;
  assign n40581 = n37798 & ~n40580;
  assign n40582 = ~n40572 & n40581;
  assign n40583 = ~n35649 & ~n40578;
  assign n40584 = pi252 & n37798;
  assign n40585 = ~n40572 & n40584;
  assign n40586 = n2793 & n40578;
  assign n40587 = pi1093 & ~n40586;
  assign n40588 = n2757 & ~n40587;
  assign n40589 = ~pi252 & n40578;
  assign n40590 = ~n40588 & ~n40589;
  assign n40591 = ~n40585 & n40590;
  assign n40592 = ~n40585 & ~n40588;
  assign n40593 = n35649 & ~n40592;
  assign n40594 = ~n40578 & ~n40593;
  assign n40595 = ~n40583 & ~n40591;
  assign n40596 = n32496 & n60689;
  assign n40597 = ~n32496 & ~n40578;
  assign n40598 = n60562 & ~n40597;
  assign n40599 = ~n40596 & n40598;
  assign n40600 = n60562 & n40582;
  assign n40601 = n60070 & n37126;
  assign n40602 = ~n4437 & ~n40601;
  assign n40603 = pi129 & n59171;
  assign n40604 = pi38 & ~n40603;
  assign n40605 = ~n6315 & ~n31488;
  assign n40606 = n31414 & ~n31447;
  assign n40607 = n2470 & ~n40606;
  assign n40608 = n31459 & ~n40607;
  assign n40609 = n28339 & ~n40608;
  assign n40610 = n28337 & ~n40609;
  assign n40611 = n28335 & ~n40610;
  assign n40612 = ~n28333 & ~n40611;
  assign n40613 = ~pi86 & ~n40612;
  assign n40614 = n28411 & ~n40613;
  assign n40615 = pi250 & ~n2682;
  assign n40616 = pi252 & n32496;
  assign n40617 = pi250 & n40616;
  assign n40618 = n37130 & n40615;
  assign n40619 = ~pi127 & ~n60691;
  assign n40620 = po740 & n60691;
  assign n40621 = ~n40619 & ~n40620;
  assign n40622 = n31412 & n40621;
  assign n40623 = ~pi97 & ~n40622;
  assign n40624 = ~n40614 & n40623;
  assign n40625 = ~n28628 & ~n40624;
  assign n40626 = ~pi108 & ~n40625;
  assign n40627 = n31410 & ~n40626;
  assign n40628 = n28449 & ~n40627;
  assign n40629 = ~n28447 & ~n40628;
  assign n40630 = n2540 & ~n40629;
  assign n40631 = ~pi97 & ~n40614;
  assign n40632 = ~n28628 & ~n40631;
  assign n40633 = ~pi108 & ~n40632;
  assign n40634 = n31410 & ~n40633;
  assign n40635 = n28449 & ~n40634;
  assign n40636 = ~n28447 & ~n40635;
  assign n40637 = n2540 & ~n40636;
  assign n40638 = n60541 & ~n40637;
  assign n40639 = po740 & n40638;
  assign n40640 = n31413 & ~n40614;
  assign n40641 = ~n28628 & ~n40640;
  assign n40642 = ~pi108 & ~n40641;
  assign n40643 = n31410 & ~n40642;
  assign n40644 = n28449 & ~n40643;
  assign n40645 = ~n28447 & ~n40644;
  assign n40646 = n2540 & ~n40645;
  assign n40647 = n60541 & ~n40646;
  assign n40648 = ~po740 & n40647;
  assign n40649 = n60691 & ~n40648;
  assign n40650 = n60691 & ~n40639;
  assign n40651 = ~n40648 & n40650;
  assign n40652 = ~n40639 & n40649;
  assign n40653 = ~pi127 & n40638;
  assign n40654 = pi127 & n40647;
  assign n40655 = ~n60691 & ~n40654;
  assign n40656 = ~n60691 & ~n40653;
  assign n40657 = ~n40654 & n40656;
  assign n40658 = ~n40653 & n40655;
  assign n40659 = ~n60692 & ~n60693;
  assign n40660 = n60541 & ~n40630;
  assign n40661 = n37380 & ~n60694;
  assign n40662 = n37379 & ~n40661;
  assign n40663 = n2592 & ~n40662;
  assign n40664 = n37377 & ~n40663;
  assign n40665 = ~pi70 & ~n40664;
  assign n40666 = ~n28320 & ~n40665;
  assign n40667 = ~pi51 & ~n40666;
  assign n40668 = n2604 & ~n40667;
  assign n40669 = n31408 & ~n40668;
  assign n40670 = ~n28318 & ~n40669;
  assign n40671 = n2620 & ~n40670;
  assign n40672 = n40605 & ~n40671;
  assign n40673 = ~pi95 & ~n40672;
  assign n40674 = ~pi39 & pi129;
  assign n40675 = ~n31400 & n40674;
  assign n40676 = ~n40673 & n40675;
  assign n40677 = pi39 & n37126;
  assign n40678 = ~pi38 & ~n40677;
  assign n40679 = ~n40676 & n40678;
  assign n40680 = ~n40604 & ~n40679;
  assign n40681 = n6305 & ~n40680;
  assign n40682 = ~n58815 & ~n30890;
  assign n40683 = n37126 & ~n40682;
  assign n40684 = ~n6305 & ~n40683;
  assign n40685 = ~pi75 & ~n40684;
  assign n40686 = ~n40681 & n40685;
  assign n40687 = pi129 & n28302;
  assign n40688 = pi75 & n40687;
  assign n40689 = ~pi92 & ~n40688;
  assign n40690 = ~n40686 & n40689;
  assign n40691 = pi92 & ~pi129;
  assign n40692 = n35283 & ~n40691;
  assign n40693 = ~n40690 & n40692;
  assign n40694 = pi54 & n60203;
  assign n40695 = n37126 & n40694;
  assign n40696 = ~pi74 & ~n40695;
  assign n40697 = ~n40693 & n40696;
  assign n40698 = n31593 & n40687;
  assign n40699 = pi74 & ~n40698;
  assign n40700 = ~pi55 & ~n40699;
  assign n40701 = ~n40697 & n40700;
  assign n40702 = pi55 & n6308;
  assign n40703 = n40687 & n40702;
  assign n40704 = ~n40701 & ~n40703;
  assign n40705 = ~pi56 & ~n40704;
  assign n40706 = pi56 & ~pi62;
  assign n40707 = ~pi56 & pi62;
  assign n40708 = ~n40706 & ~n40707;
  assign n40709 = ~n40705 & n40708;
  assign n40710 = ~n40602 & ~n40709;
  assign n40711 = n4438 & ~n40710;
  assign n40712 = n4437 & n40601;
  assign n40713 = n28292 & n37126;
  assign n40714 = ~n4438 & ~n60695;
  assign n40715 = ~n28282 & ~n40714;
  assign po284 = ~n40711 & n40715;
  assign n40717 = n2621 & n60562;
  assign n40718 = n59138 & n40717;
  assign n40719 = n60165 & n60562;
  assign n40720 = n58784 & n40563;
  assign n40721 = n2447 & n40720;
  assign n40722 = ~pi69 & n40721;
  assign n40723 = n6320 & n40722;
  assign n40724 = ~pi82 & ~pi109;
  assign n40725 = pi111 & n40724;
  assign n40726 = n58799 & n40725;
  assign n40727 = n58790 & n58799;
  assign n40728 = n40725 & n40727;
  assign n40729 = n58790 & n40725;
  assign n40730 = n58799 & n40729;
  assign n40731 = n58790 & n40726;
  assign n40732 = n40723 & n60697;
  assign n40733 = n28348 & n40732;
  assign n40734 = pi314 & n40733;
  assign n40735 = n32497 & n36413;
  assign n40736 = ~n40734 & ~n40735;
  assign po268 = n60696 & ~n40736;
  assign n40738 = ~pi70 & n38562;
  assign n40739 = ~n28320 & ~n31479;
  assign n40740 = ~n40738 & n40739;
  assign n40741 = ~pi51 & ~n40740;
  assign n40742 = n2604 & ~n40741;
  assign n40743 = n31408 & ~n40742;
  assign n40744 = ~n28318 & ~n40743;
  assign n40745 = n2620 & ~n40744;
  assign n40746 = n40605 & ~n40745;
  assign n40747 = ~pi95 & ~n40746;
  assign n40748 = ~n31400 & ~n40747;
  assign n40749 = ~pi39 & ~n40748;
  assign n40750 = ~n37419 & ~n40749;
  assign n40751 = ~pi38 & ~n40750;
  assign n40752 = n31399 & ~n40751;
  assign n40753 = n28549 & ~n28564;
  assign n40754 = n31664 & n37123;
  assign n40755 = ~pi87 & ~n60698;
  assign n40756 = ~n40752 & n40755;
  assign n40757 = n31561 & ~n40756;
  assign n40758 = ~pi250 & n40616;
  assign n40759 = n32496 & n36416;
  assign n40760 = ~pi129 & ~n60699;
  assign n40761 = po740 & n60699;
  assign n40762 = n37226 & ~n40761;
  assign n40763 = ~n40760 & n40762;
  assign n40764 = n58822 & n40763;
  assign n40765 = n2438 & ~n40764;
  assign n40766 = ~n40757 & n40765;
  assign n40767 = ~n28307 & ~n28586;
  assign n40768 = ~n40766 & n40767;
  assign n40769 = n31567 & ~n40768;
  assign n40770 = n37375 & ~n40769;
  assign n40771 = ~pi56 & ~n40770;
  assign n40772 = ~n31570 & ~n40771;
  assign n40773 = ~pi62 & ~n40772;
  assign n40774 = ~n31575 & ~n40773;
  assign n40775 = n4438 & ~n40774;
  assign po286 = n28295 & ~n40775;
  assign n40777 = ~pi51 & ~n39688;
  assign n40778 = ~pi232 & ~n40777;
  assign n40779 = n25479 & ~n40778;
  assign n40780 = ~pi51 & ~n39202;
  assign n40781 = ~n39213 & n40780;
  assign n40782 = pi169 & ~n40781;
  assign n40783 = pi162 & n29532;
  assign n40784 = ~pi169 & ~n39733;
  assign n40785 = n40783 & ~n40784;
  assign n40786 = ~n40782 & n40785;
  assign n40787 = ~n58822 & n32648;
  assign n40788 = ~n32648 & ~n39244;
  assign n40789 = ~pi162 & n29532;
  assign n40790 = ~n40788 & n40789;
  assign n40791 = ~n40787 & n40790;
  assign n40792 = ~n29532 & n39058;
  assign n40793 = ~n32648 & n40792;
  assign n40794 = pi299 & ~n40793;
  assign n40795 = ~n40791 & n40794;
  assign n40796 = ~n40786 & n40795;
  assign n40797 = ~pi51 & n39753;
  assign n40798 = pi140 & n39213;
  assign n40799 = n40797 & ~n40798;
  assign n40800 = n30958 & ~n40799;
  assign n40801 = ~pi51 & ~n39683;
  assign n40802 = pi140 & n39734;
  assign n40803 = n40801 & ~n40802;
  assign n40804 = n32690 & ~n40803;
  assign n40805 = ~n40800 & ~n40804;
  assign n40806 = ~n40796 & n40805;
  assign n40807 = pi232 & ~n40806;
  assign n40808 = n40779 & ~n40807;
  assign n40809 = ~n32698 & n39058;
  assign n40810 = ~n25479 & n40809;
  assign n40811 = ~pi100 & ~n40810;
  assign n40812 = ~n40808 & n40811;
  assign n40813 = ~n40044 & ~n40809;
  assign n40814 = pi100 & n40813;
  assign n40815 = n6311 & ~n40814;
  assign n40816 = ~n39282 & n40815;
  assign n40817 = ~n40812 & n40816;
  assign n40818 = pi87 & ~n29103;
  assign n40819 = n39286 & ~n40813;
  assign n40820 = ~n40818 & ~n40819;
  assign n40821 = ~n38944 & ~n40820;
  assign n40822 = pi130 & ~n40314;
  assign n40823 = ~pi130 & n40314;
  assign n40824 = ~n40822 & ~n40823;
  assign n40825 = ~n38935 & ~n40824;
  assign n40826 = ~n40821 & ~n40825;
  assign n40827 = ~n40817 & n40826;
  assign n40828 = ~n2829 & ~n40044;
  assign n40829 = ~n2680 & ~n39200;
  assign n40830 = ~n39569 & ~n40829;
  assign n40831 = ~pi224 & n40830;
  assign n40832 = ~n39251 & n39624;
  assign n40833 = pi224 & n40832;
  assign n40834 = n2829 & ~n40833;
  assign n40835 = pi224 & ~n40832;
  assign n40836 = ~pi224 & ~n40830;
  assign n40837 = ~n40835 & ~n40836;
  assign n40838 = n2829 & ~n40837;
  assign n40839 = ~n40831 & n40834;
  assign n40840 = ~n40828 & ~n60700;
  assign n40841 = pi140 & n40840;
  assign n40842 = n3890 & ~n40830;
  assign n40843 = ~n3890 & ~n40044;
  assign n40844 = ~n3890 & n40044;
  assign n40845 = n2829 & n40831;
  assign n40846 = ~n40844 & ~n40845;
  assign n40847 = ~n40842 & ~n40843;
  assign n40848 = ~pi140 & ~n60701;
  assign n40849 = n30958 & ~n40848;
  assign n40850 = ~n40841 & n40849;
  assign n40851 = ~n32648 & ~n39200;
  assign n40852 = pi169 & n39569;
  assign n40853 = ~n40851 & ~n40852;
  assign n40854 = ~pi216 & ~n40853;
  assign n40855 = ~pi51 & ~n39558;
  assign n40856 = ~pi169 & n40855;
  assign n40857 = pi169 & n40832;
  assign n40858 = pi162 & pi216;
  assign n40859 = ~n40857 & n40858;
  assign n40860 = ~n40856 & n40859;
  assign n40861 = ~n40854 & ~n40860;
  assign n40862 = n2852 & ~n40861;
  assign n40863 = pi169 & n39059;
  assign n40864 = ~pi51 & ~n40863;
  assign n40865 = ~n3906 & ~n40783;
  assign n40866 = ~n40864 & n40865;
  assign n40867 = ~n40862 & ~n40866;
  assign n40868 = pi299 & ~n40867;
  assign n40869 = n60632 & n39561;
  assign n40870 = ~pi51 & ~n40869;
  assign n40871 = pi140 & n40870;
  assign n40872 = ~pi51 & ~n39598;
  assign n40873 = ~pi140 & n40872;
  assign n40874 = n32690 & ~n40873;
  assign n40875 = ~n40871 & n40874;
  assign n40876 = ~n40868 & ~n40875;
  assign n40877 = ~n40850 & n40876;
  assign n40878 = pi232 & ~n40877;
  assign n40879 = n60632 & n60645;
  assign n40880 = ~pi51 & ~n40879;
  assign n40881 = ~pi232 & ~n40880;
  assign n40882 = pi39 & ~n40881;
  assign n40883 = ~n40878 & n40882;
  assign n40884 = ~pi232 & ~n39031;
  assign n40885 = ~pi39 & ~n40884;
  assign n40886 = ~n2680 & n39031;
  assign n40887 = ~n39454 & ~n40886;
  assign n40888 = ~n30960 & ~n40887;
  assign n40889 = n30960 & n39031;
  assign n40890 = pi232 & ~n40889;
  assign n40891 = ~n40888 & n40890;
  assign n40892 = n40885 & ~n40891;
  assign n40893 = ~n40883 & ~n40892;
  assign n40894 = ~pi38 & ~n40893;
  assign n40895 = pi38 & ~n40813;
  assign n40896 = ~pi100 & ~n40895;
  assign n40897 = ~n40894 & n40896;
  assign n40898 = n40815 & ~n40897;
  assign n40899 = n40820 & n40825;
  assign n40900 = ~n40898 & n40899;
  assign n40901 = ~n40827 & ~n40900;
  assign n40902 = n58992 & ~n40901;
  assign n40903 = ~pi51 & ~pi87;
  assign n40904 = ~n40863 & n40903;
  assign n40905 = n40825 & n40904;
  assign n40906 = ~pi87 & n39058;
  assign n40907 = ~pi87 & ~n30938;
  assign n40908 = n39058 & n40907;
  assign n40909 = ~n30938 & n40906;
  assign n40910 = pi87 & ~n29046;
  assign n40911 = ~n58992 & ~n40910;
  assign n40912 = ~n60702 & n40911;
  assign n40913 = ~n40905 & n40912;
  assign po287 = ~n40902 & ~n40913;
  assign n40915 = ~n2680 & ~n39106;
  assign n40916 = ~n39022 & ~n40915;
  assign n40917 = n31169 & n40916;
  assign n40918 = ~n31169 & n39106;
  assign n40919 = ~pi39 & pi176;
  assign n40920 = ~n40918 & n40919;
  assign n40921 = ~n40917 & n40920;
  assign n40922 = pi154 & pi232;
  assign n40923 = pi299 & n40922;
  assign n40924 = n40916 & n40923;
  assign n40925 = n39106 & ~n40923;
  assign n40926 = ~pi39 & ~pi176;
  assign n40927 = ~n40925 & n40926;
  assign n40928 = ~n40924 & n40927;
  assign n40929 = n2636 & n6308;
  assign n40930 = pi197 & n39213;
  assign n40931 = ~n2850 & ~n40930;
  assign n40932 = n2853 & ~n40931;
  assign n40933 = ~pi145 & ~n3890;
  assign n40934 = ~pi299 & ~n40933;
  assign n40935 = ~n39588 & n40934;
  assign n40936 = ~n40932 & ~n40935;
  assign n40937 = n58822 & ~n40936;
  assign n40938 = pi232 & ~n40937;
  assign n40939 = ~n39556 & ~n40938;
  assign n40940 = pi39 & ~n40939;
  assign n40941 = n40929 & ~n40940;
  assign n40942 = ~n40928 & n40941;
  assign n40943 = ~n40921 & n40941;
  assign n40944 = ~n40928 & n40943;
  assign n40945 = ~n40921 & n40942;
  assign n40946 = ~pi133 & ~n39409;
  assign n40947 = ~pi87 & n40946;
  assign n40948 = ~n60703 & n40947;
  assign n40949 = pi145 & n39218;
  assign n40950 = n39684 & ~n40949;
  assign n40951 = n39685 & ~n40930;
  assign n40952 = n38922 & ~n40951;
  assign n40953 = pi299 & ~n40952;
  assign n40954 = ~n40950 & ~n40953;
  assign n40955 = pi232 & ~n40954;
  assign n40956 = n39690 & ~n40955;
  assign n40957 = ~n31171 & n39001;
  assign n40958 = ~pi39 & n38922;
  assign n40959 = ~n40957 & n40958;
  assign n40960 = ~pi38 & ~n40959;
  assign n40961 = ~n40956 & n40960;
  assign n40962 = n38964 & ~n40961;
  assign n40963 = n39283 & ~n40962;
  assign n40964 = ~n39287 & ~n40963;
  assign n40965 = ~n40946 & ~n40964;
  assign n40966 = ~pi183 & ~pi299;
  assign n40967 = ~n33349 & ~n40966;
  assign n40968 = n2681 & n40967;
  assign n40969 = pi87 & ~n40968;
  assign n40970 = ~n40965 & ~n40969;
  assign n40971 = ~n40948 & n40970;
  assign n40972 = n58992 & ~n40971;
  assign n40973 = n38944 & ~n40946;
  assign n40974 = pi87 & n31185;
  assign n40975 = pi149 & n39420;
  assign n40976 = ~n58992 & ~n60704;
  assign n40977 = ~n40973 & n40976;
  assign n40978 = ~n40972 & ~n40977;
  assign n40979 = ~pi136 & n40823;
  assign n40980 = ~pi135 & n40979;
  assign n40981 = pi134 & ~n40980;
  assign n40982 = n38921 & ~n40981;
  assign n40983 = ~n58992 & n40903;
  assign n40984 = n32734 & ~n38921;
  assign n40985 = pi232 & n40984;
  assign n40986 = n40983 & ~n40985;
  assign n40987 = ~n40982 & n40986;
  assign n40988 = ~n32725 & n39058;
  assign n40989 = ~n40044 & ~n40988;
  assign n40990 = ~n2636 & n40989;
  assign n40991 = n6311 & ~n40990;
  assign n40992 = pi232 & ~n32724;
  assign n40993 = n40887 & n40992;
  assign n40994 = ~n39031 & ~n40992;
  assign n40995 = ~pi39 & ~n40994;
  assign n40996 = ~n40993 & n40995;
  assign n40997 = ~pi51 & ~n40984;
  assign n40998 = ~pi164 & pi216;
  assign n40999 = n2852 & ~n40998;
  assign n41000 = ~n40997 & ~n40999;
  assign n41001 = ~n32734 & ~n39200;
  assign n41002 = pi171 & n39569;
  assign n41003 = ~n41001 & ~n41002;
  assign n41004 = ~pi216 & ~n41003;
  assign n41005 = ~pi171 & n40855;
  assign n41006 = pi171 & n40832;
  assign n41007 = pi164 & pi216;
  assign n41008 = ~n41006 & n41007;
  assign n41009 = ~n41005 & n41008;
  assign n41010 = ~n41004 & ~n41009;
  assign n41011 = n2852 & ~n41010;
  assign n41012 = ~n41000 & ~n41011;
  assign n41013 = pi299 & ~n41012;
  assign n41014 = n32717 & n60701;
  assign n41015 = pi39 & pi186;
  assign n41016 = n32715 & ~n40872;
  assign n41017 = ~n41015 & ~n41016;
  assign n41018 = ~n41014 & n41017;
  assign n41019 = n32715 & ~n40870;
  assign n41020 = n32717 & ~n40840;
  assign n41021 = pi186 & ~n41020;
  assign n41022 = pi186 & ~n41019;
  assign n41023 = ~n41020 & n41022;
  assign n41024 = ~n41019 & n41021;
  assign n41025 = ~n41018 & ~n60705;
  assign n41026 = ~n41013 & ~n41025;
  assign n41027 = pi232 & ~n41026;
  assign n41028 = n40882 & ~n41027;
  assign n41029 = n2636 & ~n41028;
  assign n41030 = ~n40996 & n41029;
  assign n41031 = n40991 & ~n41030;
  assign n41032 = n39286 & ~n40989;
  assign n41033 = n40981 & ~n41032;
  assign n41034 = ~n41031 & n41033;
  assign n41035 = ~n39213 & n40797;
  assign n41036 = n32717 & ~n41035;
  assign n41037 = ~n39734 & n40801;
  assign n41038 = n32715 & ~n41037;
  assign n41039 = ~n41036 & ~n41038;
  assign n41040 = ~n32734 & n40792;
  assign n41041 = pi299 & ~n41040;
  assign n41042 = pi171 & ~n58822;
  assign n41043 = n2680 & n41042;
  assign n41044 = ~n32734 & ~n39244;
  assign n41045 = n29532 & ~n41044;
  assign n41046 = ~n41043 & n41045;
  assign n41047 = n41041 & ~n41046;
  assign n41048 = n41039 & ~n41047;
  assign n41049 = pi232 & ~n41048;
  assign n41050 = ~n40778 & ~n41049;
  assign n41051 = n41015 & ~n41050;
  assign n41052 = pi39 & ~pi186;
  assign n41053 = n32717 & ~n40797;
  assign n41054 = n32715 & ~n40801;
  assign n41055 = ~n41053 & ~n41054;
  assign n41056 = ~n41047 & n41055;
  assign n41057 = pi232 & ~n41056;
  assign n41058 = ~n40778 & ~n41057;
  assign n41059 = n41052 & ~n41058;
  assign n41060 = ~pi39 & ~n40988;
  assign n41061 = ~pi164 & ~n41060;
  assign n41062 = ~n41059 & n41061;
  assign n41063 = ~n41051 & n41062;
  assign n41064 = n41015 & ~n41039;
  assign n41065 = n41052 & ~n41055;
  assign n41066 = ~n41064 & ~n41065;
  assign n41067 = pi232 & ~n41066;
  assign n41068 = pi171 & ~n40781;
  assign n41069 = ~pi171 & ~n39733;
  assign n41070 = n29532 & ~n41069;
  assign n41071 = ~n41068 & n41070;
  assign n41072 = pi232 & n41041;
  assign n41073 = ~n41071 & n41072;
  assign n41074 = ~n40778 & ~n41073;
  assign n41075 = pi39 & ~n41074;
  assign n41076 = pi164 & ~n41060;
  assign n41077 = ~n41075 & n41076;
  assign n41078 = n41041 & ~n41071;
  assign n41079 = n41039 & ~n41078;
  assign n41080 = pi232 & ~n41079;
  assign n41081 = ~n40778 & ~n41080;
  assign n41082 = n41015 & ~n41081;
  assign n41083 = n41055 & ~n41078;
  assign n41084 = pi232 & ~n41083;
  assign n41085 = ~n40778 & ~n41084;
  assign n41086 = n41052 & ~n41085;
  assign n41087 = n41076 & ~n41086;
  assign n41088 = ~n41082 & n41087;
  assign n41089 = ~n41067 & n41077;
  assign n41090 = n2636 & ~n60706;
  assign n41091 = n2636 & ~n41063;
  assign n41092 = ~n60706 & n41091;
  assign n41093 = ~n41063 & n41090;
  assign n41094 = ~n40231 & n40991;
  assign n41095 = ~n60707 & n41094;
  assign n41096 = n39286 & n40988;
  assign n41097 = ~n40981 & ~n41096;
  assign n41098 = ~n41095 & n41097;
  assign n41099 = n58992 & ~n41098;
  assign n41100 = n58992 & ~n41034;
  assign n41101 = ~n41098 & n41100;
  assign n41102 = ~n41034 & n41099;
  assign n41103 = ~n40987 & ~n60708;
  assign n41104 = ~n32793 & ~n39200;
  assign n41105 = pi170 & n39569;
  assign n41106 = n3906 & ~n41105;
  assign n41107 = ~n41104 & n41106;
  assign n41108 = ~n29532 & ~n41107;
  assign n41109 = ~pi170 & n40855;
  assign n41110 = pi170 & n40832;
  assign n41111 = pi216 & ~n41110;
  assign n41112 = ~n41109 & n41111;
  assign n41113 = ~n41108 & ~n41112;
  assign n41114 = pi150 & pi299;
  assign n41115 = n32793 & ~n38921;
  assign n41116 = ~pi51 & ~n41115;
  assign n41117 = ~n2852 & n41116;
  assign n41118 = n41114 & ~n41117;
  assign n41119 = ~n41113 & n41118;
  assign n41120 = ~n3906 & n41116;
  assign n41121 = n40241 & ~n41120;
  assign n41122 = ~n41107 & n41121;
  assign n41123 = ~n41119 & ~n41122;
  assign n41124 = pi185 & n40870;
  assign n41125 = ~pi185 & n40872;
  assign n41126 = ~pi299 & ~n41125;
  assign n41127 = ~n41124 & n41126;
  assign n41128 = n41123 & ~n41127;
  assign n41129 = pi232 & ~n41128;
  assign n41130 = n40882 & ~n41129;
  assign n41131 = ~pi299 & ~n39031;
  assign n41132 = pi170 & ~n40887;
  assign n41133 = ~pi170 & n39031;
  assign n41134 = n32792 & ~n41133;
  assign n41135 = ~n41132 & n41134;
  assign n41136 = n40885 & ~n41135;
  assign n41137 = ~n41131 & n41136;
  assign n41138 = ~n41130 & ~n41137;
  assign n41139 = ~pi38 & ~n41138;
  assign n41140 = ~n32834 & n39058;
  assign n41141 = ~n40044 & ~n41140;
  assign n41142 = pi38 & ~n41141;
  assign n41143 = ~pi194 & ~n41142;
  assign n41144 = ~n41139 & n41143;
  assign n41145 = pi185 & n40840;
  assign n41146 = ~pi185 & ~n60701;
  assign n41147 = ~pi299 & ~n41146;
  assign n41148 = ~pi299 & ~n41145;
  assign n41149 = ~n41146 & n41148;
  assign n41150 = ~n41145 & n41147;
  assign n41151 = n41123 & ~n60709;
  assign n41152 = pi232 & ~n41151;
  assign n41153 = n40882 & ~n41152;
  assign n41154 = n32622 & n40887;
  assign n41155 = n41136 & ~n41154;
  assign n41156 = ~n41153 & ~n41155;
  assign n41157 = ~pi38 & ~n41156;
  assign n41158 = n32842 & n39058;
  assign n41159 = ~n40044 & ~n41158;
  assign n41160 = pi38 & ~n41159;
  assign n41161 = pi194 & ~n41160;
  assign n41162 = ~n41157 & n41161;
  assign n41163 = ~n41144 & ~n41162;
  assign n41164 = ~pi100 & ~n41163;
  assign n41165 = pi194 & n29623;
  assign n41166 = n41140 & ~n41165;
  assign n41167 = ~n40044 & ~n41166;
  assign n41168 = pi100 & n41167;
  assign n41169 = n6311 & ~n41168;
  assign n41170 = ~n41164 & n41169;
  assign n41171 = pi135 & ~n40979;
  assign n41172 = pi134 & n40980;
  assign n41173 = ~n41171 & ~n41172;
  assign n41174 = n39286 & ~n41167;
  assign n41175 = ~n41173 & ~n41174;
  assign n41176 = ~n41170 & n41175;
  assign n41177 = pi185 & n39734;
  assign n41178 = n40801 & ~n41177;
  assign n41179 = ~n25479 & n41140;
  assign n41180 = ~pi194 & ~n41179;
  assign n41181 = ~n41178 & n41180;
  assign n41182 = ~n25479 & n41158;
  assign n41183 = pi194 & ~n41182;
  assign n41184 = pi185 & n39213;
  assign n41185 = n40797 & ~n41184;
  assign n41186 = ~pi185 & n40797;
  assign n41187 = ~n41035 & n41183;
  assign n41188 = ~n41186 & n41187;
  assign n41189 = n41183 & ~n41185;
  assign n41190 = ~n41181 & ~n60710;
  assign n41191 = ~pi299 & ~n41190;
  assign n41192 = pi170 & ~n40781;
  assign n41193 = ~pi170 & ~n39733;
  assign n41194 = n29532 & ~n41193;
  assign n41195 = ~n41192 & n41194;
  assign n41196 = n41114 & ~n41195;
  assign n41197 = pi170 & ~n58822;
  assign n41198 = n2680 & n41197;
  assign n41199 = ~n32793 & ~n39244;
  assign n41200 = n29532 & ~n41199;
  assign n41201 = ~n41198 & n41200;
  assign n41202 = n40241 & ~n41201;
  assign n41203 = ~n41196 & ~n41202;
  assign n41204 = ~n32793 & n40792;
  assign n41205 = ~n41180 & ~n41183;
  assign n41206 = ~n41204 & ~n41205;
  assign n41207 = ~n41203 & n41206;
  assign n41208 = ~n41191 & ~n41207;
  assign n41209 = pi232 & ~n41208;
  assign n41210 = ~n40779 & ~n41205;
  assign n41211 = ~n41209 & ~n41210;
  assign n41212 = ~pi100 & ~n41211;
  assign n41213 = ~n39282 & n41169;
  assign n41214 = n39283 & ~n41168;
  assign n41215 = ~n41212 & n60711;
  assign n41216 = n39286 & n41166;
  assign n41217 = n41173 & ~n41216;
  assign n41218 = ~n41215 & n41217;
  assign n41219 = n58992 & ~n41218;
  assign n41220 = ~n41176 & n41219;
  assign n41221 = n38921 & n41173;
  assign n41222 = n32841 & ~n38921;
  assign n41223 = pi232 & n41115;
  assign n41224 = n40983 & ~n60712;
  assign n41225 = ~n41221 & n41224;
  assign n41226 = ~n41220 & ~n41225;
  assign n41227 = pi136 & ~n40823;
  assign n41228 = ~n40979 & ~n41227;
  assign n41229 = ~n38934 & ~n41228;
  assign n41230 = ~n39058 & n41229;
  assign n41231 = pi148 & n2681;
  assign n41232 = ~n38921 & ~n41231;
  assign n41233 = ~n41230 & ~n41232;
  assign n41234 = n40983 & ~n41233;
  assign n41235 = ~n29091 & ~n40887;
  assign n41236 = n29091 & n39031;
  assign n41237 = pi232 & ~n41236;
  assign n41238 = ~n41235 & n41237;
  assign n41239 = n40885 & ~n41238;
  assign n41240 = pi184 & n40840;
  assign n41241 = ~pi184 & ~n60701;
  assign n41242 = n29089 & ~n41241;
  assign n41243 = ~n41240 & n41242;
  assign n41244 = pi184 & n40870;
  assign n41245 = ~pi141 & ~pi299;
  assign n41246 = ~pi184 & n40872;
  assign n41247 = n41245 & ~n41246;
  assign n41248 = ~n41244 & n41247;
  assign n41249 = n3906 & ~n40830;
  assign n41250 = pi163 & n2852;
  assign n41251 = ~n40832 & n41250;
  assign n41252 = ~n3906 & ~n41250;
  assign n41253 = ~n40044 & n41252;
  assign n41254 = pi148 & ~n41253;
  assign n41255 = n40832 & n41250;
  assign n41256 = ~n2852 & n40044;
  assign n41257 = ~n3906 & ~n40044;
  assign n41258 = ~pi163 & ~n41257;
  assign n41259 = ~n41256 & ~n41258;
  assign n41260 = ~n41255 & n41259;
  assign n41261 = pi148 & ~n41260;
  assign n41262 = ~n41251 & n41254;
  assign n41263 = ~n41249 & n60713;
  assign n41264 = ~pi287 & n30546;
  assign n41265 = pi216 & ~n41264;
  assign n41266 = n2852 & ~n41265;
  assign n41267 = n60632 & n41266;
  assign n41268 = ~pi51 & ~pi148;
  assign n41269 = ~n41267 & n41268;
  assign n41270 = pi299 & ~n41269;
  assign n41271 = ~n41263 & n41270;
  assign n41272 = ~n41248 & ~n41271;
  assign n41273 = ~n41243 & n41272;
  assign n41274 = pi232 & ~n41273;
  assign n41275 = n40882 & ~n41274;
  assign n41276 = n2636 & ~n41275;
  assign n41277 = ~n41239 & n41276;
  assign n41278 = n29092 & ~n38921;
  assign n41279 = ~pi51 & ~n41278;
  assign n41280 = ~n2636 & ~n41279;
  assign n41281 = n6311 & ~n41280;
  assign n41282 = ~n41277 & n41281;
  assign n41283 = n39286 & n41279;
  assign n41284 = n41229 & ~n41283;
  assign n41285 = ~n41282 & n41284;
  assign n41286 = ~n36293 & ~n38921;
  assign n41287 = n41279 & n41286;
  assign n41288 = ~pi51 & n39685;
  assign n41289 = ~pi148 & ~n41288;
  assign n41290 = ~n41264 & ~n41289;
  assign n41291 = ~pi148 & n39058;
  assign n41292 = ~n41290 & ~n41291;
  assign n41293 = n29532 & n40780;
  assign n41294 = ~n2680 & n40792;
  assign n41295 = pi148 & ~n41294;
  assign n41296 = ~n41293 & n41295;
  assign n41297 = ~n41292 & ~n41296;
  assign n41298 = pi299 & ~n41297;
  assign n41299 = pi184 & n39213;
  assign n41300 = n40797 & ~n41299;
  assign n41301 = n29089 & ~n41300;
  assign n41302 = pi184 & n39734;
  assign n41303 = n40801 & ~n41302;
  assign n41304 = n41245 & ~n41303;
  assign n41305 = ~n41301 & ~n41304;
  assign n41306 = ~n41298 & ~n41304;
  assign n41307 = ~n41301 & n41306;
  assign n41308 = ~n41298 & n41305;
  assign n41309 = pi232 & ~n60714;
  assign n41310 = ~pi100 & n40779;
  assign n41311 = ~n41309 & n41310;
  assign n41312 = ~n41287 & ~n41311;
  assign n41313 = n6311 & ~n41312;
  assign n41314 = ~n38921 & n41283;
  assign n41315 = ~n41229 & ~n41314;
  assign n41316 = ~n41313 & n41315;
  assign n41317 = n58992 & ~n41316;
  assign n41318 = ~n41285 & n41317;
  assign n41319 = ~n41234 & ~n41318;
  assign n41320 = pi215 & pi1142;
  assign n41321 = pi299 & ~n41320;
  assign n41322 = ~pi932 & n38221;
  assign n41323 = ~pi1142 & ~n38221;
  assign n41324 = pi221 & ~n41323;
  assign n41325 = pi221 & ~n41322;
  assign n41326 = ~n41323 & n41325;
  assign n41327 = ~n41322 & n41324;
  assign n41328 = pi216 & pi277;
  assign n41329 = ~pi221 & ~n41328;
  assign n41330 = ~pi72 & ~n40742;
  assign n41331 = ~n28318 & ~n41330;
  assign n41332 = n2620 & ~n41331;
  assign n41333 = n40605 & ~n41332;
  assign n41334 = ~pi95 & ~n41333;
  assign n41335 = n38365 & ~n41334;
  assign n41336 = ~pi262 & n41335;
  assign n41337 = pi172 & ~n41336;
  assign n41338 = pi262 & n40747;
  assign n41339 = n2599 & n31407;
  assign n41340 = ~n28313 & ~n41339;
  assign n41341 = ~pi262 & n41340;
  assign n41342 = ~pi172 & ~n31400;
  assign n41343 = ~n41341 & n41342;
  assign n41344 = ~n41338 & n41343;
  assign n41345 = ~pi228 & ~n41344;
  assign n41346 = ~n31400 & ~n41340;
  assign n41347 = ~pi262 & n41346;
  assign n41348 = ~pi172 & ~n41347;
  assign n41349 = pi172 & ~pi262;
  assign n41350 = n41335 & n41349;
  assign n41351 = ~n41348 & ~n41350;
  assign n41352 = pi262 & n40748;
  assign n41353 = ~pi228 & ~n41352;
  assign n41354 = ~n41351 & n41353;
  assign n41355 = ~n41337 & n41345;
  assign n41356 = pi105 & ~n41340;
  assign n41357 = pi262 & ~n28313;
  assign n41358 = pi105 & n41357;
  assign n41359 = ~n41339 & n41358;
  assign n41360 = ~pi105 & pi172;
  assign n41361 = pi228 & ~n41360;
  assign n41362 = ~n41359 & n41361;
  assign n41363 = ~n41356 & n41362;
  assign n41364 = ~pi216 & ~n41363;
  assign n41365 = ~n60716 & n41364;
  assign n41366 = n41329 & ~n41365;
  assign n41367 = ~n60715 & ~n41366;
  assign n41368 = ~pi215 & ~n41367;
  assign n41369 = n41321 & ~n41368;
  assign n41370 = pi223 & pi1142;
  assign n41371 = ~pi299 & ~n41370;
  assign n41372 = ~pi932 & n38636;
  assign n41373 = ~pi1142 & ~n38636;
  assign n41374 = pi222 & ~n41373;
  assign n41375 = pi222 & ~n41372;
  assign n41376 = ~n41373 & n41375;
  assign n41377 = ~n41372 & n41374;
  assign n41378 = pi224 & pi277;
  assign n41379 = ~pi222 & ~n41378;
  assign n41380 = ~pi224 & ~n41341;
  assign n41381 = n41379 & ~n41380;
  assign n41382 = ~n60717 & ~n41381;
  assign n41383 = n41371 & n41382;
  assign n41384 = ~n41340 & n41379;
  assign n41385 = n41382 & ~n41384;
  assign n41386 = ~pi223 & ~n41385;
  assign n41387 = n41371 & ~n41386;
  assign n41388 = ~pi39 & ~n41387;
  assign n41389 = ~n41383 & n41388;
  assign n41390 = ~n41369 & n41389;
  assign n41391 = n28313 & n35583;
  assign n41392 = ~pi224 & n41357;
  assign n41393 = n41379 & ~n41392;
  assign n41394 = ~n60717 & ~n41393;
  assign n41395 = ~pi223 & ~n41394;
  assign n41396 = ~n41370 & ~n41395;
  assign n41397 = ~pi299 & ~n41396;
  assign n41398 = ~n41391 & n41397;
  assign n41399 = ~pi262 & n58822;
  assign n41400 = pi172 & ~pi228;
  assign n41401 = ~n31586 & ~n41400;
  assign n41402 = ~n41399 & ~n41401;
  assign n41403 = n28313 & n38211;
  assign n41404 = ~n41358 & ~n41360;
  assign n41405 = pi228 & ~n41404;
  assign n41406 = ~n41403 & ~n41405;
  assign n41407 = ~n41402 & n41406;
  assign n41408 = ~pi216 & ~n41407;
  assign n41409 = n41329 & ~n41408;
  assign n41410 = ~n60715 & ~n41409;
  assign n41411 = ~pi215 & ~n41410;
  assign n41412 = ~n41320 & ~n41411;
  assign n41413 = pi299 & ~n41412;
  assign n41414 = ~n41398 & ~n41413;
  assign n41415 = pi39 & ~n41414;
  assign n41416 = ~pi38 & ~n41415;
  assign n41417 = ~n41390 & n41416;
  assign n41418 = n35591 & n41403;
  assign n41419 = ~n41400 & ~n41405;
  assign n41420 = ~pi216 & ~n41419;
  assign n41421 = n41329 & ~n41420;
  assign n41422 = ~n60715 & ~n41421;
  assign n41423 = ~pi215 & ~n41422;
  assign n41424 = ~n41320 & ~n41423;
  assign n41425 = ~n41418 & ~n41424;
  assign n41426 = pi299 & n41425;
  assign n41427 = ~n41398 & ~n41426;
  assign n41428 = pi38 & n41427;
  assign n41429 = ~pi100 & ~n41428;
  assign n41430 = ~n41417 & n41429;
  assign n41431 = ~pi146 & ~n58822;
  assign n41432 = pi146 & ~n28550;
  assign n41433 = ~n41431 & ~n41432;
  assign n41434 = pi152 & ~n41433;
  assign n41435 = ~n37718 & n41433;
  assign n41436 = n28550 & n37718;
  assign n41437 = ~pi152 & ~n41436;
  assign n41438 = ~n41435 & n41437;
  assign n41439 = ~n41434 & ~n41438;
  assign n41440 = ~pi262 & n41439;
  assign n41441 = ~pi228 & n41439;
  assign n41442 = ~n41400 & ~n41441;
  assign n41443 = ~n41440 & ~n41442;
  assign n41444 = n41406 & ~n41443;
  assign n41445 = ~pi216 & ~n41444;
  assign n41446 = n41329 & ~n41445;
  assign n41447 = ~n60715 & ~n41446;
  assign n41448 = ~pi215 & ~n41447;
  assign n41449 = ~n41320 & ~n41448;
  assign n41450 = pi299 & ~n41449;
  assign n41451 = n2634 & ~n41398;
  assign n41452 = ~n41450 & n41451;
  assign n41453 = ~n2634 & n41427;
  assign n41454 = pi100 & ~n41453;
  assign n41455 = ~n41452 & n41454;
  assign n41456 = ~n41430 & ~n41455;
  assign n41457 = ~pi87 & ~n41456;
  assign n41458 = ~n58815 & n41427;
  assign n41459 = n58815 & n41414;
  assign n41460 = ~n41458 & ~n41459;
  assign n41461 = pi87 & n41460;
  assign n41462 = ~pi75 & ~n41461;
  assign n41463 = ~n41457 & n41462;
  assign n41464 = pi75 & n41427;
  assign n41465 = ~pi92 & ~n41464;
  assign n41466 = ~n41463 & n41465;
  assign n41467 = n6309 & ~n41460;
  assign n41468 = ~n6309 & n41427;
  assign n41469 = pi92 & ~n41468;
  assign n41470 = ~n41467 & n41469;
  assign n41471 = n6306 & ~n41470;
  assign n41472 = ~n41466 & n41471;
  assign n41473 = ~n6306 & n41427;
  assign n41474 = ~pi55 & ~n41473;
  assign n41475 = ~n41472 & n41474;
  assign n41476 = n28288 & n41412;
  assign n41477 = ~n28288 & ~n41425;
  assign n41478 = pi55 & ~n41477;
  assign n41479 = ~n41476 & n41478;
  assign n41480 = ~pi56 & ~n41479;
  assign n41481 = ~n41475 & n41480;
  assign n41482 = n60070 & ~n41412;
  assign n41483 = ~n60070 & n41425;
  assign n41484 = pi56 & ~n41483;
  assign n41485 = ~n60070 & ~n41425;
  assign n41486 = ~pi55 & n41476;
  assign n41487 = ~n41485 & ~n41486;
  assign n41488 = pi56 & ~n41487;
  assign n41489 = ~n41482 & n41484;
  assign n41490 = ~pi62 & ~n60718;
  assign n41491 = ~n41481 & n41490;
  assign n41492 = n58815 & n31573;
  assign n41493 = n41412 & n41492;
  assign n41494 = ~n41425 & ~n41492;
  assign n41495 = pi62 & ~n41494;
  assign n41496 = ~n41493 & n41495;
  assign n41497 = n4438 & ~n41496;
  assign n41498 = ~n41491 & n41497;
  assign n41499 = ~n4438 & ~n41425;
  assign n41500 = ~pi249 & ~n41499;
  assign n41501 = ~n41498 & n41500;
  assign n41502 = pi262 & n41335;
  assign n41503 = ~pi172 & ~n41502;
  assign n41504 = ~pi262 & ~n40748;
  assign n41505 = pi262 & ~n41346;
  assign n41506 = pi172 & ~n41505;
  assign n41507 = ~n41504 & n41506;
  assign n41508 = ~n41503 & ~n41507;
  assign n41509 = ~pi228 & ~n41508;
  assign n41510 = ~pi216 & ~n41362;
  assign n41511 = ~n41509 & n41510;
  assign n41512 = n41329 & ~n41511;
  assign n41513 = ~n60715 & ~n41512;
  assign n41514 = ~pi215 & ~n41513;
  assign n41515 = n41321 & ~n41514;
  assign n41516 = n41388 & ~n41515;
  assign n41517 = ~n41402 & ~n41405;
  assign n41518 = ~pi216 & ~n41517;
  assign n41519 = n41329 & ~n41518;
  assign n41520 = ~n60715 & ~n41519;
  assign n41521 = ~pi215 & ~n41520;
  assign n41522 = ~n41320 & ~n41521;
  assign n41523 = pi299 & ~n41522;
  assign n41524 = ~n41397 & ~n41523;
  assign n41525 = pi39 & ~n41524;
  assign n41526 = ~pi38 & ~n41525;
  assign n41527 = ~n41516 & n41526;
  assign n41528 = pi299 & ~n41424;
  assign n41529 = ~n41397 & ~n41528;
  assign n41530 = pi38 & n41529;
  assign n41531 = ~pi100 & ~n41530;
  assign n41532 = ~n41527 & n41531;
  assign n41533 = ~n41405 & ~n41443;
  assign n41534 = ~pi216 & ~n41533;
  assign n41535 = n41329 & ~n41534;
  assign n41536 = ~n60715 & ~n41535;
  assign n41537 = ~pi215 & ~n41536;
  assign n41538 = ~n41320 & ~n41537;
  assign n41539 = pi299 & ~n41538;
  assign n41540 = n2634 & ~n41397;
  assign n41541 = ~n41539 & n41540;
  assign n41542 = ~n2634 & n41529;
  assign n41543 = pi100 & ~n41542;
  assign n41544 = ~n41541 & n41543;
  assign n41545 = ~n41532 & ~n41544;
  assign n41546 = ~pi87 & ~n41545;
  assign n41547 = ~n58815 & n41529;
  assign n41548 = n58815 & n41524;
  assign n41549 = ~n41547 & ~n41548;
  assign n41550 = pi87 & n41549;
  assign n41551 = ~pi75 & ~n41550;
  assign n41552 = ~n41546 & n41551;
  assign n41553 = pi75 & n41529;
  assign n41554 = ~pi92 & ~n41553;
  assign n41555 = ~n41552 & n41554;
  assign n41556 = n6309 & ~n41549;
  assign n41557 = ~n6309 & n41529;
  assign n41558 = pi92 & ~n41557;
  assign n41559 = ~n41556 & n41558;
  assign n41560 = n6306 & ~n41559;
  assign n41561 = ~n41555 & n41560;
  assign n41562 = ~n6306 & n41529;
  assign n41563 = ~pi55 & ~n41562;
  assign n41564 = ~n41561 & n41563;
  assign n41565 = n28288 & n41522;
  assign n41566 = ~n28288 & n41424;
  assign n41567 = pi55 & ~n41566;
  assign n41568 = ~n41565 & n41567;
  assign n41569 = ~pi56 & ~n41568;
  assign n41570 = ~n41564 & n41569;
  assign n41571 = n60070 & ~n41522;
  assign n41572 = ~n60070 & ~n41424;
  assign n41573 = pi56 & ~n41572;
  assign n41574 = ~n60070 & n41424;
  assign n41575 = ~pi55 & n41565;
  assign n41576 = ~n41574 & ~n41575;
  assign n41577 = pi56 & ~n41576;
  assign n41578 = ~n41571 & n41573;
  assign n41579 = ~pi62 & ~n60719;
  assign n41580 = ~n41570 & n41579;
  assign n41581 = n41492 & n41522;
  assign n41582 = n41424 & ~n41492;
  assign n41583 = pi62 & ~n41582;
  assign n41584 = ~n41581 & n41583;
  assign n41585 = n4438 & ~n41584;
  assign n41586 = ~n41580 & n41585;
  assign n41587 = ~n4438 & n41424;
  assign n41588 = pi249 & ~n41587;
  assign n41589 = ~n41586 & n41588;
  assign n41590 = ~n41501 & ~n41589;
  assign n41591 = pi223 & pi1141;
  assign n41592 = ~pi299 & ~n41591;
  assign n41593 = ~pi935 & n38636;
  assign n41594 = ~pi1141 & ~n38636;
  assign n41595 = pi222 & ~n41594;
  assign n41596 = pi222 & ~n41593;
  assign n41597 = ~n41594 & n41596;
  assign n41598 = ~n41593 & n41595;
  assign n41599 = pi224 & pi270;
  assign n41600 = ~pi222 & ~n41599;
  assign n41601 = pi861 & n41340;
  assign n41602 = ~pi224 & ~n41601;
  assign n41603 = n41600 & ~n41602;
  assign n41604 = ~n60720 & ~n41603;
  assign n41605 = ~n41340 & n41600;
  assign n41606 = n41604 & ~n41605;
  assign n41607 = ~pi223 & ~n41606;
  assign n41608 = n41592 & ~n41607;
  assign n41609 = ~pi39 & ~n41608;
  assign n41610 = pi215 & pi1141;
  assign n41611 = pi299 & ~n41610;
  assign n41612 = ~pi935 & n38221;
  assign n41613 = ~pi1141 & ~n38221;
  assign n41614 = pi221 & ~n41613;
  assign n41615 = pi221 & ~n41612;
  assign n41616 = ~n41613 & n41615;
  assign n41617 = ~n41612 & n41614;
  assign n41618 = pi216 & pi270;
  assign n41619 = ~pi221 & ~n41618;
  assign n41620 = ~pi861 & n41335;
  assign n41621 = ~pi171 & ~n41620;
  assign n41622 = pi861 & ~n40748;
  assign n41623 = ~pi861 & ~n41346;
  assign n41624 = pi171 & ~n41623;
  assign n41625 = ~n41622 & n41624;
  assign n41626 = ~n41621 & ~n41625;
  assign n41627 = ~pi228 & ~n41626;
  assign n41628 = n38211 & ~n41340;
  assign n41629 = pi861 & ~n28313;
  assign n41630 = pi105 & ~n41629;
  assign n41631 = ~pi105 & pi171;
  assign n41632 = pi228 & ~n41631;
  assign n41633 = ~n41630 & n41632;
  assign n41634 = ~pi216 & ~n41633;
  assign n41635 = ~n41628 & n41634;
  assign n41636 = ~n41627 & n41635;
  assign n41637 = n41619 & ~n41636;
  assign n41638 = ~n60721 & ~n41637;
  assign n41639 = ~pi215 & ~n41638;
  assign n41640 = n41611 & ~n41639;
  assign n41641 = n41609 & ~n41640;
  assign n41642 = ~pi299 & n41391;
  assign n41643 = n28313 & n35582;
  assign n41644 = ~pi224 & ~n41629;
  assign n41645 = n41600 & ~n41644;
  assign n41646 = ~n60720 & ~n41645;
  assign n41647 = ~pi223 & ~n41646;
  assign n41648 = ~n41591 & ~n41647;
  assign n41649 = ~pi299 & ~n41648;
  assign n41650 = ~n60722 & ~n41649;
  assign n41651 = ~pi861 & n58822;
  assign n41652 = ~pi228 & ~n41042;
  assign n41653 = ~pi228 & ~n41651;
  assign n41654 = ~n41042 & n41653;
  assign n41655 = ~n41651 & n41652;
  assign n41656 = ~n41403 & n41634;
  assign n41657 = ~n60723 & n41656;
  assign n41658 = n41619 & ~n41657;
  assign n41659 = ~n60721 & ~n41658;
  assign n41660 = ~pi215 & ~n41659;
  assign n41661 = ~n41610 & ~n41660;
  assign n41662 = pi299 & ~n41661;
  assign n41663 = n41650 & ~n41662;
  assign n41664 = pi39 & ~n41663;
  assign n41665 = ~pi38 & ~n41664;
  assign n41666 = ~n41641 & n41665;
  assign n41667 = ~pi171 & ~pi228;
  assign n41668 = n41634 & ~n41667;
  assign n41669 = n41619 & ~n41668;
  assign n41670 = ~n60721 & ~n41669;
  assign n41671 = ~pi215 & ~n41670;
  assign n41672 = ~n41610 & ~n41671;
  assign n41673 = n38239 & n41403;
  assign n41674 = ~n41618 & n41673;
  assign n41675 = n41672 & ~n41674;
  assign n41676 = pi299 & ~n41675;
  assign n41677 = n41650 & ~n41676;
  assign n41678 = pi38 & n41677;
  assign n41679 = ~pi100 & ~n41678;
  assign n41680 = ~n41666 & n41679;
  assign n41681 = pi171 & ~n41439;
  assign n41682 = ~pi861 & n41439;
  assign n41683 = ~pi228 & ~n41682;
  assign n41684 = ~pi228 & ~n41681;
  assign n41685 = ~n41682 & n41684;
  assign n41686 = ~n41681 & n41683;
  assign n41687 = n41656 & ~n60724;
  assign n41688 = n41619 & ~n41687;
  assign n41689 = ~n60721 & ~n41688;
  assign n41690 = ~pi215 & ~n41689;
  assign n41691 = ~n41610 & ~n41690;
  assign n41692 = pi299 & ~n41691;
  assign n41693 = n2634 & n41650;
  assign n41694 = ~n41692 & n41693;
  assign n41695 = ~n2634 & n41677;
  assign n41696 = pi100 & ~n41695;
  assign n41697 = ~n41694 & n41696;
  assign n41698 = ~n41680 & ~n41697;
  assign n41699 = ~pi87 & ~n41698;
  assign n41700 = ~n58815 & n41677;
  assign n41701 = n58815 & n41663;
  assign n41702 = ~n41700 & ~n41701;
  assign n41703 = pi87 & n41702;
  assign n41704 = ~pi75 & ~n41703;
  assign n41705 = ~n41699 & n41704;
  assign n41706 = pi75 & n41677;
  assign n41707 = ~pi92 & ~n41706;
  assign n41708 = ~n41705 & n41707;
  assign n41709 = n6309 & ~n41702;
  assign n41710 = ~n6309 & n41677;
  assign n41711 = pi92 & ~n41710;
  assign n41712 = ~n41709 & n41711;
  assign n41713 = n6306 & ~n41712;
  assign n41714 = ~n41708 & n41713;
  assign n41715 = ~n6306 & n41677;
  assign n41716 = ~pi55 & ~n41715;
  assign n41717 = ~n41714 & n41716;
  assign n41718 = n28288 & n41661;
  assign n41719 = ~n28288 & n41675;
  assign n41720 = pi55 & ~n41719;
  assign n41721 = ~n41718 & n41720;
  assign n41722 = ~pi56 & ~n41721;
  assign n41723 = ~n41717 & n41722;
  assign n41724 = n60070 & ~n41661;
  assign n41725 = ~n60070 & ~n41675;
  assign n41726 = pi56 & ~n41725;
  assign n41727 = ~pi55 & n41718;
  assign n41728 = ~n60070 & n41675;
  assign n41729 = ~n41727 & ~n41728;
  assign n41730 = pi56 & ~n41729;
  assign n41731 = ~n41724 & n41726;
  assign n41732 = ~pi62 & ~n60725;
  assign n41733 = ~n41723 & n41732;
  assign n41734 = n41492 & n41661;
  assign n41735 = ~n41492 & n41675;
  assign n41736 = pi62 & ~n41735;
  assign n41737 = ~n41734 & n41736;
  assign n41738 = pi241 & n4438;
  assign n41739 = ~n41737 & n41738;
  assign n41740 = ~n41733 & n41739;
  assign n41741 = ~pi861 & n40747;
  assign n41742 = ~n31400 & ~n41601;
  assign n41743 = ~n41741 & n41742;
  assign n41744 = ~pi861 & n40748;
  assign n41745 = pi861 & n41346;
  assign n41746 = ~pi171 & ~n41745;
  assign n41747 = ~n41744 & n41746;
  assign n41748 = ~pi171 & ~n41743;
  assign n41749 = pi171 & pi861;
  assign n41750 = n41335 & n41749;
  assign n41751 = pi171 & n41335;
  assign n41752 = ~n41746 & ~n41751;
  assign n41753 = pi861 & ~n41752;
  assign n41754 = ~n40748 & n41746;
  assign n41755 = ~n41753 & ~n41754;
  assign n41756 = ~n60726 & ~n41750;
  assign n41757 = ~pi228 & ~n60727;
  assign n41758 = ~n41356 & n41633;
  assign n41759 = ~pi216 & ~n41758;
  assign n41760 = ~n41757 & n41759;
  assign n41761 = n41619 & ~n41760;
  assign n41762 = ~n60721 & ~n41761;
  assign n41763 = ~pi215 & ~n41762;
  assign n41764 = n41611 & ~n41763;
  assign n41765 = n41592 & n41604;
  assign n41766 = n41609 & ~n41765;
  assign n41767 = ~n41764 & n41766;
  assign n41768 = n41634 & ~n60723;
  assign n41769 = n41619 & ~n41768;
  assign n41770 = ~n60721 & ~n41769;
  assign n41771 = ~pi215 & ~n41770;
  assign n41772 = ~n41610 & ~n41771;
  assign n41773 = pi299 & ~n41772;
  assign n41774 = ~n41649 & ~n41773;
  assign n41775 = pi39 & ~n41774;
  assign n41776 = ~pi38 & ~n41775;
  assign n41777 = ~n41767 & n41776;
  assign n41778 = pi299 & ~n41672;
  assign n41779 = ~n41649 & ~n41778;
  assign n41780 = pi38 & n41779;
  assign n41781 = ~pi100 & ~n41780;
  assign n41782 = ~n41777 & n41781;
  assign n41783 = n41634 & ~n60724;
  assign n41784 = n41619 & ~n41783;
  assign n41785 = ~n60721 & ~n41784;
  assign n41786 = ~pi215 & ~n41785;
  assign n41787 = ~n41610 & ~n41786;
  assign n41788 = pi299 & ~n41787;
  assign n41789 = n2634 & ~n41649;
  assign n41790 = ~n41788 & n41789;
  assign n41791 = ~n2634 & n41779;
  assign n41792 = pi100 & ~n41791;
  assign n41793 = ~n41790 & n41792;
  assign n41794 = ~n41782 & ~n41793;
  assign n41795 = ~pi87 & ~n41794;
  assign n41796 = ~n58815 & n41779;
  assign n41797 = n58815 & n41774;
  assign n41798 = ~n41796 & ~n41797;
  assign n41799 = pi87 & n41798;
  assign n41800 = ~pi75 & ~n41799;
  assign n41801 = ~n41795 & n41800;
  assign n41802 = pi75 & n41779;
  assign n41803 = ~pi92 & ~n41802;
  assign n41804 = ~n41801 & n41803;
  assign n41805 = n6309 & ~n41798;
  assign n41806 = ~n6309 & n41779;
  assign n41807 = pi92 & ~n41806;
  assign n41808 = ~n41805 & n41807;
  assign n41809 = n6306 & ~n41808;
  assign n41810 = ~n41804 & n41809;
  assign n41811 = ~n6306 & n41779;
  assign n41812 = ~pi55 & ~n41811;
  assign n41813 = ~n41810 & n41812;
  assign n41814 = n28288 & n41772;
  assign n41815 = ~n28288 & n41672;
  assign n41816 = pi55 & ~n41815;
  assign n41817 = ~n41814 & n41816;
  assign n41818 = ~pi56 & ~n41817;
  assign n41819 = ~n41813 & n41818;
  assign n41820 = n60070 & ~n41772;
  assign n41821 = ~n60070 & ~n41672;
  assign n41822 = pi56 & ~n41821;
  assign n41823 = ~n60070 & n41672;
  assign n41824 = ~pi55 & n41814;
  assign n41825 = ~n41823 & ~n41824;
  assign n41826 = pi56 & ~n41825;
  assign n41827 = ~n41820 & n41822;
  assign n41828 = ~pi62 & ~n60728;
  assign n41829 = ~n41819 & n41828;
  assign n41830 = n41492 & n41772;
  assign n41831 = ~n41492 & n41672;
  assign n41832 = pi62 & ~n41831;
  assign n41833 = ~n41830 & n41832;
  assign n41834 = ~pi241 & n4438;
  assign n41835 = ~n41833 & n41834;
  assign n41836 = ~n41829 & n41835;
  assign n41837 = pi241 & n41674;
  assign n41838 = ~n4438 & ~n41837;
  assign n41839 = n41672 & n41838;
  assign n41840 = ~n41836 & ~n41839;
  assign n41841 = ~n41740 & ~n41839;
  assign n41842 = ~n41836 & n41841;
  assign n41843 = ~n41740 & n41840;
  assign n41844 = pi223 & pi1140;
  assign n41845 = ~pi299 & ~n41844;
  assign n41846 = ~pi921 & n38636;
  assign n41847 = ~pi1140 & ~n38636;
  assign n41848 = pi222 & ~n41847;
  assign n41849 = pi222 & ~n41846;
  assign n41850 = ~n41847 & n41849;
  assign n41851 = ~n41846 & n41848;
  assign n41852 = pi224 & pi282;
  assign n41853 = ~pi222 & ~n41852;
  assign n41854 = pi869 & n41340;
  assign n41855 = ~pi224 & ~n41854;
  assign n41856 = n41853 & ~n41855;
  assign n41857 = ~n60730 & ~n41856;
  assign n41858 = ~n41340 & n41853;
  assign n41859 = n41857 & ~n41858;
  assign n41860 = ~pi223 & ~n41859;
  assign n41861 = n41845 & ~n41860;
  assign n41862 = ~pi39 & ~n41861;
  assign n41863 = pi215 & pi1140;
  assign n41864 = pi299 & ~n41863;
  assign n41865 = ~pi921 & n38221;
  assign n41866 = ~pi1140 & ~n38221;
  assign n41867 = pi221 & ~n41866;
  assign n41868 = pi221 & ~n41865;
  assign n41869 = ~n41866 & n41868;
  assign n41870 = ~n41865 & n41867;
  assign n41871 = pi216 & pi282;
  assign n41872 = ~pi221 & ~n41871;
  assign n41873 = ~pi869 & n41335;
  assign n41874 = ~pi170 & ~n41873;
  assign n41875 = pi869 & ~n40748;
  assign n41876 = ~pi869 & ~n41346;
  assign n41877 = pi170 & ~n41876;
  assign n41878 = ~n41875 & n41877;
  assign n41879 = ~n41874 & ~n41878;
  assign n41880 = ~pi228 & ~n41879;
  assign n41881 = pi869 & ~n28313;
  assign n41882 = pi105 & ~n41881;
  assign n41883 = ~pi105 & pi170;
  assign n41884 = pi228 & ~n41883;
  assign n41885 = ~n41882 & n41884;
  assign n41886 = ~pi216 & ~n41885;
  assign n41887 = ~n41628 & n41886;
  assign n41888 = ~n41880 & n41887;
  assign n41889 = n41872 & ~n41888;
  assign n41890 = ~n60731 & ~n41889;
  assign n41891 = ~pi215 & ~n41890;
  assign n41892 = n41864 & ~n41891;
  assign n41893 = n41862 & ~n41892;
  assign n41894 = ~pi224 & ~n41881;
  assign n41895 = n41853 & ~n41894;
  assign n41896 = ~n60730 & ~n41895;
  assign n41897 = ~pi223 & ~n41896;
  assign n41898 = ~n41844 & ~n41897;
  assign n41899 = ~pi299 & ~n41898;
  assign n41900 = ~n60722 & ~n41899;
  assign n41901 = ~pi869 & n58822;
  assign n41902 = ~pi228 & ~n41197;
  assign n41903 = ~pi228 & ~n41901;
  assign n41904 = ~n41197 & n41903;
  assign n41905 = ~n41901 & n41902;
  assign n41906 = ~n41403 & n41886;
  assign n41907 = ~n60732 & n41906;
  assign n41908 = n41872 & ~n41907;
  assign n41909 = ~n60731 & ~n41908;
  assign n41910 = ~pi215 & ~n41909;
  assign n41911 = ~n41863 & ~n41910;
  assign n41912 = pi299 & ~n41911;
  assign n41913 = n41900 & ~n41912;
  assign n41914 = pi39 & ~n41913;
  assign n41915 = ~pi38 & ~n41914;
  assign n41916 = ~n41893 & n41915;
  assign n41917 = ~pi170 & ~pi228;
  assign n41918 = n41886 & ~n41917;
  assign n41919 = n41872 & ~n41918;
  assign n41920 = ~n60731 & ~n41919;
  assign n41921 = ~pi215 & ~n41920;
  assign n41922 = ~n41863 & ~n41921;
  assign n41923 = n41673 & ~n41871;
  assign n41924 = n41922 & ~n41923;
  assign n41925 = pi299 & ~n41924;
  assign n41926 = n41900 & ~n41925;
  assign n41927 = pi38 & n41926;
  assign n41928 = ~pi100 & ~n41927;
  assign n41929 = ~n41916 & n41928;
  assign n41930 = pi170 & ~n41439;
  assign n41931 = ~pi869 & n41439;
  assign n41932 = ~pi228 & ~n41931;
  assign n41933 = ~pi228 & ~n41930;
  assign n41934 = ~n41931 & n41933;
  assign n41935 = ~n41930 & n41932;
  assign n41936 = n41906 & ~n60733;
  assign n41937 = n41872 & ~n41936;
  assign n41938 = ~n60731 & ~n41937;
  assign n41939 = ~pi215 & ~n41938;
  assign n41940 = ~n41863 & ~n41939;
  assign n41941 = pi299 & ~n41940;
  assign n41942 = n2634 & n41900;
  assign n41943 = ~n41941 & n41942;
  assign n41944 = ~n2634 & n41926;
  assign n41945 = pi100 & ~n41944;
  assign n41946 = ~n41943 & n41945;
  assign n41947 = ~n41929 & ~n41946;
  assign n41948 = ~pi87 & ~n41947;
  assign n41949 = ~n58815 & n41926;
  assign n41950 = n58815 & n41913;
  assign n41951 = ~n41949 & ~n41950;
  assign n41952 = pi87 & n41951;
  assign n41953 = ~pi75 & ~n41952;
  assign n41954 = ~n41948 & n41953;
  assign n41955 = pi75 & n41926;
  assign n41956 = ~pi92 & ~n41955;
  assign n41957 = ~n41954 & n41956;
  assign n41958 = n6309 & ~n41951;
  assign n41959 = ~n6309 & n41926;
  assign n41960 = pi92 & ~n41959;
  assign n41961 = ~n41958 & n41960;
  assign n41962 = n6306 & ~n41961;
  assign n41963 = ~n41957 & n41962;
  assign n41964 = ~n6306 & n41926;
  assign n41965 = ~pi55 & ~n41964;
  assign n41966 = ~n41963 & n41965;
  assign n41967 = n28288 & n41911;
  assign n41968 = ~n28288 & n41924;
  assign n41969 = pi55 & ~n41968;
  assign n41970 = ~n41967 & n41969;
  assign n41971 = ~pi56 & ~n41970;
  assign n41972 = ~n41966 & n41971;
  assign n41973 = n60070 & ~n41911;
  assign n41974 = ~n60070 & ~n41924;
  assign n41975 = pi56 & ~n41974;
  assign n41976 = ~pi55 & n41967;
  assign n41977 = ~n60070 & n41924;
  assign n41978 = ~n41976 & ~n41977;
  assign n41979 = pi56 & ~n41978;
  assign n41980 = ~n41973 & n41975;
  assign n41981 = ~pi62 & ~n60734;
  assign n41982 = ~n41972 & n41981;
  assign n41983 = n41492 & n41911;
  assign n41984 = ~n41492 & n41924;
  assign n41985 = pi62 & ~n41984;
  assign n41986 = ~n41983 & n41985;
  assign n41987 = pi248 & n4438;
  assign n41988 = ~n41986 & n41987;
  assign n41989 = ~n41982 & n41988;
  assign n41990 = ~pi869 & n40747;
  assign n41991 = ~n31400 & ~n41854;
  assign n41992 = ~n41990 & n41991;
  assign n41993 = ~pi869 & n40748;
  assign n41994 = pi869 & n41346;
  assign n41995 = ~pi170 & ~n41994;
  assign n41996 = ~n41993 & n41995;
  assign n41997 = ~pi170 & ~n41992;
  assign n41998 = pi170 & pi869;
  assign n41999 = n41335 & n41998;
  assign n42000 = pi170 & n41335;
  assign n42001 = ~n41995 & ~n42000;
  assign n42002 = pi869 & ~n42001;
  assign n42003 = ~n40748 & n41995;
  assign n42004 = ~n42002 & ~n42003;
  assign n42005 = ~n60735 & ~n41999;
  assign n42006 = ~pi228 & ~n60736;
  assign n42007 = ~n41356 & n41885;
  assign n42008 = ~pi216 & ~n42007;
  assign n42009 = ~n42006 & n42008;
  assign n42010 = n41872 & ~n42009;
  assign n42011 = ~n60731 & ~n42010;
  assign n42012 = ~pi215 & ~n42011;
  assign n42013 = n41864 & ~n42012;
  assign n42014 = n41845 & n41857;
  assign n42015 = n41862 & ~n42014;
  assign n42016 = ~n42013 & n42015;
  assign n42017 = n41886 & ~n60732;
  assign n42018 = n41872 & ~n42017;
  assign n42019 = ~n60731 & ~n42018;
  assign n42020 = ~pi215 & ~n42019;
  assign n42021 = ~n41863 & ~n42020;
  assign n42022 = pi299 & ~n42021;
  assign n42023 = ~n41899 & ~n42022;
  assign n42024 = pi39 & ~n42023;
  assign n42025 = ~pi38 & ~n42024;
  assign n42026 = ~n42016 & n42025;
  assign n42027 = pi299 & ~n41922;
  assign n42028 = ~n41899 & ~n42027;
  assign n42029 = pi38 & n42028;
  assign n42030 = ~pi100 & ~n42029;
  assign n42031 = ~n42026 & n42030;
  assign n42032 = n41886 & ~n60733;
  assign n42033 = n41872 & ~n42032;
  assign n42034 = ~n60731 & ~n42033;
  assign n42035 = ~pi215 & ~n42034;
  assign n42036 = ~n41863 & ~n42035;
  assign n42037 = pi299 & ~n42036;
  assign n42038 = n2634 & ~n41899;
  assign n42039 = ~n42037 & n42038;
  assign n42040 = ~n2634 & n42028;
  assign n42041 = pi100 & ~n42040;
  assign n42042 = ~n42039 & n42041;
  assign n42043 = ~n42031 & ~n42042;
  assign n42044 = ~pi87 & ~n42043;
  assign n42045 = ~n58815 & n42028;
  assign n42046 = n58815 & n42023;
  assign n42047 = ~n42045 & ~n42046;
  assign n42048 = pi87 & n42047;
  assign n42049 = ~pi75 & ~n42048;
  assign n42050 = ~n42044 & n42049;
  assign n42051 = pi75 & n42028;
  assign n42052 = ~pi92 & ~n42051;
  assign n42053 = ~n42050 & n42052;
  assign n42054 = n6309 & ~n42047;
  assign n42055 = ~n6309 & n42028;
  assign n42056 = pi92 & ~n42055;
  assign n42057 = ~n42054 & n42056;
  assign n42058 = n6306 & ~n42057;
  assign n42059 = ~n42053 & n42058;
  assign n42060 = ~n6306 & n42028;
  assign n42061 = ~pi55 & ~n42060;
  assign n42062 = ~n42059 & n42061;
  assign n42063 = n28288 & n42021;
  assign n42064 = ~n28288 & n41922;
  assign n42065 = pi55 & ~n42064;
  assign n42066 = ~n42063 & n42065;
  assign n42067 = ~pi56 & ~n42066;
  assign n42068 = ~n42062 & n42067;
  assign n42069 = n60070 & ~n42021;
  assign n42070 = ~n60070 & ~n41922;
  assign n42071 = pi56 & ~n42070;
  assign n42072 = ~n60070 & n41922;
  assign n42073 = ~pi55 & n42063;
  assign n42074 = ~n42072 & ~n42073;
  assign n42075 = pi56 & ~n42074;
  assign n42076 = ~n42069 & n42071;
  assign n42077 = ~pi62 & ~n60737;
  assign n42078 = ~n42068 & n42077;
  assign n42079 = n41492 & n42021;
  assign n42080 = ~n41492 & n41922;
  assign n42081 = pi62 & ~n42080;
  assign n42082 = ~n42079 & n42081;
  assign n42083 = ~pi248 & n4438;
  assign n42084 = ~n42082 & n42083;
  assign n42085 = ~n42078 & n42084;
  assign n42086 = pi248 & n41923;
  assign n42087 = ~n4438 & ~n42086;
  assign n42088 = n41922 & n42087;
  assign n42089 = ~n42085 & ~n42088;
  assign n42090 = ~n41989 & ~n42088;
  assign n42091 = ~n42085 & n42090;
  assign n42092 = ~n41989 & n42089;
  assign n42093 = pi216 & ~pi1139;
  assign n42094 = pi833 & pi920;
  assign n42095 = ~pi833 & pi1139;
  assign n42096 = ~pi216 & ~n42095;
  assign n42097 = ~pi216 & ~n42094;
  assign n42098 = ~n42095 & n42097;
  assign n42099 = ~n42094 & n42096;
  assign n42100 = pi221 & ~n60739;
  assign n42101 = ~n42093 & n42100;
  assign n42102 = pi216 & pi281;
  assign n42103 = ~pi221 & ~n42102;
  assign n42104 = ~pi216 & ~pi862;
  assign n42105 = ~n28313 & n38211;
  assign n42106 = ~n31586 & ~n42105;
  assign n42107 = n42104 & ~n42106;
  assign n42108 = n42103 & ~n42107;
  assign n42109 = ~n42101 & ~n42108;
  assign n42110 = ~n41441 & ~n42105;
  assign n42111 = n42103 & n42110;
  assign n42112 = n42109 & ~n42111;
  assign n42113 = pi148 & ~pi215;
  assign n42114 = ~pi216 & ~n42101;
  assign n42115 = ~pi216 & ~n42100;
  assign n42116 = n42110 & n60740;
  assign n42117 = n42113 & ~n42116;
  assign n42118 = ~n42112 & n42117;
  assign n42119 = pi215 & pi1139;
  assign n42120 = ~pi148 & ~pi215;
  assign n42121 = ~n31586 & ~n38211;
  assign n42122 = pi862 & ~n41403;
  assign n42123 = ~pi216 & ~n42122;
  assign n42124 = ~n42121 & n42123;
  assign n42125 = n42103 & ~n42124;
  assign n42126 = ~n42101 & ~n42125;
  assign n42127 = ~n38211 & ~n41441;
  assign n42128 = n42103 & n42127;
  assign n42129 = n42126 & ~n42128;
  assign n42130 = n42120 & ~n42129;
  assign n42131 = ~n42119 & ~n42130;
  assign n42132 = ~n42118 & n42131;
  assign n42133 = pi299 & ~n42132;
  assign n42134 = ~pi920 & n38636;
  assign n42135 = ~pi1139 & ~n38636;
  assign n42136 = pi222 & ~n42135;
  assign n42137 = pi222 & ~n42134;
  assign n42138 = ~n42135 & n42137;
  assign n42139 = ~n42134 & n42136;
  assign n42140 = pi223 & pi1139;
  assign n42141 = ~pi224 & ~n42140;
  assign n42142 = ~n60741 & n42141;
  assign n42143 = n28313 & n42142;
  assign n42144 = ~pi862 & n42142;
  assign n42145 = pi224 & pi281;
  assign n42146 = ~pi222 & ~n42145;
  assign n42147 = ~n60741 & ~n42146;
  assign n42148 = ~pi223 & ~n42147;
  assign n42149 = ~n42140 & ~n42148;
  assign n42150 = ~pi299 & ~n42149;
  assign n42151 = ~n42144 & n42150;
  assign n42152 = ~n42143 & n42151;
  assign n42153 = n2634 & ~n42152;
  assign n42154 = ~n42133 & n42153;
  assign n42155 = n42104 & n42105;
  assign n42156 = n42103 & ~n42155;
  assign n42157 = ~n42101 & ~n42156;
  assign n42158 = pi148 & ~n38211;
  assign n42159 = n60740 & n42158;
  assign n42160 = ~pi215 & ~n42159;
  assign n42161 = ~n42157 & n42160;
  assign n42162 = ~n42119 & ~n42161;
  assign n42163 = ~n41418 & ~n42162;
  assign n42164 = pi299 & n42163;
  assign n42165 = ~n42152 & ~n42164;
  assign n42166 = ~n2634 & n42165;
  assign n42167 = pi100 & ~n42166;
  assign n42168 = ~n42154 & n42167;
  assign n42169 = ~pi228 & n40748;
  assign n42170 = ~n38211 & ~n42169;
  assign n42171 = ~pi862 & n42170;
  assign n42172 = pi228 & ~n41356;
  assign n42173 = ~pi228 & ~n41346;
  assign n42174 = ~n42172 & ~n42173;
  assign n42175 = pi862 & ~n42174;
  assign n42176 = ~pi216 & ~n42175;
  assign n42177 = ~n42171 & n42176;
  assign n42178 = n42103 & ~n42177;
  assign n42179 = ~n42101 & ~n42178;
  assign n42180 = n42120 & ~n42179;
  assign n42181 = ~pi228 & n41335;
  assign n42182 = n38211 & n41340;
  assign n42183 = ~n42181 & ~n42182;
  assign n42184 = n42104 & ~n42183;
  assign n42185 = n42103 & ~n42184;
  assign n42186 = ~n42101 & ~n42185;
  assign n42187 = n60740 & n42183;
  assign n42188 = n42113 & ~n42187;
  assign n42189 = ~n42186 & n42188;
  assign n42190 = pi299 & ~n42119;
  assign n42191 = ~n42189 & n42190;
  assign n42192 = ~n42180 & n42191;
  assign n42193 = ~n41340 & n42142;
  assign n42194 = ~n42144 & ~n42149;
  assign n42195 = ~n42193 & n42194;
  assign n42196 = ~pi299 & ~n42195;
  assign n42197 = ~pi39 & ~n42196;
  assign n42198 = ~n42192 & n42197;
  assign n42199 = n42120 & ~n42126;
  assign n42200 = n42106 & n60740;
  assign n42201 = n42113 & ~n42200;
  assign n42202 = ~n42109 & n42113;
  assign n42203 = ~n42200 & n42202;
  assign n42204 = ~n42109 & n42201;
  assign n42205 = ~n42119 & ~n60742;
  assign n42206 = ~n42199 & n42205;
  assign n42207 = pi299 & ~n42206;
  assign n42208 = ~n42152 & ~n42207;
  assign n42209 = pi39 & ~n42208;
  assign n42210 = ~pi38 & ~n42209;
  assign n42211 = ~n42198 & n42210;
  assign n42212 = pi38 & n42165;
  assign n42213 = ~pi100 & ~n42212;
  assign n42214 = ~n42211 & n42213;
  assign n42215 = ~n42168 & ~n42214;
  assign n42216 = ~pi87 & ~n42215;
  assign n42217 = ~n58815 & n42165;
  assign n42218 = n58815 & n42208;
  assign n42219 = ~n42217 & ~n42218;
  assign n42220 = pi87 & n42219;
  assign n42221 = ~pi75 & ~n42220;
  assign n42222 = ~n42216 & n42221;
  assign n42223 = pi75 & n42165;
  assign n42224 = ~pi92 & ~n42223;
  assign n42225 = ~n42222 & n42224;
  assign n42226 = n6309 & ~n42219;
  assign n42227 = ~n6309 & n42165;
  assign n42228 = pi92 & ~n42227;
  assign n42229 = ~n42226 & n42228;
  assign n42230 = n6306 & ~n42229;
  assign n42231 = ~n42225 & n42230;
  assign n42232 = ~n6306 & n42165;
  assign n42233 = ~pi55 & ~n42232;
  assign n42234 = ~n42231 & n42233;
  assign n42235 = n28288 & n42206;
  assign n42236 = ~n28288 & ~n42163;
  assign n42237 = pi55 & ~n42236;
  assign n42238 = ~n42235 & n42237;
  assign n42239 = ~pi56 & ~n42238;
  assign n42240 = ~n42234 & n42239;
  assign n42241 = n60070 & ~n42206;
  assign n42242 = ~n60070 & n42163;
  assign n42243 = pi56 & ~n42242;
  assign n42244 = ~n60070 & ~n42163;
  assign n42245 = ~pi55 & n42235;
  assign n42246 = ~n42244 & ~n42245;
  assign n42247 = pi56 & ~n42246;
  assign n42248 = ~n42241 & n42243;
  assign n42249 = ~pi62 & ~n60743;
  assign n42250 = ~n42240 & n42249;
  assign n42251 = n41492 & n42206;
  assign n42252 = ~n41492 & ~n42163;
  assign n42253 = pi62 & ~n42252;
  assign n42254 = ~n42251 & n42253;
  assign n42255 = n4438 & ~n42254;
  assign n42256 = ~n42250 & n42255;
  assign n42257 = ~n4438 & ~n42163;
  assign n42258 = ~pi247 & ~n42257;
  assign n42259 = ~n42256 & n42258;
  assign n42260 = ~n42112 & n42120;
  assign n42261 = n60740 & n42127;
  assign n42262 = n42202 & ~n42261;
  assign n42263 = ~n42119 & ~n42262;
  assign n42264 = ~n42260 & n42263;
  assign n42265 = pi299 & ~n42264;
  assign n42266 = ~n60722 & ~n42151;
  assign n42267 = n2634 & n42266;
  assign n42268 = ~n42265 & n42267;
  assign n42269 = pi299 & ~n42162;
  assign n42270 = n42266 & ~n42269;
  assign n42271 = ~n2634 & n42270;
  assign n42272 = pi100 & ~n42271;
  assign n42273 = ~n42268 & n42272;
  assign n42274 = n41340 & n42144;
  assign n42275 = n42150 & ~n42274;
  assign n42276 = pi862 & ~n42170;
  assign n42277 = ~pi862 & n42174;
  assign n42278 = ~pi216 & ~n42277;
  assign n42279 = ~n42276 & n42278;
  assign n42280 = n42103 & ~n42279;
  assign n42281 = ~n42101 & ~n42280;
  assign n42282 = n42113 & ~n42281;
  assign n42283 = n42120 & ~n42186;
  assign n42284 = ~n42119 & ~n42283;
  assign n42285 = ~n42282 & n42284;
  assign n42286 = pi299 & ~n42285;
  assign n42287 = ~n42275 & ~n42286;
  assign n42288 = ~pi39 & ~n42287;
  assign n42289 = ~n42109 & n42160;
  assign n42290 = n42205 & ~n42289;
  assign n42291 = pi299 & ~n42290;
  assign n42292 = n42266 & ~n42291;
  assign n42293 = pi39 & ~n42292;
  assign n42294 = ~pi38 & ~n42293;
  assign n42295 = ~n42288 & n42294;
  assign n42296 = pi38 & n42270;
  assign n42297 = ~pi100 & ~n42296;
  assign n42298 = ~n42295 & n42297;
  assign n42299 = ~n42273 & ~n42298;
  assign n42300 = ~pi87 & ~n42299;
  assign n42301 = ~n58815 & n42270;
  assign n42302 = n58815 & n42292;
  assign n42303 = ~n42301 & ~n42302;
  assign n42304 = pi87 & n42303;
  assign n42305 = ~pi75 & ~n42304;
  assign n42306 = ~n42300 & n42305;
  assign n42307 = pi75 & n42270;
  assign n42308 = ~pi92 & ~n42307;
  assign n42309 = ~n42306 & n42308;
  assign n42310 = n6309 & ~n42303;
  assign n42311 = ~n6309 & n42270;
  assign n42312 = pi92 & ~n42311;
  assign n42313 = ~n42310 & n42312;
  assign n42314 = n6306 & ~n42313;
  assign n42315 = ~n42309 & n42314;
  assign n42316 = ~n6306 & n42270;
  assign n42317 = ~pi55 & ~n42316;
  assign n42318 = ~n42315 & n42317;
  assign n42319 = n28288 & n42290;
  assign n42320 = ~n28288 & n42162;
  assign n42321 = pi55 & ~n42320;
  assign n42322 = ~n42319 & n42321;
  assign n42323 = ~pi56 & ~n42322;
  assign n42324 = ~n42318 & n42323;
  assign n42325 = n60070 & ~n42290;
  assign n42326 = ~n60070 & ~n42162;
  assign n42327 = pi56 & ~n42326;
  assign n42328 = ~n60070 & n42162;
  assign n42329 = ~pi55 & n42319;
  assign n42330 = ~n42328 & ~n42329;
  assign n42331 = pi56 & ~n42330;
  assign n42332 = ~n42325 & n42327;
  assign n42333 = ~pi62 & ~n60744;
  assign n42334 = ~n42324 & n42333;
  assign n42335 = n41492 & n42290;
  assign n42336 = ~n41492 & n42162;
  assign n42337 = pi62 & ~n42336;
  assign n42338 = ~n42335 & n42337;
  assign n42339 = n4438 & ~n42338;
  assign n42340 = ~n42334 & n42339;
  assign n42341 = ~n4438 & n42162;
  assign n42342 = pi247 & ~n42341;
  assign n42343 = ~n42340 & n42342;
  assign n42344 = ~n42259 & ~n42343;
  assign n42345 = pi223 & pi1138;
  assign n42346 = ~pi299 & ~n42345;
  assign n42347 = ~pi940 & n38636;
  assign n42348 = ~pi1138 & ~n38636;
  assign n42349 = pi222 & ~n42348;
  assign n42350 = pi222 & ~n42347;
  assign n42351 = ~n42348 & n42350;
  assign n42352 = ~n42347 & n42349;
  assign n42353 = pi224 & pi269;
  assign n42354 = ~pi222 & ~n42353;
  assign n42355 = pi877 & n41340;
  assign n42356 = ~pi224 & ~n42355;
  assign n42357 = n42354 & ~n42356;
  assign n42358 = ~n60745 & ~n42357;
  assign n42359 = ~n41340 & n42354;
  assign n42360 = n42358 & ~n42359;
  assign n42361 = ~pi223 & ~n42360;
  assign n42362 = n42346 & ~n42361;
  assign n42363 = ~pi39 & ~n42362;
  assign n42364 = pi215 & pi1138;
  assign n42365 = pi299 & ~n42364;
  assign n42366 = ~pi940 & n38221;
  assign n42367 = ~pi1138 & ~n38221;
  assign n42368 = pi221 & ~n42367;
  assign n42369 = pi221 & ~n42366;
  assign n42370 = ~n42367 & n42369;
  assign n42371 = ~n42366 & n42368;
  assign n42372 = pi216 & pi269;
  assign n42373 = ~pi221 & ~n42372;
  assign n42374 = ~pi877 & n41335;
  assign n42375 = ~pi169 & ~n42374;
  assign n42376 = pi877 & ~n40748;
  assign n42377 = ~pi877 & ~n41346;
  assign n42378 = pi169 & ~n42377;
  assign n42379 = ~n42376 & n42378;
  assign n42380 = ~n42375 & ~n42379;
  assign n42381 = ~pi228 & ~n42380;
  assign n42382 = pi877 & ~n28313;
  assign n42383 = pi105 & ~n42382;
  assign n42384 = ~pi105 & pi169;
  assign n42385 = pi228 & ~n42384;
  assign n42386 = ~n42383 & n42385;
  assign n42387 = ~pi216 & ~n42386;
  assign n42388 = ~n41628 & n42387;
  assign n42389 = ~n42381 & n42388;
  assign n42390 = n42373 & ~n42389;
  assign n42391 = ~n60746 & ~n42390;
  assign n42392 = ~pi215 & ~n42391;
  assign n42393 = n42365 & ~n42392;
  assign n42394 = n42363 & ~n42393;
  assign n42395 = ~pi224 & ~n42382;
  assign n42396 = n42354 & ~n42395;
  assign n42397 = ~n60745 & ~n42396;
  assign n42398 = ~pi223 & ~n42397;
  assign n42399 = ~n42345 & ~n42398;
  assign n42400 = ~pi299 & ~n42399;
  assign n42401 = ~n60722 & ~n42400;
  assign n42402 = ~pi877 & n58822;
  assign n42403 = pi169 & ~n58822;
  assign n42404 = ~pi228 & ~n42403;
  assign n42405 = ~pi228 & ~n42402;
  assign n42406 = ~n42403 & n42405;
  assign n42407 = ~n42402 & n42404;
  assign n42408 = ~n41403 & n42387;
  assign n42409 = ~n60747 & n42408;
  assign n42410 = n42373 & ~n42409;
  assign n42411 = ~n60746 & ~n42410;
  assign n42412 = ~pi215 & ~n42411;
  assign n42413 = ~n42364 & ~n42412;
  assign n42414 = pi299 & ~n42413;
  assign n42415 = n42401 & ~n42414;
  assign n42416 = pi39 & ~n42415;
  assign n42417 = ~pi38 & ~n42416;
  assign n42418 = ~n42394 & n42417;
  assign n42419 = ~pi169 & ~pi228;
  assign n42420 = n42387 & ~n42419;
  assign n42421 = n42373 & ~n42420;
  assign n42422 = ~n60746 & ~n42421;
  assign n42423 = ~pi215 & ~n42422;
  assign n42424 = ~n42364 & ~n42423;
  assign n42425 = n41673 & ~n42372;
  assign n42426 = n42424 & ~n42425;
  assign n42427 = pi299 & ~n42426;
  assign n42428 = n42401 & ~n42427;
  assign n42429 = pi38 & n42428;
  assign n42430 = ~pi100 & ~n42429;
  assign n42431 = ~n42418 & n42430;
  assign n42432 = pi169 & ~n41439;
  assign n42433 = ~pi877 & n41439;
  assign n42434 = ~pi228 & ~n42433;
  assign n42435 = ~pi228 & ~n42432;
  assign n42436 = ~n42433 & n42435;
  assign n42437 = ~n42432 & n42434;
  assign n42438 = n42408 & ~n60748;
  assign n42439 = n42373 & ~n42438;
  assign n42440 = ~n60746 & ~n42439;
  assign n42441 = ~pi215 & ~n42440;
  assign n42442 = ~n42364 & ~n42441;
  assign n42443 = pi299 & ~n42442;
  assign n42444 = n2634 & n42401;
  assign n42445 = ~n42443 & n42444;
  assign n42446 = ~n2634 & n42428;
  assign n42447 = pi100 & ~n42446;
  assign n42448 = ~n42445 & n42447;
  assign n42449 = ~n42431 & ~n42448;
  assign n42450 = ~pi87 & ~n42449;
  assign n42451 = ~n58815 & n42428;
  assign n42452 = n58815 & n42415;
  assign n42453 = ~n42451 & ~n42452;
  assign n42454 = pi87 & n42453;
  assign n42455 = ~pi75 & ~n42454;
  assign n42456 = ~n42450 & n42455;
  assign n42457 = pi75 & n42428;
  assign n42458 = ~pi92 & ~n42457;
  assign n42459 = ~n42456 & n42458;
  assign n42460 = n6309 & ~n42453;
  assign n42461 = ~n6309 & n42428;
  assign n42462 = pi92 & ~n42461;
  assign n42463 = ~n42460 & n42462;
  assign n42464 = n6306 & ~n42463;
  assign n42465 = ~n42459 & n42464;
  assign n42466 = ~n6306 & n42428;
  assign n42467 = ~pi55 & ~n42466;
  assign n42468 = ~n42465 & n42467;
  assign n42469 = n28288 & n42413;
  assign n42470 = ~n28288 & n42426;
  assign n42471 = pi55 & ~n42470;
  assign n42472 = ~n42469 & n42471;
  assign n42473 = ~pi56 & ~n42472;
  assign n42474 = ~n42468 & n42473;
  assign n42475 = n60070 & ~n42413;
  assign n42476 = ~n60070 & ~n42426;
  assign n42477 = pi56 & ~n42476;
  assign n42478 = ~pi55 & n42469;
  assign n42479 = ~n60070 & n42426;
  assign n42480 = ~n42478 & ~n42479;
  assign n42481 = pi56 & ~n42480;
  assign n42482 = ~n42475 & n42477;
  assign n42483 = ~pi62 & ~n60749;
  assign n42484 = ~n42474 & n42483;
  assign n42485 = n41492 & n42413;
  assign n42486 = ~n41492 & n42426;
  assign n42487 = pi62 & ~n42486;
  assign n42488 = ~n42485 & n42487;
  assign n42489 = pi246 & n4438;
  assign n42490 = ~n42488 & n42489;
  assign n42491 = ~n42484 & n42490;
  assign n42492 = ~pi877 & n40747;
  assign n42493 = ~n31400 & ~n42355;
  assign n42494 = ~n42492 & n42493;
  assign n42495 = ~pi877 & n40748;
  assign n42496 = pi877 & n41346;
  assign n42497 = ~pi169 & ~n42496;
  assign n42498 = ~n42495 & n42497;
  assign n42499 = ~pi169 & ~n42494;
  assign n42500 = pi169 & pi877;
  assign n42501 = n41335 & n42500;
  assign n42502 = pi169 & n41335;
  assign n42503 = ~n42497 & ~n42502;
  assign n42504 = pi877 & ~n42503;
  assign n42505 = ~n40748 & n42497;
  assign n42506 = ~n42504 & ~n42505;
  assign n42507 = ~n60750 & ~n42501;
  assign n42508 = ~pi228 & ~n60751;
  assign n42509 = ~n41356 & n42386;
  assign n42510 = ~pi216 & ~n42509;
  assign n42511 = ~n42508 & n42510;
  assign n42512 = n42373 & ~n42511;
  assign n42513 = ~n60746 & ~n42512;
  assign n42514 = ~pi215 & ~n42513;
  assign n42515 = n42365 & ~n42514;
  assign n42516 = n42346 & n42358;
  assign n42517 = n42363 & ~n42516;
  assign n42518 = ~n42515 & n42517;
  assign n42519 = n42387 & ~n60747;
  assign n42520 = n42373 & ~n42519;
  assign n42521 = ~n60746 & ~n42520;
  assign n42522 = ~pi215 & ~n42521;
  assign n42523 = ~n42364 & ~n42522;
  assign n42524 = pi299 & ~n42523;
  assign n42525 = ~n42400 & ~n42524;
  assign n42526 = pi39 & ~n42525;
  assign n42527 = ~pi38 & ~n42526;
  assign n42528 = ~n42518 & n42527;
  assign n42529 = pi299 & ~n42424;
  assign n42530 = ~n42400 & ~n42529;
  assign n42531 = pi38 & n42530;
  assign n42532 = ~pi100 & ~n42531;
  assign n42533 = ~n42528 & n42532;
  assign n42534 = n42387 & ~n60748;
  assign n42535 = n42373 & ~n42534;
  assign n42536 = ~n60746 & ~n42535;
  assign n42537 = ~pi215 & ~n42536;
  assign n42538 = ~n42364 & ~n42537;
  assign n42539 = pi299 & ~n42538;
  assign n42540 = n2634 & ~n42400;
  assign n42541 = ~n42539 & n42540;
  assign n42542 = ~n2634 & n42530;
  assign n42543 = pi100 & ~n42542;
  assign n42544 = ~n42541 & n42543;
  assign n42545 = ~n42533 & ~n42544;
  assign n42546 = ~pi87 & ~n42545;
  assign n42547 = ~n58815 & n42530;
  assign n42548 = n58815 & n42525;
  assign n42549 = ~n42547 & ~n42548;
  assign n42550 = pi87 & n42549;
  assign n42551 = ~pi75 & ~n42550;
  assign n42552 = ~n42546 & n42551;
  assign n42553 = pi75 & n42530;
  assign n42554 = ~pi92 & ~n42553;
  assign n42555 = ~n42552 & n42554;
  assign n42556 = n6309 & ~n42549;
  assign n42557 = ~n6309 & n42530;
  assign n42558 = pi92 & ~n42557;
  assign n42559 = ~n42556 & n42558;
  assign n42560 = n6306 & ~n42559;
  assign n42561 = ~n42555 & n42560;
  assign n42562 = ~n6306 & n42530;
  assign n42563 = ~pi55 & ~n42562;
  assign n42564 = ~n42561 & n42563;
  assign n42565 = n28288 & n42523;
  assign n42566 = ~n28288 & n42424;
  assign n42567 = pi55 & ~n42566;
  assign n42568 = ~n42565 & n42567;
  assign n42569 = ~pi56 & ~n42568;
  assign n42570 = ~n42564 & n42569;
  assign n42571 = n60070 & ~n42523;
  assign n42572 = ~n60070 & ~n42424;
  assign n42573 = pi56 & ~n42572;
  assign n42574 = ~n60070 & n42424;
  assign n42575 = ~pi55 & n42565;
  assign n42576 = ~n42574 & ~n42575;
  assign n42577 = pi56 & ~n42576;
  assign n42578 = ~n42571 & n42573;
  assign n42579 = ~pi62 & ~n60752;
  assign n42580 = ~n42570 & n42579;
  assign n42581 = n41492 & n42523;
  assign n42582 = ~n41492 & n42424;
  assign n42583 = pi62 & ~n42582;
  assign n42584 = ~n42581 & n42583;
  assign n42585 = ~pi246 & n4438;
  assign n42586 = ~n42584 & n42585;
  assign n42587 = ~n42580 & n42586;
  assign n42588 = pi246 & n42425;
  assign n42589 = ~n4438 & ~n42588;
  assign n42590 = n42424 & n42589;
  assign n42591 = ~n42587 & ~n42590;
  assign n42592 = ~n42491 & ~n42590;
  assign n42593 = ~n42587 & n42592;
  assign n42594 = ~n42491 & n42591;
  assign n42595 = pi223 & pi1137;
  assign n42596 = ~pi299 & ~n42595;
  assign n42597 = ~pi933 & n38636;
  assign n42598 = ~pi1137 & ~n38636;
  assign n42599 = pi222 & ~n42598;
  assign n42600 = pi222 & ~n42597;
  assign n42601 = ~n42598 & n42600;
  assign n42602 = ~n42597 & n42599;
  assign n42603 = pi224 & pi280;
  assign n42604 = ~pi222 & ~n42603;
  assign n42605 = pi878 & n41340;
  assign n42606 = ~pi224 & ~n42605;
  assign n42607 = n42604 & ~n42606;
  assign n42608 = ~n60754 & ~n42607;
  assign n42609 = ~n41340 & n42604;
  assign n42610 = n42608 & ~n42609;
  assign n42611 = ~pi223 & ~n42610;
  assign n42612 = n42596 & ~n42611;
  assign n42613 = ~pi39 & ~n42612;
  assign n42614 = pi215 & pi1137;
  assign n42615 = pi299 & ~n42614;
  assign n42616 = ~pi933 & n38221;
  assign n42617 = ~pi1137 & ~n38221;
  assign n42618 = pi221 & ~n42617;
  assign n42619 = pi221 & ~n42616;
  assign n42620 = ~n42617 & n42619;
  assign n42621 = ~n42616 & n42618;
  assign n42622 = pi216 & pi280;
  assign n42623 = ~pi221 & ~n42622;
  assign n42624 = ~pi878 & n41335;
  assign n42625 = ~pi168 & ~n42624;
  assign n42626 = pi878 & ~n40748;
  assign n42627 = ~pi878 & ~n41346;
  assign n42628 = pi168 & ~n42627;
  assign n42629 = ~n42626 & n42628;
  assign n42630 = ~n42625 & ~n42629;
  assign n42631 = ~pi228 & ~n42630;
  assign n42632 = pi878 & ~n28313;
  assign n42633 = pi105 & ~n42632;
  assign n42634 = ~pi105 & pi168;
  assign n42635 = pi228 & ~n42634;
  assign n42636 = ~n42633 & n42635;
  assign n42637 = ~pi216 & ~n42636;
  assign n42638 = ~n41628 & n42637;
  assign n42639 = ~n42631 & n42638;
  assign n42640 = n42623 & ~n42639;
  assign n42641 = ~n60755 & ~n42640;
  assign n42642 = ~pi215 & ~n42641;
  assign n42643 = n42615 & ~n42642;
  assign n42644 = n42613 & ~n42643;
  assign n42645 = ~pi224 & ~n42632;
  assign n42646 = n42604 & ~n42645;
  assign n42647 = ~n60754 & ~n42646;
  assign n42648 = ~pi223 & ~n42647;
  assign n42649 = ~n42595 & ~n42648;
  assign n42650 = ~pi299 & ~n42649;
  assign n42651 = ~n60722 & ~n42650;
  assign n42652 = pi168 & ~n58822;
  assign n42653 = ~pi878 & n58822;
  assign n42654 = ~pi228 & ~n42653;
  assign n42655 = ~pi228 & ~n42652;
  assign n42656 = ~n42653 & n42655;
  assign n42657 = ~n42652 & n42654;
  assign n42658 = ~n41403 & n42637;
  assign n42659 = ~n60756 & n42658;
  assign n42660 = n42623 & ~n42659;
  assign n42661 = ~n60755 & ~n42660;
  assign n42662 = ~pi215 & ~n42661;
  assign n42663 = ~n42614 & ~n42662;
  assign n42664 = pi299 & ~n42663;
  assign n42665 = n42651 & ~n42664;
  assign n42666 = pi39 & ~n42665;
  assign n42667 = ~pi38 & ~n42666;
  assign n42668 = ~n42644 & n42667;
  assign n42669 = ~pi168 & ~pi228;
  assign n42670 = n42637 & ~n42669;
  assign n42671 = n42623 & ~n42670;
  assign n42672 = ~n60755 & ~n42671;
  assign n42673 = ~pi215 & ~n42672;
  assign n42674 = ~n42614 & ~n42673;
  assign n42675 = n41673 & ~n42622;
  assign n42676 = n42674 & ~n42675;
  assign n42677 = pi299 & ~n42676;
  assign n42678 = n42651 & ~n42677;
  assign n42679 = pi38 & n42678;
  assign n42680 = ~pi100 & ~n42679;
  assign n42681 = ~n42668 & n42680;
  assign n42682 = pi168 & ~n41439;
  assign n42683 = ~pi878 & n41439;
  assign n42684 = ~pi228 & ~n42683;
  assign n42685 = ~pi228 & ~n42682;
  assign n42686 = ~n42683 & n42685;
  assign n42687 = ~n42682 & n42684;
  assign n42688 = n42658 & ~n60757;
  assign n42689 = n42623 & ~n42688;
  assign n42690 = ~n60755 & ~n42689;
  assign n42691 = ~pi215 & ~n42690;
  assign n42692 = ~n42614 & ~n42691;
  assign n42693 = pi299 & ~n42692;
  assign n42694 = n2634 & n42651;
  assign n42695 = ~n42693 & n42694;
  assign n42696 = ~n2634 & n42678;
  assign n42697 = pi100 & ~n42696;
  assign n42698 = ~n42695 & n42697;
  assign n42699 = ~n42681 & ~n42698;
  assign n42700 = ~pi87 & ~n42699;
  assign n42701 = ~n58815 & n42678;
  assign n42702 = n58815 & n42665;
  assign n42703 = ~n42701 & ~n42702;
  assign n42704 = pi87 & n42703;
  assign n42705 = ~pi75 & ~n42704;
  assign n42706 = ~n42700 & n42705;
  assign n42707 = pi75 & n42678;
  assign n42708 = ~pi92 & ~n42707;
  assign n42709 = ~n42706 & n42708;
  assign n42710 = n6309 & ~n42703;
  assign n42711 = ~n6309 & n42678;
  assign n42712 = pi92 & ~n42711;
  assign n42713 = ~n42710 & n42712;
  assign n42714 = n6306 & ~n42713;
  assign n42715 = ~n42709 & n42714;
  assign n42716 = ~n6306 & n42678;
  assign n42717 = ~pi55 & ~n42716;
  assign n42718 = ~n42715 & n42717;
  assign n42719 = n28288 & n42663;
  assign n42720 = ~n28288 & n42676;
  assign n42721 = pi55 & ~n42720;
  assign n42722 = ~n42719 & n42721;
  assign n42723 = ~pi56 & ~n42722;
  assign n42724 = ~n42718 & n42723;
  assign n42725 = n60070 & ~n42663;
  assign n42726 = ~n60070 & ~n42676;
  assign n42727 = pi56 & ~n42726;
  assign n42728 = ~pi55 & n42719;
  assign n42729 = ~n60070 & n42676;
  assign n42730 = ~n42728 & ~n42729;
  assign n42731 = pi56 & ~n42730;
  assign n42732 = ~n42725 & n42727;
  assign n42733 = ~pi62 & ~n60758;
  assign n42734 = ~n42724 & n42733;
  assign n42735 = n41492 & n42663;
  assign n42736 = ~n41492 & n42676;
  assign n42737 = pi62 & ~n42736;
  assign n42738 = ~n42735 & n42737;
  assign n42739 = pi240 & n4438;
  assign n42740 = ~n42738 & n42739;
  assign n42741 = ~n42734 & n42740;
  assign n42742 = ~pi878 & n40747;
  assign n42743 = ~n31400 & ~n42605;
  assign n42744 = ~n42742 & n42743;
  assign n42745 = ~pi878 & n40748;
  assign n42746 = pi878 & n41346;
  assign n42747 = ~pi168 & ~n42746;
  assign n42748 = ~n42745 & n42747;
  assign n42749 = ~pi168 & ~n42744;
  assign n42750 = pi168 & pi878;
  assign n42751 = n41335 & n42750;
  assign n42752 = pi168 & n41335;
  assign n42753 = ~n42747 & ~n42752;
  assign n42754 = pi878 & ~n42753;
  assign n42755 = ~n40748 & n42747;
  assign n42756 = ~n42754 & ~n42755;
  assign n42757 = ~n60759 & ~n42751;
  assign n42758 = ~pi228 & ~n60760;
  assign n42759 = ~n41356 & n42636;
  assign n42760 = ~pi216 & ~n42759;
  assign n42761 = ~n42758 & n42760;
  assign n42762 = n42623 & ~n42761;
  assign n42763 = ~n60755 & ~n42762;
  assign n42764 = ~pi215 & ~n42763;
  assign n42765 = n42615 & ~n42764;
  assign n42766 = n42596 & n42608;
  assign n42767 = n42613 & ~n42766;
  assign n42768 = ~n42765 & n42767;
  assign n42769 = n42637 & ~n60756;
  assign n42770 = n42623 & ~n42769;
  assign n42771 = ~n60755 & ~n42770;
  assign n42772 = ~pi215 & ~n42771;
  assign n42773 = ~n42614 & ~n42772;
  assign n42774 = pi299 & ~n42773;
  assign n42775 = ~n42650 & ~n42774;
  assign n42776 = pi39 & ~n42775;
  assign n42777 = ~pi38 & ~n42776;
  assign n42778 = ~n42768 & n42777;
  assign n42779 = pi299 & ~n42674;
  assign n42780 = ~n42650 & ~n42779;
  assign n42781 = pi38 & n42780;
  assign n42782 = ~pi100 & ~n42781;
  assign n42783 = ~n42778 & n42782;
  assign n42784 = n42637 & ~n60757;
  assign n42785 = n42623 & ~n42784;
  assign n42786 = ~n60755 & ~n42785;
  assign n42787 = ~pi215 & ~n42786;
  assign n42788 = ~n42614 & ~n42787;
  assign n42789 = pi299 & ~n42788;
  assign n42790 = n2634 & ~n42650;
  assign n42791 = ~n42789 & n42790;
  assign n42792 = ~n2634 & n42780;
  assign n42793 = pi100 & ~n42792;
  assign n42794 = ~n42791 & n42793;
  assign n42795 = ~n42783 & ~n42794;
  assign n42796 = ~pi87 & ~n42795;
  assign n42797 = ~n58815 & n42780;
  assign n42798 = n58815 & n42775;
  assign n42799 = ~n42797 & ~n42798;
  assign n42800 = pi87 & n42799;
  assign n42801 = ~pi75 & ~n42800;
  assign n42802 = ~n42796 & n42801;
  assign n42803 = pi75 & n42780;
  assign n42804 = ~pi92 & ~n42803;
  assign n42805 = ~n42802 & n42804;
  assign n42806 = n6309 & ~n42799;
  assign n42807 = ~n6309 & n42780;
  assign n42808 = pi92 & ~n42807;
  assign n42809 = ~n42806 & n42808;
  assign n42810 = n6306 & ~n42809;
  assign n42811 = ~n42805 & n42810;
  assign n42812 = ~n6306 & n42780;
  assign n42813 = ~pi55 & ~n42812;
  assign n42814 = ~n42811 & n42813;
  assign n42815 = n28288 & n42773;
  assign n42816 = ~n28288 & n42674;
  assign n42817 = pi55 & ~n42816;
  assign n42818 = ~n42815 & n42817;
  assign n42819 = ~pi56 & ~n42818;
  assign n42820 = ~n42814 & n42819;
  assign n42821 = n60070 & ~n42773;
  assign n42822 = ~n60070 & ~n42674;
  assign n42823 = pi56 & ~n42822;
  assign n42824 = ~n60070 & n42674;
  assign n42825 = ~pi55 & n42815;
  assign n42826 = ~n42824 & ~n42825;
  assign n42827 = pi56 & ~n42826;
  assign n42828 = ~n42821 & n42823;
  assign n42829 = ~pi62 & ~n60761;
  assign n42830 = ~n42820 & n42829;
  assign n42831 = n41492 & n42773;
  assign n42832 = ~n41492 & n42674;
  assign n42833 = pi62 & ~n42832;
  assign n42834 = ~n42831 & n42833;
  assign n42835 = ~pi240 & n4438;
  assign n42836 = ~n42834 & n42835;
  assign n42837 = ~n42830 & n42836;
  assign n42838 = pi240 & n42675;
  assign n42839 = ~n4438 & ~n42838;
  assign n42840 = n42674 & n42839;
  assign n42841 = ~n42837 & ~n42840;
  assign n42842 = ~n42741 & ~n42840;
  assign n42843 = ~n42837 & n42842;
  assign n42844 = ~n42741 & n42841;
  assign n42845 = ~n60087 & ~n60122;
  assign n42846 = ~pi137 & ~n42845;
  assign n42847 = n28549 & ~n42846;
  assign n42848 = n31408 & ~n35574;
  assign n42849 = ~n38279 & n42848;
  assign n42850 = n31402 & ~n42849;
  assign n42851 = n31401 & ~n42850;
  assign n42852 = ~n38290 & ~n42851;
  assign n42853 = ~pi95 & ~n42852;
  assign n42854 = ~n31400 & ~n42853;
  assign n42855 = pi137 & ~n42854;
  assign n42856 = ~n60431 & n38371;
  assign n42857 = n38372 & ~n42856;
  assign n42858 = ~pi137 & ~n42857;
  assign n42859 = ~n42855 & ~n42858;
  assign n42860 = pi332 & ~n42859;
  assign n42861 = ~n31400 & ~n38292;
  assign n42862 = pi137 & ~n42861;
  assign n42863 = ~n38374 & ~n42862;
  assign n42864 = ~pi332 & ~n42863;
  assign n42865 = ~n42860 & ~n42864;
  assign n42866 = n28553 & n42865;
  assign n42867 = pi1093 & ~n42857;
  assign n42868 = n2757 & n38372;
  assign n42869 = n2618 & ~n38304;
  assign n42870 = ~pi32 & ~n42869;
  assign n42871 = n42868 & ~n42870;
  assign n42872 = ~pi1093 & ~n42871;
  assign n42873 = ~n2757 & n42857;
  assign n42874 = n60431 & n42868;
  assign n42875 = ~n42873 & ~n42874;
  assign n42876 = n42872 & n42875;
  assign n42877 = ~n42867 & ~n42876;
  assign n42878 = n37845 & ~n42877;
  assign n42879 = ~n2757 & n38373;
  assign n42880 = n42872 & ~n42879;
  assign n42881 = n2618 & ~n38336;
  assign n42882 = ~pi32 & ~n42881;
  assign n42883 = n42868 & ~n42882;
  assign n42884 = pi1093 & ~n42879;
  assign n42885 = ~n42883 & n42884;
  assign n42886 = ~n42880 & ~n42885;
  assign n42887 = n37803 & ~n42886;
  assign n42888 = n42875 & n42887;
  assign n42889 = ~n42878 & ~n42888;
  assign n42890 = ~n42855 & n42889;
  assign n42891 = pi332 & ~n42890;
  assign n42892 = pi1093 & ~n38373;
  assign n42893 = ~n42880 & ~n42892;
  assign n42894 = n37845 & ~n42893;
  assign n42895 = ~n42887 & ~n42894;
  assign n42896 = ~n42862 & n42895;
  assign n42897 = ~pi332 & ~n42896;
  assign n42898 = ~n42891 & ~n42897;
  assign n42899 = ~n28553 & n42898;
  assign n42900 = ~pi210 & ~n42899;
  assign n42901 = ~pi210 & ~n42866;
  assign n42902 = ~n42899 & n42901;
  assign n42903 = ~n42866 & n42900;
  assign n42904 = ~n31400 & ~n38320;
  assign n42905 = pi137 & ~n42904;
  assign n42906 = ~n38378 & ~n42905;
  assign n42907 = ~pi332 & ~n42906;
  assign n42908 = ~n38314 & ~n42851;
  assign n42909 = ~pi95 & ~n42908;
  assign n42910 = n38616 & ~n42909;
  assign n42911 = ~pi137 & n38315;
  assign n42912 = ~n42856 & n42911;
  assign n42913 = pi332 & ~n42912;
  assign n42914 = ~n42910 & n42913;
  assign n42915 = ~n42907 & ~n42914;
  assign n42916 = pi210 & ~n42915;
  assign n42917 = pi299 & ~n42916;
  assign n42918 = ~n60763 & n42917;
  assign n42919 = ~n28551 & n42898;
  assign n42920 = n28551 & n42865;
  assign n42921 = ~pi198 & ~n42920;
  assign n42922 = ~pi198 & ~n42919;
  assign n42923 = ~n42920 & n42922;
  assign n42924 = ~n42919 & n42921;
  assign n42925 = pi198 & ~n42915;
  assign n42926 = ~pi299 & ~n42925;
  assign n42927 = ~n60764 & n42926;
  assign n42928 = ~n42918 & ~n42927;
  assign n42929 = ~pi39 & ~n42928;
  assign n42930 = pi39 & n38230;
  assign n42931 = ~pi38 & ~n42930;
  assign n42932 = ~n42929 & n42931;
  assign n42933 = pi38 & ~pi137;
  assign n42934 = n31399 & ~n42933;
  assign n42935 = ~n42932 & n42934;
  assign n42936 = ~n42847 & ~n42935;
  assign n42937 = ~pi87 & ~n42936;
  assign n42938 = n58815 & n38230;
  assign n42939 = pi87 & n42938;
  assign n42940 = ~pi75 & ~n42939;
  assign n42941 = ~n42937 & n42940;
  assign n42942 = n28302 & ~n42846;
  assign n42943 = pi75 & ~n42942;
  assign n42944 = ~pi92 & ~n42943;
  assign n42945 = ~n42941 & n42944;
  assign n42946 = pi92 & n6309;
  assign n42947 = n42938 & n42946;
  assign n42948 = ~pi54 & ~n42947;
  assign n42949 = ~n42945 & n42948;
  assign n42950 = n6310 & n42938;
  assign n42951 = pi54 & ~n42950;
  assign n42952 = ~pi74 & ~n42951;
  assign n42953 = ~n42949 & n42952;
  assign n42954 = pi74 & n28299;
  assign n42955 = ~pi54 & pi74;
  assign n42956 = n42950 & n42955;
  assign n42957 = n42938 & n42954;
  assign n42958 = ~pi55 & ~n60765;
  assign n42959 = ~n42953 & n42958;
  assign n42960 = n28595 & ~n42959;
  assign n42961 = pi56 & n28283;
  assign n42962 = n42938 & n42961;
  assign n42963 = ~n42960 & ~n42962;
  assign n42964 = ~pi62 & ~n42963;
  assign n42965 = n31573 & n42938;
  assign n42966 = pi62 & n42965;
  assign n42967 = n4438 & ~n42966;
  assign n42968 = ~n42964 & n42967;
  assign n42969 = ~pi62 & n42965;
  assign n42970 = ~n4438 & ~n42969;
  assign n42971 = ~n28282 & ~n42970;
  assign po382 = ~n42968 & n42971;
  assign n42973 = ~pi939 & n38636;
  assign n42974 = ~pi1146 & ~n38636;
  assign n42975 = pi222 & ~n42974;
  assign n42976 = ~n42973 & n42975;
  assign n42977 = pi276 & n26651;
  assign n42978 = ~pi223 & ~n42977;
  assign n42979 = ~pi223 & ~n42976;
  assign n42980 = ~n42977 & n42979;
  assign n42981 = ~n42976 & n42978;
  assign n42982 = pi223 & ~pi1146;
  assign n42983 = ~pi299 & ~n42982;
  assign n42984 = ~n60766 & n42983;
  assign n42985 = ~pi939 & n38221;
  assign n42986 = ~pi1146 & ~n38221;
  assign n42987 = pi221 & ~n42986;
  assign n42988 = pi221 & ~n42985;
  assign n42989 = ~n42986 & n42988;
  assign n42990 = ~n42985 & n42987;
  assign n42991 = pi215 & pi1146;
  assign n42992 = ~pi216 & ~pi228;
  assign n42993 = ~n42991 & n42992;
  assign n42994 = ~n60767 & ~n42991;
  assign n42995 = n42992 & n42994;
  assign n42996 = ~n60767 & n42993;
  assign n42997 = ~pi216 & n31586;
  assign n42998 = n42994 & n42997;
  assign n42999 = n58822 & n60768;
  assign n43000 = pi276 & n37050;
  assign n43001 = ~pi216 & ~n38211;
  assign n43002 = ~n43000 & ~n43001;
  assign n43003 = ~pi221 & ~n43002;
  assign n43004 = ~n60767 & ~n43003;
  assign n43005 = ~pi215 & ~n43004;
  assign n43006 = ~n42991 & ~n43005;
  assign n43007 = pi299 & ~n43006;
  assign n43008 = ~n60769 & n43007;
  assign n43009 = ~n42984 & ~n43008;
  assign n43010 = ~pi154 & ~n43009;
  assign n43011 = ~n60767 & ~n43000;
  assign n43012 = ~pi215 & ~n43011;
  assign n43013 = ~n42991 & ~n43012;
  assign n43014 = pi299 & ~n43013;
  assign n43015 = ~n42984 & ~n43014;
  assign n43016 = pi154 & ~n43015;
  assign n43017 = n58815 & ~n43016;
  assign n43018 = ~n43010 & n43017;
  assign n43019 = pi154 & ~n43013;
  assign n43020 = ~pi154 & ~n43006;
  assign n43021 = ~n43019 & ~n43020;
  assign n43022 = pi299 & ~n43021;
  assign n43023 = ~n42984 & ~n43022;
  assign n43024 = ~n58815 & n43023;
  assign n43025 = ~n43018 & ~n43024;
  assign n43026 = pi87 & ~n43025;
  assign n43027 = n40750 & n60768;
  assign n43028 = n43007 & ~n43027;
  assign n43029 = ~n42984 & ~n43028;
  assign n43030 = ~pi154 & ~n43029;
  assign n43031 = ~pi38 & ~n43016;
  assign n43032 = ~n43030 & n43031;
  assign n43033 = pi38 & n43023;
  assign n43034 = ~pi100 & ~n43033;
  assign n43035 = ~n43032 & n43034;
  assign n43036 = n2634 & n31168;
  assign n43037 = ~pi38 & ~pi216;
  assign n43038 = ~pi228 & n43037;
  assign n43039 = ~pi39 & n31168;
  assign n43040 = n43038 & n43039;
  assign n43041 = n42994 & n43040;
  assign n43042 = n60768 & n43036;
  assign n43043 = n41439 & n60770;
  assign n43044 = pi100 & ~n43023;
  assign n43045 = ~n43043 & n43044;
  assign n43046 = ~pi87 & ~n43045;
  assign n43047 = ~n43035 & n43046;
  assign n43048 = ~n43026 & ~n43047;
  assign n43049 = ~pi75 & ~n43048;
  assign n43050 = pi75 & n43023;
  assign n43051 = ~pi92 & ~n43050;
  assign n43052 = ~n43049 & n43051;
  assign n43053 = n6309 & n43018;
  assign n43054 = ~n60069 & n43023;
  assign n43055 = pi92 & ~n43054;
  assign n43056 = ~n43053 & n43055;
  assign n43057 = n6306 & ~n43056;
  assign n43058 = ~n43052 & n43057;
  assign n43059 = ~n6306 & n43023;
  assign n43060 = ~pi55 & ~n43059;
  assign n43061 = ~n43058 & n43060;
  assign n43062 = n28288 & n60769;
  assign n43063 = pi55 & ~n43021;
  assign n43064 = ~n43062 & n43063;
  assign n43065 = ~pi56 & ~n43064;
  assign n43066 = ~n43061 & n43065;
  assign n43067 = n60070 & ~n43021;
  assign n43068 = ~n60769 & n43067;
  assign n43069 = ~n60070 & ~n43021;
  assign n43070 = pi56 & ~n43069;
  assign n43071 = ~n43068 & n43070;
  assign n43072 = ~pi62 & ~n43071;
  assign n43073 = ~n43066 & n43072;
  assign n43074 = ~n41492 & ~n43021;
  assign n43075 = ~n43068 & ~n43074;
  assign n43076 = pi62 & ~n43075;
  assign n43077 = n4438 & ~n43076;
  assign n43078 = ~n43073 & n43077;
  assign n43079 = ~n4438 & n43021;
  assign n43080 = ~pi239 & ~n43079;
  assign n43081 = ~n43078 & n43080;
  assign n43082 = ~pi154 & ~n42183;
  assign n43083 = pi154 & ~n42174;
  assign n43084 = n35591 & ~n43083;
  assign n43085 = ~n43082 & n43084;
  assign n43086 = n43013 & ~n43085;
  assign n43087 = pi299 & ~n43086;
  assign n43088 = ~pi224 & n41340;
  assign n43089 = pi224 & ~pi276;
  assign n43090 = ~pi222 & ~n43089;
  assign n43091 = ~n43088 & n43090;
  assign n43092 = n42979 & ~n43091;
  assign n43093 = n42983 & ~n43092;
  assign n43094 = ~pi39 & ~n43093;
  assign n43095 = ~n42982 & ~n43092;
  assign n43096 = ~pi299 & ~n43095;
  assign n43097 = pi299 & n43013;
  assign n43098 = ~n43085 & n43097;
  assign n43099 = ~n43096 & ~n43098;
  assign n43100 = ~pi39 & ~n43099;
  assign n43101 = ~n43087 & n43094;
  assign n43102 = ~n41418 & n43013;
  assign n43103 = ~pi215 & ~n43102;
  assign n43104 = pi154 & ~n43102;
  assign n43105 = ~n43020 & ~n43104;
  assign n43106 = ~n43020 & ~n43103;
  assign n43107 = ~n43104 & n43106;
  assign n43108 = ~n43103 & n43105;
  assign n43109 = pi299 & ~n60772;
  assign n43110 = ~n60722 & ~n42984;
  assign n43111 = ~n43109 & n43110;
  assign n43112 = ~n60769 & ~n60772;
  assign n43113 = pi299 & ~n43112;
  assign n43114 = ~n43111 & ~n43113;
  assign n43115 = pi39 & ~n43114;
  assign n43116 = n2636 & ~n43115;
  assign n43117 = ~n60771 & n43116;
  assign n43118 = pi100 & n43043;
  assign n43119 = ~n2636 & ~n43111;
  assign n43120 = ~n43118 & n43119;
  assign n43121 = ~n43117 & ~n43120;
  assign n43122 = ~pi87 & ~n43121;
  assign n43123 = n58815 & n43113;
  assign n43124 = pi87 & ~n43111;
  assign n43125 = ~n43123 & n43124;
  assign n43126 = ~pi75 & ~n43125;
  assign n43127 = ~n43122 & n43126;
  assign n43128 = pi75 & n43111;
  assign n43129 = ~pi92 & ~n43128;
  assign n43130 = ~n43127 & n43129;
  assign n43131 = n6309 & n43123;
  assign n43132 = n60069 & n43113;
  assign n43133 = pi92 & ~n43111;
  assign n43134 = ~n60773 & n43133;
  assign n43135 = n6306 & ~n43134;
  assign n43136 = ~n43130 & n43135;
  assign n43137 = ~n6306 & n43111;
  assign n43138 = ~pi55 & ~n43137;
  assign n43139 = ~n43136 & n43138;
  assign n43140 = pi55 & ~n60772;
  assign n43141 = ~n43062 & n43140;
  assign n43142 = ~pi56 & ~n43141;
  assign n43143 = ~n43139 & n43142;
  assign n43144 = n60070 & n43112;
  assign n43145 = ~n60070 & ~n60772;
  assign n43146 = pi56 & ~n43145;
  assign n43147 = ~n43144 & n43146;
  assign n43148 = ~pi62 & ~n43147;
  assign n43149 = ~n43143 & n43148;
  assign n43150 = n41492 & n60769;
  assign n43151 = pi62 & ~n60772;
  assign n43152 = ~n41492 & ~n60772;
  assign n43153 = ~pi56 & n43144;
  assign n43154 = ~n43152 & ~n43153;
  assign n43155 = pi62 & ~n43154;
  assign n43156 = ~n43150 & n43151;
  assign n43157 = n4438 & ~n60774;
  assign n43158 = ~n43149 & n43157;
  assign n43159 = ~n4438 & n60772;
  assign n43160 = pi239 & ~n43159;
  assign n43161 = ~n43158 & n43160;
  assign n43162 = ~n43081 & ~n43161;
  assign n43163 = ~pi927 & n38221;
  assign n43164 = ~pi1145 & ~n38221;
  assign n43165 = pi221 & ~n43164;
  assign n43166 = pi221 & ~n43163;
  assign n43167 = ~n43164 & n43166;
  assign n43168 = ~n43163 & n43165;
  assign n43169 = pi216 & pi274;
  assign n43170 = ~pi221 & ~n43169;
  assign n43171 = ~pi151 & n42183;
  assign n43172 = pi151 & n42174;
  assign n43173 = ~pi216 & ~n43172;
  assign n43174 = ~n43171 & n43173;
  assign n43175 = n43170 & ~n43174;
  assign n43176 = ~n60775 & ~n43175;
  assign n43177 = ~pi215 & ~n43176;
  assign n43178 = pi215 & pi1145;
  assign n43179 = pi299 & ~n43178;
  assign n43180 = ~n43177 & n43179;
  assign n43181 = ~pi927 & n38636;
  assign n43182 = ~pi1145 & ~n38636;
  assign n43183 = pi222 & ~n43182;
  assign n43184 = pi222 & ~n43181;
  assign n43185 = ~n43182 & n43184;
  assign n43186 = ~n43181 & n43183;
  assign n43187 = pi224 & pi274;
  assign n43188 = ~pi222 & ~n43187;
  assign n43189 = ~n43088 & n43188;
  assign n43190 = ~n60776 & ~n43189;
  assign n43191 = ~pi223 & ~n43190;
  assign n43192 = pi223 & pi1145;
  assign n43193 = ~pi299 & ~n43192;
  assign n43194 = ~n43191 & n43193;
  assign n43195 = ~pi39 & ~n43194;
  assign n43196 = ~n43180 & n43195;
  assign n43197 = n26651 & ~n43187;
  assign n43198 = ~n60776 & ~n43197;
  assign n43199 = ~pi223 & ~n43198;
  assign n43200 = ~n43192 & ~n43199;
  assign n43201 = ~pi299 & ~n43200;
  assign n43202 = ~n60722 & ~n43201;
  assign n43203 = ~pi151 & ~n38211;
  assign n43204 = ~n41403 & ~n43203;
  assign n43205 = ~pi151 & n31586;
  assign n43206 = ~n43204 & ~n43205;
  assign n43207 = ~pi216 & ~n43206;
  assign n43208 = n43170 & ~n43207;
  assign n43209 = ~n60775 & ~n43208;
  assign n43210 = ~pi215 & ~n43209;
  assign n43211 = ~n43178 & ~n43210;
  assign n43212 = pi299 & ~n43211;
  assign n43213 = n43202 & ~n43212;
  assign n43214 = pi39 & ~n43213;
  assign n43215 = ~pi38 & ~n43214;
  assign n43216 = ~n43196 & n43215;
  assign n43217 = ~pi216 & ~n43203;
  assign n43218 = n43170 & ~n43217;
  assign n43219 = ~n60775 & ~n43218;
  assign n43220 = ~pi215 & ~n43219;
  assign n43221 = ~n43178 & ~n43220;
  assign n43222 = n41673 & ~n43169;
  assign n43223 = n43221 & ~n43222;
  assign n43224 = pi299 & ~n43223;
  assign n43225 = n43202 & ~n43224;
  assign n43226 = pi38 & n43225;
  assign n43227 = ~pi100 & ~n43226;
  assign n43228 = ~n43216 & n43227;
  assign n43229 = ~pi151 & n42110;
  assign n43230 = n43207 & ~n43229;
  assign n43231 = n43170 & ~n43230;
  assign n43232 = ~n60775 & ~n43231;
  assign n43233 = ~pi215 & ~n43232;
  assign n43234 = ~n43178 & ~n43233;
  assign n43235 = pi299 & ~n43234;
  assign n43236 = n2634 & n43202;
  assign n43237 = ~n43235 & n43236;
  assign n43238 = ~n2634 & n43225;
  assign n43239 = pi100 & ~n43238;
  assign n43240 = ~n43237 & n43239;
  assign n43241 = ~n43228 & ~n43240;
  assign n43242 = ~pi87 & ~n43241;
  assign n43243 = ~n58815 & n43225;
  assign n43244 = n58815 & n43213;
  assign n43245 = ~n43243 & ~n43244;
  assign n43246 = pi87 & n43245;
  assign n43247 = ~pi75 & ~n43246;
  assign n43248 = ~n43242 & n43247;
  assign n43249 = pi75 & n43225;
  assign n43250 = ~pi92 & ~n43249;
  assign n43251 = ~n43248 & n43250;
  assign n43252 = n6309 & ~n43245;
  assign n43253 = ~n6309 & n43225;
  assign n43254 = pi92 & ~n43253;
  assign n43255 = ~n43252 & n43254;
  assign n43256 = n6306 & ~n43255;
  assign n43257 = ~n43251 & n43256;
  assign n43258 = ~n6306 & n43225;
  assign n43259 = ~pi55 & ~n43258;
  assign n43260 = ~n43257 & n43259;
  assign n43261 = n28288 & n43211;
  assign n43262 = ~n28288 & n43223;
  assign n43263 = pi55 & ~n43262;
  assign n43264 = ~n43261 & n43263;
  assign n43265 = ~pi56 & ~n43264;
  assign n43266 = ~n43260 & n43265;
  assign n43267 = n60070 & ~n43211;
  assign n43268 = ~n60070 & ~n43223;
  assign n43269 = pi56 & ~n43268;
  assign n43270 = ~n60070 & n43223;
  assign n43271 = ~pi55 & n43261;
  assign n43272 = ~n43270 & ~n43271;
  assign n43273 = pi56 & ~n43272;
  assign n43274 = ~n43267 & n43269;
  assign n43275 = ~pi62 & ~n60777;
  assign n43276 = ~n43266 & n43275;
  assign n43277 = n41492 & n43211;
  assign n43278 = ~n41492 & n43223;
  assign n43279 = pi62 & ~n43278;
  assign n43280 = ~n43277 & n43279;
  assign n43281 = pi235 & n4438;
  assign n43282 = ~n43280 & n43281;
  assign n43283 = ~n43276 & n43282;
  assign n43284 = n42992 & ~n43178;
  assign n43285 = ~n60775 & n43284;
  assign n43286 = ~n60775 & ~n43178;
  assign n43287 = n42997 & n43286;
  assign n43288 = n58822 & n43285;
  assign n43289 = pi299 & ~n43221;
  assign n43290 = ~n60778 & n43289;
  assign n43291 = n58815 & ~n43201;
  assign n43292 = ~n43290 & n43291;
  assign n43293 = ~n43201 & ~n43289;
  assign n43294 = ~n58815 & n43293;
  assign n43295 = ~n43292 & ~n43294;
  assign n43296 = pi87 & ~n43295;
  assign n43297 = ~pi100 & n40750;
  assign n43298 = ~pi39 & pi100;
  assign n43299 = n41439 & n43298;
  assign n43300 = ~n43297 & ~n43299;
  assign n43301 = n43038 & n43286;
  assign n43302 = ~pi38 & n43285;
  assign n43303 = ~n43300 & n60779;
  assign n43304 = n43289 & ~n43303;
  assign n43305 = ~pi87 & ~n43201;
  assign n43306 = ~n43304 & n43305;
  assign n43307 = ~n43296 & ~n43306;
  assign n43308 = ~pi75 & ~n43307;
  assign n43309 = pi75 & n43293;
  assign n43310 = ~pi92 & ~n43309;
  assign n43311 = ~n43308 & n43310;
  assign n43312 = n6309 & n43292;
  assign n43313 = ~n60069 & n43293;
  assign n43314 = pi92 & ~n43313;
  assign n43315 = ~n43312 & n43314;
  assign n43316 = n6306 & ~n43315;
  assign n43317 = ~n43311 & n43316;
  assign n43318 = ~n6306 & n43293;
  assign n43319 = ~pi55 & ~n43318;
  assign n43320 = ~n43317 & n43319;
  assign n43321 = n28288 & n60778;
  assign n43322 = pi55 & ~n43221;
  assign n43323 = ~n43321 & n43322;
  assign n43324 = ~pi56 & ~n43323;
  assign n43325 = ~n43320 & n43324;
  assign n43326 = ~pi55 & n43321;
  assign n43327 = n60070 & n60778;
  assign n43328 = ~n43221 & ~n60780;
  assign n43329 = pi56 & ~n43328;
  assign n43330 = ~pi62 & ~n43329;
  assign n43331 = ~n43325 & n43330;
  assign n43332 = ~pi56 & n60780;
  assign n43333 = n41492 & n60778;
  assign n43334 = pi62 & ~n43221;
  assign n43335 = ~n60781 & n43334;
  assign n43336 = ~pi235 & n4438;
  assign n43337 = ~n43335 & n43336;
  assign n43338 = ~n43331 & n43337;
  assign n43339 = pi235 & n43222;
  assign n43340 = ~n4438 & ~n43339;
  assign n43341 = n43221 & n43340;
  assign n43342 = ~n43338 & ~n43341;
  assign po155 = ~n43283 & n43342;
  assign n43344 = pi223 & pi1143;
  assign n43345 = ~pi299 & ~n43344;
  assign n43346 = ~pi944 & n38636;
  assign n43347 = ~pi1143 & ~n38636;
  assign n43348 = pi222 & ~n43347;
  assign n43349 = pi222 & ~n43346;
  assign n43350 = ~n43347 & n43349;
  assign n43351 = ~n43346 & n43348;
  assign n43352 = pi224 & pi264;
  assign n43353 = ~pi222 & ~n43352;
  assign n43354 = ~pi284 & n41340;
  assign n43355 = ~pi224 & ~n43354;
  assign n43356 = n43353 & ~n43355;
  assign n43357 = ~n60782 & ~n43356;
  assign n43358 = ~n41340 & n43353;
  assign n43359 = n43357 & ~n43358;
  assign n43360 = ~pi223 & ~n43359;
  assign n43361 = n43345 & ~n43360;
  assign n43362 = ~pi39 & ~n43361;
  assign n43363 = pi215 & pi1143;
  assign n43364 = pi299 & ~n43363;
  assign n43365 = ~pi944 & n38221;
  assign n43366 = ~pi1143 & ~n38221;
  assign n43367 = pi221 & ~n43366;
  assign n43368 = pi221 & ~n43365;
  assign n43369 = ~n43366 & n43368;
  assign n43370 = ~n43365 & n43367;
  assign n43371 = pi216 & pi264;
  assign n43372 = ~pi221 & ~n43371;
  assign n43373 = pi284 & ~n28313;
  assign n43374 = pi105 & ~n43373;
  assign n43375 = ~pi105 & pi146;
  assign n43376 = pi228 & ~n43375;
  assign n43377 = ~n43374 & n43376;
  assign n43378 = ~n41356 & n43377;
  assign n43379 = pi146 & ~n41335;
  assign n43380 = ~pi146 & n41346;
  assign n43381 = pi284 & ~n43380;
  assign n43382 = ~n43379 & n43381;
  assign n43383 = ~pi146 & ~pi284;
  assign n43384 = ~n40748 & n43383;
  assign n43385 = ~n43382 & ~n43384;
  assign n43386 = ~pi228 & ~n43385;
  assign n43387 = ~n43378 & ~n43386;
  assign n43388 = ~pi216 & ~n43387;
  assign n43389 = n43372 & ~n43388;
  assign n43390 = ~n60783 & ~n43389;
  assign n43391 = ~pi215 & ~n43390;
  assign n43392 = n43364 & ~n43391;
  assign n43393 = n43362 & ~n43392;
  assign n43394 = ~pi224 & n43373;
  assign n43395 = n43353 & ~n43394;
  assign n43396 = ~n60782 & ~n43395;
  assign n43397 = ~pi223 & ~n43396;
  assign n43398 = ~n43344 & ~n43397;
  assign n43399 = ~pi299 & ~n43398;
  assign n43400 = ~pi284 & n58822;
  assign n43401 = pi146 & ~n58822;
  assign n43402 = ~pi228 & ~n43401;
  assign n43403 = pi284 & n58822;
  assign n43404 = ~n41431 & ~n43403;
  assign n43405 = ~pi228 & ~n43404;
  assign n43406 = ~n43400 & n43402;
  assign n43407 = ~n43377 & ~n60784;
  assign n43408 = ~pi216 & ~n43407;
  assign n43409 = n43372 & ~n43408;
  assign n43410 = ~n60783 & ~n43409;
  assign n43411 = ~pi215 & ~n43410;
  assign n43412 = ~n43363 & ~n43411;
  assign n43413 = pi299 & ~n43412;
  assign n43414 = ~n43399 & ~n43413;
  assign n43415 = pi39 & ~n43414;
  assign n43416 = ~pi38 & ~n43415;
  assign n43417 = ~n43393 & n43416;
  assign n43418 = ~n41403 & ~n43377;
  assign n43419 = ~pi146 & ~pi228;
  assign n43420 = n43418 & ~n43419;
  assign n43421 = ~pi216 & ~n43420;
  assign n43422 = n43372 & ~n43421;
  assign n43423 = ~n60783 & ~n43422;
  assign n43424 = ~pi215 & ~n43423;
  assign n43425 = ~n43363 & ~n43424;
  assign n43426 = n41673 & ~n43371;
  assign n43427 = n43425 & ~n43426;
  assign n43428 = pi299 & ~n43427;
  assign n43429 = ~n43399 & ~n43428;
  assign n43430 = pi38 & n43429;
  assign n43431 = ~pi100 & ~n43430;
  assign n43432 = ~n43417 & n43431;
  assign n43433 = pi252 & n2677;
  assign n43434 = ~pi284 & ~n43433;
  assign n43435 = n43400 & ~n43433;
  assign n43436 = n58822 & n43434;
  assign n43437 = ~pi228 & ~n60785;
  assign n43438 = ~pi228 & ~n41432;
  assign n43439 = ~n60785 & n43438;
  assign n43440 = ~n41432 & n43437;
  assign n43441 = ~n43377 & ~n60786;
  assign n43442 = ~pi216 & ~n43441;
  assign n43443 = n43372 & ~n43442;
  assign n43444 = ~n60783 & ~n43443;
  assign n43445 = ~pi215 & ~n43444;
  assign n43446 = ~n43363 & ~n43445;
  assign n43447 = pi299 & ~n43446;
  assign n43448 = n2634 & ~n43399;
  assign n43449 = ~n43447 & n43448;
  assign n43450 = ~n2634 & n43429;
  assign n43451 = pi100 & ~n43450;
  assign n43452 = ~n43449 & n43451;
  assign n43453 = ~n43432 & ~n43452;
  assign n43454 = ~pi87 & ~n43453;
  assign n43455 = ~n58815 & n43429;
  assign n43456 = n58815 & n43414;
  assign n43457 = ~n43455 & ~n43456;
  assign n43458 = pi87 & n43457;
  assign n43459 = ~pi75 & ~n43458;
  assign n43460 = ~n43454 & n43459;
  assign n43461 = pi75 & n43429;
  assign n43462 = ~pi92 & ~n43461;
  assign n43463 = ~n43460 & n43462;
  assign n43464 = n6309 & ~n43457;
  assign n43465 = ~n6309 & n43429;
  assign n43466 = pi92 & ~n43465;
  assign n43467 = ~n43464 & n43466;
  assign n43468 = n6306 & ~n43467;
  assign n43469 = ~n43463 & n43468;
  assign n43470 = ~n6306 & n43429;
  assign n43471 = ~pi55 & ~n43470;
  assign n43472 = ~n43469 & n43471;
  assign n43473 = n28288 & n43412;
  assign n43474 = ~n28288 & n43427;
  assign n43475 = pi55 & ~n43474;
  assign n43476 = ~n43473 & n43475;
  assign n43477 = ~pi56 & ~n43476;
  assign n43478 = ~n43472 & n43477;
  assign n43479 = n60070 & ~n43412;
  assign n43480 = ~n60070 & ~n43427;
  assign n43481 = pi56 & ~n43480;
  assign n43482 = ~pi55 & n43473;
  assign n43483 = ~n60070 & n43427;
  assign n43484 = ~n43482 & ~n43483;
  assign n43485 = pi56 & ~n43484;
  assign n43486 = ~n43479 & n43481;
  assign n43487 = ~pi62 & ~n60787;
  assign n43488 = ~n43478 & n43487;
  assign n43489 = n41492 & n43412;
  assign n43490 = ~n41492 & n43427;
  assign n43491 = pi62 & ~n43490;
  assign n43492 = ~n43489 & n43491;
  assign n43493 = pi238 & n4438;
  assign n43494 = ~n43492 & n43493;
  assign n43495 = ~n43488 & n43494;
  assign n43496 = ~pi146 & ~n41335;
  assign n43497 = pi146 & n41346;
  assign n43498 = ~pi284 & ~n43497;
  assign n43499 = ~n43496 & n43498;
  assign n43500 = pi146 & pi284;
  assign n43501 = ~n40748 & n43500;
  assign n43502 = ~pi228 & ~n43501;
  assign n43503 = pi146 & ~n40748;
  assign n43504 = pi284 & ~n43503;
  assign n43505 = ~pi146 & n41335;
  assign n43506 = pi146 & ~n41346;
  assign n43507 = ~pi284 & ~n43506;
  assign n43508 = ~n43505 & n43507;
  assign n43509 = ~n43498 & ~n43501;
  assign n43510 = ~n43496 & ~n43509;
  assign n43511 = ~n43504 & ~n43508;
  assign n43512 = ~pi228 & ~n60788;
  assign n43513 = ~n43499 & n43502;
  assign n43514 = ~n41628 & ~n43377;
  assign n43515 = ~n60789 & n43514;
  assign n43516 = ~pi216 & ~n43515;
  assign n43517 = n43372 & ~n43516;
  assign n43518 = ~n60783 & ~n43517;
  assign n43519 = ~pi215 & ~n43518;
  assign n43520 = n43364 & ~n43519;
  assign n43521 = n43345 & n43357;
  assign n43522 = n43362 & ~n43521;
  assign n43523 = ~n43520 & n43522;
  assign n43524 = ~n41391 & n43399;
  assign n43525 = ~n60784 & n43418;
  assign n43526 = ~pi216 & ~n43525;
  assign n43527 = n43372 & ~n43526;
  assign n43528 = ~n60783 & ~n43527;
  assign n43529 = ~pi215 & ~n43528;
  assign n43530 = ~n43363 & ~n43529;
  assign n43531 = pi299 & ~n43530;
  assign n43532 = ~n43524 & ~n43531;
  assign n43533 = pi39 & ~n43532;
  assign n43534 = ~pi38 & ~n43533;
  assign n43535 = ~n43523 & n43534;
  assign n43536 = pi299 & ~n43425;
  assign n43537 = ~n43524 & ~n43536;
  assign n43538 = pi38 & n43537;
  assign n43539 = ~pi100 & ~n43538;
  assign n43540 = ~n43535 & n43539;
  assign n43541 = n43418 & ~n60786;
  assign n43542 = ~pi216 & ~n43541;
  assign n43543 = n43372 & ~n43542;
  assign n43544 = ~n60783 & ~n43543;
  assign n43545 = ~pi215 & ~n43544;
  assign n43546 = ~n43363 & ~n43545;
  assign n43547 = pi299 & ~n43546;
  assign n43548 = n2634 & ~n43524;
  assign n43549 = ~n43547 & n43548;
  assign n43550 = ~n2634 & n43537;
  assign n43551 = pi100 & ~n43550;
  assign n43552 = ~n43549 & n43551;
  assign n43553 = ~n43540 & ~n43552;
  assign n43554 = ~pi87 & ~n43553;
  assign n43555 = ~n58815 & n43537;
  assign n43556 = n58815 & n43532;
  assign n43557 = ~n43555 & ~n43556;
  assign n43558 = pi87 & n43557;
  assign n43559 = ~pi75 & ~n43558;
  assign n43560 = ~n43554 & n43559;
  assign n43561 = pi75 & n43537;
  assign n43562 = ~pi92 & ~n43561;
  assign n43563 = ~n43560 & n43562;
  assign n43564 = n6309 & ~n43557;
  assign n43565 = ~n6309 & n43537;
  assign n43566 = pi92 & ~n43565;
  assign n43567 = ~n43564 & n43566;
  assign n43568 = n6306 & ~n43567;
  assign n43569 = ~n43563 & n43568;
  assign n43570 = ~n6306 & n43537;
  assign n43571 = ~pi55 & ~n43570;
  assign n43572 = ~n43569 & n43571;
  assign n43573 = n28288 & n43530;
  assign n43574 = ~n28288 & n43425;
  assign n43575 = pi55 & ~n43574;
  assign n43576 = ~n43573 & n43575;
  assign n43577 = ~pi56 & ~n43576;
  assign n43578 = ~n43572 & n43577;
  assign n43579 = n60070 & ~n43530;
  assign n43580 = ~n60070 & ~n43425;
  assign n43581 = pi56 & ~n43580;
  assign n43582 = ~n60070 & n43425;
  assign n43583 = ~pi55 & n43573;
  assign n43584 = ~n43582 & ~n43583;
  assign n43585 = pi56 & ~n43584;
  assign n43586 = ~n43579 & n43581;
  assign n43587 = ~pi62 & ~n60790;
  assign n43588 = ~n43578 & n43587;
  assign n43589 = n41492 & n43530;
  assign n43590 = ~n41492 & n43425;
  assign n43591 = pi62 & ~n43590;
  assign n43592 = ~n43589 & n43591;
  assign n43593 = ~pi238 & n4438;
  assign n43594 = ~n43592 & n43593;
  assign n43595 = ~n43588 & n43594;
  assign n43596 = pi238 & n43426;
  assign n43597 = ~n4438 & ~n43596;
  assign n43598 = n43425 & n43597;
  assign n43599 = ~n43595 & ~n43598;
  assign po156 = ~n43495 & n43599;
  assign n43601 = ~pi928 & n38221;
  assign n43602 = ~pi1136 & ~n38221;
  assign n43603 = pi221 & ~n43602;
  assign n43604 = pi221 & ~n43601;
  assign n43605 = ~n43602 & n43604;
  assign n43606 = ~n43601 & n43603;
  assign n43607 = pi216 & pi266;
  assign n43608 = ~pi166 & ~n41335;
  assign n43609 = pi166 & n41346;
  assign n43610 = pi875 & ~n43609;
  assign n43611 = ~n43608 & n43610;
  assign n43612 = pi166 & ~pi875;
  assign n43613 = ~n40748 & n43612;
  assign n43614 = ~pi228 & ~n43613;
  assign n43615 = ~n43611 & n43614;
  assign n43616 = pi875 & ~n28313;
  assign n43617 = pi105 & ~n43616;
  assign n43618 = ~pi105 & ~pi166;
  assign n43619 = ~n43617 & ~n43618;
  assign n43620 = n42172 & ~n43619;
  assign n43621 = ~pi216 & ~n43620;
  assign n43622 = ~n41628 & n43621;
  assign n43623 = ~n43611 & ~n43613;
  assign n43624 = ~pi228 & ~n43623;
  assign n43625 = ~n42172 & ~n43624;
  assign n43626 = n43621 & ~n43625;
  assign n43627 = ~n43615 & n43622;
  assign n43628 = ~n43607 & ~n60792;
  assign n43629 = ~pi221 & ~n43628;
  assign n43630 = ~n60791 & ~n43629;
  assign n43631 = ~pi215 & ~n43630;
  assign n43632 = pi215 & pi1136;
  assign n43633 = pi299 & ~n43632;
  assign n43634 = ~n43631 & n43633;
  assign n43635 = ~pi224 & ~pi875;
  assign n43636 = ~n28313 & n43635;
  assign n43637 = pi224 & ~pi266;
  assign n43638 = ~pi222 & ~n43637;
  assign n43639 = ~n43636 & n43638;
  assign n43640 = n6544 & ~n41340;
  assign n43641 = n43639 & ~n43640;
  assign n43642 = ~pi928 & n38636;
  assign n43643 = ~pi1136 & ~n38636;
  assign n43644 = pi222 & ~n43643;
  assign n43645 = pi222 & ~n43642;
  assign n43646 = ~n43643 & n43645;
  assign n43647 = ~n43642 & n43644;
  assign n43648 = pi223 & pi1136;
  assign n43649 = ~pi299 & ~n43648;
  assign n43650 = ~n60793 & n43649;
  assign n43651 = ~n43641 & n43650;
  assign n43652 = ~n43639 & ~n60793;
  assign n43653 = ~n43640 & n43652;
  assign n43654 = ~pi223 & ~n43653;
  assign n43655 = n43649 & ~n43654;
  assign n43656 = ~pi39 & ~n43655;
  assign n43657 = ~n43651 & n43656;
  assign n43658 = ~n43634 & n43657;
  assign n43659 = ~pi223 & ~n43652;
  assign n43660 = ~n43648 & ~n43659;
  assign n43661 = ~pi299 & ~n43660;
  assign n43662 = n35583 & ~n43616;
  assign n43663 = n43661 & ~n43662;
  assign n43664 = pi228 & n43619;
  assign n43665 = ~pi875 & n58822;
  assign n43666 = ~pi166 & ~n58822;
  assign n43667 = ~pi228 & ~n43666;
  assign n43668 = ~pi228 & ~n43665;
  assign n43669 = ~n43666 & n43668;
  assign n43670 = ~n43665 & n43667;
  assign n43671 = ~n43664 & ~n60794;
  assign n43672 = ~pi216 & ~n43671;
  assign n43673 = ~n43607 & ~n43672;
  assign n43674 = ~pi221 & ~n43673;
  assign n43675 = ~n60791 & ~n43674;
  assign n43676 = ~pi215 & ~n43675;
  assign n43677 = ~n43632 & ~n43676;
  assign n43678 = pi299 & ~n43677;
  assign n43679 = ~n43663 & ~n43678;
  assign n43680 = pi39 & ~n43679;
  assign n43681 = ~pi38 & ~n43680;
  assign n43682 = ~n43658 & n43681;
  assign n43683 = pi166 & ~pi228;
  assign n43684 = ~n43664 & ~n43683;
  assign n43685 = ~pi216 & ~n43684;
  assign n43686 = ~n43607 & ~n43685;
  assign n43687 = ~pi221 & ~n43686;
  assign n43688 = ~n60791 & ~n43687;
  assign n43689 = ~pi215 & ~n43688;
  assign n43690 = ~n43632 & ~n43689;
  assign n43691 = pi299 & ~n43690;
  assign n43692 = ~n43663 & ~n43691;
  assign n43693 = pi38 & n43692;
  assign n43694 = ~pi100 & ~n43693;
  assign n43695 = ~n43682 & n43694;
  assign n43696 = ~pi875 & n41433;
  assign n43697 = pi166 & ~n43696;
  assign n43698 = ~n2676 & ~n41433;
  assign n43699 = n2676 & ~n28550;
  assign n43700 = pi875 & ~n43699;
  assign n43701 = ~n43698 & n43700;
  assign n43702 = ~n43697 & ~n43701;
  assign n43703 = ~pi228 & ~n43702;
  assign n43704 = ~n43664 & ~n43703;
  assign n43705 = ~pi216 & ~n43704;
  assign n43706 = ~n43607 & ~n43705;
  assign n43707 = ~pi221 & ~n43706;
  assign n43708 = ~n60791 & ~n43707;
  assign n43709 = ~pi215 & ~n43708;
  assign n43710 = ~n43632 & ~n43709;
  assign n43711 = pi299 & ~n43710;
  assign n43712 = n2634 & ~n43663;
  assign n43713 = ~n43711 & n43712;
  assign n43714 = ~n2634 & n43692;
  assign n43715 = pi100 & ~n43714;
  assign n43716 = ~n43713 & n43715;
  assign n43717 = ~n43695 & ~n43716;
  assign n43718 = ~pi87 & ~n43717;
  assign n43719 = ~n58815 & n43692;
  assign n43720 = n58815 & n43679;
  assign n43721 = ~n43719 & ~n43720;
  assign n43722 = pi87 & n43721;
  assign n43723 = ~pi75 & ~n43722;
  assign n43724 = ~n43718 & n43723;
  assign n43725 = pi75 & n43692;
  assign n43726 = ~pi92 & ~n43725;
  assign n43727 = ~n43724 & n43726;
  assign n43728 = n6309 & ~n43721;
  assign n43729 = ~n6309 & n43692;
  assign n43730 = pi92 & ~n43729;
  assign n43731 = ~n43728 & n43730;
  assign n43732 = n6306 & ~n43731;
  assign n43733 = ~n43727 & n43732;
  assign n43734 = ~n6306 & n43692;
  assign n43735 = ~pi55 & ~n43734;
  assign n43736 = ~n43733 & n43735;
  assign n43737 = n28288 & n43677;
  assign n43738 = ~n28288 & n43690;
  assign n43739 = pi55 & ~n43738;
  assign n43740 = ~n43737 & n43739;
  assign n43741 = ~pi56 & ~n43740;
  assign n43742 = ~n43736 & n43741;
  assign n43743 = n60070 & ~n43677;
  assign n43744 = ~n60070 & ~n43690;
  assign n43745 = pi56 & ~n43744;
  assign n43746 = ~n60070 & n43690;
  assign n43747 = ~pi55 & n43737;
  assign n43748 = ~n43746 & ~n43747;
  assign n43749 = pi56 & ~n43748;
  assign n43750 = ~n43743 & n43745;
  assign n43751 = ~pi62 & ~n60795;
  assign n43752 = ~n43742 & n43751;
  assign n43753 = n41492 & n43677;
  assign n43754 = ~n41492 & n43690;
  assign n43755 = pi62 & ~n43754;
  assign n43756 = ~n43753 & n43755;
  assign n43757 = n4438 & ~n43756;
  assign n43758 = ~n43752 & n43757;
  assign n43759 = ~n4438 & n43690;
  assign n43760 = ~pi245 & ~n43759;
  assign n43761 = ~n43758 & n43760;
  assign n43762 = ~pi166 & ~n40748;
  assign n43763 = pi875 & ~n43762;
  assign n43764 = pi166 & n41335;
  assign n43765 = ~pi166 & ~n41346;
  assign n43766 = ~pi875 & ~n43765;
  assign n43767 = ~n43764 & n43766;
  assign n43768 = ~pi228 & ~n43767;
  assign n43769 = ~pi228 & ~n43763;
  assign n43770 = ~n43767 & n43769;
  assign n43771 = ~n43763 & n43768;
  assign n43772 = n43621 & ~n60796;
  assign n43773 = ~n43607 & ~n43772;
  assign n43774 = ~pi221 & ~n43773;
  assign n43775 = ~n60791 & ~n43774;
  assign n43776 = ~pi215 & ~n43775;
  assign n43777 = n43633 & ~n43776;
  assign n43778 = n43656 & ~n43777;
  assign n43779 = ~n41403 & ~n43664;
  assign n43780 = ~n60794 & n43779;
  assign n43781 = ~pi216 & ~n43780;
  assign n43782 = ~n43607 & ~n43781;
  assign n43783 = ~pi221 & ~n43782;
  assign n43784 = ~n60791 & ~n43783;
  assign n43785 = ~pi215 & ~n43784;
  assign n43786 = ~n43632 & ~n43785;
  assign n43787 = pi299 & ~n43786;
  assign n43788 = ~n43661 & ~n43787;
  assign n43789 = pi39 & ~n43788;
  assign n43790 = ~pi38 & ~n43789;
  assign n43791 = ~n43778 & n43790;
  assign n43792 = ~n41418 & n43690;
  assign n43793 = pi299 & ~n43792;
  assign n43794 = ~n43661 & ~n43793;
  assign n43795 = pi38 & n43794;
  assign n43796 = ~pi100 & ~n43795;
  assign n43797 = ~n43791 & n43796;
  assign n43798 = ~n43703 & n43779;
  assign n43799 = ~pi216 & ~n43798;
  assign n43800 = ~n43607 & ~n43799;
  assign n43801 = ~pi221 & ~n43800;
  assign n43802 = ~n60791 & ~n43801;
  assign n43803 = ~pi215 & ~n43802;
  assign n43804 = ~n43632 & ~n43803;
  assign n43805 = pi299 & ~n43804;
  assign n43806 = n2634 & ~n43661;
  assign n43807 = ~n43805 & n43806;
  assign n43808 = ~n2634 & n43794;
  assign n43809 = pi100 & ~n43808;
  assign n43810 = ~n43807 & n43809;
  assign n43811 = ~n43797 & ~n43810;
  assign n43812 = ~pi87 & ~n43811;
  assign n43813 = ~n58815 & n43794;
  assign n43814 = n58815 & n43788;
  assign n43815 = ~n43813 & ~n43814;
  assign n43816 = pi87 & n43815;
  assign n43817 = ~pi75 & ~n43816;
  assign n43818 = ~n43812 & n43817;
  assign n43819 = pi75 & n43794;
  assign n43820 = ~pi92 & ~n43819;
  assign n43821 = ~n43818 & n43820;
  assign n43822 = n6309 & ~n43815;
  assign n43823 = ~n6309 & n43794;
  assign n43824 = pi92 & ~n43823;
  assign n43825 = ~n43822 & n43824;
  assign n43826 = n6306 & ~n43825;
  assign n43827 = ~n43821 & n43826;
  assign n43828 = ~n6306 & n43794;
  assign n43829 = ~pi55 & ~n43828;
  assign n43830 = ~n43827 & n43829;
  assign n43831 = n28288 & n43786;
  assign n43832 = ~n28288 & n43792;
  assign n43833 = pi55 & ~n43832;
  assign n43834 = ~n43831 & n43833;
  assign n43835 = ~pi56 & ~n43834;
  assign n43836 = ~n43830 & n43835;
  assign n43837 = n60070 & ~n43786;
  assign n43838 = ~n60070 & ~n43792;
  assign n43839 = pi56 & ~n43838;
  assign n43840 = ~pi55 & n43831;
  assign n43841 = ~n60070 & n43792;
  assign n43842 = ~n43840 & ~n43841;
  assign n43843 = pi56 & ~n43842;
  assign n43844 = ~n43837 & n43839;
  assign n43845 = ~pi62 & ~n60797;
  assign n43846 = ~n43836 & n43845;
  assign n43847 = n41492 & n43786;
  assign n43848 = ~n41492 & n43792;
  assign n43849 = pi62 & ~n43848;
  assign n43850 = ~n43847 & n43849;
  assign n43851 = n4438 & ~n43850;
  assign n43852 = ~n43846 & n43851;
  assign n43853 = ~n4438 & n43792;
  assign n43854 = pi245 & ~n43853;
  assign n43855 = ~n43852 & n43854;
  assign n43856 = ~n43761 & ~n43855;
  assign n43857 = ~pi938 & n38221;
  assign n43858 = ~pi1135 & ~n38221;
  assign n43859 = pi221 & ~n43858;
  assign n43860 = pi221 & ~n43857;
  assign n43861 = ~n43858 & n43860;
  assign n43862 = ~n43857 & n43859;
  assign n43863 = pi216 & pi279;
  assign n43864 = ~pi161 & ~n41335;
  assign n43865 = pi161 & n41346;
  assign n43866 = pi879 & ~n43865;
  assign n43867 = ~n43864 & n43866;
  assign n43868 = pi161 & ~pi879;
  assign n43869 = ~n40748 & n43868;
  assign n43870 = ~pi228 & ~n43869;
  assign n43871 = ~n43867 & n43870;
  assign n43872 = pi879 & ~n28313;
  assign n43873 = pi105 & ~n43872;
  assign n43874 = ~pi105 & ~pi161;
  assign n43875 = ~n43873 & ~n43874;
  assign n43876 = n42172 & ~n43875;
  assign n43877 = ~pi216 & ~n43876;
  assign n43878 = ~n41628 & n43877;
  assign n43879 = ~n43867 & ~n43869;
  assign n43880 = ~pi228 & ~n43879;
  assign n43881 = ~n42172 & ~n43880;
  assign n43882 = n43877 & ~n43881;
  assign n43883 = ~n43871 & n43878;
  assign n43884 = ~n43863 & ~n60799;
  assign n43885 = ~pi221 & ~n43884;
  assign n43886 = ~n60798 & ~n43885;
  assign n43887 = ~pi215 & ~n43886;
  assign n43888 = pi215 & pi1135;
  assign n43889 = pi299 & ~n43888;
  assign n43890 = ~n43887 & n43889;
  assign n43891 = pi223 & pi1135;
  assign n43892 = ~pi299 & ~n43891;
  assign n43893 = ~pi938 & n38636;
  assign n43894 = ~pi1135 & ~n38636;
  assign n43895 = pi222 & ~n43894;
  assign n43896 = pi222 & ~n43893;
  assign n43897 = ~n43894 & n43896;
  assign n43898 = ~n43893 & n43895;
  assign n43899 = ~pi224 & ~pi879;
  assign n43900 = ~n28313 & n43899;
  assign n43901 = pi224 & ~pi279;
  assign n43902 = ~pi222 & ~n43901;
  assign n43903 = ~n43900 & n43902;
  assign n43904 = ~n60800 & ~n43903;
  assign n43905 = ~pi223 & ~n43904;
  assign n43906 = ~n43640 & n43905;
  assign n43907 = n43892 & ~n43906;
  assign n43908 = ~pi39 & ~n43907;
  assign n43909 = ~n43890 & n43908;
  assign n43910 = ~n43891 & ~n43905;
  assign n43911 = ~pi299 & ~n43910;
  assign n43912 = n35583 & ~n43872;
  assign n43913 = n43911 & ~n43912;
  assign n43914 = pi228 & n43875;
  assign n43915 = ~pi879 & n58822;
  assign n43916 = pi161 & ~pi228;
  assign n43917 = ~n31586 & ~n43916;
  assign n43918 = ~n43915 & ~n43917;
  assign n43919 = ~n43914 & ~n43918;
  assign n43920 = ~pi216 & ~n43919;
  assign n43921 = ~n43863 & ~n43920;
  assign n43922 = ~pi221 & ~n43921;
  assign n43923 = ~n60798 & ~n43922;
  assign n43924 = ~pi215 & ~n43923;
  assign n43925 = ~n43888 & ~n43924;
  assign n43926 = pi299 & ~n43925;
  assign n43927 = ~n43913 & ~n43926;
  assign n43928 = pi39 & ~n43927;
  assign n43929 = ~pi38 & ~n43928;
  assign n43930 = ~n43909 & n43929;
  assign n43931 = ~n43914 & ~n43916;
  assign n43932 = ~pi216 & ~n43931;
  assign n43933 = ~n43863 & ~n43932;
  assign n43934 = ~pi221 & ~n43933;
  assign n43935 = ~n60798 & ~n43934;
  assign n43936 = ~pi215 & ~n43935;
  assign n43937 = ~n43888 & ~n43936;
  assign n43938 = pi299 & ~n43937;
  assign n43939 = ~n43913 & ~n43938;
  assign n43940 = pi38 & n43939;
  assign n43941 = ~pi100 & ~n43940;
  assign n43942 = ~n43930 & n43941;
  assign n43943 = ~pi879 & n41433;
  assign n43944 = pi161 & ~n43943;
  assign n43945 = ~pi152 & ~pi166;
  assign n43946 = ~n41433 & ~n43945;
  assign n43947 = ~n28550 & n43945;
  assign n43948 = pi879 & ~n43947;
  assign n43949 = ~n43946 & n43948;
  assign n43950 = ~n43944 & ~n43949;
  assign n43951 = ~pi228 & ~n43950;
  assign n43952 = ~n43914 & ~n43951;
  assign n43953 = ~pi216 & ~n43952;
  assign n43954 = ~n43863 & ~n43953;
  assign n43955 = ~pi221 & ~n43954;
  assign n43956 = ~n60798 & ~n43955;
  assign n43957 = ~pi215 & ~n43956;
  assign n43958 = ~n43888 & ~n43957;
  assign n43959 = pi299 & ~n43958;
  assign n43960 = n2634 & ~n43913;
  assign n43961 = ~n43959 & n43960;
  assign n43962 = ~n2634 & n43939;
  assign n43963 = pi100 & ~n43962;
  assign n43964 = ~n43961 & n43963;
  assign n43965 = ~n43942 & ~n43964;
  assign n43966 = ~pi87 & ~n43965;
  assign n43967 = ~n58815 & n43939;
  assign n43968 = n58815 & n43927;
  assign n43969 = ~n43967 & ~n43968;
  assign n43970 = pi87 & n43969;
  assign n43971 = ~pi75 & ~n43970;
  assign n43972 = ~n43966 & n43971;
  assign n43973 = pi75 & n43939;
  assign n43974 = ~pi92 & ~n43973;
  assign n43975 = ~n43972 & n43974;
  assign n43976 = n6309 & ~n43969;
  assign n43977 = ~n6309 & n43939;
  assign n43978 = pi92 & ~n43977;
  assign n43979 = ~n43976 & n43978;
  assign n43980 = n6306 & ~n43979;
  assign n43981 = ~n43975 & n43980;
  assign n43982 = ~n6306 & n43939;
  assign n43983 = ~pi55 & ~n43982;
  assign n43984 = ~n43981 & n43983;
  assign n43985 = n28288 & n43925;
  assign n43986 = ~n28288 & n43937;
  assign n43987 = pi55 & ~n43986;
  assign n43988 = ~n43985 & n43987;
  assign n43989 = ~pi56 & ~n43988;
  assign n43990 = ~n43984 & n43989;
  assign n43991 = n60070 & ~n43925;
  assign n43992 = ~n60070 & ~n43937;
  assign n43993 = pi56 & ~n43992;
  assign n43994 = ~n60070 & n43937;
  assign n43995 = ~pi55 & n43985;
  assign n43996 = ~n43994 & ~n43995;
  assign n43997 = pi56 & ~n43996;
  assign n43998 = ~n43991 & n43993;
  assign n43999 = ~pi62 & ~n60801;
  assign n44000 = ~n43990 & n43999;
  assign n44001 = n41492 & n43925;
  assign n44002 = ~n41492 & n43937;
  assign n44003 = pi62 & ~n44002;
  assign n44004 = ~n44001 & n44003;
  assign n44005 = n4438 & ~n44004;
  assign n44006 = ~n44000 & n44005;
  assign n44007 = ~n4438 & n43937;
  assign n44008 = ~pi244 & ~n44007;
  assign n44009 = ~n44006 & n44008;
  assign n44010 = ~pi161 & ~n40748;
  assign n44011 = pi879 & ~n44010;
  assign n44012 = pi161 & n41335;
  assign n44013 = ~pi161 & ~n41346;
  assign n44014 = ~pi879 & ~n44013;
  assign n44015 = ~n44012 & n44014;
  assign n44016 = ~pi228 & ~n44015;
  assign n44017 = ~pi228 & ~n44011;
  assign n44018 = ~n44015 & n44017;
  assign n44019 = ~n44011 & n44016;
  assign n44020 = n43877 & ~n60802;
  assign n44021 = ~n43863 & ~n44020;
  assign n44022 = ~pi221 & ~n44021;
  assign n44023 = ~n60798 & ~n44022;
  assign n44024 = ~pi215 & ~n44023;
  assign n44025 = n43889 & ~n44024;
  assign n44026 = ~n43640 & n43904;
  assign n44027 = ~pi223 & ~n44026;
  assign n44028 = n43892 & ~n44027;
  assign n44029 = ~pi39 & ~n44028;
  assign n44030 = ~n44025 & n44029;
  assign n44031 = ~n41403 & ~n43914;
  assign n44032 = ~n43918 & n44031;
  assign n44033 = ~pi216 & ~n44032;
  assign n44034 = ~n43863 & ~n44033;
  assign n44035 = ~pi221 & ~n44034;
  assign n44036 = ~n60798 & ~n44035;
  assign n44037 = ~pi215 & ~n44036;
  assign n44038 = ~n43888 & ~n44037;
  assign n44039 = pi299 & ~n44038;
  assign n44040 = ~n43911 & ~n44039;
  assign n44041 = pi39 & ~n44040;
  assign n44042 = ~pi38 & ~n44041;
  assign n44043 = ~n44030 & n44042;
  assign n44044 = ~n41418 & n43937;
  assign n44045 = pi299 & ~n44044;
  assign n44046 = ~n43911 & ~n44045;
  assign n44047 = pi38 & n44046;
  assign n44048 = ~pi100 & ~n44047;
  assign n44049 = ~n44043 & n44048;
  assign n44050 = ~n43951 & n44031;
  assign n44051 = ~pi216 & ~n44050;
  assign n44052 = ~n43863 & ~n44051;
  assign n44053 = ~pi221 & ~n44052;
  assign n44054 = ~n60798 & ~n44053;
  assign n44055 = ~pi215 & ~n44054;
  assign n44056 = ~n43888 & ~n44055;
  assign n44057 = pi299 & ~n44056;
  assign n44058 = n2634 & ~n43911;
  assign n44059 = ~n44057 & n44058;
  assign n44060 = ~n2634 & n44046;
  assign n44061 = pi100 & ~n44060;
  assign n44062 = ~n44059 & n44061;
  assign n44063 = ~n44049 & ~n44062;
  assign n44064 = ~pi87 & ~n44063;
  assign n44065 = ~n58815 & n44046;
  assign n44066 = n58815 & n44040;
  assign n44067 = ~n44065 & ~n44066;
  assign n44068 = pi87 & n44067;
  assign n44069 = ~pi75 & ~n44068;
  assign n44070 = ~n44064 & n44069;
  assign n44071 = pi75 & n44046;
  assign n44072 = ~pi92 & ~n44071;
  assign n44073 = ~n44070 & n44072;
  assign n44074 = n6309 & ~n44067;
  assign n44075 = ~n6309 & n44046;
  assign n44076 = pi92 & ~n44075;
  assign n44077 = ~n44074 & n44076;
  assign n44078 = n6306 & ~n44077;
  assign n44079 = ~n44073 & n44078;
  assign n44080 = ~n6306 & n44046;
  assign n44081 = ~pi55 & ~n44080;
  assign n44082 = ~n44079 & n44081;
  assign n44083 = n28288 & n44038;
  assign n44084 = ~n28288 & n44044;
  assign n44085 = pi55 & ~n44084;
  assign n44086 = ~n44083 & n44085;
  assign n44087 = ~pi56 & ~n44086;
  assign n44088 = ~n44082 & n44087;
  assign n44089 = n60070 & ~n44038;
  assign n44090 = ~n60070 & ~n44044;
  assign n44091 = pi56 & ~n44090;
  assign n44092 = ~pi55 & n44083;
  assign n44093 = ~n60070 & n44044;
  assign n44094 = ~n44092 & ~n44093;
  assign n44095 = pi56 & ~n44094;
  assign n44096 = ~n44089 & n44091;
  assign n44097 = ~pi62 & ~n60803;
  assign n44098 = ~n44088 & n44097;
  assign n44099 = n41492 & n44038;
  assign n44100 = ~n41492 & n44044;
  assign n44101 = pi62 & ~n44100;
  assign n44102 = ~n44099 & n44101;
  assign n44103 = n4438 & ~n44102;
  assign n44104 = ~n44098 & n44103;
  assign n44105 = ~n4438 & n44044;
  assign n44106 = pi244 & ~n44105;
  assign n44107 = ~n44104 & n44106;
  assign n44108 = ~n44009 & ~n44107;
  assign n44109 = pi833 & ~pi930;
  assign n44110 = n2850 & n44109;
  assign n44111 = pi216 & pi278;
  assign n44112 = ~pi221 & ~n44111;
  assign n44113 = ~pi105 & pi152;
  assign n44114 = pi228 & ~n44113;
  assign n44115 = ~pi846 & n41340;
  assign n44116 = pi105 & ~n44115;
  assign n44117 = n44114 & ~n44116;
  assign n44118 = ~pi216 & ~n44117;
  assign n44119 = pi152 & ~n41335;
  assign n44120 = ~pi152 & n41346;
  assign n44121 = ~pi846 & ~n44120;
  assign n44122 = ~n44119 & n44121;
  assign n44123 = ~pi152 & pi846;
  assign n44124 = ~n40748 & n44123;
  assign n44125 = ~n44122 & ~n44124;
  assign n44126 = ~pi228 & ~n44125;
  assign n44127 = n44118 & ~n44126;
  assign n44128 = n44112 & ~n44127;
  assign n44129 = ~n44110 & ~n44128;
  assign n44130 = pi221 & ~n38221;
  assign n44131 = n2851 & ~n44130;
  assign n44132 = n44129 & n44131;
  assign n44133 = pi224 & pi278;
  assign n44134 = ~pi222 & ~n44133;
  assign n44135 = ~pi224 & ~n44115;
  assign n44136 = n44134 & ~n44135;
  assign n44137 = n2827 & n44109;
  assign n44138 = n2828 & ~n38637;
  assign n44139 = ~n44137 & n44138;
  assign n44140 = ~n44136 & ~n44137;
  assign n44141 = n44138 & n44140;
  assign n44142 = ~n44136 & n44139;
  assign n44143 = ~pi39 & ~n60804;
  assign n44144 = ~n44132 & n44143;
  assign n44145 = pi846 & ~n28313;
  assign n44146 = ~pi224 & n44145;
  assign n44147 = n44134 & ~n44146;
  assign n44148 = n38638 & ~n44137;
  assign n44149 = ~n44147 & n44148;
  assign n44150 = ~pi299 & ~n44149;
  assign n44151 = ~n41391 & n44150;
  assign n44152 = ~pi215 & ~n44130;
  assign n44153 = ~n44110 & n44152;
  assign n44154 = pi105 & n44145;
  assign n44155 = ~n44113 & ~n44154;
  assign n44156 = pi228 & ~n44155;
  assign n44157 = ~n41403 & ~n44156;
  assign n44158 = ~pi846 & n58822;
  assign n44159 = ~pi152 & ~n58822;
  assign n44160 = ~pi228 & ~n44159;
  assign n44161 = ~pi228 & ~n44158;
  assign n44162 = ~n44159 & n44161;
  assign n44163 = ~n44158 & n44160;
  assign n44164 = n44157 & ~n60805;
  assign n44165 = ~pi216 & ~n44164;
  assign n44166 = n44112 & ~n44165;
  assign n44167 = n44153 & ~n44166;
  assign n44168 = pi299 & ~n44167;
  assign n44169 = ~n44151 & ~n44168;
  assign n44170 = pi39 & ~n44169;
  assign n44171 = ~pi38 & ~n44170;
  assign n44172 = ~n44144 & n44171;
  assign n44173 = pi152 & ~pi228;
  assign n44174 = ~n44156 & ~n44173;
  assign n44175 = ~pi216 & ~n44174;
  assign n44176 = n44112 & ~n44175;
  assign n44177 = n44153 & ~n44176;
  assign n44178 = ~n41418 & ~n44177;
  assign n44179 = pi299 & n44178;
  assign n44180 = ~n44151 & ~n44179;
  assign n44181 = pi38 & n44180;
  assign n44182 = ~pi100 & ~n44181;
  assign n44183 = ~n44172 & n44182;
  assign n44184 = pi846 & ~n41438;
  assign n44185 = ~n41434 & ~n44184;
  assign n44186 = ~pi228 & ~n44185;
  assign n44187 = n44157 & ~n44186;
  assign n44188 = ~pi216 & ~n44187;
  assign n44189 = n44112 & ~n44188;
  assign n44190 = n44153 & ~n44189;
  assign n44191 = pi299 & ~n44190;
  assign n44192 = n2634 & ~n44151;
  assign n44193 = ~n44191 & n44192;
  assign n44194 = ~n2634 & n44180;
  assign n44195 = pi100 & ~n44194;
  assign n44196 = ~n44193 & n44195;
  assign n44197 = ~n44183 & ~n44196;
  assign n44198 = ~pi87 & ~n44197;
  assign n44199 = ~n58815 & n44180;
  assign n44200 = n58815 & n44169;
  assign n44201 = ~n44199 & ~n44200;
  assign n44202 = pi87 & n44201;
  assign n44203 = ~pi75 & ~n44202;
  assign n44204 = ~n44198 & n44203;
  assign n44205 = pi75 & n44180;
  assign n44206 = ~pi92 & ~n44205;
  assign n44207 = ~n44204 & n44206;
  assign n44208 = n6309 & ~n44201;
  assign n44209 = ~n6309 & n44180;
  assign n44210 = pi92 & ~n44209;
  assign n44211 = ~n44208 & n44210;
  assign n44212 = n6306 & ~n44211;
  assign n44213 = ~n44207 & n44212;
  assign n44214 = ~n6306 & n44180;
  assign n44215 = ~pi55 & ~n44214;
  assign n44216 = ~n44213 & n44215;
  assign n44217 = n28288 & n44167;
  assign n44218 = ~n28288 & ~n44178;
  assign n44219 = pi55 & ~n44218;
  assign n44220 = ~n44217 & n44219;
  assign n44221 = ~pi56 & ~n44220;
  assign n44222 = ~n44216 & n44221;
  assign n44223 = n60070 & ~n44167;
  assign n44224 = ~n60070 & n44178;
  assign n44225 = pi56 & ~n44224;
  assign n44226 = ~n60070 & ~n44178;
  assign n44227 = ~pi55 & n44217;
  assign n44228 = ~n44226 & ~n44227;
  assign n44229 = pi56 & ~n44228;
  assign n44230 = ~n44223 & n44225;
  assign n44231 = ~pi62 & ~n60806;
  assign n44232 = ~n44222 & n44231;
  assign n44233 = n41492 & n44167;
  assign n44234 = ~n41492 & ~n44178;
  assign n44235 = pi62 & ~n44234;
  assign n44236 = ~n44233 & n44235;
  assign n44237 = n4438 & ~n44236;
  assign n44238 = ~n44232 & n44237;
  assign n44239 = ~n4438 & ~n44178;
  assign n44240 = pi242 & ~n44239;
  assign n44241 = ~n44238 & n44240;
  assign n44242 = ~pi152 & ~n41335;
  assign n44243 = pi152 & n41346;
  assign n44244 = pi846 & ~n44243;
  assign n44245 = ~n44242 & n44244;
  assign n44246 = pi152 & ~pi846;
  assign n44247 = ~n40748 & n44246;
  assign n44248 = ~pi228 & ~n44247;
  assign n44249 = ~n44245 & n44248;
  assign n44250 = ~n41340 & n44114;
  assign n44251 = n44118 & ~n44250;
  assign n44252 = ~n44249 & n44251;
  assign n44253 = n44112 & ~n44252;
  assign n44254 = ~n44110 & ~n44253;
  assign n44255 = n44131 & n44254;
  assign n44256 = ~n41339 & n44146;
  assign n44257 = n44134 & ~n44256;
  assign n44258 = n44139 & ~n44257;
  assign n44259 = ~pi39 & ~n44258;
  assign n44260 = ~n44255 & n44259;
  assign n44261 = ~n44156 & ~n60805;
  assign n44262 = ~pi216 & ~n44261;
  assign n44263 = n44112 & ~n44262;
  assign n44264 = n44153 & ~n44263;
  assign n44265 = pi299 & ~n44264;
  assign n44266 = ~n44150 & ~n44265;
  assign n44267 = pi39 & ~n44266;
  assign n44268 = ~pi38 & ~n44267;
  assign n44269 = ~n44260 & n44268;
  assign n44270 = pi299 & ~n44177;
  assign n44271 = ~n44150 & ~n44270;
  assign n44272 = pi38 & n44271;
  assign n44273 = ~pi100 & ~n44272;
  assign n44274 = ~n44269 & n44273;
  assign n44275 = ~n44156 & ~n44186;
  assign n44276 = ~pi216 & ~n44275;
  assign n44277 = n44112 & ~n44276;
  assign n44278 = n44153 & ~n44277;
  assign n44279 = pi299 & ~n44278;
  assign n44280 = n2634 & ~n44150;
  assign n44281 = ~n44279 & n44280;
  assign n44282 = ~n2634 & n44271;
  assign n44283 = pi100 & ~n44282;
  assign n44284 = ~n44281 & n44283;
  assign n44285 = ~n44274 & ~n44284;
  assign n44286 = ~pi87 & ~n44285;
  assign n44287 = ~n58815 & n44271;
  assign n44288 = n58815 & n44266;
  assign n44289 = ~n44287 & ~n44288;
  assign n44290 = pi87 & n44289;
  assign n44291 = ~pi75 & ~n44290;
  assign n44292 = ~n44286 & n44291;
  assign n44293 = pi75 & n44271;
  assign n44294 = ~pi92 & ~n44293;
  assign n44295 = ~n44292 & n44294;
  assign n44296 = n6309 & ~n44289;
  assign n44297 = ~n6309 & n44271;
  assign n44298 = pi92 & ~n44297;
  assign n44299 = ~n44296 & n44298;
  assign n44300 = n6306 & ~n44299;
  assign n44301 = ~n44295 & n44300;
  assign n44302 = ~n6306 & n44271;
  assign n44303 = ~pi55 & ~n44302;
  assign n44304 = ~n44301 & n44303;
  assign n44305 = n28288 & n44264;
  assign n44306 = ~n28288 & n44177;
  assign n44307 = pi55 & ~n44306;
  assign n44308 = ~n44305 & n44307;
  assign n44309 = ~pi56 & ~n44308;
  assign n44310 = ~n44304 & n44309;
  assign n44311 = n60070 & ~n44264;
  assign n44312 = ~n60070 & ~n44177;
  assign n44313 = pi56 & ~n44312;
  assign n44314 = ~n60070 & n44177;
  assign n44315 = ~pi55 & n44305;
  assign n44316 = ~n44314 & ~n44315;
  assign n44317 = pi56 & ~n44316;
  assign n44318 = ~n44311 & n44313;
  assign n44319 = ~pi62 & ~n60807;
  assign n44320 = ~n44310 & n44319;
  assign n44321 = n41492 & n44264;
  assign n44322 = ~n41492 & n44177;
  assign n44323 = pi62 & ~n44322;
  assign n44324 = ~n44321 & n44323;
  assign n44325 = n4438 & ~n44324;
  assign n44326 = ~n44320 & n44325;
  assign n44327 = ~n4438 & n44177;
  assign n44328 = ~pi242 & ~n44327;
  assign n44329 = ~n44326 & n44328;
  assign n44330 = ~n44241 & ~n44329;
  assign n44331 = ~pi1134 & ~n44330;
  assign n44332 = n2828 & ~n44140;
  assign n44333 = ~pi39 & ~n44332;
  assign n44334 = n2851 & ~n44129;
  assign n44335 = n44333 & ~n44334;
  assign n44336 = n38638 & n44151;
  assign n44337 = ~pi299 & ~n44336;
  assign n44338 = ~n44110 & ~n44166;
  assign n44339 = ~pi215 & ~n44338;
  assign n44340 = pi299 & ~n44339;
  assign n44341 = ~n44337 & ~n44340;
  assign n44342 = pi39 & ~n44341;
  assign n44343 = ~pi38 & ~n44342;
  assign n44344 = ~n44335 & n44343;
  assign n44345 = ~n44110 & ~n44176;
  assign n44346 = ~pi215 & ~n44345;
  assign n44347 = ~n41418 & n44346;
  assign n44348 = pi299 & ~n44347;
  assign n44349 = ~n44337 & ~n44348;
  assign n44350 = pi38 & n44349;
  assign n44351 = ~pi100 & ~n44350;
  assign n44352 = ~n44344 & n44351;
  assign n44353 = ~n44110 & ~n44189;
  assign n44354 = ~pi215 & ~n44353;
  assign n44355 = pi299 & ~n44354;
  assign n44356 = n2634 & ~n44337;
  assign n44357 = ~n44355 & n44356;
  assign n44358 = ~n2634 & n44349;
  assign n44359 = pi100 & ~n44358;
  assign n44360 = ~n44357 & n44359;
  assign n44361 = ~n44352 & ~n44360;
  assign n44362 = ~pi87 & ~n44361;
  assign n44363 = ~n58815 & n44349;
  assign n44364 = n58815 & n44341;
  assign n44365 = ~n44363 & ~n44364;
  assign n44366 = pi87 & n44365;
  assign n44367 = ~pi75 & ~n44366;
  assign n44368 = ~n44362 & n44367;
  assign n44369 = pi75 & n44349;
  assign n44370 = ~pi92 & ~n44369;
  assign n44371 = ~n44368 & n44370;
  assign n44372 = n6309 & ~n44365;
  assign n44373 = ~n6309 & n44349;
  assign n44374 = pi92 & ~n44373;
  assign n44375 = ~n44372 & n44374;
  assign n44376 = n6306 & ~n44375;
  assign n44377 = ~n44371 & n44376;
  assign n44378 = ~n6306 & n44349;
  assign n44379 = ~pi55 & ~n44378;
  assign n44380 = ~n44377 & n44379;
  assign n44381 = n28288 & n44339;
  assign n44382 = ~n28288 & n44347;
  assign n44383 = pi55 & ~n44382;
  assign n44384 = ~n44381 & n44383;
  assign n44385 = ~pi56 & ~n44384;
  assign n44386 = ~n44380 & n44385;
  assign n44387 = n60070 & ~n44339;
  assign n44388 = ~n60070 & ~n44347;
  assign n44389 = pi56 & ~n44388;
  assign n44390 = ~pi55 & n44381;
  assign n44391 = ~n60070 & n44347;
  assign n44392 = ~n44390 & ~n44391;
  assign n44393 = pi56 & ~n44392;
  assign n44394 = ~n44387 & n44389;
  assign n44395 = ~pi62 & ~n60808;
  assign n44396 = ~n44386 & n44395;
  assign n44397 = n41492 & n44339;
  assign n44398 = ~n41492 & n44347;
  assign n44399 = pi62 & ~n44398;
  assign n44400 = ~n44397 & n44399;
  assign n44401 = n4438 & ~n44400;
  assign n44402 = ~n44396 & n44401;
  assign n44403 = ~n4438 & n44347;
  assign n44404 = pi242 & ~n44403;
  assign n44405 = ~n44402 & n44404;
  assign n44406 = n2851 & ~n44254;
  assign n44407 = n2828 & n44257;
  assign n44408 = n44333 & ~n44407;
  assign n44409 = ~n44406 & n44408;
  assign n44410 = ~pi223 & n44147;
  assign n44411 = n44337 & ~n44410;
  assign n44412 = ~n44110 & ~n44263;
  assign n44413 = ~pi215 & ~n44412;
  assign n44414 = pi299 & ~n44413;
  assign n44415 = ~n44411 & ~n44414;
  assign n44416 = pi39 & ~n44415;
  assign n44417 = ~pi38 & ~n44416;
  assign n44418 = ~n44409 & n44417;
  assign n44419 = pi299 & ~n44346;
  assign n44420 = ~n44411 & ~n44419;
  assign n44421 = pi38 & n44420;
  assign n44422 = ~pi100 & ~n44421;
  assign n44423 = ~n44418 & n44422;
  assign n44424 = ~n44110 & ~n44277;
  assign n44425 = ~pi215 & ~n44424;
  assign n44426 = pi299 & ~n44425;
  assign n44427 = n2634 & ~n44411;
  assign n44428 = ~n44426 & n44427;
  assign n44429 = ~n2634 & n44420;
  assign n44430 = pi100 & ~n44429;
  assign n44431 = ~n44428 & n44430;
  assign n44432 = ~n44423 & ~n44431;
  assign n44433 = ~pi87 & ~n44432;
  assign n44434 = ~n58815 & n44420;
  assign n44435 = n58815 & n44415;
  assign n44436 = ~n44434 & ~n44435;
  assign n44437 = pi87 & n44436;
  assign n44438 = ~pi75 & ~n44437;
  assign n44439 = ~n44433 & n44438;
  assign n44440 = pi75 & n44420;
  assign n44441 = ~pi92 & ~n44440;
  assign n44442 = ~n44439 & n44441;
  assign n44443 = n6309 & ~n44436;
  assign n44444 = ~n6309 & n44420;
  assign n44445 = pi92 & ~n44444;
  assign n44446 = ~n44443 & n44445;
  assign n44447 = n6306 & ~n44446;
  assign n44448 = ~n44442 & n44447;
  assign n44449 = ~n6306 & n44420;
  assign n44450 = ~pi55 & ~n44449;
  assign n44451 = ~n44448 & n44450;
  assign n44452 = n28288 & n44413;
  assign n44453 = ~n28288 & n44346;
  assign n44454 = pi55 & ~n44453;
  assign n44455 = ~n44452 & n44454;
  assign n44456 = ~pi56 & ~n44455;
  assign n44457 = ~n44451 & n44456;
  assign n44458 = n60070 & ~n44413;
  assign n44459 = ~n60070 & ~n44346;
  assign n44460 = pi56 & ~n44459;
  assign n44461 = ~n60070 & n44346;
  assign n44462 = ~pi55 & n44452;
  assign n44463 = ~n44461 & ~n44462;
  assign n44464 = pi56 & ~n44463;
  assign n44465 = ~n44458 & n44460;
  assign n44466 = ~pi62 & ~n60809;
  assign n44467 = ~n44457 & n44466;
  assign n44468 = n41492 & n44413;
  assign n44469 = ~n41492 & n44346;
  assign n44470 = pi62 & ~n44469;
  assign n44471 = ~n44468 & n44470;
  assign n44472 = n4438 & ~n44471;
  assign n44473 = ~n44467 & n44472;
  assign n44474 = ~n4438 & n44346;
  assign n44475 = ~pi242 & ~n44474;
  assign n44476 = ~n44473 & n44475;
  assign n44477 = pi1134 & ~n44476;
  assign n44478 = ~n44405 & n44477;
  assign po165 = ~n44331 & ~n44478;
  assign n44480 = ~pi39 & ~n39068;
  assign n44481 = pi39 & ~n39688;
  assign n44482 = n2636 & ~n44481;
  assign n44483 = ~n44480 & n44482;
  assign n44484 = ~n40231 & ~n44483;
  assign n44485 = ~pi87 & ~n44484;
  assign n44486 = n60561 & ~n44485;
  assign n44487 = ~n60561 & ~n38944;
  assign n44488 = n38939 & ~n44487;
  assign n44489 = n38938 & n44488;
  assign n44490 = ~n60561 & n38944;
  assign n44491 = n6310 & n32859;
  assign n44492 = ~n44484 & n44491;
  assign n44493 = ~n44490 & ~n44492;
  assign n44494 = n38938 & n38939;
  assign n44495 = ~n44493 & n44494;
  assign n44496 = ~n44486 & n44489;
  assign n44497 = n28288 & ~n36439;
  assign n44498 = ~n3871 & n44497;
  assign n44499 = pi286 & n44498;
  assign n44500 = pi288 & pi289;
  assign n44501 = n44499 & n44500;
  assign n44502 = pi285 & n44497;
  assign n44503 = ~n44501 & ~n44502;
  assign n44504 = pi285 & n44501;
  assign n44505 = n58992 & ~n44504;
  assign n44506 = ~n44503 & n44505;
  assign n44507 = n58992 & n44501;
  assign n44508 = ~pi286 & n3871;
  assign n44509 = ~pi288 & n44508;
  assign n44510 = ~pi289 & n44509;
  assign n44511 = pi285 & ~n44510;
  assign n44512 = ~n44507 & n44511;
  assign n44513 = ~n44506 & ~n44512;
  assign po442 = ~pi793 & ~n44513;
  assign n44515 = ~pi286 & ~n44498;
  assign n44516 = pi288 & ~n44499;
  assign n44517 = ~n44515 & n44516;
  assign n44518 = ~pi288 & ~n3212;
  assign n44519 = n3871 & ~n44497;
  assign n44520 = pi286 & ~n44519;
  assign n44521 = ~n44497 & n44508;
  assign n44522 = ~n44520 & ~n44521;
  assign n44523 = n44518 & ~n44522;
  assign n44524 = n58992 & ~n44523;
  assign n44525 = ~n44517 & n44524;
  assign n44526 = n3871 & n44518;
  assign n44527 = ~pi286 & n44526;
  assign n44528 = pi286 & ~n44526;
  assign n44529 = ~n58992 & ~n44528;
  assign n44530 = ~n44527 & n44529;
  assign n44531 = ~pi793 & ~n44530;
  assign po443 = ~n44525 & n44531;
  assign n44533 = pi288 & ~n3871;
  assign n44534 = ~n44526 & ~n44533;
  assign n44535 = n58992 & n44497;
  assign n44536 = ~n36439 & n60562;
  assign n44537 = n44534 & ~po637;
  assign n44538 = ~n44534 & po637;
  assign n44539 = ~pi793 & ~n44538;
  assign po445 = ~n44537 & n44539;
  assign n44541 = pi289 & ~n44521;
  assign n44542 = pi285 & ~pi289;
  assign n44543 = n44521 & n44542;
  assign n44544 = ~pi288 & ~n44543;
  assign n44545 = ~n44541 & n44544;
  assign n44546 = ~pi289 & n44516;
  assign n44547 = ~n44501 & ~n44546;
  assign n44548 = ~n44545 & n44547;
  assign n44549 = n58992 & ~n44548;
  assign n44550 = n44509 & n44542;
  assign n44551 = pi289 & ~n44509;
  assign n44552 = ~n58992 & ~n44551;
  assign n44553 = ~n44550 & n44552;
  assign n44554 = ~pi793 & ~n44553;
  assign po446 = ~n44549 & n44554;
  assign n44556 = pi233 & pi237;
  assign n44557 = ~pi332 & ~n2778;
  assign n44558 = ~pi947 & ~n44557;
  assign n44559 = pi96 & pi210;
  assign n44560 = pi332 & n44559;
  assign n44561 = ~pi32 & pi70;
  assign n44562 = ~pi70 & ~pi841;
  assign n44563 = pi32 & n44562;
  assign n44564 = ~n44561 & ~n44563;
  assign n44565 = ~pi210 & ~n44564;
  assign n44566 = ~pi32 & ~pi96;
  assign n44567 = pi70 & n44566;
  assign n44568 = ~pi332 & ~n44567;
  assign n44569 = ~n44565 & n44568;
  assign n44570 = ~n44560 & ~n44569;
  assign n44571 = ~n2680 & n44570;
  assign n44572 = n2778 & ~n44571;
  assign n44573 = n44558 & ~n44572;
  assign n44574 = pi332 & pi468;
  assign n44575 = ~pi468 & ~n44569;
  assign n44576 = ~n44574 & ~n44575;
  assign n44577 = ~n2778 & n44576;
  assign n44578 = n2778 & ~n44570;
  assign n44579 = pi947 & ~n44578;
  assign n44580 = ~n44577 & n44579;
  assign n44581 = ~n44573 & ~n44580;
  assign n44582 = ~n28288 & n44581;
  assign n44583 = ~pi95 & n60582;
  assign n44584 = ~pi70 & ~n44583;
  assign n44585 = n44566 & ~n44584;
  assign n44586 = pi210 & n44585;
  assign n44587 = ~pi95 & n2597;
  assign n44588 = pi32 & ~n44562;
  assign n44589 = ~pi96 & ~n44588;
  assign n44590 = ~pi95 & n2601;
  assign n44591 = ~n44588 & n44590;
  assign n44592 = n44587 & n44589;
  assign n44593 = n6343 & n60812;
  assign n44594 = n58807 & n44593;
  assign n44595 = n44564 & ~n44594;
  assign n44596 = ~pi210 & ~n44595;
  assign n44597 = ~pi332 & ~n44596;
  assign n44598 = ~n44586 & n44597;
  assign n44599 = ~n44560 & ~n44598;
  assign n44600 = ~n2680 & n44599;
  assign n44601 = n2778 & ~n44600;
  assign n44602 = n44558 & ~n44601;
  assign n44603 = ~pi468 & ~n44598;
  assign n44604 = ~n44574 & ~n44603;
  assign n44605 = ~n2778 & n44604;
  assign n44606 = n2778 & ~n44599;
  assign n44607 = pi947 & ~n44606;
  assign n44608 = ~n44605 & n44607;
  assign n44609 = ~n44602 & ~n44608;
  assign n44610 = n28288 & n44609;
  assign n44611 = ~n44582 & ~n44610;
  assign n44612 = n4440 & ~n44611;
  assign n44613 = ~n4440 & n44581;
  assign n44614 = pi59 & ~n44613;
  assign n44615 = ~n44612 & n44614;
  assign n44616 = n2614 & n38298;
  assign n44617 = n44587 & n44616;
  assign n44618 = ~pi70 & ~n44617;
  assign n44619 = n44566 & ~n44618;
  assign n44620 = pi210 & n44619;
  assign n44621 = n60812 & n44616;
  assign n44622 = n44564 & ~n44621;
  assign n44623 = ~pi210 & ~n44622;
  assign n44624 = ~pi332 & ~n44623;
  assign n44625 = ~n44620 & n44624;
  assign n44626 = ~n44560 & ~n44625;
  assign n44627 = ~n2680 & n44626;
  assign n44628 = n2778 & ~n44627;
  assign n44629 = n44558 & ~n44628;
  assign n44630 = ~pi468 & ~n44625;
  assign n44631 = ~n44574 & ~n44630;
  assign n44632 = ~n2778 & n44631;
  assign n44633 = n2778 & ~n44626;
  assign n44634 = pi947 & ~n44633;
  assign n44635 = ~n44632 & n44634;
  assign n44636 = n31592 & ~n44635;
  assign n44637 = ~n44629 & n44636;
  assign n44638 = n40694 & n44609;
  assign n44639 = pi299 & ~n44638;
  assign n44640 = ~n44637 & n44639;
  assign n44641 = pi96 & pi198;
  assign n44642 = pi332 & n44641;
  assign n44643 = pi198 & n44619;
  assign n44644 = ~pi198 & ~n44622;
  assign n44645 = ~pi332 & ~n44644;
  assign n44646 = ~n44643 & n44645;
  assign n44647 = ~n44642 & ~n44646;
  assign n44648 = n2778 & ~n44647;
  assign n44649 = ~pi468 & ~n44646;
  assign n44650 = ~n2778 & ~n44574;
  assign n44651 = ~n44649 & n44650;
  assign n44652 = pi587 & ~n44651;
  assign n44653 = ~pi587 & ~n44557;
  assign n44654 = n2680 & n2778;
  assign n44655 = n44653 & ~n44654;
  assign n44656 = ~n44652 & ~n44655;
  assign n44657 = ~n44648 & ~n44656;
  assign n44658 = n31592 & ~n44657;
  assign n44659 = pi198 & n44585;
  assign n44660 = ~pi198 & ~n44595;
  assign n44661 = ~pi332 & ~n44660;
  assign n44662 = ~n44659 & n44661;
  assign n44663 = ~n44642 & ~n44662;
  assign n44664 = n2778 & ~n44663;
  assign n44665 = ~pi468 & ~n44662;
  assign n44666 = n44650 & ~n44665;
  assign n44667 = pi587 & ~n44666;
  assign n44668 = pi587 & ~n44664;
  assign n44669 = ~n44666 & n44668;
  assign n44670 = ~n44664 & n44667;
  assign n44671 = ~n2680 & n44663;
  assign n44672 = n2778 & ~n44671;
  assign n44673 = n44653 & ~n44672;
  assign n44674 = n40694 & ~n44673;
  assign n44675 = ~n60813 & n44674;
  assign n44676 = ~pi299 & ~n44675;
  assign n44677 = ~n44658 & n44676;
  assign n44678 = ~pi74 & ~n44677;
  assign n44679 = pi299 & ~n44635;
  assign n44680 = pi299 & ~n44629;
  assign n44681 = ~n44635 & n44680;
  assign n44682 = ~n44629 & n44679;
  assign n44683 = ~n2680 & n44647;
  assign n44684 = n2778 & ~n44683;
  assign n44685 = n44653 & ~n44684;
  assign n44686 = pi587 & ~n44648;
  assign n44687 = ~n44651 & n44686;
  assign n44688 = ~pi299 & ~n44687;
  assign n44689 = ~pi299 & ~n44685;
  assign n44690 = ~n44687 & n44689;
  assign n44691 = ~n44685 & n44688;
  assign n44692 = ~n60814 & ~n60815;
  assign n44693 = n31592 & ~n44692;
  assign n44694 = pi299 & ~n44609;
  assign n44695 = ~n60813 & ~n44673;
  assign n44696 = ~pi299 & ~n44695;
  assign n44697 = n40694 & ~n44696;
  assign n44698 = n40694 & ~n44694;
  assign n44699 = ~n44696 & n44698;
  assign n44700 = ~n44694 & n44697;
  assign n44701 = ~n44693 & ~n60816;
  assign n44702 = ~pi74 & ~n44701;
  assign n44703 = ~n44640 & n44678;
  assign n44704 = pi299 & ~n44581;
  assign n44705 = ~pi74 & n60203;
  assign n44706 = ~pi198 & ~n44564;
  assign n44707 = n44568 & ~n44706;
  assign n44708 = n31740 & ~n44707;
  assign n44709 = n44557 & ~n44708;
  assign n44710 = ~n44642 & ~n44707;
  assign n44711 = n2778 & ~n44710;
  assign n44712 = ~pi299 & ~n31739;
  assign n44713 = ~n44711 & n44712;
  assign n44714 = ~n44709 & n44713;
  assign n44715 = ~n44705 & ~n44714;
  assign n44716 = ~n44704 & n44715;
  assign n44717 = ~pi55 & ~n44716;
  assign n44718 = ~n60817 & n44717;
  assign n44719 = pi55 & n44611;
  assign n44720 = n4437 & ~n44719;
  assign n44721 = ~n44718 & n44720;
  assign n44722 = ~n4437 & n44581;
  assign n44723 = ~pi59 & ~n44722;
  assign n44724 = ~n44721 & n44723;
  assign n44725 = ~n44615 & ~n44724;
  assign n44726 = ~pi57 & ~n44725;
  assign n44727 = pi57 & ~n44581;
  assign n44728 = ~n44726 & ~n44727;
  assign n44729 = n44556 & ~n44728;
  assign n44730 = pi57 & pi332;
  assign n44731 = pi332 & ~n4437;
  assign n44732 = ~pi59 & ~n44731;
  assign n44733 = pi74 & pi332;
  assign n44734 = ~pi55 & ~n44733;
  assign n44735 = n32914 & n38298;
  assign n44736 = pi468 & ~n2778;
  assign n44737 = ~pi299 & pi587;
  assign n44738 = ~pi468 & ~n33129;
  assign n44739 = ~n44737 & n44738;
  assign n44740 = pi468 & n2778;
  assign n44741 = ~n33129 & ~n44737;
  assign n44742 = ~pi468 & ~n44741;
  assign n44743 = ~n44740 & ~n44742;
  assign n44744 = ~n44736 & ~n44739;
  assign n44745 = n44735 & ~n60818;
  assign n44746 = ~pi332 & ~n44745;
  assign n44747 = n31592 & ~n44746;
  assign n44748 = n58822 & n31783;
  assign n44749 = ~pi332 & ~n44748;
  assign n44750 = n40694 & ~n44749;
  assign n44751 = pi332 & ~n60203;
  assign n44752 = ~n44750 & ~n44751;
  assign n44753 = ~n44747 & n44752;
  assign n44754 = ~pi74 & ~n44753;
  assign n44755 = n44734 & ~n44754;
  assign n44756 = n28288 & n31736;
  assign n44757 = n60090 & n31736;
  assign n44758 = n58822 & n44756;
  assign n44759 = ~pi332 & ~n60819;
  assign n44760 = pi55 & n44759;
  assign n44761 = n4437 & ~n44760;
  assign n44762 = ~n44755 & n44761;
  assign n44763 = n44732 & ~n44762;
  assign n44764 = n4440 & ~n44759;
  assign n44765 = pi332 & ~n4440;
  assign n44766 = pi59 & ~n44765;
  assign n44767 = ~n44764 & n44766;
  assign n44768 = ~pi57 & ~n44767;
  assign n44769 = ~n44763 & n44768;
  assign n44770 = ~n44730 & ~n44769;
  assign n44771 = ~n44556 & ~n44770;
  assign n44772 = ~n44729 & ~n44771;
  assign n44773 = ~pi201 & ~n44772;
  assign n44774 = ~pi299 & n58992;
  assign n44775 = n31740 & n44641;
  assign n44776 = n44774 & ~n44775;
  assign n44777 = ~n31736 & ~n44774;
  assign n44778 = ~n44559 & ~n44774;
  assign n44779 = ~n44777 & ~n44778;
  assign n44780 = ~n44776 & ~n44777;
  assign n44781 = ~n44778 & n44780;
  assign n44782 = ~n44776 & n44779;
  assign n44783 = n44556 & n60820;
  assign n44784 = pi201 & ~n44783;
  assign po358 = ~n44773 & ~n44784;
  assign n44786 = ~pi233 & pi237;
  assign n44787 = ~n44728 & n44786;
  assign n44788 = ~n44770 & ~n44786;
  assign n44789 = ~n44787 & ~n44788;
  assign n44790 = ~pi202 & ~n44789;
  assign n44791 = n60820 & n44786;
  assign n44792 = pi202 & ~n44791;
  assign po359 = ~n44790 & ~n44792;
  assign n44794 = ~pi233 & ~pi237;
  assign n44795 = ~n44728 & n44794;
  assign n44796 = ~n44770 & ~n44794;
  assign n44797 = ~n44795 & ~n44796;
  assign n44798 = ~pi203 & ~n44797;
  assign n44799 = n60820 & n44794;
  assign n44800 = pi203 & ~n44799;
  assign po360 = ~n44798 & ~n44800;
  assign n44802 = ~pi332 & ~n2781;
  assign n44803 = ~pi907 & ~n44802;
  assign n44804 = n2781 & ~n44571;
  assign n44805 = n44803 & ~n44804;
  assign n44806 = ~n2781 & n44576;
  assign n44807 = n2781 & ~n44570;
  assign n44808 = pi907 & ~n44807;
  assign n44809 = ~n44806 & n44808;
  assign n44810 = ~n44805 & ~n44809;
  assign n44811 = pi57 & ~n44810;
  assign n44812 = ~n28288 & n44810;
  assign n44813 = ~n2781 & n44604;
  assign n44814 = n2781 & ~n44599;
  assign n44815 = pi907 & ~n44814;
  assign n44816 = ~n44813 & n44815;
  assign n44817 = pi332 & ~n6518;
  assign n44818 = pi680 & ~n44817;
  assign n44819 = ~n44600 & n44818;
  assign n44820 = n44803 & ~n44819;
  assign n44821 = ~n44816 & ~n44820;
  assign n44822 = n28288 & n44821;
  assign n44823 = ~n44812 & ~n44822;
  assign n44824 = n4440 & ~n44823;
  assign n44825 = ~n4440 & n44810;
  assign n44826 = pi59 & ~n44825;
  assign n44827 = ~n44824 & n44826;
  assign n44828 = pi299 & n44821;
  assign n44829 = n2781 & n44641;
  assign n44830 = pi332 & ~n44829;
  assign n44831 = ~pi299 & ~n44830;
  assign n44832 = n31605 & n44663;
  assign n44833 = n44831 & ~n44832;
  assign n44834 = ~n44828 & ~n44833;
  assign n44835 = n40694 & ~n44834;
  assign n44836 = n31605 & n44647;
  assign n44837 = n44831 & ~n44836;
  assign n44838 = ~n2781 & n44631;
  assign n44839 = n2781 & ~n44626;
  assign n44840 = pi907 & ~n44839;
  assign n44841 = ~n44838 & n44840;
  assign n44842 = n2781 & ~n44627;
  assign n44843 = n44803 & ~n44842;
  assign n44844 = pi299 & ~n44843;
  assign n44845 = pi299 & ~n44841;
  assign n44846 = ~n44843 & n44845;
  assign n44847 = ~n44841 & n44844;
  assign n44848 = ~n44837 & ~n60821;
  assign n44849 = n31592 & ~n44848;
  assign n44850 = ~n44835 & ~n44849;
  assign n44851 = ~pi74 & ~n44850;
  assign n44852 = pi299 & ~n44810;
  assign n44853 = ~pi468 & pi602;
  assign n44854 = pi468 & n2781;
  assign n44855 = ~n44853 & ~n44854;
  assign n44856 = n44710 & ~n44855;
  assign n44857 = ~n44830 & ~n44856;
  assign n44858 = ~pi299 & ~n44857;
  assign n44859 = ~n44705 & ~n44858;
  assign n44860 = ~n44852 & n44859;
  assign n44861 = ~pi55 & ~n44860;
  assign n44862 = ~n44851 & n44861;
  assign n44863 = pi55 & n44823;
  assign n44864 = n4437 & ~n44863;
  assign n44865 = ~n44862 & n44864;
  assign n44866 = ~n4437 & n44810;
  assign n44867 = ~pi59 & ~n44866;
  assign n44868 = ~n44865 & n44867;
  assign n44869 = ~n44827 & ~n44868;
  assign n44870 = ~pi57 & ~n44869;
  assign n44871 = ~n44811 & ~n44870;
  assign n44872 = n44556 & ~n44871;
  assign n44873 = ~pi299 & ~n44855;
  assign n44874 = ~n31654 & ~n44873;
  assign n44875 = n58822 & ~n44874;
  assign n44876 = ~pi332 & ~n44875;
  assign n44877 = n40694 & ~n44876;
  assign n44878 = pi299 & ~pi907;
  assign n44879 = ~pi299 & ~pi602;
  assign n44880 = ~pi468 & ~n44879;
  assign n44881 = ~pi468 & ~n44878;
  assign n44882 = ~n44879 & n44881;
  assign n44883 = ~n44878 & n44880;
  assign n44884 = ~n44854 & ~n60822;
  assign n44885 = n44735 & ~n44884;
  assign n44886 = ~pi332 & ~n44885;
  assign n44887 = n31592 & ~n44886;
  assign n44888 = ~n44877 & ~n44887;
  assign n44889 = ~pi74 & ~n44888;
  assign n44890 = n44734 & ~n44751;
  assign n44891 = ~n44889 & n44890;
  assign n44892 = n28288 & n31584;
  assign n44893 = n60090 & n31584;
  assign n44894 = n58822 & n44892;
  assign n44895 = ~pi332 & ~n60823;
  assign n44896 = pi55 & n44895;
  assign n44897 = n4437 & ~n44896;
  assign n44898 = ~n44891 & n44897;
  assign n44899 = n44732 & ~n44898;
  assign n44900 = n4440 & ~n44895;
  assign n44901 = n44766 & ~n44900;
  assign n44902 = ~pi57 & ~n44901;
  assign n44903 = ~n44899 & n44902;
  assign n44904 = ~n44730 & ~n44903;
  assign n44905 = ~n44556 & ~n44904;
  assign n44906 = ~n44872 & ~n44905;
  assign n44907 = ~pi204 & ~n44906;
  assign n44908 = n31605 & n44641;
  assign n44909 = n44774 & ~n44908;
  assign n44910 = ~n31584 & ~n44774;
  assign n44911 = ~n44778 & ~n44910;
  assign n44912 = ~n44909 & n44911;
  assign n44913 = n44556 & n44912;
  assign n44914 = pi204 & ~n44913;
  assign po361 = ~n44907 & ~n44914;
  assign n44916 = n44786 & ~n44871;
  assign n44917 = ~n44786 & ~n44904;
  assign n44918 = ~n44916 & ~n44917;
  assign n44919 = ~pi205 & ~n44918;
  assign n44920 = n44786 & n44912;
  assign n44921 = pi205 & ~n44920;
  assign po362 = ~n44919 & ~n44921;
  assign n44923 = pi233 & ~pi237;
  assign n44924 = ~n44871 & n44923;
  assign n44925 = ~n44904 & ~n44923;
  assign n44926 = ~n44924 & ~n44925;
  assign n44927 = ~pi206 & ~n44926;
  assign n44928 = n44912 & n44923;
  assign n44929 = pi206 & ~n44928;
  assign po363 = ~n44927 & ~n44929;
  assign n44931 = n44794 & ~n44871;
  assign n44932 = ~n44794 & ~n44904;
  assign n44933 = ~n44931 & ~n44932;
  assign n44934 = ~pi218 & ~n44933;
  assign n44935 = n44794 & n44912;
  assign n44936 = pi218 & ~n44935;
  assign po375 = ~n44934 & ~n44936;
  assign n44938 = ~n44728 & n44923;
  assign n44939 = ~n44770 & ~n44923;
  assign n44940 = ~n44938 & ~n44939;
  assign n44941 = ~pi220 & ~n44940;
  assign n44942 = n60820 & n44923;
  assign n44943 = pi220 & ~n44942;
  assign po377 = ~n44941 & ~n44943;
  assign n44945 = ~pi96 & ~pi1093;
  assign n44946 = n2727 & n44945;
  assign n44947 = n28288 & ~n44946;
  assign n44948 = ~pi96 & ~n60122;
  assign n44949 = pi479 & ~n44948;
  assign n44950 = n35649 & ~n44949;
  assign n44951 = n44947 & n44950;
  assign n44952 = n58812 & n44951;
  assign n44953 = ~n36310 & n44951;
  assign n44954 = n58812 & n44953;
  assign n44955 = ~n36310 & n44952;
  assign n44956 = n31487 & n35576;
  assign n44957 = n60280 & n35616;
  assign n44958 = n28317 & n35575;
  assign n44959 = n59291 & n60825;
  assign n44960 = pi74 & n31593;
  assign n44961 = n9189 & n60825;
  assign n44962 = ~pi54 & n44961;
  assign n44963 = pi74 & n44962;
  assign n44964 = n44959 & n44960;
  assign n44965 = ~n60824 & ~n60826;
  assign po232 = n58992 & ~n44965;
  assign n44967 = ~pi39 & pi137;
  assign n44968 = n59292 & n36455;
  assign n44969 = ~pi210 & n37864;
  assign n44970 = pi299 & n44969;
  assign n44971 = n29185 & n37864;
  assign n44972 = ~pi198 & n37879;
  assign n44973 = n44774 & n44972;
  assign n44974 = ~n60827 & ~n44973;
  assign n44975 = ~n44968 & ~n44974;
  assign n44976 = ~n58992 & n44969;
  assign n44977 = ~n44975 & ~n44976;
  assign n44978 = n31239 & ~n44977;
  assign n44979 = ~n44967 & ~n44978;
  assign n44980 = n31573 & n32934;
  assign n44981 = n31586 & n41492;
  assign n44982 = ~n38211 & ~n60828;
  assign n44983 = pi62 & ~n44982;
  assign n44984 = ~pi100 & n42169;
  assign n44985 = n58822 & ~n31676;
  assign n44986 = ~pi299 & ~n44985;
  assign n44987 = pi299 & ~n41439;
  assign n44988 = ~n44986 & ~n44987;
  assign n44989 = pi100 & n31586;
  assign n44990 = n44988 & n44989;
  assign n44991 = ~pi39 & ~n44990;
  assign n44992 = ~n44984 & n44991;
  assign n44993 = pi39 & ~n31588;
  assign n44994 = ~pi38 & ~n44993;
  assign n44995 = ~n44992 & n44994;
  assign n44996 = ~n38211 & ~n44995;
  assign n44997 = ~pi87 & ~n44996;
  assign n44998 = ~n32934 & ~n38211;
  assign n44999 = pi87 & ~n44998;
  assign n45000 = ~pi75 & ~n44999;
  assign n45001 = ~n44997 & n45000;
  assign n45002 = pi75 & ~n38211;
  assign n45003 = ~pi92 & ~n45002;
  assign n45004 = ~n45001 & n45003;
  assign n45005 = ~n60282 & ~n38211;
  assign n45006 = pi92 & ~n45005;
  assign n45007 = n6306 & ~n45006;
  assign n45008 = ~n45004 & n45007;
  assign n45009 = ~n6306 & ~n38211;
  assign n45010 = ~pi55 & ~n45009;
  assign n45011 = ~n45008 & n45010;
  assign n45012 = ~n60248 & ~n38211;
  assign n45013 = pi55 & ~n45012;
  assign n45014 = ~pi56 & ~n45013;
  assign n45015 = ~n45011 & n45014;
  assign n45016 = n28283 & n32934;
  assign n45017 = n60070 & n31586;
  assign n45018 = pi56 & ~n38211;
  assign n45019 = ~n60829 & n45018;
  assign n45020 = ~pi62 & ~n45019;
  assign n45021 = ~n45015 & n45020;
  assign n45022 = ~n44983 & ~n45021;
  assign n45023 = n4438 & ~n45022;
  assign n45024 = ~n4438 & n38211;
  assign n45025 = ~n45023 & ~n45024;
  assign n45026 = pi40 & ~pi287;
  assign n45027 = n37260 & n45026;
  assign n45028 = ~n37420 & n45027;
  assign n45029 = ~n60562 & ~n45028;
  assign n45030 = n31439 & n37181;
  assign n45031 = ~pi102 & ~n45030;
  assign n45032 = n59134 & n60165;
  assign n45033 = n6317 & n45032;
  assign n45034 = n6317 & n59134;
  assign n45035 = n60165 & n45034;
  assign n45036 = n37798 & n40275;
  assign n45037 = ~n45031 & n60830;
  assign n45038 = n6336 & n45037;
  assign n45039 = ~n45027 & ~n45038;
  assign n45040 = ~n2443 & n45039;
  assign n45041 = n2443 & ~n45038;
  assign n45042 = ~n2443 & ~n45039;
  assign n45043 = n2443 & n45038;
  assign n45044 = ~n45042 & ~n45043;
  assign n45045 = ~n45040 & ~n45041;
  assign n45046 = ~n2880 & ~n60831;
  assign n45047 = n2880 & ~n45039;
  assign n45048 = pi1091 & ~n45047;
  assign n45049 = ~n45046 & n45048;
  assign n45050 = ~pi1093 & ~n60831;
  assign n45051 = ~n2727 & n45039;
  assign n45052 = n2727 & ~n45038;
  assign n45053 = pi1093 & ~n45052;
  assign n45054 = ~n2727 & ~n45039;
  assign n45055 = n2727 & n45038;
  assign n45056 = ~n45054 & ~n45055;
  assign n45057 = pi1093 & ~n45056;
  assign n45058 = ~n45051 & n45053;
  assign n45059 = ~pi1091 & ~n60832;
  assign n45060 = ~pi1091 & ~n45050;
  assign n45061 = ~n60832 & n45060;
  assign n45062 = ~n45050 & n45059;
  assign n45063 = ~n45049 & ~n60833;
  assign n45064 = n60562 & ~n45063;
  assign po624 = ~n45029 & ~n45064;
  assign n45066 = n37086 & n60557;
  assign n45067 = n2727 & n45066;
  assign n45068 = ~pi1093 & ~n45067;
  assign n45069 = pi1093 & ~n40281;
  assign n45070 = ~n6416 & n28288;
  assign n45071 = ~n45069 & n45070;
  assign n45072 = ~n45068 & n45071;
  assign n45073 = n3213 & ~n45072;
  assign n45074 = ~pi1093 & n2597;
  assign n45075 = ~pi1093 & n60280;
  assign n45076 = n32908 & n45074;
  assign n45077 = ~pi1093 & n2599;
  assign n45078 = n28288 & n45077;
  assign n45079 = n59292 & n60834;
  assign n45080 = n37101 & n60835;
  assign n45081 = n36278 & n45080;
  assign n45082 = n36281 & n45080;
  assign n45083 = n6389 & n45081;
  assign n45084 = ~n3213 & ~n60836;
  assign n45085 = n58992 & ~n45084;
  assign po246 = ~n45073 & n45085;
  assign n45087 = pi1092 & ~n2797;
  assign n45088 = ~pi340 & n44497;
  assign n45089 = n58992 & n45088;
  assign n45090 = ~pi340 & po637;
  assign n45091 = ~pi330 & ~po637;
  assign n45092 = ~n60837 & ~n45091;
  assign n45093 = ~n58992 & n45087;
  assign n45094 = ~pi330 & n45093;
  assign n45095 = pi330 & ~n44497;
  assign n45096 = n58992 & n45087;
  assign n45097 = pi340 & n44497;
  assign n45098 = n45096 & ~n45097;
  assign n45099 = ~pi330 & ~n44497;
  assign n45100 = ~n45088 & ~n45099;
  assign n45101 = n45096 & ~n45100;
  assign n45102 = ~n45095 & n45098;
  assign n45103 = ~n45094 & ~n60838;
  assign n45104 = n45087 & ~n45092;
  assign n45105 = ~pi341 & n44497;
  assign n45106 = n58992 & n45105;
  assign n45107 = ~pi341 & po637;
  assign n45108 = ~pi331 & ~po637;
  assign n45109 = ~n60840 & ~n45108;
  assign n45110 = ~pi331 & n45093;
  assign n45111 = pi331 & ~n44497;
  assign n45112 = pi341 & n44497;
  assign n45113 = n45096 & ~n45112;
  assign n45114 = ~pi331 & ~n44497;
  assign n45115 = ~n45105 & ~n45114;
  assign n45116 = n45096 & ~n45115;
  assign n45117 = ~n45111 & n45113;
  assign n45118 = ~n45110 & ~n60841;
  assign n45119 = n45087 & ~n45109;
  assign n45120 = ~pi340 & ~po637;
  assign n45121 = ~pi331 & n44497;
  assign n45122 = n58992 & n45121;
  assign n45123 = ~pi331 & po637;
  assign n45124 = n45096 & ~n45121;
  assign n45125 = ~n45093 & ~n45124;
  assign n45126 = n45087 & ~n60843;
  assign n45127 = pi340 & n45093;
  assign n45128 = ~pi340 & ~n44497;
  assign n45129 = n45096 & ~n45128;
  assign n45130 = ~n45121 & n45129;
  assign n45131 = ~n45127 & ~n45130;
  assign n45132 = pi340 & ~n60844;
  assign n45133 = n44497 & n45124;
  assign n45134 = ~n45132 & ~n45133;
  assign n45135 = ~n45120 & ~n60844;
  assign n45136 = ~pi330 & po637;
  assign n45137 = ~pi341 & ~po637;
  assign n45138 = ~n45136 & ~n45137;
  assign po498 = n45087 & ~n45138;
  assign n45140 = n35617 & n36552;
  assign n45141 = n35650 & n38480;
  assign n45142 = pi96 & n2620;
  assign n45143 = n2444 & n45142;
  assign n45144 = ~n35650 & n45143;
  assign n45145 = n38284 & n45144;
  assign n45146 = ~n45141 & ~n45145;
  assign n45147 = ~pi95 & ~n45146;
  assign n45148 = ~n45140 & ~n45147;
  assign po254 = n60562 & ~n45148;
  assign n45150 = n43298 & n44988;
  assign n45151 = ~n43297 & ~n45150;
  assign n45152 = ~pi38 & ~n45151;
  assign n45153 = ~pi87 & ~n45152;
  assign n45154 = n31561 & ~n45153;
  assign n45155 = ~pi92 & ~n45154;
  assign n45156 = ~pi74 & n35283;
  assign n45157 = ~n45155 & n45156;
  assign n45158 = ~pi55 & ~n45157;
  assign n45159 = ~n28594 & ~n45158;
  assign n45160 = ~pi56 & ~n45159;
  assign n45161 = ~n31570 & ~n45160;
  assign n45162 = ~pi62 & ~n45161;
  assign n45163 = ~pi57 & n31576;
  assign po275 = ~n45162 & n45163;
  assign n45165 = ~pi58 & n2732;
  assign n45166 = n2530 & n37093;
  assign n45167 = ~n45165 & ~n45166;
  assign n45168 = n60165 & ~n45167;
  assign n45169 = n2880 & ~n45168;
  assign n45170 = ~n2441 & n45168;
  assign n45171 = n6547 & n45066;
  assign n45172 = pi829 & ~n45171;
  assign n45173 = ~n45170 & n45172;
  assign n45174 = ~n2692 & n45173;
  assign n45175 = ~n45169 & ~n45174;
  assign n45176 = pi1091 & ~n45175;
  assign n45177 = ~n2727 & n45168;
  assign n45178 = ~pi829 & ~n45177;
  assign n45179 = ~n45173 & ~n45178;
  assign n45180 = ~pi1093 & ~n45179;
  assign n45181 = ~n37057 & ~n45165;
  assign n45182 = n40279 & ~n45181;
  assign n45183 = ~n2878 & ~n28504;
  assign n45184 = ~n45182 & ~n45183;
  assign n45185 = ~n45177 & n45184;
  assign n45186 = n60562 & ~n45185;
  assign n45187 = ~n45180 & n45186;
  assign po205 = ~n45176 & n45187;
  assign n45189 = pi1093 & n35646;
  assign n45190 = ~pi96 & ~n45189;
  assign n45191 = n2672 & ~n31503;
  assign n45192 = n58837 & n45191;
  assign n45193 = pi96 & ~pi1093;
  assign n45194 = n2798 & ~n36310;
  assign n45195 = ~n45193 & ~n45194;
  assign n45196 = n2672 & ~n45195;
  assign n45197 = n58837 & n45196;
  assign n45198 = ~n45190 & n45192;
  assign n45199 = ~pi75 & ~n60846;
  assign n45200 = pi75 & ~n44959;
  assign n45201 = n37304 & ~n45200;
  assign po233 = ~n45199 & n45201;
  assign n45203 = pi315 & ~n60837;
  assign n45204 = pi1080 & n60837;
  assign n45205 = ~n45203 & ~n45204;
  assign n45206 = pi316 & ~n60837;
  assign n45207 = pi1047 & n60837;
  assign n45208 = ~n45206 & ~n45207;
  assign n45209 = pi317 & ~n45136;
  assign n45210 = pi1078 & n45136;
  assign n45211 = ~n45209 & ~n45210;
  assign n45212 = pi318 & ~n60840;
  assign n45213 = pi1074 & n60840;
  assign n45214 = ~n45212 & ~n45213;
  assign n45215 = pi319 & ~n60840;
  assign n45216 = pi1072 & n60840;
  assign n45217 = ~n45215 & ~n45216;
  assign n45218 = pi320 & ~n60837;
  assign n45219 = pi1048 & n60837;
  assign n45220 = ~n45218 & ~n45219;
  assign n45221 = pi321 & ~n60837;
  assign n45222 = pi1058 & n60837;
  assign n45223 = ~n45221 & ~n45222;
  assign n45224 = pi322 & ~n60837;
  assign n45225 = pi1051 & n60837;
  assign n45226 = ~n45224 & ~n45225;
  assign n45227 = pi323 & ~n60837;
  assign n45228 = pi1065 & n60837;
  assign n45229 = ~n45227 & ~n45228;
  assign n45230 = pi324 & ~n60840;
  assign n45231 = pi1086 & n60840;
  assign n45232 = ~n45230 & ~n45231;
  assign n45233 = pi325 & ~n60840;
  assign n45234 = pi1063 & n60840;
  assign n45235 = ~n45233 & ~n45234;
  assign n45236 = pi326 & ~n60840;
  assign n45237 = pi1057 & n60840;
  assign n45238 = ~n45236 & ~n45237;
  assign n45239 = pi327 & ~n60837;
  assign n45240 = pi1040 & n60837;
  assign n45241 = ~n45239 & ~n45240;
  assign n45242 = pi328 & ~n60840;
  assign n45243 = pi1058 & n60840;
  assign n45244 = ~n45242 & ~n45243;
  assign n45245 = pi329 & ~n60840;
  assign n45246 = pi1043 & n60840;
  assign n45247 = ~n45245 & ~n45246;
  assign n45248 = pi333 & ~n60840;
  assign n45249 = pi1040 & n60840;
  assign n45250 = ~n45248 & ~n45249;
  assign n45251 = pi334 & ~n60840;
  assign n45252 = pi1065 & n60840;
  assign n45253 = ~n45251 & ~n45252;
  assign n45254 = pi335 & ~n60840;
  assign n45255 = pi1069 & n60840;
  assign n45256 = ~n45254 & ~n45255;
  assign n45257 = pi338 & ~n45136;
  assign n45258 = pi1072 & n45136;
  assign n45259 = ~n45257 & ~n45258;
  assign n45260 = pi339 & ~n45136;
  assign n45261 = pi1086 & n45136;
  assign n45262 = ~n45260 & ~n45261;
  assign n45263 = pi344 & ~n60837;
  assign n45264 = pi1069 & n60837;
  assign n45265 = ~n45263 & ~n45264;
  assign n45266 = pi349 & ~n60837;
  assign n45267 = pi1043 & n60837;
  assign n45268 = ~n45266 & ~n45267;
  assign n45269 = pi352 & ~n60837;
  assign n45270 = pi1078 & n60837;
  assign n45271 = ~n45269 & ~n45270;
  assign n45272 = pi353 & ~n60837;
  assign n45273 = pi1063 & n60837;
  assign n45274 = ~n45272 & ~n45273;
  assign n45275 = pi365 & ~n45136;
  assign n45276 = pi1065 & n45136;
  assign n45277 = ~n45275 & ~n45276;
  assign n45278 = pi366 & ~n45136;
  assign n45279 = pi1069 & n45136;
  assign n45280 = ~n45278 & ~n45279;
  assign n45281 = pi369 & ~n45136;
  assign n45282 = pi1080 & n45136;
  assign n45283 = ~n45281 & ~n45282;
  assign n45284 = pi371 & ~n45136;
  assign n45285 = pi1051 & n45136;
  assign n45286 = ~n45284 & ~n45285;
  assign n45287 = pi372 & ~n45136;
  assign n45288 = pi1048 & n45136;
  assign n45289 = ~n45287 & ~n45288;
  assign n45290 = pi375 & ~n45136;
  assign n45291 = pi1047 & n45136;
  assign n45292 = ~n45290 & ~n45291;
  assign n45293 = pi377 & ~n45136;
  assign n45294 = pi1074 & n45136;
  assign n45295 = ~n45293 & ~n45294;
  assign n45296 = pi378 & ~n45136;
  assign n45297 = pi1063 & n45136;
  assign n45298 = ~n45296 & ~n45297;
  assign n45299 = pi394 & ~n60840;
  assign n45300 = pi1080 & n60840;
  assign n45301 = ~n45299 & ~n45300;
  assign n45302 = pi396 & ~n60840;
  assign n45303 = pi1051 & n60840;
  assign n45304 = ~n45302 & ~n45303;
  assign n45305 = pi397 & ~n60840;
  assign n45306 = pi1048 & n60840;
  assign n45307 = ~n45305 & ~n45306;
  assign n45308 = pi399 & ~n60840;
  assign n45309 = pi1047 & n60840;
  assign n45310 = ~n45308 & ~n45309;
  assign n45311 = pi402 & ~n60840;
  assign n45312 = pi1078 & n60840;
  assign n45313 = ~n45311 & ~n45312;
  assign n45314 = pi416 & ~n60843;
  assign n45315 = pi1069 & n60843;
  assign n45316 = ~n45314 & ~n45315;
  assign n45317 = pi419 & ~n60843;
  assign n45318 = pi1080 & n60843;
  assign n45319 = ~n45317 & ~n45318;
  assign n45320 = pi421 & ~n60843;
  assign n45321 = pi1051 & n60843;
  assign n45322 = ~n45320 & ~n45321;
  assign n45323 = pi422 & ~n60843;
  assign n45324 = pi1048 & n60843;
  assign n45325 = ~n45323 & ~n45324;
  assign n45326 = pi424 & ~n60843;
  assign n45327 = pi1047 & n60843;
  assign n45328 = ~n45326 & ~n45327;
  assign n45329 = pi427 & ~n60843;
  assign n45330 = pi1078 & n60843;
  assign n45331 = ~n45329 & ~n45330;
  assign n45332 = pi439 & ~n45136;
  assign n45333 = pi1057 & n45136;
  assign n45334 = ~n45332 & ~n45333;
  assign n45335 = pi440 & ~n45136;
  assign n45336 = pi1043 & n45136;
  assign n45337 = ~n45335 & ~n45336;
  assign n45338 = pi442 & ~n45136;
  assign n45339 = pi1058 & n45136;
  assign n45340 = ~n45338 & ~n45339;
  assign n45341 = pi444 & ~n60843;
  assign n45342 = pi1072 & n60843;
  assign n45343 = ~n45341 & ~n45342;
  assign n45344 = pi446 & ~n60843;
  assign n45345 = pi1086 & n60843;
  assign n45346 = ~n45344 & ~n45345;
  assign n45347 = pi447 & ~n45136;
  assign n45348 = pi1040 & n45136;
  assign n45349 = ~n45347 & ~n45348;
  assign n45350 = pi448 & ~n60843;
  assign n45351 = pi1074 & n60843;
  assign n45352 = ~n45350 & ~n45351;
  assign n45353 = pi449 & ~n60843;
  assign n45354 = pi1057 & n60843;
  assign n45355 = ~n45353 & ~n45354;
  assign n45356 = pi451 & ~n60843;
  assign n45357 = pi1063 & n60843;
  assign n45358 = ~n45356 & ~n45357;
  assign n45359 = pi453 & ~n60843;
  assign n45360 = pi1040 & n60843;
  assign n45361 = ~n45359 & ~n45360;
  assign n45362 = pi454 & ~n60843;
  assign n45363 = pi1043 & n60843;
  assign n45364 = ~n45362 & ~n45363;
  assign n45365 = pi458 & ~n60837;
  assign n45366 = pi1072 & n60837;
  assign n45367 = ~n45365 & ~n45366;
  assign n45368 = pi459 & ~n60843;
  assign n45369 = pi1058 & n60843;
  assign n45370 = ~n45368 & ~n45369;
  assign n45371 = pi460 & ~n60837;
  assign n45372 = pi1086 & n60837;
  assign n45373 = ~n45371 & ~n45372;
  assign n45374 = pi461 & ~n60837;
  assign n45375 = pi1057 & n60837;
  assign n45376 = ~n45374 & ~n45375;
  assign n45377 = pi462 & ~n60837;
  assign n45378 = pi1074 & n60837;
  assign n45379 = ~n45377 & ~n45378;
  assign n45380 = pi464 & ~n60843;
  assign n45381 = pi1065 & n60843;
  assign n45382 = ~n45380 & ~n45381;
  assign n45383 = ~pi97 & n58805;
  assign n45384 = ~pi108 & ~n45383;
  assign n45385 = n2531 & ~n45384;
  assign n45386 = n60477 & n45385;
  assign n45387 = ~pi314 & ~n45386;
  assign n45388 = pi314 & ~n2583;
  assign n45389 = n2581 & ~n36247;
  assign n45390 = ~n45388 & n45389;
  assign n45391 = ~n45387 & n45390;
  assign n45392 = n2581 & n36247;
  assign n45393 = n45386 & n45392;
  assign n45394 = ~pi51 & ~n45393;
  assign n45395 = ~n45391 & n45394;
  assign n45396 = n58810 & n58815;
  assign n45397 = ~n45395 & n45396;
  assign n45398 = ~pi87 & ~n45397;
  assign n45399 = n31561 & n37304;
  assign po266 = ~n45398 & n45399;
  assign n45401 = pi39 & ~pi979;
  assign n45402 = ~n2802 & n45401;
  assign n45403 = n2803 & n45402;
  assign n45404 = n2801 & n45403;
  assign n45405 = n32632 & n45404;
  assign n45406 = n24385 & n59928;
  assign n45407 = n58826 & n45406;
  assign n45408 = pi468 & ~n45407;
  assign n45409 = ~n45405 & ~n45408;
  assign n45410 = n2516 & n59134;
  assign n45411 = pi24 & n60165;
  assign n45412 = ~pi39 & n45411;
  assign n45413 = n45410 & n45412;
  assign n45414 = n28334 & n45413;
  assign n45415 = ~n45404 & ~n45414;
  assign po218 = n32632 & ~n45415;
  assign n45417 = po740 & n60696;
  assign po194 = ~n45181 & n45417;
  assign n45419 = n2461 & n28371;
  assign n45420 = n37080 & n45419;
  assign n45421 = ~pi64 & n6325;
  assign n45422 = n45420 & n45421;
  assign n45423 = ~pi81 & ~n45422;
  assign n45424 = ~pi199 & pi200;
  assign n45425 = ~pi299 & n45424;
  assign n45426 = pi211 & ~pi219;
  assign n45427 = pi299 & n45426;
  assign n45428 = ~n45425 & ~n45427;
  assign n45429 = pi314 & ~n45428;
  assign n45430 = n60165 & n45429;
  assign n45431 = ~n45423 & n45430;
  assign n45432 = n60263 & n45431;
  assign n45433 = pi314 & n58783;
  assign n45434 = n60557 & n45433;
  assign n45435 = n60521 & n45428;
  assign n45436 = n45434 & n45435;
  assign n45437 = n45420 & n45436;
  assign n45438 = ~n45432 & ~n45437;
  assign po229 = n60562 & ~n45438;
  assign n45440 = pi81 & ~pi102;
  assign n45441 = n45434 & n45440;
  assign n45442 = n2520 & n45441;
  assign n45443 = n28288 & n45442;
  assign n45444 = ~pi299 & n36719;
  assign n45445 = ~pi211 & pi299;
  assign n45446 = ~pi219 & n45445;
  assign n45447 = pi211 & pi299;
  assign n45448 = pi219 & pi299;
  assign n45449 = ~n45447 & ~n45448;
  assign n45450 = ~n36720 & n45449;
  assign n45451 = ~n45444 & ~n45446;
  assign n45452 = n58992 & n60847;
  assign po242 = n45443 & n45452;
  assign n45454 = ~n36413 & ~n40733;
  assign n45455 = ~pi314 & n40733;
  assign n45456 = po740 & ~n45455;
  assign n45457 = n60696 & ~n45456;
  assign n45458 = ~n45454 & n45457;
  assign n45459 = pi53 & n2501;
  assign n45460 = pi53 & n60623;
  assign n45461 = n58798 & n45459;
  assign n45462 = n60075 & n60848;
  assign n45463 = n45411 & n45462;
  assign n45464 = ~pi39 & ~n45463;
  assign n45465 = ~pi287 & ~pi979;
  assign n45466 = n2802 & n45465;
  assign n45467 = pi39 & ~n45466;
  assign n45468 = n32632 & ~n45467;
  assign n45469 = ~n45464 & n45468;
  assign n45470 = ~n37419 & n45468;
  assign n45471 = ~n45464 & n45470;
  assign n45472 = ~n37419 & n45469;
  assign n45473 = ~n38255 & ~n38440;
  assign n45474 = ~pi70 & ~n45473;
  assign n45475 = ~pi51 & ~n45474;
  assign n45476 = n2604 & ~n45475;
  assign n45477 = n31408 & ~n45476;
  assign n45478 = n31402 & ~n45477;
  assign n45479 = n31401 & ~n45478;
  assign n45480 = ~n31498 & ~n45479;
  assign n45481 = ~pi95 & ~n45480;
  assign n45482 = n38365 & ~n45481;
  assign n45483 = ~pi39 & ~n45482;
  assign n45484 = ~pi38 & ~n37419;
  assign n45485 = ~n45483 & n45484;
  assign n45486 = ~pi100 & n45485;
  assign n45487 = n37429 & ~n45486;
  assign n45488 = ~n31560 & ~n45487;
  assign n45489 = ~pi75 & ~n45488;
  assign n45490 = ~n28303 & ~n45489;
  assign n45491 = ~pi92 & ~n45490;
  assign n45492 = n35283 & ~n45491;
  assign n45493 = ~pi74 & ~n45492;
  assign n45494 = n31398 & ~n45493;
  assign n45495 = ~pi56 & ~n45494;
  assign n45496 = ~n31570 & ~n45495;
  assign n45497 = ~pi62 & ~n45496;
  assign po393 = n45163 & ~n45497;
  assign n45499 = ~n58992 & n45426;
  assign n45500 = pi71 & n45499;
  assign n45501 = pi71 & ~n45428;
  assign n45502 = pi84 & n29129;
  assign n45503 = n38966 & n45502;
  assign n45504 = n2447 & n45503;
  assign n45505 = n58790 & n40720;
  assign n45506 = n2532 & n45505;
  assign n45507 = n58797 & n40720;
  assign n45508 = n45428 & n60850;
  assign n45509 = n60278 & ~n45428;
  assign n45510 = n60262 & n45509;
  assign n45511 = ~n45508 & ~n45510;
  assign n45512 = n28288 & n60165;
  assign n45513 = ~n45511 & n45512;
  assign n45514 = n45504 & n45513;
  assign n45515 = ~n45501 & ~n45514;
  assign n45516 = n58992 & ~n45515;
  assign n45517 = ~n45500 & ~n45516;
  assign n45518 = ~pi199 & ~pi299;
  assign n45519 = n45443 & ~n45518;
  assign n45520 = pi219 & ~n45519;
  assign n45521 = pi199 & ~pi299;
  assign n45522 = n2671 & n45521;
  assign n45523 = n40929 & n45522;
  assign n45524 = n45442 & n45523;
  assign n45525 = ~pi219 & ~n45524;
  assign n45526 = n58992 & ~n45525;
  assign po224 = ~n45520 & n45526;
  assign n45528 = pi54 & n58822;
  assign n45529 = ~pi49 & ~pi76;
  assign n45530 = n6323 & n45529;
  assign n45531 = ~pi60 & ~pi85;
  assign n45532 = pi106 & n45531;
  assign n45533 = n2457 & n36224;
  assign n45534 = n45532 & n45533;
  assign n45535 = n45530 & n45534;
  assign n45536 = n6322 & n37189;
  assign n45537 = n40563 & n45536;
  assign n45538 = n45535 & n45536;
  assign n45539 = n40563 & n45538;
  assign n45540 = n45535 & n45537;
  assign n45541 = ~pi53 & ~n60851;
  assign n45542 = n29725 & ~n45541;
  assign n45543 = ~pi54 & n37798;
  assign n45544 = n45542 & n45543;
  assign n45545 = ~n45528 & ~n45544;
  assign n45546 = n9189 & n60412;
  assign n45547 = ~n45545 & n45546;
  assign n45548 = ~pi39 & ~n45547;
  assign po456 = ~n45467 & ~n45548;
  assign n45550 = pi38 & ~n60825;
  assign n45551 = pi332 & n35633;
  assign n45552 = ~pi64 & ~n45551;
  assign n45553 = ~pi39 & ~pi81;
  assign n45554 = ~pi841 & n45553;
  assign n45555 = n2482 & n45554;
  assign n45556 = n60557 & n45555;
  assign n45557 = ~n45552 & n45556;
  assign n45558 = ~pi81 & ~n31415;
  assign n45559 = ~pi39 & ~pi841;
  assign n45560 = n2482 & n45559;
  assign n45561 = n60557 & n45560;
  assign n45562 = ~n45552 & n45560;
  assign n45563 = n60557 & n45562;
  assign n45564 = ~n45552 & n45561;
  assign n45565 = n45558 & n60852;
  assign n45566 = ~n31415 & n45557;
  assign n45567 = ~pi38 & ~n60853;
  assign n45568 = n59928 & ~n45567;
  assign po196 = ~n45550 & n45568;
  assign n45570 = pi979 & n37049;
  assign po203 = n2801 & n45570;
  assign n45572 = n35619 & n40565;
  assign n45573 = n45530 & n45572;
  assign n45574 = pi61 & ~pi82;
  assign n45575 = ~pi83 & ~pi89;
  assign n45576 = n45574 & n45575;
  assign n45577 = n2471 & n37186;
  assign n45578 = n45576 & n45577;
  assign n45579 = n37185 & n45578;
  assign n45580 = n36230 & n45579;
  assign n45581 = n45573 & n45580;
  assign n45582 = n58797 & n45581;
  assign n45583 = ~pi841 & n45582;
  assign n45584 = n2532 & n60074;
  assign n45585 = pi24 & n45584;
  assign n45586 = ~n45583 & ~n45585;
  assign po204 = n60696 & ~n45586;
  assign n45588 = pi74 & ~n58826;
  assign n45589 = pi841 & n2641;
  assign n45590 = n2579 & n45589;
  assign n45591 = ~pi70 & pi841;
  assign n45592 = ~pi72 & pi841;
  assign n45593 = n2641 & n45592;
  assign n45594 = n2600 & n45591;
  assign n45595 = n30008 & n60854;
  assign n45596 = n2579 & n60854;
  assign n45597 = n2621 & n45596;
  assign n45598 = n2599 & n45590;
  assign n45599 = n60688 & n60855;
  assign n45600 = ~pi74 & ~n45599;
  assign n45601 = n37907 & ~n45600;
  assign po207 = ~n45588 & n45601;
  assign n45603 = pi54 & ~n44961;
  assign n45604 = n45410 & n60851;
  assign n45605 = n6343 & n60203;
  assign n45606 = n40577 & n45605;
  assign n45607 = n45604 & n45606;
  assign n45608 = ~pi54 & ~n45607;
  assign n45609 = n60412 & ~n45608;
  assign po212 = ~n45603 & n45609;
  assign n45611 = pi55 & n37250;
  assign n45612 = ~n40706 & ~n45611;
  assign n45613 = n2598 & n60070;
  assign n45614 = n31495 & n45613;
  assign n45615 = pi56 & ~n45614;
  assign n45616 = n4438 & ~n45615;
  assign po214 = ~n45612 & n45616;
  assign n45618 = pi841 & n45582;
  assign n45619 = ~pi24 & n45410;
  assign n45620 = n2516 & n60615;
  assign n45621 = n28334 & n60856;
  assign n45622 = ~n45618 & ~n45621;
  assign po219 = n60696 & ~n45622;
  assign n45624 = pi57 & ~n37251;
  assign n45625 = n40707 & n45614;
  assign n45626 = ~pi57 & ~n45625;
  assign n45627 = ~pi59 & ~n45626;
  assign n45628 = ~pi59 & ~n45624;
  assign n45629 = ~n45626 & n45628;
  assign n45630 = ~n45624 & n45627;
  assign n45631 = pi841 & n2581;
  assign n45632 = n35634 & n45631;
  assign n45633 = ~pi24 & pi70;
  assign n45634 = n2593 & n45633;
  assign n45635 = ~n45632 & ~n45634;
  assign n45636 = n58821 & n60562;
  assign n45637 = pi70 & ~n2687;
  assign n45638 = pi841 & n2580;
  assign n45639 = n35634 & n45638;
  assign n45640 = ~pi70 & ~n45639;
  assign n45641 = n45636 & ~n45640;
  assign n45642 = ~n45637 & n45641;
  assign n45643 = ~n45635 & n45636;
  assign n45644 = ~pi1050 & n29751;
  assign n45645 = ~pi90 & ~n45644;
  assign n45646 = ~pi93 & n32914;
  assign n45647 = n2444 & n45636;
  assign n45648 = n32914 & n60562;
  assign n45649 = ~pi93 & n60859;
  assign n45650 = n60562 & n45646;
  assign n45651 = ~n45645 & n60860;
  assign n45652 = ~n45645 & n60859;
  assign n45653 = n32527 & n45652;
  assign n45654 = ~n28325 & n45651;
  assign po248 = ~n2555 & n60861;
  assign n45656 = ~pi1050 & n58822;
  assign n45657 = pi92 & ~n45656;
  assign n45658 = pi93 & n32914;
  assign n45659 = n28322 & n45658;
  assign n45660 = ~pi92 & ~n45659;
  assign n45661 = n37905 & ~n45660;
  assign po251 = ~n45657 & n45661;
  assign n45663 = ~pi92 & n60166;
  assign n45664 = ~n36301 & ~n45663;
  assign n45665 = pi314 & pi1050;
  assign n45666 = n37905 & n45665;
  assign po256 = ~n45664 & n45666;
  assign n45668 = pi24 & n45604;
  assign n45669 = n38979 & n45542;
  assign n45670 = ~n45668 & ~n45669;
  assign n45671 = pi841 & ~n45670;
  assign n45672 = n37331 & n45462;
  assign n45673 = ~n45671 & ~n45672;
  assign po264 = n60696 & ~n45673;
  assign n45675 = pi72 & n36552;
  assign n45676 = n59138 & n45455;
  assign n45677 = ~n45675 & ~n45676;
  assign po269 = n40717 & ~n45677;
  assign n45679 = n35636 & n45584;
  assign n45680 = ~n35634 & ~n45584;
  assign n45681 = n2580 & ~n45680;
  assign n45682 = ~pi70 & ~n45681;
  assign n45683 = pi332 & n29717;
  assign n45684 = ~n45682 & n45683;
  assign n45685 = ~n45679 & ~n45684;
  assign n45686 = ~pi39 & ~n45685;
  assign n45687 = pi39 & n36455;
  assign n45688 = ~pi38 & ~n45687;
  assign n45689 = ~n45686 & n45688;
  assign po489 = n36085 & ~n45689;
  assign n45691 = ~pi93 & pi102;
  assign n45692 = pi102 & n2589;
  assign n45693 = n2445 & n45691;
  assign n45694 = pi102 & n58783;
  assign n45695 = n2589 & n45694;
  assign n45696 = n58783 & n60862;
  assign n45697 = n58823 & n60863;
  assign n45698 = n58792 & n45697;
  assign n45699 = n2521 & n45698;
  assign n45700 = ~pi40 & ~n45699;
  assign n45701 = n6316 & ~n45700;
  assign n45702 = ~pi1082 & ~n45701;
  assign n45703 = n2621 & n45699;
  assign n45704 = pi1082 & ~n45703;
  assign n45705 = n60562 & ~n45704;
  assign po198 = ~n45702 & n45705;
  assign n45707 = pi841 & n60562;
  assign n45708 = n36237 & n45707;
  assign n45709 = ~pi51 & n60854;
  assign n45710 = n36237 & n45709;
  assign n45711 = n60562 & n45710;
  assign n45712 = n37815 & n45711;
  assign n45713 = n60557 & n45708;
  assign n45714 = n6306 & n44961;
  assign n45715 = ~pi74 & n44962;
  assign n45716 = n59292 & n60825;
  assign n45717 = pi55 & ~n60865;
  assign n45718 = n2482 & n28288;
  assign n45719 = n60557 & n45718;
  assign n45720 = n6333 & n45719;
  assign n45721 = ~pi55 & ~n45720;
  assign n45722 = n4439 & ~n45721;
  assign n45723 = pi55 & n60865;
  assign n45724 = n2482 & n60557;
  assign n45725 = n6333 & n60070;
  assign n45726 = n45724 & n45725;
  assign n45727 = ~n45723 & ~n45726;
  assign n45728 = n4439 & ~n45727;
  assign n45729 = ~n45717 & n45722;
  assign po216 = n2555 & n60860;
  assign n45731 = n2530 & n60696;
  assign n45732 = n58796 & n45731;
  assign n45733 = n58797 & n60696;
  assign n45734 = ~pi107 & pi841;
  assign n45735 = pi64 & ~n45734;
  assign n45736 = ~pi64 & ~pi107;
  assign n45737 = ~pi63 & ~pi81;
  assign n45738 = ~n45736 & n45737;
  assign n45739 = ~n45735 & n45738;
  assign n45740 = n2482 & n45739;
  assign n45741 = n60867 & n45740;
  assign n45742 = ~pi63 & pi107;
  assign n45743 = n2486 & n45742;
  assign n45744 = ~pi64 & ~n45743;
  assign n45745 = n2482 & ~n45744;
  assign n45746 = n45558 & n45745;
  assign n45747 = pi841 & ~n45746;
  assign n45748 = n58786 & n45742;
  assign n45749 = ~pi841 & ~n45748;
  assign n45750 = n60867 & ~n45749;
  assign n45751 = ~n45747 & n45750;
  assign n45752 = n2486 & n45741;
  assign n45753 = pi83 & ~pi103;
  assign n45754 = n40720 & n45753;
  assign n45755 = n60562 & n45754;
  assign n45756 = n45434 & n45755;
  assign n45757 = n58782 & n45755;
  assign n45758 = n45434 & n45757;
  assign n45759 = n58782 & n45756;
  assign n45760 = pi69 & n6321;
  assign n45761 = n32871 & n45760;
  assign n45762 = ~pi71 & ~n45761;
  assign n45763 = ~pi81 & ~pi314;
  assign n45764 = n2482 & n45763;
  assign n45765 = n28390 & n45764;
  assign n45766 = ~n45762 & n45765;
  assign n45767 = pi71 & pi314;
  assign n45768 = n2471 & n45767;
  assign n45769 = n60278 & n45768;
  assign n45770 = n2469 & n45769;
  assign n45771 = ~n45766 & ~n45770;
  assign po227 = n60867 & ~n45771;
  assign n45773 = ~pi314 & ~n39013;
  assign n45774 = pi314 & ~n39011;
  assign n45775 = n60696 & ~n45774;
  assign po235 = ~n45773 & n45775;
  assign n45777 = n58992 & n45719;
  assign n45778 = n60562 & n45724;
  assign n45779 = pi81 & ~pi314;
  assign n45780 = n2520 & n45779;
  assign n45781 = pi68 & ~pi81;
  assign n45782 = n2458 & n45781;
  assign n45783 = n37080 & n45782;
  assign n45784 = n45421 & n45783;
  assign n45785 = n28345 & n45784;
  assign n45786 = ~n45780 & ~n45785;
  assign po239 = n60870 & ~n45786;
  assign n45788 = pi69 & pi314;
  assign n45789 = n2466 & n45788;
  assign n45790 = pi66 & ~pi73;
  assign n45791 = n2465 & n45790;
  assign n45792 = n2459 & n45791;
  assign n45793 = n2462 & n45791;
  assign n45794 = n2455 & n45792;
  assign n45795 = ~n45789 & ~n60871;
  assign n45796 = n40721 & n60867;
  assign po240 = ~n45795 & n45796;
  assign n45798 = ~pi83 & ~n45503;
  assign n45799 = n28342 & n60850;
  assign n45800 = n60850 & ~n45798;
  assign n45801 = n28342 & n45800;
  assign n45802 = ~n45798 & n45799;
  assign n45803 = ~pi314 & ~n60872;
  assign n45804 = n45504 & n60850;
  assign n45805 = pi314 & ~n45804;
  assign n45806 = n60696 & ~n45805;
  assign po241 = ~n45803 & n45806;
  assign n45808 = n28382 & n40722;
  assign n45809 = ~pi314 & n40723;
  assign n45810 = n45419 & n45809;
  assign n45811 = ~n45808 & ~n45810;
  assign po243 = n60867 & ~n45811;
  assign n45813 = n60077 & n40720;
  assign n45814 = pi314 & n60696;
  assign n45815 = n58797 & n45814;
  assign n45816 = pi314 & n60867;
  assign n45817 = n58790 & n45813;
  assign n45818 = n60077 & n45505;
  assign n45819 = n2532 & n45814;
  assign n45820 = n60874 & n45819;
  assign n45821 = n45813 & n60873;
  assign n45822 = pi109 & n58794;
  assign n45823 = ~pi109 & ~pi314;
  assign n45824 = n45813 & n45823;
  assign n45825 = ~n45822 & ~n45824;
  assign n45826 = n60696 & n40727;
  assign n45827 = ~pi109 & ~n60874;
  assign n45828 = n28448 & ~n45827;
  assign n45829 = ~pi314 & ~n45828;
  assign n45830 = pi109 & n2540;
  assign n45831 = n2548 & n45830;
  assign n45832 = pi314 & ~n45831;
  assign n45833 = n45731 & ~n45832;
  assign n45834 = ~n45829 & n45833;
  assign n45835 = ~n45825 & n45826;
  assign n45836 = n39101 & n60696;
  assign n45837 = n60624 & n45814;
  assign n45838 = n58815 & n60555;
  assign n45839 = ~n28549 & ~n45838;
  assign n45840 = ~pi75 & ~n45839;
  assign n45841 = n28575 & n37225;
  assign n45842 = ~n45840 & ~n45841;
  assign n45843 = ~pi87 & ~pi250;
  assign n45844 = n37304 & n45843;
  assign po407 = ~n45842 & n45844;
  assign n45846 = n40723 & n60867;
  assign n45847 = n60076 & n40723;
  assign n45848 = n60867 & n45847;
  assign n45849 = n60076 & n45846;
  assign po260 = n45030 & n60870;
  assign n45851 = ~n31605 & n44774;
  assign n45852 = ~n44910 & ~n45851;
  assign n45853 = ~pi205 & n45852;
  assign n45854 = n58992 & n31782;
  assign n45855 = ~n44777 & ~n45854;
  assign n45856 = ~pi202 & n45855;
  assign n45857 = ~pi233 & ~n45856;
  assign n45858 = ~pi233 & ~n45853;
  assign n45859 = ~n45856 & n45858;
  assign n45860 = ~n45853 & n45857;
  assign n45861 = ~pi204 & n45852;
  assign n45862 = ~pi201 & n45855;
  assign n45863 = pi233 & ~n45862;
  assign n45864 = pi233 & ~n45861;
  assign n45865 = ~n45862 & n45864;
  assign n45866 = ~n45861 & n45863;
  assign n45867 = ~n60879 & ~n60880;
  assign n45868 = pi237 & ~n45867;
  assign n45869 = ~pi218 & n45852;
  assign n45870 = ~pi203 & n45855;
  assign n45871 = ~pi233 & ~n45870;
  assign n45872 = ~pi233 & ~n45869;
  assign n45873 = ~n45870 & n45872;
  assign n45874 = ~n45869 & n45871;
  assign n45875 = ~pi206 & n45852;
  assign n45876 = ~pi220 & n45855;
  assign n45877 = pi233 & ~n45876;
  assign n45878 = pi233 & ~n45875;
  assign n45879 = ~n45876 & n45878;
  assign n45880 = ~n45875 & n45877;
  assign n45881 = ~n60881 & ~n60882;
  assign n45882 = ~pi237 & ~n45881;
  assign po746 = ~n45868 & ~n45882;
  assign n45884 = ~pi211 & ~n58992;
  assign n45885 = ~pi219 & n45884;
  assign n45886 = ~n58992 & n36679;
  assign n45887 = ~n45452 & ~n60883;
  assign po635 = pi71 & ~n45887;
  assign n45889 = ~pi270 & ~pi277;
  assign n45890 = ~pi282 & n45889;
  assign n45891 = pi266 & ~pi269;
  assign n45892 = pi278 & pi279;
  assign n45893 = ~pi280 & n45892;
  assign n45894 = n45891 & n45893;
  assign n45895 = ~pi281 & n45894;
  assign n45896 = n45890 & n45895;
  assign n45897 = pi264 & ~n45896;
  assign n45898 = ~pi264 & n45896;
  assign po953 = ~n45897 & ~n45898;
  assign n45900 = n5138 & n28759;
  assign n45901 = ~n28604 & ~n45900;
  assign n45902 = ~pi982 & ~n6416;
  assign n45903 = n2878 & n5138;
  assign n45904 = ~n45902 & ~n45903;
  assign po981 = n2441 & ~n45904;
  assign po997 = ~pi33 & n30925;
  assign n45907 = n2797 & n5138;
  assign n45908 = pi951 & ~n45907;
  assign po986 = pi1092 & ~n45908;
  assign n45910 = ~pi832 & pi1091;
  assign n45911 = pi1162 & n45910;
  assign po989 = n5142 & n45911;
  assign n45913 = pi281 & ~n45894;
  assign po987 = ~n45895 & ~n45913;
  assign n45915 = pi833 & ~n2794;
  assign n45916 = ~n59143 & ~n45915;
  assign po1107 = n2761 & ~n2878;
  assign n45918 = ~pi786 & pi954;
  assign n45919 = ~pi24 & ~pi954;
  assign n45920 = pi24 & ~pi954;
  assign n45921 = pi786 & pi954;
  assign n45922 = ~n45920 & ~n45921;
  assign n45923 = ~n45918 & ~n45919;
  assign n45924 = ~pi920 & ~pi1093;
  assign n45925 = pi1093 & ~pi1139;
  assign n45926 = pi1093 & pi1139;
  assign n45927 = pi920 & ~pi1093;
  assign n45928 = ~n45926 & ~n45927;
  assign n45929 = ~n45924 & ~n45925;
  assign n45930 = pi1093 & pi1140;
  assign n45931 = pi921 & ~pi1093;
  assign n45932 = ~n45930 & ~n45931;
  assign n45933 = pi1093 & pi1145;
  assign n45934 = pi927 & ~pi1093;
  assign n45935 = ~pi927 & ~pi1093;
  assign n45936 = pi1093 & ~pi1145;
  assign n45937 = ~n45935 & ~n45936;
  assign n45938 = ~n45933 & ~n45934;
  assign n45939 = pi1093 & ~pi1136;
  assign n45940 = ~pi928 & ~pi1093;
  assign po1084 = ~n45939 & ~n45940;
  assign n45942 = pi1093 & pi1144;
  assign n45943 = pi929 & ~pi1093;
  assign n45944 = ~pi929 & ~pi1093;
  assign n45945 = pi1093 & ~pi1144;
  assign n45946 = ~n45944 & ~n45945;
  assign n45947 = ~n45942 & ~n45943;
  assign n45948 = pi1093 & pi1134;
  assign n45949 = pi930 & ~pi1093;
  assign n45950 = ~pi930 & ~pi1093;
  assign n45951 = pi1093 & ~pi1134;
  assign n45952 = ~n45950 & ~n45951;
  assign n45953 = ~n45948 & ~n45949;
  assign n45954 = pi1093 & pi1142;
  assign n45955 = pi932 & ~pi1093;
  assign n45956 = ~n45954 & ~n45955;
  assign n45957 = pi1093 & pi1137;
  assign n45958 = pi933 & ~pi1093;
  assign n45959 = ~n45957 & ~n45958;
  assign n45960 = pi1093 & pi1141;
  assign n45961 = pi935 & ~pi1093;
  assign n45962 = ~n45960 & ~n45961;
  assign n45963 = pi1093 & pi1135;
  assign n45964 = pi938 & ~pi1093;
  assign n45965 = ~n45963 & ~n45964;
  assign n45966 = pi1093 & pi1146;
  assign n45967 = pi939 & ~pi1093;
  assign n45968 = ~pi939 & ~pi1093;
  assign n45969 = pi1093 & ~pi1146;
  assign n45970 = ~n45968 & ~n45969;
  assign n45971 = ~n45966 & ~n45967;
  assign n45972 = pi1093 & pi1138;
  assign n45973 = pi940 & ~pi1093;
  assign n45974 = ~n45972 & ~n45973;
  assign n45975 = ~pi944 & ~pi1093;
  assign n45976 = pi1093 & ~pi1143;
  assign n45977 = pi1093 & pi1143;
  assign n45978 = pi944 & ~pi1093;
  assign n45979 = ~n45977 & ~n45978;
  assign n45980 = ~n45975 & ~n45976;
  assign n45981 = pi957 & pi1092;
  assign n45982 = ~pi31 & ~n45981;
  assign po1135 = pi824 & pi1092;
  assign n45984 = ~pi567 & pi1092;
  assign n45985 = ~pi1093 & n45984;
  assign n45986 = pi680 & n7433;
  assign n45987 = ~n59304 & n45986;
  assign n45988 = ~n45985 & ~n45987;
  assign n45989 = n9554 & ~n45988;
  assign n45990 = pi788 & ~n7983;
  assign n45991 = ~n7716 & n45990;
  assign n45992 = n45989 & n45991;
  assign n45993 = ~n45985 & ~n45992;
  assign n45994 = ~n7913 & ~n45993;
  assign n45995 = pi603 & n6731;
  assign n45996 = ~n59346 & n45995;
  assign n45997 = pi603 & ~n7597;
  assign n45998 = n6731 & ~n59346;
  assign n45999 = ~n59347 & n45998;
  assign n46000 = n45997 & n45999;
  assign n46001 = n10748 & n45996;
  assign n46002 = n10740 & n60891;
  assign n46003 = n7716 & ~n45985;
  assign n46004 = ~pi619 & n60891;
  assign n46005 = ~n45985 & ~n46004;
  assign n46006 = ~pi1159 & ~n46005;
  assign n46007 = pi619 & n60891;
  assign n46008 = ~n45985 & ~n46007;
  assign n46009 = pi1159 & ~n46008;
  assign n46010 = pi789 & ~n46009;
  assign n46011 = pi789 & ~n46006;
  assign n46012 = ~n46009 & n46011;
  assign n46013 = ~n46006 & n46010;
  assign n46014 = ~n7715 & n60892;
  assign n46015 = ~n46002 & n46003;
  assign n46016 = n59242 & n45989;
  assign n46017 = ~n60893 & n46016;
  assign n46018 = ~n10741 & n60891;
  assign n46019 = ~pi789 & ~n45985;
  assign n46020 = ~n60891 & n46019;
  assign n46021 = ~n60892 & ~n46020;
  assign n46022 = ~n45985 & ~n46018;
  assign n46023 = ~n8054 & n60894;
  assign n46024 = ~n46017 & ~n46023;
  assign n46025 = n45989 & ~n60893;
  assign n46026 = ~n60894 & ~n46025;
  assign n46027 = n59242 & ~n46026;
  assign n46028 = n12139 & n60894;
  assign n46029 = ~n7716 & n45989;
  assign n46030 = pi641 & n46029;
  assign n46031 = ~n45985 & ~n46030;
  assign n46032 = n7911 & ~n46031;
  assign n46033 = ~pi641 & n46029;
  assign n46034 = ~n45985 & ~n46033;
  assign n46035 = n7912 & ~n46034;
  assign n46036 = ~n46032 & ~n46035;
  assign n46037 = ~n46028 & n46036;
  assign n46038 = pi788 & ~n46037;
  assign n46039 = ~n46027 & ~n46038;
  assign n46040 = ~n45994 & n46024;
  assign n46041 = ~n59357 & ~n60895;
  assign n46042 = n9651 & n45989;
  assign n46043 = ~n7762 & n46029;
  assign n46044 = n9652 & ~n45988;
  assign n46045 = pi628 & n60896;
  assign n46046 = ~n45985 & ~n46045;
  assign n46047 = pi1156 & ~n46046;
  assign n46048 = n8054 & ~n45985;
  assign n46049 = n8054 & n45985;
  assign n46050 = ~n46023 & ~n46049;
  assign n46051 = n60894 & ~n46048;
  assign n46052 = n7958 & ~n60897;
  assign n46053 = ~pi629 & ~n46052;
  assign n46054 = ~pi629 & ~n46047;
  assign n46055 = ~n46052 & n46054;
  assign n46056 = ~n46047 & n46053;
  assign n46057 = ~pi628 & n60896;
  assign n46058 = ~n45985 & ~n46057;
  assign n46059 = ~pi1156 & ~n46058;
  assign n46060 = n7957 & ~n60897;
  assign n46061 = pi629 & ~n46060;
  assign n46062 = pi629 & ~n46059;
  assign n46063 = ~n46060 & n46062;
  assign n46064 = ~n46059 & n46061;
  assign n46065 = pi792 & ~n60899;
  assign n46066 = pi792 & ~n60898;
  assign n46067 = ~n60899 & n46066;
  assign n46068 = ~n60898 & n46065;
  assign n46069 = ~n46041 & ~n60900;
  assign n46070 = ~pi647 & ~n46069;
  assign n46071 = n7793 & ~n45985;
  assign n46072 = ~n7793 & ~n60897;
  assign n46073 = n7793 & n45985;
  assign n46074 = ~n46072 & ~n46073;
  assign n46075 = ~n7793 & n60897;
  assign n46076 = ~n46071 & ~n46075;
  assign n46077 = ~n60897 & ~n46071;
  assign n46078 = pi647 & ~n60901;
  assign n46079 = ~pi1157 & ~n46078;
  assign n46080 = ~n46070 & n46079;
  assign n46081 = ~n59240 & n60896;
  assign n46082 = pi647 & n46081;
  assign n46083 = pi1157 & ~n45985;
  assign n46084 = ~n46082 & n46083;
  assign n46085 = ~pi630 & ~n46084;
  assign n46086 = ~n46080 & n46085;
  assign n46087 = pi647 & ~n46069;
  assign n46088 = ~pi647 & ~n60901;
  assign n46089 = pi1157 & ~n46088;
  assign n46090 = ~n46087 & n46089;
  assign n46091 = ~pi647 & n46081;
  assign n46092 = ~pi1157 & ~n45985;
  assign n46093 = ~n46091 & n46092;
  assign n46094 = pi630 & ~n46093;
  assign n46095 = ~n46090 & n46094;
  assign n46096 = ~n46086 & ~n46095;
  assign n46097 = pi787 & ~n46096;
  assign n46098 = ~pi787 & ~n46069;
  assign n46099 = ~n46097 & ~n46098;
  assign n46100 = ~pi644 & ~n46099;
  assign n46101 = ~n9743 & n46081;
  assign n46102 = ~n45985 & ~n46101;
  assign n46103 = pi644 & ~n46102;
  assign n46104 = ~pi715 & ~n46103;
  assign n46105 = ~n46100 & n46104;
  assign n46106 = ~n7835 & n46072;
  assign n46107 = n11491 & ~n60897;
  assign n46108 = ~pi644 & n60902;
  assign n46109 = pi715 & ~n45985;
  assign n46110 = ~n46108 & n46109;
  assign n46111 = ~pi1160 & ~n46110;
  assign n46112 = ~n46105 & n46111;
  assign n46113 = pi644 & ~n46099;
  assign n46114 = ~pi644 & ~n46102;
  assign n46115 = pi715 & ~n46114;
  assign n46116 = ~n46113 & n46115;
  assign n46117 = pi644 & n60902;
  assign n46118 = ~pi715 & ~n45985;
  assign n46119 = ~n46117 & n46118;
  assign n46120 = pi1160 & ~n46119;
  assign n46121 = ~n46116 & n46120;
  assign n46122 = ~n46112 & ~n46121;
  assign n46123 = ~n46105 & ~n46110;
  assign n46124 = ~pi1160 & ~n46123;
  assign n46125 = pi644 & n46099;
  assign n46126 = ~pi644 & n46102;
  assign n46127 = pi715 & ~n46126;
  assign n46128 = ~n46125 & n46127;
  assign n46129 = ~n45985 & ~n46117;
  assign n46130 = ~pi715 & ~n46129;
  assign n46131 = pi1160 & ~n46130;
  assign n46132 = ~n46128 & n46131;
  assign n46133 = pi790 & ~n46132;
  assign n46134 = ~n46124 & n46133;
  assign n46135 = pi790 & ~n46122;
  assign n46136 = ~pi790 & ~n46099;
  assign n46137 = ~n60903 & ~n46136;
  assign n46138 = pi230 & ~n46137;
  assign n46139 = ~pi230 & n45984;
  assign n46140 = ~n46138 & ~n46139;
  assign n46141 = pi243 & ~pi1091;
  assign n46142 = ~pi83 & ~pi85;
  assign n46143 = pi314 & ~n46142;
  assign n46144 = pi802 & n46143;
  assign n46145 = pi276 & n46144;
  assign n46146 = ~pi1091 & ~n46145;
  assign n46147 = pi271 & ~n46146;
  assign n46148 = ~pi1091 & ~n46147;
  assign n46149 = pi273 & ~n46148;
  assign n46150 = ~pi1091 & ~n46149;
  assign n46151 = ~pi200 & ~n46150;
  assign n46152 = pi199 & ~n46150;
  assign n46153 = ~pi81 & n46142;
  assign n46154 = pi314 & ~n46153;
  assign n46155 = pi802 & n46154;
  assign n46156 = pi276 & n46155;
  assign n46157 = ~pi1091 & n46156;
  assign n46158 = pi271 & n46157;
  assign n46159 = pi273 & n46158;
  assign n46160 = ~n46149 & ~n46159;
  assign n46161 = ~pi1091 & n46160;
  assign n46162 = ~pi199 & ~n46161;
  assign n46163 = ~n46152 & ~n46162;
  assign n46164 = n46157 & ~n46163;
  assign n46165 = ~pi299 & ~n46164;
  assign n46166 = ~n46152 & n46165;
  assign n46167 = ~n46151 & n46166;
  assign n46168 = pi299 & ~n46159;
  assign n46169 = ~n46167 & ~n46168;
  assign n46170 = ~n46141 & ~n46169;
  assign n46171 = pi299 & n46150;
  assign n46172 = ~n46159 & n46171;
  assign n46173 = ~pi200 & ~n46157;
  assign n46174 = ~n46163 & ~n46173;
  assign n46175 = ~pi299 & ~n46174;
  assign n46176 = ~n46162 & n46175;
  assign n46177 = ~n46167 & ~n46176;
  assign n46178 = ~n46172 & n46177;
  assign n46179 = ~pi243 & ~n46178;
  assign n46180 = ~n46152 & n46175;
  assign n46181 = ~n46168 & ~n46180;
  assign n46182 = ~n46151 & n46165;
  assign n46183 = ~n46162 & n46182;
  assign n46184 = pi243 & ~n46183;
  assign n46185 = n46181 & n46184;
  assign n46186 = ~n46179 & ~n46185;
  assign n46187 = ~pi1155 & ~n46186;
  assign n46188 = ~pi1091 & n46145;
  assign n46189 = pi271 & n46188;
  assign n46190 = pi273 & n46189;
  assign n46191 = pi299 & ~n46190;
  assign n46192 = ~n46183 & ~n46191;
  assign n46193 = ~n46180 & n46192;
  assign n46194 = ~n46171 & ~n46182;
  assign n46195 = pi243 & ~n46194;
  assign n46196 = ~n46193 & n46195;
  assign n46197 = pi1155 & ~n46196;
  assign n46198 = ~n46172 & ~n46183;
  assign n46199 = pi1155 & n46198;
  assign n46200 = ~n46197 & ~n46199;
  assign n46201 = ~n46168 & ~n46175;
  assign n46202 = ~pi243 & n46201;
  assign n46203 = ~n46172 & ~n46175;
  assign n46204 = n46169 & n46203;
  assign n46205 = ~n46167 & n46201;
  assign n46206 = ~pi243 & n60904;
  assign n46207 = ~n46167 & n46202;
  assign n46208 = ~n46200 & ~n60905;
  assign n46209 = ~n46187 & ~n46208;
  assign n46210 = ~n46170 & n46209;
  assign n46211 = pi1156 & ~n46210;
  assign n46212 = ~n46171 & ~n46176;
  assign n46213 = ~pi243 & ~n46212;
  assign n46214 = ~pi1155 & ~n46213;
  assign n46215 = ~n46165 & ~n46168;
  assign n46216 = ~pi1155 & n46215;
  assign n46217 = ~n46214 & ~n46216;
  assign n46218 = ~n46168 & ~n46182;
  assign n46219 = pi243 & n46218;
  assign n46220 = ~n46166 & ~n46168;
  assign n46221 = ~n46182 & n46220;
  assign n46222 = pi243 & n46221;
  assign n46223 = ~n46166 & n46219;
  assign n46224 = ~n46217 & ~n60906;
  assign n46225 = ~pi1156 & ~n46224;
  assign n46226 = ~pi243 & ~n46203;
  assign n46227 = pi1155 & ~n46226;
  assign n46228 = ~n46219 & n46227;
  assign n46229 = n46225 & ~n46228;
  assign n46230 = pi1157 & ~n46229;
  assign n46231 = ~n46211 & n46230;
  assign n46232 = pi243 & n46215;
  assign n46233 = ~pi243 & ~pi1091;
  assign n46234 = ~n46165 & ~n46191;
  assign n46235 = n46233 & ~n46234;
  assign n46236 = ~pi1155 & ~n46235;
  assign n46237 = ~n46216 & ~n46236;
  assign n46238 = ~n46232 & ~n46237;
  assign n46239 = ~pi1156 & ~n46238;
  assign n46240 = pi1155 & ~n46141;
  assign n46241 = n46152 & n46240;
  assign n46242 = ~n46228 & ~n46241;
  assign n46243 = n46239 & n46242;
  assign n46244 = ~n46162 & n46165;
  assign n46245 = ~n46172 & ~n46244;
  assign n46246 = pi243 & ~n46245;
  assign n46247 = ~pi243 & n46220;
  assign n46248 = ~n46246 & ~n46247;
  assign n46249 = ~pi1155 & n46218;
  assign n46250 = ~n46157 & n46249;
  assign n46251 = pi1156 & ~n46250;
  assign n46252 = n46248 & n46251;
  assign n46253 = ~pi1157 & ~n46252;
  assign n46254 = ~n46243 & n46253;
  assign n46255 = pi211 & ~n46254;
  assign n46256 = ~n46231 & n46255;
  assign n46257 = pi1156 & ~n46209;
  assign n46258 = ~n46172 & ~n46182;
  assign n46259 = pi243 & ~n46258;
  assign n46260 = ~n46202 & ~n46259;
  assign n46261 = n46225 & n46260;
  assign n46262 = pi1157 & ~n46261;
  assign n46263 = ~n46257 & n46262;
  assign n46264 = n46248 & n46260;
  assign n46265 = pi1155 & ~n46264;
  assign n46266 = n46239 & ~n46265;
  assign n46267 = ~pi1155 & n46258;
  assign n46268 = ~n46201 & n46267;
  assign n46269 = n46252 & ~n46268;
  assign n46270 = ~pi1157 & ~n46269;
  assign n46271 = ~n46266 & n46270;
  assign n46272 = ~pi211 & ~n46271;
  assign n46273 = ~n46263 & n46272;
  assign n46274 = ~pi219 & ~n46273;
  assign n46275 = ~n46256 & n46274;
  assign n46276 = pi253 & pi254;
  assign n46277 = pi267 & n46276;
  assign n46278 = ~pi263 & n46277;
  assign n46279 = ~n46167 & ~n46171;
  assign n46280 = ~pi243 & n46279;
  assign n46281 = ~n46175 & ~n46191;
  assign n46282 = n46280 & n46281;
  assign n46283 = n46197 & ~n46282;
  assign n46284 = pi243 & ~n46193;
  assign n46285 = ~n46280 & ~n46284;
  assign n46286 = ~n46170 & ~n46213;
  assign n46287 = ~n46285 & n46286;
  assign n46288 = ~pi1155 & ~n46287;
  assign n46289 = ~n46283 & ~n46288;
  assign n46290 = pi1156 & ~n46289;
  assign n46291 = ~pi211 & pi1157;
  assign n46292 = ~n46176 & ~n46191;
  assign n46293 = ~pi243 & ~n46292;
  assign n46294 = pi243 & ~n46166;
  assign n46295 = ~pi1155 & ~n46294;
  assign n46296 = ~n46293 & n46295;
  assign n46297 = ~pi243 & pi1155;
  assign n46298 = n46281 & n46297;
  assign n46299 = ~pi1156 & ~n46298;
  assign n46300 = ~n46195 & n46299;
  assign n46301 = ~n46296 & n46300;
  assign n46302 = n46291 & ~n46301;
  assign n46303 = ~n46290 & n46302;
  assign n46304 = pi243 & n46192;
  assign n46305 = n46227 & ~n46304;
  assign n46306 = ~n46214 & ~n46305;
  assign n46307 = ~n46285 & ~n46306;
  assign n46308 = pi1156 & ~n46307;
  assign n46309 = pi211 & pi1157;
  assign n46310 = ~n46182 & ~n46191;
  assign n46311 = pi243 & n46310;
  assign n46312 = ~n46226 & ~n46311;
  assign n46313 = pi1155 & ~n46312;
  assign n46314 = ~n46166 & n46310;
  assign n46315 = pi243 & n46314;
  assign n46316 = n46294 & n46310;
  assign n46317 = ~n46213 & ~n60907;
  assign n46318 = ~n46313 & n46317;
  assign n46319 = ~pi1156 & ~n46318;
  assign n46320 = n46309 & ~n46319;
  assign n46321 = ~n46308 & n46320;
  assign n46322 = ~n46191 & ~n46244;
  assign n46323 = pi1155 & n46322;
  assign n46324 = ~n46175 & n46322;
  assign n46325 = ~n46323 & ~n46324;
  assign n46326 = pi243 & ~n46325;
  assign n46327 = ~n46166 & ~n46171;
  assign n46328 = ~pi243 & ~n46327;
  assign n46329 = ~n46250 & n46328;
  assign n46330 = ~n46326 & ~n46329;
  assign n46331 = pi1156 & ~n46330;
  assign n46332 = ~n46244 & n46311;
  assign n46333 = ~n46171 & ~n46180;
  assign n46334 = ~pi243 & ~n46333;
  assign n46335 = pi1155 & ~n46334;
  assign n46336 = ~n46332 & n46335;
  assign n46337 = pi243 & n46234;
  assign n46338 = n46236 & ~n46337;
  assign n46339 = ~pi1156 & ~n46338;
  assign n46340 = ~n46336 & n46339;
  assign n46341 = ~pi1157 & ~n46340;
  assign n46342 = ~n46331 & n46341;
  assign n46343 = ~n46321 & ~n46342;
  assign n46344 = ~n46303 & n46343;
  assign n46345 = pi219 & ~n46344;
  assign n46346 = n46278 & ~n46345;
  assign n46347 = ~n46275 & n46346;
  assign n46348 = pi199 & pi200;
  assign n46349 = ~pi1155 & n36719;
  assign n46350 = ~n46348 & ~n60908;
  assign n46351 = ~pi299 & pi1091;
  assign n46352 = n46350 & n46351;
  assign n46353 = ~n46233 & ~n46352;
  assign n46354 = pi199 & pi1091;
  assign n46355 = ~pi299 & n46354;
  assign n46356 = n46240 & ~n46355;
  assign n46357 = pi1156 & ~n46356;
  assign n46358 = n46353 & n46357;
  assign n46359 = pi199 & ~pi200;
  assign n46360 = ~pi299 & n46359;
  assign n46361 = pi1091 & ~n46360;
  assign n46362 = ~n46141 & ~n46361;
  assign n46363 = ~pi1155 & n46362;
  assign n46364 = pi200 & pi1091;
  assign n46365 = pi200 & ~pi299;
  assign n46366 = pi1091 & n46365;
  assign n46367 = ~pi299 & n46364;
  assign n46368 = n46240 & ~n60909;
  assign n46369 = ~pi1156 & ~n46368;
  assign n46370 = ~n46363 & n46369;
  assign n46371 = ~n46358 & ~n46370;
  assign n46372 = pi1157 & ~n46371;
  assign n46373 = ~pi1155 & ~n46141;
  assign n46374 = pi1091 & ~n45425;
  assign n46375 = n46373 & ~n46374;
  assign n46376 = ~n46356 & ~n46375;
  assign n46377 = pi200 & ~pi1156;
  assign n46378 = n46351 & n46377;
  assign n46379 = ~n46376 & ~n46378;
  assign n46380 = ~pi1157 & ~n46379;
  assign n46381 = ~pi211 & ~n46380;
  assign n46382 = ~n46372 & n46381;
  assign n46383 = pi1156 & ~n46353;
  assign n46384 = ~pi299 & n46348;
  assign n46385 = pi1156 & ~n46384;
  assign n46386 = pi1091 & ~n45444;
  assign n46387 = n46385 & n46386;
  assign n46388 = ~n46383 & ~n46387;
  assign n46389 = ~pi200 & ~pi299;
  assign n46390 = ~pi1155 & ~n46233;
  assign n46391 = ~n46141 & ~n46390;
  assign n46392 = n46389 & n46391;
  assign n46393 = ~n46362 & ~n46392;
  assign n46394 = ~pi1156 & ~n46393;
  assign n46395 = pi1157 & ~n46394;
  assign n46396 = n46388 & n46395;
  assign n46397 = ~n45424 & n46351;
  assign n46398 = n46373 & ~n46397;
  assign n46399 = n46357 & ~n46398;
  assign n46400 = ~n46386 & n46391;
  assign n46401 = ~pi1156 & ~n46400;
  assign n46402 = ~n46399 & ~n46401;
  assign n46403 = ~pi1157 & ~n46402;
  assign n46404 = pi211 & ~n46403;
  assign n46405 = n46388 & ~n46394;
  assign n46406 = pi1157 & ~n46405;
  assign n46407 = ~pi1157 & ~n46399;
  assign n46408 = ~pi1157 & ~n46401;
  assign n46409 = ~n46399 & n46408;
  assign n46410 = ~n46401 & n46407;
  assign n46411 = ~n46406 & ~n60910;
  assign n46412 = pi211 & ~n46411;
  assign n46413 = ~n46396 & n46404;
  assign n46414 = ~n46382 & ~n60911;
  assign n46415 = ~pi219 & ~n46414;
  assign n46416 = pi299 & pi1091;
  assign n46417 = n46379 & ~n46416;
  assign n46418 = ~pi1157 & ~n46417;
  assign n46419 = pi219 & ~n46418;
  assign n46420 = n46309 & ~n46383;
  assign n46421 = ~n46394 & n46420;
  assign n46422 = ~pi299 & ~n46359;
  assign n46423 = pi1091 & n46422;
  assign n46424 = n46373 & ~n46423;
  assign n46425 = ~n46368 & ~n46424;
  assign n46426 = ~pi1156 & ~n46425;
  assign n46427 = n46291 & ~n46426;
  assign n46428 = n46388 & n46427;
  assign n46429 = ~n46421 & ~n46428;
  assign n46430 = pi219 & ~n46421;
  assign n46431 = ~n46418 & ~n46428;
  assign n46432 = n46430 & n46431;
  assign n46433 = n46419 & n46429;
  assign n46434 = ~n46415 & ~n60912;
  assign n46435 = ~n46278 & ~n46434;
  assign n46436 = n58992 & ~n46435;
  assign n46437 = ~n46347 & n46436;
  assign n46438 = pi272 & pi283;
  assign n46439 = pi275 & n46438;
  assign n46440 = pi268 & n46439;
  assign n46441 = pi243 & n46161;
  assign n46442 = n46141 & n46160;
  assign n46443 = pi211 & pi1156;
  assign n46444 = ~pi211 & pi1155;
  assign n46445 = ~n46443 & ~n46444;
  assign n46446 = pi1091 & n46445;
  assign n46447 = ~pi243 & n46159;
  assign n46448 = ~n46446 & ~n46447;
  assign n46449 = ~n60913 & n46448;
  assign n46450 = ~pi219 & ~n46449;
  assign n46451 = ~pi243 & n46150;
  assign n46452 = pi243 & n46190;
  assign n46453 = ~n46141 & n46291;
  assign n46454 = ~n46188 & n46453;
  assign n46455 = pi219 & ~n46454;
  assign n46456 = ~n46452 & n46455;
  assign n46457 = ~n46451 & n46456;
  assign n46458 = n46278 & ~n46457;
  assign n46459 = ~n46452 & ~n46454;
  assign n46460 = ~n46451 & n46459;
  assign n46461 = pi219 & ~n46460;
  assign n46462 = ~pi219 & ~n46446;
  assign n46463 = ~n46447 & n46462;
  assign n46464 = ~n60913 & n46463;
  assign n46465 = ~n46461 & ~n46464;
  assign n46466 = n46278 & ~n46465;
  assign n46467 = ~n46450 & n46458;
  assign n46468 = ~pi219 & ~n46445;
  assign n46469 = pi1157 & n36681;
  assign n46470 = pi219 & n46291;
  assign n46471 = ~n46468 & ~n60915;
  assign n46472 = pi1091 & ~n46471;
  assign n46473 = ~n46233 & ~n46472;
  assign n46474 = ~n46278 & ~n46473;
  assign n46475 = ~n58992 & ~n46474;
  assign n46476 = ~n60914 & n46475;
  assign n46477 = n46440 & ~n46476;
  assign n46478 = ~n46437 & n46477;
  assign n46479 = n58992 & n46434;
  assign n46480 = ~n58992 & n46473;
  assign n46481 = ~n46440 & ~n46480;
  assign n46482 = ~n46479 & n46481;
  assign n46483 = ~pi230 & ~n46482;
  assign n46484 = ~n46478 & n46483;
  assign n46485 = ~pi200 & pi1157;
  assign n46486 = pi199 & ~n46485;
  assign n46487 = ~n60908 & ~n46377;
  assign n46488 = ~n46486 & n46487;
  assign n46489 = n44774 & n46488;
  assign n46490 = ~n44774 & ~n46471;
  assign n46491 = pi230 & ~n46490;
  assign n46492 = pi230 & ~n46489;
  assign n46493 = ~n46490 & n46492;
  assign n46494 = ~n46489 & n46491;
  assign po400 = ~n46484 & ~n60916;
  assign n46496 = pi1154 & ~n36720;
  assign n46497 = pi200 & ~pi1155;
  assign n46498 = ~n36719 & ~n46348;
  assign n46499 = ~pi299 & n46498;
  assign n46500 = ~pi1156 & ~n46365;
  assign n46501 = n46499 & ~n46500;
  assign n46502 = ~n46497 & n46501;
  assign n46503 = ~n46496 & ~n46502;
  assign n46504 = ~pi211 & ~n46503;
  assign n46505 = ~pi219 & ~n46504;
  assign n46506 = pi299 & pi1155;
  assign n46507 = ~pi199 & pi1155;
  assign n46508 = pi200 & ~n46507;
  assign n46509 = ~pi299 & ~n46508;
  assign n46510 = ~pi199 & pi1154;
  assign n46511 = pi199 & pi1156;
  assign n46512 = ~pi200 & ~n46511;
  assign n46513 = ~n46510 & n46512;
  assign n46514 = pi1156 & n46359;
  assign n46515 = ~pi200 & ~pi1154;
  assign n46516 = ~pi199 & ~n46497;
  assign n46517 = ~n46515 & n46516;
  assign n46518 = ~n46514 & ~n46517;
  assign n46519 = ~pi299 & ~n46518;
  assign n46520 = n46365 & n46507;
  assign n46521 = ~pi1154 & ~n46520;
  assign n46522 = n45518 & ~n46497;
  assign n46523 = ~n46521 & n46522;
  assign n46524 = ~pi1156 & ~n46523;
  assign n46525 = ~pi199 & ~pi1154;
  assign n46526 = ~pi200 & n46525;
  assign n46527 = n46509 & ~n60918;
  assign n46528 = ~n46524 & n46527;
  assign n46529 = n46509 & ~n46513;
  assign n46530 = ~n46506 & ~n60917;
  assign n46531 = pi211 & ~n46530;
  assign n46532 = n46505 & ~n46531;
  assign n46533 = pi1156 & n45445;
  assign n46534 = pi219 & ~n46533;
  assign n46535 = pi1154 & ~n46508;
  assign n46536 = pi1156 & ~n46535;
  assign n46537 = ~pi299 & ~n46536;
  assign n46538 = n36720 & ~n46508;
  assign n46539 = ~pi1154 & n46538;
  assign n46540 = ~n45445 & ~n46539;
  assign n46541 = ~n46537 & n46540;
  assign n46542 = pi1156 & ~n46541;
  assign n46543 = ~n46496 & ~n46520;
  assign n46544 = n46537 & ~n46543;
  assign n46545 = pi219 & ~n46544;
  assign n46546 = ~n46542 & n46545;
  assign n46547 = ~n60917 & n46534;
  assign n46548 = n58992 & ~n60919;
  assign n46549 = ~n46532 & n46548;
  assign n46550 = ~pi211 & pi1156;
  assign n46551 = pi219 & ~n46550;
  assign n46552 = ~pi211 & pi1154;
  assign n46553 = pi211 & pi1155;
  assign n46554 = ~pi219 & ~n46553;
  assign n46555 = ~n46552 & n46554;
  assign n46556 = ~n46551 & ~n46555;
  assign n46557 = ~n58992 & n46556;
  assign n46558 = pi230 & ~n46557;
  assign n46559 = ~n46549 & n46558;
  assign n46560 = ~pi1091 & ~n46322;
  assign n46561 = ~pi1155 & n46560;
  assign n46562 = ~n46245 & n46561;
  assign n46563 = pi1155 & ~n46169;
  assign n46564 = ~pi1154 & ~n46563;
  assign n46565 = ~n46562 & n46564;
  assign n46566 = ~pi1156 & ~n46565;
  assign n46567 = pi1155 & ~n46279;
  assign n46568 = ~pi1154 & ~n46567;
  assign n46569 = ~n46561 & n46568;
  assign n46570 = pi1155 & ~n46220;
  assign n46571 = pi1154 & ~n46570;
  assign n46572 = n46181 & n46571;
  assign n46573 = ~n46569 & ~n46572;
  assign n46574 = n46566 & n46573;
  assign n46575 = ~pi1155 & n46212;
  assign n46576 = ~n46168 & n46177;
  assign n46577 = ~n46575 & ~n46576;
  assign n46578 = ~pi1154 & ~n46577;
  assign n46579 = pi1156 & ~n46578;
  assign n46580 = n46212 & n46568;
  assign n46581 = ~n46173 & n46572;
  assign n46582 = ~n46580 & ~n46581;
  assign n46583 = n46579 & n46582;
  assign n46584 = ~pi211 & ~n46583;
  assign n46585 = ~pi211 & ~n46574;
  assign n46586 = ~n46583 & n46585;
  assign n46587 = ~n46574 & n46584;
  assign n46588 = n46203 & n46571;
  assign n46589 = n46579 & ~n46588;
  assign n46590 = ~n46172 & ~n46180;
  assign n46591 = n46571 & n46590;
  assign n46592 = n46566 & ~n46591;
  assign n46593 = pi211 & ~n46592;
  assign n46594 = pi211 & ~n46589;
  assign n46595 = ~n46592 & n46594;
  assign n46596 = ~n46589 & n46593;
  assign n46597 = ~pi219 & ~n60921;
  assign n46598 = ~pi219 & ~n60920;
  assign n46599 = ~n60921 & n46598;
  assign n46600 = ~n60920 & n46597;
  assign n46601 = pi1155 & n46167;
  assign n46602 = pi1154 & n46333;
  assign n46603 = ~n46601 & n46602;
  assign n46604 = ~n46569 & ~n46603;
  assign n46605 = ~pi1156 & ~n46604;
  assign n46606 = ~n46175 & n46603;
  assign n46607 = ~n46580 & ~n46606;
  assign n46608 = n46443 & ~n46607;
  assign n46609 = ~pi1154 & n46322;
  assign n46610 = ~n46281 & ~n46609;
  assign n46611 = n46550 & ~n46601;
  assign n46612 = ~n46610 & n46611;
  assign n46613 = pi219 & ~n46612;
  assign n46614 = ~n46608 & n46613;
  assign n46615 = ~n46605 & n46613;
  assign n46616 = ~n46608 & n46615;
  assign n46617 = ~n46605 & n46614;
  assign n46618 = ~pi263 & ~n60923;
  assign n46619 = ~n60922 & n46618;
  assign n46620 = ~n46199 & ~n46267;
  assign n46621 = ~n46176 & ~n46620;
  assign n46622 = ~pi1156 & ~n46621;
  assign n46623 = pi211 & n46249;
  assign n46624 = ~pi211 & n46267;
  assign n46625 = ~n46199 & ~n46624;
  assign n46626 = ~n46623 & n46625;
  assign n46627 = pi1154 & ~n46626;
  assign n46628 = ~n46622 & n46627;
  assign n46629 = pi1156 & n46221;
  assign n46630 = ~n46175 & n46245;
  assign n46631 = n46553 & n46630;
  assign n46632 = n46201 & ~n46244;
  assign n46633 = n46444 & n46632;
  assign n46634 = ~n46216 & ~n46633;
  assign n46635 = ~n46631 & n46634;
  assign n46636 = ~n46629 & n46635;
  assign n46637 = ~pi1154 & ~n46636;
  assign n46638 = ~n46628 & ~n46637;
  assign n46639 = pi1154 & ~n46199;
  assign n46640 = ~n46249 & n46639;
  assign n46641 = ~pi1154 & ~n46216;
  assign n46642 = pi1155 & n46630;
  assign n46643 = n46641 & ~n46642;
  assign n46644 = ~n46267 & n46639;
  assign n46645 = pi1154 & n46176;
  assign n46646 = ~pi1156 & ~n46645;
  assign n46647 = ~n46644 & n46646;
  assign n46648 = ~pi1156 & ~n46647;
  assign n46649 = ~n46643 & ~n46648;
  assign n46650 = ~n46629 & ~n46649;
  assign n46651 = ~n46640 & ~n46650;
  assign n46652 = pi211 & ~n46651;
  assign n46653 = pi1155 & n46632;
  assign n46654 = n46641 & ~n46653;
  assign n46655 = n46647 & ~n46654;
  assign n46656 = ~n46221 & n46654;
  assign n46657 = pi1156 & ~n46656;
  assign n46658 = ~n46644 & n46657;
  assign n46659 = ~pi211 & ~n46658;
  assign n46660 = ~n46655 & n46659;
  assign n46661 = ~pi219 & ~n46660;
  assign n46662 = ~n46652 & n46661;
  assign n46663 = ~pi219 & ~n46638;
  assign n46664 = ~n46183 & n46333;
  assign n46665 = pi1155 & ~n46664;
  assign n46666 = ~n46182 & n46327;
  assign n46667 = ~pi1155 & ~n46666;
  assign n46668 = ~pi1154 & ~n46667;
  assign n46669 = ~pi1154 & ~n46665;
  assign n46670 = ~n46667 & n46669;
  assign n46671 = ~n46665 & n46668;
  assign n46672 = ~n46194 & ~n46323;
  assign n46673 = pi1154 & ~n46672;
  assign n46674 = n46550 & ~n46673;
  assign n46675 = ~n60925 & n46674;
  assign n46676 = pi1154 & n46180;
  assign n46677 = ~n46193 & ~n46676;
  assign n46678 = ~pi1156 & n46244;
  assign n46679 = ~n46672 & ~n46678;
  assign n46680 = ~n46677 & n46679;
  assign n46681 = ~n46550 & ~n46680;
  assign n46682 = pi219 & ~n46681;
  assign n46683 = ~n46672 & ~n46677;
  assign n46684 = ~n46244 & n46683;
  assign n46685 = ~pi1156 & ~n46684;
  assign n46686 = n46443 & ~n46683;
  assign n46687 = pi219 & ~n46686;
  assign n46688 = pi219 & ~n46675;
  assign n46689 = ~n46686 & n46688;
  assign n46690 = ~n46675 & n46687;
  assign n46691 = ~n46685 & n60926;
  assign n46692 = ~n46675 & n46682;
  assign n46693 = pi263 & ~n60927;
  assign n46694 = ~n60924 & n46693;
  assign n46695 = n46277 & ~n46694;
  assign n46696 = n46277 & ~n46619;
  assign n46697 = ~n46694 & n46696;
  assign n46698 = ~n46619 & n46695;
  assign n46699 = pi1155 & ~n46384;
  assign n46700 = n60909 & ~n46699;
  assign n46701 = pi1091 & ~n46499;
  assign n46702 = ~pi1154 & n46701;
  assign n46703 = ~n46700 & ~n46702;
  assign n46704 = ~pi211 & ~n46703;
  assign n46705 = ~pi299 & ~n45424;
  assign n46706 = pi1155 & ~n46705;
  assign n46707 = pi211 & pi1091;
  assign n46708 = n46389 & ~n46525;
  assign n46709 = n46707 & ~n46708;
  assign n46710 = ~n46706 & n46709;
  assign n46711 = pi1156 & ~n46710;
  assign n46712 = ~n46704 & n46711;
  assign n46713 = pi1091 & ~pi1154;
  assign n46714 = ~n46386 & ~n46713;
  assign n46715 = ~n46706 & ~n46714;
  assign n46716 = pi211 & n46715;
  assign n46717 = ~pi211 & pi1091;
  assign n46718 = ~n46520 & n46717;
  assign n46719 = n46543 & n46717;
  assign n46720 = ~n46496 & n46718;
  assign n46721 = ~pi1156 & ~n60929;
  assign n46722 = ~n46716 & n46721;
  assign n46723 = ~n46712 & ~n46722;
  assign n46724 = ~n46704 & ~n46710;
  assign n46725 = pi1156 & ~n46724;
  assign n46726 = ~n46716 & ~n60929;
  assign n46727 = ~pi1156 & ~n46726;
  assign n46728 = ~pi219 & ~n46727;
  assign n46729 = ~n46725 & n46728;
  assign n46730 = ~pi219 & ~n46723;
  assign n46731 = ~n46416 & n46703;
  assign n46732 = n46443 & ~n46731;
  assign n46733 = ~pi1156 & ~n46520;
  assign n46734 = ~n46714 & n46733;
  assign n46735 = pi200 & n46507;
  assign n46736 = ~pi299 & ~n46498;
  assign n46737 = pi1155 & ~n46736;
  assign n46738 = ~pi1155 & ~n46422;
  assign n46739 = ~n46737 & ~n46738;
  assign n46740 = n46422 & ~n46735;
  assign n46741 = ~pi1154 & ~n60931;
  assign n46742 = n46365 & ~n46507;
  assign n46743 = pi1154 & ~n46742;
  assign n46744 = pi1091 & n46550;
  assign n46745 = ~n46743 & n46744;
  assign n46746 = ~n46741 & n46745;
  assign n46747 = pi219 & ~n46746;
  assign n46748 = pi219 & ~n46734;
  assign n46749 = ~n46746 & n46748;
  assign n46750 = ~n46734 & n46747;
  assign n46751 = ~n46732 & n60932;
  assign n46752 = ~n60930 & ~n46751;
  assign n46753 = ~pi263 & ~n46752;
  assign n46754 = ~pi1155 & ~n36720;
  assign n46755 = n46741 & ~n46754;
  assign n46756 = pi1155 & ~n45521;
  assign n46757 = ~n46389 & ~n46756;
  assign n46758 = pi1154 & ~n46757;
  assign n46759 = pi1156 & ~n46758;
  assign n46760 = ~n46755 & n46759;
  assign n46761 = ~pi1156 & n46715;
  assign n46762 = pi211 & ~n46761;
  assign n46763 = ~n46760 & n46762;
  assign n46764 = n46505 & ~n46763;
  assign n46765 = pi263 & pi1091;
  assign n46766 = ~n60919 & n46765;
  assign n46767 = ~n46764 & n46766;
  assign n46768 = ~n46753 & ~n46767;
  assign n46769 = ~n46277 & ~n46768;
  assign n46770 = n58992 & ~n46769;
  assign n46771 = ~n60928 & n46770;
  assign n46772 = pi211 & n46150;
  assign n46773 = ~pi211 & ~n46713;
  assign n46774 = ~n46553 & ~n46773;
  assign n46775 = ~n46772 & n46774;
  assign n46776 = ~n46159 & ~n46775;
  assign n46777 = ~pi219 & ~n46776;
  assign n46778 = pi219 & ~n46150;
  assign n46779 = ~pi211 & ~n46188;
  assign n46780 = n46778 & ~n46779;
  assign n46781 = ~pi263 & ~n46780;
  assign n46782 = ~n46777 & n46781;
  assign n46783 = ~pi219 & ~n46159;
  assign n46784 = pi1154 & n46717;
  assign n46785 = ~n46553 & ~n46784;
  assign n46786 = ~n46772 & ~n46785;
  assign n46787 = n46783 & ~n46786;
  assign n46788 = ~pi211 & ~n46150;
  assign n46789 = pi211 & n46190;
  assign n46790 = pi219 & ~n46789;
  assign n46791 = ~n46788 & n46790;
  assign n46792 = pi263 & ~n46791;
  assign n46793 = ~n46787 & n46792;
  assign n46794 = ~n46782 & ~n46793;
  assign n46795 = pi1091 & n46551;
  assign n46796 = n46277 & ~n46795;
  assign n46797 = ~n46794 & n46796;
  assign n46798 = pi1091 & ~n46556;
  assign n46799 = pi263 & ~pi1091;
  assign n46800 = ~n46798 & ~n46799;
  assign n46801 = ~n46277 & n46800;
  assign n46802 = ~n58992 & ~n46801;
  assign n46803 = ~n46797 & n46802;
  assign n46804 = n46440 & ~n46803;
  assign n46805 = ~n46771 & n46804;
  assign n46806 = n58992 & n46768;
  assign n46807 = ~n58992 & ~n46800;
  assign n46808 = ~n46440 & ~n46807;
  assign n46809 = ~n46806 & n46808;
  assign n46810 = ~pi230 & ~n46809;
  assign n46811 = ~n46805 & n46810;
  assign po420 = ~n46559 & ~n46811;
  assign n46813 = ~pi1153 & n46245;
  assign n46814 = ~n46590 & ~n46813;
  assign n46815 = n46279 & ~n46814;
  assign n46816 = n46169 & ~n46815;
  assign n46817 = n46665 & ~n46816;
  assign n46818 = pi1154 & ~n46817;
  assign n46819 = ~pi1153 & ~n46220;
  assign n46820 = ~pi1154 & ~n46819;
  assign n46821 = pi1155 & ~n46820;
  assign n46822 = n46218 & ~n46821;
  assign n46823 = ~n46818 & ~n46822;
  assign n46824 = ~pi1153 & ~n46234;
  assign n46825 = ~n46182 & n46322;
  assign n46826 = ~n46824 & n46825;
  assign n46827 = ~pi1155 & ~n46630;
  assign n46828 = ~pi1155 & ~n46826;
  assign n46829 = ~n46630 & n46828;
  assign n46830 = ~n46826 & n46827;
  assign n46831 = pi211 & ~n60933;
  assign n46832 = ~n46823 & n46831;
  assign n46833 = ~pi1153 & ~n46215;
  assign n46834 = ~n46182 & ~n46833;
  assign n46835 = ~pi1154 & n46834;
  assign n46836 = pi1153 & pi1154;
  assign n46837 = ~n46835 & ~n46836;
  assign n46838 = pi1153 & ~n46245;
  assign n46839 = ~pi1155 & ~n46838;
  assign n46840 = ~n46837 & n46839;
  assign n46841 = pi1153 & n46194;
  assign n46842 = ~n46221 & ~n46841;
  assign n46843 = pi1155 & ~n46842;
  assign n46844 = pi1153 & ~pi1155;
  assign n46845 = pi1154 & ~n46844;
  assign n46846 = n46632 & n46845;
  assign n46847 = ~n46843 & ~n46846;
  assign n46848 = ~n46840 & n46847;
  assign n46849 = ~pi1153 & ~n46632;
  assign n46850 = n46839 & ~n46849;
  assign n46851 = pi1154 & ~n46653;
  assign n46852 = ~n46850 & n46851;
  assign n46853 = ~n46843 & n46851;
  assign n46854 = ~n46850 & n46853;
  assign n46855 = ~n46843 & n46852;
  assign n46856 = n46834 & n46839;
  assign n46857 = ~pi1154 & ~n46843;
  assign n46858 = ~n46856 & n46857;
  assign n46859 = ~pi211 & ~n46858;
  assign n46860 = ~n60934 & n46859;
  assign n46861 = ~pi211 & ~n60934;
  assign n46862 = ~n46858 & n46861;
  assign n46863 = ~pi211 & ~n46848;
  assign n46864 = ~pi267 & ~n60935;
  assign n46865 = ~n46832 & n46864;
  assign n46866 = ~pi1153 & n46258;
  assign n46867 = ~n46220 & ~n46866;
  assign n46868 = ~pi1155 & n46169;
  assign n46869 = ~n46867 & n46868;
  assign n46870 = pi1153 & ~n46203;
  assign n46871 = pi1155 & ~n46870;
  assign n46872 = n46576 & n46871;
  assign n46873 = pi1154 & ~n46872;
  assign n46874 = pi1154 & ~n46869;
  assign n46875 = ~n46872 & n46874;
  assign n46876 = ~n46869 & n46873;
  assign n46877 = ~pi1154 & ~n46813;
  assign n46878 = ~n46181 & n46877;
  assign n46879 = ~pi1155 & ~n46878;
  assign n46880 = ~n46203 & n46877;
  assign n46881 = ~n46879 & n46880;
  assign n46882 = ~n60936 & ~n46881;
  assign n46883 = pi211 & ~n46882;
  assign n46884 = pi1154 & n46867;
  assign n46885 = n46879 & ~n46884;
  assign n46886 = ~pi1153 & n46212;
  assign n46887 = ~n46201 & ~n46886;
  assign n46888 = pi1154 & n46167;
  assign n46889 = pi1155 & ~n46888;
  assign n46890 = ~n46887 & n46889;
  assign n46891 = ~pi211 & ~n46890;
  assign n46892 = ~n46885 & n46891;
  assign n46893 = pi267 & ~n46892;
  assign n46894 = ~n46883 & n46893;
  assign n46895 = ~pi219 & ~n46894;
  assign n46896 = ~n46865 & n46895;
  assign n46897 = ~pi1154 & ~n46314;
  assign n46898 = ~n46826 & n46897;
  assign n46899 = pi1153 & n46192;
  assign n46900 = pi1154 & pi1155;
  assign n46901 = ~n46193 & n46900;
  assign n46902 = ~n46899 & n46901;
  assign n46903 = ~n46898 & ~n46902;
  assign n46904 = pi211 & ~n46903;
  assign n46905 = pi1154 & ~n46175;
  assign n46906 = pi1154 & n46324;
  assign n46907 = n46322 & n46905;
  assign n46908 = ~pi1155 & ~n60937;
  assign n46909 = n46828 & ~n60937;
  assign n46910 = ~n46826 & n46908;
  assign n46911 = pi1154 & n46664;
  assign n46912 = n46444 & ~n46666;
  assign n46913 = ~n46841 & n46912;
  assign n46914 = ~n46911 & n46913;
  assign n46915 = ~n60938 & ~n46914;
  assign n46916 = ~n46904 & n46915;
  assign n46917 = ~pi267 & ~n46916;
  assign n46918 = pi1154 & ~n46815;
  assign n46919 = ~pi1153 & ~n46560;
  assign n46920 = ~pi1154 & ~n46333;
  assign n46921 = ~n46919 & n46920;
  assign n46922 = ~pi1155 & ~n46921;
  assign n46923 = ~n46918 & n46922;
  assign n46924 = ~pi211 & ~n46159;
  assign n46925 = ~pi211 & n46168;
  assign n46926 = pi299 & n46924;
  assign n46927 = n46590 & ~n60939;
  assign n46928 = ~n46167 & n46212;
  assign n46929 = n46927 & n46928;
  assign n46930 = ~n46292 & ~n46929;
  assign n46931 = n46167 & ~n46609;
  assign n46932 = n46871 & ~n46931;
  assign n46933 = ~n46930 & n46932;
  assign n46934 = ~n46923 & ~n46933;
  assign n46935 = pi267 & ~n46934;
  assign n46936 = pi219 & ~n46935;
  assign n46937 = ~pi267 & ~n60938;
  assign n46938 = ~n46914 & n46937;
  assign n46939 = ~n46904 & n46938;
  assign n46940 = pi267 & ~n46933;
  assign n46941 = ~n46923 & n46940;
  assign n46942 = ~n46939 & ~n46941;
  assign n46943 = pi219 & ~n46942;
  assign n46944 = ~n46917 & n46936;
  assign n46945 = ~n46896 & ~n60940;
  assign n46946 = n46276 & ~n46945;
  assign n46947 = pi1153 & ~n60909;
  assign n46948 = pi1155 & ~n46947;
  assign n46949 = n46701 & n46948;
  assign n46950 = ~pi1153 & ~n46374;
  assign n46951 = pi1153 & ~n46355;
  assign n46952 = ~pi1155 & ~n46951;
  assign n46953 = ~n46950 & n46952;
  assign n46954 = pi1154 & ~n46953;
  assign n46955 = ~n46949 & n46954;
  assign n46956 = ~pi1153 & ~n46361;
  assign n46957 = n46948 & ~n46956;
  assign n46958 = pi1153 & ~n36720;
  assign n46959 = ~pi1155 & ~n46958;
  assign n46960 = pi1091 & n46959;
  assign n46961 = ~pi1154 & ~n46960;
  assign n46962 = ~n46957 & n46961;
  assign n46963 = ~n46955 & ~n46962;
  assign n46964 = ~n46949 & ~n46953;
  assign n46965 = pi1154 & ~n46964;
  assign n46966 = ~n46957 & ~n46960;
  assign n46967 = ~pi1154 & ~n46966;
  assign n46968 = ~pi219 & ~n46967;
  assign n46969 = ~n46965 & n46968;
  assign n46970 = ~pi219 & ~n46965;
  assign n46971 = ~n46967 & n46970;
  assign n46972 = ~pi219 & ~n46963;
  assign n46973 = ~pi1153 & ~n46386;
  assign n46974 = pi1091 & n46699;
  assign n46975 = ~n46973 & n46974;
  assign n46976 = pi1154 & ~n46975;
  assign n46977 = ~pi200 & ~pi1153;
  assign n46978 = ~pi199 & ~n46977;
  assign n46979 = ~pi299 & n46978;
  assign n46980 = pi1091 & ~n46979;
  assign n46981 = n46976 & n46980;
  assign n46982 = pi1153 & ~n46365;
  assign n46983 = ~pi1153 & ~n46422;
  assign n46984 = ~n46982 & ~n46983;
  assign n46985 = pi1155 & ~n46984;
  assign n46986 = pi1153 & n45444;
  assign n46987 = ~pi1154 & ~n46986;
  assign n46988 = pi1091 & n46987;
  assign n46989 = n46713 & ~n46986;
  assign n46990 = ~n46985 & n60942;
  assign n46991 = pi219 & ~n46990;
  assign n46992 = ~n46981 & n46991;
  assign n46993 = ~n60941 & ~n46992;
  assign n46994 = ~pi211 & ~n46993;
  assign n46995 = ~pi299 & ~n46978;
  assign n46996 = ~pi1155 & ~n46995;
  assign n46997 = ~n46737 & ~n46996;
  assign n46998 = ~n45448 & ~n46997;
  assign n46999 = ~pi299 & ~n46348;
  assign n47000 = ~pi1153 & n36719;
  assign n47001 = n46999 & ~n47000;
  assign n47002 = pi1155 & n47001;
  assign n47003 = pi1154 & ~n47002;
  assign n47004 = pi1091 & n47003;
  assign n47005 = ~n46998 & n47004;
  assign n47006 = n46360 & ~n46738;
  assign n47007 = ~n46361 & ~n46738;
  assign n47008 = n60942 & ~n47007;
  assign n47009 = n60942 & ~n47006;
  assign n47010 = pi211 & ~n60943;
  assign n47011 = ~n47005 & n47010;
  assign n47012 = ~n46994 & ~n47011;
  assign n47013 = pi267 & ~n47012;
  assign n47014 = ~pi1153 & ~n36720;
  assign n47015 = ~pi200 & pi1155;
  assign n47016 = n45521 & ~n47015;
  assign n47017 = ~pi1154 & n46365;
  assign n47018 = ~n47016 & ~n47017;
  assign n47019 = ~n47014 & n47018;
  assign n47020 = pi1091 & n47019;
  assign n47021 = ~pi211 & ~n47020;
  assign n47022 = pi211 & pi1154;
  assign n47023 = pi1091 & ~pi1155;
  assign n47024 = ~n46995 & n47023;
  assign n47025 = n47022 & ~n47024;
  assign n47026 = ~n46975 & n47025;
  assign n47027 = ~pi219 & ~n47026;
  assign n47028 = ~pi219 & ~n47021;
  assign n47029 = ~n47026 & n47028;
  assign n47030 = ~n47021 & n47027;
  assign n47031 = n46979 & n47023;
  assign n47032 = n46976 & ~n47031;
  assign n47033 = pi1154 & ~n47032;
  assign n47034 = n46713 & ~n46738;
  assign n47035 = ~n46984 & n47034;
  assign n47036 = ~pi211 & ~n47035;
  assign n47037 = ~n47033 & n47036;
  assign n47038 = n46699 & n47003;
  assign n47039 = ~n47032 & ~n47038;
  assign n47040 = pi211 & ~n47039;
  assign n47041 = pi219 & ~n47040;
  assign n47042 = pi219 & ~n47037;
  assign n47043 = ~n47040 & n47042;
  assign n47044 = ~n47037 & n47041;
  assign n47045 = ~n60944 & ~n60945;
  assign n47046 = pi1091 & ~pi1153;
  assign n47047 = n46360 & n47046;
  assign n47048 = pi1091 & pi1153;
  assign n47049 = n46389 & n47048;
  assign n47050 = ~n47047 & ~n47049;
  assign n47051 = ~n46959 & ~n47050;
  assign n47052 = pi211 & ~pi1154;
  assign n47053 = ~n47051 & n47052;
  assign n47054 = ~pi267 & ~n47053;
  assign n47055 = ~n47045 & n47054;
  assign n47056 = ~n47013 & ~n47055;
  assign n47057 = ~n46276 & ~n47056;
  assign n47058 = n58992 & ~n47057;
  assign n47059 = ~n46946 & n47058;
  assign n47060 = ~pi219 & n46159;
  assign n47061 = ~n46780 & ~n47060;
  assign n47062 = pi267 & n47061;
  assign n47063 = ~pi267 & ~n46161;
  assign n47064 = ~n46791 & n47063;
  assign n47065 = n46276 & ~n47064;
  assign n47066 = ~n47062 & n47065;
  assign n47067 = pi219 & ~n46444;
  assign n47068 = ~pi211 & pi1153;
  assign n47069 = ~pi219 & ~n47022;
  assign n47070 = ~n47068 & n47069;
  assign n47071 = ~n47067 & ~n47070;
  assign n47072 = pi1091 & ~n47071;
  assign n47073 = ~pi267 & ~pi1091;
  assign n47074 = ~n46276 & n47073;
  assign n47075 = ~n47072 & ~n47074;
  assign n47076 = ~n47066 & n47075;
  assign n47077 = ~n58992 & ~n47076;
  assign n47078 = n46440 & ~n47077;
  assign n47079 = ~n47059 & n47078;
  assign n47080 = n58992 & n47056;
  assign n47081 = ~n47072 & ~n47073;
  assign n47082 = ~n58992 & ~n47081;
  assign n47083 = ~n46440 & ~n47082;
  assign n47084 = ~n47080 & n47083;
  assign n47085 = ~pi230 & ~n47084;
  assign n47086 = ~n47079 & n47085;
  assign n47087 = ~pi199 & ~pi1153;
  assign n47088 = n46389 & ~n47087;
  assign n47089 = pi1155 & n47088;
  assign n47090 = ~n46987 & ~n46995;
  assign n47091 = ~pi1155 & n46986;
  assign n47092 = ~pi1154 & ~n47091;
  assign n47093 = ~n46995 & ~n47092;
  assign n47094 = ~n47089 & ~n47093;
  assign n47095 = ~n47089 & ~n47090;
  assign n47096 = pi219 & ~n47001;
  assign n47097 = pi211 & ~n47096;
  assign n47098 = ~n60946 & n47097;
  assign n47099 = ~pi219 & ~n47019;
  assign n47100 = pi200 & ~n46510;
  assign n47101 = ~pi1155 & ~n45518;
  assign n47102 = ~n47000 & ~n47101;
  assign n47103 = ~n47100 & n47102;
  assign n47104 = pi219 & ~n46506;
  assign n47105 = ~n47103 & n47104;
  assign n47106 = ~pi211 & ~n47105;
  assign n47107 = ~n47099 & n47106;
  assign n47108 = ~n47098 & ~n47107;
  assign n47109 = ~n60946 & ~n47096;
  assign n47110 = pi211 & ~n47109;
  assign n47111 = ~n46506 & ~n47103;
  assign n47112 = pi219 & ~n47111;
  assign n47113 = ~pi219 & n47019;
  assign n47114 = ~pi211 & ~n47113;
  assign n47115 = ~n47112 & n47114;
  assign n47116 = n58992 & ~n47115;
  assign n47117 = ~n47110 & n47116;
  assign n47118 = n58992 & ~n47108;
  assign n47119 = ~n58992 & n47071;
  assign n47120 = pi230 & ~n47119;
  assign n47121 = ~n60947 & n47120;
  assign po424 = ~n47086 & ~n47121;
  assign n47123 = pi1153 & ~pi1154;
  assign n47124 = ~n46705 & n47123;
  assign n47125 = ~pi1153 & ~n46389;
  assign n47126 = ~n46736 & ~n47125;
  assign n47127 = pi1154 & n47126;
  assign n47128 = ~n47124 & ~n47127;
  assign n47129 = n45426 & ~n47128;
  assign n47130 = ~pi199 & pi1153;
  assign n47131 = pi200 & n47130;
  assign n47132 = pi1153 & n45424;
  assign n47133 = ~pi299 & n60948;
  assign n47134 = ~pi1154 & ~n47133;
  assign n47135 = pi299 & n36681;
  assign n47136 = n46499 & ~n47087;
  assign n47137 = ~n45426 & n47136;
  assign n47138 = ~n47135 & ~n47137;
  assign n47139 = ~n47134 & ~n47138;
  assign n47140 = ~n47129 & ~n47139;
  assign n47141 = n58992 & ~n47140;
  assign n47142 = pi219 & ~n46552;
  assign n47143 = pi211 & pi1153;
  assign n47144 = ~pi219 & ~n47143;
  assign n47145 = ~n47142 & ~n47144;
  assign n47146 = ~n58992 & n47145;
  assign n47147 = ~pi1152 & ~n47146;
  assign n47148 = ~n47141 & n47147;
  assign n47149 = ~n45445 & ~n46389;
  assign n47150 = pi1154 & ~n47149;
  assign n47151 = pi200 & ~pi1153;
  assign n47152 = n45518 & ~n47151;
  assign n47153 = pi219 & ~n47152;
  assign n47154 = pi1153 & ~n46999;
  assign n47155 = ~n47125 & ~n47154;
  assign n47156 = n47022 & ~n47155;
  assign n47157 = pi1154 & n46365;
  assign n47158 = ~n47130 & n47157;
  assign n47159 = ~pi1154 & ~n47152;
  assign n47160 = ~n47158 & ~n47159;
  assign n47161 = ~n47156 & n47160;
  assign n47162 = pi219 & ~n47161;
  assign n47163 = ~n47150 & n47153;
  assign n47164 = ~pi200 & pi1154;
  assign n47165 = n45521 & ~n47164;
  assign n47166 = ~n45445 & n47125;
  assign n47167 = ~n47165 & ~n47166;
  assign n47168 = ~pi219 & ~n47167;
  assign n47169 = n58992 & ~n47168;
  assign n47170 = ~n60949 & n47169;
  assign n47171 = ~n58992 & ~n47142;
  assign n47172 = n45426 & ~n47143;
  assign n47173 = n47171 & ~n47172;
  assign n47174 = pi1152 & ~n47173;
  assign n47175 = ~n47170 & n47174;
  assign n47176 = ~n47148 & ~n47175;
  assign n47177 = pi230 & ~n47176;
  assign n47178 = ~n46172 & ~n46176;
  assign n47179 = ~pi1153 & ~n47178;
  assign n47180 = ~n46183 & n46927;
  assign n47181 = ~n47179 & n47180;
  assign n47182 = ~pi1153 & n47181;
  assign n47183 = ~n46220 & ~n47182;
  assign n47184 = ~pi1154 & ~n47183;
  assign n47185 = pi1153 & ~n60904;
  assign n47186 = n46905 & n46927;
  assign n47187 = ~n47185 & n47186;
  assign n47188 = pi254 & ~n47187;
  assign n47189 = ~n47184 & n47188;
  assign n47190 = ~n46245 & ~n46911;
  assign n47191 = pi211 & n46168;
  assign n47192 = ~n46182 & ~n47191;
  assign n47193 = ~pi1153 & ~n47192;
  assign n47194 = ~pi254 & ~n47193;
  assign n47195 = ~n47190 & n47194;
  assign n47196 = ~n47189 & ~n47195;
  assign n47197 = ~pi219 & ~n47196;
  assign n47198 = ~n46281 & ~n46929;
  assign n47199 = pi1153 & ~n46929;
  assign n47200 = pi1154 & ~n47199;
  assign n47201 = ~n47198 & n47200;
  assign n47202 = pi1153 & ~n46327;
  assign n47203 = ~pi1153 & ~n46333;
  assign n47204 = ~pi1154 & ~n47203;
  assign n47205 = ~n47202 & n47204;
  assign n47206 = pi254 & ~n47205;
  assign n47207 = ~n47201 & n47206;
  assign n47208 = n46324 & ~n46824;
  assign n47209 = ~pi1154 & ~n47208;
  assign n47210 = ~n46825 & n47209;
  assign n47211 = ~pi1153 & ~n46327;
  assign n47212 = n46664 & ~n47211;
  assign n47213 = n46552 & ~n47212;
  assign n47214 = ~n46151 & n47213;
  assign n47215 = ~n46310 & n47022;
  assign n47216 = ~n46899 & n47215;
  assign n47217 = ~pi254 & ~n47216;
  assign n47218 = ~n47214 & n47217;
  assign n47219 = ~n47210 & n47218;
  assign n47220 = ~n47207 & ~n47219;
  assign n47221 = pi219 & ~n47220;
  assign n47222 = pi253 & ~n47221;
  assign n47223 = ~n47197 & n47222;
  assign n47224 = pi219 & pi1091;
  assign n47225 = ~n46784 & ~n47224;
  assign n47226 = ~n47161 & ~n47225;
  assign n47227 = ~pi211 & n47014;
  assign n47228 = ~pi1154 & ~n46951;
  assign n47229 = ~n46973 & n47228;
  assign n47230 = ~n47227 & n47229;
  assign n47231 = pi1153 & ~n45521;
  assign n47232 = pi1091 & n47022;
  assign n47233 = ~n46389 & n47232;
  assign n47234 = ~n47231 & n47233;
  assign n47235 = ~n47230 & ~n47234;
  assign n47236 = ~pi219 & ~n47235;
  assign n47237 = ~n47226 & ~n47236;
  assign n47238 = pi254 & ~n47237;
  assign n47239 = ~pi254 & ~pi1091;
  assign n47240 = ~n60949 & ~n47168;
  assign n47241 = ~pi254 & ~n47240;
  assign n47242 = ~n47239 & ~n47241;
  assign n47243 = ~n47238 & n47242;
  assign n47244 = ~pi253 & ~n47243;
  assign n47245 = n58992 & ~n47244;
  assign n47246 = ~n47223 & n47245;
  assign n47247 = ~pi219 & n46717;
  assign n47248 = ~pi219 & ~n46161;
  assign n47249 = ~n46924 & n47248;
  assign n47250 = ~pi219 & ~n47249;
  assign n47251 = ~n58992 & n47250;
  assign n47252 = ~n46150 & n47251;
  assign n47253 = ~n58992 & n47247;
  assign n47254 = pi1091 & ~n47145;
  assign n47255 = ~n58992 & ~n47239;
  assign n47256 = ~n47239 & ~n47254;
  assign n47257 = ~n58992 & n47256;
  assign n47258 = ~n47254 & n47255;
  assign n47259 = pi253 & ~n58992;
  assign n47260 = ~pi253 & ~n47256;
  assign n47261 = ~n58992 & ~n47260;
  assign n47262 = ~n60951 & ~n47259;
  assign n47263 = ~n60950 & ~n60951;
  assign n47264 = ~n47259 & n47263;
  assign n47265 = ~n60950 & ~n60952;
  assign n47266 = pi1091 & n47142;
  assign n47267 = n45426 & n47046;
  assign n47268 = pi254 & ~n47267;
  assign n47269 = ~n47266 & n47268;
  assign n47270 = n47061 & n47269;
  assign n47271 = n46783 & ~n46788;
  assign n47272 = ~n47048 & n47271;
  assign n47273 = ~pi254 & ~n47266;
  assign n47274 = ~n46791 & n47273;
  assign n47275 = ~n47272 & n47274;
  assign n47276 = pi253 & ~n47275;
  assign n47277 = pi253 & ~n47270;
  assign n47278 = ~n47275 & n47277;
  assign n47279 = ~n47270 & n47276;
  assign n47280 = ~n60953 & ~n60954;
  assign n47281 = pi1152 & ~n47280;
  assign n47282 = ~n47246 & n47281;
  assign n47283 = ~pi211 & n46666;
  assign n47284 = ~n46169 & ~n47283;
  assign n47285 = ~n46886 & n47284;
  assign n47286 = ~pi219 & ~n46645;
  assign n47287 = ~n47285 & n47286;
  assign n47288 = ~pi1154 & ~n46897;
  assign n47289 = ~pi1154 & n46314;
  assign n47290 = ~n46886 & ~n46928;
  assign n47291 = ~n60955 & n47290;
  assign n47292 = ~n46292 & n46552;
  assign n47293 = pi219 & ~n47292;
  assign n47294 = ~n47291 & n47293;
  assign n47295 = ~n47287 & ~n47294;
  assign n47296 = pi254 & ~n47295;
  assign n47297 = n46193 & ~n47211;
  assign n47298 = n47022 & ~n47297;
  assign n47299 = pi219 & ~n47213;
  assign n47300 = ~n47209 & n47299;
  assign n47301 = ~n47298 & n47300;
  assign n47302 = n46630 & ~n46833;
  assign n47303 = pi1154 & n46221;
  assign n47304 = ~n47302 & ~n47303;
  assign n47305 = ~n46168 & ~n46676;
  assign n47306 = ~pi211 & ~n47305;
  assign n47307 = ~pi219 & ~n47306;
  assign n47308 = pi1154 & ~n46221;
  assign n47309 = ~n47302 & n47308;
  assign n47310 = ~pi1154 & ~n47302;
  assign n47311 = n47307 & ~n47310;
  assign n47312 = ~n47309 & n47311;
  assign n47313 = ~n47304 & n47307;
  assign n47314 = ~pi254 & ~n60956;
  assign n47315 = ~n47301 & n47314;
  assign n47316 = ~n47296 & ~n47315;
  assign n47317 = pi253 & ~n47316;
  assign n47318 = pi1153 & ~n46736;
  assign n47319 = pi1091 & n47318;
  assign n47320 = ~n47047 & ~n47319;
  assign n47321 = pi211 & ~n47228;
  assign n47322 = ~n47320 & n47321;
  assign n47323 = pi1091 & n47136;
  assign n47324 = pi1154 & ~n47323;
  assign n47325 = pi1091 & n47133;
  assign n47326 = n45425 & n47048;
  assign n47327 = ~pi1154 & ~n60957;
  assign n47328 = ~pi211 & ~n47327;
  assign n47329 = ~n47324 & n47328;
  assign n47330 = ~n47322 & ~n47329;
  assign n47331 = ~pi219 & ~n47330;
  assign n47332 = pi211 & n47324;
  assign n47333 = pi1091 & n46983;
  assign n47334 = n46552 & ~n47333;
  assign n47335 = ~n47319 & n47334;
  assign n47336 = pi219 & ~n47327;
  assign n47337 = ~n47335 & n47336;
  assign n47338 = ~n47332 & n47337;
  assign n47339 = ~n47331 & ~n47338;
  assign n47340 = ~pi254 & ~n47339;
  assign n47341 = pi1091 & ~n45426;
  assign n47342 = ~n47133 & n47341;
  assign n47343 = ~pi1154 & ~n47342;
  assign n47344 = ~n36681 & ~n45426;
  assign n47345 = n46351 & ~n46498;
  assign n47346 = pi1153 & ~n47345;
  assign n47347 = ~n46956 & ~n47346;
  assign n47348 = ~n46701 & ~n47347;
  assign n47349 = n47344 & ~n47348;
  assign n47350 = n36681 & ~n47346;
  assign n47351 = n46423 & n47350;
  assign n47352 = pi1154 & ~n47351;
  assign n47353 = ~n47349 & n47352;
  assign n47354 = ~n47343 & ~n47353;
  assign n47355 = ~pi1154 & n46397;
  assign n47356 = n46705 & n46713;
  assign n47357 = ~n47347 & ~n60958;
  assign n47358 = n45426 & ~n47357;
  assign n47359 = pi254 & ~n47358;
  assign n47360 = ~n47354 & n47359;
  assign n47361 = ~n47340 & ~n47360;
  assign n47362 = ~pi253 & n47361;
  assign n47363 = n58992 & ~n47362;
  assign n47364 = ~n47317 & n47363;
  assign n47365 = ~n47250 & n47275;
  assign n47366 = n47248 & ~n47271;
  assign n47367 = n47270 & ~n47366;
  assign n47368 = pi253 & ~n47367;
  assign n47369 = pi253 & ~n47365;
  assign n47370 = ~n47367 & n47369;
  assign n47371 = ~n47365 & n47368;
  assign n47372 = n60952 & ~n60959;
  assign n47373 = ~pi1152 & ~n47372;
  assign n47374 = ~n47364 & n47373;
  assign n47375 = n46440 & ~n47374;
  assign n47376 = ~n47282 & n47375;
  assign n47377 = n58992 & ~n47361;
  assign n47378 = ~pi1152 & ~n60951;
  assign n47379 = ~n47377 & n47378;
  assign n47380 = n58992 & n47243;
  assign n47381 = pi1152 & ~n60950;
  assign n47382 = pi1152 & n47263;
  assign n47383 = ~n60951 & n47381;
  assign n47384 = ~n47380 & n60960;
  assign n47385 = ~n46440 & ~n47384;
  assign n47386 = ~n47379 & n47385;
  assign n47387 = ~pi230 & ~n47386;
  assign n47388 = ~n47376 & n47387;
  assign po411 = ~n47177 & ~n47388;
  assign n47390 = ~pi230 & pi587;
  assign n47391 = pi230 & n6701;
  assign n47392 = ~n59346 & n47391;
  assign n47393 = ~n25407 & n47392;
  assign n47394 = n59348 & n47393;
  assign n47395 = n12602 & n47394;
  assign n47396 = ~n47390 & ~n47395;
  assign n47397 = ~pi230 & pi602;
  assign n47398 = pi790 & ~n23532;
  assign n47399 = pi790 & ~n23534;
  assign n47400 = ~n23532 & n47399;
  assign n47401 = ~n23534 & n47398;
  assign n47402 = ~n59304 & ~n9743;
  assign n47403 = ~n60961 & n47402;
  assign n47404 = pi230 & n7054;
  assign n47405 = ~n59240 & n47404;
  assign n47406 = n9554 & n47405;
  assign n47407 = n9651 & n47405;
  assign n47408 = n9554 & n47407;
  assign n47409 = n9651 & n47406;
  assign n47410 = n47403 & n47405;
  assign n47411 = n9652 & n47410;
  assign n47412 = n47403 & n60962;
  assign n47413 = ~n47397 & ~n60963;
  assign n47414 = ~pi219 & pi299;
  assign n47415 = ~n45447 & ~n47414;
  assign n47416 = ~n46422 & n47415;
  assign n47417 = n58992 & n47416;
  assign n47418 = pi219 & n45884;
  assign n47419 = ~n47417 & ~n47418;
  assign n47420 = ~pi1151 & pi1153;
  assign n47421 = ~n47419 & n47420;
  assign n47422 = ~n46982 & ~n47014;
  assign n47423 = n36679 & n47422;
  assign n47424 = pi199 & ~pi1153;
  assign n47425 = n46389 & ~n47424;
  assign n47426 = pi211 & ~n47425;
  assign n47427 = ~n47423 & ~n47426;
  assign n47428 = pi1151 & n58992;
  assign n47429 = ~pi1153 & ~n45518;
  assign n47430 = ~n46365 & ~n47429;
  assign n47431 = n36681 & ~n47430;
  assign n47432 = n47428 & ~n47431;
  assign n47433 = n47427 & n47432;
  assign n47434 = ~n47421 & ~n47433;
  assign n47435 = ~pi1152 & ~n47434;
  assign n47436 = pi219 & ~n47068;
  assign n47437 = ~pi219 & ~n58992;
  assign n47438 = pi1153 & n45884;
  assign n47439 = ~n47437 & ~n47438;
  assign n47440 = ~n58992 & ~n47436;
  assign n47441 = pi1152 & ~n36679;
  assign n47442 = pi1151 & ~n45426;
  assign n47443 = ~n47441 & ~n47442;
  assign n47444 = ~n60964 & ~n47443;
  assign n47445 = n36681 & n47318;
  assign n47446 = n46499 & ~n47424;
  assign n47447 = ~pi1151 & ~n45427;
  assign n47448 = ~n47446 & n47447;
  assign n47449 = ~n47445 & n47448;
  assign n47450 = pi1152 & n58992;
  assign n47451 = pi1153 & ~n47149;
  assign n47452 = ~n45518 & ~n47414;
  assign n47453 = pi1151 & n47452;
  assign n47454 = ~n47451 & n47453;
  assign n47455 = n47450 & ~n47454;
  assign n47456 = ~n47449 & n47455;
  assign n47457 = pi230 & ~n47456;
  assign n47458 = ~n47444 & n47457;
  assign n47459 = pi1153 & ~n47419;
  assign n47460 = ~pi1151 & ~n47459;
  assign n47461 = n58992 & ~n47431;
  assign n47462 = n47427 & n47461;
  assign n47463 = ~n45426 & ~n60964;
  assign n47464 = pi1151 & ~n47463;
  assign n47465 = pi1151 & ~n47462;
  assign n47466 = ~n47463 & n47465;
  assign n47467 = ~n47462 & n47464;
  assign n47468 = ~n47460 & ~n60965;
  assign n47469 = ~pi1152 & ~n47468;
  assign n47470 = n58992 & ~n47454;
  assign n47471 = ~n47449 & n47470;
  assign n47472 = ~pi1151 & n36679;
  assign n47473 = ~n47436 & ~n47472;
  assign n47474 = ~n60964 & ~n47472;
  assign n47475 = ~n58992 & n47473;
  assign n47476 = pi1152 & ~n60966;
  assign n47477 = pi1152 & ~n47471;
  assign n47478 = ~n60966 & n47477;
  assign n47479 = ~n47471 & n47476;
  assign n47480 = ~n47469 & ~n60967;
  assign n47481 = pi230 & ~n47480;
  assign n47482 = ~n47435 & n47458;
  assign n47483 = pi219 & ~n47211;
  assign n47484 = ~n47199 & n47483;
  assign n47485 = ~pi219 & ~n46819;
  assign n47486 = ~n47185 & n47485;
  assign n47487 = pi253 & ~n47486;
  assign n47488 = ~n47484 & n47487;
  assign n47489 = ~n46192 & ~n47283;
  assign n47490 = pi1153 & ~n47489;
  assign n47491 = ~n46322 & ~n47490;
  assign n47492 = pi219 & n47491;
  assign n47493 = pi1153 & n46198;
  assign n47494 = ~pi219 & ~n46813;
  assign n47495 = ~n47493 & n47494;
  assign n47496 = ~pi253 & ~n47495;
  assign n47497 = ~n47492 & n47496;
  assign n47498 = ~n47488 & ~n47497;
  assign n47499 = n58992 & ~n47498;
  assign n47500 = pi253 & ~n46190;
  assign n47501 = ~n47248 & n47500;
  assign n47502 = ~pi253 & ~n46783;
  assign n47503 = ~n46791 & n47502;
  assign n47504 = ~n47501 & ~n47503;
  assign n47505 = ~n47068 & n47224;
  assign n47506 = ~n58992 & ~n47505;
  assign n47507 = ~n46783 & ~n47505;
  assign n47508 = ~n46791 & n47507;
  assign n47509 = ~pi253 & ~n47508;
  assign n47510 = ~n46190 & ~n47505;
  assign n47511 = ~n47248 & n47510;
  assign n47512 = pi253 & ~n47511;
  assign n47513 = ~n58992 & ~n47512;
  assign n47514 = ~n47509 & n47513;
  assign n47515 = ~n47504 & n47506;
  assign n47516 = pi1151 & ~n60950;
  assign n47517 = pi1151 & ~n60969;
  assign n47518 = ~n60950 & n47517;
  assign n47519 = ~n60969 & n47516;
  assign n47520 = ~n47499 & n60970;
  assign n47521 = ~pi219 & ~n47181;
  assign n47522 = pi219 & n46180;
  assign n47523 = ~n47521 & ~n47522;
  assign n47524 = ~n47492 & n47523;
  assign n47525 = ~pi253 & ~n47524;
  assign n47526 = n47248 & ~n47284;
  assign n47527 = ~n46177 & ~n47179;
  assign n47528 = n47526 & ~n47527;
  assign n47529 = pi219 & n46279;
  assign n47530 = ~n46292 & n47199;
  assign n47531 = n47529 & ~n47530;
  assign n47532 = ~n47528 & ~n47531;
  assign n47533 = pi253 & ~n47532;
  assign n47534 = n58992 & ~n47533;
  assign n47535 = ~n47525 & n47534;
  assign n47536 = ~pi1151 & ~n47535;
  assign n47537 = ~n47520 & ~n47536;
  assign n47538 = ~n58992 & ~n46778;
  assign n47539 = ~n47366 & n47538;
  assign n47540 = ~n46150 & n47539;
  assign n47541 = ~n60969 & ~n47540;
  assign n47542 = ~n47537 & n47541;
  assign n47543 = pi1152 & ~n47542;
  assign n47544 = pi219 & ~n47491;
  assign n47545 = ~n47495 & n47526;
  assign n47546 = ~n47544 & ~n47545;
  assign n47547 = ~n46182 & ~n47546;
  assign n47548 = ~pi253 & ~n47547;
  assign n47549 = n46927 & n47248;
  assign n47550 = ~n46870 & n47549;
  assign n47551 = pi1153 & n47198;
  assign n47552 = pi219 & ~n47203;
  assign n47553 = ~n47551 & n47552;
  assign n47554 = ~n47550 & ~n47553;
  assign n47555 = pi253 & ~n47554;
  assign n47556 = n58992 & ~n47555;
  assign n47557 = ~n47548 & n47556;
  assign n47558 = n60970 & ~n47557;
  assign n47559 = ~n46166 & n47544;
  assign n47560 = ~pi219 & n46220;
  assign n47561 = n46834 & n47560;
  assign n47562 = ~pi253 & ~n47561;
  assign n47563 = ~n47559 & n47562;
  assign n47564 = ~pi219 & n47178;
  assign n47565 = ~n46919 & ~n47564;
  assign n47566 = n46930 & n47565;
  assign n47567 = pi253 & ~n47566;
  assign n47568 = n58992 & ~n47567;
  assign n47569 = ~n47563 & n47568;
  assign n47570 = ~pi1151 & ~n60969;
  assign n47571 = ~n47569 & n47570;
  assign n47572 = ~pi1152 & ~n47571;
  assign n47573 = ~n47558 & n47572;
  assign n47574 = ~n47543 & ~n47573;
  assign n47575 = n46440 & ~n47574;
  assign n47576 = ~pi253 & ~pi1091;
  assign n47577 = ~n58992 & ~n47576;
  assign n47578 = ~n47505 & n47577;
  assign n47579 = pi219 & n47578;
  assign n47580 = n47048 & n47417;
  assign n47581 = pi253 & ~pi1091;
  assign n47582 = ~pi1151 & ~n47581;
  assign n47583 = ~n47580 & n47582;
  assign n47584 = ~n47579 & n47583;
  assign n47585 = pi1091 & ~n47427;
  assign n47586 = n36681 & ~n46947;
  assign n47587 = ~n46973 & n47586;
  assign n47588 = ~n47585 & ~n47587;
  assign n47589 = pi253 & ~n47588;
  assign n47590 = ~n60847 & ~n47451;
  assign n47591 = pi1091 & ~n47590;
  assign n47592 = ~pi253 & ~n47591;
  assign n47593 = n58992 & ~n47592;
  assign n47594 = ~n47589 & n47593;
  assign n47595 = pi219 & n47046;
  assign n47596 = ~n46707 & ~n47595;
  assign n47597 = n47577 & n47596;
  assign n47598 = pi1151 & ~n47597;
  assign n47599 = ~n47594 & n47598;
  assign n47600 = ~n47584 & ~n47599;
  assign n47601 = ~pi1152 & ~n47600;
  assign n47602 = ~n46950 & n47350;
  assign n47603 = n45426 & n46351;
  assign n47604 = ~n47446 & n47603;
  assign n47605 = pi253 & ~n47604;
  assign n47606 = ~n47602 & n47605;
  assign n47607 = pi1091 & n47446;
  assign n47608 = pi211 & ~n46416;
  assign n47609 = ~n47607 & n47608;
  assign n47610 = n60909 & n47087;
  assign n47611 = n36681 & ~n47610;
  assign n47612 = ~n47319 & n47611;
  assign n47613 = ~pi253 & ~n47612;
  assign n47614 = ~n47609 & n47613;
  assign n47615 = ~n47606 & ~n47614;
  assign n47616 = ~pi57 & ~pi1151;
  assign n47617 = ~pi1151 & n58992;
  assign n47618 = n4441 & n47616;
  assign n47619 = n47344 & ~n47581;
  assign n47620 = ~n47607 & n47619;
  assign n47621 = n60971 & ~n47620;
  assign n47622 = ~n47615 & n47621;
  assign n47623 = ~pi1151 & n47247;
  assign n47624 = n47578 & ~n47623;
  assign n47625 = n47149 & ~n47581;
  assign n47626 = ~n47046 & ~n47625;
  assign n47627 = n47452 & ~n47626;
  assign n47628 = n47428 & ~n47576;
  assign n47629 = ~n47627 & n47628;
  assign n47630 = pi1152 & ~n47629;
  assign n47631 = n58992 & ~n47576;
  assign n47632 = ~n47627 & n47631;
  assign n47633 = ~n47578 & ~n47632;
  assign n47634 = pi1151 & ~n47633;
  assign n47635 = ~n47247 & n47578;
  assign n47636 = pi1152 & ~n47635;
  assign n47637 = ~n47634 & n47636;
  assign n47638 = ~n47624 & n47630;
  assign n47639 = ~n47622 & n60972;
  assign n47640 = ~n46440 & ~n47639;
  assign n47641 = ~n47601 & n47640;
  assign n47642 = ~pi230 & ~n47641;
  assign n47643 = ~n47575 & n47642;
  assign po410 = ~n60968 & ~n47643;
  assign n47645 = ~pi1137 & ~pi1138;
  assign n47646 = ~pi1134 & n47645;
  assign n47647 = ~pi680 & pi1135;
  assign n47648 = ~pi603 & ~pi1135;
  assign n47649 = pi1136 & ~n47648;
  assign n47650 = pi1136 & ~n47647;
  assign n47651 = ~n47648 & n47650;
  assign n47652 = ~n47647 & n47649;
  assign n47653 = ~pi778 & pi1135;
  assign n47654 = ~pi981 & ~pi1135;
  assign n47655 = ~pi1136 & ~n47654;
  assign n47656 = ~pi1136 & ~n47653;
  assign n47657 = ~n47654 & n47656;
  assign n47658 = ~n47653 & n47655;
  assign n47659 = ~n60973 & ~n60974;
  assign n47660 = n47646 & ~n47659;
  assign n47661 = pi1135 & n47645;
  assign n47662 = pi1136 & ~n47661;
  assign n47663 = ~pi759 & n47662;
  assign n47664 = pi1135 & ~pi1136;
  assign n47665 = pi1134 & n47645;
  assign n47666 = ~n47664 & n47665;
  assign n47667 = ~pi696 & pi1135;
  assign n47668 = ~pi837 & ~pi1136;
  assign n47669 = ~n47667 & ~n47668;
  assign n47670 = n47666 & n47669;
  assign n47671 = ~n47663 & n47670;
  assign n47672 = ~n47660 & ~n47671;
  assign n47673 = ~n5138 & ~n47672;
  assign n47674 = ~pi590 & pi592;
  assign n47675 = ~pi588 & ~n47674;
  assign n47676 = ~pi590 & pi591;
  assign n47677 = pi390 & n47676;
  assign n47678 = n47675 & ~n47677;
  assign n47679 = pi363 & ~pi591;
  assign n47680 = pi592 & ~n47679;
  assign n47681 = ~n47678 & ~n47680;
  assign n47682 = pi590 & ~pi591;
  assign n47683 = ~pi592 & n47682;
  assign n47684 = pi342 & n47683;
  assign n47685 = ~n47681 & ~n47684;
  assign n47686 = ~pi223 & ~pi224;
  assign n47687 = pi414 & n5089;
  assign n47688 = pi588 & ~n47687;
  assign n47689 = n47686 & ~n47688;
  assign n47690 = ~n47685 & n47689;
  assign n47691 = pi199 & ~pi1049;
  assign n47692 = ~pi199 & ~pi291;
  assign n47693 = ~n47686 & ~n47692;
  assign n47694 = ~n47686 & ~n47691;
  assign n47695 = ~n47692 & n47694;
  assign n47696 = ~n47691 & n47693;
  assign n47697 = ~n47690 & ~n60975;
  assign n47698 = n5138 & ~n47697;
  assign n47699 = ~n47673 & ~n47698;
  assign n47700 = ~pi661 & pi1135;
  assign n47701 = ~pi616 & ~pi1135;
  assign n47702 = pi1136 & ~n47701;
  assign n47703 = pi1136 & ~n47700;
  assign n47704 = ~n47701 & n47703;
  assign n47705 = ~n47700 & n47702;
  assign n47706 = ~pi781 & pi1135;
  assign n47707 = ~pi808 & ~pi1135;
  assign n47708 = ~pi1136 & ~n47707;
  assign n47709 = ~pi1136 & ~n47706;
  assign n47710 = ~n47707 & n47709;
  assign n47711 = ~n47706 & n47708;
  assign n47712 = ~n60976 & ~n60977;
  assign n47713 = n47646 & ~n47712;
  assign n47714 = ~pi758 & n47662;
  assign n47715 = ~pi736 & pi1135;
  assign n47716 = ~pi850 & ~pi1136;
  assign n47717 = ~n47715 & ~n47716;
  assign n47718 = n47666 & n47717;
  assign n47719 = ~n47714 & n47718;
  assign n47720 = ~n47713 & ~n47719;
  assign n47721 = ~n5138 & ~n47720;
  assign n47722 = pi397 & n47676;
  assign n47723 = n47675 & ~n47722;
  assign n47724 = pi372 & ~pi591;
  assign n47725 = pi592 & ~n47724;
  assign n47726 = ~n47723 & ~n47725;
  assign n47727 = pi320 & n47683;
  assign n47728 = ~n47726 & ~n47727;
  assign n47729 = pi422 & n5089;
  assign n47730 = pi588 & ~n47729;
  assign n47731 = n47686 & ~n47730;
  assign n47732 = ~n47728 & n47731;
  assign n47733 = pi199 & ~pi1048;
  assign n47734 = ~pi199 & ~pi290;
  assign n47735 = ~n47686 & ~n47734;
  assign n47736 = ~n47686 & ~n47733;
  assign n47737 = ~n47734 & n47736;
  assign n47738 = ~n47733 & n47735;
  assign n47739 = ~n47732 & ~n60978;
  assign n47740 = n5138 & ~n47739;
  assign n47741 = ~n47721 & ~n47740;
  assign n47742 = ~pi637 & pi1135;
  assign n47743 = ~pi617 & ~pi1135;
  assign n47744 = pi1136 & ~n47743;
  assign n47745 = pi1136 & ~n47742;
  assign n47746 = ~n47743 & n47745;
  assign n47747 = ~n47742 & n47744;
  assign n47748 = pi814 & ~pi1135;
  assign n47749 = ~pi788 & pi1135;
  assign n47750 = ~pi1136 & ~n47749;
  assign n47751 = ~pi1136 & ~n47748;
  assign n47752 = ~n47749 & n47751;
  assign n47753 = ~n47748 & n47750;
  assign n47754 = ~n60979 & ~n60980;
  assign n47755 = n47646 & ~n47754;
  assign n47756 = ~pi749 & n47662;
  assign n47757 = ~pi706 & pi1135;
  assign n47758 = ~pi866 & ~pi1136;
  assign n47759 = ~n47757 & ~n47758;
  assign n47760 = n47666 & n47759;
  assign n47761 = ~n47756 & n47760;
  assign n47762 = ~n47755 & ~n47761;
  assign n47763 = ~n5138 & ~n47762;
  assign n47764 = pi411 & n47676;
  assign n47765 = n47675 & ~n47764;
  assign n47766 = pi387 & ~pi591;
  assign n47767 = pi592 & ~n47766;
  assign n47768 = ~n47765 & ~n47767;
  assign n47769 = pi452 & n47683;
  assign n47770 = ~n47768 & ~n47769;
  assign n47771 = pi435 & n5089;
  assign n47772 = pi588 & ~n47771;
  assign n47773 = n47686 & ~n47772;
  assign n47774 = ~n47770 & n47773;
  assign n47775 = pi199 & ~pi1053;
  assign n47776 = ~pi199 & ~pi295;
  assign n47777 = ~n47686 & ~n47776;
  assign n47778 = ~n47686 & ~n47775;
  assign n47779 = ~n47776 & n47778;
  assign n47780 = ~n47775 & n47777;
  assign n47781 = ~n47774 & ~n60981;
  assign n47782 = n5138 & ~n47781;
  assign n47783 = ~n47763 & ~n47782;
  assign n47784 = pi199 & ~pi1070;
  assign n47785 = ~pi199 & ~pi256;
  assign n47786 = ~n47686 & ~n47785;
  assign n47787 = ~n47686 & ~n47784;
  assign n47788 = ~n47785 & n47787;
  assign n47789 = ~n47784 & n47786;
  assign n47790 = ~pi591 & pi592;
  assign n47791 = pi336 & n47790;
  assign n47792 = pi463 & pi591;
  assign n47793 = ~pi592 & n47792;
  assign n47794 = ~n47791 & ~n47793;
  assign n47795 = ~pi590 & ~n47794;
  assign n47796 = pi362 & n47683;
  assign n47797 = ~pi588 & ~n47796;
  assign n47798 = ~n47795 & n47797;
  assign n47799 = pi437 & n5089;
  assign n47800 = pi588 & ~n47799;
  assign n47801 = n47686 & ~n47800;
  assign n47802 = ~n47798 & n47801;
  assign n47803 = ~n60982 & ~n47802;
  assign n47804 = n5138 & ~n47803;
  assign n47805 = pi639 & pi1135;
  assign n47806 = pi622 & ~pi1135;
  assign n47807 = pi1136 & ~n47806;
  assign n47808 = pi1136 & ~n47805;
  assign n47809 = ~n47806 & n47808;
  assign n47810 = ~n47805 & n47807;
  assign n47811 = pi783 & pi1135;
  assign n47812 = pi804 & ~pi1135;
  assign n47813 = ~pi1136 & ~n47812;
  assign n47814 = ~pi1136 & ~n47811;
  assign n47815 = ~n47812 & n47814;
  assign n47816 = ~n47811 & n47813;
  assign n47817 = ~n60983 & ~n60984;
  assign n47818 = ~pi1134 & ~n47817;
  assign n47819 = ~n5138 & n47645;
  assign n47820 = ~pi735 & pi1135;
  assign n47821 = ~pi743 & ~pi1135;
  assign n47822 = pi1136 & ~n47821;
  assign n47823 = pi1136 & ~n47820;
  assign n47824 = ~n47821 & n47823;
  assign n47825 = ~n47820 & n47822;
  assign n47826 = ~pi1135 & ~pi1136;
  assign n47827 = pi859 & n47826;
  assign n47828 = pi1134 & ~n47827;
  assign n47829 = ~n60985 & n47828;
  assign n47830 = n47819 & ~n47829;
  assign n47831 = ~n47818 & n47830;
  assign n47832 = ~n47804 & ~n47831;
  assign n47833 = pi876 & n47826;
  assign n47834 = ~pi730 & pi1135;
  assign n47835 = ~pi748 & ~pi1135;
  assign n47836 = pi1136 & ~n47835;
  assign n47837 = pi1136 & ~n47834;
  assign n47838 = ~n47835 & n47837;
  assign n47839 = ~n47834 & n47836;
  assign n47840 = ~n47833 & ~n60986;
  assign n47841 = n47665 & ~n47840;
  assign n47842 = ~pi710 & pi1135;
  assign n47843 = pi1136 & ~n47842;
  assign n47844 = ~pi803 & ~pi1135;
  assign n47845 = pi789 & n47664;
  assign n47846 = ~n47844 & ~n47845;
  assign n47847 = pi803 & ~pi1136;
  assign n47848 = ~pi1135 & ~n47847;
  assign n47849 = pi710 & pi1136;
  assign n47850 = ~n47845 & ~n47849;
  assign n47851 = ~n47848 & n47850;
  assign n47852 = ~n47843 & n47846;
  assign n47853 = ~pi623 & n47662;
  assign n47854 = n47646 & ~n47853;
  assign n47855 = ~n60987 & n47854;
  assign n47856 = ~n47841 & ~n47855;
  assign n47857 = ~n5138 & ~n47856;
  assign n47858 = pi199 & ~pi1037;
  assign n47859 = ~pi199 & ~pi296;
  assign n47860 = ~n47686 & ~n47859;
  assign n47861 = ~n47686 & ~n47858;
  assign n47862 = ~n47859 & n47861;
  assign n47863 = ~n47858 & n47860;
  assign n47864 = pi412 & n47676;
  assign n47865 = n47675 & ~n47864;
  assign n47866 = pi388 & ~pi591;
  assign n47867 = pi592 & ~n47866;
  assign n47868 = ~n47865 & ~n47867;
  assign n47869 = pi455 & n47683;
  assign n47870 = ~n47868 & ~n47869;
  assign n47871 = pi436 & n5089;
  assign n47872 = pi588 & ~n47871;
  assign n47873 = n47686 & ~n47872;
  assign n47874 = ~n47870 & n47873;
  assign n47875 = ~n60988 & ~n47874;
  assign n47876 = n5138 & ~n47875;
  assign n47877 = ~n47857 & ~n47876;
  assign n47878 = ~pi643 & pi1135;
  assign n47879 = ~pi606 & ~pi1135;
  assign n47880 = pi1136 & ~n47879;
  assign n47881 = pi1136 & ~n47878;
  assign n47882 = ~n47879 & n47881;
  assign n47883 = ~n47878 & n47880;
  assign n47884 = pi812 & ~pi1135;
  assign n47885 = ~pi787 & pi1135;
  assign n47886 = ~pi1136 & ~n47885;
  assign n47887 = ~pi1136 & ~n47884;
  assign n47888 = ~n47885 & n47887;
  assign n47889 = ~n47884 & n47886;
  assign n47890 = ~n60989 & ~n60990;
  assign n47891 = n47646 & ~n47890;
  assign n47892 = ~pi746 & n47662;
  assign n47893 = ~pi729 & pi1135;
  assign n47894 = ~pi881 & ~pi1136;
  assign n47895 = ~n47893 & ~n47894;
  assign n47896 = n47666 & n47895;
  assign n47897 = ~n47892 & n47896;
  assign n47898 = ~n47891 & ~n47897;
  assign n47899 = ~n5138 & ~n47898;
  assign n47900 = pi410 & n47676;
  assign n47901 = n47675 & ~n47900;
  assign n47902 = pi386 & ~pi591;
  assign n47903 = pi592 & ~n47902;
  assign n47904 = ~n47901 & ~n47903;
  assign n47905 = pi361 & n47683;
  assign n47906 = ~n47904 & ~n47905;
  assign n47907 = pi434 & n5089;
  assign n47908 = pi588 & ~n47907;
  assign n47909 = n47686 & ~n47908;
  assign n47910 = ~n47906 & n47909;
  assign n47911 = pi199 & ~pi1059;
  assign n47912 = ~pi199 & ~pi293;
  assign n47913 = ~n47686 & ~n47912;
  assign n47914 = ~n47686 & ~n47911;
  assign n47915 = ~n47912 & n47914;
  assign n47916 = ~n47911 & n47913;
  assign n47917 = ~n47910 & ~n60991;
  assign n47918 = n5138 & ~n47917;
  assign n47919 = ~n47899 & ~n47918;
  assign n47920 = pi199 & ~pi1036;
  assign n47921 = ~pi199 & ~pi255;
  assign n47922 = ~n47686 & ~n47921;
  assign n47923 = ~n47686 & ~n47920;
  assign n47924 = ~n47921 & n47923;
  assign n47925 = ~n47920 & n47922;
  assign n47926 = pi389 & n47790;
  assign n47927 = pi413 & pi591;
  assign n47928 = ~pi592 & n47927;
  assign n47929 = ~n47926 & ~n47928;
  assign n47930 = ~pi590 & ~n47929;
  assign n47931 = pi450 & n47683;
  assign n47932 = ~pi588 & ~n47931;
  assign n47933 = ~n47930 & n47932;
  assign n47934 = pi438 & n5089;
  assign n47935 = pi588 & ~n47934;
  assign n47936 = n47686 & ~n47935;
  assign n47937 = ~n47933 & n47936;
  assign n47938 = ~n60992 & ~n47937;
  assign n47939 = n5138 & ~n47938;
  assign n47940 = ~pi665 & pi1136;
  assign n47941 = ~pi791 & ~pi1136;
  assign n47942 = pi1135 & ~n47941;
  assign n47943 = pi1135 & ~n47940;
  assign n47944 = ~n47941 & n47943;
  assign n47945 = ~n47940 & n47942;
  assign n47946 = ~pi621 & pi1136;
  assign n47947 = ~pi810 & ~pi1136;
  assign n47948 = ~pi1135 & ~n47947;
  assign n47949 = ~pi1135 & ~n47946;
  assign n47950 = ~n47947 & n47949;
  assign n47951 = ~n47946 & n47948;
  assign n47952 = ~n60993 & ~n60994;
  assign n47953 = n47646 & ~n47952;
  assign n47954 = ~pi739 & n47662;
  assign n47955 = ~pi874 & ~pi1136;
  assign n47956 = ~pi690 & pi1135;
  assign n47957 = ~n47955 & ~n47956;
  assign n47958 = n47666 & n47957;
  assign n47959 = ~n47954 & n47958;
  assign n47960 = ~n47953 & ~n47959;
  assign n47961 = ~n5138 & ~n47960;
  assign n47962 = ~n47939 & ~n47961;
  assign n47963 = pi590 & ~pi592;
  assign n47964 = pi357 & n47963;
  assign n47965 = pi382 & n47674;
  assign n47966 = ~n47964 & ~n47965;
  assign n47967 = ~pi591 & ~n47966;
  assign n47968 = pi406 & ~pi592;
  assign n47969 = n47676 & n47968;
  assign n47970 = ~n47967 & ~n47969;
  assign n47971 = ~pi588 & ~n47970;
  assign n47972 = ~pi591 & ~pi592;
  assign n47973 = pi588 & ~pi590;
  assign n47974 = pi430 & n47973;
  assign n47975 = pi430 & n47972;
  assign n47976 = n47973 & n47975;
  assign n47977 = n47972 & n47974;
  assign n47978 = ~n47971 & ~n60995;
  assign n47979 = n47686 & ~n47978;
  assign n47980 = pi200 & pi1067;
  assign n47981 = ~pi200 & pi1044;
  assign n47982 = ~pi199 & ~n47981;
  assign n47983 = ~pi199 & ~n47980;
  assign n47984 = ~n47981 & n47983;
  assign n47985 = ~n47980 & n47982;
  assign n47986 = pi199 & ~pi1076;
  assign n47987 = ~n47686 & ~n47986;
  assign n47988 = ~n60996 & n47987;
  assign n47989 = ~n47979 & ~n47988;
  assign n47990 = n5138 & ~n47989;
  assign n47991 = pi860 & n47826;
  assign n47992 = pi728 & pi1135;
  assign n47993 = pi744 & ~pi1135;
  assign n47994 = pi1136 & ~n47993;
  assign n47995 = pi1136 & ~n47992;
  assign n47996 = ~n47993 & n47995;
  assign n47997 = ~n47992 & n47994;
  assign n47998 = ~n47991 & ~n60997;
  assign n47999 = n47665 & ~n47998;
  assign n48000 = pi1136 & ~n47645;
  assign n48001 = ~pi1134 & ~n48000;
  assign n48002 = pi657 & pi1135;
  assign n48003 = ~pi652 & ~pi1135;
  assign n48004 = pi1136 & ~n48003;
  assign n48005 = pi1136 & ~n48002;
  assign n48006 = ~n48003 & n48005;
  assign n48007 = ~n48002 & n48004;
  assign n48008 = pi813 & n47645;
  assign n48009 = n47826 & n48008;
  assign n48010 = ~n60998 & ~n48009;
  assign n48011 = n48001 & ~n48010;
  assign n48012 = ~n47999 & ~n48011;
  assign n48013 = ~n5138 & ~n48012;
  assign n48014 = ~n47990 & ~n48013;
  assign n48015 = pi351 & n47963;
  assign n48016 = pi376 & n47674;
  assign n48017 = ~n48015 & ~n48016;
  assign n48018 = ~pi591 & ~n48017;
  assign n48019 = pi401 & ~pi592;
  assign n48020 = n47676 & n48019;
  assign n48021 = ~n48018 & ~n48020;
  assign n48022 = ~pi588 & ~n48021;
  assign n48023 = pi426 & n47973;
  assign n48024 = pi426 & n47972;
  assign n48025 = n47973 & n48024;
  assign n48026 = n47972 & n48023;
  assign n48027 = ~n48022 & ~n60999;
  assign n48028 = n47686 & ~n48027;
  assign n48029 = pi200 & ~pi1036;
  assign n48030 = ~pi200 & ~pi1049;
  assign n48031 = ~pi200 & pi1049;
  assign n48032 = pi200 & pi1036;
  assign n48033 = ~n48031 & ~n48032;
  assign n48034 = ~n48029 & ~n48030;
  assign n48035 = ~pi199 & n61000;
  assign n48036 = pi199 & ~pi1079;
  assign n48037 = ~n47686 & ~n48036;
  assign n48038 = ~n48035 & n48037;
  assign n48039 = ~n48028 & ~n48038;
  assign n48040 = n5138 & ~n48039;
  assign n48041 = pi798 & n47826;
  assign n48042 = pi655 & pi1135;
  assign n48043 = ~pi658 & ~pi1135;
  assign n48044 = pi1136 & ~n48043;
  assign n48045 = pi1136 & ~n48042;
  assign n48046 = ~n48043 & n48045;
  assign n48047 = ~n48042 & n48044;
  assign n48048 = ~n48041 & ~n61001;
  assign n48049 = n47646 & ~n48048;
  assign n48050 = pi752 & n47662;
  assign n48051 = ~pi703 & pi1135;
  assign n48052 = ~pi843 & ~pi1136;
  assign n48053 = ~n48051 & ~n48052;
  assign n48054 = n47666 & n48053;
  assign n48055 = ~n48050 & n48054;
  assign n48056 = ~n48049 & ~n48055;
  assign n48057 = ~n5138 & ~n48056;
  assign n48058 = ~n48040 & ~n48057;
  assign n48059 = pi352 & n47963;
  assign n48060 = pi317 & n47674;
  assign n48061 = ~n48059 & ~n48060;
  assign n48062 = ~pi591 & ~n48061;
  assign n48063 = pi402 & ~pi592;
  assign n48064 = n47676 & n48063;
  assign n48065 = ~n48062 & ~n48064;
  assign n48066 = ~pi588 & ~n48065;
  assign n48067 = pi427 & n47973;
  assign n48068 = pi427 & n47972;
  assign n48069 = n47973 & n48068;
  assign n48070 = n47972 & n48067;
  assign n48071 = ~n48066 & ~n61002;
  assign n48072 = n47686 & ~n48071;
  assign n48073 = pi200 & ~pi1065;
  assign n48074 = ~pi200 & ~pi1084;
  assign n48075 = ~pi200 & pi1084;
  assign n48076 = pi200 & pi1065;
  assign n48077 = ~n48075 & ~n48076;
  assign n48078 = ~n48073 & ~n48074;
  assign n48079 = ~pi199 & n61003;
  assign n48080 = pi199 & ~pi1078;
  assign n48081 = ~n47686 & ~n48080;
  assign n48082 = ~n48079 & n48081;
  assign n48083 = ~n48072 & ~n48082;
  assign n48084 = n5138 & ~n48083;
  assign n48085 = pi649 & pi1135;
  assign n48086 = ~pi656 & ~pi1135;
  assign n48087 = pi1136 & ~n48086;
  assign n48088 = pi1136 & ~n48085;
  assign n48089 = ~n48086 & n48088;
  assign n48090 = ~n48085 & n48087;
  assign n48091 = pi801 & n47826;
  assign n48092 = ~pi1134 & ~n48091;
  assign n48093 = ~n61004 & n48092;
  assign n48094 = pi770 & ~pi1135;
  assign n48095 = ~pi726 & pi1135;
  assign n48096 = pi1136 & ~n48095;
  assign n48097 = pi1136 & ~n48094;
  assign n48098 = ~n48095 & n48097;
  assign n48099 = ~n48094 & n48096;
  assign n48100 = pi844 & n47826;
  assign n48101 = pi1134 & ~n48100;
  assign n48102 = ~n61005 & n48101;
  assign n48103 = n47819 & ~n48102;
  assign n48104 = ~n48093 & n48103;
  assign n48105 = ~n48084 & ~n48104;
  assign n48106 = pi753 & n47662;
  assign n48107 = ~pi847 & ~pi1136;
  assign n48108 = pi702 & pi1135;
  assign n48109 = ~n48107 & ~n48108;
  assign n48110 = n47666 & n48109;
  assign n48111 = ~n48106 & n48110;
  assign n48112 = pi1136 & n47645;
  assign n48113 = ~pi618 & ~pi1135;
  assign n48114 = ~pi627 & pi1135;
  assign n48115 = ~pi1134 & ~n48114;
  assign n48116 = ~pi1134 & ~n48113;
  assign n48117 = ~n48114 & n48116;
  assign n48118 = ~n48113 & n48115;
  assign n48119 = n48112 & n61006;
  assign n48120 = ~n5138 & ~n48119;
  assign n48121 = ~n48111 & n48120;
  assign n48122 = pi370 & n47790;
  assign n48123 = pi395 & pi591;
  assign n48124 = ~pi592 & n48123;
  assign n48125 = ~n48122 & ~n48124;
  assign n48126 = ~pi590 & ~n48125;
  assign n48127 = pi347 & n47683;
  assign n48128 = ~n48126 & ~n48127;
  assign n48129 = ~pi588 & n47686;
  assign n48130 = ~n48128 & n48129;
  assign n48131 = ~pi200 & ~pi304;
  assign n48132 = pi200 & ~pi1048;
  assign n48133 = ~n48131 & ~n48132;
  assign n48134 = pi200 & pi1048;
  assign n48135 = ~pi200 & pi304;
  assign n48136 = ~pi199 & ~n48135;
  assign n48137 = ~n48134 & n48136;
  assign n48138 = ~pi199 & ~n48133;
  assign n48139 = pi199 & ~pi1055;
  assign n48140 = ~n47686 & ~n48139;
  assign n48141 = ~n61007 & n48140;
  assign n48142 = n5089 & n47686;
  assign n48143 = pi420 & pi588;
  assign n48144 = n48142 & n48143;
  assign n48145 = n5138 & ~n48144;
  assign n48146 = ~n48141 & n48145;
  assign n48147 = ~n48130 & n48146;
  assign n48148 = ~n48141 & ~n48144;
  assign n48149 = ~n48130 & n48148;
  assign n48150 = n5138 & ~n48149;
  assign n48151 = ~n48111 & ~n48119;
  assign n48152 = ~n5138 & ~n48151;
  assign n48153 = ~n48150 & ~n48152;
  assign n48154 = ~n48121 & ~n48147;
  assign n48155 = n47686 & n47790;
  assign n48156 = pi442 & n48155;
  assign n48157 = ~pi592 & n47686;
  assign n48158 = pi328 & pi591;
  assign n48159 = n48157 & n48158;
  assign n48160 = ~n48156 & ~n48159;
  assign n48161 = ~pi590 & ~n48160;
  assign n48162 = pi321 & n47686;
  assign n48163 = n47683 & n48162;
  assign n48164 = ~n48161 & ~n48163;
  assign n48165 = ~pi588 & ~n48164;
  assign n48166 = ~pi200 & ~pi305;
  assign n48167 = pi200 & ~pi1084;
  assign n48168 = ~n48166 & ~n48167;
  assign n48169 = pi200 & pi1084;
  assign n48170 = ~pi200 & pi305;
  assign n48171 = ~pi199 & ~n48170;
  assign n48172 = ~n48169 & n48171;
  assign n48173 = ~pi199 & ~n48168;
  assign n48174 = pi199 & ~pi1058;
  assign n48175 = ~n47686 & ~n48174;
  assign n48176 = ~n61009 & n48175;
  assign n48177 = n47686 & n47972;
  assign n48178 = pi459 & n47973;
  assign n48179 = n48177 & n48178;
  assign n48180 = n5138 & ~n48179;
  assign n48181 = ~n48176 & n48180;
  assign n48182 = ~n48165 & n48181;
  assign n48183 = pi754 & n47662;
  assign n48184 = pi709 & pi1135;
  assign n48185 = ~pi857 & ~pi1136;
  assign n48186 = ~n48184 & ~n48185;
  assign n48187 = n47645 & ~n47664;
  assign n48188 = pi1134 & ~n48184;
  assign n48189 = ~n48185 & n48188;
  assign n48190 = n48187 & n48189;
  assign n48191 = n47666 & n48186;
  assign n48192 = ~n48183 & n61010;
  assign n48193 = ~pi609 & ~pi1135;
  assign n48194 = ~pi660 & pi1135;
  assign n48195 = ~pi1134 & ~n48194;
  assign n48196 = ~pi1134 & ~n48193;
  assign n48197 = ~n48194 & n48196;
  assign n48198 = ~n48193 & n48195;
  assign n48199 = n48112 & n61011;
  assign n48200 = ~n5138 & ~n48199;
  assign n48201 = ~n48192 & n48200;
  assign po865 = ~n48182 & ~n48201;
  assign n48203 = pi755 & n47662;
  assign n48204 = ~pi858 & ~pi1136;
  assign n48205 = pi725 & pi1135;
  assign n48206 = ~n48204 & ~n48205;
  assign n48207 = n47666 & n48206;
  assign n48208 = ~n48203 & n48207;
  assign n48209 = ~pi630 & ~pi1135;
  assign n48210 = ~pi647 & pi1135;
  assign n48211 = ~pi1134 & ~n48210;
  assign n48212 = ~pi1134 & ~n48209;
  assign n48213 = ~n48210 & n48212;
  assign n48214 = ~n48209 & n48211;
  assign n48215 = n48112 & n61012;
  assign n48216 = ~n5138 & ~n48215;
  assign n48217 = ~n48208 & n48216;
  assign n48218 = pi373 & n47790;
  assign n48219 = pi398 & pi591;
  assign n48220 = ~pi592 & n48219;
  assign n48221 = ~n48218 & ~n48220;
  assign n48222 = ~pi590 & ~n48221;
  assign n48223 = pi348 & n47683;
  assign n48224 = ~n48222 & ~n48223;
  assign n48225 = n48129 & ~n48224;
  assign n48226 = ~pi200 & ~pi306;
  assign n48227 = pi200 & ~pi1059;
  assign n48228 = ~n48226 & ~n48227;
  assign n48229 = pi200 & pi1059;
  assign n48230 = ~pi200 & pi306;
  assign n48231 = ~pi199 & ~n48230;
  assign n48232 = ~n48229 & n48231;
  assign n48233 = ~pi199 & ~n48228;
  assign n48234 = pi199 & ~pi1087;
  assign n48235 = ~n47686 & ~n48234;
  assign n48236 = ~n61013 & n48235;
  assign n48237 = pi423 & pi588;
  assign n48238 = n48142 & n48237;
  assign n48239 = n5138 & ~n48238;
  assign n48240 = ~n48236 & n48239;
  assign n48241 = ~n48225 & n48240;
  assign n48242 = ~n48236 & ~n48238;
  assign n48243 = ~n48225 & n48242;
  assign n48244 = n5138 & ~n48243;
  assign n48245 = ~n48208 & ~n48215;
  assign n48246 = ~n5138 & ~n48245;
  assign n48247 = ~n48244 & ~n48246;
  assign n48248 = ~n48217 & ~n48241;
  assign n48249 = ~pi644 & ~pi1135;
  assign n48250 = ~pi715 & pi1135;
  assign n48251 = ~pi1134 & ~n48250;
  assign n48252 = ~pi1134 & ~n48249;
  assign n48253 = ~n48250 & n48252;
  assign n48254 = ~n48249 & n48251;
  assign n48255 = n48112 & n61015;
  assign n48256 = pi751 & n47662;
  assign n48257 = ~pi842 & ~pi1136;
  assign n48258 = pi701 & pi1135;
  assign n48259 = ~n48257 & ~n48258;
  assign n48260 = pi1134 & ~n48258;
  assign n48261 = ~n48257 & n48260;
  assign n48262 = n48187 & n48261;
  assign n48263 = n47666 & n48259;
  assign n48264 = ~n48256 & n61016;
  assign n48265 = ~n48255 & ~n48264;
  assign n48266 = ~n5138 & ~n48265;
  assign n48267 = pi374 & n47790;
  assign n48268 = pi400 & pi591;
  assign n48269 = ~pi592 & n48268;
  assign n48270 = ~n48267 & ~n48269;
  assign n48271 = ~pi590 & ~n48270;
  assign n48272 = pi350 & n47683;
  assign n48273 = ~n48271 & ~n48272;
  assign n48274 = ~pi588 & ~n48273;
  assign n48275 = pi425 & n47973;
  assign n48276 = pi425 & n47972;
  assign n48277 = n47973 & n48276;
  assign n48278 = n47972 & n48275;
  assign n48279 = n47686 & ~n61017;
  assign n48280 = ~n48274 & n48279;
  assign n48281 = pi298 & n36719;
  assign n48282 = pi1044 & n45424;
  assign n48283 = pi199 & pi1035;
  assign n48284 = ~n47686 & ~n48283;
  assign n48285 = ~n48282 & n48284;
  assign n48286 = ~n48281 & n48284;
  assign n48287 = ~n48282 & n48286;
  assign n48288 = ~n48281 & n48285;
  assign n48289 = n5138 & ~n61018;
  assign n48290 = ~n48280 & n48289;
  assign n48291 = ~n48266 & ~n48290;
  assign n48292 = pi756 & n47662;
  assign n48293 = ~pi854 & ~pi1136;
  assign n48294 = pi734 & pi1135;
  assign n48295 = ~n48293 & ~n48294;
  assign n48296 = n47666 & n48295;
  assign n48297 = ~n48292 & n48296;
  assign n48298 = ~pi629 & ~pi1135;
  assign n48299 = ~pi628 & pi1135;
  assign n48300 = ~pi1134 & ~n48299;
  assign n48301 = ~pi1134 & ~n48298;
  assign n48302 = ~n48299 & n48301;
  assign n48303 = ~n48298 & n48300;
  assign n48304 = n48112 & n61019;
  assign n48305 = ~n5138 & ~n48304;
  assign n48306 = ~n48297 & n48305;
  assign n48307 = pi371 & n47790;
  assign n48308 = pi396 & pi591;
  assign n48309 = ~pi592 & n48308;
  assign n48310 = ~n48307 & ~n48309;
  assign n48311 = ~pi590 & ~n48310;
  assign n48312 = pi322 & n47683;
  assign n48313 = ~n48311 & ~n48312;
  assign n48314 = n48129 & ~n48313;
  assign n48315 = ~pi200 & ~pi309;
  assign n48316 = pi200 & ~pi1072;
  assign n48317 = ~n48315 & ~n48316;
  assign n48318 = pi200 & pi1072;
  assign n48319 = ~pi200 & pi309;
  assign n48320 = ~pi199 & ~n48319;
  assign n48321 = ~n48318 & n48320;
  assign n48322 = ~pi199 & ~n48317;
  assign n48323 = pi199 & ~pi1051;
  assign n48324 = ~n47686 & ~n48323;
  assign n48325 = ~n61020 & n48324;
  assign n48326 = pi421 & pi588;
  assign n48327 = n48142 & n48326;
  assign n48328 = n5138 & ~n48327;
  assign n48329 = ~n48325 & n48328;
  assign n48330 = ~n48314 & n48329;
  assign n48331 = ~n48325 & ~n48327;
  assign n48332 = ~n48314 & n48331;
  assign n48333 = n5138 & ~n48332;
  assign n48334 = ~n48297 & ~n48304;
  assign n48335 = ~n5138 & ~n48334;
  assign n48336 = ~n48333 & ~n48335;
  assign n48337 = ~n48306 & ~n48330;
  assign n48338 = pi461 & n47963;
  assign n48339 = pi439 & n47674;
  assign n48340 = ~n48338 & ~n48339;
  assign n48341 = ~pi591 & ~n48340;
  assign n48342 = pi326 & ~pi592;
  assign n48343 = n47676 & n48342;
  assign n48344 = ~n48341 & ~n48343;
  assign n48345 = ~pi588 & ~n48344;
  assign n48346 = pi449 & n47973;
  assign n48347 = pi449 & n47972;
  assign n48348 = n47973 & n48347;
  assign n48349 = n47972 & n48346;
  assign n48350 = ~n48345 & ~n61022;
  assign n48351 = n47686 & ~n48350;
  assign n48352 = pi200 & pi1039;
  assign n48353 = ~pi200 & pi1053;
  assign n48354 = ~pi199 & ~n48353;
  assign n48355 = ~pi199 & ~n48352;
  assign n48356 = ~n48353 & n48355;
  assign n48357 = ~n48352 & n48354;
  assign n48358 = pi199 & ~pi1057;
  assign n48359 = ~n47686 & ~n48358;
  assign n48360 = ~n61023 & n48359;
  assign n48361 = ~n48351 & ~n48360;
  assign n48362 = n5138 & ~n48361;
  assign n48363 = pi867 & n47826;
  assign n48364 = pi697 & pi1135;
  assign n48365 = pi762 & ~pi1135;
  assign n48366 = pi1136 & ~n48365;
  assign n48367 = pi1136 & ~n48364;
  assign n48368 = ~n48365 & n48367;
  assign n48369 = ~n48364 & n48366;
  assign n48370 = ~n48363 & ~n61024;
  assign n48371 = n47665 & ~n48370;
  assign n48372 = pi693 & pi1135;
  assign n48373 = ~pi653 & ~pi1135;
  assign n48374 = pi1136 & ~n48373;
  assign n48375 = pi1136 & ~n48372;
  assign n48376 = ~n48373 & n48375;
  assign n48377 = ~n48372 & n48374;
  assign n48378 = pi816 & n47645;
  assign n48379 = n47826 & n48378;
  assign n48380 = ~n61025 & ~n48379;
  assign n48381 = n48001 & ~n48380;
  assign n48382 = ~n48371 & ~n48381;
  assign n48383 = ~n5138 & ~n48382;
  assign n48384 = ~n48362 & ~n48383;
  assign n48385 = pi440 & n48155;
  assign n48386 = pi329 & pi591;
  assign n48387 = n48157 & n48386;
  assign n48388 = ~n48385 & ~n48387;
  assign n48389 = ~pi590 & ~n48388;
  assign n48390 = pi349 & n47686;
  assign n48391 = n47683 & n48390;
  assign n48392 = ~n48389 & ~n48391;
  assign n48393 = ~pi588 & ~n48392;
  assign n48394 = ~pi200 & ~pi307;
  assign n48395 = pi200 & ~pi1053;
  assign n48396 = ~n48394 & ~n48395;
  assign n48397 = pi200 & pi1053;
  assign n48398 = ~pi200 & pi307;
  assign n48399 = ~pi199 & ~n48398;
  assign n48400 = ~n48397 & n48399;
  assign n48401 = ~pi199 & ~n48396;
  assign n48402 = pi199 & ~pi1043;
  assign n48403 = ~n47686 & ~n48402;
  assign n48404 = ~n61026 & n48403;
  assign n48405 = pi454 & n47973;
  assign n48406 = n48177 & n48405;
  assign n48407 = n5138 & ~n48406;
  assign n48408 = ~n48404 & n48407;
  assign n48409 = ~n48393 & n48408;
  assign n48410 = pi761 & n47662;
  assign n48411 = pi738 & pi1135;
  assign n48412 = ~pi845 & ~pi1136;
  assign n48413 = ~n48411 & ~n48412;
  assign n48414 = pi1134 & ~n48411;
  assign n48415 = ~n48412 & n48414;
  assign n48416 = n48187 & n48415;
  assign n48417 = n47666 & n48413;
  assign n48418 = ~n48410 & n61027;
  assign n48419 = ~pi626 & ~pi1135;
  assign n48420 = ~pi641 & pi1135;
  assign n48421 = ~pi1134 & ~n48420;
  assign n48422 = ~pi1134 & ~n48419;
  assign n48423 = ~n48420 & n48422;
  assign n48424 = ~n48419 & n48421;
  assign n48425 = n48112 & n61028;
  assign n48426 = ~n5138 & ~n48425;
  assign n48427 = ~n48418 & n48426;
  assign po873 = ~n48409 & ~n48427;
  assign n48429 = pi318 & pi591;
  assign n48430 = ~pi592 & n48429;
  assign n48431 = ~pi591 & n3707;
  assign n48432 = ~n48430 & ~n48431;
  assign n48433 = ~pi590 & ~n48432;
  assign n48434 = pi462 & n47683;
  assign n48435 = ~n48433 & ~n48434;
  assign n48436 = n48129 & ~n48435;
  assign n48437 = pi200 & ~pi1070;
  assign n48438 = ~pi200 & ~pi1048;
  assign n48439 = ~pi200 & pi1048;
  assign n48440 = pi200 & pi1070;
  assign n48441 = ~n48439 & ~n48440;
  assign n48442 = ~n48437 & ~n48438;
  assign n48443 = ~pi199 & n61029;
  assign n48444 = pi199 & ~pi1074;
  assign n48445 = ~n47686 & ~n48444;
  assign n48446 = ~n48443 & n48445;
  assign n48447 = pi448 & pi588;
  assign n48448 = n48142 & n48447;
  assign n48449 = ~n48446 & ~n48448;
  assign n48450 = ~n48436 & n48449;
  assign n48451 = n5138 & ~n48450;
  assign n48452 = pi800 & n47826;
  assign n48453 = pi669 & pi1135;
  assign n48454 = ~pi645 & ~pi1135;
  assign n48455 = pi1136 & ~n48454;
  assign n48456 = pi1136 & ~n48453;
  assign n48457 = ~n48454 & n48456;
  assign n48458 = ~n48453 & n48455;
  assign n48459 = ~n48452 & ~n61030;
  assign n48460 = n47646 & ~n48459;
  assign n48461 = pi768 & n47662;
  assign n48462 = ~pi839 & ~pi1136;
  assign n48463 = ~pi705 & pi1135;
  assign n48464 = ~n48462 & ~n48463;
  assign n48465 = pi1134 & ~n48463;
  assign n48466 = ~n48462 & n48465;
  assign n48467 = n48187 & n48466;
  assign n48468 = n47666 & n48464;
  assign n48469 = ~n48461 & n61031;
  assign n48470 = ~n48460 & ~n48469;
  assign n48471 = ~n5138 & ~n48470;
  assign n48472 = ~n48451 & ~n48471;
  assign n48473 = pi369 & n48155;
  assign n48474 = pi394 & pi591;
  assign n48475 = n48157 & n48474;
  assign n48476 = ~n48473 & ~n48475;
  assign n48477 = ~pi590 & ~n48476;
  assign n48478 = pi315 & n47686;
  assign n48479 = n47683 & n48478;
  assign n48480 = ~n48477 & ~n48479;
  assign n48481 = ~pi588 & ~n48480;
  assign n48482 = ~pi200 & ~pi303;
  assign n48483 = pi200 & ~pi1049;
  assign n48484 = ~n48482 & ~n48483;
  assign n48485 = pi200 & pi1049;
  assign n48486 = ~pi200 & pi303;
  assign n48487 = ~pi199 & ~n48486;
  assign n48488 = ~n48485 & n48487;
  assign n48489 = ~pi199 & ~n48484;
  assign n48490 = pi199 & ~pi1080;
  assign n48491 = ~n47686 & ~n48490;
  assign n48492 = ~n61032 & n48491;
  assign n48493 = pi419 & n47973;
  assign n48494 = n48177 & n48493;
  assign n48495 = n5138 & ~n48494;
  assign n48496 = ~n48492 & n48495;
  assign n48497 = ~n48481 & n48496;
  assign n48498 = pi767 & n47662;
  assign n48499 = pi698 & pi1135;
  assign n48500 = ~pi853 & ~pi1136;
  assign n48501 = ~n48499 & ~n48500;
  assign n48502 = pi1134 & ~n48499;
  assign n48503 = ~n48500 & n48502;
  assign n48504 = n48187 & n48503;
  assign n48505 = n47666 & n48501;
  assign n48506 = ~n48498 & n61033;
  assign n48507 = ~pi608 & ~pi1135;
  assign n48508 = ~pi625 & pi1135;
  assign n48509 = ~pi1134 & ~n48508;
  assign n48510 = ~pi1134 & ~n48507;
  assign n48511 = ~n48508 & n48510;
  assign n48512 = ~n48507 & n48509;
  assign n48513 = n48112 & n61034;
  assign n48514 = ~n5138 & ~n48513;
  assign n48515 = ~n48506 & n48514;
  assign po875 = ~n48497 & ~n48515;
  assign n48517 = pi378 & n47790;
  assign n48518 = pi325 & pi591;
  assign n48519 = ~pi592 & n48518;
  assign n48520 = ~n48517 & ~n48519;
  assign n48521 = ~pi590 & ~n48520;
  assign n48522 = pi353 & n47683;
  assign n48523 = ~n48521 & ~n48522;
  assign n48524 = n48129 & ~n48523;
  assign n48525 = pi200 & ~pi1062;
  assign n48526 = ~pi200 & ~pi1072;
  assign n48527 = ~pi200 & pi1072;
  assign n48528 = pi200 & pi1062;
  assign n48529 = ~n48527 & ~n48528;
  assign n48530 = ~n48525 & ~n48526;
  assign n48531 = ~pi199 & n61035;
  assign n48532 = pi199 & ~pi1063;
  assign n48533 = ~n47686 & ~n48532;
  assign n48534 = ~n48531 & n48533;
  assign n48535 = pi451 & pi588;
  assign n48536 = n48142 & n48535;
  assign n48537 = ~n48534 & ~n48536;
  assign n48538 = ~n48524 & n48537;
  assign n48539 = n5138 & ~n48538;
  assign n48540 = pi807 & n47826;
  assign n48541 = pi650 & pi1135;
  assign n48542 = ~pi636 & ~pi1135;
  assign n48543 = pi1136 & ~n48542;
  assign n48544 = pi1136 & ~n48541;
  assign n48545 = ~n48542 & n48544;
  assign n48546 = ~n48541 & n48543;
  assign n48547 = ~n48540 & ~n61036;
  assign n48548 = n47646 & ~n48547;
  assign n48549 = pi774 & n47662;
  assign n48550 = ~pi868 & ~pi1136;
  assign n48551 = ~pi687 & pi1135;
  assign n48552 = ~n48550 & ~n48551;
  assign n48553 = pi1134 & ~n48551;
  assign n48554 = ~n48550 & n48553;
  assign n48555 = n48187 & n48554;
  assign n48556 = n47666 & n48552;
  assign n48557 = ~n48549 & n61037;
  assign n48558 = ~n48548 & ~n48557;
  assign n48559 = ~n5138 & ~n48558;
  assign n48560 = ~n48539 & ~n48559;
  assign n48561 = pi356 & n47963;
  assign n48562 = pi381 & n47674;
  assign n48563 = ~n48561 & ~n48562;
  assign n48564 = ~pi591 & ~n48563;
  assign n48565 = pi405 & ~pi592;
  assign n48566 = n47676 & n48565;
  assign n48567 = ~n48564 & ~n48566;
  assign n48568 = ~pi588 & ~n48567;
  assign n48569 = pi445 & n47973;
  assign n48570 = pi445 & n47972;
  assign n48571 = n47973 & n48570;
  assign n48572 = n47972 & n48569;
  assign n48573 = ~n48568 & ~n61038;
  assign n48574 = n47686 & ~n48573;
  assign n48575 = pi200 & pi1040;
  assign n48576 = ~pi200 & pi1037;
  assign n48577 = ~pi199 & ~n48576;
  assign n48578 = ~pi199 & ~n48575;
  assign n48579 = ~n48576 & n48578;
  assign n48580 = ~n48575 & n48577;
  assign n48581 = pi199 & ~pi1081;
  assign n48582 = ~n47686 & ~n48581;
  assign n48583 = ~n61039 & n48582;
  assign n48584 = ~n48574 & ~n48583;
  assign n48585 = n5138 & ~n48584;
  assign n48586 = pi880 & n47826;
  assign n48587 = pi684 & pi1135;
  assign n48588 = pi750 & ~pi1135;
  assign n48589 = pi1136 & ~n48588;
  assign n48590 = pi1136 & ~n48587;
  assign n48591 = ~n48588 & n48590;
  assign n48592 = ~n48587 & n48589;
  assign n48593 = ~n48586 & ~n61040;
  assign n48594 = n47665 & ~n48593;
  assign n48595 = pi654 & pi1135;
  assign n48596 = ~pi651 & ~pi1135;
  assign n48597 = pi1136 & ~n48596;
  assign n48598 = pi1136 & ~n48595;
  assign n48599 = ~n48596 & n48598;
  assign n48600 = ~n48595 & n48597;
  assign n48601 = pi794 & n47645;
  assign n48602 = n47826 & n48601;
  assign n48603 = ~n61041 & ~n48602;
  assign n48604 = n48001 & ~n48603;
  assign n48605 = ~n48594 & ~n48604;
  assign n48606 = ~n5138 & ~n48605;
  assign n48607 = ~n48585 & ~n48606;
  assign n48608 = pi379 & n47790;
  assign n48609 = pi403 & pi591;
  assign n48610 = ~pi592 & n48609;
  assign n48611 = ~n48608 & ~n48610;
  assign n48612 = ~pi590 & ~n48611;
  assign n48613 = pi354 & n47683;
  assign n48614 = ~n48612 & ~n48613;
  assign n48615 = n48129 & ~n48614;
  assign n48616 = pi200 & ~pi1069;
  assign n48617 = ~pi200 & ~pi1059;
  assign n48618 = ~pi200 & pi1059;
  assign n48619 = pi200 & pi1069;
  assign n48620 = ~n48618 & ~n48619;
  assign n48621 = ~n48616 & ~n48617;
  assign n48622 = ~pi199 & n61042;
  assign n48623 = pi199 & ~pi1045;
  assign n48624 = ~n47686 & ~n48623;
  assign n48625 = ~n48622 & n48624;
  assign n48626 = pi428 & pi588;
  assign n48627 = n48142 & n48626;
  assign n48628 = ~n48625 & ~n48627;
  assign n48629 = ~n48615 & n48628;
  assign n48630 = n5138 & ~n48629;
  assign n48631 = ~pi851 & pi1134;
  assign n48632 = ~pi795 & ~pi1134;
  assign n48633 = ~pi1136 & ~n48632;
  assign n48634 = ~pi1136 & ~n48631;
  assign n48635 = ~n48632 & n48634;
  assign n48636 = ~n48631 & n48633;
  assign n48637 = pi776 & pi1134;
  assign n48638 = ~pi640 & ~pi1134;
  assign n48639 = pi1136 & ~n48638;
  assign n48640 = pi1136 & ~n48637;
  assign n48641 = ~n48638 & n48640;
  assign n48642 = ~n48637 & n48639;
  assign n48643 = ~n61043 & ~n61044;
  assign n48644 = ~pi1135 & ~n48643;
  assign n48645 = pi732 & ~pi1134;
  assign n48646 = pi694 & pi1134;
  assign n48647 = pi1135 & pi1136;
  assign n48648 = ~n48646 & n48647;
  assign n48649 = ~n48645 & n48648;
  assign n48650 = ~n48644 & ~n48649;
  assign n48651 = n47819 & ~n48650;
  assign n48652 = ~n48630 & ~n48651;
  assign n48653 = pi199 & ~pi1065;
  assign n48654 = ~pi199 & ~pi257;
  assign n48655 = ~n47686 & ~n48654;
  assign n48656 = ~n48653 & n48655;
  assign n48657 = pi365 & n47790;
  assign n48658 = pi334 & pi591;
  assign n48659 = ~pi592 & n48658;
  assign n48660 = ~n48657 & ~n48659;
  assign n48661 = ~pi590 & ~n48660;
  assign n48662 = pi323 & n47683;
  assign n48663 = ~pi588 & ~n48662;
  assign n48664 = ~n48661 & n48663;
  assign n48665 = pi464 & n5089;
  assign n48666 = pi588 & ~n48665;
  assign n48667 = n47686 & ~n48666;
  assign n48668 = ~n48664 & n48667;
  assign n48669 = ~n48656 & ~n48668;
  assign n48670 = n5138 & ~n48669;
  assign n48671 = ~pi634 & pi1136;
  assign n48672 = ~pi784 & ~pi1136;
  assign n48673 = pi1135 & ~n48672;
  assign n48674 = pi1135 & ~n48671;
  assign n48675 = ~n48672 & n48674;
  assign n48676 = ~n48671 & n48673;
  assign n48677 = ~pi633 & pi1136;
  assign n48678 = ~pi815 & ~pi1136;
  assign n48679 = ~pi1135 & ~n48678;
  assign n48680 = ~pi1135 & ~n48677;
  assign n48681 = ~n48678 & n48680;
  assign n48682 = ~n48677 & n48679;
  assign n48683 = ~n61045 & ~n61046;
  assign n48684 = n47646 & ~n48683;
  assign n48685 = ~pi766 & n47662;
  assign n48686 = ~pi855 & ~pi1136;
  assign n48687 = ~pi700 & pi1135;
  assign n48688 = ~n48686 & ~n48687;
  assign n48689 = n47666 & n48688;
  assign n48690 = ~n48685 & n48689;
  assign n48691 = ~n48684 & ~n48690;
  assign n48692 = ~n5138 & ~n48691;
  assign n48693 = ~n48670 & ~n48692;
  assign n48694 = pi404 & n47676;
  assign n48695 = n47675 & ~n48694;
  assign n48696 = pi380 & ~pi591;
  assign n48697 = pi592 & ~n48696;
  assign n48698 = ~n48695 & ~n48697;
  assign n48699 = pi355 & n47683;
  assign n48700 = ~n48698 & ~n48699;
  assign n48701 = pi429 & n5089;
  assign n48702 = pi588 & ~n48701;
  assign n48703 = n47686 & ~n48702;
  assign n48704 = ~n48700 & n48703;
  assign n48705 = pi199 & ~pi1084;
  assign n48706 = ~pi199 & ~pi292;
  assign n48707 = ~n47686 & ~n48706;
  assign n48708 = ~n47686 & ~n48705;
  assign n48709 = ~n48706 & n48708;
  assign n48710 = ~n48705 & n48707;
  assign n48711 = ~n48704 & ~n61047;
  assign n48712 = n5138 & ~n48711;
  assign n48713 = pi662 & pi1135;
  assign n48714 = pi614 & ~pi1135;
  assign n48715 = pi1136 & ~n48714;
  assign n48716 = pi1136 & ~n48713;
  assign n48717 = ~n48714 & n48716;
  assign n48718 = ~n48713 & n48715;
  assign n48719 = pi785 & pi1135;
  assign n48720 = pi811 & ~pi1135;
  assign n48721 = ~pi1136 & ~n48720;
  assign n48722 = ~pi1136 & ~n48719;
  assign n48723 = ~n48720 & n48722;
  assign n48724 = ~n48719 & n48721;
  assign n48725 = ~n61048 & ~n61049;
  assign n48726 = ~pi1134 & ~n48725;
  assign n48727 = ~pi727 & pi1135;
  assign n48728 = ~pi772 & ~pi1135;
  assign n48729 = pi1136 & ~n48728;
  assign n48730 = pi1136 & ~n48727;
  assign n48731 = ~n48728 & n48730;
  assign n48732 = ~n48727 & n48729;
  assign n48733 = pi872 & n47826;
  assign n48734 = pi1134 & ~n48733;
  assign n48735 = ~n61050 & n48734;
  assign n48736 = n47819 & ~n48735;
  assign n48737 = ~n48726 & n48736;
  assign n48738 = ~n48712 & ~n48737;
  assign n48739 = ~pi638 & pi1135;
  assign n48740 = ~pi607 & ~pi1135;
  assign n48741 = pi1136 & ~n48740;
  assign n48742 = pi1136 & ~n48739;
  assign n48743 = ~n48740 & n48742;
  assign n48744 = ~n48739 & n48741;
  assign n48745 = pi799 & ~pi1135;
  assign n48746 = ~pi790 & pi1135;
  assign n48747 = ~pi1136 & ~n48746;
  assign n48748 = ~pi1136 & ~n48745;
  assign n48749 = ~n48746 & n48748;
  assign n48750 = ~n48745 & n48747;
  assign n48751 = ~n61051 & ~n61052;
  assign n48752 = n47646 & ~n48751;
  assign n48753 = ~pi764 & n47662;
  assign n48754 = ~pi691 & pi1135;
  assign n48755 = ~pi873 & ~pi1136;
  assign n48756 = ~n48754 & ~n48755;
  assign n48757 = n47666 & n48756;
  assign n48758 = ~n48753 & n48757;
  assign n48759 = ~n48752 & ~n48758;
  assign n48760 = ~n5138 & ~n48759;
  assign n48761 = pi456 & n47676;
  assign n48762 = n47675 & ~n48761;
  assign n48763 = pi337 & ~pi591;
  assign n48764 = pi592 & ~n48763;
  assign n48765 = ~n48762 & ~n48764;
  assign n48766 = pi441 & n47683;
  assign n48767 = ~n48765 & ~n48766;
  assign n48768 = pi443 & n5089;
  assign n48769 = pi588 & ~n48768;
  assign n48770 = n47686 & ~n48769;
  assign n48771 = ~n48767 & n48770;
  assign n48772 = pi199 & ~pi1044;
  assign n48773 = ~pi199 & ~pi297;
  assign n48774 = ~n47686 & ~n48773;
  assign n48775 = ~n47686 & ~n48772;
  assign n48776 = ~n48773 & n48775;
  assign n48777 = ~n48772 & n48774;
  assign n48778 = ~n48771 & ~n61053;
  assign n48779 = n5138 & ~n48778;
  assign n48780 = ~n48760 & ~n48779;
  assign n48781 = pi319 & n47676;
  assign n48782 = n47675 & ~n48781;
  assign n48783 = pi338 & ~pi591;
  assign n48784 = pi592 & ~n48783;
  assign n48785 = ~n48782 & ~n48784;
  assign n48786 = pi458 & n47683;
  assign n48787 = ~n48785 & ~n48786;
  assign n48788 = pi444 & n5089;
  assign n48789 = pi588 & ~n48788;
  assign n48790 = n47686 & ~n48789;
  assign n48791 = ~n48787 & n48790;
  assign n48792 = pi199 & ~pi1072;
  assign n48793 = ~pi199 & ~pi294;
  assign n48794 = ~n47686 & ~n48793;
  assign n48795 = ~n47686 & ~n48792;
  assign n48796 = ~n48793 & n48795;
  assign n48797 = ~n48792 & n48794;
  assign n48798 = ~n48791 & ~n61054;
  assign n48799 = n5138 & ~n48798;
  assign n48800 = pi681 & pi1136;
  assign n48801 = pi792 & ~pi1136;
  assign n48802 = pi1135 & ~n48801;
  assign n48803 = pi1135 & ~n48800;
  assign n48804 = ~n48801 & n48803;
  assign n48805 = ~n48800 & n48802;
  assign n48806 = pi642 & pi1136;
  assign n48807 = ~pi809 & ~pi1136;
  assign n48808 = ~pi1135 & ~n48807;
  assign n48809 = ~pi1135 & ~n48806;
  assign n48810 = ~n48807 & n48809;
  assign n48811 = ~n48806 & n48808;
  assign n48812 = ~n61055 & ~n61056;
  assign n48813 = ~pi1134 & ~n48812;
  assign n48814 = ~pi699 & pi1135;
  assign n48815 = ~pi763 & ~pi1135;
  assign n48816 = pi1136 & ~n48815;
  assign n48817 = pi1136 & ~n48814;
  assign n48818 = ~n48815 & n48817;
  assign n48819 = ~n48814 & n48816;
  assign n48820 = pi871 & n47826;
  assign n48821 = pi1134 & ~n48820;
  assign n48822 = ~n61057 & n48821;
  assign n48823 = n47819 & ~n48822;
  assign n48824 = ~n48813 & n48823;
  assign n48825 = ~n48799 & ~n48824;
  assign n48826 = pi199 & ~pi1062;
  assign n48827 = ~pi199 & ~pi258;
  assign n48828 = ~n47686 & ~n48827;
  assign n48829 = ~n47686 & ~n48826;
  assign n48830 = ~n48827 & n48829;
  assign n48831 = ~n48826 & n48828;
  assign n48832 = pi364 & n47790;
  assign n48833 = pi391 & pi591;
  assign n48834 = ~pi592 & n48833;
  assign n48835 = ~n48832 & ~n48834;
  assign n48836 = ~pi590 & ~n48835;
  assign n48837 = pi343 & n47683;
  assign n48838 = ~pi588 & ~n48837;
  assign n48839 = ~n48836 & n48838;
  assign n48840 = pi415 & n5089;
  assign n48841 = pi588 & ~n48840;
  assign n48842 = n47686 & ~n48841;
  assign n48843 = ~n48839 & n48842;
  assign n48844 = ~n61058 & ~n48843;
  assign n48845 = n5138 & ~n48844;
  assign n48846 = ~pi612 & ~pi1135;
  assign n48847 = pi695 & pi1135;
  assign n48848 = ~pi1134 & ~n48847;
  assign n48849 = ~pi1134 & ~n48846;
  assign n48850 = ~n48847 & n48849;
  assign n48851 = ~n48846 & n48848;
  assign n48852 = n48112 & n61059;
  assign n48853 = pi745 & n47662;
  assign n48854 = pi723 & pi1135;
  assign n48855 = ~pi852 & ~pi1136;
  assign n48856 = ~n48854 & ~n48855;
  assign n48857 = n47666 & n48856;
  assign n48858 = ~n48853 & n48857;
  assign n48859 = ~n48852 & ~n48858;
  assign n48860 = ~n5138 & ~n48859;
  assign n48861 = ~n48845 & ~n48860;
  assign n48862 = pi199 & ~pi1040;
  assign n48863 = ~pi199 & ~pi261;
  assign n48864 = ~n47686 & ~n48863;
  assign n48865 = ~n47686 & ~n48862;
  assign n48866 = ~n48863 & n48865;
  assign n48867 = ~n48862 & n48864;
  assign n48868 = pi447 & n47790;
  assign n48869 = pi333 & pi591;
  assign n48870 = ~pi592 & n48869;
  assign n48871 = ~n48868 & ~n48870;
  assign n48872 = ~pi590 & ~n48871;
  assign n48873 = pi327 & n47683;
  assign n48874 = ~pi588 & ~n48873;
  assign n48875 = ~n48872 & n48874;
  assign n48876 = pi453 & n5089;
  assign n48877 = pi588 & ~n48876;
  assign n48878 = n47686 & ~n48877;
  assign n48879 = ~n48875 & n48878;
  assign n48880 = ~n61060 & ~n48879;
  assign n48881 = n5138 & ~n48880;
  assign n48882 = ~pi611 & ~pi1135;
  assign n48883 = pi646 & pi1135;
  assign n48884 = ~pi1134 & ~n48883;
  assign n48885 = ~pi1134 & ~n48882;
  assign n48886 = ~n48883 & n48885;
  assign n48887 = ~n48882 & n48884;
  assign n48888 = n48112 & n61061;
  assign n48889 = pi741 & n47662;
  assign n48890 = pi724 & pi1135;
  assign n48891 = ~pi865 & ~pi1136;
  assign n48892 = ~n48890 & ~n48891;
  assign n48893 = n47666 & n48892;
  assign n48894 = ~n48889 & n48893;
  assign n48895 = ~n48888 & ~n48894;
  assign n48896 = ~n5138 & ~n48895;
  assign n48897 = ~n48881 & ~n48896;
  assign n48898 = pi199 & ~pi1069;
  assign n48899 = ~pi199 & ~pi259;
  assign n48900 = ~n47686 & ~n48899;
  assign n48901 = ~n47686 & ~n48898;
  assign n48902 = ~n48899 & n48901;
  assign n48903 = ~n48898 & n48900;
  assign n48904 = pi366 & n47790;
  assign n48905 = pi335 & pi591;
  assign n48906 = ~pi592 & n48905;
  assign n48907 = ~n48904 & ~n48906;
  assign n48908 = ~pi590 & ~n48907;
  assign n48909 = pi344 & n47683;
  assign n48910 = ~pi588 & ~n48909;
  assign n48911 = ~n48908 & n48910;
  assign n48912 = pi416 & n5089;
  assign n48913 = pi588 & ~n48912;
  assign n48914 = n47686 & ~n48913;
  assign n48915 = ~n48911 & n48914;
  assign n48916 = ~n61062 & ~n48915;
  assign n48917 = n5138 & ~n48916;
  assign n48918 = ~pi620 & ~pi1135;
  assign n48919 = pi635 & pi1135;
  assign n48920 = ~pi1134 & ~n48919;
  assign n48921 = ~pi1134 & ~n48918;
  assign n48922 = ~n48919 & n48921;
  assign n48923 = ~n48918 & n48920;
  assign n48924 = n48112 & n61063;
  assign n48925 = pi742 & n47662;
  assign n48926 = pi704 & pi1135;
  assign n48927 = ~pi870 & ~pi1136;
  assign n48928 = ~n48926 & ~n48927;
  assign n48929 = n47666 & n48928;
  assign n48930 = ~n48925 & n48929;
  assign n48931 = ~n48924 & ~n48930;
  assign n48932 = ~n5138 & ~n48931;
  assign n48933 = ~n48917 & ~n48932;
  assign n48934 = pi199 & ~pi1067;
  assign n48935 = ~pi199 & ~pi260;
  assign n48936 = ~n47686 & ~n48935;
  assign n48937 = ~n47686 & ~n48934;
  assign n48938 = ~n48935 & n48937;
  assign n48939 = ~n48934 & n48936;
  assign n48940 = pi368 & n47790;
  assign n48941 = pi393 & pi591;
  assign n48942 = ~pi592 & n48941;
  assign n48943 = ~n48940 & ~n48942;
  assign n48944 = ~pi590 & ~n48943;
  assign n48945 = pi346 & n47683;
  assign n48946 = ~pi588 & ~n48945;
  assign n48947 = ~n48944 & n48946;
  assign n48948 = pi418 & n5089;
  assign n48949 = pi588 & ~n48948;
  assign n48950 = n47686 & ~n48949;
  assign n48951 = ~n48947 & n48950;
  assign n48952 = ~n61064 & ~n48951;
  assign n48953 = n5138 & ~n48952;
  assign n48954 = ~pi613 & ~pi1135;
  assign n48955 = pi632 & pi1135;
  assign n48956 = ~pi1134 & ~n48955;
  assign n48957 = ~pi1134 & ~n48954;
  assign n48958 = ~n48955 & n48957;
  assign n48959 = ~n48954 & n48956;
  assign n48960 = n48112 & n61065;
  assign n48961 = pi760 & n47662;
  assign n48962 = pi688 & pi1135;
  assign n48963 = ~pi856 & ~pi1136;
  assign n48964 = ~n48962 & ~n48963;
  assign n48965 = n47666 & n48964;
  assign n48966 = ~n48961 & n48965;
  assign n48967 = ~n48960 & ~n48966;
  assign n48968 = ~n5138 & ~n48967;
  assign n48969 = ~n48953 & ~n48968;
  assign n48970 = pi199 & ~pi1039;
  assign n48971 = ~pi199 & ~pi251;
  assign n48972 = ~n47686 & ~n48971;
  assign n48973 = ~n47686 & ~n48970;
  assign n48974 = ~n48971 & n48973;
  assign n48975 = ~n48970 & n48972;
  assign n48976 = pi367 & n47790;
  assign n48977 = pi392 & pi591;
  assign n48978 = ~pi592 & n48977;
  assign n48979 = ~n48976 & ~n48978;
  assign n48980 = ~pi590 & ~n48979;
  assign n48981 = pi345 & n47683;
  assign n48982 = ~pi588 & ~n48981;
  assign n48983 = ~n48980 & n48982;
  assign n48984 = pi417 & n5089;
  assign n48985 = pi588 & ~n48984;
  assign n48986 = n47686 & ~n48985;
  assign n48987 = ~n48983 & n48986;
  assign n48988 = ~n61066 & ~n48987;
  assign n48989 = n5138 & ~n48988;
  assign n48990 = ~pi610 & ~pi1135;
  assign n48991 = pi631 & pi1135;
  assign n48992 = ~pi1134 & ~n48991;
  assign n48993 = ~pi1134 & ~n48990;
  assign n48994 = ~n48991 & n48993;
  assign n48995 = ~n48990 & n48992;
  assign n48996 = n48112 & n61067;
  assign n48997 = pi757 & n47662;
  assign n48998 = pi686 & pi1135;
  assign n48999 = ~pi848 & ~pi1136;
  assign n49000 = ~n48998 & ~n48999;
  assign n49001 = n47666 & n49000;
  assign n49002 = ~n48997 & n49001;
  assign n49003 = ~n48996 & ~n49002;
  assign n49004 = ~n5138 & ~n49003;
  assign n49005 = ~n48989 & ~n49004;
  assign n49006 = pi897 & n36719;
  assign n49007 = ~pi476 & n45424;
  assign n49008 = ~n49006 & ~n49007;
  assign n49009 = ~n61023 & ~n49008;
  assign n49010 = pi251 & n49008;
  assign n49011 = ~n49009 & ~n49010;
  assign n49012 = ~n61000 & ~n49008;
  assign n49013 = pi255 & n49008;
  assign n49014 = n61000 & ~n49008;
  assign n49015 = ~pi255 & n49008;
  assign n49016 = ~n49014 & ~n49015;
  assign n49017 = ~n49012 & ~n49013;
  assign n49018 = ~n61029 & ~n49008;
  assign n49019 = pi256 & n49008;
  assign n49020 = n61029 & ~n49008;
  assign n49021 = ~pi256 & n49008;
  assign n49022 = ~n49020 & ~n49021;
  assign n49023 = ~n49018 & ~n49019;
  assign n49024 = ~n61003 & ~n49008;
  assign n49025 = pi257 & n49008;
  assign n49026 = n61003 & ~n49008;
  assign n49027 = ~pi257 & n49008;
  assign n49028 = ~n49026 & ~n49027;
  assign n49029 = ~n49024 & ~n49025;
  assign n49030 = ~n61035 & ~n49008;
  assign n49031 = pi258 & n49008;
  assign n49032 = n61035 & ~n49008;
  assign n49033 = ~pi258 & n49008;
  assign n49034 = ~n49032 & ~n49033;
  assign n49035 = ~n49030 & ~n49031;
  assign n49036 = ~n61042 & ~n49008;
  assign n49037 = pi259 & n49008;
  assign n49038 = n61042 & ~n49008;
  assign n49039 = ~pi259 & n49008;
  assign n49040 = ~n49038 & ~n49039;
  assign n49041 = ~n49036 & ~n49037;
  assign n49042 = ~n60996 & ~n49008;
  assign n49043 = pi260 & n49008;
  assign n49044 = ~n49042 & ~n49043;
  assign n49045 = ~n61039 & ~n49008;
  assign n49046 = pi261 & n49008;
  assign n49047 = ~n49045 & ~n49046;
  assign n49048 = ~pi476 & pi1048;
  assign n49049 = pi290 & pi476;
  assign n49050 = ~pi290 & pi476;
  assign n49051 = ~pi476 & ~pi1048;
  assign n49052 = ~n49050 & ~n49051;
  assign n49053 = ~n49048 & ~n49049;
  assign n49054 = ~pi476 & pi1049;
  assign n49055 = pi291 & pi476;
  assign n49056 = ~pi291 & pi476;
  assign n49057 = ~pi476 & ~pi1049;
  assign n49058 = ~n49056 & ~n49057;
  assign n49059 = ~n49054 & ~n49055;
  assign n49060 = ~pi476 & pi1084;
  assign n49061 = pi292 & pi476;
  assign n49062 = ~pi292 & pi476;
  assign n49063 = ~pi476 & ~pi1084;
  assign n49064 = ~n49062 & ~n49063;
  assign n49065 = ~n49060 & ~n49061;
  assign n49066 = ~pi476 & pi1059;
  assign n49067 = pi293 & pi476;
  assign n49068 = ~pi293 & pi476;
  assign n49069 = ~pi476 & ~pi1059;
  assign n49070 = ~n49068 & ~n49069;
  assign n49071 = ~n49066 & ~n49067;
  assign n49072 = ~pi476 & pi1072;
  assign n49073 = pi294 & pi476;
  assign n49074 = ~pi294 & pi476;
  assign n49075 = ~pi476 & ~pi1072;
  assign n49076 = ~n49074 & ~n49075;
  assign n49077 = ~n49072 & ~n49073;
  assign n49078 = ~pi476 & pi1053;
  assign n49079 = pi295 & pi476;
  assign n49080 = ~pi295 & pi476;
  assign n49081 = ~pi476 & ~pi1053;
  assign n49082 = ~n49080 & ~n49081;
  assign n49083 = ~n49078 & ~n49079;
  assign n49084 = ~pi476 & pi1037;
  assign n49085 = pi296 & pi476;
  assign n49086 = ~pi296 & pi476;
  assign n49087 = ~pi476 & ~pi1037;
  assign n49088 = ~n49086 & ~n49087;
  assign n49089 = ~n49084 & ~n49085;
  assign n49090 = ~pi476 & pi1044;
  assign n49091 = pi297 & pi476;
  assign n49092 = ~pi297 & pi476;
  assign n49093 = ~pi476 & ~pi1044;
  assign n49094 = ~n49092 & ~n49093;
  assign n49095 = ~n49090 & ~n49091;
  assign n49096 = pi375 & n48155;
  assign n49097 = pi399 & pi591;
  assign n49098 = n48157 & n49097;
  assign n49099 = ~n49096 & ~n49098;
  assign n49100 = ~pi590 & ~n49099;
  assign n49101 = pi316 & n47686;
  assign n49102 = n47683 & n49101;
  assign n49103 = ~n49100 & ~n49102;
  assign n49104 = ~pi588 & ~n49103;
  assign n49105 = ~pi200 & ~pi308;
  assign n49106 = pi200 & ~pi1037;
  assign n49107 = ~n49105 & ~n49106;
  assign n49108 = pi200 & pi1037;
  assign n49109 = ~pi200 & pi308;
  assign n49110 = ~pi199 & ~n49109;
  assign n49111 = ~n49108 & n49110;
  assign n49112 = ~pi199 & ~n49107;
  assign n49113 = pi199 & ~pi1047;
  assign n49114 = ~n47686 & ~n49113;
  assign n49115 = ~n61081 & n49114;
  assign n49116 = pi424 & n47973;
  assign n49117 = n48177 & n49116;
  assign n49118 = n5138 & ~n49117;
  assign n49119 = ~n49115 & n49118;
  assign n49120 = ~n49104 & n49119;
  assign n49121 = pi777 & n47662;
  assign n49122 = pi737 & pi1135;
  assign n49123 = ~pi838 & ~pi1136;
  assign n49124 = ~n49122 & ~n49123;
  assign n49125 = pi1134 & ~n49122;
  assign n49126 = ~n49123 & n49125;
  assign n49127 = n48187 & n49126;
  assign n49128 = n47666 & n49124;
  assign n49129 = ~n49121 & n61082;
  assign n49130 = ~pi619 & ~pi1135;
  assign n49131 = ~pi648 & pi1135;
  assign n49132 = ~pi1134 & ~n49131;
  assign n49133 = ~pi1134 & ~n49130;
  assign n49134 = ~n49131 & n49133;
  assign n49135 = ~n49130 & n49132;
  assign n49136 = n48112 & n61083;
  assign n49137 = ~n5138 & ~n49136;
  assign n49138 = ~n49129 & n49137;
  assign po890 = ~n49120 & ~n49138;
  assign n49140 = ~n58992 & ~n46791;
  assign n49141 = ~n46783 & n49140;
  assign n49142 = pi219 & ~n47489;
  assign n49143 = ~pi219 & n46198;
  assign n49144 = ~n49142 & ~n49143;
  assign n49145 = n58992 & ~n49144;
  assign n49146 = ~pi219 & ~n46218;
  assign n49147 = ~n46166 & ~n49146;
  assign n49148 = n49145 & n49147;
  assign n49149 = ~n49141 & ~n49148;
  assign n49150 = ~pi1151 & ~n49149;
  assign n49151 = ~n47250 & n49140;
  assign n49152 = ~n46180 & n49142;
  assign n49153 = ~n46183 & n47549;
  assign n49154 = ~n49152 & ~n49153;
  assign n49155 = n58992 & ~n49154;
  assign n49156 = ~n49151 & ~n49155;
  assign n49157 = pi1151 & ~n49156;
  assign n49158 = ~pi268 & ~n49157;
  assign n49159 = ~n49150 & n49158;
  assign n49160 = ~n58992 & ~n46780;
  assign n49161 = ~n47366 & n49160;
  assign n49162 = pi219 & ~n46930;
  assign n49163 = ~n47526 & ~n49162;
  assign n49164 = n46177 & ~n49163;
  assign n49165 = n58992 & ~n49164;
  assign n49166 = ~n49161 & ~n49165;
  assign n49167 = pi1151 & ~n49166;
  assign n49168 = ~n47248 & n49160;
  assign n49169 = n58992 & ~n47564;
  assign n49170 = ~n49162 & n49169;
  assign n49171 = ~n49168 & ~n49170;
  assign n49172 = ~pi1151 & ~n49171;
  assign n49173 = pi268 & ~n49172;
  assign n49174 = ~n49167 & n49173;
  assign n49175 = ~pi1150 & ~n49174;
  assign n49176 = ~n49159 & n49175;
  assign n49177 = ~n47249 & n49160;
  assign n49178 = ~n46281 & ~n47564;
  assign n49179 = ~n49154 & ~n49178;
  assign n49180 = n58992 & ~n49179;
  assign n49181 = ~n46190 & ~n47198;
  assign n49182 = n49180 & ~n49181;
  assign n49183 = ~n49177 & ~n49182;
  assign n49184 = ~pi1151 & ~n49183;
  assign n49185 = n58992 & ~n46929;
  assign n49186 = ~n46146 & n49185;
  assign n49187 = ~n47060 & n49160;
  assign n49188 = n58992 & ~n47560;
  assign n49189 = pi219 & n46327;
  assign n49190 = n49188 & ~n49189;
  assign n49191 = ~n49187 & ~n49190;
  assign n49192 = ~n49186 & n49191;
  assign n49193 = pi1151 & ~n49192;
  assign n49194 = pi268 & ~n49193;
  assign n49195 = ~n49184 & n49194;
  assign n49196 = ~n47271 & n49140;
  assign n49197 = pi219 & ~n46191;
  assign n49198 = ~n47526 & ~n49197;
  assign n49199 = ~n46182 & ~n49198;
  assign n49200 = ~n47283 & ~n49199;
  assign n49201 = n58992 & ~n49200;
  assign n49202 = ~n49196 & ~n49201;
  assign n49203 = ~pi1151 & ~n49202;
  assign n49204 = ~n49168 & n49196;
  assign n49205 = ~n49151 & ~n49204;
  assign n49206 = ~n49145 & n49205;
  assign n49207 = pi1151 & ~n49206;
  assign n49208 = ~pi268 & ~n49207;
  assign n49209 = ~n49203 & n49208;
  assign n49210 = pi1150 & ~n49209;
  assign n49211 = ~n49195 & n49210;
  assign n49212 = ~n49176 & ~n49211;
  assign n49213 = pi1152 & ~n49212;
  assign n49214 = pi219 & ~n58992;
  assign n49215 = ~n46190 & n49214;
  assign n49216 = ~n47251 & ~n49215;
  assign n49217 = ~n49180 & n49216;
  assign n49218 = pi1151 & n49217;
  assign n49219 = ~n46234 & n49188;
  assign n49220 = ~n46783 & ~n49215;
  assign n49221 = ~n49219 & n49220;
  assign n49222 = ~pi1151 & n49221;
  assign n49223 = ~pi268 & ~n49222;
  assign n49224 = ~n49218 & n49223;
  assign n49225 = n58992 & ~n47529;
  assign n49226 = ~n47526 & n49225;
  assign n49227 = ~n47539 & ~n49226;
  assign n49228 = pi1151 & ~n49227;
  assign n49229 = ~n47060 & n47538;
  assign n49230 = ~n49190 & ~n49229;
  assign n49231 = n46150 & ~n49230;
  assign n49232 = ~pi1151 & n49231;
  assign n49233 = pi268 & ~n49232;
  assign n49234 = ~n49228 & n49233;
  assign n49235 = ~n49224 & ~n49234;
  assign n49236 = ~pi1150 & ~n49235;
  assign n49237 = n58992 & ~n46244;
  assign n49238 = n49199 & n49237;
  assign n49239 = ~n49204 & ~n49238;
  assign n49240 = ~pi1151 & n49239;
  assign n49241 = ~n46150 & ~n49230;
  assign n49242 = ~n49221 & ~n49241;
  assign n49243 = pi1151 & n49242;
  assign n49244 = ~pi268 & ~n49243;
  assign n49245 = pi1151 & ~n49242;
  assign n49246 = ~pi1151 & ~n49239;
  assign n49247 = ~n49245 & ~n49246;
  assign n49248 = ~pi268 & ~n49247;
  assign n49249 = ~n49240 & n49244;
  assign n49250 = ~n47249 & n47538;
  assign n49251 = n49154 & n49185;
  assign n49252 = ~n49250 & ~n49251;
  assign n49253 = ~pi1151 & n49252;
  assign n49254 = pi1151 & n49230;
  assign n49255 = pi268 & ~n49254;
  assign n49256 = ~pi1151 & ~n49252;
  assign n49257 = pi1151 & ~n49230;
  assign n49258 = ~n49256 & ~n49257;
  assign n49259 = pi268 & ~n49258;
  assign n49260 = ~n49253 & n49255;
  assign n49261 = pi1150 & ~n61085;
  assign n49262 = ~n61084 & n49261;
  assign n49263 = ~pi1152 & ~n49262;
  assign n49264 = ~n49236 & n49263;
  assign n49265 = ~n61084 & ~n61085;
  assign n49266 = ~pi1152 & ~n49265;
  assign n49267 = pi1152 & ~n49209;
  assign n49268 = ~n49195 & n49267;
  assign n49269 = ~n49266 & ~n49268;
  assign n49270 = pi1150 & ~n49269;
  assign n49271 = pi1152 & ~n49157;
  assign n49272 = pi1152 & ~n49150;
  assign n49273 = ~n49157 & n49272;
  assign n49274 = ~n49150 & n49271;
  assign n49275 = ~pi1152 & ~n49222;
  assign n49276 = ~n49218 & n49275;
  assign n49277 = ~n61086 & ~n49276;
  assign n49278 = ~pi268 & ~n49277;
  assign n49279 = pi1151 & n49166;
  assign n49280 = ~pi1151 & n49171;
  assign n49281 = pi1152 & ~n49280;
  assign n49282 = ~n49279 & n49281;
  assign n49283 = pi1151 & n49227;
  assign n49284 = ~pi1151 & ~n49231;
  assign n49285 = ~pi1152 & ~n49284;
  assign n49286 = ~n49283 & n49285;
  assign n49287 = pi268 & ~n49286;
  assign n49288 = ~n49282 & n49287;
  assign n49289 = ~pi1150 & ~n49288;
  assign n49290 = ~n49278 & n49289;
  assign n49291 = ~n49270 & ~n49290;
  assign n49292 = ~n49213 & ~n49264;
  assign n49293 = n46439 & ~n61087;
  assign n49294 = pi268 & pi1152;
  assign n49295 = ~pi219 & ~n44774;
  assign n49296 = ~pi199 & n44774;
  assign n49297 = ~n49295 & ~n49296;
  assign n49298 = ~pi211 & ~n44774;
  assign n49299 = n58992 & n46389;
  assign n49300 = ~n49298 & ~n49299;
  assign n49301 = pi1152 & ~n49300;
  assign n49302 = n49297 & ~n49301;
  assign n49303 = ~pi1151 & n49300;
  assign n49304 = pi1150 & ~n49303;
  assign n49305 = ~pi1152 & n49297;
  assign n49306 = pi1151 & ~n49297;
  assign n49307 = n49300 & ~n49306;
  assign n49308 = pi1150 & ~n49307;
  assign n49309 = ~n49305 & n49308;
  assign n49310 = ~n49302 & n49304;
  assign n49311 = ~n49294 & n61088;
  assign n49312 = ~n44774 & n47344;
  assign n49313 = n58992 & n46736;
  assign n49314 = ~n44774 & ~n47344;
  assign n49315 = n44774 & ~n46348;
  assign n49316 = ~n36719 & n61089;
  assign n49317 = ~n49314 & ~n49316;
  assign n49318 = ~n49312 & ~n49313;
  assign n49319 = pi1151 & n61090;
  assign n49320 = pi1152 & n49319;
  assign n49321 = n58992 & ~n45428;
  assign n49322 = ~n45499 & ~n49321;
  assign n49323 = pi1151 & ~n49322;
  assign n49324 = ~pi1152 & ~n49323;
  assign n49325 = ~pi1151 & n47419;
  assign n49326 = ~pi1150 & ~n49325;
  assign n49327 = ~n49324 & n49326;
  assign n49328 = ~n49320 & n49327;
  assign n49329 = ~n49311 & ~n49328;
  assign n49330 = pi1091 & ~n49329;
  assign n49331 = pi1152 & n61088;
  assign n49332 = pi1152 & n49308;
  assign n49333 = pi1091 & ~n61091;
  assign n49334 = pi268 & ~n49333;
  assign n49335 = ~n49330 & ~n49334;
  assign n49336 = ~n46439 & ~n49335;
  assign n49337 = ~pi230 & ~n49336;
  assign n49338 = ~n49293 & n49337;
  assign n49339 = pi230 & ~n61088;
  assign n49340 = ~n49328 & n49339;
  assign po425 = ~n49338 & ~n49340;
  assign po1102 = pi230 & n2794;
  assign n49343 = ~pi212 & ~pi214;
  assign n49344 = ~pi211 & ~n49343;
  assign n49345 = pi219 & ~n49344;
  assign n49346 = ~n58992 & ~n49345;
  assign n49347 = pi1142 & ~n36624;
  assign n49348 = pi211 & pi1143;
  assign n49349 = ~pi211 & pi1144;
  assign n49350 = ~n49348 & ~n49349;
  assign n49351 = ~pi212 & pi214;
  assign n49352 = pi212 & ~pi214;
  assign n49353 = ~n49351 & ~n49352;
  assign n49354 = ~n36621 & ~n49343;
  assign n49355 = ~n36621 & ~n49350;
  assign n49356 = ~n49343 & n49355;
  assign n49357 = ~n49350 & ~n61092;
  assign n49358 = ~pi211 & pi1143;
  assign n49359 = n36621 & n49358;
  assign n49360 = ~n61093 & ~n49359;
  assign n49361 = ~pi219 & ~n49360;
  assign n49362 = ~n49347 & ~n49361;
  assign n49363 = n49346 & ~n49362;
  assign n49364 = pi199 & pi1142;
  assign n49365 = ~pi200 & ~n49364;
  assign n49366 = ~pi199 & pi1144;
  assign n49367 = n49365 & ~n49366;
  assign n49368 = ~pi199 & pi1143;
  assign n49369 = pi200 & ~n49368;
  assign n49370 = ~n49367 & ~n49369;
  assign n49371 = ~pi299 & ~n49370;
  assign n49372 = ~pi207 & ~n49371;
  assign n49373 = n49365 & ~n49368;
  assign n49374 = pi207 & ~pi299;
  assign n49375 = ~pi199 & pi1142;
  assign n49376 = pi200 & ~n49375;
  assign n49377 = n49374 & ~n49376;
  assign n49378 = ~n49373 & n49377;
  assign n49379 = ~n49372 & ~n49378;
  assign n49380 = pi208 & ~n49379;
  assign n49381 = pi207 & ~pi208;
  assign n49382 = n49370 & n49381;
  assign n49383 = ~n49380 & ~n49382;
  assign n49384 = ~pi299 & ~n49383;
  assign n49385 = pi211 & pi1142;
  assign n49386 = n36621 & n49385;
  assign n49387 = ~n49359 & ~n49386;
  assign n49388 = ~n49355 & n49387;
  assign n49389 = ~pi219 & n49388;
  assign n49390 = ~pi211 & pi1142;
  assign n49391 = pi219 & ~n49390;
  assign n49392 = pi299 & ~n49343;
  assign n49393 = ~n49391 & n49392;
  assign n49394 = ~n49389 & n49393;
  assign n49395 = ~n49384 & ~n49394;
  assign n49396 = pi299 & ~n49350;
  assign n49397 = ~n49384 & ~n49396;
  assign n49398 = ~pi214 & ~n49384;
  assign n49399 = ~pi212 & ~n49398;
  assign n49400 = ~n49397 & n49399;
  assign n49401 = ~n49396 & n49398;
  assign n49402 = ~n49358 & ~n49385;
  assign n49403 = pi299 & ~n49402;
  assign n49404 = pi214 & ~n49403;
  assign n49405 = ~n49384 & n49404;
  assign n49406 = pi212 & ~n49405;
  assign n49407 = ~n49401 & n49406;
  assign n49408 = ~pi219 & ~n49407;
  assign n49409 = ~n49400 & n49408;
  assign n49410 = ~pi299 & n49383;
  assign n49411 = pi299 & ~pi1142;
  assign n49412 = n49344 & ~n49411;
  assign n49413 = ~n49410 & n49412;
  assign n49414 = ~n49344 & n49384;
  assign n49415 = pi219 & ~n49414;
  assign n49416 = ~n49413 & n49415;
  assign n49417 = n58992 & ~n49416;
  assign n49418 = ~n49409 & n49417;
  assign n49419 = n58992 & ~n49395;
  assign n49420 = ~n49363 & ~n61094;
  assign n49421 = pi213 & n49420;
  assign n49422 = ~n46550 & ~n46553;
  assign n49423 = ~pi214 & n49422;
  assign n49424 = ~n46444 & ~n47022;
  assign n49425 = pi214 & n49424;
  assign n49426 = pi212 & ~n49425;
  assign n49427 = ~pi214 & ~n49422;
  assign n49428 = pi214 & ~n49424;
  assign n49429 = ~n49427 & ~n49428;
  assign n49430 = pi212 & ~n49429;
  assign n49431 = pi212 & ~n49423;
  assign n49432 = ~n49425 & n49431;
  assign n49433 = ~n49423 & n49426;
  assign n49434 = ~n46291 & ~n46443;
  assign n49435 = pi214 & ~n49434;
  assign n49436 = ~pi212 & n49435;
  assign n49437 = n49351 & ~n49434;
  assign n49438 = ~pi219 & ~n61096;
  assign n49439 = ~pi212 & ~n49435;
  assign n49440 = pi212 & n49429;
  assign n49441 = ~n49439 & ~n49440;
  assign n49442 = ~n61095 & ~n61096;
  assign n49443 = ~pi219 & ~n61097;
  assign n49444 = ~n61095 & n49438;
  assign n49445 = ~pi211 & pi214;
  assign n49446 = pi1155 & n49445;
  assign n49447 = ~pi212 & ~n49446;
  assign n49448 = ~pi214 & ~n46552;
  assign n49449 = n36621 & ~n47068;
  assign n49450 = ~n49448 & ~n49449;
  assign n49451 = ~n49447 & n49450;
  assign n49452 = pi219 & ~n49451;
  assign n49453 = ~n58992 & ~n49452;
  assign n49454 = ~n61098 & n49453;
  assign n49455 = ~pi213 & ~n49454;
  assign n49456 = n47414 & n61097;
  assign n49457 = n46506 & n49351;
  assign n49458 = pi299 & pi1154;
  assign n49459 = ~pi214 & n49458;
  assign n49460 = pi214 & pi299;
  assign n49461 = pi1153 & n49460;
  assign n49462 = ~n49459 & ~n49461;
  assign n49463 = ~pi214 & ~n49458;
  assign n49464 = pi299 & pi1153;
  assign n49465 = pi214 & ~n49464;
  assign n49466 = pi212 & ~n49465;
  assign n49467 = ~n49463 & n49466;
  assign n49468 = pi212 & ~n49463;
  assign n49469 = ~n49465 & n49468;
  assign n49470 = pi212 & ~n49462;
  assign n49471 = ~n49457 & ~n61099;
  assign n49472 = n36681 & ~n49471;
  assign n49473 = ~n49456 & ~n49472;
  assign n49474 = ~n49384 & n49473;
  assign n49475 = n58992 & ~n49474;
  assign n49476 = n49455 & ~n49475;
  assign n49477 = pi209 & ~n49476;
  assign n49478 = ~n49421 & n49477;
  assign n49479 = pi199 & n47015;
  assign n49480 = pi1155 & n46359;
  assign n49481 = ~pi299 & n61100;
  assign n49482 = pi1155 & n46360;
  assign n49483 = ~pi1156 & ~n61101;
  assign n49484 = pi199 & ~pi1155;
  assign n49485 = ~pi200 & ~pi1155;
  assign n49486 = n46499 & ~n49485;
  assign n49487 = n46499 & ~n49484;
  assign n49488 = ~n49483 & n61102;
  assign n49489 = pi207 & n49488;
  assign n49490 = ~pi208 & ~n49489;
  assign n49491 = pi1154 & ~n47154;
  assign n49492 = n45518 & n47015;
  assign n49493 = pi1154 & n46498;
  assign n49494 = ~n47429 & n49493;
  assign n49495 = ~n49492 & ~n49494;
  assign n49496 = n49491 & ~n49495;
  assign n49497 = ~pi199 & ~pi1155;
  assign n49498 = ~pi1154 & ~n49497;
  assign n49499 = n47425 & n49498;
  assign n49500 = pi1155 & ~n47422;
  assign n49501 = ~pi1155 & n46360;
  assign n49502 = n45521 & n49485;
  assign n49503 = pi1153 & n61103;
  assign n49504 = ~n49500 & ~n49503;
  assign n49505 = ~pi1154 & ~n49504;
  assign n49506 = ~n46756 & ~n47446;
  assign n49507 = pi1154 & ~n49506;
  assign n49508 = ~n49505 & ~n49507;
  assign n49509 = ~pi299 & ~n49508;
  assign n49510 = ~n49496 & ~n49499;
  assign n49511 = pi207 & n61104;
  assign n49512 = pi1156 & n45518;
  assign n49513 = pi1156 & n46522;
  assign n49514 = ~n46497 & n49512;
  assign n49515 = ~n46521 & n46538;
  assign n49516 = ~n61105 & ~n49515;
  assign n49517 = ~pi207 & ~n49516;
  assign n49518 = pi208 & ~n49517;
  assign n49519 = pi207 & ~n61104;
  assign n49520 = ~pi207 & n49516;
  assign n49521 = ~n49519 & ~n49520;
  assign n49522 = pi208 & ~n49521;
  assign n49523 = ~n49511 & n49518;
  assign n49524 = ~n49490 & ~n61106;
  assign n49525 = ~pi1157 & ~n49524;
  assign n49526 = pi1156 & ~n49484;
  assign n49527 = n46999 & n49526;
  assign n49528 = ~pi1156 & n46389;
  assign n49529 = ~pi1156 & ~n49484;
  assign n49530 = n46389 & n49529;
  assign n49531 = ~n49484 & n49528;
  assign n49532 = ~n49527 & ~n61107;
  assign n49533 = pi207 & ~n49532;
  assign n49534 = ~pi208 & ~n49533;
  assign n49535 = ~n61106 & ~n49534;
  assign n49536 = pi1157 & ~n49535;
  assign n49537 = ~n49525 & ~n49536;
  assign n49538 = pi211 & ~n49537;
  assign n49539 = ~pi214 & ~n49537;
  assign n49540 = ~pi212 & ~n49539;
  assign n49541 = pi207 & n49508;
  assign n49542 = ~pi207 & ~n46506;
  assign n49543 = n49516 & n49542;
  assign n49544 = pi208 & ~n49543;
  assign n49545 = ~n49541 & n49544;
  assign n49546 = pi1155 & ~n46365;
  assign n49547 = ~n45518 & ~n49546;
  assign n49548 = pi1156 & ~n49547;
  assign n49549 = n46500 & ~n46738;
  assign n49550 = ~n49548 & ~n49549;
  assign n49551 = pi207 & n49550;
  assign n49552 = ~pi208 & pi1157;
  assign n49553 = ~pi208 & ~n49542;
  assign n49554 = pi1157 & n49553;
  assign n49555 = ~n49542 & n49552;
  assign n49556 = ~n49551 & n61108;
  assign n49557 = ~pi299 & n49483;
  assign n49558 = ~n46736 & ~n47101;
  assign n49559 = ~n49557 & n49558;
  assign n49560 = n49553 & n49559;
  assign n49561 = ~n49556 & ~n49560;
  assign n49562 = ~n49545 & n49561;
  assign n49563 = n49445 & n49562;
  assign n49564 = n49540 & ~n49563;
  assign n49565 = ~pi211 & ~pi214;
  assign n49566 = pi1154 & ~n60931;
  assign n49567 = n49516 & ~n49566;
  assign n49568 = ~pi207 & ~n49567;
  assign n49569 = ~pi299 & n49506;
  assign n49570 = pi1154 & ~n49569;
  assign n49571 = ~n49499 & ~n49570;
  assign n49572 = pi207 & ~n49571;
  assign n49573 = ~n49568 & ~n49572;
  assign n49574 = pi208 & ~n49573;
  assign n49575 = ~n46754 & ~n49546;
  assign n49576 = ~pi1156 & ~n49575;
  assign n49577 = pi1156 & ~n47016;
  assign n49578 = ~n49576 & ~n49577;
  assign n49579 = ~n49527 & n49575;
  assign n49580 = pi207 & n61109;
  assign n49581 = ~pi207 & ~pi299;
  assign n49582 = ~pi208 & ~n49581;
  assign n49583 = ~n49580 & n49582;
  assign n49584 = pi299 & ~pi1154;
  assign n49585 = pi1157 & ~n49584;
  assign n49586 = n49583 & n49585;
  assign n49587 = ~n49458 & ~n49489;
  assign n49588 = ~pi208 & ~n49587;
  assign n49589 = ~pi1157 & n49588;
  assign n49590 = ~n49586 & ~n49589;
  assign n49591 = ~n49574 & n49590;
  assign n49592 = n49565 & n49591;
  assign n49593 = pi1157 & ~n49583;
  assign n49594 = pi1156 & ~n61100;
  assign n49595 = n46705 & n49594;
  assign n49596 = ~n49483 & ~n49595;
  assign n49597 = pi207 & n49596;
  assign n49598 = ~pi299 & ~n49597;
  assign n49599 = ~pi208 & ~n49598;
  assign n49600 = ~pi1157 & ~n49599;
  assign n49601 = ~n49593 & ~n49600;
  assign n49602 = pi299 & ~pi1153;
  assign n49603 = ~n49600 & ~n49602;
  assign n49604 = ~n49593 & n49603;
  assign n49605 = n49601 & ~n49602;
  assign n49606 = pi1153 & ~n46422;
  assign n49607 = n49495 & ~n49606;
  assign n49608 = pi207 & ~n49607;
  assign n49609 = ~n46754 & ~n46756;
  assign n49610 = pi1156 & ~n49609;
  assign n49611 = pi299 & ~pi1155;
  assign n49612 = ~n46706 & ~n49611;
  assign n49613 = ~pi299 & ~n46735;
  assign n49614 = ~n49610 & n61111;
  assign n49615 = ~n49566 & ~n49610;
  assign n49616 = n61111 & n49615;
  assign n49617 = ~n49566 & n49614;
  assign n49618 = ~pi207 & ~n49602;
  assign n49619 = ~n61112 & n49618;
  assign n49620 = ~n49608 & ~n49619;
  assign n49621 = pi208 & ~n49620;
  assign n49622 = n49445 & ~n49621;
  assign n49623 = ~n61110 & n49622;
  assign n49624 = pi212 & ~n49623;
  assign n49625 = pi212 & ~n49592;
  assign n49626 = ~n49623 & n49625;
  assign n49627 = ~n49592 & n49624;
  assign n49628 = ~n49564 & ~n61113;
  assign n49629 = ~n49538 & ~n49628;
  assign n49630 = pi219 & ~n49629;
  assign n49631 = ~pi1154 & ~pi1156;
  assign n49632 = ~n61111 & n49631;
  assign n49633 = ~pi207 & ~n49566;
  assign n49634 = ~n49632 & n49633;
  assign n49635 = ~pi207 & n61112;
  assign n49636 = ~n49610 & n49634;
  assign n49637 = n49374 & n49508;
  assign n49638 = n49374 & n49607;
  assign n49639 = pi208 & ~n61115;
  assign n49640 = ~n61114 & n49639;
  assign n49641 = n49593 & ~n49640;
  assign n49642 = ~pi211 & ~n49641;
  assign n49643 = ~pi211 & ~n49525;
  assign n49644 = ~n49641 & n49643;
  assign n49645 = ~n49525 & n49642;
  assign n49646 = pi299 & pi1156;
  assign n49647 = pi207 & ~n49646;
  assign n49648 = ~n49515 & ~n49610;
  assign n49649 = ~pi207 & n49648;
  assign n49650 = ~pi207 & ~n49648;
  assign n49651 = pi207 & n49646;
  assign n49652 = ~n49650 & ~n49651;
  assign n49653 = ~n49647 & ~n49649;
  assign n49654 = ~n49511 & n61117;
  assign n49655 = pi208 & ~n49654;
  assign n49656 = ~n49483 & n49599;
  assign n49657 = ~n49533 & ~n49646;
  assign n49658 = n49552 & ~n49657;
  assign n49659 = ~n49656 & ~n49658;
  assign n49660 = ~n49655 & n49659;
  assign n49661 = pi211 & ~n49660;
  assign n49662 = pi214 & ~n49661;
  assign n49663 = ~n61116 & n49662;
  assign n49664 = n49540 & ~n49663;
  assign n49665 = n36620 & ~n49591;
  assign n49666 = ~n36620 & ~n49565;
  assign n49667 = ~n49562 & n49666;
  assign n49668 = n49565 & ~n49660;
  assign n49669 = ~n49667 & ~n49668;
  assign n49670 = ~n49665 & n49669;
  assign n49671 = pi212 & ~n49670;
  assign n49672 = ~pi219 & ~n49671;
  assign n49673 = ~n49664 & n49672;
  assign n49674 = n58992 & ~n49673;
  assign n49675 = ~n49630 & n49674;
  assign n49676 = n49455 & ~n49675;
  assign n49677 = pi299 & ~pi1143;
  assign n49678 = n46737 & ~n49677;
  assign n49679 = pi299 & pi1143;
  assign n49680 = ~pi1155 & n49679;
  assign n49681 = pi1154 & ~n61103;
  assign n49682 = ~n49680 & n49681;
  assign n49683 = ~n49678 & n49682;
  assign n49684 = n46521 & ~n49679;
  assign n49685 = ~pi1156 & ~n49684;
  assign n49686 = ~n49683 & n49685;
  assign n49687 = ~n49609 & ~n49677;
  assign n49688 = ~pi1154 & ~n49687;
  assign n49689 = pi1154 & ~n46509;
  assign n49690 = ~n49679 & n49689;
  assign n49691 = pi1156 & ~n49690;
  assign n49692 = ~n49688 & n49691;
  assign n49693 = ~n49686 & ~n49692;
  assign n49694 = ~pi207 & n49693;
  assign n49695 = n49519 & ~n49679;
  assign n49696 = pi208 & ~n49695;
  assign n49697 = pi208 & ~n49694;
  assign n49698 = ~n49695 & n49697;
  assign n49699 = ~n49694 & n49696;
  assign n49700 = ~pi1157 & n49599;
  assign n49701 = ~n49677 & n49700;
  assign n49702 = pi207 & ~n49677;
  assign n49703 = ~n61109 & n49702;
  assign n49704 = ~n49679 & ~n49703;
  assign n49705 = n49552 & ~n49704;
  assign n49706 = ~pi211 & n36621;
  assign n49707 = pi211 & ~n61092;
  assign n49708 = pi211 & n49351;
  assign n49709 = pi212 & n49666;
  assign n49710 = ~n49708 & ~n49709;
  assign n49711 = ~n49706 & ~n49707;
  assign n49712 = ~n49705 & ~n61119;
  assign n49713 = ~n49701 & n49712;
  assign n49714 = ~n61118 & n49713;
  assign n49715 = pi299 & pi1144;
  assign n49716 = n49519 & ~n49715;
  assign n49717 = pi299 & ~pi1144;
  assign n49718 = n46737 & ~n49717;
  assign n49719 = ~pi1155 & n49715;
  assign n49720 = n49681 & ~n49719;
  assign n49721 = ~n49718 & n49720;
  assign n49722 = n46521 & ~n49715;
  assign n49723 = ~pi1156 & ~n49722;
  assign n49724 = ~n49721 & n49723;
  assign n49725 = ~n49609 & ~n49717;
  assign n49726 = ~pi1154 & ~n49725;
  assign n49727 = n49689 & ~n49715;
  assign n49728 = pi1156 & ~n49727;
  assign n49729 = ~n49726 & n49728;
  assign n49730 = ~n49724 & ~n49729;
  assign n49731 = ~pi207 & n49730;
  assign n49732 = pi208 & ~n49731;
  assign n49733 = pi208 & ~n49716;
  assign n49734 = ~n49731 & n49733;
  assign n49735 = ~n49716 & n49732;
  assign n49736 = n49700 & ~n49717;
  assign n49737 = pi207 & ~n49717;
  assign n49738 = ~n61109 & n49737;
  assign n49739 = ~n49715 & ~n49738;
  assign n49740 = n49552 & ~n49739;
  assign n49741 = ~pi211 & ~n61092;
  assign n49742 = n36678 & ~n49343;
  assign n49743 = ~n49740 & n61121;
  assign n49744 = ~n49736 & n49743;
  assign n49745 = ~n61120 & n49744;
  assign n49746 = ~n49701 & ~n49705;
  assign n49747 = ~n61118 & n49746;
  assign n49748 = n49706 & n49747;
  assign n49749 = pi211 & ~n49747;
  assign n49750 = ~n49736 & ~n49740;
  assign n49751 = ~n61120 & n49750;
  assign n49752 = ~pi211 & ~n49751;
  assign n49753 = ~n61092 & ~n49752;
  assign n49754 = ~n61092 & ~n49749;
  assign n49755 = ~n49752 & n49754;
  assign n49756 = ~n49749 & n49753;
  assign n49757 = ~n49748 & ~n61122;
  assign n49758 = ~n49714 & ~n49745;
  assign n49759 = ~pi219 & ~n61123;
  assign n49760 = ~pi219 & ~n49343;
  assign n49761 = ~n49344 & ~n49760;
  assign n49762 = ~n49537 & n49761;
  assign n49763 = ~n49411 & ~n49600;
  assign n49764 = ~n49593 & n49763;
  assign n49765 = ~n49411 & n49601;
  assign n49766 = pi208 & ~n49411;
  assign n49767 = ~n61114 & n49766;
  assign n49768 = pi299 & pi1142;
  assign n49769 = pi207 & ~n49768;
  assign n49770 = ~n61104 & n49769;
  assign n49771 = ~n49411 & ~n49615;
  assign n49772 = ~n46520 & ~n49768;
  assign n49773 = n49631 & ~n49772;
  assign n49774 = ~pi207 & ~n49773;
  assign n49775 = ~n49771 & n49774;
  assign n49776 = pi208 & ~n49775;
  assign n49777 = ~n49770 & n49776;
  assign n49778 = ~n61115 & n49767;
  assign n49779 = ~n36624 & ~n49761;
  assign n49780 = ~n61125 & n49779;
  assign n49781 = ~n61124 & n49779;
  assign n49782 = ~n61125 & n49781;
  assign n49783 = ~n61124 & n49780;
  assign n49784 = n58992 & ~n61126;
  assign n49785 = n58992 & ~n49762;
  assign n49786 = ~n61126 & n49785;
  assign n49787 = ~n49762 & n49784;
  assign n49788 = ~n49759 & n61127;
  assign n49789 = pi213 & ~n49363;
  assign n49790 = ~n49788 & n49789;
  assign n49791 = ~pi209 & ~n49790;
  assign n49792 = ~n49676 & n49791;
  assign n49793 = ~n49478 & ~n49792;
  assign n49794 = pi230 & ~n49793;
  assign n49795 = ~pi230 & ~pi233;
  assign n49796 = ~n49794 & ~n49795;
  assign n49797 = ~pi211 & pi1145;
  assign n49798 = pi211 & pi1144;
  assign n49799 = ~n49797 & ~n49798;
  assign n49800 = ~n36621 & n49799;
  assign n49801 = n36621 & n49350;
  assign n49802 = ~n49343 & ~n49801;
  assign n49803 = ~n49343 & ~n49800;
  assign n49804 = ~n49801 & n49803;
  assign n49805 = ~n49800 & n49802;
  assign n49806 = ~pi219 & ~n61128;
  assign n49807 = pi219 & ~n49358;
  assign n49808 = n49346 & ~n49807;
  assign n49809 = ~n49806 & n49808;
  assign n49810 = n47414 & n61128;
  assign n49811 = pi199 & pi1143;
  assign n49812 = ~pi200 & ~n49811;
  assign n49813 = ~n49366 & n49812;
  assign n49814 = pi208 & n49374;
  assign n49815 = ~n49369 & n49814;
  assign n49816 = ~n49813 & n49815;
  assign n49817 = ~pi199 & pi1145;
  assign n49818 = n49812 & ~n49817;
  assign n49819 = ~pi207 & ~pi208;
  assign n49820 = ~n36320 & ~n49819;
  assign n49821 = pi200 & ~n49366;
  assign n49822 = n49820 & ~n49821;
  assign n49823 = ~n49818 & n49822;
  assign n49824 = ~n49816 & ~n49823;
  assign n49825 = ~pi299 & ~n49824;
  assign n49826 = pi219 & ~n49343;
  assign n49827 = pi299 & n49358;
  assign n49828 = ~pi211 & n49679;
  assign n49829 = pi299 & n49826;
  assign n49830 = n49358 & n49829;
  assign n49831 = n49826 & n61129;
  assign n49832 = ~n49825 & ~n61130;
  assign n49833 = ~n49810 & n49832;
  assign n49834 = n58992 & ~n49833;
  assign n49835 = ~n49809 & ~n49834;
  assign n49836 = pi213 & n49835;
  assign n49837 = pi214 & n49422;
  assign n49838 = ~pi214 & n49434;
  assign n49839 = pi212 & ~n49838;
  assign n49840 = pi214 & ~n49422;
  assign n49841 = ~pi214 & ~n49434;
  assign n49842 = ~n49840 & ~n49841;
  assign n49843 = pi212 & ~n49842;
  assign n49844 = ~n49837 & n49839;
  assign n49845 = ~pi211 & pi1158;
  assign n49846 = ~n46309 & ~n49845;
  assign n49847 = n49351 & ~n49846;
  assign n49848 = ~pi219 & ~n49847;
  assign n49849 = ~pi219 & ~n61131;
  assign n49850 = ~n49847 & n49849;
  assign n49851 = ~n61131 & n49848;
  assign n49852 = n46550 & n49351;
  assign n49853 = ~n58992 & n49852;
  assign n49854 = ~n47437 & ~n49853;
  assign n49855 = pi214 & n46552;
  assign n49856 = pi1155 & n49565;
  assign n49857 = ~n49855 & ~n49856;
  assign n49858 = pi212 & ~n58992;
  assign n49859 = pi214 & ~n46552;
  assign n49860 = ~pi214 & ~n46444;
  assign n49861 = pi212 & ~n49860;
  assign n49862 = pi212 & ~n49857;
  assign n49863 = ~n49859 & n49861;
  assign n49864 = ~n58992 & n61133;
  assign n49865 = ~n49857 & n49858;
  assign n49866 = n49854 & ~n61134;
  assign n49867 = ~n61132 & ~n49866;
  assign n49868 = ~pi213 & ~n49867;
  assign n49869 = n47414 & ~n61132;
  assign n49870 = n49351 & n49646;
  assign n49871 = ~pi214 & n46506;
  assign n49872 = pi1154 & n49460;
  assign n49873 = ~n49871 & ~n49872;
  assign n49874 = ~pi214 & ~n46506;
  assign n49875 = pi214 & ~n49458;
  assign n49876 = pi212 & ~n49875;
  assign n49877 = ~n49874 & n49876;
  assign n49878 = pi212 & ~n49874;
  assign n49879 = ~n49875 & n49878;
  assign n49880 = pi212 & ~n49873;
  assign n49881 = ~n49870 & ~n61135;
  assign n49882 = n36681 & ~n49881;
  assign n49883 = ~n49825 & ~n49882;
  assign n49884 = ~n49869 & n49883;
  assign n49885 = n58992 & ~n49884;
  assign n49886 = n49868 & ~n49885;
  assign n49887 = pi209 & ~n49886;
  assign n49888 = ~n49836 & n49887;
  assign n49889 = n46389 & n49381;
  assign n49890 = pi1158 & n45444;
  assign n49891 = ~pi199 & ~pi1158;
  assign n49892 = pi1156 & ~n49891;
  assign n49893 = ~pi1156 & ~n45444;
  assign n49894 = pi1158 & ~n49893;
  assign n49895 = ~n46511 & ~n49894;
  assign n49896 = ~n49890 & ~n49892;
  assign n49897 = n49889 & ~n61136;
  assign n49898 = pi207 & n49516;
  assign n49899 = ~pi207 & ~n49488;
  assign n49900 = pi208 & ~n49899;
  assign n49901 = ~n49898 & n49900;
  assign n49902 = ~n49897 & ~n49901;
  assign n49903 = ~pi1157 & ~n49902;
  assign n49904 = ~pi200 & ~pi1158;
  assign n49905 = ~pi199 & ~n49904;
  assign n49906 = ~n46514 & ~n49905;
  assign n49907 = ~pi1158 & ~n46499;
  assign n49908 = n46385 & ~n49907;
  assign n49909 = ~n49905 & ~n49908;
  assign n49910 = n49374 & ~n49909;
  assign n49911 = n49374 & ~n49906;
  assign n49912 = ~pi208 & n61137;
  assign n49913 = ~pi207 & n49532;
  assign n49914 = pi208 & ~n49913;
  assign n49915 = ~n49898 & n49914;
  assign n49916 = ~n49912 & ~n49915;
  assign n49917 = pi1157 & ~n49916;
  assign n49918 = ~n49903 & ~n49917;
  assign n49919 = ~pi214 & n49918;
  assign n49920 = ~pi212 & ~n49919;
  assign n49921 = ~pi299 & n49906;
  assign n49922 = n49582 & ~n49921;
  assign n49923 = pi207 & n61111;
  assign n49924 = pi207 & n49614;
  assign n49925 = ~n49610 & n49923;
  assign n49926 = n49615 & n49923;
  assign n49927 = ~n49566 & n61138;
  assign n49928 = ~pi207 & n61109;
  assign n49929 = pi208 & ~n49928;
  assign n49930 = ~n61139 & n49929;
  assign n49931 = ~n49922 & ~n49930;
  assign n49932 = pi1157 & ~n49931;
  assign n49933 = ~n49903 & ~n49932;
  assign n49934 = pi211 & n49933;
  assign n49935 = pi1158 & n61112;
  assign n49936 = ~pi1158 & n49516;
  assign n49937 = pi207 & ~n49936;
  assign n49938 = ~n49935 & n49937;
  assign n49939 = ~pi299 & ~n49596;
  assign n49940 = pi299 & ~pi1158;
  assign n49941 = ~pi207 & ~n49940;
  assign n49942 = ~n49939 & n49941;
  assign n49943 = pi208 & ~n49942;
  assign n49944 = ~n49938 & n49943;
  assign n49945 = pi207 & ~n36720;
  assign n49946 = ~pi299 & ~n49945;
  assign n49947 = pi1158 & ~n49946;
  assign n49948 = n46514 & n49374;
  assign n49949 = ~pi208 & ~n49948;
  assign n49950 = ~n49947 & n49949;
  assign n49951 = ~pi1157 & ~n49950;
  assign n49952 = ~n49944 & n49951;
  assign n49953 = pi208 & pi1157;
  assign n49954 = ~pi207 & ~n61109;
  assign n49955 = ~n49940 & n49954;
  assign n49956 = ~n49938 & ~n49955;
  assign n49957 = n49953 & ~n49956;
  assign n49958 = pi1157 & ~n49890;
  assign n49959 = ~n46501 & n49958;
  assign n49960 = pi207 & ~n49959;
  assign n49961 = ~n49947 & ~n49960;
  assign n49962 = n49552 & ~n49961;
  assign n49963 = ~pi211 & ~n49962;
  assign n49964 = ~n49957 & n49963;
  assign n49965 = ~n49952 & n49963;
  assign n49966 = ~n49957 & n49965;
  assign n49967 = ~n49952 & n49964;
  assign n49968 = ~n49934 & ~n61140;
  assign n49969 = pi214 & ~n49968;
  assign n49970 = n49920 & ~n49969;
  assign n49971 = ~pi207 & n49559;
  assign n49972 = ~n46506 & n49516;
  assign n49973 = pi207 & ~n49972;
  assign n49974 = ~n49971 & ~n49973;
  assign n49975 = pi208 & ~n49974;
  assign n49976 = ~pi208 & n46506;
  assign n49977 = ~n49897 & ~n49976;
  assign n49978 = ~n49975 & n49977;
  assign n49979 = ~pi1157 & ~n49978;
  assign n49980 = ~pi207 & ~n49550;
  assign n49981 = ~n49973 & ~n49980;
  assign n49982 = n49953 & ~n49981;
  assign n49983 = ~n46506 & ~n61137;
  assign n49984 = n49552 & ~n49983;
  assign n49985 = ~n49982 & ~n49984;
  assign n49986 = ~n49979 & n49985;
  assign n49987 = n36620 & ~n49986;
  assign n49988 = n49565 & ~n49933;
  assign n49989 = pi207 & ~n49648;
  assign n49990 = ~pi207 & n49596;
  assign n49991 = pi208 & ~n49990;
  assign n49992 = ~n49989 & n49991;
  assign n49993 = ~pi208 & ~n49646;
  assign n49994 = ~pi200 & pi207;
  assign n49995 = ~n61136 & n49994;
  assign n49996 = n49993 & ~n49995;
  assign n49997 = ~pi1157 & ~n49996;
  assign n49998 = ~n49992 & n49997;
  assign n49999 = ~n61107 & ~n49577;
  assign n50000 = ~pi207 & ~n49999;
  assign n50001 = ~n49989 & ~n50000;
  assign n50002 = n49953 & ~n50001;
  assign n50003 = ~n49646 & ~n61137;
  assign n50004 = n49552 & ~n50003;
  assign n50005 = ~n50002 & ~n50004;
  assign n50006 = ~n49998 & n50005;
  assign n50007 = n49666 & ~n50006;
  assign n50008 = ~n49988 & ~n50007;
  assign n50009 = ~n49987 & ~n50007;
  assign n50010 = ~n49988 & n50009;
  assign n50011 = ~n49987 & n50008;
  assign n50012 = pi212 & ~n61141;
  assign n50013 = ~pi219 & ~n50012;
  assign n50014 = ~n49970 & n50013;
  assign n50015 = ~n49344 & n49918;
  assign n50016 = n49351 & n50006;
  assign n50017 = ~pi214 & ~n49986;
  assign n50018 = ~n49584 & n49954;
  assign n50019 = pi1157 & ~n50018;
  assign n50020 = pi1154 & ~n49595;
  assign n50021 = ~n61102 & ~n50020;
  assign n50022 = ~pi207 & ~n49557;
  assign n50023 = ~n50021 & n50022;
  assign n50024 = ~pi1157 & ~n49897;
  assign n50025 = ~n50023 & n50024;
  assign n50026 = ~n50019 & ~n50025;
  assign n50027 = pi207 & ~n49567;
  assign n50028 = pi208 & ~n50027;
  assign n50029 = ~n50026 & n50028;
  assign n50030 = n61137 & ~n50024;
  assign n50031 = ~pi208 & ~n49458;
  assign n50032 = ~n50030 & n50031;
  assign n50033 = pi214 & ~n50032;
  assign n50034 = ~n50029 & n50033;
  assign n50035 = pi212 & ~n50034;
  assign n50036 = ~n50017 & n50035;
  assign n50037 = ~n50016 & ~n50036;
  assign n50038 = ~pi211 & ~n50037;
  assign n50039 = ~n50015 & ~n50038;
  assign n50040 = pi219 & ~n50039;
  assign n50041 = n58992 & ~n50040;
  assign n50042 = ~n50014 & n50041;
  assign n50043 = n49868 & ~n50042;
  assign n50044 = pi299 & ~pi1145;
  assign n50045 = ~n60931 & ~n50044;
  assign n50046 = pi1154 & ~n50045;
  assign n50047 = pi299 & pi1145;
  assign n50048 = n46521 & ~n50047;
  assign n50049 = ~pi1156 & ~n50048;
  assign n50050 = ~n50046 & n50049;
  assign n50051 = ~n49609 & ~n50044;
  assign n50052 = ~pi1154 & ~n50051;
  assign n50053 = n49689 & ~n50047;
  assign n50054 = pi1156 & ~n50053;
  assign n50055 = ~n50052 & n50054;
  assign n50056 = ~n50050 & ~n50055;
  assign n50057 = pi207 & ~n50056;
  assign n50058 = ~pi199 & n46485;
  assign n50059 = n49939 & ~n50058;
  assign n50060 = ~pi207 & ~n50044;
  assign n50061 = ~n50059 & n50060;
  assign n50062 = pi208 & ~n50061;
  assign n50063 = ~n50057 & n50062;
  assign n50064 = ~pi299 & n46514;
  assign n50065 = n46389 & n46511;
  assign n50066 = ~pi1157 & ~n61142;
  assign n50067 = ~pi1157 & ~n49890;
  assign n50068 = ~n61142 & n50067;
  assign n50069 = ~n49890 & n50066;
  assign n50070 = n49960 & ~n61143;
  assign n50071 = ~pi208 & ~n50047;
  assign n50072 = ~n50070 & n50071;
  assign n50073 = ~n50063 & ~n50072;
  assign n50074 = ~pi211 & ~n50073;
  assign n50075 = ~pi1157 & ~n49995;
  assign n50076 = ~pi208 & ~n50075;
  assign n50077 = n61137 & n50076;
  assign n50078 = n49912 & ~n50024;
  assign n50079 = ~pi208 & ~n61144;
  assign n50080 = ~n49715 & n50079;
  assign n50081 = pi207 & ~n49730;
  assign n50082 = ~pi207 & ~n49717;
  assign n50083 = ~n50059 & n50082;
  assign n50084 = pi208 & ~n50083;
  assign n50085 = ~n50081 & n50084;
  assign n50086 = ~n50080 & ~n50085;
  assign n50087 = pi211 & ~n50086;
  assign n50088 = ~n50074 & ~n50087;
  assign n50089 = ~pi214 & ~n50088;
  assign n50090 = ~n49679 & n50079;
  assign n50091 = pi207 & ~n49693;
  assign n50092 = ~pi207 & ~n49677;
  assign n50093 = ~n50059 & n50092;
  assign n50094 = pi208 & ~n50093;
  assign n50095 = ~n50091 & n50094;
  assign n50096 = ~n50090 & ~n50095;
  assign n50097 = pi211 & n50096;
  assign n50098 = ~pi211 & n50086;
  assign n50099 = pi214 & ~n50098;
  assign n50100 = ~n50097 & n50099;
  assign n50101 = pi212 & ~n50100;
  assign n50102 = ~n50089 & n50101;
  assign n50103 = pi214 & ~n50088;
  assign n50104 = n49920 & ~n50103;
  assign n50105 = ~pi219 & ~n50104;
  assign n50106 = ~pi219 & ~n50102;
  assign n50107 = ~n50104 & n50106;
  assign n50108 = ~n50102 & n50105;
  assign n50109 = n49344 & ~n50096;
  assign n50110 = ~n50015 & ~n50109;
  assign n50111 = pi219 & ~n50110;
  assign n50112 = n58992 & ~n50111;
  assign n50113 = ~n61145 & n50112;
  assign n50114 = pi213 & ~n49809;
  assign n50115 = ~n50113 & n50114;
  assign n50116 = ~pi209 & ~n50115;
  assign n50117 = ~n50043 & n50116;
  assign n50118 = ~n49888 & ~n50117;
  assign n50119 = pi230 & ~n50118;
  assign n50120 = ~pi230 & ~pi237;
  assign n50121 = ~n50119 & ~n50120;
  assign n50122 = pi1150 & ~n49192;
  assign n50123 = ~pi1150 & ~n49183;
  assign n50124 = ~n50122 & ~n50123;
  assign n50125 = pi1151 & ~n50124;
  assign n50126 = ~pi1150 & ~n49252;
  assign n50127 = pi1150 & ~n49230;
  assign n50128 = ~n50126 & ~n50127;
  assign n50129 = ~pi1151 & ~n50128;
  assign n50130 = pi275 & ~n50129;
  assign n50131 = ~n50125 & n50130;
  assign n50132 = pi1151 & ~n49202;
  assign n50133 = ~n49246 & ~n50132;
  assign n50134 = ~pi1150 & ~n50133;
  assign n50135 = ~pi1151 & ~n49242;
  assign n50136 = ~n49207 & ~n50135;
  assign n50137 = pi1150 & ~n50136;
  assign n50138 = ~pi275 & ~n50137;
  assign n50139 = ~n50134 & n50138;
  assign n50140 = pi1149 & ~n50139;
  assign n50141 = ~n50131 & n50140;
  assign n50142 = ~pi1150 & n49149;
  assign n50143 = pi1150 & n49156;
  assign n50144 = pi1151 & ~n50143;
  assign n50145 = ~n50142 & n50144;
  assign n50146 = pi1150 & ~n49217;
  assign n50147 = ~pi1150 & ~n49221;
  assign n50148 = ~pi1151 & ~n50147;
  assign n50149 = ~n50146 & n50148;
  assign n50150 = ~pi275 & ~n50149;
  assign n50151 = ~n50145 & n50150;
  assign n50152 = pi1150 & n49166;
  assign n50153 = ~pi1150 & n49171;
  assign n50154 = pi1151 & ~n50153;
  assign n50155 = ~n50152 & n50154;
  assign n50156 = pi1150 & n49227;
  assign n50157 = ~pi1150 & ~n49231;
  assign n50158 = ~pi1151 & ~n50157;
  assign n50159 = ~n50156 & n50158;
  assign n50160 = pi275 & ~n50159;
  assign n50161 = ~n50155 & n50160;
  assign n50162 = ~pi1149 & ~n50161;
  assign n50163 = ~n50151 & n50162;
  assign n50164 = n46438 & ~n50163;
  assign n50165 = ~n50141 & n50164;
  assign n50166 = ~pi1151 & n45887;
  assign n50167 = pi1149 & ~n49300;
  assign n50168 = ~n50166 & n50167;
  assign n50169 = ~pi1149 & pi1151;
  assign n50170 = ~n47419 & n50169;
  assign n50171 = ~n50168 & ~n50170;
  assign n50172 = ~pi1150 & ~n50171;
  assign n50173 = n58992 & n46999;
  assign n50174 = ~pi1149 & n49319;
  assign n50175 = pi1151 & ~n49300;
  assign n50176 = pi1149 & n49297;
  assign n50177 = ~n50175 & n50176;
  assign n50178 = pi1150 & ~n50177;
  assign n50179 = ~n50174 & n50178;
  assign n50180 = pi1091 & ~n50179;
  assign n50181 = ~n50174 & ~n50177;
  assign n50182 = pi1150 & ~n50181;
  assign n50183 = ~pi1150 & ~n50170;
  assign n50184 = ~n50168 & n50183;
  assign n50185 = ~n50182 & ~n50184;
  assign n50186 = pi1091 & ~n50185;
  assign n50187 = ~n50172 & n50180;
  assign n50188 = ~n44774 & n47341;
  assign n50189 = n58992 & n46397;
  assign n50190 = ~n50188 & ~n50189;
  assign n50191 = ~pi1149 & pi1150;
  assign n50192 = ~pi1151 & n50191;
  assign n50193 = ~n50190 & n50192;
  assign n50194 = pi275 & ~n50193;
  assign n50195 = ~n61146 & n50194;
  assign n50196 = ~pi1151 & n49322;
  assign n50197 = pi1150 & ~n50196;
  assign n50198 = ~n49319 & n50197;
  assign n50199 = ~pi1150 & pi1151;
  assign n50200 = ~n47419 & n50199;
  assign n50201 = ~pi1149 & ~n50200;
  assign n50202 = ~n50198 & n50201;
  assign n50203 = pi1149 & ~pi1150;
  assign n50204 = n49300 & n50203;
  assign n50205 = ~n50177 & ~n50204;
  assign n50206 = ~n50202 & n50205;
  assign n50207 = ~pi275 & pi1091;
  assign n50208 = n50206 & n50207;
  assign n50209 = ~n46438 & ~n50208;
  assign n50210 = ~n50195 & n50209;
  assign n50211 = ~n61146 & ~n50193;
  assign n50212 = pi275 & ~n50211;
  assign n50213 = pi1091 & n50206;
  assign n50214 = ~pi275 & ~n50213;
  assign n50215 = ~n46438 & ~n50214;
  assign n50216 = ~n50212 & n50215;
  assign n50217 = ~n50145 & ~n50149;
  assign n50218 = ~pi275 & ~n50217;
  assign n50219 = ~n50152 & ~n50153;
  assign n50220 = pi1151 & ~n50219;
  assign n50221 = ~n50156 & ~n50157;
  assign n50222 = ~pi1151 & ~n50221;
  assign n50223 = pi275 & ~n50222;
  assign n50224 = ~n50220 & n50223;
  assign n50225 = ~pi1149 & ~n50224;
  assign n50226 = ~n50218 & n50225;
  assign n50227 = pi1151 & ~n49183;
  assign n50228 = ~pi1150 & ~n49256;
  assign n50229 = ~n50227 & n50228;
  assign n50230 = ~pi1151 & ~n49230;
  assign n50231 = pi1150 & ~n50230;
  assign n50232 = ~n49193 & n50231;
  assign n50233 = pi275 & ~n50232;
  assign n50234 = ~n50229 & n50233;
  assign n50235 = ~pi1150 & ~n49202;
  assign n50236 = pi1150 & ~n49206;
  assign n50237 = pi1151 & ~n50236;
  assign n50238 = ~n50235 & n50237;
  assign n50239 = ~pi1150 & ~n49239;
  assign n50240 = pi1150 & ~n49242;
  assign n50241 = ~pi1151 & ~n50240;
  assign n50242 = ~n50239 & n50241;
  assign n50243 = ~pi275 & ~n50242;
  assign n50244 = ~n50238 & n50243;
  assign n50245 = pi1149 & ~n50244;
  assign n50246 = ~n50234 & n50245;
  assign n50247 = n46438 & ~n50246;
  assign n50248 = n46438 & ~n50226;
  assign n50249 = ~n50246 & n50248;
  assign n50250 = ~n50226 & n50247;
  assign n50251 = ~n50216 & ~n61147;
  assign n50252 = ~n50165 & ~n50210;
  assign n50253 = ~pi230 & n61148;
  assign n50254 = pi230 & ~n50206;
  assign n50255 = ~pi230 & ~n61148;
  assign n50256 = pi230 & n50206;
  assign n50257 = ~n50255 & ~n50256;
  assign n50258 = ~n50253 & ~n50254;
  assign n50259 = pi1150 & ~n49183;
  assign n50260 = ~pi1149 & ~n50126;
  assign n50261 = ~n50259 & n50260;
  assign n50262 = ~pi1150 & ~n49230;
  assign n50263 = pi1149 & ~n50262;
  assign n50264 = ~n50122 & n50263;
  assign n50265 = pi1150 & n49192;
  assign n50266 = ~pi1150 & n49230;
  assign n50267 = pi1149 & ~n50266;
  assign n50268 = ~n50265 & n50267;
  assign n50269 = pi1150 & n49183;
  assign n50270 = ~pi1150 & n49252;
  assign n50271 = ~pi1149 & ~n50270;
  assign n50272 = ~n50269 & n50271;
  assign n50273 = ~n50268 & ~n50272;
  assign n50274 = ~n50261 & ~n50264;
  assign n50275 = pi1148 & ~n61150;
  assign n50276 = ~pi1150 & n49227;
  assign n50277 = pi1149 & ~n50276;
  assign n50278 = ~n50152 & n50277;
  assign n50279 = pi1150 & n49171;
  assign n50280 = ~pi1149 & ~n50157;
  assign n50281 = ~n50279 & n50280;
  assign n50282 = ~n50278 & ~n50281;
  assign n50283 = ~pi1148 & ~n50282;
  assign n50284 = pi283 & ~n50283;
  assign n50285 = pi1148 & n61150;
  assign n50286 = ~pi1148 & ~n50281;
  assign n50287 = ~n50278 & n50286;
  assign n50288 = ~n50285 & ~n50287;
  assign n50289 = pi283 & ~n50288;
  assign n50290 = ~n50275 & n50284;
  assign n50291 = pi1091 & n61090;
  assign n50292 = pi1150 & ~n50291;
  assign n50293 = ~pi1150 & n50190;
  assign n50294 = ~pi1148 & pi1149;
  assign n50295 = ~n50293 & n50294;
  assign n50296 = ~n50292 & n50295;
  assign n50297 = ~pi1150 & n45887;
  assign n50298 = ~n49300 & ~n50297;
  assign n50299 = ~pi1149 & ~n50298;
  assign n50300 = ~n49300 & ~n50203;
  assign n50301 = n49297 & ~n50300;
  assign n50302 = pi1148 & ~n50301;
  assign n50303 = ~n49295 & ~n49298;
  assign n50304 = ~n49295 & ~n61089;
  assign n50305 = ~n49298 & n50304;
  assign n50306 = ~n61089 & n50303;
  assign n50307 = pi1150 & ~n61152;
  assign n50308 = pi1149 & ~n50307;
  assign n50309 = n49297 & n50308;
  assign n50310 = pi1148 & ~n50299;
  assign n50311 = ~n50309 & n50310;
  assign n50312 = ~n50299 & n50302;
  assign n50313 = pi1150 & ~n47419;
  assign n50314 = ~pi1149 & ~n50313;
  assign n50315 = ~pi1148 & ~n50314;
  assign n50316 = pi1091 & ~n50315;
  assign n50317 = ~n61153 & n50316;
  assign n50318 = ~n50296 & ~n50317;
  assign n50319 = pi1149 & ~n50293;
  assign n50320 = ~n50292 & n50319;
  assign n50321 = pi1091 & n50314;
  assign n50322 = ~pi1148 & ~n50321;
  assign n50323 = ~n50320 & n50322;
  assign n50324 = ~n50299 & ~n50301;
  assign n50325 = pi1091 & ~n50324;
  assign n50326 = pi1148 & ~n50325;
  assign n50327 = ~pi283 & ~n50326;
  assign n50328 = ~n50323 & n50327;
  assign n50329 = ~pi283 & ~n50323;
  assign n50330 = ~n50326 & n50329;
  assign n50331 = ~pi283 & ~n50318;
  assign n50332 = pi272 & ~n61154;
  assign n50333 = ~n61151 & n50332;
  assign n50334 = pi1150 & n49149;
  assign n50335 = ~pi1149 & ~n50147;
  assign n50336 = ~n50334 & n50335;
  assign n50337 = ~pi1150 & ~n49217;
  assign n50338 = pi1149 & ~n50143;
  assign n50339 = ~n50337 & n50338;
  assign n50340 = ~n50336 & ~n50339;
  assign n50341 = ~pi1148 & ~n50340;
  assign n50342 = pi1150 & ~n49202;
  assign n50343 = ~pi1149 & ~n50239;
  assign n50344 = ~n50342 & n50343;
  assign n50345 = ~pi1150 & ~n49242;
  assign n50346 = pi1149 & ~n50345;
  assign n50347 = ~n50236 & n50346;
  assign n50348 = pi1148 & ~n50347;
  assign n50349 = ~n50344 & n50348;
  assign n50350 = pi283 & ~n50349;
  assign n50351 = ~n50344 & ~n50347;
  assign n50352 = pi1148 & ~n50351;
  assign n50353 = ~pi1148 & ~n50336;
  assign n50354 = ~n50339 & n50353;
  assign n50355 = ~n50352 & ~n50354;
  assign n50356 = pi283 & ~n50355;
  assign n50357 = ~n50341 & n50350;
  assign n50358 = pi1091 & n61153;
  assign n50359 = pi1150 & ~n61090;
  assign n50360 = ~pi1150 & ~n49322;
  assign n50361 = pi1149 & ~n50360;
  assign n50362 = pi1149 & n61090;
  assign n50363 = ~n50308 & ~n50362;
  assign n50364 = ~n50360 & ~n50363;
  assign n50365 = ~n50359 & n50361;
  assign n50366 = pi1091 & ~n61156;
  assign n50367 = pi1091 & n50315;
  assign n50368 = ~n61156 & n50367;
  assign n50369 = n50315 & n50366;
  assign n50370 = ~pi283 & ~n61157;
  assign n50371 = ~n50358 & n50370;
  assign n50372 = ~pi272 & ~n50371;
  assign n50373 = ~n61155 & n50372;
  assign n50374 = ~pi230 & ~n50373;
  assign n50375 = ~pi230 & ~n50333;
  assign n50376 = ~n50373 & n50375;
  assign n50377 = ~n50333 & n50374;
  assign n50378 = n50315 & ~n61156;
  assign n50379 = pi230 & ~n61153;
  assign n50380 = ~n50378 & n50379;
  assign po429 = ~n61158 & ~n50380;
  assign n50382 = ~pi1147 & ~n49217;
  assign n50383 = pi1147 & n49242;
  assign n50384 = ~pi1149 & ~n50383;
  assign n50385 = ~n50382 & n50384;
  assign n50386 = ~pi1147 & n49156;
  assign n50387 = pi1147 & n49206;
  assign n50388 = pi1149 & ~n50387;
  assign n50389 = ~n50386 & n50388;
  assign n50390 = pi1148 & ~n50389;
  assign n50391 = ~n50385 & n50390;
  assign n50392 = pi1147 & n49202;
  assign n50393 = ~pi1147 & n49149;
  assign n50394 = pi1149 & ~n50393;
  assign n50395 = ~n50392 & n50394;
  assign n50396 = pi1147 & n49239;
  assign n50397 = ~pi1147 & ~n49221;
  assign n50398 = ~pi1149 & ~n50397;
  assign n50399 = ~n50396 & n50398;
  assign n50400 = ~pi1148 & ~n50399;
  assign n50401 = ~n50395 & n50400;
  assign n50402 = ~pi283 & ~n50401;
  assign n50403 = ~n50391 & n50402;
  assign n50404 = pi1147 & n49183;
  assign n50405 = ~pi1147 & n49171;
  assign n50406 = ~pi1148 & ~n50405;
  assign n50407 = ~n50404 & n50406;
  assign n50408 = ~pi1147 & n49166;
  assign n50409 = pi1147 & n49192;
  assign n50410 = pi1148 & ~n50409;
  assign n50411 = ~n50408 & n50410;
  assign n50412 = pi1149 & ~n50411;
  assign n50413 = ~n50407 & n50412;
  assign n50414 = pi1147 & n49252;
  assign n50415 = ~pi1147 & ~n49231;
  assign n50416 = ~pi1148 & ~n50415;
  assign n50417 = ~n50414 & n50416;
  assign n50418 = ~pi1147 & n49227;
  assign n50419 = pi1147 & n49230;
  assign n50420 = pi1148 & ~n50419;
  assign n50421 = ~n50418 & n50420;
  assign n50422 = ~pi1149 & ~n50421;
  assign n50423 = ~n50417 & n50422;
  assign n50424 = pi283 & ~n50423;
  assign n50425 = ~n50413 & n50424;
  assign n50426 = ~pi230 & ~n50425;
  assign n50427 = ~n50385 & ~n50389;
  assign n50428 = pi1148 & ~n50427;
  assign n50429 = ~n50395 & ~n50399;
  assign n50430 = ~pi1148 & ~n50429;
  assign n50431 = ~pi283 & ~n50430;
  assign n50432 = ~n50428 & n50431;
  assign n50433 = pi1147 & ~n49183;
  assign n50434 = ~pi1147 & ~n49171;
  assign n50435 = ~pi1148 & ~n50434;
  assign n50436 = ~n50433 & n50435;
  assign n50437 = ~pi1147 & ~n49166;
  assign n50438 = pi1147 & ~n49192;
  assign n50439 = pi1148 & ~n50438;
  assign n50440 = ~n50437 & n50439;
  assign n50441 = pi1149 & ~n50440;
  assign n50442 = ~n50436 & n50441;
  assign n50443 = pi1147 & ~n49252;
  assign n50444 = ~pi1147 & n49231;
  assign n50445 = ~pi1148 & ~n50444;
  assign n50446 = ~n50443 & n50445;
  assign n50447 = ~pi1147 & ~n49227;
  assign n50448 = pi1147 & ~n49230;
  assign n50449 = pi1148 & ~n50448;
  assign n50450 = ~n50447 & n50449;
  assign n50451 = ~pi1149 & ~n50450;
  assign n50452 = ~n50446 & n50451;
  assign n50453 = pi283 & ~n50452;
  assign n50454 = ~n50442 & n50453;
  assign n50455 = ~n50432 & ~n50454;
  assign n50456 = ~pi230 & ~n50455;
  assign n50457 = ~n50403 & n50426;
  assign n50458 = pi1147 & ~n45887;
  assign n50459 = n50362 & ~n50458;
  assign n50460 = pi1147 & ~n49297;
  assign n50461 = ~pi1149 & n49322;
  assign n50462 = ~n50460 & n50461;
  assign n50463 = pi1148 & ~n50462;
  assign n50464 = pi1148 & ~n50459;
  assign n50465 = ~n50462 & n50464;
  assign n50466 = ~n50459 & n50463;
  assign n50467 = pi1149 & ~n47419;
  assign n50468 = ~n50458 & ~n50467;
  assign n50469 = ~pi1148 & ~n50468;
  assign n50470 = pi230 & ~n50469;
  assign n50471 = ~n61160 & n50470;
  assign po440 = ~n61159 & ~n50471;
  assign n50473 = pi1153 & ~n49565;
  assign n50474 = ~n49445 & ~n49448;
  assign n50475 = ~n50473 & ~n50474;
  assign n50476 = pi212 & ~n50475;
  assign n50477 = ~n46552 & ~n47143;
  assign n50478 = n49351 & ~n50477;
  assign n50479 = ~pi219 & ~n50478;
  assign n50480 = ~n50476 & n50479;
  assign n50481 = n49346 & ~n50480;
  assign n50482 = pi1152 & ~n50481;
  assign n50483 = ~n36320 & n49516;
  assign n50484 = ~pi1154 & ~n49492;
  assign n50485 = ~pi199 & n49485;
  assign n50486 = ~n60908 & n46999;
  assign n50487 = ~n50484 & n50486;
  assign n50488 = pi207 & n50487;
  assign n50489 = ~n49820 & ~n50488;
  assign n50490 = ~n50483 & ~n50489;
  assign n50491 = ~pi214 & ~n50490;
  assign n50492 = ~pi212 & ~n50491;
  assign n50493 = ~pi207 & n49458;
  assign n50494 = ~n50027 & ~n50493;
  assign n50495 = ~pi208 & ~n50494;
  assign n50496 = ~pi299 & ~n46350;
  assign n50497 = ~n50484 & ~n50496;
  assign n50498 = pi207 & n50497;
  assign n50499 = ~n49568 & ~n50498;
  assign n50500 = pi208 & ~n50499;
  assign n50501 = ~n50495 & ~n50500;
  assign n50502 = ~pi211 & ~n50501;
  assign n50503 = n49582 & ~n61139;
  assign n50504 = n49374 & ~n50497;
  assign n50505 = pi208 & ~n50504;
  assign n50506 = ~n61114 & n50505;
  assign n50507 = ~n50503 & ~n50506;
  assign n50508 = ~n49602 & ~n50507;
  assign n50509 = pi211 & n50508;
  assign n50510 = ~n50502 & ~n50509;
  assign n50511 = pi214 & n50510;
  assign n50512 = n50492 & ~n50511;
  assign n50513 = ~pi219 & ~n50512;
  assign n50514 = ~pi214 & ~n50510;
  assign n50515 = ~pi211 & ~pi1153;
  assign n50516 = pi299 & n50515;
  assign n50517 = ~pi211 & n49602;
  assign n50518 = pi214 & ~n61161;
  assign n50519 = ~pi211 & ~n50508;
  assign n50520 = pi214 & ~n50519;
  assign n50521 = ~n50507 & n50520;
  assign n50522 = ~n50507 & n50518;
  assign n50523 = ~n50514 & ~n61162;
  assign n50524 = pi212 & ~n50523;
  assign n50525 = n50513 & ~n50524;
  assign n50526 = ~n49344 & n50490;
  assign n50527 = pi219 & ~n50526;
  assign n50528 = n49344 & ~n50507;
  assign n50529 = n50527 & ~n50528;
  assign n50530 = n58992 & ~n50529;
  assign n50531 = ~n50525 & n50530;
  assign n50532 = n50482 & ~n50531;
  assign n50533 = ~n36621 & n50477;
  assign n50534 = n49760 & ~n50533;
  assign n50535 = ~n49449 & n50534;
  assign n50536 = ~n58992 & n50535;
  assign n50537 = ~pi1152 & ~n50536;
  assign n50538 = pi211 & ~n50490;
  assign n50539 = pi214 & ~n50538;
  assign n50540 = n50520 & ~n50538;
  assign n50541 = ~n50519 & n50539;
  assign n50542 = ~n50514 & ~n61163;
  assign n50543 = pi212 & ~n50542;
  assign n50544 = n50513 & ~n50543;
  assign n50545 = pi219 & ~n50490;
  assign n50546 = n58992 & ~n50545;
  assign n50547 = ~n50544 & n50546;
  assign n50548 = n50537 & ~n50547;
  assign n50549 = ~pi213 & ~n50548;
  assign n50550 = ~pi213 & ~n50532;
  assign n50551 = ~n50548 & n50550;
  assign n50552 = ~n50532 & n50549;
  assign n50553 = ~n49646 & ~n49989;
  assign n50554 = ~pi208 & ~n50553;
  assign n50555 = n61117 & ~n50488;
  assign n50556 = pi208 & ~n50555;
  assign n50557 = ~n50554 & ~n50556;
  assign n50558 = ~pi211 & ~n50557;
  assign n50559 = n49553 & ~n49972;
  assign n50560 = pi207 & ~n46506;
  assign n50561 = ~n50487 & n50560;
  assign n50562 = pi208 & ~n50561;
  assign n50563 = n49544 & ~n50561;
  assign n50564 = ~n49543 & n50562;
  assign n50565 = ~n50559 & ~n61165;
  assign n50566 = pi211 & ~n50565;
  assign n50567 = ~n50558 & ~n50566;
  assign n50568 = pi214 & n50567;
  assign n50569 = n50492 & ~n50568;
  assign n50570 = ~pi214 & n50567;
  assign n50571 = pi211 & ~n50501;
  assign n50572 = ~pi211 & ~n50565;
  assign n50573 = pi214 & ~n50572;
  assign n50574 = ~n50571 & n50573;
  assign n50575 = pi212 & ~n50574;
  assign n50576 = ~n50570 & n50575;
  assign n50577 = ~pi219 & ~n50576;
  assign n50578 = ~pi219 & ~n50569;
  assign n50579 = ~n50576 & n50578;
  assign n50580 = ~n50569 & n50577;
  assign n50581 = ~n49343 & n50502;
  assign n50582 = n50527 & ~n50581;
  assign n50583 = n35344 & ~n50582;
  assign n50584 = ~n61166 & n50583;
  assign n50585 = pi209 & ~n50584;
  assign n50586 = ~n61164 & n50585;
  assign n50587 = ~pi1153 & ~n45444;
  assign n50588 = n49491 & ~n50587;
  assign n50589 = ~n47136 & ~n50588;
  assign n50590 = ~n36320 & n50589;
  assign n50591 = n36320 & ~n47001;
  assign n50592 = ~n49819 & ~n50591;
  assign n50593 = ~n50590 & n50592;
  assign n50594 = pi211 & ~n50593;
  assign n50595 = ~n47134 & ~n47158;
  assign n50596 = n46422 & ~n50595;
  assign n50597 = n49582 & ~n50596;
  assign n50598 = ~pi207 & n50596;
  assign n50599 = ~n46359 & n46995;
  assign n50600 = pi207 & n50599;
  assign n50601 = pi208 & ~n50600;
  assign n50602 = ~n50598 & n50601;
  assign n50603 = ~n50597 & ~n50602;
  assign n50604 = ~pi211 & n50603;
  assign n50605 = ~pi211 & ~n50603;
  assign n50606 = pi211 & n50593;
  assign n50607 = ~n50605 & ~n50606;
  assign n50608 = ~n50594 & ~n50604;
  assign n50609 = ~n49343 & ~n61167;
  assign n50610 = pi219 & ~n50593;
  assign n50611 = ~n49826 & ~n50610;
  assign n50612 = ~n50609 & ~n50611;
  assign n50613 = n58992 & ~n50612;
  assign n50614 = ~pi214 & ~n50593;
  assign n50615 = ~pi212 & ~n50614;
  assign n50616 = pi207 & ~n50589;
  assign n50617 = ~n49458 & ~n50616;
  assign n50618 = ~pi208 & ~n50617;
  assign n50619 = pi207 & ~n50599;
  assign n50620 = ~n49584 & n50619;
  assign n50621 = ~n46496 & ~n50588;
  assign n50622 = ~n47136 & n50621;
  assign n50623 = ~pi207 & ~n50622;
  assign n50624 = ~n50620 & ~n50623;
  assign n50625 = pi208 & ~n50624;
  assign n50626 = ~n50618 & ~n50625;
  assign n50627 = ~pi211 & ~n50626;
  assign n50628 = ~pi207 & n49464;
  assign n50629 = pi1154 & ~n45521;
  assign n50630 = ~n47125 & n50629;
  assign n50631 = ~n47126 & ~n50630;
  assign n50632 = pi207 & ~n50631;
  assign n50633 = ~n50628 & ~n50632;
  assign n50634 = ~pi208 & ~n50633;
  assign n50635 = ~pi207 & ~n50631;
  assign n50636 = pi207 & ~n46384;
  assign n50637 = ~n47014 & n50636;
  assign n50638 = ~n50635 & ~n50637;
  assign n50639 = pi208 & ~n50638;
  assign n50640 = ~n50634 & ~n50639;
  assign n50641 = pi211 & ~n50640;
  assign n50642 = ~n50627 & ~n50641;
  assign n50643 = pi214 & n50642;
  assign n50644 = n50615 & ~n50643;
  assign n50645 = ~pi214 & n50642;
  assign n50646 = pi211 & ~n50603;
  assign n50647 = ~pi211 & ~n50640;
  assign n50648 = pi214 & ~n50647;
  assign n50649 = ~n50646 & n50648;
  assign n50650 = pi212 & ~n50649;
  assign n50651 = ~n50645 & n50650;
  assign n50652 = ~pi219 & ~n50651;
  assign n50653 = ~pi219 & ~n50644;
  assign n50654 = ~n50651 & n50653;
  assign n50655 = ~n50644 & n50652;
  assign n50656 = n50613 & ~n61168;
  assign n50657 = n50482 & ~n50656;
  assign n50658 = ~n47124 & ~n50630;
  assign n50659 = pi207 & ~n50658;
  assign n50660 = ~n50628 & ~n50659;
  assign n50661 = ~pi208 & ~n50660;
  assign n50662 = ~pi207 & ~n50658;
  assign n50663 = pi1153 & n49945;
  assign n50664 = ~n50662 & ~n50663;
  assign n50665 = pi208 & ~n50664;
  assign n50666 = ~n61119 & ~n50665;
  assign n50667 = ~n50661 & n50666;
  assign n50668 = ~n47014 & ~n47231;
  assign n50669 = pi1154 & ~n50668;
  assign n50670 = ~n47133 & ~n50669;
  assign n50671 = pi207 & ~n50670;
  assign n50672 = ~n50493 & ~n50671;
  assign n50673 = ~pi208 & ~n50672;
  assign n50674 = ~pi207 & n50670;
  assign n50675 = ~pi299 & ~pi1153;
  assign n50676 = ~n36720 & ~n50675;
  assign n50677 = ~n49584 & n50676;
  assign n50678 = pi207 & ~n50677;
  assign n50679 = pi208 & ~n50678;
  assign n50680 = ~n50674 & n50679;
  assign n50681 = ~n50673 & ~n50680;
  assign n50682 = n61121 & n50681;
  assign n50683 = ~n50661 & ~n50665;
  assign n50684 = n49706 & n50683;
  assign n50685 = ~pi211 & n50681;
  assign n50686 = pi211 & n50683;
  assign n50687 = ~n50685 & ~n50686;
  assign n50688 = ~n61092 & ~n50687;
  assign n50689 = ~n50684 & ~n50688;
  assign n50690 = ~n50667 & ~n50682;
  assign n50691 = ~pi219 & ~n61169;
  assign n50692 = pi1154 & ~n47152;
  assign n50693 = ~n47134 & ~n50692;
  assign n50694 = n49820 & n50693;
  assign n50695 = n46958 & n49814;
  assign n50696 = ~n50694 & ~n50695;
  assign n50697 = pi219 & n50696;
  assign n50698 = n58992 & ~n50697;
  assign n50699 = n61092 & ~n49445;
  assign n50700 = n50696 & n50699;
  assign n50701 = n50698 & ~n50700;
  assign n50702 = ~n50691 & n50701;
  assign n50703 = n50537 & ~n50702;
  assign n50704 = ~n50657 & ~n50703;
  assign n50705 = ~pi213 & n50704;
  assign n50706 = ~n49344 & n50593;
  assign n50707 = ~n49343 & n50627;
  assign n50708 = ~n50706 & ~n50707;
  assign n50709 = pi219 & ~n50708;
  assign n50710 = pi211 & ~n50626;
  assign n50711 = n49553 & ~n50596;
  assign n50712 = ~n50602 & ~n50711;
  assign n50713 = ~pi1154 & n36719;
  assign n50714 = n60918 & n49581;
  assign n50715 = ~n49611 & ~n50714;
  assign n50716 = ~n50712 & n50715;
  assign n50717 = ~pi211 & n50716;
  assign n50718 = n36621 & ~n50717;
  assign n50719 = ~n50710 & n50718;
  assign n50720 = pi211 & n50716;
  assign n50721 = ~n49646 & n50589;
  assign n50722 = ~pi207 & ~n50721;
  assign n50723 = pi299 & ~pi1156;
  assign n50724 = n50619 & ~n50723;
  assign n50725 = pi208 & ~n50724;
  assign n50726 = ~n50722 & n50725;
  assign n50727 = n49993 & ~n50616;
  assign n50728 = ~pi211 & ~n50727;
  assign n50729 = ~n50726 & n50728;
  assign n50730 = ~n61092 & ~n50729;
  assign n50731 = ~n50720 & n50730;
  assign n50732 = ~pi212 & n50614;
  assign n50733 = ~pi219 & ~n50732;
  assign n50734 = ~n50731 & n50733;
  assign n50735 = ~n50719 & n50734;
  assign n50736 = ~n50709 & ~n50735;
  assign n50737 = n47450 & ~n50736;
  assign n50738 = ~pi1152 & n58992;
  assign n50739 = ~pi299 & ~n60948;
  assign n50740 = ~pi1154 & ~n50739;
  assign n50741 = ~n49611 & n50740;
  assign n50742 = ~n47101 & n50669;
  assign n50743 = ~n50741 & ~n50742;
  assign n50744 = pi207 & n50743;
  assign n50745 = n49553 & ~n50744;
  assign n50746 = ~pi207 & n50743;
  assign n50747 = ~n49611 & n50676;
  assign n50748 = pi207 & ~n50747;
  assign n50749 = pi208 & ~n50748;
  assign n50750 = ~n50746 & n50749;
  assign n50751 = ~n50745 & ~n50750;
  assign n50752 = ~pi211 & n50751;
  assign n50753 = pi211 & n50681;
  assign n50754 = n36621 & ~n50753;
  assign n50755 = n36621 & ~n50752;
  assign n50756 = ~n50753 & n50755;
  assign n50757 = ~n50752 & n50754;
  assign n50758 = pi211 & n50751;
  assign n50759 = ~pi211 & ~n49646;
  assign n50760 = n50696 & n50759;
  assign n50761 = ~n61092 & ~n50760;
  assign n50762 = ~n50758 & n50761;
  assign n50763 = ~n61170 & ~n50762;
  assign n50764 = ~pi219 & ~n50763;
  assign n50765 = n49343 & ~n50696;
  assign n50766 = pi211 & n50696;
  assign n50767 = n49826 & ~n50766;
  assign n50768 = ~n50685 & n50767;
  assign n50769 = ~n50765 & ~n50768;
  assign n50770 = ~n50764 & n50769;
  assign n50771 = n50738 & ~n50770;
  assign n50772 = ~n50737 & ~n50771;
  assign n50773 = pi213 & ~n50772;
  assign n50774 = ~pi209 & ~n50773;
  assign n50775 = ~n50705 & n50774;
  assign n50776 = ~n50586 & ~n50775;
  assign n50777 = ~pi212 & n49840;
  assign n50778 = n49351 & ~n49422;
  assign n50779 = ~pi219 & ~n61171;
  assign n50780 = ~n61095 & n50779;
  assign n50781 = pi213 & ~n47142;
  assign n50782 = n49346 & n50781;
  assign n50783 = ~n50780 & n50782;
  assign n50784 = ~n50776 & ~n50783;
  assign n50785 = pi230 & ~n50784;
  assign n50786 = ~pi230 & pi234;
  assign n50787 = ~n50785 & ~n50786;
  assign n50788 = ~pi230 & ~pi235;
  assign n50789 = ~n46706 & ~n61105;
  assign n50790 = pi207 & ~n50789;
  assign n50791 = ~n49971 & ~n50790;
  assign n50792 = pi208 & ~n50791;
  assign n50793 = ~n49560 & ~n50792;
  assign n50794 = ~pi1157 & ~n50793;
  assign n50795 = ~n49980 & ~n50790;
  assign n50796 = n49953 & ~n50795;
  assign n50797 = ~n49556 & ~n50796;
  assign n50798 = ~n50794 & n50797;
  assign n50799 = pi211 & ~n50798;
  assign n50800 = ~pi1156 & n46520;
  assign n50801 = ~n49610 & ~n50800;
  assign n50802 = pi207 & ~n50801;
  assign n50803 = ~n49990 & ~n50802;
  assign n50804 = pi208 & ~n50803;
  assign n50805 = ~n49656 & ~n50804;
  assign n50806 = ~pi1157 & ~n50805;
  assign n50807 = ~n50000 & ~n50802;
  assign n50808 = n49953 & ~n50807;
  assign n50809 = ~n49658 & ~n50808;
  assign n50810 = ~n50806 & n50809;
  assign n50811 = ~pi211 & ~n50810;
  assign n50812 = n36621 & ~n50811;
  assign n50813 = n36621 & ~n50799;
  assign n50814 = ~n50811 & n50813;
  assign n50815 = ~n50799 & n50812;
  assign n50816 = n36320 & ~n61105;
  assign n50817 = ~n50800 & n50816;
  assign n50818 = ~n49899 & ~n50817;
  assign n50819 = ~n49490 & n50818;
  assign n50820 = ~pi1157 & ~n50819;
  assign n50821 = ~n49913 & ~n50817;
  assign n50822 = ~n49534 & n50821;
  assign n50823 = pi1157 & ~n50822;
  assign n50824 = ~n50820 & ~n50823;
  assign n50825 = n49343 & ~n50824;
  assign n50826 = pi211 & ~n50810;
  assign n50827 = ~n61138 & n49929;
  assign n50828 = ~n49583 & ~n50827;
  assign n50829 = pi1157 & n50828;
  assign n50830 = n49593 & ~n50827;
  assign n50831 = ~pi211 & ~n50820;
  assign n50832 = ~n61173 & n50831;
  assign n50833 = ~n61092 & ~n50832;
  assign n50834 = ~n50826 & n50833;
  assign n50835 = ~n50825 & ~n50834;
  assign n50836 = ~n61172 & n50835;
  assign n50837 = ~pi219 & ~n50836;
  assign n50838 = ~pi211 & n50798;
  assign n50839 = pi211 & ~n50824;
  assign n50840 = ~n61092 & ~n50839;
  assign n50841 = ~n50838 & n50840;
  assign n50842 = n61092 & n50824;
  assign n50843 = pi219 & ~n50842;
  assign n50844 = ~n50841 & n50843;
  assign n50845 = pi209 & ~n50844;
  assign n50846 = ~n50837 & n50845;
  assign n50847 = ~n49508 & n49553;
  assign n50848 = ~pi207 & n49508;
  assign n50849 = pi208 & ~n50744;
  assign n50850 = ~n50848 & n50849;
  assign n50851 = ~n50847 & ~n50850;
  assign n50852 = pi211 & n50851;
  assign n50853 = n36320 & ~n50693;
  assign n50854 = n61104 & ~n49819;
  assign n50855 = ~n36320 & ~n50854;
  assign n50856 = ~n50853 & ~n50855;
  assign n50857 = n50759 & ~n50856;
  assign n50858 = ~n50852 & ~n50857;
  assign n50859 = ~n49646 & ~n50856;
  assign n50860 = ~pi211 & ~n50859;
  assign n50861 = pi211 & ~n50851;
  assign n50862 = n36621 & ~n50861;
  assign n50863 = ~n50860 & n50862;
  assign n50864 = n36621 & ~n50858;
  assign n50865 = n49343 & ~n50856;
  assign n50866 = pi211 & n49646;
  assign n50867 = ~n46291 & ~n50866;
  assign n50868 = ~n50856 & n50867;
  assign n50869 = ~n50669 & ~n50740;
  assign n50870 = pi207 & n50869;
  assign n50871 = n49581 & n49607;
  assign n50872 = pi208 & ~n50871;
  assign n50873 = ~n50870 & n50872;
  assign n50874 = n49582 & ~n61115;
  assign n50875 = pi1157 & n49344;
  assign n50876 = ~n50874 & n50875;
  assign n50877 = ~n50873 & n50876;
  assign n50878 = ~n50868 & ~n50877;
  assign n50879 = ~n36621 & ~n50878;
  assign n50880 = ~n50865 & ~n50879;
  assign n50881 = ~n50873 & ~n50874;
  assign n50882 = pi1157 & ~n50881;
  assign n50883 = ~pi1157 & n50856;
  assign n50884 = ~pi211 & ~n50883;
  assign n50885 = ~pi211 & ~n50882;
  assign n50886 = ~n50883 & n50885;
  assign n50887 = ~n50882 & n50884;
  assign n50888 = pi211 & n50859;
  assign n50889 = ~n61175 & ~n50888;
  assign n50890 = ~n61092 & ~n50889;
  assign n50891 = ~n61174 & ~n50865;
  assign n50892 = ~n50890 & n50891;
  assign n50893 = ~n61174 & n50880;
  assign n50894 = ~pi219 & ~n61176;
  assign n50895 = ~pi211 & n50851;
  assign n50896 = pi211 & ~n50856;
  assign n50897 = ~n61092 & ~n50896;
  assign n50898 = ~n50895 & n50897;
  assign n50899 = n61092 & n50856;
  assign n50900 = pi219 & ~n50899;
  assign n50901 = ~n50898 & n50900;
  assign n50902 = ~pi209 & ~n50901;
  assign n50903 = ~n50894 & n50902;
  assign n50904 = ~n50846 & ~n50903;
  assign n50905 = n58992 & ~n50904;
  assign n50906 = ~n61096 & n49849;
  assign n50907 = n49438 & ~n61131;
  assign n50908 = pi219 & n61092;
  assign n50909 = ~n58992 & ~n47067;
  assign n50910 = ~n47067 & ~n50908;
  assign n50911 = ~n58992 & n50910;
  assign n50912 = ~n50908 & n50909;
  assign n50913 = ~n61177 & n61178;
  assign n50914 = pi213 & ~n50913;
  assign n50915 = ~n50905 & n50914;
  assign n50916 = ~pi299 & ~pi1157;
  assign n50917 = ~n50806 & n50916;
  assign n50918 = n50805 & n50916;
  assign n50919 = ~n49602 & ~n61173;
  assign n50920 = pi1157 & ~n50828;
  assign n50921 = pi299 & ~pi1157;
  assign n50922 = ~n50806 & ~n50921;
  assign n50923 = ~n50920 & n50922;
  assign n50924 = ~n49602 & ~n50923;
  assign n50925 = ~n61179 & n50919;
  assign n50926 = ~pi211 & ~n61180;
  assign n50927 = n50840 & ~n50926;
  assign n50928 = n50843 & ~n50927;
  assign n50929 = pi211 & n61180;
  assign n50930 = ~n46521 & ~n61111;
  assign n50931 = ~n49584 & ~n61111;
  assign n50932 = ~n61105 & ~n61181;
  assign n50933 = pi207 & ~n50932;
  assign n50934 = ~n50023 & ~n50933;
  assign n50935 = pi208 & ~n50934;
  assign n50936 = ~n49588 & ~n50935;
  assign n50937 = ~pi1157 & ~n50936;
  assign n50938 = n49585 & ~n50828;
  assign n50939 = ~n50937 & ~n50938;
  assign n50940 = ~pi211 & ~n50939;
  assign n50941 = n36621 & ~n50940;
  assign n50942 = ~n50929 & n50941;
  assign n50943 = pi211 & n50939;
  assign n50944 = ~n50838 & ~n50943;
  assign n50945 = ~n61092 & ~n50944;
  assign n50946 = ~n50825 & ~n50945;
  assign n50947 = ~n50942 & n50946;
  assign n50948 = ~pi219 & ~n50947;
  assign n50949 = ~n50928 & ~n50948;
  assign n50950 = pi209 & ~n50949;
  assign n50951 = ~n49608 & ~n50628;
  assign n50952 = ~pi208 & ~n50951;
  assign n50953 = ~pi207 & ~n49607;
  assign n50954 = ~n50659 & ~n50953;
  assign n50955 = pi208 & ~n50954;
  assign n50956 = ~n50952 & ~n50955;
  assign n50957 = ~pi211 & n50956;
  assign n50958 = n50897 & ~n50957;
  assign n50959 = n50900 & ~n50958;
  assign n50960 = ~n49572 & ~n50493;
  assign n50961 = ~pi208 & ~n50960;
  assign n50962 = ~pi207 & ~n49571;
  assign n50963 = ~n50671 & ~n50962;
  assign n50964 = pi208 & ~n50963;
  assign n50965 = ~n61119 & ~n50964;
  assign n50966 = ~n50961 & n50965;
  assign n50967 = n61121 & n50851;
  assign n50968 = n60503 & n50956;
  assign n50969 = ~n50865 & ~n50968;
  assign n50970 = ~n50967 & n50969;
  assign n50971 = ~n50961 & ~n50964;
  assign n50972 = pi211 & n50971;
  assign n50973 = ~n50895 & ~n50972;
  assign n50974 = ~n61092 & ~n50973;
  assign n50975 = ~pi211 & ~n50971;
  assign n50976 = pi211 & ~n50956;
  assign n50977 = n36621 & ~n50976;
  assign n50978 = ~n50975 & n50977;
  assign n50979 = ~n50865 & ~n50978;
  assign n50980 = ~n50974 & n50979;
  assign n50981 = ~n50966 & n50970;
  assign n50982 = ~pi219 & ~n61182;
  assign n50983 = ~n50959 & ~n50982;
  assign n50984 = ~pi209 & ~n50983;
  assign n50985 = n58992 & ~n50984;
  assign n50986 = ~n50950 & n50985;
  assign n50987 = ~n61092 & ~n49424;
  assign n50988 = n36621 & ~n50477;
  assign n50989 = ~pi219 & ~n50988;
  assign n50990 = ~pi219 & ~n50987;
  assign n50991 = ~n50988 & n50990;
  assign n50992 = ~n50987 & n50989;
  assign n50993 = ~n60964 & ~n50908;
  assign n50994 = ~n50908 & ~n61183;
  assign n50995 = ~n60964 & n50994;
  assign n50996 = ~n61183 & n50993;
  assign n50997 = ~pi213 & ~n61184;
  assign n50998 = ~n50986 & n50997;
  assign n50999 = ~n50915 & ~n50998;
  assign n51000 = pi230 & ~n50999;
  assign po392 = ~n50788 & ~n51000;
  assign n51002 = ~pi230 & pi238;
  assign n51003 = n46499 & n47123;
  assign n51004 = n50621 & ~n51003;
  assign n51005 = pi207 & ~n51004;
  assign n51006 = ~n50962 & ~n51005;
  assign n51007 = pi208 & ~n51006;
  assign n51008 = ~n50961 & ~n51007;
  assign n51009 = pi211 & ~n51008;
  assign n51010 = ~n46999 & n50748;
  assign n51011 = ~pi1154 & ~n50675;
  assign n51012 = ~n46736 & n51011;
  assign n51013 = pi207 & ~n51012;
  assign n51014 = n50621 & n51013;
  assign n51015 = pi208 & ~n51014;
  assign n51016 = ~n51010 & n51015;
  assign n51017 = ~n50848 & n51016;
  assign n51018 = ~n50847 & ~n51017;
  assign n51019 = ~pi211 & ~n51018;
  assign n51020 = n49351 & ~n51019;
  assign n51021 = ~n51009 & n51020;
  assign n51022 = n49666 & ~n51008;
  assign n51023 = n49565 & ~n51018;
  assign n51024 = ~n47318 & ~n50588;
  assign n51025 = pi207 & ~n51024;
  assign n51026 = ~n50953 & ~n51025;
  assign n51027 = pi208 & ~n51026;
  assign n51028 = ~n50952 & ~n51027;
  assign n51029 = n36620 & ~n51028;
  assign n51030 = pi212 & ~n51029;
  assign n51031 = ~n51023 & n51030;
  assign n51032 = ~n51022 & n51031;
  assign n51033 = ~n51021 & ~n51032;
  assign n51034 = ~pi219 & ~n51033;
  assign n51035 = n36320 & ~n51003;
  assign n51036 = ~n50588 & n51035;
  assign n51037 = ~n50855 & ~n51036;
  assign n51038 = pi211 & n51037;
  assign n51039 = ~pi211 & ~n51028;
  assign n51040 = ~n51038 & ~n51039;
  assign n51041 = n49826 & n51040;
  assign n51042 = ~pi214 & ~n51037;
  assign n51043 = ~pi212 & n51042;
  assign n51044 = pi209 & n58992;
  assign n51045 = ~n51043 & n51044;
  assign n51046 = ~n51041 & n51045;
  assign n51047 = ~n51034 & n51046;
  assign n51048 = ~pi207 & ~n46995;
  assign n51049 = ~n49945 & ~n51048;
  assign n51050 = pi208 & ~n51049;
  assign n51051 = ~n46995 & n49582;
  assign n51052 = ~n51050 & ~n51051;
  assign n51053 = ~pi211 & ~n49584;
  assign n51054 = ~n51052 & n51053;
  assign n51055 = ~n45425 & ~n47231;
  assign n51056 = pi207 & ~n51055;
  assign n51057 = ~n50628 & ~n51056;
  assign n51058 = ~pi208 & ~n51057;
  assign n51059 = pi200 & pi207;
  assign n51060 = ~pi199 & ~n51059;
  assign n51061 = ~pi299 & ~n51060;
  assign n51062 = pi208 & ~n51061;
  assign n51063 = ~pi207 & n36719;
  assign n51064 = ~pi299 & ~n51063;
  assign n51065 = ~pi1153 & ~n51064;
  assign n51066 = n51062 & ~n51065;
  assign n51067 = ~n51058 & ~n51066;
  assign n51068 = pi211 & ~n51067;
  assign n51069 = ~n51054 & ~n51068;
  assign n51070 = n36621 & ~n51069;
  assign n51071 = ~n61092 & ~n51052;
  assign n51072 = pi299 & n49424;
  assign n51073 = n51071 & ~n51072;
  assign n51074 = ~n51070 & ~n51073;
  assign n51075 = ~pi219 & ~n51074;
  assign n51076 = ~n36320 & n46977;
  assign n51077 = ~n49820 & ~n49994;
  assign n51078 = n45518 & ~n51077;
  assign n51079 = ~n51076 & n51078;
  assign n51080 = ~pi211 & n49464;
  assign n51081 = ~n49343 & n51080;
  assign n51082 = ~n51079 & ~n51081;
  assign n51083 = ~n49760 & ~n51082;
  assign n51084 = ~n51075 & ~n51083;
  assign n51085 = n60971 & ~n51084;
  assign n51086 = n50599 & ~n50636;
  assign n51087 = pi208 & ~n51086;
  assign n51088 = n49582 & ~n50600;
  assign n51089 = ~n51087 & ~n51088;
  assign n51090 = ~pi211 & ~n51089;
  assign n51091 = ~n49611 & n51090;
  assign n51092 = pi211 & ~n51089;
  assign n51093 = ~n49584 & n51092;
  assign n51094 = ~n51091 & ~n51093;
  assign n51095 = ~n61092 & ~n51094;
  assign n51096 = n36719 & n49820;
  assign n51097 = ~pi299 & ~n51096;
  assign n51098 = n47143 & ~n51097;
  assign n51099 = n46498 & n49374;
  assign n51100 = pi208 & n46999;
  assign n51101 = ~n51063 & n51100;
  assign n51102 = ~n51099 & ~n51101;
  assign n51103 = ~n51098 & n51102;
  assign n51104 = ~n51054 & n51103;
  assign n51105 = n36621 & ~n51104;
  assign n51106 = n45444 & n49820;
  assign n51107 = pi1153 & n51106;
  assign n51108 = n51102 & ~n51107;
  assign n51109 = ~pi214 & n51102;
  assign n51110 = ~n51107 & n51109;
  assign n51111 = ~pi212 & ~n51110;
  assign n51112 = ~pi214 & n51111;
  assign n51113 = n49343 & ~n51108;
  assign n51114 = ~pi219 & ~n61185;
  assign n51115 = ~n51105 & n51114;
  assign n51116 = ~n51095 & n51115;
  assign n51117 = ~n45447 & ~n51097;
  assign n51118 = ~pi214 & ~n51106;
  assign n51119 = ~pi212 & n51118;
  assign n51120 = n51117 & ~n51119;
  assign n51121 = pi1153 & n51120;
  assign n51122 = pi219 & n51102;
  assign n51123 = ~n51121 & n51122;
  assign n51124 = n47428 & ~n51123;
  assign n51125 = ~n51116 & n51124;
  assign n51126 = pi1152 & ~n51125;
  assign n51127 = ~n51085 & n51126;
  assign n51128 = ~n36320 & n46389;
  assign n51129 = ~n49819 & n51128;
  assign n51130 = n46498 & n49814;
  assign n51131 = ~n46498 & n49374;
  assign n51132 = pi208 & ~n51131;
  assign n51133 = pi200 & n49581;
  assign n51134 = n51132 & ~n51133;
  assign n51135 = ~pi299 & n51134;
  assign n51136 = ~n49889 & ~n51135;
  assign n51137 = ~n51129 & ~n51130;
  assign n51138 = ~n46985 & ~n47088;
  assign n51139 = ~n49553 & ~n51132;
  assign n51140 = ~n51138 & ~n51139;
  assign n51141 = ~n51130 & ~n51140;
  assign n51142 = ~pi299 & ~n51141;
  assign n51143 = ~n47000 & ~n61186;
  assign n51144 = ~pi214 & ~n61187;
  assign n51145 = ~pi212 & ~n51144;
  assign n51146 = pi299 & ~n49424;
  assign n51147 = pi214 & ~n51146;
  assign n51148 = ~n61187 & n51147;
  assign n51149 = n51145 & ~n51148;
  assign n51150 = n49565 & n51141;
  assign n51151 = ~pi299 & ~n49994;
  assign n51152 = ~pi208 & ~n51151;
  assign n51153 = ~n51134 & ~n51152;
  assign n51154 = ~n47014 & ~n51153;
  assign n51155 = n36620 & ~n51154;
  assign n51156 = ~n49458 & n49666;
  assign n51157 = ~n61187 & n51156;
  assign n51158 = pi212 & ~n51157;
  assign n51159 = ~n51155 & n51158;
  assign n51160 = ~n51150 & n51159;
  assign n51161 = ~pi219 & ~n51160;
  assign n51162 = ~n51149 & n51161;
  assign n51163 = ~pi211 & ~n51153;
  assign n51164 = pi211 & ~n61186;
  assign n51165 = ~n51163 & ~n51164;
  assign n51166 = ~n47014 & ~n51165;
  assign n51167 = n49343 & ~n61187;
  assign n51168 = n51166 & ~n51167;
  assign n51169 = pi219 & ~n51168;
  assign n51170 = n47428 & ~n51169;
  assign n51171 = ~n51162 & n51170;
  assign n51172 = ~n49458 & ~n51107;
  assign n51173 = ~pi211 & ~n51172;
  assign n51174 = n36621 & ~n51098;
  assign n51175 = ~n51173 & n51174;
  assign n51176 = ~n61092 & ~n51146;
  assign n51177 = ~n51107 & n51176;
  assign n51178 = ~n51175 & ~n51177;
  assign n51179 = ~pi219 & ~n51178;
  assign n51180 = ~n49760 & ~n51121;
  assign n51181 = n60971 & ~n51180;
  assign n51182 = ~n51179 & n51181;
  assign n51183 = ~pi1152 & ~n51182;
  assign n51184 = ~n51171 & n51183;
  assign n51185 = ~pi209 & ~n51184;
  assign n51186 = ~n51127 & n51185;
  assign n51187 = pi219 & n50515;
  assign n51188 = ~pi1153 & n36681;
  assign n51189 = n49346 & ~n61188;
  assign n51190 = ~n61183 & n51189;
  assign n51191 = ~n51186 & ~n51190;
  assign n51192 = ~n51127 & ~n51184;
  assign n51193 = ~pi209 & ~n51192;
  assign n51194 = n58992 & ~n51043;
  assign n51195 = ~n51041 & n51194;
  assign n51196 = ~n51034 & n51195;
  assign n51197 = pi209 & ~n51196;
  assign n51198 = ~n51193 & ~n51197;
  assign n51199 = ~n51190 & ~n51198;
  assign n51200 = ~n51047 & n51191;
  assign n51201 = pi213 & ~n61189;
  assign n51202 = ~n60503 & n49760;
  assign n51203 = ~n58992 & n51202;
  assign n51204 = ~pi1153 & n36678;
  assign n51205 = ~n36621 & n50515;
  assign n51206 = ~n36621 & ~n50515;
  assign n51207 = ~n36682 & ~n47068;
  assign n51208 = ~n60503 & ~n61190;
  assign n51209 = ~n49706 & ~n51206;
  assign n51210 = n51203 & ~n61191;
  assign n51211 = n51203 & ~n61190;
  assign n51212 = ~pi1151 & ~n61192;
  assign n51213 = ~n50871 & n51015;
  assign n51214 = ~n50874 & ~n51213;
  assign n51215 = pi211 & ~n51214;
  assign n51216 = ~n51039 & ~n51215;
  assign n51217 = pi214 & n51216;
  assign n51218 = ~pi212 & ~n51042;
  assign n51219 = ~n51217 & n51218;
  assign n51220 = ~pi219 & ~n51219;
  assign n51221 = ~pi214 & ~n51216;
  assign n51222 = ~pi211 & ~n51214;
  assign n51223 = ~n51038 & ~n51222;
  assign n51224 = pi214 & ~n51223;
  assign n51225 = ~n51221 & ~n51224;
  assign n51226 = pi212 & ~n51225;
  assign n51227 = n51220 & ~n51226;
  assign n51228 = pi219 & ~n51037;
  assign n51229 = n58992 & ~n51228;
  assign n51230 = ~n51227 & n51229;
  assign n51231 = n51212 & ~n51230;
  assign n51232 = ~n36624 & n49346;
  assign n51233 = pi1151 & ~n51232;
  assign n51234 = ~n61192 & n51233;
  assign n51235 = ~n49343 & n51223;
  assign n51236 = ~n51043 & ~n51235;
  assign n51237 = pi219 & ~n51236;
  assign n51238 = n58992 & ~n51237;
  assign n51239 = pi214 & ~n51214;
  assign n51240 = ~n51221 & ~n51239;
  assign n51241 = pi212 & ~n51240;
  assign n51242 = n51220 & ~n51241;
  assign n51243 = n51238 & ~n51242;
  assign n51244 = n51234 & ~n51243;
  assign n51245 = pi1152 & ~n51244;
  assign n51246 = pi1152 & ~n51231;
  assign n51247 = ~n51244 & n51246;
  assign n51248 = ~n51231 & n51245;
  assign n51249 = pi1153 & n61121;
  assign n51250 = n47068 & ~n61092;
  assign n51251 = n36624 & ~n61194;
  assign n51252 = n49346 & ~n51251;
  assign n51253 = pi1151 & ~n51252;
  assign n51254 = pi214 & n51040;
  assign n51255 = ~n51042 & ~n51254;
  assign n51256 = ~pi212 & ~n51255;
  assign n51257 = ~pi214 & ~n51040;
  assign n51258 = ~pi211 & n51037;
  assign n51259 = ~n51215 & ~n51258;
  assign n51260 = pi214 & ~n51259;
  assign n51261 = pi212 & ~n51260;
  assign n51262 = pi212 & ~n51257;
  assign n51263 = ~n51260 & n51262;
  assign n51264 = ~n51257 & n51261;
  assign n51265 = ~n51256 & ~n61195;
  assign n51266 = ~pi219 & ~n51265;
  assign n51267 = n51238 & ~n51266;
  assign n51268 = n51253 & ~n51267;
  assign n51269 = n36678 & n49760;
  assign n51270 = n60512 & ~n49343;
  assign n51271 = n36679 & ~n61092;
  assign n51272 = ~pi219 & ~n61092;
  assign n51273 = n45884 & n51272;
  assign n51274 = n36624 & ~n61121;
  assign n51275 = n51203 & ~n51274;
  assign n51276 = n61121 & n51203;
  assign n51277 = ~n58992 & n61196;
  assign n51278 = n47437 & n61194;
  assign n51279 = pi1153 & n61197;
  assign n51280 = ~pi1151 & ~n61198;
  assign n51281 = n51040 & n51272;
  assign n51282 = ~n51037 & ~n51272;
  assign n51283 = n58992 & ~n51282;
  assign n51284 = ~n51281 & n51283;
  assign n51285 = n51280 & ~n51284;
  assign n51286 = ~pi1152 & ~n51285;
  assign n51287 = ~n51268 & n51286;
  assign n51288 = pi209 & ~n51287;
  assign n51289 = ~n51268 & ~n51285;
  assign n51290 = ~pi1152 & ~n51289;
  assign n51291 = ~n51231 & ~n51244;
  assign n51292 = pi1152 & ~n51291;
  assign n51293 = ~n51290 & ~n51292;
  assign n51294 = pi209 & ~n51293;
  assign n51295 = pi209 & ~n61193;
  assign n51296 = ~n51287 & n51295;
  assign n51297 = ~n61193 & n51288;
  assign n51298 = ~pi214 & n51166;
  assign n51299 = ~n45447 & ~n51107;
  assign n51300 = ~n61187 & n51299;
  assign n51301 = pi214 & ~n51300;
  assign n51302 = pi212 & ~n51301;
  assign n51303 = ~n51298 & n51302;
  assign n51304 = ~pi212 & ~n51168;
  assign n51305 = ~n51303 & ~n51304;
  assign n51306 = ~pi219 & ~n51305;
  assign n51307 = ~n45445 & ~n51107;
  assign n51308 = ~n61187 & n51307;
  assign n51309 = ~n51167 & ~n51308;
  assign n51310 = pi219 & ~n51309;
  assign n51311 = n58992 & ~n51310;
  assign n51312 = ~n51306 & n51311;
  assign n51313 = n51253 & ~n51312;
  assign n51314 = n51118 & n51121;
  assign n51315 = pi212 & ~n51118;
  assign n51316 = ~n51299 & n51315;
  assign n51317 = ~pi219 & ~n51316;
  assign n51318 = n49351 & n51080;
  assign n51319 = ~n51106 & ~n51318;
  assign n51320 = n51317 & n51319;
  assign n51321 = ~n51314 & n51320;
  assign n51322 = pi219 & ~n51106;
  assign n51323 = n58992 & ~n51322;
  assign n51324 = n51121 & n51323;
  assign n51325 = ~n51321 & n51324;
  assign n51326 = n51280 & ~n51325;
  assign n51327 = ~pi1152 & ~n51326;
  assign n51328 = ~n51313 & n51327;
  assign n51329 = ~n51090 & n51108;
  assign n51330 = pi214 & n51329;
  assign n51331 = ~n51110 & ~n51330;
  assign n51332 = ~pi212 & ~n51331;
  assign n51333 = ~n51329 & ~n51332;
  assign n51334 = pi219 & ~n51333;
  assign n51335 = n58992 & ~n51334;
  assign n51336 = pi1153 & ~n51097;
  assign n51337 = ~n51092 & ~n51336;
  assign n51338 = n51109 & n51337;
  assign n51339 = pi214 & n51089;
  assign n51340 = pi212 & ~n51339;
  assign n51341 = ~n51338 & n51340;
  assign n51342 = pi214 & n51102;
  assign n51343 = n51337 & n51342;
  assign n51344 = n51111 & ~n51343;
  assign n51345 = ~pi219 & ~n51344;
  assign n51346 = ~n51341 & n51345;
  assign n51347 = n51335 & ~n51346;
  assign n51348 = n51234 & ~n51347;
  assign n51349 = pi219 & ~n51079;
  assign n51350 = n58992 & ~n51349;
  assign n51351 = ~pi211 & n51067;
  assign n51352 = n51071 & ~n51351;
  assign n51353 = n61092 & n51079;
  assign n51354 = pi299 & n49706;
  assign n51355 = ~pi219 & ~n51354;
  assign n51356 = ~n51353 & n51355;
  assign n51357 = ~n51352 & n51356;
  assign n51358 = n51350 & ~n51357;
  assign n51359 = n51212 & ~n51358;
  assign n51360 = pi1152 & ~n51359;
  assign n51361 = ~n51348 & n51360;
  assign n51362 = ~n51348 & ~n51359;
  assign n51363 = pi1152 & ~n51362;
  assign n51364 = ~n51313 & ~n51326;
  assign n51365 = ~pi1152 & ~n51364;
  assign n51366 = ~n51363 & ~n51365;
  assign n51367 = ~n51328 & ~n51361;
  assign n51368 = ~pi209 & ~n61200;
  assign n51369 = ~pi213 & ~n51368;
  assign n51370 = ~n61199 & n51369;
  assign n51371 = ~n51201 & ~n51370;
  assign n51372 = pi230 & ~n51371;
  assign n51373 = ~n51002 & ~n51372;
  assign n51374 = n49381 & ~n49516;
  assign n51375 = ~pi214 & n51374;
  assign n51376 = ~pi212 & ~n51375;
  assign n51377 = ~pi219 & n51376;
  assign n51378 = ~n50554 & n50759;
  assign n51379 = pi211 & ~n46506;
  assign n51380 = ~n50559 & n51379;
  assign n51381 = pi214 & ~n51380;
  assign n51382 = ~n51378 & n51381;
  assign n51383 = n51377 & ~n51382;
  assign n51384 = pi212 & ~n51374;
  assign n51385 = n58992 & ~n51384;
  assign n51386 = pi219 & n51376;
  assign n51387 = pi211 & ~n51374;
  assign n51388 = pi214 & ~n51387;
  assign n51389 = ~n49458 & ~n50495;
  assign n51390 = n51388 & ~n51389;
  assign n51391 = n51386 & ~n51390;
  assign n51392 = n51385 & ~n51391;
  assign n51393 = ~n51383 & n51385;
  assign n51394 = ~n51391 & n51393;
  assign n51395 = ~n51383 & n51392;
  assign n51396 = ~pi209 & ~n61201;
  assign n51397 = ~pi214 & n61144;
  assign n51398 = ~pi212 & ~n51397;
  assign n51399 = pi219 & n51398;
  assign n51400 = ~pi211 & ~n49458;
  assign n51401 = ~n61144 & n51400;
  assign n51402 = pi211 & ~n61144;
  assign n51403 = pi214 & ~n51402;
  assign n51404 = ~n51401 & n51403;
  assign n51405 = n51399 & ~n51404;
  assign n51406 = pi212 & ~n61144;
  assign n51407 = n58992 & ~n51406;
  assign n51408 = ~pi219 & n51398;
  assign n51409 = ~n61144 & n50759;
  assign n51410 = pi214 & ~n51409;
  assign n51411 = ~n61144 & n51379;
  assign n51412 = n51410 & ~n51411;
  assign n51413 = n51408 & ~n51412;
  assign n51414 = n51407 & ~n51413;
  assign n51415 = ~n51405 & n51414;
  assign n51416 = pi209 & ~n51415;
  assign n51417 = ~n51396 & ~n51416;
  assign n51418 = n49351 & ~n50779;
  assign n51419 = n47171 & n51418;
  assign n51420 = ~pi213 & ~n51419;
  assign n51421 = ~n51417 & n51420;
  assign n51422 = pi299 & pi1158;
  assign n51423 = ~n49381 & n51422;
  assign n51424 = ~pi208 & n49938;
  assign n51425 = ~n51423 & ~n51424;
  assign n51426 = ~pi211 & ~n51425;
  assign n51427 = pi208 & pi299;
  assign n51428 = pi1157 & ~n51427;
  assign n51429 = ~n50503 & n51428;
  assign n51430 = ~pi1157 & ~n51374;
  assign n51431 = pi211 & ~n51430;
  assign n51432 = ~n51429 & n51431;
  assign n51433 = ~n51426 & ~n51432;
  assign n51434 = pi214 & ~n51433;
  assign n51435 = n51377 & ~n51434;
  assign n51436 = ~n51378 & n51388;
  assign n51437 = n51386 & ~n51436;
  assign n51438 = ~pi209 & n51385;
  assign n51439 = ~n51437 & n51438;
  assign n51440 = ~n51435 & n51439;
  assign n51441 = pi208 & ~n51422;
  assign n51442 = ~n49552 & ~n51441;
  assign n51443 = ~n49950 & n51442;
  assign n51444 = n49963 & ~n51443;
  assign n51445 = ~n49922 & n51428;
  assign n51446 = ~n50024 & ~n51445;
  assign n51447 = pi211 & ~n51446;
  assign n51448 = pi214 & ~n51447;
  assign n51449 = ~n51444 & n51448;
  assign n51450 = n51408 & ~n51449;
  assign n51451 = ~n51402 & n51410;
  assign n51452 = n51399 & ~n51451;
  assign n51453 = pi209 & n51407;
  assign n51454 = ~n51452 & n51453;
  assign n51455 = ~n51450 & n51453;
  assign n51456 = ~n51452 & n51455;
  assign n51457 = ~n51450 & n51454;
  assign n51458 = ~n49848 & ~n49854;
  assign n51459 = pi213 & ~n51458;
  assign n51460 = ~n61202 & n51459;
  assign n51461 = ~n51440 & n51460;
  assign n51462 = ~n51421 & ~n51461;
  assign n51463 = pi230 & ~n51462;
  assign n51464 = ~pi230 & ~pi239;
  assign po396 = ~n51463 & ~n51464;
  assign n51466 = n49346 & ~n51274;
  assign n51467 = pi211 & ~n51153;
  assign n51468 = ~pi211 & ~n61186;
  assign n51469 = pi214 & ~n51468;
  assign n51470 = pi214 & ~n51467;
  assign n51471 = ~n51468 & n51470;
  assign n51472 = ~n51467 & n51469;
  assign n51473 = n36621 & ~n61203;
  assign n51474 = ~pi214 & n61186;
  assign n51475 = ~pi212 & ~n51474;
  assign n51476 = pi214 & n51165;
  assign n51477 = n51475 & ~n51476;
  assign n51478 = ~pi219 & ~n51477;
  assign n51479 = pi212 & ~n61203;
  assign n51480 = ~n51165 & n51479;
  assign n51481 = n51478 & ~n51480;
  assign n51482 = ~n51473 & n51481;
  assign n51483 = pi212 & ~n51165;
  assign n51484 = pi219 & ~n51483;
  assign n51485 = ~n51477 & n51484;
  assign n51486 = n58992 & ~n51485;
  assign n51487 = ~n51482 & n51486;
  assign n51488 = ~n51466 & ~n51487;
  assign n51489 = pi1147 & n51488;
  assign n51490 = n44774 & n51096;
  assign n51491 = n49295 & n61121;
  assign n51492 = ~n51490 & ~n51491;
  assign n51493 = ~pi1147 & n51492;
  assign n51494 = pi1149 & ~n51493;
  assign n51495 = ~n51489 & n51494;
  assign n51496 = pi299 & n36620;
  assign n51497 = ~pi212 & ~n51496;
  assign n51498 = n51102 & n51497;
  assign n51499 = ~n45445 & n51102;
  assign n51500 = ~n51109 & ~n51499;
  assign n51501 = ~pi214 & n45447;
  assign n51502 = pi212 & ~n51501;
  assign n51503 = ~n51500 & n51502;
  assign n51504 = ~n51498 & ~n51503;
  assign n51505 = ~pi219 & ~n51504;
  assign n51506 = n46422 & ~n51059;
  assign n51507 = pi208 & ~n51506;
  assign n51508 = ~pi199 & ~n51507;
  assign n51509 = ~n51102 & ~n51508;
  assign n51510 = ~pi299 & ~n51509;
  assign n51511 = ~pi219 & n51510;
  assign n51512 = ~n51505 & ~n51511;
  assign n51513 = ~pi211 & ~n51512;
  assign n51514 = ~pi214 & n51499;
  assign n51515 = pi212 & ~n51514;
  assign n51516 = ~n45447 & n51342;
  assign n51517 = n51515 & ~n51516;
  assign n51518 = ~pi212 & n51500;
  assign n51519 = ~pi219 & ~n51518;
  assign n51520 = ~n51517 & n51519;
  assign n51521 = n58992 & ~n51102;
  assign n51522 = n58992 & ~n49345;
  assign n51523 = pi219 & ~n45445;
  assign n51524 = n51522 & ~n51523;
  assign n51525 = ~n51521 & ~n51524;
  assign n51526 = ~n51520 & ~n51525;
  assign n51527 = ~n51510 & n51526;
  assign n51528 = ~n51513 & n51527;
  assign n51529 = ~n51232 & ~n51528;
  assign n51530 = pi1147 & ~pi1149;
  assign n51531 = ~n51529 & n51530;
  assign n51532 = ~n51495 & ~n51531;
  assign n51533 = ~pi1148 & ~n51532;
  assign n51534 = pi212 & ~n49565;
  assign n51535 = ~pi219 & ~n51534;
  assign n51536 = ~pi219 & ~n49708;
  assign n51537 = ~n51534 & n51536;
  assign n51538 = ~n49708 & n51535;
  assign n51539 = n49346 & ~n61204;
  assign n51540 = pi1147 & ~n51539;
  assign n51541 = n49392 & n51522;
  assign n51542 = ~n61204 & n51541;
  assign n51543 = ~n51521 & ~n51542;
  assign n51544 = ~n51521 & ~n51539;
  assign n51545 = ~n51542 & n51544;
  assign n51546 = ~n51539 & n51543;
  assign n51547 = pi1147 & n61205;
  assign n51548 = n51540 & n51543;
  assign n51549 = ~n49820 & ~n49945;
  assign n51550 = ~n36320 & n46705;
  assign n51551 = ~n51549 & ~n51550;
  assign n51552 = n51064 & n51551;
  assign n51553 = ~n51496 & ~n51552;
  assign n51554 = ~pi212 & ~n51553;
  assign n51555 = ~pi219 & ~n51554;
  assign n51556 = ~pi299 & ~n51551;
  assign n51557 = pi214 & ~n51556;
  assign n51558 = ~pi214 & n51552;
  assign n51559 = ~pi212 & ~n51558;
  assign n51560 = ~n51557 & n51559;
  assign n51561 = ~pi214 & ~n51556;
  assign n51562 = pi211 & ~n51064;
  assign n51563 = ~pi211 & ~n51556;
  assign n51564 = ~n51552 & ~n51563;
  assign n51565 = ~n51556 & ~n51562;
  assign n51566 = pi214 & ~n61207;
  assign n51567 = pi212 & ~n51566;
  assign n51568 = ~n51561 & n51567;
  assign n51569 = ~n51560 & ~n51568;
  assign n51570 = ~n45447 & ~n51552;
  assign n51571 = ~n51557 & n51570;
  assign n51572 = pi212 & ~n51571;
  assign n51573 = n51569 & n51572;
  assign n51574 = n51555 & ~n51573;
  assign n51575 = pi219 & ~n51552;
  assign n51576 = n58992 & ~n51575;
  assign n51577 = ~n51574 & n51576;
  assign n51578 = n47437 & ~n61119;
  assign n51579 = ~pi1147 & ~n51578;
  assign n51580 = ~n51577 & ~n51578;
  assign n51581 = ~pi1147 & n51580;
  assign n51582 = ~n51577 & n51579;
  assign n51583 = ~n61206 & ~n61208;
  assign n51584 = ~pi1149 & ~n51583;
  assign n51585 = n58992 & n51078;
  assign n51586 = ~n51323 & ~n51585;
  assign n51587 = ~pi214 & ~n51078;
  assign n51588 = ~pi212 & ~n51587;
  assign n51589 = n45518 & n49381;
  assign n51590 = ~pi299 & ~n51589;
  assign n51591 = ~n45521 & n49582;
  assign n51592 = ~n51062 & ~n51591;
  assign n51593 = ~n51062 & n51590;
  assign n51594 = pi214 & n61209;
  assign n51595 = n51588 & ~n51594;
  assign n51596 = ~pi219 & ~n51595;
  assign n51597 = ~pi211 & ~n61209;
  assign n51598 = pi211 & n51078;
  assign n51599 = pi214 & ~n51598;
  assign n51600 = ~n51597 & n51599;
  assign n51601 = pi212 & ~n51600;
  assign n51602 = ~n61209 & n51601;
  assign n51603 = n51596 & ~n51602;
  assign n51604 = ~n51586 & ~n51603;
  assign n51605 = ~n51203 & ~n51604;
  assign n51606 = ~pi1147 & ~n51605;
  assign n51607 = n46999 & ~n49819;
  assign n51608 = n58992 & n51607;
  assign n51609 = ~n51541 & ~n51608;
  assign n51610 = ~n45884 & ~n47437;
  assign n51611 = ~n49343 & ~n51610;
  assign n51612 = n51609 & ~n51611;
  assign n51613 = pi1147 & ~n51612;
  assign n51614 = pi1149 & ~n51613;
  assign n51615 = ~n51606 & n51614;
  assign n51616 = pi1148 & ~n51615;
  assign n51617 = ~pi1147 & n51605;
  assign n51618 = pi1147 & n51612;
  assign n51619 = pi1149 & ~n51618;
  assign n51620 = ~n51617 & n51619;
  assign n51621 = ~pi1149 & ~n61206;
  assign n51622 = ~n61208 & n51621;
  assign n51623 = ~n51620 & ~n51622;
  assign n51624 = pi1148 & ~n51623;
  assign n51625 = ~n51584 & n51616;
  assign n51626 = ~n51533 & ~n61210;
  assign n51627 = pi213 & n51626;
  assign n51628 = ~pi211 & n50047;
  assign n51629 = pi219 & ~n51628;
  assign n51630 = n51522 & ~n51629;
  assign n51631 = pi219 & n61186;
  assign n51632 = n58992 & ~n51631;
  assign n51633 = ~n51630 & ~n51632;
  assign n51634 = pi299 & pi1146;
  assign n51635 = n61186 & ~n51634;
  assign n51636 = pi211 & ~n51635;
  assign n51637 = ~n51163 & ~n51636;
  assign n51638 = ~pi214 & n51637;
  assign n51639 = ~pi211 & pi1146;
  assign n51640 = pi211 & pi1145;
  assign n51641 = ~n51639 & ~n51640;
  assign n51642 = pi299 & ~n51641;
  assign n51643 = pi214 & ~n51642;
  assign n51644 = n61186 & n51643;
  assign n51645 = pi212 & ~n51644;
  assign n51646 = ~n51638 & n51645;
  assign n51647 = pi214 & n51637;
  assign n51648 = n51475 & ~n51647;
  assign n51649 = ~pi219 & ~n51648;
  assign n51650 = ~pi219 & ~n51646;
  assign n51651 = ~n51648 & n51650;
  assign n51652 = ~n51646 & n51649;
  assign n51653 = ~n51633 & ~n61211;
  assign n51654 = pi214 & ~n51641;
  assign n51655 = pi211 & pi1146;
  assign n51656 = ~pi214 & n51655;
  assign n51657 = ~n51654 & ~n51656;
  assign n51658 = pi212 & ~n51657;
  assign n51659 = n49351 & n51655;
  assign n51660 = ~n51658 & ~n51659;
  assign n51661 = ~n49826 & n51660;
  assign n51662 = ~n58992 & n49797;
  assign n51663 = ~n47437 & ~n51662;
  assign n51664 = ~n51661 & ~n51663;
  assign n51665 = pi1147 & ~n61197;
  assign n51666 = ~n51664 & n51665;
  assign n51667 = ~n51653 & n51666;
  assign n51668 = ~pi1147 & ~n51664;
  assign n51669 = pi219 & n51630;
  assign n51670 = pi299 & ~n51660;
  assign n51671 = n35404 & n51670;
  assign n51672 = ~n51669 & ~n51671;
  assign n51673 = n51668 & n51672;
  assign n51674 = ~n51490 & n51673;
  assign n51675 = ~pi1148 & ~n51674;
  assign n51676 = ~n51667 & n51675;
  assign n51677 = ~n49343 & n51597;
  assign n51678 = ~n49344 & n51078;
  assign n51679 = pi219 & ~n51678;
  assign n51680 = ~n51677 & n51679;
  assign n51681 = n58992 & ~n51680;
  assign n51682 = n45518 & n51681;
  assign n51683 = ~n51630 & ~n51682;
  assign n51684 = pi211 & n51634;
  assign n51685 = ~n51078 & ~n51684;
  assign n51686 = n51588 & ~n51685;
  assign n51687 = pi212 & ~n61209;
  assign n51688 = ~n51078 & n51657;
  assign n51689 = n51687 & ~n51688;
  assign n51690 = ~pi219 & ~n51689;
  assign n51691 = ~pi219 & ~n51686;
  assign n51692 = ~n51689 & n51691;
  assign n51693 = ~n51686 & n51690;
  assign n51694 = ~n51683 & ~n61212;
  assign n51695 = n51668 & ~n51694;
  assign n51696 = pi219 & ~n51607;
  assign n51697 = n58992 & ~n51696;
  assign n51698 = ~pi299 & ~n51607;
  assign n51699 = pi299 & n51534;
  assign n51700 = pi212 & ~n51699;
  assign n51701 = pi212 & ~n51698;
  assign n51702 = ~n51699 & n51701;
  assign n51703 = ~n51698 & n51700;
  assign n51704 = ~pi211 & n49460;
  assign n51705 = ~n51607 & ~n51704;
  assign n51706 = pi211 & ~n51607;
  assign n51707 = ~n49460 & ~n51607;
  assign n51708 = ~pi212 & ~n51707;
  assign n51709 = ~n51706 & n51708;
  assign n51710 = ~pi212 & ~n51705;
  assign n51711 = ~pi219 & ~n61214;
  assign n51712 = ~pi219 & ~n61213;
  assign n51713 = ~n61214 & n51712;
  assign n51714 = ~n61213 & n51711;
  assign n51715 = n51697 & ~n61215;
  assign n51716 = n51672 & ~n51715;
  assign n51717 = n51666 & n51672;
  assign n51718 = ~n51715 & n51717;
  assign n51719 = n51666 & n51716;
  assign n51720 = pi1148 & ~n61216;
  assign n51721 = ~n51695 & n51720;
  assign n51722 = pi1149 & ~n51721;
  assign n51723 = ~n51676 & n51722;
  assign n51724 = ~n51521 & ~n51630;
  assign n51725 = ~n45445 & ~n51684;
  assign n51726 = n51102 & n51725;
  assign n51727 = ~n61092 & ~n51726;
  assign n51728 = n51102 & ~n51642;
  assign n51729 = n36621 & ~n51728;
  assign n51730 = n49343 & ~n51102;
  assign n51731 = ~pi219 & ~n51730;
  assign n51732 = ~n51729 & n51731;
  assign n51733 = ~n51727 & n51732;
  assign n51734 = ~n51724 & ~n51733;
  assign n51735 = n51666 & ~n51734;
  assign n51736 = n58992 & n51552;
  assign n51737 = n51673 & ~n51736;
  assign n51738 = pi1148 & ~n51737;
  assign n51739 = pi1148 & ~n51735;
  assign n51740 = ~n51737 & n51739;
  assign n51741 = ~n51735 & n51738;
  assign n51742 = ~pi1146 & n45447;
  assign n51743 = ~n61092 & ~n51742;
  assign n51744 = ~n51729 & ~n51743;
  assign n51745 = ~pi219 & ~n51510;
  assign n51746 = ~n51744 & n51745;
  assign n51747 = n49797 & n49829;
  assign n51748 = n49826 & n51628;
  assign n51749 = ~n49760 & n51509;
  assign n51750 = ~n61218 & ~n51749;
  assign n51751 = ~n51743 & ~n51749;
  assign n51752 = ~n51729 & n51751;
  assign n51753 = pi219 & ~n51509;
  assign n51754 = ~n51510 & ~n51753;
  assign n51755 = ~n51752 & n51754;
  assign n51756 = ~n61218 & ~n51755;
  assign n51757 = ~n51746 & n51750;
  assign n51758 = n58992 & ~n61219;
  assign n51759 = n51666 & ~n51758;
  assign n51760 = ~pi1148 & ~n51673;
  assign n51761 = ~n51759 & n51760;
  assign n51762 = ~pi1149 & ~n51761;
  assign n51763 = ~pi1148 & ~n51759;
  assign n51764 = ~n51739 & ~n51763;
  assign n51765 = ~n51673 & ~n51764;
  assign n51766 = n51736 & n51739;
  assign n51767 = ~pi1149 & ~n51766;
  assign n51768 = ~n51765 & n51767;
  assign n51769 = ~n61217 & n51762;
  assign n51770 = ~n61217 & ~n51761;
  assign n51771 = ~pi1149 & ~n51770;
  assign n51772 = ~n51676 & ~n51721;
  assign n51773 = pi1149 & ~n51772;
  assign n51774 = ~n51771 & ~n51773;
  assign n51775 = ~n51723 & ~n61220;
  assign n51776 = ~pi213 & n61221;
  assign n51777 = pi209 & ~n51776;
  assign n51778 = ~n51627 & n51777;
  assign n51779 = ~pi199 & pi1146;
  assign n51780 = pi199 & pi1145;
  assign n51781 = ~pi200 & ~n51780;
  assign n51782 = ~n51779 & n51781;
  assign n51783 = pi200 & ~n49817;
  assign n51784 = n49374 & ~n51783;
  assign n51785 = ~n51782 & n51784;
  assign n51786 = ~n49820 & ~n51785;
  assign n51787 = pi200 & ~n51779;
  assign n51788 = ~pi299 & ~n51787;
  assign n51789 = n46359 & ~n51780;
  assign n51790 = n51788 & ~n51789;
  assign n51791 = ~n36320 & ~n51790;
  assign n51792 = ~n51786 & ~n51791;
  assign n51793 = ~n49344 & n51792;
  assign n51794 = pi219 & ~n51793;
  assign n51795 = n49381 & n51790;
  assign n51796 = ~pi207 & n51790;
  assign n51797 = ~n51634 & ~n51785;
  assign n51798 = ~n51796 & n51797;
  assign n51799 = pi208 & ~n51798;
  assign n51800 = ~n51795 & ~n51799;
  assign n51801 = ~pi299 & n51800;
  assign n51802 = ~pi211 & ~n51801;
  assign n51803 = ~n49343 & n51802;
  assign n51804 = n51794 & ~n51803;
  assign n51805 = n58992 & ~n51804;
  assign n51806 = pi211 & ~n51801;
  assign n51807 = n51781 & n51796;
  assign n51808 = n51799 & ~n51807;
  assign n51809 = ~n51781 & n51788;
  assign n51810 = n49381 & n51809;
  assign n51811 = ~n51808 & ~n51810;
  assign n51812 = ~pi299 & n51811;
  assign n51813 = pi214 & ~n51812;
  assign n51814 = ~n51806 & ~n51813;
  assign n51815 = pi212 & ~n51814;
  assign n51816 = n36620 & ~n51801;
  assign n51817 = ~pi219 & ~n51792;
  assign n51818 = ~n51816 & n51817;
  assign n51819 = ~n51815 & n51818;
  assign n51820 = n51805 & ~n51819;
  assign n51821 = ~n49666 & ~n51801;
  assign n51822 = ~n51792 & ~n51821;
  assign n51823 = ~pi214 & ~n51792;
  assign n51824 = ~n51802 & n51823;
  assign n51825 = pi214 & ~n51792;
  assign n51826 = ~n51806 & n51825;
  assign n51827 = pi212 & ~n51826;
  assign n51828 = ~n51824 & n51827;
  assign n51829 = pi212 & ~n51822;
  assign n51830 = ~n51792 & ~n51802;
  assign n51831 = ~pi212 & ~n51823;
  assign n51832 = ~n51830 & n51831;
  assign n51833 = ~pi219 & ~n51832;
  assign n51834 = ~n61222 & n51833;
  assign n51835 = n51820 & ~n51834;
  assign n51836 = ~n51232 & ~n51835;
  assign n51837 = pi1147 & ~n51836;
  assign n51838 = ~n36320 & ~n51809;
  assign n51839 = ~pi299 & ~n51811;
  assign n51840 = ~n51786 & ~n51838;
  assign n51841 = ~pi57 & ~pi1147;
  assign n51842 = ~pi1147 & n58992;
  assign n51843 = n4441 & n51841;
  assign n51844 = n61223 & n61224;
  assign n51845 = ~pi1149 & ~n51844;
  assign n51846 = ~n51837 & n51845;
  assign n51847 = n51805 & ~n51834;
  assign n51848 = ~n51466 & ~n51847;
  assign n51849 = pi1147 & ~n51848;
  assign n51850 = ~pi1147 & n61196;
  assign n51851 = ~n51844 & ~n51850;
  assign n51852 = n44774 & n61196;
  assign n51853 = n51811 & n51852;
  assign n51854 = ~n51851 & ~n51853;
  assign n51855 = pi1149 & ~n51854;
  assign n51856 = ~n51849 & n51855;
  assign n51857 = ~pi1148 & ~n51856;
  assign n51858 = ~n51846 & n51857;
  assign n51859 = ~n49343 & n51812;
  assign n51860 = n36621 & n51830;
  assign n51861 = ~n51859 & ~n51860;
  assign n51862 = ~pi219 & ~n51861;
  assign n51863 = ~n49760 & ~n61223;
  assign n51864 = n58992 & ~n51863;
  assign n51865 = pi214 & n51830;
  assign n51866 = ~n51812 & ~n51865;
  assign n51867 = pi212 & ~n51866;
  assign n51868 = ~pi214 & n61223;
  assign n51869 = ~pi212 & ~n51868;
  assign n51870 = ~n51813 & n51869;
  assign n51871 = ~n51867 & ~n51870;
  assign n51872 = ~pi219 & ~n51871;
  assign n51873 = pi219 & ~n61223;
  assign n51874 = n58992 & ~n51873;
  assign n51875 = ~n51872 & n51874;
  assign n51876 = ~n51862 & n51864;
  assign n51877 = ~pi1147 & ~n51203;
  assign n51878 = ~n61225 & n51877;
  assign n51879 = ~n49392 & n51817;
  assign n51880 = n51805 & ~n51879;
  assign n51881 = pi1147 & ~n51611;
  assign n51882 = ~n51880 & n51881;
  assign n51883 = pi1149 & ~n51882;
  assign n51884 = ~n51878 & n51883;
  assign n51885 = ~n51819 & n61225;
  assign n51886 = n51579 & ~n51885;
  assign n51887 = n51540 & ~n51820;
  assign n51888 = ~pi1149 & ~n51887;
  assign n51889 = ~n51886 & n51888;
  assign n51890 = ~n51884 & ~n51889;
  assign n51891 = pi1148 & ~n51890;
  assign n51892 = pi213 & ~n51891;
  assign n51893 = ~n51858 & n51892;
  assign n51894 = ~n50044 & n51806;
  assign n51895 = n51643 & n51800;
  assign n51896 = ~n51816 & ~n51895;
  assign n51897 = ~n51894 & ~n51896;
  assign n51898 = ~pi214 & n51725;
  assign n51899 = n51800 & n51898;
  assign n51900 = pi212 & ~n51899;
  assign n51901 = ~n51897 & n51900;
  assign n51902 = ~n51684 & ~n61223;
  assign n51903 = ~pi214 & ~n61223;
  assign n51904 = ~pi212 & ~n51903;
  assign n51905 = ~n51902 & n51904;
  assign n51906 = ~pi219 & ~n51905;
  assign n51907 = ~n51832 & n51906;
  assign n51908 = ~n51901 & ~n51905;
  assign n51909 = n51833 & n51908;
  assign n51910 = ~n51901 & n51907;
  assign n51911 = ~n50044 & n51802;
  assign n51912 = ~n49343 & n51911;
  assign n51913 = n51794 & ~n51912;
  assign n51914 = n58992 & ~n51913;
  assign n51915 = ~n61226 & n51914;
  assign n51916 = n51666 & ~n51915;
  assign n51917 = n51643 & ~n61223;
  assign n51918 = ~pi214 & n51902;
  assign n51919 = pi212 & ~n51918;
  assign n51920 = ~n51917 & n51919;
  assign n51921 = n51906 & ~n51920;
  assign n51922 = n49343 & n61223;
  assign n51923 = pi219 & ~n51922;
  assign n51924 = ~n49343 & n61223;
  assign n51925 = ~n49344 & ~n51924;
  assign n51926 = ~pi211 & ~n50047;
  assign n51927 = ~n61223 & n51926;
  assign n51928 = ~n51925 & ~n51927;
  assign n51929 = n51923 & ~n51928;
  assign n51930 = n58992 & ~n51929;
  assign n51931 = ~n51921 & n51930;
  assign n51932 = n51668 & ~n51931;
  assign n51933 = ~n51916 & ~n51932;
  assign n51934 = ~pi213 & ~n51933;
  assign n51935 = ~pi209 & ~n51934;
  assign n51936 = ~n51893 & n51935;
  assign n51937 = pi213 & ~n51626;
  assign n51938 = ~pi213 & ~n61220;
  assign n51939 = ~pi213 & ~n61221;
  assign n51940 = ~n51723 & n51938;
  assign n51941 = pi209 & ~n61227;
  assign n51942 = ~n51937 & n51941;
  assign n51943 = ~n51837 & ~n51844;
  assign n51944 = ~pi1149 & ~n51943;
  assign n51945 = ~n51849 & ~n51854;
  assign n51946 = pi1149 & ~n51945;
  assign n51947 = ~pi1148 & ~n51946;
  assign n51948 = ~n51944 & n51947;
  assign n51949 = pi1148 & ~n51884;
  assign n51950 = ~n51889 & n51949;
  assign n51951 = pi213 & ~n51950;
  assign n51952 = ~n51948 & n51951;
  assign n51953 = ~pi213 & n51933;
  assign n51954 = ~pi209 & ~n51953;
  assign n51955 = ~n51952 & n51954;
  assign n51956 = ~n51942 & ~n51955;
  assign n51957 = ~n51778 & ~n51936;
  assign n51958 = pi230 & n61228;
  assign n51959 = ~pi230 & pi240;
  assign n51960 = pi230 & ~n61228;
  assign n51961 = ~pi230 & ~pi240;
  assign n51962 = ~n51960 & ~n51961;
  assign n51963 = ~n51958 & ~n51959;
  assign n51964 = n51111 & ~n51339;
  assign n51965 = ~pi219 & ~n51964;
  assign n51966 = pi212 & ~n51089;
  assign n51967 = n51965 & ~n51966;
  assign n51968 = pi1152 & ~n51967;
  assign n51969 = n51335 & n51968;
  assign n51970 = pi1151 & ~n51611;
  assign n51971 = ~pi1152 & n51311;
  assign n51972 = ~pi299 & ~n51154;
  assign n51973 = ~n51167 & ~n51972;
  assign n51974 = ~pi219 & ~n51973;
  assign n51975 = n51971 & ~n51974;
  assign n51976 = n51970 & ~n51975;
  assign n51977 = ~n51969 & n51976;
  assign n51978 = ~pi1151 & ~n51539;
  assign n51979 = pi219 & ~n51107;
  assign n51980 = n58992 & ~n51979;
  assign n51981 = ~n51524 & ~n51980;
  assign n51982 = ~n51350 & n51981;
  assign n51983 = n36621 & n51052;
  assign n51984 = ~n51119 & ~n51299;
  assign n51985 = ~n36621 & ~n51079;
  assign n51986 = ~n51984 & n51985;
  assign n51987 = ~n51983 & ~n51986;
  assign n51988 = ~pi219 & ~n51987;
  assign n51989 = ~n51982 & ~n51988;
  assign n51990 = pi1152 & ~n51989;
  assign n51991 = ~pi212 & ~n51097;
  assign n51992 = ~n51118 & n51991;
  assign n51993 = ~n45445 & n51992;
  assign n51994 = ~pi219 & ~n51993;
  assign n51995 = ~pi211 & n51118;
  assign n51996 = pi212 & ~n51097;
  assign n51997 = ~n51995 & n51996;
  assign n51998 = pi214 & ~n51117;
  assign n51999 = n51997 & ~n51998;
  assign n52000 = n51994 & ~n51999;
  assign n52001 = ~n51107 & n51317;
  assign n52002 = ~pi299 & n52001;
  assign n52003 = ~n52000 & ~n52002;
  assign n52004 = n51980 & n52003;
  assign n52005 = ~pi1152 & ~n52004;
  assign n52006 = ~n51981 & ~n52001;
  assign n52007 = n52005 & ~n52006;
  assign n52008 = ~n51990 & ~n52007;
  assign n52009 = n51978 & ~n52008;
  assign n52010 = pi1150 & ~n52009;
  assign n52011 = ~n51977 & n52010;
  assign n52012 = ~n49666 & ~n51089;
  assign n52013 = pi212 & n51108;
  assign n52014 = ~n52012 & n52013;
  assign n52015 = ~n51332 & ~n52014;
  assign n52016 = ~pi219 & ~n52015;
  assign n52017 = pi1152 & ~n52016;
  assign n52018 = n51335 & n52017;
  assign n52019 = pi1151 & ~n51466;
  assign n52020 = ~pi214 & ~n51308;
  assign n52021 = n51302 & ~n52020;
  assign n52022 = ~pi212 & ~n51309;
  assign n52023 = ~n52021 & ~n52022;
  assign n52024 = ~pi219 & ~n52023;
  assign n52025 = n51971 & ~n52024;
  assign n52026 = n52019 & ~n52025;
  assign n52027 = ~n52018 & n52026;
  assign n52028 = ~pi1151 & ~n51232;
  assign n52029 = ~pi1152 & ~n52006;
  assign n52030 = pi1152 & ~n51079;
  assign n52031 = n51317 & n52030;
  assign n52032 = ~n51982 & ~n52031;
  assign n52033 = ~n52029 & n52032;
  assign n52034 = ~n51079 & n51317;
  assign n52035 = pi1152 & ~n51982;
  assign n52036 = ~n52034 & n52035;
  assign n52037 = ~pi1152 & n52006;
  assign n52038 = n52028 & ~n52037;
  assign n52039 = ~n52036 & n52038;
  assign n52040 = n52028 & ~n52033;
  assign n52041 = ~pi1150 & ~n61230;
  assign n52042 = ~n52027 & n52041;
  assign n52043 = pi1149 & ~n52042;
  assign n52044 = pi1149 & ~n52011;
  assign n52045 = ~n52042 & n52044;
  assign n52046 = ~n52011 & n52043;
  assign n52047 = pi1151 & ~n51203;
  assign n52048 = ~pi214 & n51153;
  assign n52049 = pi212 & ~n52048;
  assign n52050 = ~n51476 & n52049;
  assign n52051 = ~n51145 & ~n52050;
  assign n52052 = ~n51972 & ~n52051;
  assign n52053 = ~pi219 & ~n52052;
  assign n52054 = ~n51631 & ~n52053;
  assign n52055 = ~pi1152 & ~n52054;
  assign n52056 = ~n51521 & ~n51980;
  assign n52057 = ~pi214 & n51089;
  assign n52058 = pi212 & ~n52057;
  assign n52059 = ~n51330 & n52058;
  assign n52060 = pi1152 & n51965;
  assign n52061 = ~n52059 & n52060;
  assign n52062 = ~n52056 & ~n52061;
  assign n52063 = n51965 & ~n52059;
  assign n52064 = pi1152 & ~n52063;
  assign n52065 = ~pi1152 & ~n51631;
  assign n52066 = ~n52053 & n52065;
  assign n52067 = ~n52064 & ~n52066;
  assign n52068 = ~n52056 & ~n52067;
  assign n52069 = ~n52055 & n52062;
  assign n52070 = n52047 & ~n61232;
  assign n52071 = ~pi1151 & ~n51578;
  assign n52072 = ~n51079 & ~n52003;
  assign n52073 = n51350 & ~n52072;
  assign n52074 = pi1152 & ~n52073;
  assign n52075 = ~n52005 & ~n52074;
  assign n52076 = n52071 & ~n52075;
  assign n52077 = pi1150 & ~n52076;
  assign n52078 = ~n52070 & n52077;
  assign n52079 = pi1152 & n51079;
  assign n52080 = ~pi1152 & n51107;
  assign n52081 = ~n52079 & ~n52080;
  assign n52082 = n60971 & ~n52081;
  assign n52083 = n51090 & n51272;
  assign n52084 = ~n51089 & n61196;
  assign n52085 = pi1152 & n51108;
  assign n52086 = ~n61233 & n52085;
  assign n52087 = n47414 & n61121;
  assign n52088 = ~pi1152 & ~n52087;
  assign n52089 = ~n61187 & n52088;
  assign n52090 = ~n52086 & ~n52089;
  assign n52091 = n58992 & ~n52090;
  assign n52092 = ~n58992 & ~n61196;
  assign n52093 = pi1151 & ~n52092;
  assign n52094 = ~n52091 & n52093;
  assign n52095 = n51108 & ~n61233;
  assign n52096 = pi1152 & ~n52095;
  assign n52097 = n58992 & ~n52096;
  assign n52098 = n52093 & ~n52097;
  assign n52099 = n60971 & n51107;
  assign n52100 = ~n61187 & ~n52087;
  assign n52101 = n52093 & ~n52100;
  assign n52102 = ~n52099 & ~n52101;
  assign n52103 = ~pi1152 & ~n52102;
  assign n52104 = pi1152 & n60971;
  assign n52105 = n51079 & n52104;
  assign n52106 = ~n52103 & ~n52105;
  assign n52107 = ~n52098 & n52106;
  assign n52108 = ~n52082 & ~n52094;
  assign n52109 = ~pi1150 & ~n61234;
  assign n52110 = ~pi1149 & ~n52109;
  assign n52111 = ~n52078 & n52110;
  assign n52112 = ~pi213 & ~n52111;
  assign n52113 = ~n52078 & ~n52109;
  assign n52114 = ~pi1149 & ~n52113;
  assign n52115 = ~n52011 & ~n52042;
  assign n52116 = pi1149 & ~n52115;
  assign n52117 = ~n52114 & ~n52116;
  assign n52118 = ~n61231 & ~n52111;
  assign n52119 = ~pi213 & ~n61235;
  assign n52120 = ~n61231 & n52112;
  assign n52121 = pi213 & n61200;
  assign n52122 = pi209 & ~n52121;
  assign n52123 = ~n61236 & n52122;
  assign n52124 = ~n61161 & ~n51556;
  assign n52125 = pi214 & n52124;
  assign n52126 = n51559 & ~n52125;
  assign n52127 = ~pi214 & n52124;
  assign n52128 = n51567 & ~n52127;
  assign n52129 = ~n52126 & ~n52128;
  assign n52130 = ~pi219 & ~n52129;
  assign n52131 = n51576 & ~n52130;
  assign n52132 = n51212 & ~n52131;
  assign n52133 = pi211 & ~n61209;
  assign n52134 = ~pi211 & ~n49602;
  assign n52135 = ~n61209 & n52134;
  assign n52136 = ~n52133 & ~n52135;
  assign n52137 = ~pi214 & n52136;
  assign n52138 = n51687 & ~n52137;
  assign n52139 = pi214 & n52136;
  assign n52140 = n51588 & ~n52139;
  assign n52141 = ~pi219 & ~n52140;
  assign n52142 = ~pi219 & ~n52138;
  assign n52143 = ~n52140 & n52142;
  assign n52144 = ~n52138 & n52141;
  assign n52145 = n51681 & ~n61237;
  assign n52146 = n51234 & ~n52145;
  assign n52147 = pi1152 & ~n52146;
  assign n52148 = ~n52132 & n52147;
  assign n52149 = ~n51272 & n51552;
  assign n52150 = ~n49602 & ~n51556;
  assign n52151 = ~pi211 & ~n52150;
  assign n52152 = n51272 & ~n61207;
  assign n52153 = ~n52151 & n52152;
  assign n52154 = ~n52149 & ~n52153;
  assign n52155 = n58992 & ~n52154;
  assign n52156 = n51280 & ~n52155;
  assign n52157 = ~n49666 & ~n61209;
  assign n52158 = ~n51078 & ~n52157;
  assign n52159 = ~n51078 & ~n52133;
  assign n52160 = pi214 & n52159;
  assign n52161 = n51587 & ~n51597;
  assign n52162 = pi212 & ~n52161;
  assign n52163 = ~n52160 & n52162;
  assign n52164 = pi212 & ~n52158;
  assign n52165 = ~n52136 & n61238;
  assign n52166 = ~n51598 & ~n52135;
  assign n52167 = n51588 & ~n52166;
  assign n52168 = ~pi219 & ~n52167;
  assign n52169 = ~n52165 & n52168;
  assign n52170 = n51681 & ~n52169;
  assign n52171 = n51253 & ~n52170;
  assign n52172 = ~pi1152 & ~n52171;
  assign n52173 = ~pi1152 & ~n52156;
  assign n52174 = ~n52171 & n52173;
  assign n52175 = ~n52156 & n52172;
  assign n52176 = pi1150 & ~n61239;
  assign n52177 = ~n52148 & n52176;
  assign n52178 = pi219 & ~n51120;
  assign n52179 = n58992 & ~n52178;
  assign n52180 = n51994 & ~n51997;
  assign n52181 = n52179 & ~n52180;
  assign n52182 = ~n51321 & n52179;
  assign n52183 = n51234 & ~n52182;
  assign n52184 = ~n52181 & n52183;
  assign n52185 = pi299 & n51202;
  assign n52186 = n36624 & n49392;
  assign n52187 = ~n61191 & n61240;
  assign n52188 = ~n61190 & n61240;
  assign n52189 = n51212 & ~n61241;
  assign n52190 = pi1152 & ~n52189;
  assign n52191 = ~n52184 & n52190;
  assign n52192 = pi1153 & n52087;
  assign n52193 = n51080 & n51272;
  assign n52194 = n47414 & n61194;
  assign n52195 = n51280 & ~n61242;
  assign n52196 = ~pi1152 & ~n52195;
  assign n52197 = n51253 & ~n52182;
  assign n52198 = n52196 & ~n52197;
  assign n52199 = ~pi1150 & ~n52198;
  assign n52200 = ~n52191 & n52199;
  assign n52201 = ~n52177 & ~n52200;
  assign n52202 = ~pi1149 & ~n52201;
  assign n52203 = ~n61203 & ~n51474;
  assign n52204 = ~pi219 & ~n52203;
  assign n52205 = ~n51168 & ~n51699;
  assign n52206 = ~pi219 & ~n51699;
  assign n52207 = ~n51168 & n52206;
  assign n52208 = ~n52203 & n52207;
  assign n52209 = n52204 & n52205;
  assign n52210 = n51486 & ~n61243;
  assign n52211 = n51234 & ~n52210;
  assign n52212 = ~n49392 & ~n51509;
  assign n52213 = ~n46499 & n61191;
  assign n52214 = ~n52212 & ~n52213;
  assign n52215 = ~pi219 & ~n52214;
  assign n52216 = n4441 & ~n51753;
  assign n52217 = ~pi57 & n52216;
  assign n52218 = n58992 & ~n51753;
  assign n52219 = ~n52215 & n61244;
  assign n52220 = n51212 & ~n52219;
  assign n52221 = pi1152 & ~n52220;
  assign n52222 = ~n52211 & n52221;
  assign n52223 = ~n51475 & ~n51479;
  assign n52224 = ~n49602 & n51163;
  assign n52225 = ~n51153 & n52134;
  assign n52226 = ~n51164 & ~n61245;
  assign n52227 = ~n51473 & n52226;
  assign n52228 = ~n52223 & ~n52227;
  assign n52229 = ~pi219 & ~n52228;
  assign n52230 = n51486 & ~n52229;
  assign n52231 = n51253 & ~n52230;
  assign n52232 = ~n51509 & ~n52087;
  assign n52233 = n58992 & ~n52232;
  assign n52234 = ~n61161 & n52233;
  assign n52235 = n51280 & ~n52234;
  assign n52236 = ~pi1152 & ~n52235;
  assign n52237 = ~n52231 & n52236;
  assign n52238 = ~n52222 & ~n52237;
  assign n52239 = ~pi1150 & ~n52238;
  assign n52240 = ~pi219 & ~n51607;
  assign n52241 = ~n51699 & n52240;
  assign n52242 = ~pi1153 & n52241;
  assign n52243 = pi212 & n51496;
  assign n52244 = pi299 & n60503;
  assign n52245 = ~pi219 & ~n61246;
  assign n52246 = n51524 & ~n52245;
  assign n52247 = ~n51715 & ~n52246;
  assign n52248 = ~n52242 & ~n52247;
  assign n52249 = n51253 & ~n52248;
  assign n52250 = ~pi1151 & ~n51521;
  assign n52251 = ~pi1152 & ~n52250;
  assign n52252 = ~n52196 & ~n52251;
  assign n52253 = ~n52249 & ~n52252;
  assign n52254 = n4441 & ~n51122;
  assign n52255 = ~pi57 & n52254;
  assign n52256 = n58992 & ~n51122;
  assign n52257 = ~pi299 & n51102;
  assign n52258 = ~n61092 & ~n61161;
  assign n52259 = ~n52257 & n52258;
  assign n52260 = n36621 & ~n51499;
  assign n52261 = n51731 & ~n52260;
  assign n52262 = ~n52259 & n52261;
  assign n52263 = n61247 & ~n52262;
  assign n52264 = n51212 & ~n52263;
  assign n52265 = ~pi211 & n52241;
  assign n52266 = ~n51609 & ~n52265;
  assign n52267 = n51234 & ~n52266;
  assign n52268 = ~n52248 & n52267;
  assign n52269 = pi1152 & ~n52268;
  assign n52270 = pi1152 & ~n52264;
  assign n52271 = ~n52268 & n52270;
  assign n52272 = ~n52264 & n52269;
  assign n52273 = ~n52253 & ~n61248;
  assign n52274 = pi1150 & ~n52273;
  assign n52275 = pi1149 & ~n52274;
  assign n52276 = ~n52239 & n52275;
  assign n52277 = ~pi1150 & ~n52222;
  assign n52278 = ~n52237 & n52277;
  assign n52279 = pi1150 & ~n52253;
  assign n52280 = ~n61248 & n52279;
  assign n52281 = pi1149 & ~n52280;
  assign n52282 = ~n52278 & n52281;
  assign n52283 = ~pi1149 & ~n52200;
  assign n52284 = ~n52177 & n52283;
  assign n52285 = ~n52282 & ~n52284;
  assign n52286 = ~n52202 & ~n52276;
  assign n52287 = pi213 & ~n61249;
  assign n52288 = ~n51577 & n52071;
  assign n52289 = ~n51604 & n52047;
  assign n52290 = pi1150 & ~n52289;
  assign n52291 = ~n52288 & n52290;
  assign n52292 = n50199 & ~n51492;
  assign n52293 = ~pi1149 & ~n52292;
  assign n52294 = ~n52291 & n52293;
  assign n52295 = ~n51487 & n52019;
  assign n52296 = ~n51528 & n52028;
  assign n52297 = ~pi1150 & ~n52296;
  assign n52298 = ~n52295 & n52297;
  assign n52299 = ~n51542 & n51978;
  assign n52300 = ~pi1151 & n61205;
  assign n52301 = ~n51521 & n52299;
  assign n52302 = n51609 & n51970;
  assign n52303 = pi1150 & ~n52302;
  assign n52304 = ~n61250 & n52303;
  assign n52305 = pi1149 & ~n52304;
  assign n52306 = ~n52298 & n52305;
  assign n52307 = ~n52294 & ~n52306;
  assign n52308 = ~pi213 & n52307;
  assign n52309 = ~pi209 & ~n52308;
  assign n52310 = ~pi209 & ~n52287;
  assign n52311 = ~n52308 & n52310;
  assign n52312 = ~n52287 & n52309;
  assign n52313 = pi213 & n61249;
  assign n52314 = ~pi213 & ~n52307;
  assign n52315 = ~pi209 & ~n52314;
  assign n52316 = ~n52313 & n52315;
  assign n52317 = ~pi213 & n61235;
  assign n52318 = pi213 & ~n61200;
  assign n52319 = pi209 & ~n52318;
  assign n52320 = ~n52317 & n52319;
  assign n52321 = ~n52316 & ~n52320;
  assign n52322 = ~n52123 & ~n61251;
  assign n52323 = pi230 & ~n61252;
  assign n52324 = ~pi230 & pi241;
  assign n52325 = pi230 & n61252;
  assign n52326 = ~pi230 & ~pi241;
  assign n52327 = ~n52325 & ~n52326;
  assign n52328 = ~n52323 & ~n52324;
  assign n52329 = ~pi230 & ~pi242;
  assign n52330 = pi214 & ~n49799;
  assign n52331 = ~pi214 & ~n51641;
  assign n52332 = ~n52330 & ~n52331;
  assign n52333 = pi212 & ~n52332;
  assign n52334 = ~pi212 & n51654;
  assign n52335 = ~pi219 & ~n52334;
  assign n52336 = ~n52333 & n52335;
  assign n52337 = pi219 & ~n49349;
  assign n52338 = n49346 & ~n52337;
  assign n52339 = ~n52336 & n52338;
  assign n52340 = pi199 & pi1144;
  assign n52341 = ~pi200 & ~n52340;
  assign n52342 = ~n51779 & n52341;
  assign n52343 = ~pi299 & ~n51783;
  assign n52344 = ~n52342 & n52343;
  assign n52345 = ~pi207 & ~n52344;
  assign n52346 = ~pi299 & ~n49821;
  assign n52347 = ~n49817 & n52341;
  assign n52348 = n52346 & ~n52347;
  assign n52349 = pi207 & ~n52348;
  assign n52350 = pi208 & ~n52349;
  assign n52351 = pi208 & ~n52345;
  assign n52352 = ~n52349 & n52351;
  assign n52353 = ~n52345 & n52350;
  assign n52354 = n49381 & n52344;
  assign n52355 = ~n50047 & ~n52354;
  assign n52356 = ~n61254 & n52355;
  assign n52357 = ~pi211 & ~n52356;
  assign n52358 = ~n49715 & ~n52354;
  assign n52359 = ~n61254 & n52358;
  assign n52360 = pi211 & ~n52359;
  assign n52361 = pi214 & ~n52360;
  assign n52362 = pi214 & ~n52357;
  assign n52363 = ~n52360 & n52362;
  assign n52364 = ~n52357 & n52361;
  assign n52365 = ~n51634 & ~n52354;
  assign n52366 = ~n61254 & n52365;
  assign n52367 = ~pi211 & ~n52366;
  assign n52368 = pi211 & ~n52356;
  assign n52369 = ~n52367 & ~n52368;
  assign n52370 = ~pi214 & n52369;
  assign n52371 = pi212 & ~n52370;
  assign n52372 = pi212 & ~n61255;
  assign n52373 = ~n52370 & n52372;
  assign n52374 = ~n61255 & n52371;
  assign n52375 = n49820 & n52344;
  assign n52376 = ~pi299 & ~n52369;
  assign n52377 = ~n61254 & ~n52375;
  assign n52378 = ~pi214 & ~n61257;
  assign n52379 = ~pi212 & ~n52378;
  assign n52380 = pi214 & n52369;
  assign n52381 = n52379 & ~n52380;
  assign n52382 = ~pi219 & ~n52381;
  assign n52383 = ~n61256 & n52382;
  assign n52384 = ~n49344 & n61257;
  assign n52385 = pi219 & ~n52384;
  assign n52386 = n49344 & ~n52359;
  assign n52387 = n52385 & ~n52386;
  assign n52388 = n58992 & ~n52387;
  assign n52389 = ~n52383 & n52388;
  assign n52390 = ~n52339 & ~n52389;
  assign n52391 = pi213 & n52390;
  assign n52392 = pi211 & ~n52375;
  assign n52393 = n49344 & ~n49768;
  assign n52394 = ~n52354 & n52393;
  assign n52395 = ~n52392 & ~n52394;
  assign n52396 = pi219 & ~n52395;
  assign n52397 = n49343 & ~n52375;
  assign n52398 = pi299 & ~n49388;
  assign n52399 = n49760 & ~n52354;
  assign n52400 = n36621 & ~n49403;
  assign n52401 = ~n61092 & ~n49396;
  assign n52402 = ~n52400 & ~n52401;
  assign n52403 = ~pi219 & ~n52354;
  assign n52404 = ~n52402 & n52403;
  assign n52405 = ~n52398 & n52399;
  assign n52406 = ~n52397 & ~n61258;
  assign n52407 = ~n52396 & n52406;
  assign n52408 = ~n61254 & ~n52407;
  assign n52409 = n58992 & ~n52408;
  assign n52410 = ~pi213 & ~n49363;
  assign n52411 = ~n52409 & n52410;
  assign n52412 = ~n52391 & ~n52411;
  assign n52413 = pi209 & ~n52412;
  assign n52414 = ~pi213 & ~n49420;
  assign n52415 = ~n49343 & n49349;
  assign n52416 = pi219 & n49343;
  assign n52417 = ~n52337 & ~n52416;
  assign n52418 = pi219 & ~n52415;
  assign n52419 = ~n52336 & n61259;
  assign n52420 = pi299 & ~n52419;
  assign n52421 = n58992 & ~n52420;
  assign n52422 = pi299 & n61259;
  assign n52423 = ~n52336 & n52422;
  assign n52424 = ~n49384 & ~n52423;
  assign n52425 = n58992 & ~n52424;
  assign n52426 = ~n49410 & n52421;
  assign n52427 = ~n52339 & ~n61260;
  assign n52428 = pi213 & ~n52427;
  assign n52429 = ~pi209 & ~n52428;
  assign n52430 = ~pi209 & ~n52414;
  assign n52431 = ~n52428 & n52430;
  assign n52432 = ~n52414 & n52429;
  assign n52433 = ~n52413 & ~n61261;
  assign n52434 = pi230 & ~n52433;
  assign po399 = ~n52329 & ~n52434;
  assign n52436 = ~pi230 & ~pi244;
  assign n52437 = pi213 & ~n51933;
  assign n52438 = ~n49717 & n51806;
  assign n52439 = ~n51911 & ~n52438;
  assign n52440 = ~n51812 & ~n52439;
  assign n52441 = pi214 & ~n52440;
  assign n52442 = n51904 & ~n52441;
  assign n52443 = ~pi214 & n52439;
  assign n52444 = n49350 & n49460;
  assign n52445 = pi212 & ~n52444;
  assign n52446 = ~n52443 & n52445;
  assign n52447 = ~n51812 & n52446;
  assign n52448 = ~pi219 & ~n52447;
  assign n52449 = ~pi219 & ~n52442;
  assign n52450 = ~n52447 & n52449;
  assign n52451 = ~n52442 & n52448;
  assign n52452 = ~pi211 & ~n49679;
  assign n52453 = ~n61223 & n52452;
  assign n52454 = ~n51925 & ~n52453;
  assign n52455 = n51923 & ~n52454;
  assign n52456 = n61224 & ~n52455;
  assign n52457 = ~n61262 & n52456;
  assign n52458 = ~n51801 & n52446;
  assign n52459 = pi214 & n52439;
  assign n52460 = n51831 & ~n52459;
  assign n52461 = ~pi219 & ~n52460;
  assign n52462 = ~n52458 & n52461;
  assign n52463 = pi299 & n49807;
  assign n52464 = pi1147 & ~n52463;
  assign n52465 = n51805 & n52464;
  assign n52466 = ~n52462 & n52465;
  assign n52467 = ~pi213 & ~n49809;
  assign n52468 = ~n52466 & n52467;
  assign n52469 = ~n52457 & n52468;
  assign n52470 = ~n52437 & ~n52469;
  assign n52471 = ~n49809 & ~n52466;
  assign n52472 = ~n52457 & n52471;
  assign n52473 = ~pi213 & ~n52472;
  assign n52474 = pi213 & n51933;
  assign n52475 = pi209 & ~n52474;
  assign n52476 = ~n52473 & n52475;
  assign n52477 = pi209 & ~n52470;
  assign n52478 = n51668 & ~n51671;
  assign n52479 = ~n51666 & ~n52478;
  assign n52480 = n51668 & ~n51670;
  assign n52481 = n36621 & ~n51642;
  assign n52482 = ~n36621 & n51725;
  assign n52483 = n49760 & ~n52482;
  assign n52484 = n49760 & ~n52481;
  assign n52485 = ~n52482 & n52484;
  assign n52486 = ~n52481 & n52483;
  assign n52487 = ~n52480 & n61264;
  assign n52488 = ~n49825 & ~n61218;
  assign n52489 = ~n52487 & n52488;
  assign n52490 = n58992 & ~n52489;
  assign n52491 = ~n52479 & ~n52490;
  assign n52492 = pi213 & ~n52491;
  assign n52493 = ~pi213 & ~n49835;
  assign n52494 = ~pi209 & ~n52493;
  assign n52495 = ~n52492 & n52494;
  assign n52496 = ~n61263 & ~n52495;
  assign n52497 = pi230 & ~n52496;
  assign po401 = ~n52436 & ~n52497;
  assign n52499 = ~n49343 & n52367;
  assign n52500 = n49344 & ~n52366;
  assign n52501 = n52385 & ~n61265;
  assign n52502 = n58992 & ~n52501;
  assign n52503 = ~pi299 & n52356;
  assign n52504 = ~pi211 & ~n52503;
  assign n52505 = pi211 & ~n52366;
  assign n52506 = ~n52504 & ~n52505;
  assign n52507 = pi214 & ~n52506;
  assign n52508 = ~pi214 & ~n52503;
  assign n52509 = ~n52507 & ~n52508;
  assign n52510 = pi212 & ~n52509;
  assign n52511 = n52379 & ~n52503;
  assign n52512 = ~pi219 & ~n52511;
  assign n52513 = ~n52510 & n52512;
  assign n52514 = n52502 & ~n52513;
  assign n52515 = pi1146 & n51232;
  assign n52516 = pi1147 & ~n51203;
  assign n52517 = ~n52515 & n52516;
  assign n52518 = ~n52514 & n52517;
  assign n52519 = ~pi1147 & ~n52515;
  assign n52520 = ~n61197 & n52519;
  assign n52521 = pi214 & ~n51684;
  assign n52522 = ~n61257 & n52521;
  assign n52523 = pi212 & ~n52522;
  assign n52524 = ~n61257 & ~n52504;
  assign n52525 = ~pi214 & n52524;
  assign n52526 = n52523 & ~n52525;
  assign n52527 = n52379 & ~n52524;
  assign n52528 = ~pi219 & ~n52527;
  assign n52529 = ~n52526 & n52528;
  assign n52530 = n52502 & ~n52529;
  assign n52531 = n52520 & ~n52530;
  assign n52532 = pi1148 & ~n52531;
  assign n52533 = pi1148 & ~n52518;
  assign n52534 = ~n52531 & n52533;
  assign n52535 = ~n52518 & n52532;
  assign n52536 = ~n51540 & ~n52517;
  assign n52537 = ~n45447 & ~n61257;
  assign n52538 = ~pi214 & ~n52537;
  assign n52539 = ~n52507 & ~n52538;
  assign n52540 = pi212 & ~n52539;
  assign n52541 = n52379 & ~n52537;
  assign n52542 = ~pi219 & ~n52541;
  assign n52543 = ~n52540 & n52542;
  assign n52544 = n52502 & ~n52543;
  assign n52545 = ~n52536 & ~n52544;
  assign n52546 = ~n52378 & n52523;
  assign n52547 = ~pi212 & n61257;
  assign n52548 = ~pi219 & ~n52547;
  assign n52549 = ~n52546 & n52548;
  assign n52550 = n52502 & ~n52549;
  assign n52551 = n52519 & ~n52550;
  assign n52552 = ~pi1148 & ~n52551;
  assign n52553 = ~pi1148 & ~n52545;
  assign n52554 = ~n52551 & n52553;
  assign n52555 = ~n52545 & n52552;
  assign n52556 = ~n52518 & ~n52531;
  assign n52557 = pi1148 & ~n52556;
  assign n52558 = ~n52545 & ~n52551;
  assign n52559 = ~pi1148 & ~n52558;
  assign n52560 = ~n52557 & ~n52559;
  assign n52561 = ~n61266 & ~n61267;
  assign n52562 = pi213 & ~n61268;
  assign n52563 = ~pi213 & n52390;
  assign n52564 = ~pi209 & ~n52563;
  assign n52565 = ~n52562 & n52564;
  assign n52566 = pi199 & pi1146;
  assign n52567 = ~pi200 & ~n52566;
  assign n52568 = n51788 & ~n52567;
  assign n52569 = pi207 & n52568;
  assign n52570 = pi1146 & ~n46422;
  assign n52571 = ~n52569 & ~n52570;
  assign n52572 = pi208 & ~n52571;
  assign n52573 = n46359 & ~n52566;
  assign n52574 = n51788 & ~n52573;
  assign n52575 = pi208 & n52574;
  assign n52576 = ~pi207 & ~n52575;
  assign n52577 = n51128 & ~n52573;
  assign n52578 = ~n52576 & n52577;
  assign n52579 = ~n52572 & ~n52578;
  assign n52580 = ~pi208 & n51634;
  assign n52581 = ~n52572 & ~n52580;
  assign n52582 = ~n52578 & n52581;
  assign n52583 = ~n52578 & ~n52580;
  assign n52584 = ~n52572 & n52583;
  assign n52585 = n52579 & ~n52580;
  assign n52586 = ~pi299 & ~n61269;
  assign n52587 = ~pi299 & ~n52579;
  assign n52588 = ~pi214 & ~n61270;
  assign n52589 = ~pi212 & ~n52588;
  assign n52590 = ~n36320 & ~n51129;
  assign n52591 = n52568 & ~n52590;
  assign n52592 = pi211 & ~n52591;
  assign n52593 = ~pi299 & ~n52568;
  assign n52594 = ~n61269 & ~n52593;
  assign n52595 = ~pi299 & ~n52594;
  assign n52596 = ~pi211 & n52595;
  assign n52597 = ~n52592 & ~n52596;
  assign n52598 = ~n61270 & ~n52597;
  assign n52599 = n52589 & ~n52598;
  assign n52600 = ~pi219 & ~n52599;
  assign n52601 = n52521 & ~n61270;
  assign n52602 = ~pi214 & n52598;
  assign n52603 = pi212 & ~n52602;
  assign n52604 = ~n52601 & n52603;
  assign n52605 = n52600 & ~n52604;
  assign n52606 = ~n49344 & n61270;
  assign n52607 = pi219 & ~n52606;
  assign n52608 = n49344 & ~n61269;
  assign n52609 = n52607 & ~n52608;
  assign n52610 = n58992 & ~n52609;
  assign n52611 = ~n52605 & n52610;
  assign n52612 = n52520 & ~n52611;
  assign n52613 = pi200 & n36320;
  assign n52614 = ~pi199 & ~n52613;
  assign n52615 = ~pi1146 & ~n52614;
  assign n52616 = n46999 & ~n52573;
  assign n52617 = ~n36320 & ~n52616;
  assign n52618 = pi207 & n52574;
  assign n52619 = ~n49820 & ~n52618;
  assign n52620 = ~n52617 & ~n52619;
  assign n52621 = n46999 & ~n52567;
  assign n52622 = ~pi207 & n52621;
  assign n52623 = ~n51634 & ~n52622;
  assign n52624 = ~n52618 & n52623;
  assign n52625 = pi208 & ~n52624;
  assign n52626 = ~pi299 & n52625;
  assign n52627 = n49381 & n52616;
  assign n52628 = ~n52575 & ~n52627;
  assign n52629 = ~n52626 & n52628;
  assign n52630 = n51607 & ~n52615;
  assign n52631 = ~pi214 & ~n61271;
  assign n52632 = ~pi212 & ~n52631;
  assign n52633 = ~pi299 & ~n61271;
  assign n52634 = n52632 & ~n52633;
  assign n52635 = ~pi219 & ~n52634;
  assign n52636 = pi212 & ~n52633;
  assign n52637 = ~n51634 & ~n61271;
  assign n52638 = n36620 & n52637;
  assign n52639 = n52636 & ~n52638;
  assign n52640 = n52635 & ~n52639;
  assign n52641 = ~n49344 & n61271;
  assign n52642 = pi219 & ~n52641;
  assign n52643 = n49344 & ~n52637;
  assign n52644 = n52642 & ~n52643;
  assign n52645 = n58992 & ~n52644;
  assign n52646 = ~n52640 & n52645;
  assign n52647 = n52517 & ~n52646;
  assign n52648 = pi1148 & ~n52647;
  assign n52649 = ~n52612 & n52648;
  assign n52650 = ~n36320 & ~n52621;
  assign n52651 = ~n52619 & ~n52650;
  assign n52652 = ~n45447 & ~n52651;
  assign n52653 = pi214 & ~n52652;
  assign n52654 = ~pi214 & n52651;
  assign n52655 = ~pi212 & ~n52654;
  assign n52656 = ~n52653 & n52655;
  assign n52657 = ~pi214 & ~n52652;
  assign n52658 = n49381 & n52621;
  assign n52659 = ~n52625 & ~n52658;
  assign n52660 = ~n52580 & ~n52658;
  assign n52661 = ~n52580 & n52659;
  assign n52662 = ~n52625 & n52660;
  assign n52663 = ~pi299 & n61272;
  assign n52664 = ~pi299 & n52659;
  assign n52665 = pi214 & ~n61273;
  assign n52666 = ~pi211 & ~n52633;
  assign n52667 = ~n61271 & ~n52666;
  assign n52668 = n52665 & ~n52667;
  assign n52669 = pi212 & ~n52668;
  assign n52670 = ~n52657 & n52669;
  assign n52671 = ~n52656 & ~n52670;
  assign n52672 = ~pi219 & ~n52671;
  assign n52673 = ~pi1146 & ~n49666;
  assign n52674 = n51699 & ~n52673;
  assign n52675 = n52672 & ~n52674;
  assign n52676 = ~n49343 & n52651;
  assign n52677 = ~n49344 & ~n52676;
  assign n52678 = ~n61272 & ~n52677;
  assign n52679 = ~pi212 & n52654;
  assign n52680 = pi219 & ~n52679;
  assign n52681 = ~n52678 & n52680;
  assign n52682 = n58992 & ~n52681;
  assign n52683 = ~n52675 & n52682;
  assign n52684 = ~n52536 & ~n52683;
  assign n52685 = pi219 & ~n52591;
  assign n52686 = ~n49826 & ~n52685;
  assign n52687 = ~n49343 & ~n52592;
  assign n52688 = n52594 & n52687;
  assign n52689 = ~n52686 & ~n52688;
  assign n52690 = ~n61246 & ~n61270;
  assign n52691 = ~n52571 & ~n52690;
  assign n52692 = ~pi219 & ~n52691;
  assign n52693 = n58992 & ~n52692;
  assign n52694 = n58992 & ~n52689;
  assign n52695 = ~n52692 & n52694;
  assign n52696 = ~n52689 & n52693;
  assign n52697 = n52519 & ~n61274;
  assign n52698 = ~pi1148 & ~n52697;
  assign n52699 = ~n52684 & n52698;
  assign n52700 = ~n52649 & ~n52699;
  assign n52701 = pi213 & n52700;
  assign n52702 = ~n51642 & ~n61270;
  assign n52703 = n52589 & ~n52702;
  assign n52704 = pi299 & ~n52332;
  assign n52705 = ~n61270 & ~n52704;
  assign n52706 = pi212 & ~n52705;
  assign n52707 = ~pi219 & ~n52706;
  assign n52708 = ~n52703 & n52707;
  assign n52709 = ~pi299 & n61269;
  assign n52710 = ~pi299 & n52579;
  assign n52711 = n49344 & ~n61275;
  assign n52712 = ~n49717 & n52711;
  assign n52713 = n52607 & ~n52712;
  assign n52714 = n61224 & ~n52713;
  assign n52715 = ~n52708 & n52714;
  assign n52716 = ~n51642 & ~n61271;
  assign n52717 = pi214 & n52716;
  assign n52718 = n52632 & ~n52717;
  assign n52719 = ~n61271 & ~n52704;
  assign n52720 = pi212 & ~n52719;
  assign n52721 = ~pi219 & ~n52720;
  assign n52722 = ~n52718 & n52721;
  assign n52723 = ~pi57 & pi1147;
  assign n52724 = pi1147 & n58992;
  assign n52725 = n4441 & n52723;
  assign n52726 = ~n49715 & ~n61271;
  assign n52727 = n49344 & ~n52726;
  assign n52728 = n52642 & ~n52727;
  assign n52729 = n61276 & ~n52728;
  assign n52730 = ~n52722 & n52729;
  assign n52731 = pi1148 & ~n52339;
  assign n52732 = ~n52730 & n52731;
  assign n52733 = ~n52715 & n52732;
  assign n52734 = ~pi214 & n52591;
  assign n52735 = pi214 & ~n52595;
  assign n52736 = ~n52702 & n52735;
  assign n52737 = ~n52734 & ~n52736;
  assign n52738 = ~pi212 & ~n52737;
  assign n52739 = ~n52593 & n52706;
  assign n52740 = ~pi219 & ~n52739;
  assign n52741 = ~n52738 & n52740;
  assign n52742 = ~n49717 & ~n52595;
  assign n52743 = ~pi211 & ~n52742;
  assign n52744 = n52687 & ~n52743;
  assign n52745 = ~n52686 & ~n52744;
  assign n52746 = n61224 & ~n52745;
  assign n52747 = ~n52741 & n52746;
  assign n52748 = n52665 & ~n52716;
  assign n52749 = ~n52654 & ~n52748;
  assign n52750 = ~pi212 & ~n52749;
  assign n52751 = ~n61273 & n52720;
  assign n52752 = ~pi219 & ~n52751;
  assign n52753 = ~n52750 & n52752;
  assign n52754 = ~n61273 & ~n52726;
  assign n52755 = ~pi211 & ~n52754;
  assign n52756 = ~n52677 & ~n52755;
  assign n52757 = n52680 & ~n52756;
  assign n52758 = n61276 & ~n52757;
  assign n52759 = n61276 & ~n52753;
  assign n52760 = ~n52757 & n52759;
  assign n52761 = ~n52753 & n52758;
  assign n52762 = ~pi1148 & ~n52339;
  assign n52763 = ~n61277 & n52762;
  assign n52764 = ~n52747 & n52763;
  assign n52765 = ~n52733 & ~n52764;
  assign n52766 = ~pi213 & ~n52765;
  assign n52767 = pi209 & ~n52766;
  assign n52768 = ~n52701 & n52767;
  assign n52769 = pi213 & n61268;
  assign n52770 = ~pi213 & ~n52390;
  assign n52771 = ~pi209 & ~n52770;
  assign n52772 = ~n52769 & n52771;
  assign n52773 = pi213 & ~n52700;
  assign n52774 = ~pi213 & ~n52733;
  assign n52775 = ~n52764 & n52774;
  assign n52776 = pi209 & ~n52775;
  assign n52777 = ~n52773 & n52776;
  assign n52778 = ~n52772 & ~n52777;
  assign n52779 = ~n52565 & ~n52768;
  assign n52780 = pi230 & n61278;
  assign n52781 = ~pi230 & pi245;
  assign n52782 = pi230 & ~n61278;
  assign n52783 = ~pi230 & ~pi245;
  assign n52784 = ~n52782 & ~n52783;
  assign n52785 = ~n52780 & ~n52781;
  assign n52786 = ~pi209 & n52700;
  assign n52787 = pi219 & ~n51634;
  assign n52788 = n51522 & ~n52787;
  assign n52789 = ~n51632 & ~n52788;
  assign n52790 = ~n51647 & n52049;
  assign n52791 = ~pi212 & ~n61186;
  assign n52792 = ~pi219 & ~n52791;
  assign n52793 = ~n51992 & n52792;
  assign n52794 = ~n52790 & n52793;
  assign n52795 = ~n52789 & ~n52794;
  assign n52796 = n52517 & ~n52795;
  assign n52797 = n51469 & ~n51636;
  assign n52798 = ~pi214 & n51165;
  assign n52799 = pi212 & ~n52798;
  assign n52800 = ~n52797 & n52799;
  assign n52801 = n51478 & ~n52800;
  assign n52802 = ~n52789 & ~n52801;
  assign n52803 = n52520 & ~n52802;
  assign n52804 = ~n52796 & ~n52803;
  assign n52805 = pi1150 & ~n52804;
  assign n52806 = ~n51511 & ~n51520;
  assign n52807 = n52520 & ~n52806;
  assign n52808 = ~n51508 & n51521;
  assign n52809 = ~n52788 & ~n52808;
  assign n52810 = n61092 & n51742;
  assign n52811 = ~n51510 & ~n51742;
  assign n52812 = n61092 & ~n52811;
  assign n52813 = ~n52212 & ~n52812;
  assign n52814 = ~n52212 & ~n52810;
  assign n52815 = ~pi219 & ~n61280;
  assign n52816 = ~n52809 & ~n52815;
  assign n52817 = ~n52807 & n52816;
  assign n52818 = ~n52517 & ~n52520;
  assign n52819 = ~pi1150 & ~n52818;
  assign n52820 = ~n52817 & n52819;
  assign n52821 = pi1148 & ~n52820;
  assign n52822 = ~n52816 & ~n52818;
  assign n52823 = ~pi1150 & ~n52807;
  assign n52824 = ~n52822 & n52823;
  assign n52825 = pi1150 & ~n52803;
  assign n52826 = ~n52796 & n52825;
  assign n52827 = ~n52824 & ~n52826;
  assign n52828 = pi1148 & ~n52827;
  assign n52829 = ~n52805 & n52821;
  assign n52830 = ~pi219 & ~n51655;
  assign n52831 = ~n52245 & ~n52830;
  assign n52832 = n52788 & n52831;
  assign n52833 = n52519 & ~n52832;
  assign n52834 = ~n52536 & ~n52788;
  assign n52835 = ~n52833 & ~n52834;
  assign n52836 = pi1150 & n51490;
  assign n52837 = ~n52835 & ~n52836;
  assign n52838 = pi1150 & n51106;
  assign n52839 = pi299 & n49708;
  assign n52840 = ~pi219 & ~n52839;
  assign n52841 = ~n52674 & n52840;
  assign n52842 = ~n52838 & n52841;
  assign n52843 = ~n52536 & n52842;
  assign n52844 = ~pi1148 & ~n52843;
  assign n52845 = ~n52837 & n52844;
  assign n52846 = ~n61281 & ~n52845;
  assign n52847 = ~pi1149 & ~n52846;
  assign n52848 = ~pi214 & n52159;
  assign n52849 = n51601 & ~n52848;
  assign n52850 = ~pi219 & ~n52849;
  assign n52851 = ~n51587 & ~n52159;
  assign n52852 = ~pi212 & n52851;
  assign n52853 = n52850 & ~n52852;
  assign n52854 = ~pi299 & n51062;
  assign n52855 = ~n51589 & ~n51634;
  assign n52856 = ~n52854 & n52855;
  assign n52857 = n52853 & n52856;
  assign n52858 = ~n51682 & ~n52788;
  assign n52859 = n52850 & ~n52851;
  assign n52860 = ~n52858 & ~n52859;
  assign n52861 = ~n52857 & n52860;
  assign n52862 = n51588 & ~n51600;
  assign n52863 = ~pi219 & ~n61238;
  assign n52864 = ~pi219 & ~n52862;
  assign n52865 = ~n61238 & n52864;
  assign n52866 = ~n52862 & n52863;
  assign n52867 = n51681 & ~n61282;
  assign n52868 = pi1150 & n52867;
  assign n52869 = n52861 & n52868;
  assign n52870 = n51522 & ~n51556;
  assign n52871 = ~n51576 & ~n52870;
  assign n52872 = ~n51553 & ~n51991;
  assign n52873 = ~pi219 & ~n52872;
  assign n52874 = ~n52871 & ~n52873;
  assign n52875 = ~pi1146 & ~n51552;
  assign n52876 = ~pi1150 & ~n52875;
  assign n52877 = n52874 & n52876;
  assign n52878 = n52519 & ~n52877;
  assign n52879 = ~n52869 & n52878;
  assign n52880 = n49460 & n51655;
  assign n52881 = ~n51552 & ~n52880;
  assign n52882 = n51574 & n52881;
  assign n52883 = ~pi1146 & n51575;
  assign n52884 = ~pi1150 & ~n52883;
  assign n52885 = ~n52871 & n52884;
  assign n52886 = ~n52882 & n52885;
  assign n52887 = pi1150 & n52861;
  assign n52888 = ~n52536 & ~n52887;
  assign n52889 = ~n52886 & n52888;
  assign n52890 = ~n52879 & ~n52889;
  assign n52891 = ~n52871 & ~n52883;
  assign n52892 = ~n52882 & n52891;
  assign n52893 = ~n52536 & ~n52892;
  assign n52894 = n52874 & ~n52875;
  assign n52895 = n52519 & ~n52894;
  assign n52896 = ~pi1150 & ~n52895;
  assign n52897 = ~n52893 & n52896;
  assign n52898 = n52861 & n52867;
  assign n52899 = n52519 & ~n52898;
  assign n52900 = ~n52536 & ~n52861;
  assign n52901 = pi1150 & ~n52900;
  assign n52902 = ~n52899 & n52901;
  assign n52903 = ~pi1148 & ~n52902;
  assign n52904 = ~n52897 & n52903;
  assign n52905 = ~pi1148 & ~n52890;
  assign n52906 = ~n51521 & ~n52788;
  assign n52907 = ~n51499 & n51517;
  assign n52908 = ~n51504 & ~n52907;
  assign n52909 = ~n52520 & ~n52908;
  assign n52910 = n51102 & n52521;
  assign n52911 = n51515 & ~n52910;
  assign n52912 = n51519 & ~n52911;
  assign n52913 = ~n52909 & n52912;
  assign n52914 = ~n52906 & ~n52913;
  assign n52915 = ~n52818 & ~n52914;
  assign n52916 = ~pi1150 & ~n52915;
  assign n52917 = ~n51715 & ~n52832;
  assign n52918 = ~n61197 & ~n51715;
  assign n52919 = n52833 & n52918;
  assign n52920 = n52520 & n52917;
  assign n52921 = pi1146 & n51541;
  assign n52922 = ~n51607 & ~n61240;
  assign n52923 = pi214 & n51706;
  assign n52924 = n51701 & ~n52923;
  assign n52925 = ~pi219 & ~n51708;
  assign n52926 = ~n52924 & n52925;
  assign n52927 = n51697 & ~n52926;
  assign n52928 = n58992 & ~n52922;
  assign n52929 = ~n52921 & ~n61285;
  assign n52930 = n52517 & ~n52921;
  assign n52931 = ~n61285 & n52930;
  assign n52932 = n52517 & n52929;
  assign n52933 = pi1150 & ~n61286;
  assign n52934 = ~n61284 & n52933;
  assign n52935 = pi1148 & ~n52934;
  assign n52936 = ~n52916 & n52935;
  assign n52937 = pi1149 & ~n52936;
  assign n52938 = ~n61283 & n52937;
  assign n52939 = ~n61283 & ~n52936;
  assign n52940 = pi1149 & ~n52939;
  assign n52941 = ~pi1149 & ~n52845;
  assign n52942 = ~n61281 & n52941;
  assign n52943 = ~n52940 & ~n52942;
  assign n52944 = ~n52847 & ~n52938;
  assign n52945 = pi209 & ~n61287;
  assign n52946 = ~pi213 & ~n52945;
  assign n52947 = ~n52786 & n52946;
  assign n52948 = ~pi212 & ~n52734;
  assign n52949 = ~n45447 & ~n52591;
  assign n52950 = pi214 & ~n52949;
  assign n52951 = n52948 & ~n52950;
  assign n52952 = pi214 & n52597;
  assign n52953 = pi212 & ~n52952;
  assign n52954 = ~pi214 & ~n52949;
  assign n52955 = n52953 & ~n52954;
  assign n52956 = ~n52951 & ~n52955;
  assign n52957 = ~pi219 & ~n52956;
  assign n52958 = n61224 & ~n52685;
  assign n52959 = ~n52957 & n52958;
  assign n52960 = ~pi1150 & ~n51578;
  assign n52961 = pi219 & ~n52651;
  assign n52962 = n61276 & ~n52961;
  assign n52963 = ~n52672 & n52962;
  assign n52964 = n52960 & ~n52963;
  assign n52965 = ~n52959 & n52964;
  assign n52966 = ~n52735 & n52948;
  assign n52967 = ~pi214 & ~n52595;
  assign n52968 = n52953 & ~n52967;
  assign n52969 = ~n52966 & ~n52968;
  assign n52970 = ~pi219 & ~n52969;
  assign n52971 = ~n52685 & ~n52970;
  assign n52972 = ~pi1147 & ~n52971;
  assign n52973 = n52655 & ~n52665;
  assign n52974 = ~pi214 & ~n61273;
  assign n52975 = n52669 & ~n52974;
  assign n52976 = ~n52973 & ~n52975;
  assign n52977 = ~pi219 & ~n52976;
  assign n52978 = ~n52961 & ~n52977;
  assign n52979 = pi1147 & ~n52978;
  assign n52980 = n58992 & ~n52979;
  assign n52981 = ~n52972 & n52980;
  assign n52982 = pi1150 & ~n51203;
  assign n52983 = ~n52981 & n52982;
  assign n52984 = ~n52965 & ~n52983;
  assign n52985 = pi1149 & ~n52984;
  assign n52986 = pi1150 & n61196;
  assign n52987 = ~pi1147 & n52594;
  assign n52988 = n44774 & ~n52987;
  assign n52989 = n52986 & ~n52988;
  assign n52990 = pi1147 & ~n52651;
  assign n52991 = n52591 & ~n52986;
  assign n52992 = ~pi1147 & ~n52991;
  assign n52993 = n58992 & ~n52992;
  assign n52994 = ~n52990 & n52993;
  assign n52995 = ~pi1149 & ~n52994;
  assign n52996 = ~n52989 & n52995;
  assign n52997 = ~pi1148 & ~n52996;
  assign n52998 = ~n52985 & n52997;
  assign n52999 = n52607 & ~n52711;
  assign n53000 = n61224 & ~n52999;
  assign n53001 = ~pi219 & ~n61270;
  assign n53002 = ~pi219 & n52690;
  assign n53003 = ~n61246 & n53001;
  assign n53004 = n53000 & ~n61288;
  assign n53005 = ~n49343 & n52666;
  assign n53006 = n52642 & ~n53005;
  assign n53007 = n4441 & ~n53006;
  assign n53008 = n52723 & n53007;
  assign n53009 = n61276 & ~n53006;
  assign n53010 = pi214 & ~n45447;
  assign n53011 = ~n61271 & n53010;
  assign n53012 = pi212 & ~n53011;
  assign n53013 = ~n52631 & n53012;
  assign n53014 = ~pi212 & n61271;
  assign n53015 = ~pi219 & ~n53014;
  assign n53016 = ~n53013 & n53015;
  assign n53017 = n61289 & ~n53016;
  assign n53018 = ~pi1150 & ~n51232;
  assign n53019 = ~n53017 & n53018;
  assign n53020 = ~n53004 & n53018;
  assign n53021 = ~n53017 & n53020;
  assign n53022 = ~n53004 & n53019;
  assign n53023 = pi214 & n52949;
  assign n53024 = ~n61270 & n52949;
  assign n53025 = pi214 & n53024;
  assign n53026 = ~n61270 & n53023;
  assign n53027 = n52603 & ~n61291;
  assign n53028 = n52600 & ~n53027;
  assign n53029 = n53000 & ~n53028;
  assign n53030 = ~pi214 & n52667;
  assign n53031 = n53012 & ~n53030;
  assign n53032 = n52632 & ~n52667;
  assign n53033 = ~pi219 & ~n53032;
  assign n53034 = ~pi219 & ~n53031;
  assign n53035 = ~n53032 & n53034;
  assign n53036 = ~n53031 & n53033;
  assign n53037 = n61289 & ~n61292;
  assign n53038 = pi1150 & ~n51466;
  assign n53039 = ~n53037 & n53038;
  assign n53040 = ~n53029 & n53039;
  assign n53041 = ~n61290 & ~n53040;
  assign n53042 = ~pi1149 & ~n53041;
  assign n53043 = pi212 & n52735;
  assign n53044 = ~n49343 & ~n52949;
  assign n53045 = n53001 & ~n53044;
  assign n53046 = ~n52735 & n53024;
  assign n53047 = pi212 & ~n53046;
  assign n53048 = n52589 & ~n61291;
  assign n53049 = ~pi219 & ~n53048;
  assign n53050 = ~n53047 & n53049;
  assign n53051 = ~n53043 & n53045;
  assign n53052 = n53000 & ~n61293;
  assign n53053 = n52635 & ~n52636;
  assign n53054 = ~n53006 & ~n53053;
  assign n53055 = n4441 & n53054;
  assign n53056 = n53007 & ~n53053;
  assign n53057 = ~n52265 & n52723;
  assign n53058 = ~n52265 & n61276;
  assign n53059 = n53054 & n53058;
  assign n53060 = n61294 & n53057;
  assign n53061 = ~n51539 & ~n61295;
  assign n53062 = ~n53052 & n53061;
  assign n53063 = ~pi1150 & ~n53062;
  assign n53064 = ~n4441 & ~n49761;
  assign n53065 = n52723 & ~n53064;
  assign n53066 = ~n61294 & n53065;
  assign n53067 = n4441 & ~n49760;
  assign n53068 = n52606 & n53067;
  assign n53069 = ~n49761 & ~n61275;
  assign n53070 = n51841 & ~n53064;
  assign n53071 = ~n53069 & n53070;
  assign n53072 = ~n53068 & n53071;
  assign n53073 = pi57 & n49761;
  assign n53074 = pi1150 & ~n53073;
  assign n53075 = ~n53072 & n53074;
  assign n53076 = ~n53066 & n53075;
  assign n53077 = pi1149 & ~n53076;
  assign n53078 = ~n53063 & n53077;
  assign n53079 = pi1148 & ~n53078;
  assign n53080 = ~n53042 & n53079;
  assign n53081 = ~pi209 & ~n53080;
  assign n53082 = ~n52998 & n53081;
  assign n53083 = n50191 & ~n51492;
  assign n53084 = ~pi1150 & n51580;
  assign n53085 = ~n51577 & n52960;
  assign n53086 = pi1150 & n51605;
  assign n53087 = pi1149 & ~n53086;
  assign n53088 = ~n61296 & n53087;
  assign n53089 = ~n53083 & ~n53088;
  assign n53090 = ~pi1148 & ~n53089;
  assign n53091 = pi1150 & ~n51488;
  assign n53092 = ~pi1150 & ~n51529;
  assign n53093 = ~pi1149 & ~n53092;
  assign n53094 = ~n53091 & n53093;
  assign n53095 = ~pi1150 & ~n61205;
  assign n53096 = pi1150 & ~n51612;
  assign n53097 = pi1149 & ~n53096;
  assign n53098 = ~n53095 & n53097;
  assign n53099 = pi1148 & ~n53098;
  assign n53100 = ~pi1150 & n61205;
  assign n53101 = pi1150 & n51612;
  assign n53102 = pi1149 & ~n53101;
  assign n53103 = pi1149 & ~n53100;
  assign n53104 = ~n53101 & n53103;
  assign n53105 = ~n53100 & n53102;
  assign n53106 = pi1150 & n51488;
  assign n53107 = ~pi1150 & n51529;
  assign n53108 = ~pi1149 & ~n53107;
  assign n53109 = ~n53106 & n53108;
  assign n53110 = ~n61297 & ~n53109;
  assign n53111 = pi1148 & ~n53110;
  assign n53112 = ~n53094 & n53099;
  assign n53113 = ~n53090 & ~n61298;
  assign n53114 = pi209 & n53113;
  assign n53115 = pi213 & ~n53114;
  assign n53116 = ~n53082 & n53115;
  assign n53117 = ~pi213 & n61287;
  assign n53118 = pi213 & ~n53113;
  assign n53119 = pi209 & ~n53118;
  assign n53120 = ~n53117 & n53119;
  assign n53121 = ~n52985 & ~n52996;
  assign n53122 = ~pi1148 & ~n53121;
  assign n53123 = ~pi1149 & ~n61290;
  assign n53124 = ~n53040 & n53123;
  assign n53125 = ~pi1150 & ~n51539;
  assign n53126 = ~n61295 & n53125;
  assign n53127 = ~n53052 & n53126;
  assign n53128 = ~n53072 & ~n53073;
  assign n53129 = ~n53066 & n53128;
  assign n53130 = pi1150 & ~n53129;
  assign n53131 = pi1149 & ~n53130;
  assign n53132 = pi1149 & ~n53127;
  assign n53133 = ~n53130 & n53132;
  assign n53134 = ~n53127 & n53131;
  assign n53135 = pi1148 & ~n61299;
  assign n53136 = ~n53124 & n53135;
  assign n53137 = pi213 & ~n53136;
  assign n53138 = ~n53122 & n53137;
  assign n53139 = ~pi213 & ~n52700;
  assign n53140 = ~pi209 & ~n53139;
  assign n53141 = ~n53138 & n53140;
  assign n53142 = ~n53120 & ~n53141;
  assign n53143 = ~n52947 & ~n53116;
  assign n53144 = pi230 & n61300;
  assign n53145 = ~pi230 & pi246;
  assign n53146 = pi230 & ~n61300;
  assign n53147 = ~pi230 & ~pi246;
  assign n53148 = ~n53146 & ~n53147;
  assign n53149 = ~n53144 & ~n53145;
  assign n53150 = ~pi1147 & ~n52288;
  assign n53151 = pi1151 & ~n51578;
  assign n53152 = ~n51586 & ~n52853;
  assign n53153 = n53151 & ~n53152;
  assign n53154 = n53150 & ~n53153;
  assign n53155 = n51555 & ~n51572;
  assign n53156 = ~n52871 & ~n53155;
  assign n53157 = ~n51539 & ~n53156;
  assign n53158 = ~pi1151 & n53157;
  assign n53159 = n51681 & ~n52859;
  assign n53160 = pi1151 & ~n51539;
  assign n53161 = ~n53159 & n53160;
  assign n53162 = pi1147 & ~n53161;
  assign n53163 = ~n53158 & n53162;
  assign n53164 = ~pi1149 & ~n53163;
  assign n53165 = ~n53154 & n53164;
  assign n53166 = ~pi1151 & ~n51203;
  assign n53167 = n51519 & ~n52907;
  assign n53168 = n61247 & ~n53167;
  assign n53169 = ~n51505 & n61247;
  assign n53170 = ~n53168 & ~n53169;
  assign n53171 = n53166 & n53170;
  assign n53172 = n52047 & ~n61285;
  assign n53173 = ~pi1147 & ~n53172;
  assign n53174 = ~n53171 & n53173;
  assign n53175 = pi1147 & ~n52302;
  assign n53176 = ~n51541 & ~n51611;
  assign n53177 = n52250 & n53176;
  assign n53178 = n53175 & ~n53177;
  assign n53179 = pi1149 & ~n53178;
  assign n53180 = ~n53174 & n53179;
  assign n53181 = pi1150 & ~n53180;
  assign n53182 = ~n53165 & n53181;
  assign n53183 = pi212 & ~n51153;
  assign n53184 = n52793 & ~n53183;
  assign n53185 = n51486 & ~n53184;
  assign n53186 = n51970 & ~n53185;
  assign n53187 = pi1147 & ~n53186;
  assign n53188 = n61092 & ~n51500;
  assign n53189 = ~n51510 & ~n53188;
  assign n53190 = ~n51510 & n61244;
  assign n53191 = ~n53188 & n53190;
  assign n53192 = n61244 & n53189;
  assign n53193 = ~pi1151 & ~n51611;
  assign n53194 = ~n61302 & n53193;
  assign n53195 = ~n51527 & n53194;
  assign n53196 = n53187 & ~n53195;
  assign n53197 = ~n52050 & n52793;
  assign n53198 = n51632 & ~n53197;
  assign n53199 = ~n51203 & ~n53198;
  assign n53200 = pi1151 & n53199;
  assign n53201 = n52047 & ~n53198;
  assign n53202 = n53166 & ~n61302;
  assign n53203 = ~pi1147 & ~n53202;
  assign n53204 = ~n61303 & n53203;
  assign n53205 = pi1149 & ~n53204;
  assign n53206 = ~n53196 & n53205;
  assign n53207 = ~n52181 & n53160;
  assign n53208 = pi1147 & ~n52299;
  assign n53209 = ~n53207 & n53208;
  assign n53210 = n49295 & ~n61119;
  assign n53211 = ~pi1151 & ~n53210;
  assign n53212 = ~pi1147 & ~n53211;
  assign n53213 = n51323 & ~n52000;
  assign n53214 = n53151 & ~n53213;
  assign n53215 = n53212 & ~n53214;
  assign n53216 = ~pi1149 & ~n53215;
  assign n53217 = ~n53209 & n53216;
  assign n53218 = ~pi1150 & ~n53217;
  assign n53219 = ~n53206 & n53218;
  assign n53220 = ~n53182 & ~n53219;
  assign n53221 = pi1148 & ~n53220;
  assign n53222 = pi1147 & ~n52295;
  assign n53223 = ~pi1151 & ~n51466;
  assign n53224 = ~n51527 & n53223;
  assign n53225 = n53222 & ~n53224;
  assign n53226 = pi1151 & ~n61197;
  assign n53227 = ~n51481 & n51632;
  assign n53228 = ~n61197 & ~n53227;
  assign n53229 = pi1151 & n53228;
  assign n53230 = n53226 & ~n53227;
  assign n53231 = ~pi1151 & ~n61197;
  assign n53232 = ~n52233 & n53231;
  assign n53233 = ~pi1147 & ~n53232;
  assign n53234 = ~n61304 & n53233;
  assign n53235 = ~n53225 & ~n53234;
  assign n53236 = ~pi1150 & ~n53235;
  assign n53237 = n52019 & n52247;
  assign n53238 = pi1147 & ~n53237;
  assign n53239 = ~n51466 & ~n51526;
  assign n53240 = ~pi1151 & n53239;
  assign n53241 = n53238 & ~n53240;
  assign n53242 = ~n53168 & n53231;
  assign n53243 = ~n51715 & n53226;
  assign n53244 = ~pi1147 & ~n53243;
  assign n53245 = ~n53242 & n53244;
  assign n53246 = ~n53241 & ~n53245;
  assign n53247 = pi1150 & ~n53246;
  assign n53248 = pi1149 & ~n53247;
  assign n53249 = ~pi1150 & ~n53234;
  assign n53250 = ~n53225 & n53249;
  assign n53251 = pi1150 & ~n53245;
  assign n53252 = pi1150 & ~n53241;
  assign n53253 = ~n53245 & n53252;
  assign n53254 = ~n53241 & n53251;
  assign n53255 = ~n53250 & ~n61305;
  assign n53256 = pi1149 & ~n53255;
  assign n53257 = ~n53236 & n53248;
  assign n53258 = ~n61282 & n53159;
  assign n53259 = n51233 & ~n53258;
  assign n53260 = ~n51232 & ~n52874;
  assign n53261 = ~pi1151 & n53260;
  assign n53262 = pi1147 & ~n53261;
  assign n53263 = ~n53259 & n53262;
  assign n53264 = ~pi1151 & ~n51736;
  assign n53265 = ~pi1147 & ~n53264;
  assign n53266 = pi1151 & ~n51585;
  assign n53267 = n53265 & ~n53266;
  assign n53268 = pi1150 & ~n53267;
  assign n53269 = ~n53263 & n53268;
  assign n53270 = ~n51106 & n52245;
  assign n53271 = n52179 & ~n53270;
  assign n53272 = n51233 & ~n53271;
  assign n53273 = n52028 & ~n52246;
  assign n53274 = pi1147 & ~n53273;
  assign n53275 = ~n53272 & n53274;
  assign n53276 = ~pi1147 & pi1151;
  assign n53277 = n51490 & n53276;
  assign n53278 = ~pi1150 & ~n53277;
  assign n53279 = ~n53275 & n53278;
  assign n53280 = ~n53269 & ~n53279;
  assign n53281 = ~pi1149 & ~n53280;
  assign n53282 = ~pi1148 & ~n53281;
  assign n53283 = ~n61306 & n53282;
  assign n53284 = ~n61306 & ~n53281;
  assign n53285 = ~pi1148 & ~n53284;
  assign n53286 = pi1148 & ~n53219;
  assign n53287 = ~n53182 & n53286;
  assign n53288 = ~n53285 & ~n53287;
  assign n53289 = ~n53221 & ~n53283;
  assign n53290 = ~pi213 & ~n61307;
  assign n53291 = pi213 & ~n52307;
  assign n53292 = pi209 & ~n53291;
  assign n53293 = ~n53290 & n53292;
  assign n53294 = ~pi219 & ~n51997;
  assign n53295 = ~n51997 & n52204;
  assign n53296 = ~n52203 & n53294;
  assign n53297 = n51486 & ~n61308;
  assign n53298 = ~n51482 & n53297;
  assign n53299 = n52028 & ~n53298;
  assign n53300 = n53222 & ~n53299;
  assign n53301 = n51120 & n51323;
  assign n53302 = ~n36621 & n53301;
  assign n53303 = ~n53271 & ~n53302;
  assign n53304 = n52019 & n53303;
  assign n53305 = n52028 & ~n53271;
  assign n53306 = ~pi1147 & ~n53305;
  assign n53307 = ~n53304 & n53306;
  assign n53308 = ~pi1150 & ~n53307;
  assign n53309 = ~n53300 & n53308;
  assign n53310 = ~n51539 & ~n53297;
  assign n53311 = ~pi1151 & n53310;
  assign n53312 = n53187 & ~n53311;
  assign n53313 = n51970 & ~n53301;
  assign n53314 = ~n52181 & n53313;
  assign n53315 = n51978 & ~n52181;
  assign n53316 = ~pi1147 & ~n53315;
  assign n53317 = ~pi1147 & ~n53314;
  assign n53318 = ~n53315 & n53317;
  assign n53319 = ~n53314 & n53316;
  assign n53320 = pi1150 & ~n61309;
  assign n53321 = ~n53312 & n53320;
  assign n53322 = ~n53309 & ~n53321;
  assign n53323 = pi1149 & ~n53322;
  assign n53324 = ~n61197 & ~n52233;
  assign n53325 = ~pi1151 & ~n52808;
  assign n53326 = pi1147 & ~n53325;
  assign n53327 = ~n53324 & n53326;
  assign n53328 = n51491 & n53276;
  assign n53329 = ~pi1150 & ~n53328;
  assign n53330 = ~n53327 & n53329;
  assign n53331 = n51512 & n61244;
  assign n53332 = ~n51578 & ~n53331;
  assign n53333 = ~pi1151 & n53332;
  assign n53334 = n52071 & ~n53331;
  assign n53335 = n52047 & ~n61302;
  assign n53336 = pi1147 & ~n53335;
  assign n53337 = ~n61310 & n53336;
  assign n53338 = ~n44774 & n51202;
  assign n53339 = pi1151 & ~n53338;
  assign n53340 = n53212 & ~n53339;
  assign n53341 = pi1150 & ~n53340;
  assign n53342 = ~n53337 & n53341;
  assign n53343 = ~n53330 & ~n53342;
  assign n53344 = ~pi1149 & ~n53343;
  assign n53345 = ~pi1148 & ~n53344;
  assign n53346 = ~n53323 & n53345;
  assign n53347 = n51569 & n51576;
  assign n53348 = n52047 & ~n53347;
  assign n53349 = n53150 & ~n53348;
  assign n53350 = n52047 & n53170;
  assign n53351 = n52071 & ~n53169;
  assign n53352 = pi1147 & ~n53351;
  assign n53353 = ~n53350 & n53352;
  assign n53354 = pi1150 & ~n53353;
  assign n53355 = ~n53349 & n53354;
  assign n53356 = ~n53168 & n53226;
  assign n53357 = pi1147 & ~n52250;
  assign n53358 = ~n53356 & n53357;
  assign n53359 = n58992 & ~n52149;
  assign n53360 = ~n52152 & n53359;
  assign n53361 = ~n52092 & ~n53360;
  assign n53362 = n53265 & n53361;
  assign n53363 = ~pi1150 & ~n53362;
  assign n53364 = ~n53358 & n53363;
  assign n53365 = ~pi1149 & ~n53364;
  assign n53366 = ~n53355 & n53365;
  assign n53367 = n52028 & ~n53258;
  assign n53368 = ~n51466 & ~n52867;
  assign n53369 = pi1151 & n53368;
  assign n53370 = ~pi1147 & ~n53369;
  assign n53371 = ~n53367 & n53370;
  assign n53372 = ~n51608 & n53273;
  assign n53373 = n53238 & ~n53372;
  assign n53374 = ~pi1150 & ~n53373;
  assign n53375 = ~n53371 & n53374;
  assign n53376 = n51978 & ~n53159;
  assign n53377 = n51596 & ~n51687;
  assign n53378 = n51681 & ~n53377;
  assign n53379 = n51970 & ~n53378;
  assign n53380 = ~pi1147 & ~n53379;
  assign n53381 = ~n53376 & n53380;
  assign n53382 = ~n51539 & ~n52266;
  assign n53383 = ~pi1151 & n53382;
  assign n53384 = n53175 & ~n53383;
  assign n53385 = pi1150 & ~n53384;
  assign n53386 = ~n53381 & n53385;
  assign n53387 = pi1149 & ~n53386;
  assign n53388 = ~n53375 & n53387;
  assign n53389 = ~n53366 & ~n53388;
  assign n53390 = ~n53355 & ~n53364;
  assign n53391 = ~pi1149 & ~n53390;
  assign n53392 = ~n53375 & ~n53386;
  assign n53393 = pi1149 & ~n53392;
  assign n53394 = pi1148 & ~n53393;
  assign n53395 = ~n53391 & n53394;
  assign n53396 = pi1148 & ~n53389;
  assign n53397 = pi213 & ~n61311;
  assign n53398 = ~n53346 & n53397;
  assign n53399 = ~pi213 & n51626;
  assign n53400 = ~pi209 & ~n53399;
  assign n53401 = ~n53398 & n53400;
  assign n53402 = ~pi213 & n61307;
  assign n53403 = pi213 & n52307;
  assign n53404 = pi209 & ~n53403;
  assign n53405 = ~n53402 & n53404;
  assign n53406 = ~n53346 & ~n61311;
  assign n53407 = pi213 & ~n53406;
  assign n53408 = ~pi213 & ~n51626;
  assign n53409 = ~pi209 & ~n53408;
  assign n53410 = ~n53407 & n53409;
  assign n53411 = ~n53405 & ~n53410;
  assign n53412 = ~n53293 & ~n53401;
  assign n53413 = pi230 & n61312;
  assign n53414 = ~pi230 & pi247;
  assign n53415 = pi230 & ~n61312;
  assign n53416 = ~pi230 & ~pi247;
  assign n53417 = ~n53415 & ~n53416;
  assign n53418 = ~n53413 & ~n53414;
  assign n53419 = ~n51577 & n53151;
  assign n53420 = ~pi1152 & ~n53419;
  assign n53421 = ~n53211 & n53420;
  assign n53422 = n52071 & ~n53213;
  assign n53423 = pi1152 & ~n53422;
  assign n53424 = ~n53153 & n53423;
  assign n53425 = ~pi1150 & ~n53424;
  assign n53426 = ~n53421 & n53425;
  assign n53427 = ~pi1152 & ~n53202;
  assign n53428 = ~n53350 & n53427;
  assign n53429 = ~pi1151 & n53199;
  assign n53430 = n53166 & ~n53198;
  assign n53431 = pi1152 & ~n53172;
  assign n53432 = ~n61314 & n53431;
  assign n53433 = pi1150 & ~n53432;
  assign n53434 = pi1150 & ~n53428;
  assign n53435 = ~n53432 & n53434;
  assign n53436 = ~n53428 & n53433;
  assign n53437 = ~pi1148 & ~n61315;
  assign n53438 = ~n53426 & n53437;
  assign n53439 = pi1152 & ~n52302;
  assign n53440 = ~n53185 & n53193;
  assign n53441 = n53439 & ~n53440;
  assign n53442 = pi1151 & ~n51521;
  assign n53443 = n53176 & n53442;
  assign n53444 = ~pi1152 & ~n53443;
  assign n53445 = ~n53195 & n53444;
  assign n53446 = pi1150 & ~n53445;
  assign n53447 = ~n53441 & n53446;
  assign n53448 = pi1151 & n53157;
  assign n53449 = ~pi1152 & ~n52299;
  assign n53450 = ~n53448 & n53449;
  assign n53451 = pi1152 & ~n53315;
  assign n53452 = ~n53161 & n53451;
  assign n53453 = ~pi1150 & ~n53452;
  assign n53454 = ~pi1150 & ~n53450;
  assign n53455 = ~n53452 & n53454;
  assign n53456 = ~n53450 & n53453;
  assign n53457 = pi1148 & ~n61316;
  assign n53458 = pi1148 & ~n53447;
  assign n53459 = ~n61316 & n53458;
  assign n53460 = ~n53447 & n53457;
  assign n53461 = ~n53438 & ~n61317;
  assign n53462 = pi1149 & ~n53461;
  assign n53463 = ~pi1151 & n51488;
  assign n53464 = ~n51487 & n53223;
  assign n53465 = pi1152 & ~n61318;
  assign n53466 = ~n53237 & n53465;
  assign n53467 = pi1151 & n53239;
  assign n53468 = ~pi1152 & ~n53224;
  assign n53469 = ~n53467 & n53468;
  assign n53470 = ~n53466 & ~n53469;
  assign n53471 = pi1150 & ~n53470;
  assign n53472 = ~n53259 & ~n53305;
  assign n53473 = pi1152 & ~n53472;
  assign n53474 = pi1151 & n53260;
  assign n53475 = ~n53273 & ~n53474;
  assign n53476 = ~pi1152 & ~n53475;
  assign n53477 = ~pi1150 & ~n53476;
  assign n53478 = ~n53473 & n53477;
  assign n53479 = pi1148 & ~n53478;
  assign n53480 = ~n53471 & n53479;
  assign n53481 = ~pi1151 & n53228;
  assign n53482 = ~n53227 & n53231;
  assign n53483 = pi1152 & ~n53243;
  assign n53484 = ~n61319 & n53483;
  assign n53485 = ~pi1152 & ~n53232;
  assign n53486 = ~n53356 & n53485;
  assign n53487 = pi1150 & ~n53486;
  assign n53488 = ~n53484 & n53487;
  assign n53489 = pi1151 & ~pi1152;
  assign n53490 = n51736 & n53489;
  assign n53491 = ~pi1151 & ~n51490;
  assign n53492 = pi1152 & ~n53266;
  assign n53493 = ~n53491 & n53492;
  assign n53494 = ~pi1150 & ~n53493;
  assign n53495 = ~pi1150 & ~n53490;
  assign n53496 = ~n53493 & n53495;
  assign n53497 = ~n53490 & n53494;
  assign n53498 = ~n53488 & ~n61320;
  assign n53499 = ~pi1148 & ~n53498;
  assign n53500 = ~pi1149 & ~n53499;
  assign n53501 = ~n53480 & n53500;
  assign n53502 = ~n53471 & ~n53478;
  assign n53503 = pi1148 & ~n53502;
  assign n53504 = ~pi1148 & ~n61320;
  assign n53505 = ~n53488 & n53504;
  assign n53506 = ~pi1149 & ~n53505;
  assign n53507 = ~n53503 & n53506;
  assign n53508 = pi1149 & ~n61317;
  assign n53509 = ~n53438 & n53508;
  assign n53510 = ~n53507 & ~n53509;
  assign n53511 = ~n53462 & ~n53501;
  assign n53512 = ~pi213 & ~n61321;
  assign n53513 = ~n51580 & n53489;
  assign n53514 = ~pi1151 & ~n51491;
  assign n53515 = ~n51490 & n53514;
  assign n53516 = pi1152 & ~n53515;
  assign n53517 = ~n52289 & n53516;
  assign n53518 = ~pi1150 & ~n53517;
  assign n53519 = ~n53513 & n53518;
  assign n53520 = ~n52302 & n53465;
  assign n53521 = n53439 & ~n61318;
  assign n53522 = pi1151 & n61205;
  assign n53523 = ~pi1152 & ~n53522;
  assign n53524 = ~n52296 & n53523;
  assign n53525 = pi1150 & ~n53524;
  assign n53526 = ~n61322 & n53525;
  assign n53527 = ~n53513 & ~n53517;
  assign n53528 = ~pi1150 & ~n53527;
  assign n53529 = ~n61322 & ~n53524;
  assign n53530 = pi1150 & ~n53529;
  assign n53531 = ~n53528 & ~n53530;
  assign n53532 = ~n53519 & ~n53526;
  assign n53533 = pi213 & n61323;
  assign n53534 = pi209 & ~n53533;
  assign n53535 = ~n53512 & n53534;
  assign n53536 = ~n53186 & n53465;
  assign n53537 = pi1151 & n53310;
  assign n53538 = ~pi1152 & ~n53299;
  assign n53539 = ~n53537 & n53538;
  assign n53540 = ~n53536 & ~n53539;
  assign n53541 = pi1150 & ~n53540;
  assign n53542 = pi1151 & n53332;
  assign n53543 = n53151 & ~n53331;
  assign n53544 = ~pi1152 & ~n53325;
  assign n53545 = ~n61324 & n53544;
  assign n53546 = pi1152 & ~n53232;
  assign n53547 = ~n53335 & n53546;
  assign n53548 = ~n53545 & ~n53547;
  assign n53549 = ~pi1150 & ~n53548;
  assign n53550 = ~pi1149 & ~n53549;
  assign n53551 = ~n53541 & n53550;
  assign n53552 = pi1152 & ~n53242;
  assign n53553 = ~n53350 & n53552;
  assign n53554 = n53151 & ~n53169;
  assign n53555 = n52251 & ~n53554;
  assign n53556 = ~pi1150 & ~n53555;
  assign n53557 = ~n53553 & n53556;
  assign n53558 = n52247 & n53223;
  assign n53559 = n53439 & ~n53558;
  assign n53560 = pi1151 & n53382;
  assign n53561 = ~pi1152 & ~n53372;
  assign n53562 = ~n53560 & n53561;
  assign n53563 = pi1150 & ~n53562;
  assign n53564 = ~n53559 & n53563;
  assign n53565 = ~n53557 & ~n53564;
  assign n53566 = pi1149 & ~n53565;
  assign n53567 = pi1148 & ~n53566;
  assign n53568 = ~n53551 & n53567;
  assign n53569 = n53223 & n53303;
  assign n53570 = pi1152 & ~n53314;
  assign n53571 = ~n53569 & n53570;
  assign n53572 = ~pi1152 & ~n53305;
  assign n53573 = ~n53207 & n53572;
  assign n53574 = pi1150 & ~n53573;
  assign n53575 = ~n53571 & n53574;
  assign n53576 = pi1152 & ~n53339;
  assign n53577 = ~n53514 & n53576;
  assign n53578 = n53210 & n53489;
  assign n53579 = ~pi1150 & ~n53578;
  assign n53580 = ~n53577 & n53579;
  assign n53581 = ~pi1149 & ~n53580;
  assign n53582 = ~n53575 & n53581;
  assign n53583 = ~n53264 & n53420;
  assign n53584 = ~pi1151 & ~n53361;
  assign n53585 = pi1152 & ~n53584;
  assign n53586 = ~n53348 & n53585;
  assign n53587 = ~pi1150 & ~n53586;
  assign n53588 = ~n53583 & n53587;
  assign n53589 = ~pi1152 & ~n53161;
  assign n53590 = ~n53367 & n53589;
  assign n53591 = ~pi1151 & n53368;
  assign n53592 = pi1152 & ~n53379;
  assign n53593 = ~n53591 & n53592;
  assign n53594 = pi1150 & ~n53593;
  assign n53595 = ~n53590 & n53594;
  assign n53596 = pi1149 & ~n53595;
  assign n53597 = ~n53588 & n53596;
  assign n53598 = ~n53582 & ~n53597;
  assign n53599 = ~pi1148 & ~n53598;
  assign n53600 = pi213 & ~n53599;
  assign n53601 = ~n53568 & n53600;
  assign n53602 = ~pi213 & n53113;
  assign n53603 = ~pi209 & ~n53602;
  assign n53604 = ~n53601 & n53603;
  assign n53605 = ~pi213 & n61321;
  assign n53606 = pi213 & ~n61323;
  assign n53607 = pi209 & ~n53606;
  assign n53608 = ~n53605 & n53607;
  assign n53609 = pi1150 & ~n53539;
  assign n53610 = pi1150 & ~n53536;
  assign n53611 = ~n53539 & n53610;
  assign n53612 = ~n53536 & n53609;
  assign n53613 = ~pi1150 & ~n53547;
  assign n53614 = ~n53545 & n53613;
  assign n53615 = ~pi1149 & ~n53614;
  assign n53616 = ~n61325 & n53615;
  assign n53617 = pi1149 & ~n53564;
  assign n53618 = ~n53557 & n53617;
  assign n53619 = pi1148 & ~n53618;
  assign n53620 = ~n53616 & n53619;
  assign n53621 = ~pi1148 & ~n53582;
  assign n53622 = ~n53597 & n53621;
  assign n53623 = pi213 & ~n53622;
  assign n53624 = pi213 & ~n53620;
  assign n53625 = ~n53622 & n53624;
  assign n53626 = ~n53620 & n53623;
  assign n53627 = ~pi213 & ~n53113;
  assign n53628 = ~pi209 & ~n53627;
  assign n53629 = ~n61326 & n53628;
  assign n53630 = ~n53608 & ~n53629;
  assign n53631 = ~n53535 & ~n53604;
  assign n53632 = pi230 & n61327;
  assign n53633 = ~pi230 & pi248;
  assign n53634 = pi230 & ~n61327;
  assign n53635 = ~pi230 & ~pi248;
  assign n53636 = ~n53634 & ~n53635;
  assign n53637 = ~n53632 & ~n53633;
  assign n53638 = pi209 & ~n50704;
  assign n53639 = pi57 & ~n50535;
  assign n53640 = pi299 & n50477;
  assign n53641 = ~n52257 & ~n53640;
  assign n53642 = ~pi214 & ~n53641;
  assign n53643 = ~n51080 & n51342;
  assign n53644 = pi212 & ~n53643;
  assign n53645 = ~n53642 & n53644;
  assign n53646 = pi214 & ~n53641;
  assign n53647 = ~pi212 & ~n51109;
  assign n53648 = ~n53646 & n53647;
  assign n53649 = ~pi219 & ~n53648;
  assign n53650 = ~pi219 & ~n53645;
  assign n53651 = ~n53648 & n53650;
  assign n53652 = ~n53645 & n53649;
  assign n53653 = n52254 & ~n61329;
  assign n53654 = ~n4441 & n50535;
  assign n53655 = ~pi57 & pi1151;
  assign n53656 = ~n53654 & n53655;
  assign n53657 = ~n53653 & n53656;
  assign n53658 = pi1151 & ~n53653;
  assign n53659 = ~pi57 & ~n53658;
  assign n53660 = ~n50536 & ~n53659;
  assign n53661 = ~n53639 & ~n53657;
  assign n53662 = ~n51510 & ~n53640;
  assign n53663 = ~n51109 & n53662;
  assign n53664 = ~pi212 & ~n53663;
  assign n53665 = ~pi214 & n53662;
  assign n53666 = ~n45445 & ~n51509;
  assign n53667 = n50518 & ~n53666;
  assign n53668 = pi212 & ~n53667;
  assign n53669 = ~n53665 & n53668;
  assign n53670 = ~n53664 & ~n53669;
  assign n53671 = ~pi219 & ~n53670;
  assign n53672 = n52216 & ~n53671;
  assign n53673 = n47616 & ~n53654;
  assign n53674 = ~n53672 & n53673;
  assign n53675 = ~n61330 & ~n53674;
  assign n53676 = ~pi1152 & ~n53675;
  assign n53677 = ~pi214 & ~n53640;
  assign n53678 = ~n50518 & ~n53677;
  assign n53679 = n51470 & ~n61245;
  assign n53680 = ~n51153 & ~n53640;
  assign n53681 = ~pi214 & ~n53680;
  assign n53682 = pi212 & ~n53681;
  assign n53683 = ~n53679 & n53682;
  assign n53684 = n53183 & ~n53678;
  assign n53685 = n51992 & ~n53640;
  assign n53686 = n52792 & ~n53685;
  assign n53687 = ~n61331 & n53686;
  assign n53688 = ~pi1151 & ~n53687;
  assign n53689 = n51486 & n53688;
  assign n53690 = pi299 & ~n50477;
  assign n53691 = ~n36621 & n53690;
  assign n53692 = ~n50476 & ~n53691;
  assign n53693 = n49392 & ~n53692;
  assign n53694 = n52240 & ~n53693;
  assign n53695 = ~n51524 & ~n51697;
  assign n53696 = pi1151 & ~n53695;
  assign n53697 = ~n53694 & n53696;
  assign n53698 = n50482 & ~n53697;
  assign n53699 = ~n53689 & n53698;
  assign n53700 = pi1150 & ~n53699;
  assign n53701 = ~n53676 & n53700;
  assign n53702 = n36621 & n52151;
  assign n53703 = n50699 & ~n51552;
  assign n53704 = ~n51556 & ~n53640;
  assign n53705 = pi211 & n52150;
  assign n53706 = ~n49584 & n51563;
  assign n53707 = ~n61092 & ~n53706;
  assign n53708 = ~n53705 & n53707;
  assign n53709 = ~n61092 & ~n53705;
  assign n53710 = ~n53706 & n53709;
  assign n53711 = ~n61092 & ~n53704;
  assign n53712 = ~n53703 & ~n61332;
  assign n53713 = ~n53702 & ~n53703;
  assign n53714 = ~n61332 & n53713;
  assign n53715 = ~n53702 & n53712;
  assign n53716 = ~pi219 & ~n61333;
  assign n53717 = pi1151 & n51576;
  assign n53718 = ~n53716 & n53717;
  assign n53719 = ~n51080 & ~n53691;
  assign n53720 = n60971 & n50534;
  assign n53721 = ~n53719 & n53720;
  assign n53722 = n50537 & ~n53721;
  assign n53723 = ~n53718 & n53722;
  assign n53724 = n51587 & ~n53690;
  assign n53725 = pi212 & ~n53724;
  assign n53726 = ~n52139 & n53725;
  assign n53727 = ~pi212 & n51078;
  assign n53728 = ~pi219 & ~n53727;
  assign n53729 = ~n53685 & n53728;
  assign n53730 = ~n53726 & n53729;
  assign n53731 = pi1151 & n51681;
  assign n53732 = n47428 & ~n51680;
  assign n53733 = ~n53730 & n61334;
  assign n53734 = ~pi1151 & n53271;
  assign n53735 = n50482 & ~n53721;
  assign n53736 = ~n53734 & n53735;
  assign n53737 = ~n53733 & n53736;
  assign n53738 = ~pi1150 & ~n53737;
  assign n53739 = ~n53723 & n53738;
  assign n53740 = ~pi209 & ~n53739;
  assign n53741 = ~n53701 & n53740;
  assign n53742 = pi213 & ~n53741;
  assign n53743 = ~n53638 & n53742;
  assign n53744 = ~n36620 & ~n50696;
  assign n53745 = n49582 & ~n50870;
  assign n53746 = ~pi207 & n50869;
  assign n53747 = pi207 & ~n49602;
  assign n53748 = ~n46958 & n53747;
  assign n53749 = pi208 & ~n53748;
  assign n53750 = ~n53746 & n53749;
  assign n53751 = ~n53745 & ~n53750;
  assign n53752 = pi211 & ~n53751;
  assign n53753 = pi214 & n53752;
  assign n53754 = ~n53744 & ~n53753;
  assign n53755 = ~pi212 & ~n53754;
  assign n53756 = ~pi219 & ~n53755;
  assign n53757 = ~pi211 & n53751;
  assign n53758 = ~n50766 & ~n53757;
  assign n53759 = pi214 & ~n53758;
  assign n53760 = ~pi211 & ~n50696;
  assign n53761 = ~pi214 & ~n53760;
  assign n53762 = ~n53752 & n53761;
  assign n53763 = pi212 & ~n53762;
  assign n53764 = ~n53759 & n53763;
  assign n53765 = n53756 & ~n53764;
  assign n53766 = n50698 & ~n53765;
  assign n53767 = n53151 & ~n53766;
  assign n53768 = ~n50696 & n50738;
  assign n53769 = ~n53489 & ~n53768;
  assign n53770 = ~n53767 & ~n53769;
  assign n53771 = pi214 & n50603;
  assign n53772 = n50615 & ~n53771;
  assign n53773 = ~pi219 & ~n53772;
  assign n53774 = pi214 & n61167;
  assign n53775 = ~pi214 & n50603;
  assign n53776 = pi212 & ~n53775;
  assign n53777 = ~n53774 & n53776;
  assign n53778 = n53773 & ~n53777;
  assign n53779 = n58992 & ~n50610;
  assign n53780 = ~n53778 & n53779;
  assign n53781 = n52047 & ~n53780;
  assign n53782 = n61167 & n51272;
  assign n53783 = ~n50593 & ~n51272;
  assign n53784 = n58992 & ~n53783;
  assign n53785 = ~n53782 & n53784;
  assign n53786 = n53231 & ~n53785;
  assign n53787 = pi1152 & ~n53786;
  assign n53788 = ~n53781 & n53787;
  assign n53789 = ~pi1150 & ~n53788;
  assign n53790 = ~n53770 & n53789;
  assign n53791 = ~n50614 & ~n53774;
  assign n53792 = ~pi212 & ~n53791;
  assign n53793 = ~pi211 & n50593;
  assign n53794 = ~n50646 & ~n53793;
  assign n53795 = pi214 & ~n53794;
  assign n53796 = ~pi214 & ~n61167;
  assign n53797 = pi212 & ~n53796;
  assign n53798 = pi212 & ~n53795;
  assign n53799 = ~n53796 & n53798;
  assign n53800 = ~n53795 & n53797;
  assign n53801 = ~n53792 & ~n61335;
  assign n53802 = ~pi219 & ~n53801;
  assign n53803 = n50613 & ~n53802;
  assign n53804 = n53223 & ~n53803;
  assign n53805 = pi212 & ~n50603;
  assign n53806 = n53773 & ~n53805;
  assign n53807 = n50613 & ~n53806;
  assign n53808 = n51970 & ~n53807;
  assign n53809 = pi1152 & ~n53808;
  assign n53810 = ~n53804 & n53809;
  assign n53811 = ~n49343 & n53758;
  assign n53812 = pi219 & ~n50765;
  assign n53813 = ~n53811 & n53812;
  assign n53814 = n58992 & ~n53813;
  assign n53815 = pi214 & n53751;
  assign n53816 = n53763 & ~n53815;
  assign n53817 = n53756 & ~n53816;
  assign n53818 = n53814 & ~n53817;
  assign n53819 = n53160 & ~n53818;
  assign n53820 = pi212 & ~n53754;
  assign n53821 = ~pi212 & ~n50696;
  assign n53822 = ~pi219 & ~n53821;
  assign n53823 = ~n53820 & n53822;
  assign n53824 = n53814 & ~n53823;
  assign n53825 = n52028 & ~n53824;
  assign n53826 = ~pi1152 & ~n53825;
  assign n53827 = ~n53819 & n53826;
  assign n53828 = pi1150 & ~n53827;
  assign n53829 = ~n53810 & n53828;
  assign n53830 = ~n53770 & ~n53788;
  assign n53831 = ~pi1150 & ~n53830;
  assign n53832 = ~n53810 & ~n53827;
  assign n53833 = pi1150 & ~n53832;
  assign n53834 = ~n53831 & ~n53833;
  assign n53835 = ~n53790 & ~n53829;
  assign n53836 = pi209 & n61336;
  assign n53837 = ~pi209 & n61323;
  assign n53838 = ~pi213 & ~n53837;
  assign n53839 = ~n53836 & n53838;
  assign n53840 = ~pi213 & ~n61323;
  assign n53841 = ~n53701 & ~n53739;
  assign n53842 = pi213 & ~n53841;
  assign n53843 = ~pi209 & ~n53842;
  assign n53844 = ~n53840 & n53843;
  assign n53845 = ~pi213 & ~n53790;
  assign n53846 = ~pi213 & ~n61336;
  assign n53847 = ~n53829 & n53845;
  assign n53848 = pi213 & n50704;
  assign n53849 = pi209 & ~n53848;
  assign n53850 = ~n61337 & n53849;
  assign n53851 = ~n53844 & ~n53850;
  assign n53852 = ~n53743 & ~n53839;
  assign n53853 = pi230 & n61338;
  assign n53854 = ~pi230 & pi249;
  assign n53855 = pi230 & ~n61338;
  assign n53856 = ~pi230 & ~pi249;
  assign n53857 = ~n53855 & ~n53856;
  assign n53858 = ~n53853 & ~n53854;
  assign n53859 = ~pi273 & ~n46189;
  assign n53860 = ~n46149 & ~n53859;
  assign n53861 = pi219 & ~n53860;
  assign n53862 = ~pi273 & ~n46158;
  assign n53863 = n46160 & ~n53862;
  assign n53864 = pi1091 & pi1146;
  assign n53865 = ~pi211 & n53864;
  assign n53866 = ~pi219 & ~n53865;
  assign n53867 = ~n53863 & n53866;
  assign n53868 = ~n53861 & ~n53867;
  assign n53869 = pi299 & n53868;
  assign n53870 = ~pi200 & n53864;
  assign n53871 = ~pi199 & ~n53870;
  assign n53872 = ~n53863 & n53871;
  assign n53873 = pi199 & ~n53860;
  assign n53874 = ~pi299 & ~n53873;
  assign n53875 = ~n53872 & n53874;
  assign n53876 = ~n53869 & ~n53875;
  assign n53877 = ~n45427 & ~n46324;
  assign n53878 = pi1091 & ~n53877;
  assign n53879 = n53876 & ~n53878;
  assign n53880 = n58992 & ~n53879;
  assign n53881 = pi1091 & n47539;
  assign n53882 = ~n53880 & ~n53881;
  assign n53883 = pi1147 & ~n53882;
  assign n53884 = ~n58992 & n53868;
  assign n53885 = n61224 & ~n53876;
  assign n53886 = ~pi1148 & ~n53885;
  assign n53887 = pi1091 & n36681;
  assign n53888 = ~n53868 & ~n53887;
  assign n53889 = pi299 & ~n53888;
  assign n53890 = ~pi271 & ~n46188;
  assign n53891 = ~n46147 & ~n53890;
  assign n53892 = pi199 & ~n53891;
  assign n53893 = ~pi1091 & ~n46156;
  assign n53894 = pi271 & ~n53893;
  assign n53895 = ~pi271 & ~n46157;
  assign n53896 = ~n53894 & ~n53895;
  assign n53897 = ~n53864 & ~n53896;
  assign n53898 = ~pi199 & n53897;
  assign n53899 = ~n53892 & ~n53898;
  assign n53900 = pi200 & ~n53899;
  assign n53901 = n46355 & ~n53900;
  assign n53902 = ~n53875 & ~n53901;
  assign n53903 = ~n53889 & n53902;
  assign n53904 = n58992 & ~n53903;
  assign n53905 = n45884 & n47224;
  assign n53906 = pi1148 & ~n53905;
  assign n53907 = ~n53904 & n53906;
  assign n53908 = ~n53886 & ~n53907;
  assign n53909 = ~n53884 & ~n53908;
  assign n53910 = ~n53883 & n53909;
  assign n53911 = ~pi230 & ~n53910;
  assign n53912 = ~pi1146 & n36679;
  assign n53913 = pi1147 & n49295;
  assign n53914 = ~n49298 & ~n53913;
  assign n53915 = ~n53912 & ~n53914;
  assign n53916 = ~pi1146 & n36719;
  assign n53917 = ~pi199 & pi1147;
  assign n53918 = pi200 & ~n53917;
  assign n53919 = ~n53916 & ~n53918;
  assign n53920 = n44774 & n53919;
  assign n53921 = pi1148 & ~n53920;
  assign n53922 = ~n53915 & n53921;
  assign n53923 = ~pi211 & ~n51634;
  assign n53924 = n49295 & ~n53923;
  assign n53925 = n49296 & ~n53916;
  assign n53926 = ~n53924 & ~n53925;
  assign n53927 = pi1147 & ~n53926;
  assign n53928 = pi1146 & ~n61276;
  assign n53929 = ~n45887 & n53928;
  assign n53930 = ~pi1148 & ~n53929;
  assign n53931 = ~n53927 & n53930;
  assign n53932 = pi230 & ~n53931;
  assign n53933 = pi230 & ~n53922;
  assign n53934 = ~n53931 & n53933;
  assign n53935 = ~n53922 & n53932;
  assign n53936 = ~n53911 & ~n61340;
  assign n53937 = pi1147 & n46354;
  assign n53938 = pi1091 & pi1145;
  assign n53939 = n36719 & ~n53938;
  assign n53940 = ~n53896 & n53939;
  assign n53941 = ~n53892 & ~n53940;
  assign n53942 = ~n53937 & ~n53941;
  assign n53943 = ~pi199 & ~n53938;
  assign n53944 = ~n53896 & n53943;
  assign n53945 = ~n53892 & ~n53944;
  assign n53946 = ~pi200 & ~n53937;
  assign n53947 = ~n53945 & n53946;
  assign n53948 = ~n53900 & ~n53947;
  assign n53949 = ~n53900 & ~n53942;
  assign n53950 = n44774 & ~n61341;
  assign n53951 = pi219 & ~n53891;
  assign n53952 = ~n53865 & ~n53897;
  assign n53953 = pi1091 & n49797;
  assign n53954 = ~pi219 & ~n53953;
  assign n53955 = ~n53952 & n53954;
  assign n53956 = ~n53951 & ~n53955;
  assign n53957 = ~pi211 & pi1147;
  assign n53958 = n47224 & n53957;
  assign n53959 = ~n44774 & ~n53958;
  assign n53960 = ~n53956 & n53959;
  assign n53961 = ~n53950 & ~n53960;
  assign n53962 = ~pi230 & ~n53961;
  assign n53963 = ~pi200 & ~n49817;
  assign n53964 = n51788 & ~n53963;
  assign n53965 = ~n51628 & ~n51684;
  assign n53966 = ~pi219 & ~n53965;
  assign n53967 = pi1147 & n47416;
  assign n53968 = ~n53966 & ~n53967;
  assign n53969 = ~n53964 & n53968;
  assign n53970 = n58992 & ~n53969;
  assign n53971 = ~n49797 & n52830;
  assign n53972 = pi219 & ~n53957;
  assign n53973 = ~n58992 & ~n53972;
  assign n53974 = ~n53971 & ~n53972;
  assign n53975 = ~n58992 & n53974;
  assign n53976 = ~n53971 & n53973;
  assign n53977 = pi230 & ~n61342;
  assign n53978 = ~n53970 & n53977;
  assign po428 = ~n53962 & ~n53978;
  assign n53980 = pi264 & ~n46154;
  assign n53981 = ~pi796 & n46154;
  assign n53982 = ~pi1091 & ~n53981;
  assign n53983 = ~pi1091 & ~n53980;
  assign n53984 = ~n53981 & n53983;
  assign n53985 = ~n53980 & n53982;
  assign n53986 = pi1091 & pi1141;
  assign n53987 = ~n61343 & ~n53986;
  assign n53988 = ~pi200 & ~n53987;
  assign n53989 = pi1091 & pi1142;
  assign n53990 = ~n61343 & ~n53989;
  assign n53991 = pi200 & ~n53990;
  assign n53992 = ~pi199 & ~n53991;
  assign n53993 = ~pi199 & ~n53988;
  assign n53994 = ~n53991 & n53993;
  assign n53995 = ~n53988 & n53992;
  assign n53996 = pi264 & ~n46143;
  assign n53997 = ~pi796 & n46143;
  assign n53998 = ~pi1091 & ~n53997;
  assign n53999 = ~pi1091 & ~n53996;
  assign n54000 = ~n53997 & n53999;
  assign n54001 = ~n53996 & n53998;
  assign n54002 = pi1091 & pi1143;
  assign n54003 = ~pi200 & n54002;
  assign n54004 = pi199 & ~n54003;
  assign n54005 = ~n61345 & n54004;
  assign n54006 = n44774 & ~n54005;
  assign n54007 = ~n61344 & n54006;
  assign n54008 = ~pi211 & ~n53987;
  assign n54009 = pi211 & ~n53990;
  assign n54010 = ~pi219 & ~n54009;
  assign n54011 = ~pi219 & ~n54008;
  assign n54012 = ~n54009 & n54011;
  assign n54013 = ~n54008 & n54010;
  assign n54014 = pi219 & ~n46717;
  assign n54015 = ~n49807 & ~n54014;
  assign n54016 = ~n61345 & ~n54015;
  assign n54017 = ~n44774 & ~n54016;
  assign n54018 = ~n61346 & n54017;
  assign n54019 = ~n54007 & ~n54018;
  assign n54020 = ~pi230 & ~n54019;
  assign n54021 = ~pi199 & pi1141;
  assign n54022 = n49812 & ~n54021;
  assign n54023 = ~n49376 & ~n54022;
  assign n54024 = n44774 & ~n54023;
  assign n54025 = ~pi211 & pi1141;
  assign n54026 = ~pi219 & ~n49385;
  assign n54027 = ~n54025 & n54026;
  assign n54028 = ~n49807 & ~n54027;
  assign n54029 = ~n44774 & ~n54028;
  assign n54030 = pi230 & ~n54029;
  assign n54031 = pi230 & ~n54024;
  assign n54032 = ~n54029 & n54031;
  assign n54033 = ~n54024 & n54030;
  assign n54034 = ~n54020 & ~n61347;
  assign n54035 = pi265 & ~n46154;
  assign n54036 = ~pi819 & n46154;
  assign n54037 = ~pi1091 & ~n54036;
  assign n54038 = ~pi1091 & ~n54035;
  assign n54039 = ~n54036 & n54038;
  assign n54040 = ~n54035 & n54037;
  assign n54041 = ~n53989 & ~n61348;
  assign n54042 = ~pi200 & ~n54041;
  assign n54043 = ~n54002 & ~n61348;
  assign n54044 = pi200 & ~n54043;
  assign n54045 = ~pi199 & ~n54044;
  assign n54046 = ~pi199 & ~n54042;
  assign n54047 = ~n54044 & n54046;
  assign n54048 = ~n54042 & n54045;
  assign n54049 = pi265 & ~n46143;
  assign n54050 = ~pi819 & n46143;
  assign n54051 = ~pi1091 & ~n54050;
  assign n54052 = ~pi1091 & ~n54049;
  assign n54053 = ~n54050 & n54052;
  assign n54054 = ~n54049 & n54051;
  assign n54055 = pi1091 & pi1144;
  assign n54056 = ~pi200 & n54055;
  assign n54057 = pi199 & ~n54056;
  assign n54058 = ~n61350 & n54057;
  assign n54059 = n44774 & ~n54058;
  assign n54060 = ~n61349 & n54059;
  assign n54061 = ~pi211 & ~n54041;
  assign n54062 = pi211 & ~n54043;
  assign n54063 = ~pi219 & ~n54062;
  assign n54064 = ~pi219 & ~n54061;
  assign n54065 = ~n54062 & n54064;
  assign n54066 = ~n54061 & n54063;
  assign n54067 = ~n52337 & ~n54014;
  assign n54068 = ~n61350 & ~n54067;
  assign n54069 = ~n44774 & ~n54068;
  assign n54070 = ~n61351 & n54069;
  assign n54071 = ~n54060 & ~n54070;
  assign n54072 = ~pi230 & ~n54071;
  assign n54073 = ~pi219 & ~n49348;
  assign n54074 = ~n49390 & n54073;
  assign n54075 = ~n52337 & ~n54074;
  assign n54076 = ~n44774 & ~n54075;
  assign n54077 = ~n49375 & n52341;
  assign n54078 = ~n49369 & ~n54077;
  assign n54079 = n44774 & ~n54078;
  assign n54080 = pi230 & ~n54079;
  assign n54081 = pi230 & ~n54076;
  assign n54082 = ~n54079 & n54081;
  assign n54083 = ~n54076 & n54080;
  assign n54084 = ~n54072 & ~n61352;
  assign n54085 = ~pi211 & pi1136;
  assign n54086 = pi219 & ~n54085;
  assign n54087 = pi211 & ~pi1135;
  assign n54088 = ~n54086 & ~n54087;
  assign n54089 = ~n36679 & n54088;
  assign n54090 = pi299 & n54089;
  assign n54091 = ~pi199 & pi1135;
  assign n54092 = pi200 & ~n54091;
  assign n54093 = pi199 & pi1136;
  assign n54094 = ~pi200 & ~n54093;
  assign n54095 = ~pi299 & ~n54094;
  assign n54096 = ~pi299 & ~n54092;
  assign n54097 = ~n54094 & n54096;
  assign n54098 = ~n54092 & n54095;
  assign n54099 = ~n54090 & ~n61353;
  assign n54100 = n58992 & ~n54099;
  assign n54101 = ~n58992 & n54089;
  assign n54102 = pi230 & ~n54101;
  assign n54103 = ~n54100 & n54102;
  assign n54104 = ~pi948 & n46154;
  assign n54105 = ~pi266 & ~n46154;
  assign n54106 = ~pi1091 & ~n54105;
  assign n54107 = ~pi1091 & ~n54104;
  assign n54108 = ~n54105 & n54107;
  assign n54109 = ~n54104 & n54106;
  assign n54110 = ~pi199 & ~n61354;
  assign n54111 = pi1091 & pi1136;
  assign n54112 = ~pi948 & n46143;
  assign n54113 = ~pi266 & ~n46143;
  assign n54114 = ~pi1091 & ~n54113;
  assign n54115 = ~pi1091 & ~n54112;
  assign n54116 = ~n54113 & n54115;
  assign n54117 = ~n54112 & n54114;
  assign n54118 = pi199 & ~n61355;
  assign n54119 = ~n54111 & n54118;
  assign n54120 = ~n54110 & ~n54119;
  assign n54121 = ~pi200 & n54120;
  assign n54122 = pi1091 & pi1135;
  assign n54123 = n54110 & ~n54122;
  assign n54124 = pi200 & ~n54118;
  assign n54125 = ~n54123 & n54124;
  assign n54126 = ~n54121 & ~n54125;
  assign n54127 = n44774 & ~n54126;
  assign n54128 = ~n54014 & ~n54086;
  assign n54129 = ~n61355 & ~n54128;
  assign n54130 = ~n44774 & ~n54129;
  assign n54131 = ~pi219 & ~n61354;
  assign n54132 = pi1135 & n46707;
  assign n54133 = n54131 & ~n54132;
  assign n54134 = n54130 & ~n54133;
  assign n54135 = ~pi230 & ~n54134;
  assign n54136 = ~n54127 & n54135;
  assign n54137 = ~n54103 & ~n54136;
  assign n54138 = ~pi1134 & ~n54137;
  assign n54139 = n46359 & ~n54093;
  assign n54140 = ~n54092 & ~n54139;
  assign n54141 = n44774 & n54140;
  assign n54142 = ~n44774 & n54088;
  assign n54143 = pi230 & ~n54142;
  assign n54144 = pi230 & ~n54141;
  assign n54145 = ~n54142 & n54144;
  assign n54146 = ~n54141 & n54143;
  assign n54147 = ~pi199 & pi1091;
  assign n54148 = ~n54120 & ~n54147;
  assign n54149 = ~pi200 & ~n54148;
  assign n54150 = ~n54125 & ~n54149;
  assign n54151 = n44774 & ~n54150;
  assign n54152 = pi1091 & ~n54087;
  assign n54153 = n54131 & ~n54152;
  assign n54154 = n54130 & ~n54153;
  assign n54155 = ~pi230 & ~n54154;
  assign n54156 = ~n54151 & n54155;
  assign n54157 = ~n61356 & ~n54156;
  assign n54158 = pi1134 & ~n54157;
  assign po423 = ~n54138 & ~n54158;
  assign n54160 = pi211 & pi1137;
  assign n54161 = ~n54085 & ~n54160;
  assign n54162 = pi1091 & ~n54161;
  assign n54163 = n49295 & ~n54162;
  assign n54164 = ~pi200 & n54111;
  assign n54165 = pi1137 & n46364;
  assign n54166 = ~n54164 & ~n54165;
  assign n54167 = n49296 & n54166;
  assign n54168 = ~n54163 & ~n54167;
  assign n54169 = pi269 & ~n46154;
  assign n54170 = ~pi817 & n46154;
  assign n54171 = ~pi1091 & ~n54170;
  assign n54172 = ~pi1091 & ~n54169;
  assign n54173 = ~n54170 & n54172;
  assign n54174 = ~n54169 & n54171;
  assign n54175 = ~n54168 & ~n61357;
  assign n54176 = pi219 & ~n44774;
  assign n54177 = pi1138 & n46717;
  assign n54178 = n54176 & ~n54177;
  assign n54179 = ~pi200 & pi1091;
  assign n54180 = pi1138 & n54179;
  assign n54181 = pi199 & ~n54180;
  assign n54182 = n44774 & n54181;
  assign n54183 = ~n54178 & ~n54182;
  assign n54184 = pi269 & ~n46143;
  assign n54185 = ~pi817 & n46143;
  assign n54186 = ~pi1091 & ~n54185;
  assign n54187 = ~pi1091 & ~n54184;
  assign n54188 = ~n54185 & n54187;
  assign n54189 = ~n54184 & n54186;
  assign n54190 = ~n54183 & ~n61358;
  assign n54191 = ~n54175 & ~n54190;
  assign n54192 = ~pi230 & ~n54191;
  assign n54193 = ~pi199 & pi1137;
  assign n54194 = pi200 & ~n54193;
  assign n54195 = ~pi199 & pi1136;
  assign n54196 = pi199 & pi1138;
  assign n54197 = ~pi200 & ~n54196;
  assign n54198 = ~pi200 & ~n54195;
  assign n54199 = ~n54196 & n54198;
  assign n54200 = ~n54195 & n54197;
  assign n54201 = ~n54194 & ~n61359;
  assign n54202 = n44774 & ~n54201;
  assign n54203 = ~pi219 & ~n54161;
  assign n54204 = ~pi211 & pi1138;
  assign n54205 = pi219 & n54204;
  assign n54206 = ~n54203 & ~n54205;
  assign n54207 = ~n44774 & n54206;
  assign n54208 = ~n54202 & ~n54207;
  assign n54209 = pi230 & ~n54208;
  assign po426 = ~n54192 & ~n54209;
  assign n54211 = n46717 & n54025;
  assign n54212 = pi1091 & n54025;
  assign n54213 = n54176 & ~n61360;
  assign n54214 = ~pi200 & n53986;
  assign n54215 = pi199 & ~n54214;
  assign n54216 = n44774 & n54215;
  assign n54217 = ~n54213 & ~n54216;
  assign n54218 = pi270 & ~n46143;
  assign n54219 = ~pi805 & n46143;
  assign n54220 = ~pi1091 & ~n54219;
  assign n54221 = ~pi1091 & ~n54218;
  assign n54222 = ~n54219 & n54221;
  assign n54223 = ~n54218 & n54220;
  assign n54224 = ~n54217 & ~n61361;
  assign n54225 = ~pi211 & pi1139;
  assign n54226 = pi211 & pi1140;
  assign n54227 = ~n54225 & ~n54226;
  assign n54228 = pi1091 & ~n54227;
  assign n54229 = n49295 & ~n54228;
  assign n54230 = pi1091 & pi1140;
  assign n54231 = pi200 & n54230;
  assign n54232 = pi1140 & n46364;
  assign n54233 = pi1139 & n54179;
  assign n54234 = ~n61362 & ~n54233;
  assign n54235 = n49296 & n54234;
  assign n54236 = ~n54229 & ~n54235;
  assign n54237 = pi270 & ~n46154;
  assign n54238 = ~pi805 & n46154;
  assign n54239 = ~pi1091 & ~n54238;
  assign n54240 = ~pi1091 & ~n54237;
  assign n54241 = ~n54238 & n54240;
  assign n54242 = ~n54237 & n54239;
  assign n54243 = ~n54236 & ~n61363;
  assign n54244 = ~pi230 & ~n54243;
  assign n54245 = ~pi230 & ~n54224;
  assign n54246 = ~n54243 & n54245;
  assign n54247 = ~n54224 & n54244;
  assign n54248 = ~pi199 & pi1140;
  assign n54249 = pi200 & ~n54248;
  assign n54250 = ~pi199 & pi1139;
  assign n54251 = pi199 & pi1141;
  assign n54252 = ~pi200 & ~n54251;
  assign n54253 = ~pi200 & ~n54250;
  assign n54254 = ~n54251 & n54253;
  assign n54255 = ~n54250 & n54252;
  assign n54256 = ~n54249 & ~n61365;
  assign n54257 = n44774 & ~n54256;
  assign n54258 = ~pi219 & ~n54227;
  assign n54259 = pi1141 & n36681;
  assign n54260 = pi219 & n54025;
  assign n54261 = pi219 & ~n54025;
  assign n54262 = ~pi219 & n54227;
  assign n54263 = ~n54261 & ~n54262;
  assign n54264 = ~n54258 & ~n61366;
  assign n54265 = ~n44774 & ~n61367;
  assign n54266 = pi230 & ~n54265;
  assign n54267 = pi230 & ~n54257;
  assign n54268 = ~n54265 & n54267;
  assign n54269 = ~n54257 & n54266;
  assign n54270 = ~n61364 & ~n61368;
  assign n54271 = pi274 & ~n46154;
  assign n54272 = ~pi659 & n46154;
  assign n54273 = ~pi1091 & ~n54272;
  assign n54274 = ~pi1091 & ~n54271;
  assign n54275 = ~n54272 & n54274;
  assign n54276 = ~n54271 & n54273;
  assign n54277 = ~n54055 & ~n61369;
  assign n54278 = pi211 & ~n54277;
  assign n54279 = ~n54002 & ~n61369;
  assign n54280 = ~pi211 & ~n54279;
  assign n54281 = ~pi219 & ~n54280;
  assign n54282 = ~pi219 & ~n54278;
  assign n54283 = ~n54280 & n54282;
  assign n54284 = ~n54278 & n54281;
  assign n54285 = pi274 & ~n46143;
  assign n54286 = ~pi659 & n46143;
  assign n54287 = ~pi1091 & ~n54286;
  assign n54288 = ~pi1091 & ~n54285;
  assign n54289 = ~n54286 & n54288;
  assign n54290 = ~n54285 & n54287;
  assign n54291 = pi219 & ~n53953;
  assign n54292 = ~n61371 & n54291;
  assign n54293 = ~n44774 & ~n54292;
  assign n54294 = ~n61370 & n54293;
  assign n54295 = pi200 & ~n54277;
  assign n54296 = ~pi200 & ~n54279;
  assign n54297 = ~pi199 & ~n54296;
  assign n54298 = ~pi199 & ~n54295;
  assign n54299 = ~n54296 & n54298;
  assign n54300 = ~n54295 & n54297;
  assign n54301 = ~pi200 & n53938;
  assign n54302 = pi199 & ~n54301;
  assign n54303 = ~n61371 & n54302;
  assign n54304 = n44774 & ~n54303;
  assign n54305 = ~n61372 & n54304;
  assign n54306 = ~pi230 & ~n54305;
  assign n54307 = ~n54294 & n54306;
  assign n54308 = ~pi219 & ~n49358;
  assign n54309 = ~n49798 & n54308;
  assign n54310 = ~n51663 & ~n54309;
  assign n54311 = ~n47414 & ~n51628;
  assign n54312 = ~n54309 & ~n54311;
  assign n54313 = ~n49368 & n51781;
  assign n54314 = n52346 & ~n54313;
  assign n54315 = ~n54312 & ~n54314;
  assign n54316 = n58992 & ~n54315;
  assign n54317 = pi230 & ~n54316;
  assign n54318 = ~n54310 & n54317;
  assign po431 = ~n54307 & ~n54318;
  assign n54320 = ~pi276 & ~n46144;
  assign n54321 = n46146 & ~n54320;
  assign n54322 = ~n53865 & n54176;
  assign n54323 = pi199 & ~n53870;
  assign n54324 = n44774 & n54323;
  assign n54325 = ~n54322 & ~n54324;
  assign n54326 = ~n54321 & ~n54325;
  assign n54327 = ~pi276 & ~n46155;
  assign n54328 = n53893 & ~n54327;
  assign n54329 = ~n49349 & ~n51640;
  assign n54330 = pi1091 & ~n54329;
  assign n54331 = n49295 & ~n54330;
  assign n54332 = pi1145 & n46364;
  assign n54333 = ~n54056 & ~n54332;
  assign n54334 = n49296 & n54333;
  assign n54335 = ~n54331 & ~n54334;
  assign n54336 = ~n54328 & ~n54335;
  assign n54337 = ~pi230 & ~n54336;
  assign n54338 = ~pi230 & ~n54326;
  assign n54339 = ~n54336 & n54338;
  assign n54340 = ~n54326 & n54337;
  assign n54341 = pi1146 & n36681;
  assign n54342 = pi219 & n51639;
  assign n54343 = ~pi219 & ~n54329;
  assign n54344 = ~n61374 & ~n54343;
  assign n54345 = ~n44774 & n54344;
  assign n54346 = ~n49366 & n52567;
  assign n54347 = ~n51783 & ~n54346;
  assign n54348 = n44774 & ~n54347;
  assign n54349 = pi230 & ~n54348;
  assign n54350 = pi230 & ~n54345;
  assign n54351 = ~n54348 & n54350;
  assign n54352 = ~n54345 & n54349;
  assign n54353 = ~n61373 & ~n61375;
  assign n54354 = pi277 & ~n46154;
  assign n54355 = ~pi820 & n46154;
  assign n54356 = ~pi1091 & ~n54355;
  assign n54357 = ~pi1091 & ~n54354;
  assign n54358 = ~n54355 & n54357;
  assign n54359 = ~n54354 & n54356;
  assign n54360 = ~n54230 & ~n61376;
  assign n54361 = ~pi200 & ~n54360;
  assign n54362 = ~n53986 & ~n61376;
  assign n54363 = pi200 & ~n54362;
  assign n54364 = ~pi199 & ~n54363;
  assign n54365 = ~pi199 & ~n54361;
  assign n54366 = ~n54363 & n54365;
  assign n54367 = ~n54361 & n54364;
  assign n54368 = pi277 & ~n46143;
  assign n54369 = ~pi820 & n46143;
  assign n54370 = ~pi1091 & ~n54369;
  assign n54371 = ~pi1091 & ~n54368;
  assign n54372 = ~n54369 & n54371;
  assign n54373 = ~n54368 & n54370;
  assign n54374 = ~pi200 & n53989;
  assign n54375 = pi199 & ~n54374;
  assign n54376 = ~n61378 & n54375;
  assign n54377 = n44774 & ~n54376;
  assign n54378 = ~n61377 & n54377;
  assign n54379 = ~pi211 & ~n54360;
  assign n54380 = pi211 & ~n54362;
  assign n54381 = ~pi219 & ~n54380;
  assign n54382 = ~pi219 & ~n54379;
  assign n54383 = ~n54380 & n54382;
  assign n54384 = ~n54379 & n54381;
  assign n54385 = ~n49391 & ~n54014;
  assign n54386 = ~n61378 & ~n54385;
  assign n54387 = ~n44774 & ~n54386;
  assign n54388 = ~n61379 & n54387;
  assign n54389 = ~n54378 & ~n54388;
  assign n54390 = ~pi230 & ~n54389;
  assign n54391 = n49365 & ~n54248;
  assign n54392 = pi200 & ~n54021;
  assign n54393 = ~n54391 & ~n54392;
  assign n54394 = n44774 & ~n54393;
  assign n54395 = pi211 & pi1141;
  assign n54396 = ~pi211 & pi1140;
  assign n54397 = ~pi219 & ~n54396;
  assign n54398 = ~pi219 & ~n54395;
  assign n54399 = ~n54396 & n54398;
  assign n54400 = ~n54395 & n54397;
  assign n54401 = ~n49391 & ~n61380;
  assign n54402 = ~n44774 & ~n54401;
  assign n54403 = pi230 & ~n54402;
  assign n54404 = pi230 & ~n54394;
  assign n54405 = ~n54402 & n54404;
  assign n54406 = ~n54394 & n54403;
  assign n54407 = ~n54390 & ~n61381;
  assign n54408 = ~pi976 & n46143;
  assign n54409 = ~pi278 & ~n46143;
  assign n54410 = ~pi1091 & ~n54409;
  assign n54411 = ~pi1091 & ~n54408;
  assign n54412 = ~n54409 & n54411;
  assign n54413 = ~n54408 & n54410;
  assign n54414 = pi199 & ~n61382;
  assign n54415 = pi1091 & ~pi1132;
  assign n54416 = pi278 & ~n46154;
  assign n54417 = pi976 & n46154;
  assign n54418 = ~pi1091 & ~n54417;
  assign n54419 = ~pi1091 & ~n54416;
  assign n54420 = ~n54417 & n54419;
  assign n54421 = ~n54416 & n54418;
  assign n54422 = ~n54415 & ~n61383;
  assign n54423 = ~pi199 & ~n54422;
  assign n54424 = ~n54414 & ~n54423;
  assign n54425 = ~pi200 & ~n54424;
  assign n54426 = pi1091 & ~pi1133;
  assign n54427 = ~n61383 & ~n54426;
  assign n54428 = ~pi199 & ~n54427;
  assign n54429 = ~n54414 & ~n54428;
  assign n54430 = pi200 & ~n54429;
  assign n54431 = ~pi299 & ~n54430;
  assign n54432 = ~n54425 & n54431;
  assign n54433 = pi219 & ~n61382;
  assign n54434 = ~pi211 & pi1132;
  assign n54435 = pi211 & pi1133;
  assign n54436 = pi211 & ~pi1133;
  assign n54437 = ~pi211 & ~pi1132;
  assign n54438 = ~n54436 & ~n54437;
  assign n54439 = ~n54434 & ~n54435;
  assign n54440 = pi1091 & ~n61384;
  assign n54441 = ~n61383 & ~n54440;
  assign n54442 = ~pi219 & ~n54441;
  assign n54443 = ~n54433 & ~n54442;
  assign n54444 = pi299 & n54443;
  assign n54445 = ~n54432 & ~n54444;
  assign n54446 = n58992 & ~n54445;
  assign n54447 = ~n58992 & n54443;
  assign n54448 = ~pi230 & ~n54447;
  assign n54449 = ~n54446 & n54448;
  assign n54450 = ~pi199 & pi1132;
  assign n54451 = ~pi200 & ~n54450;
  assign n54452 = ~pi199 & pi1133;
  assign n54453 = pi200 & ~n54452;
  assign n54454 = ~pi299 & ~n54453;
  assign n54455 = ~n54451 & n54454;
  assign n54456 = n47414 & n61384;
  assign n54457 = ~n54455 & ~n54456;
  assign n54458 = n58992 & ~n54457;
  assign n54459 = n47437 & n61384;
  assign n54460 = pi230 & ~n54459;
  assign n54461 = ~n54458 & n54460;
  assign n54462 = ~n54449 & ~n54461;
  assign n54463 = ~pi1134 & ~n54462;
  assign n54464 = ~pi219 & ~n61384;
  assign n54465 = ~n51610 & ~n54464;
  assign n54466 = n36719 & ~n54450;
  assign n54467 = n54454 & ~n54466;
  assign n54468 = ~n47135 & ~n54456;
  assign n54469 = ~n54467 & n54468;
  assign n54470 = n58992 & ~n54469;
  assign n54471 = pi230 & ~n54470;
  assign n54472 = ~n54465 & n54471;
  assign n54473 = ~n46354 & n54425;
  assign n54474 = n54431 & ~n54473;
  assign n54475 = n45448 & n46717;
  assign n54476 = ~n54444 & ~n54475;
  assign n54477 = ~n54474 & n54476;
  assign n54478 = n58992 & ~n54477;
  assign n54479 = ~n53905 & n54448;
  assign n54480 = ~n54478 & n54479;
  assign n54481 = ~n54472 & ~n54480;
  assign n54482 = pi1134 & ~n54481;
  assign po435 = ~n54463 & ~n54482;
  assign n54484 = ~pi958 & n46143;
  assign n54485 = ~pi279 & ~n46143;
  assign n54486 = ~pi1091 & ~n54485;
  assign n54487 = ~pi1091 & ~n54484;
  assign n54488 = ~n54485 & n54487;
  assign n54489 = ~n54484 & n54486;
  assign n54490 = pi1135 & n54179;
  assign n54491 = ~n61385 & ~n54490;
  assign n54492 = pi199 & ~n54491;
  assign n54493 = pi279 & ~n46154;
  assign n54494 = pi958 & n46154;
  assign n54495 = ~pi1091 & ~n54494;
  assign n54496 = ~pi1091 & ~n54493;
  assign n54497 = ~n54494 & n54496;
  assign n54498 = ~n54493 & n54495;
  assign n54499 = ~pi1133 & n54179;
  assign n54500 = ~pi199 & ~n54499;
  assign n54501 = ~n61386 & n54500;
  assign n54502 = ~n54492 & ~n54501;
  assign n54503 = n44774 & ~n54502;
  assign n54504 = ~n46364 & n54503;
  assign n54505 = ~n46707 & ~n54426;
  assign n54506 = ~n61386 & n54505;
  assign n54507 = ~pi219 & ~n54506;
  assign n54508 = pi1135 & n46717;
  assign n54509 = pi219 & ~n54508;
  assign n54510 = ~n61385 & n54509;
  assign n54511 = ~n44774 & ~n54510;
  assign n54512 = ~n54507 & n54511;
  assign n54513 = ~pi230 & ~n54512;
  assign n54514 = ~n54504 & n54513;
  assign n54515 = pi199 & pi1135;
  assign n54516 = ~n54452 & ~n54515;
  assign n54517 = n46389 & ~n54516;
  assign n54518 = pi1135 & n36681;
  assign n54519 = ~pi211 & ~pi1133;
  assign n54520 = ~pi219 & ~n54519;
  assign n54521 = ~pi211 & n54520;
  assign n54522 = ~n54518 & ~n54521;
  assign n54523 = pi299 & ~n54522;
  assign n54524 = ~n54517 & ~n54523;
  assign n54525 = n58992 & ~n54524;
  assign n54526 = ~n58992 & ~n54522;
  assign n54527 = pi230 & ~n54526;
  assign n54528 = ~n54525 & n54527;
  assign n54529 = ~n54514 & ~n54528;
  assign n54530 = ~pi1134 & ~n54529;
  assign n54531 = ~pi1133 & n36719;
  assign n54532 = ~pi200 & pi1135;
  assign n54533 = pi199 & ~n54532;
  assign n54534 = ~n54531 & ~n54533;
  assign n54535 = n44774 & ~n54534;
  assign n54536 = ~n54518 & ~n54520;
  assign n54537 = ~n44774 & n54536;
  assign n54538 = ~n54535 & ~n54537;
  assign n54539 = pi230 & ~n54538;
  assign n54540 = pi1091 & ~n54519;
  assign n54541 = n49295 & n54540;
  assign n54542 = ~n54503 & ~n54541;
  assign n54543 = n54513 & n54542;
  assign n54544 = ~n54539 & ~n54543;
  assign n54545 = pi1134 & ~n54544;
  assign po436 = ~n54530 & ~n54545;
  assign n54547 = pi1137 & n54179;
  assign n54548 = pi280 & ~n46143;
  assign n54549 = ~pi914 & n46143;
  assign n54550 = ~pi1091 & ~n54549;
  assign n54551 = ~pi1091 & ~n54548;
  assign n54552 = ~n54549 & n54551;
  assign n54553 = ~n54548 & n54550;
  assign n54554 = ~n54547 & ~n61387;
  assign n54555 = pi199 & ~n54554;
  assign n54556 = pi914 & n46154;
  assign n54557 = ~pi280 & ~n46154;
  assign n54558 = ~pi1091 & ~n54557;
  assign n54559 = ~pi1091 & ~n54556;
  assign n54560 = ~n54557 & n54559;
  assign n54561 = ~n54556 & n54558;
  assign n54562 = pi200 & pi1136;
  assign n54563 = pi1091 & ~n54532;
  assign n54564 = ~n54562 & n54563;
  assign n54565 = ~pi199 & ~n54564;
  assign n54566 = ~n61388 & n54565;
  assign n54567 = ~n54555 & ~n54566;
  assign n54568 = n44774 & ~n54567;
  assign n54569 = ~pi211 & pi1135;
  assign n54570 = pi211 & pi1136;
  assign n54571 = ~n54569 & ~n54570;
  assign n54572 = pi1091 & n54571;
  assign n54573 = ~n61388 & ~n54572;
  assign n54574 = ~pi219 & ~n54573;
  assign n54575 = ~pi211 & pi1137;
  assign n54576 = pi219 & ~n54575;
  assign n54577 = ~n54014 & ~n54576;
  assign n54578 = ~n61387 & ~n54577;
  assign n54579 = ~n44774 & ~n54578;
  assign n54580 = ~n54574 & n54579;
  assign n54581 = ~n54574 & ~n54578;
  assign n54582 = ~n44774 & ~n54581;
  assign n54583 = n44774 & ~n54566;
  assign n54584 = n44774 & ~n54555;
  assign n54585 = ~n54566 & n54584;
  assign n54586 = ~n54555 & n54583;
  assign n54587 = ~n54582 & ~n61389;
  assign n54588 = ~n54568 & ~n54580;
  assign n54589 = ~pi230 & n61390;
  assign n54590 = pi200 & ~n54195;
  assign n54591 = pi199 & pi1137;
  assign n54592 = ~pi200 & ~n54091;
  assign n54593 = ~n54591 & n54592;
  assign n54594 = ~n54590 & ~n54593;
  assign n54595 = n44774 & ~n54594;
  assign n54596 = ~pi219 & n54571;
  assign n54597 = ~n54576 & ~n54596;
  assign n54598 = ~n44774 & ~n54597;
  assign n54599 = pi230 & ~n54598;
  assign n54600 = ~n54595 & n54599;
  assign n54601 = ~pi230 & ~n61390;
  assign n54602 = n44774 & n54594;
  assign n54603 = ~n44774 & n54597;
  assign n54604 = pi230 & ~n54603;
  assign n54605 = pi230 & ~n54602;
  assign n54606 = ~n54603 & n54605;
  assign n54607 = ~n54602 & n54604;
  assign n54608 = ~n54601 & ~n61391;
  assign n54609 = ~n54589 & ~n54600;
  assign n54610 = pi211 & pi1138;
  assign n54611 = ~n54575 & ~n54610;
  assign n54612 = pi1091 & ~n54611;
  assign n54613 = n49295 & ~n54612;
  assign n54614 = pi1138 & n46364;
  assign n54615 = ~n54547 & ~n54614;
  assign n54616 = n49296 & n54615;
  assign n54617 = ~n54613 & ~n54616;
  assign n54618 = pi281 & ~n46154;
  assign n54619 = ~pi830 & n46154;
  assign n54620 = ~pi1091 & ~n54619;
  assign n54621 = ~pi1091 & ~n54618;
  assign n54622 = ~n54619 & n54621;
  assign n54623 = ~n54618 & n54620;
  assign n54624 = ~n54617 & ~n61393;
  assign n54625 = pi1139 & n46717;
  assign n54626 = n54176 & ~n54625;
  assign n54627 = pi199 & ~n54233;
  assign n54628 = n44774 & n54627;
  assign n54629 = ~n54626 & ~n54628;
  assign n54630 = pi281 & ~n46143;
  assign n54631 = ~pi830 & n46143;
  assign n54632 = ~pi1091 & ~n54631;
  assign n54633 = ~pi1091 & ~n54630;
  assign n54634 = ~n54631 & n54633;
  assign n54635 = ~n54630 & n54632;
  assign n54636 = ~n54629 & ~n61394;
  assign n54637 = ~n54624 & ~n54636;
  assign n54638 = ~pi230 & ~n54637;
  assign n54639 = ~pi199 & pi1138;
  assign n54640 = pi200 & ~n54639;
  assign n54641 = pi199 & pi1139;
  assign n54642 = ~pi200 & ~n54193;
  assign n54643 = ~n54641 & n54642;
  assign n54644 = ~n54640 & ~n54643;
  assign n54645 = n44774 & ~n54644;
  assign n54646 = pi219 & n54225;
  assign n54647 = ~pi219 & ~n54611;
  assign n54648 = ~n54646 & ~n54647;
  assign n54649 = ~n44774 & n54648;
  assign n54650 = ~n54645 & ~n54649;
  assign n54651 = pi230 & ~n54650;
  assign po438 = ~n54638 & ~n54651;
  assign n54653 = pi211 & pi1139;
  assign n54654 = ~n54204 & ~n54653;
  assign n54655 = pi1091 & ~n54654;
  assign n54656 = n49295 & ~n54655;
  assign n54657 = pi1139 & n46364;
  assign n54658 = ~n54180 & ~n54657;
  assign n54659 = n49296 & n54658;
  assign n54660 = ~n54656 & ~n54659;
  assign n54661 = pi282 & ~n46154;
  assign n54662 = ~pi836 & n46154;
  assign n54663 = ~pi1091 & ~n54662;
  assign n54664 = ~pi1091 & ~n54661;
  assign n54665 = ~n54662 & n54664;
  assign n54666 = ~n54661 & n54663;
  assign n54667 = ~n54660 & ~n61395;
  assign n54668 = pi1140 & n46717;
  assign n54669 = n54176 & ~n54668;
  assign n54670 = ~pi200 & n54230;
  assign n54671 = pi199 & ~n54670;
  assign n54672 = n44774 & n54671;
  assign n54673 = ~n54669 & ~n54672;
  assign n54674 = pi282 & ~n46143;
  assign n54675 = ~pi836 & n46143;
  assign n54676 = ~pi1091 & ~n54675;
  assign n54677 = ~pi1091 & ~n54674;
  assign n54678 = ~n54675 & n54677;
  assign n54679 = ~n54674 & n54676;
  assign n54680 = ~n54673 & ~n61396;
  assign n54681 = ~n54667 & ~n54680;
  assign n54682 = ~pi230 & ~n54681;
  assign n54683 = pi200 & ~n54250;
  assign n54684 = pi199 & pi1140;
  assign n54685 = ~pi200 & ~n54639;
  assign n54686 = ~n54684 & n54685;
  assign n54687 = ~n54683 & ~n54686;
  assign n54688 = n44774 & ~n54687;
  assign n54689 = pi219 & n54396;
  assign n54690 = ~pi219 & ~n54654;
  assign n54691 = ~n54689 & ~n54690;
  assign n54692 = ~n44774 & n54691;
  assign n54693 = ~n54688 & ~n54692;
  assign n54694 = pi230 & ~n54693;
  assign po439 = ~n54682 & ~n54694;
  assign n54696 = n58992 & n60068;
  assign n54697 = n60068 & ~n36439;
  assign n54698 = n58992 & n54697;
  assign n54699 = ~n36439 & n60563;
  assign n54700 = ~pi330 & n61397;
  assign n54701 = pi336 & ~n54700;
  assign n54702 = pi1070 & n54700;
  assign n54703 = ~n54701 & ~n54702;
  assign n54704 = pi337 & ~n54700;
  assign n54705 = pi1044 & n54700;
  assign n54706 = ~n54704 & ~n54705;
  assign n54707 = ~pi340 & n54697;
  assign n54708 = n58992 & n54707;
  assign n54709 = ~pi340 & n61397;
  assign n54710 = pi342 & ~n61398;
  assign n54711 = pi1049 & n61398;
  assign n54712 = ~n54710 & ~n54711;
  assign n54713 = pi343 & ~n61398;
  assign n54714 = pi1062 & n61398;
  assign n54715 = ~n54713 & ~n54714;
  assign n54716 = pi345 & ~n61398;
  assign n54717 = pi1039 & n61398;
  assign n54718 = ~n54716 & ~n54717;
  assign n54719 = pi346 & ~n61398;
  assign n54720 = pi1067 & n61398;
  assign n54721 = ~n54719 & ~n54720;
  assign n54722 = pi347 & ~n61398;
  assign n54723 = pi1055 & n61398;
  assign n54724 = ~n54722 & ~n54723;
  assign n54725 = pi348 & ~n61398;
  assign n54726 = pi1087 & n61398;
  assign n54727 = ~n54725 & ~n54726;
  assign n54728 = pi350 & ~n61398;
  assign n54729 = pi1035 & n61398;
  assign n54730 = ~n54728 & ~n54729;
  assign n54731 = pi351 & ~n61398;
  assign n54732 = pi1079 & n61398;
  assign n54733 = ~n54731 & ~n54732;
  assign n54734 = pi354 & ~n61398;
  assign n54735 = pi1045 & n61398;
  assign n54736 = ~n54734 & ~n54735;
  assign n54737 = pi355 & ~n61398;
  assign n54738 = pi1084 & n61398;
  assign n54739 = ~n54737 & ~n54738;
  assign n54740 = pi356 & ~n61398;
  assign n54741 = pi1081 & n61398;
  assign n54742 = ~n54740 & ~n54741;
  assign n54743 = pi357 & ~n61398;
  assign n54744 = pi1076 & n61398;
  assign n54745 = ~n54743 & ~n54744;
  assign n54746 = pi358 & ~n61398;
  assign n54747 = pi1071 & n61398;
  assign n54748 = ~n54746 & ~n54747;
  assign n54749 = pi359 & ~n61398;
  assign n54750 = pi1068 & n61398;
  assign n54751 = ~n54749 & ~n54750;
  assign n54752 = pi360 & ~n61398;
  assign n54753 = pi1042 & n61398;
  assign n54754 = ~n54752 & ~n54753;
  assign n54755 = pi361 & ~n61398;
  assign n54756 = pi1059 & n61398;
  assign n54757 = ~n54755 & ~n54756;
  assign n54758 = pi362 & ~n61398;
  assign n54759 = pi1070 & n61398;
  assign n54760 = ~n54758 & ~n54759;
  assign n54761 = pi363 & ~n54700;
  assign n54762 = pi1049 & n54700;
  assign n54763 = ~n54761 & ~n54762;
  assign n54764 = pi364 & ~n54700;
  assign n54765 = pi1062 & n54700;
  assign n54766 = ~n54764 & ~n54765;
  assign n54767 = pi367 & ~n54700;
  assign n54768 = pi1039 & n54700;
  assign n54769 = ~n54767 & ~n54768;
  assign n54770 = pi368 & ~n54700;
  assign n54771 = pi1067 & n54700;
  assign n54772 = ~n54770 & ~n54771;
  assign n54773 = pi370 & ~n54700;
  assign n54774 = pi1055 & n54700;
  assign n54775 = ~n54773 & ~n54774;
  assign n54776 = pi373 & ~n54700;
  assign n54777 = pi1087 & n54700;
  assign n54778 = ~n54776 & ~n54777;
  assign n54779 = pi374 & ~n54700;
  assign n54780 = pi1035 & n54700;
  assign n54781 = ~n54779 & ~n54780;
  assign n54782 = pi376 & ~n54700;
  assign n54783 = pi1079 & n54700;
  assign n54784 = ~n54782 & ~n54783;
  assign n54785 = pi379 & ~n54700;
  assign n54786 = pi1045 & n54700;
  assign n54787 = ~n54785 & ~n54786;
  assign n54788 = pi380 & ~n54700;
  assign n54789 = pi1084 & n54700;
  assign n54790 = ~n54788 & ~n54789;
  assign n54791 = pi381 & ~n54700;
  assign n54792 = pi1081 & n54700;
  assign n54793 = ~n54791 & ~n54792;
  assign n54794 = pi382 & ~n54700;
  assign n54795 = pi1076 & n54700;
  assign n54796 = ~n54794 & ~n54795;
  assign n54797 = pi383 & ~n54700;
  assign n54798 = pi1071 & n54700;
  assign n54799 = ~n54797 & ~n54798;
  assign n54800 = pi384 & ~n54700;
  assign n54801 = pi1068 & n54700;
  assign n54802 = ~n54800 & ~n54801;
  assign n54803 = pi385 & ~n54700;
  assign n54804 = pi1042 & n54700;
  assign n54805 = ~n54803 & ~n54804;
  assign n54806 = pi386 & ~n54700;
  assign n54807 = pi1059 & n54700;
  assign n54808 = ~n54806 & ~n54807;
  assign n54809 = pi387 & ~n54700;
  assign n54810 = pi1053 & n54700;
  assign n54811 = ~n54809 & ~n54810;
  assign n54812 = pi388 & ~n54700;
  assign n54813 = pi1037 & n54700;
  assign n54814 = ~n54812 & ~n54813;
  assign n54815 = pi389 & ~n54700;
  assign n54816 = pi1036 & n54700;
  assign n54817 = ~n54815 & ~n54816;
  assign n54818 = ~pi341 & n54697;
  assign n54819 = n58992 & n54818;
  assign n54820 = ~pi341 & n61397;
  assign n54821 = pi390 & ~n61399;
  assign n54822 = pi1049 & n61399;
  assign n54823 = ~n54821 & ~n54822;
  assign n54824 = pi391 & ~n61399;
  assign n54825 = pi1062 & n61399;
  assign n54826 = ~n54824 & ~n54825;
  assign n54827 = pi392 & ~n61399;
  assign n54828 = pi1039 & n61399;
  assign n54829 = ~n54827 & ~n54828;
  assign n54830 = pi393 & ~n61399;
  assign n54831 = pi1067 & n61399;
  assign n54832 = ~n54830 & ~n54831;
  assign n54833 = pi395 & ~n61399;
  assign n54834 = pi1055 & n61399;
  assign n54835 = ~n54833 & ~n54834;
  assign n54836 = pi398 & ~n61399;
  assign n54837 = pi1087 & n61399;
  assign n54838 = ~n54836 & ~n54837;
  assign n54839 = pi400 & ~n61399;
  assign n54840 = pi1035 & n61399;
  assign n54841 = ~n54839 & ~n54840;
  assign n54842 = pi401 & ~n61399;
  assign n54843 = pi1079 & n61399;
  assign n54844 = ~n54842 & ~n54843;
  assign n54845 = pi403 & ~n61399;
  assign n54846 = pi1045 & n61399;
  assign n54847 = ~n54845 & ~n54846;
  assign n54848 = pi404 & ~n61399;
  assign n54849 = pi1084 & n61399;
  assign n54850 = ~n54848 & ~n54849;
  assign n54851 = pi405 & ~n61399;
  assign n54852 = pi1081 & n61399;
  assign n54853 = ~n54851 & ~n54852;
  assign n54854 = pi406 & ~n61399;
  assign n54855 = pi1076 & n61399;
  assign n54856 = ~n54854 & ~n54855;
  assign n54857 = pi407 & ~n61399;
  assign n54858 = pi1071 & n61399;
  assign n54859 = ~n54857 & ~n54858;
  assign n54860 = pi408 & ~n61399;
  assign n54861 = pi1068 & n61399;
  assign n54862 = ~n54860 & ~n54861;
  assign n54863 = pi409 & ~n61399;
  assign n54864 = pi1042 & n61399;
  assign n54865 = ~n54863 & ~n54864;
  assign n54866 = pi410 & ~n61399;
  assign n54867 = pi1059 & n61399;
  assign n54868 = ~n54866 & ~n54867;
  assign n54869 = pi411 & ~n61399;
  assign n54870 = pi1053 & n61399;
  assign n54871 = ~n54869 & ~n54870;
  assign n54872 = pi412 & ~n61399;
  assign n54873 = pi1037 & n61399;
  assign n54874 = ~n54872 & ~n54873;
  assign n54875 = pi413 & ~n61399;
  assign n54876 = pi1036 & n61399;
  assign n54877 = ~n54875 & ~n54876;
  assign n54878 = ~pi331 & n54697;
  assign n54879 = n58992 & n54878;
  assign n54880 = ~pi331 & n61397;
  assign n54881 = pi414 & ~n61400;
  assign n54882 = pi1049 & n61400;
  assign n54883 = ~n54881 & ~n54882;
  assign n54884 = pi415 & ~n61400;
  assign n54885 = pi1062 & n61400;
  assign n54886 = ~n54884 & ~n54885;
  assign n54887 = pi417 & ~n61400;
  assign n54888 = pi1039 & n61400;
  assign n54889 = ~n54887 & ~n54888;
  assign n54890 = pi418 & ~n61400;
  assign n54891 = pi1067 & n61400;
  assign n54892 = ~n54890 & ~n54891;
  assign n54893 = pi420 & ~n61400;
  assign n54894 = pi1055 & n61400;
  assign n54895 = ~n54893 & ~n54894;
  assign n54896 = pi423 & ~n61400;
  assign n54897 = pi1087 & n61400;
  assign n54898 = ~n54896 & ~n54897;
  assign n54899 = pi425 & ~n61400;
  assign n54900 = pi1035 & n61400;
  assign n54901 = ~n54899 & ~n54900;
  assign n54902 = pi426 & ~n61400;
  assign n54903 = pi1079 & n61400;
  assign n54904 = ~n54902 & ~n54903;
  assign n54905 = pi428 & ~n61400;
  assign n54906 = pi1045 & n61400;
  assign n54907 = ~n54905 & ~n54906;
  assign n54908 = pi429 & ~n61400;
  assign n54909 = pi1084 & n61400;
  assign n54910 = ~n54908 & ~n54909;
  assign n54911 = pi430 & ~n61400;
  assign n54912 = pi1076 & n61400;
  assign n54913 = ~n54911 & ~n54912;
  assign n54914 = pi431 & ~n61400;
  assign n54915 = pi1071 & n61400;
  assign n54916 = ~n54914 & ~n54915;
  assign n54917 = pi432 & ~n61400;
  assign n54918 = pi1068 & n61400;
  assign n54919 = ~n54917 & ~n54918;
  assign n54920 = pi433 & ~n61400;
  assign n54921 = pi1042 & n61400;
  assign n54922 = ~n54920 & ~n54921;
  assign n54923 = pi434 & ~n61400;
  assign n54924 = pi1059 & n61400;
  assign n54925 = ~n54923 & ~n54924;
  assign n54926 = pi435 & ~n61400;
  assign n54927 = pi1053 & n61400;
  assign n54928 = ~n54926 & ~n54927;
  assign n54929 = pi436 & ~n61400;
  assign n54930 = pi1037 & n61400;
  assign n54931 = ~n54929 & ~n54930;
  assign n54932 = pi437 & ~n61400;
  assign n54933 = pi1070 & n61400;
  assign n54934 = ~n54932 & ~n54933;
  assign n54935 = pi438 & ~n61400;
  assign n54936 = pi1036 & n61400;
  assign n54937 = ~n54935 & ~n54936;
  assign n54938 = pi441 & ~n61398;
  assign n54939 = pi1044 & n61398;
  assign n54940 = ~n54938 & ~n54939;
  assign n54941 = pi443 & ~n61400;
  assign n54942 = pi1044 & n61400;
  assign n54943 = ~n54941 & ~n54942;
  assign n54944 = pi445 & ~n61400;
  assign n54945 = pi1081 & n61400;
  assign n54946 = ~n54944 & ~n54945;
  assign n54947 = pi450 & ~n61398;
  assign n54948 = pi1036 & n61398;
  assign n54949 = ~n54947 & ~n54948;
  assign n54950 = pi452 & ~n61398;
  assign n54951 = pi1053 & n61398;
  assign n54952 = ~n54950 & ~n54951;
  assign n54953 = pi455 & ~n61398;
  assign n54954 = pi1037 & n61398;
  assign n54955 = ~n54953 & ~n54954;
  assign n54956 = pi456 & ~n61399;
  assign n54957 = pi1044 & n61399;
  assign n54958 = ~n54956 & ~n54957;
  assign n54959 = pi463 & ~n61399;
  assign n54960 = pi1070 & n61399;
  assign n54961 = ~n54959 & ~n54960;
  assign n54962 = n60165 & n60563;
  assign n54963 = n2621 & n60563;
  assign n54964 = n59138 & n54963;
  assign n54965 = ~n45456 & n54964;
  assign n54966 = ~n45456 & n54962;
  assign n54967 = ~n45454 & n61401;
  assign n54968 = ~pi954 & ~n54967;
  assign n54969 = pi313 & pi954;
  assign po470 = ~n54968 & ~n54969;
  assign n54971 = pi228 & pi231;
  assign n54972 = ~pi228 & n45485;
  assign n54973 = ~n54971 & ~n54972;
  assign n54974 = ~pi100 & ~n54973;
  assign n54975 = ~n31587 & ~n54971;
  assign n54976 = pi100 & ~n54975;
  assign n54977 = ~pi87 & ~n54976;
  assign n54978 = ~n54974 & n54977;
  assign n54979 = pi87 & ~n54971;
  assign n54980 = ~n32934 & n54979;
  assign n54981 = ~pi75 & ~n54980;
  assign n54982 = ~n54978 & n54981;
  assign n54983 = ~n60247 & ~n54971;
  assign n54984 = pi75 & ~n54983;
  assign n54985 = ~pi92 & ~n54984;
  assign n54986 = ~n54982 & n54985;
  assign n54987 = pi92 & ~n54971;
  assign n54988 = ~n60282 & n54987;
  assign n54989 = ~n54986 & ~n54988;
  assign n54990 = ~pi54 & ~n54989;
  assign n54991 = pi54 & ~n54971;
  assign n54992 = ~pi74 & ~n54991;
  assign n54993 = ~n54990 & n54992;
  assign n54994 = ~n60249 & ~n54971;
  assign n54995 = ~n31593 & ~n54971;
  assign n54996 = pi74 & ~n54995;
  assign n54997 = ~n54983 & n54996;
  assign n54998 = pi74 & ~n54994;
  assign n54999 = ~pi55 & ~n61402;
  assign n55000 = ~n54993 & n54999;
  assign n55001 = pi55 & ~n54971;
  assign n55002 = ~pi56 & ~n55001;
  assign n55003 = ~n55000 & n55002;
  assign n55004 = ~n60829 & ~n54971;
  assign n55005 = pi56 & ~n55004;
  assign n55006 = ~pi62 & ~n55005;
  assign n55007 = ~n55003 & n55006;
  assign n55008 = pi62 & ~n54971;
  assign n55009 = ~n60828 & n55008;
  assign n55010 = ~n55007 & ~n55009;
  assign n55011 = n4438 & ~n55010;
  assign n55012 = ~n4438 & ~n54971;
  assign po383 = ~n55011 & ~n55012;
  assign n55014 = n4437 & n60068;
  assign n55015 = n58826 & n55014;
  assign n55016 = pi57 & ~pi59;
  assign n55017 = n55015 & n55016;
  assign n55018 = ~pi312 & n55017;
  assign n55019 = ~pi300 & pi301;
  assign n55020 = ~pi55 & n55019;
  assign n55021 = ~pi300 & n55018;
  assign n55022 = ~pi55 & pi301;
  assign n55023 = n55021 & n55022;
  assign n55024 = n55018 & n55020;
  assign n55025 = ~pi55 & ~pi311;
  assign n55026 = ~n61403 & ~n55025;
  assign n55027 = ~pi311 & n61403;
  assign n55028 = pi311 & ~n61403;
  assign n55029 = ~pi55 & ~n61403;
  assign n55030 = ~pi311 & ~n55029;
  assign n55031 = ~n55028 & ~n55030;
  assign n55032 = ~n55026 & ~n55027;
  assign n55033 = ~pi55 & ~n55021;
  assign n55034 = ~pi301 & n55033;
  assign n55035 = ~n61403 & ~n55034;
  assign n55036 = n6426 & n45613;
  assign n55037 = ~pi924 & n40707;
  assign n55038 = ~n40706 & ~n55037;
  assign n55039 = n55036 & ~n55038;
  assign n55040 = ~pi57 & ~n55039;
  assign n55041 = n4440 & n60865;
  assign n55042 = pi57 & ~n55041;
  assign n55043 = ~pi59 & ~n55042;
  assign n55044 = ~pi59 & ~n55040;
  assign n55045 = ~n55042 & n55044;
  assign n55046 = ~n55040 & n55043;
  assign n55047 = pi924 & n40707;
  assign n55048 = n55036 & n55047;
  assign n55049 = ~pi59 & ~n55048;
  assign n55050 = pi59 & ~n55041;
  assign n55051 = ~pi57 & ~n55050;
  assign n55052 = ~pi57 & ~n55049;
  assign n55053 = ~n55050 & n55052;
  assign n55054 = ~n55049 & n55051;
  assign n55055 = pi300 & ~n55018;
  assign n55056 = n55033 & ~n55055;
  assign n55057 = n58797 & n31449;
  assign n55058 = n2547 & n31450;
  assign n55059 = n58786 & n55057;
  assign n55060 = pi999 & n61407;
  assign n55061 = ~pi24 & n45584;
  assign n55062 = ~n55060 & ~n55061;
  assign n55063 = n54964 & ~n55062;
  assign n55064 = n54962 & ~n55062;
  assign n55065 = pi312 & ~n55017;
  assign n55066 = ~n55018 & ~n55065;
  assign po469 = ~pi55 & ~n55066;
  assign n55068 = ~pi999 & n54964;
  assign n55069 = ~pi999 & n54962;
  assign po265 = n61407 & n61409;
  assign n55071 = pi481 & ~n44783;
  assign n55072 = pi248 & n44783;
  assign n55073 = ~n55071 & ~n55072;
  assign n55074 = pi482 & ~n44799;
  assign n55075 = pi249 & n44799;
  assign n55076 = ~n55074 & ~n55075;
  assign n55077 = pi483 & ~n44928;
  assign n55078 = pi242 & n44928;
  assign n55079 = ~n55077 & ~n55078;
  assign n55080 = pi484 & ~n44928;
  assign n55081 = pi249 & n44928;
  assign n55082 = ~n55080 & ~n55081;
  assign n55083 = pi485 & ~n44935;
  assign n55084 = pi234 & n44935;
  assign n55085 = ~n55083 & ~n55084;
  assign n55086 = pi486 & ~n44935;
  assign n55087 = pi244 & n44935;
  assign n55088 = ~n55086 & ~n55087;
  assign n55089 = pi487 & ~n44783;
  assign n55090 = pi246 & n44783;
  assign n55091 = ~n55089 & ~n55090;
  assign n55092 = pi488 & ~n44783;
  assign n55093 = ~pi239 & n44783;
  assign po645 = ~n55092 & ~n55093;
  assign n55095 = pi489 & ~n44935;
  assign n55096 = pi242 & n44935;
  assign n55097 = ~n55095 & ~n55096;
  assign n55098 = pi490 & ~n44928;
  assign n55099 = pi241 & n44928;
  assign n55100 = ~n55098 & ~n55099;
  assign n55101 = pi491 & ~n44928;
  assign n55102 = pi238 & n44928;
  assign n55103 = ~n55101 & ~n55102;
  assign n55104 = pi492 & ~n44928;
  assign n55105 = pi240 & n44928;
  assign n55106 = ~n55104 & ~n55105;
  assign n55107 = pi493 & ~n44928;
  assign n55108 = pi244 & n44928;
  assign n55109 = ~n55107 & ~n55108;
  assign n55110 = pi494 & ~n44928;
  assign n55111 = ~pi239 & n44928;
  assign po651 = ~n55110 & ~n55111;
  assign n55113 = pi495 & ~n44928;
  assign n55114 = pi235 & n44928;
  assign n55115 = ~n55113 & ~n55114;
  assign n55116 = pi496 & ~n44920;
  assign n55117 = pi249 & n44920;
  assign n55118 = ~n55116 & ~n55117;
  assign n55119 = pi497 & ~n44920;
  assign n55120 = ~pi239 & n44920;
  assign po654 = ~n55119 & ~n55120;
  assign n55122 = pi498 & ~n44799;
  assign n55123 = pi238 & n44799;
  assign n55124 = ~n55122 & ~n55123;
  assign n55125 = pi499 & ~n44920;
  assign n55126 = pi246 & n44920;
  assign n55127 = ~n55125 & ~n55126;
  assign n55128 = pi500 & ~n44920;
  assign n55129 = pi241 & n44920;
  assign n55130 = ~n55128 & ~n55129;
  assign n55131 = pi501 & ~n44920;
  assign n55132 = pi248 & n44920;
  assign n55133 = ~n55131 & ~n55132;
  assign n55134 = pi502 & ~n44920;
  assign n55135 = pi247 & n44920;
  assign n55136 = ~n55134 & ~n55135;
  assign n55137 = pi503 & ~n44920;
  assign n55138 = pi245 & n44920;
  assign n55139 = ~n55137 & ~n55138;
  assign n55140 = pi504 & ~n44913;
  assign n55141 = pi242 & n44913;
  assign n55142 = ~n55140 & ~n55141;
  assign n55143 = pi505 & ~n44920;
  assign n55144 = pi234 & n44912;
  assign n55145 = n44786 & n55144;
  assign n55146 = ~pi234 & n45852;
  assign n55147 = n44920 & n55146;
  assign n55148 = pi505 & ~n55147;
  assign n55149 = ~pi505 & n44786;
  assign n55150 = n55144 & n55149;
  assign n55151 = ~n55148 & ~n55150;
  assign n55152 = ~n55143 & ~n55145;
  assign n55153 = pi506 & ~n44913;
  assign n55154 = pi241 & n44913;
  assign n55155 = ~n55153 & ~n55154;
  assign n55156 = pi507 & ~n44913;
  assign n55157 = pi238 & n44913;
  assign n55158 = ~n55156 & ~n55157;
  assign n55159 = pi508 & ~n44913;
  assign n55160 = pi247 & n44913;
  assign n55161 = ~n55159 & ~n55160;
  assign n55162 = pi509 & ~n44913;
  assign n55163 = pi245 & n44913;
  assign n55164 = ~n55162 & ~n55163;
  assign n55165 = pi510 & ~n44783;
  assign n55166 = pi242 & n44783;
  assign n55167 = ~n55165 & ~n55166;
  assign n55168 = ~pi234 & n45855;
  assign n55169 = n44783 & ~n55168;
  assign n55170 = pi511 & ~n44783;
  assign n55171 = ~n55169 & ~n55170;
  assign n55172 = pi512 & ~n44783;
  assign n55173 = pi235 & n44783;
  assign n55174 = ~n55172 & ~n55173;
  assign n55175 = pi513 & ~n44783;
  assign n55176 = pi244 & n44783;
  assign n55177 = ~n55175 & ~n55176;
  assign n55178 = pi514 & ~n44783;
  assign n55179 = pi245 & n44783;
  assign n55180 = ~n55178 & ~n55179;
  assign n55181 = pi515 & ~n44783;
  assign n55182 = pi240 & n44783;
  assign n55183 = ~n55181 & ~n55182;
  assign n55184 = pi516 & ~n44783;
  assign n55185 = pi247 & n44783;
  assign n55186 = ~n55184 & ~n55185;
  assign n55187 = pi517 & ~n44783;
  assign n55188 = pi238 & n44783;
  assign n55189 = ~n55187 & ~n55188;
  assign n55190 = pi518 & ~n44791;
  assign n55191 = pi234 & n60820;
  assign n55192 = n44786 & n55191;
  assign n55193 = n44791 & n55168;
  assign n55194 = pi518 & ~n55193;
  assign n55195 = ~pi518 & n44786;
  assign n55196 = n55191 & n55195;
  assign n55197 = ~n55194 & ~n55196;
  assign n55198 = ~n55190 & ~n55192;
  assign n55199 = pi519 & ~n44791;
  assign n55200 = ~pi239 & n44791;
  assign po676 = ~n55199 & ~n55200;
  assign n55202 = pi520 & ~n44791;
  assign n55203 = pi246 & n44791;
  assign n55204 = ~n55202 & ~n55203;
  assign n55205 = pi521 & ~n44791;
  assign n55206 = pi248 & n44791;
  assign n55207 = ~n55205 & ~n55206;
  assign n55208 = pi522 & ~n44791;
  assign n55209 = pi238 & n44791;
  assign n55210 = ~n55208 & ~n55209;
  assign n55211 = pi523 & ~n44942;
  assign n55212 = n44923 & n55191;
  assign n55213 = n44942 & n55168;
  assign n55214 = pi523 & ~n55213;
  assign n55215 = ~pi523 & n44923;
  assign n55216 = n55191 & n55215;
  assign n55217 = ~n55214 & ~n55216;
  assign n55218 = ~n55211 & ~n55212;
  assign n55219 = pi524 & ~n44942;
  assign n55220 = ~pi239 & n44942;
  assign po681 = ~n55219 & ~n55220;
  assign n55222 = pi525 & ~n44942;
  assign n55223 = pi245 & n44942;
  assign n55224 = ~n55222 & ~n55223;
  assign n55225 = pi526 & ~n44942;
  assign n55226 = pi246 & n44942;
  assign n55227 = ~n55225 & ~n55226;
  assign n55228 = pi527 & ~n44942;
  assign n55229 = pi247 & n44942;
  assign n55230 = ~n55228 & ~n55229;
  assign n55231 = pi528 & ~n44942;
  assign n55232 = pi249 & n44942;
  assign n55233 = ~n55231 & ~n55232;
  assign n55234 = pi529 & ~n44942;
  assign n55235 = pi238 & n44942;
  assign n55236 = ~n55234 & ~n55235;
  assign n55237 = pi530 & ~n44942;
  assign n55238 = pi240 & n44942;
  assign n55239 = ~n55237 & ~n55238;
  assign n55240 = pi531 & ~n44799;
  assign n55241 = pi235 & n44799;
  assign n55242 = ~n55240 & ~n55241;
  assign n55243 = pi532 & ~n44799;
  assign n55244 = pi247 & n44799;
  assign n55245 = ~n55243 & ~n55244;
  assign n55246 = pi533 & ~n44913;
  assign n55247 = pi235 & n44913;
  assign n55248 = ~n55246 & ~n55247;
  assign n55249 = ~pi123 & pi228;
  assign n55250 = ~pi228 & pi1093;
  assign n55251 = ~pi228 & ~pi1093;
  assign n55252 = pi123 & pi228;
  assign n55253 = ~n55251 & ~n55252;
  assign n55254 = ~n55249 & ~n55250;
  assign n55255 = pi199 & n61413;
  assign n55256 = ~pi262 & ~pi1093;
  assign n55257 = ~n45954 & ~n55256;
  assign n55258 = ~pi228 & ~n55257;
  assign n55259 = pi123 & pi262;
  assign n55260 = ~pi123 & ~pi1142;
  assign n55261 = pi228 & ~n55260;
  assign n55262 = pi228 & ~n55259;
  assign n55263 = ~n55260 & n55262;
  assign n55264 = ~n55259 & n55261;
  assign n55265 = ~n55258 & ~n61414;
  assign n55266 = n51059 & n61413;
  assign n55267 = ~n55265 & ~n55266;
  assign n55268 = pi208 & ~n55267;
  assign n55269 = ~n55255 & ~n55268;
  assign n55270 = ~pi299 & ~n55269;
  assign n55271 = ~n49381 & ~n61240;
  assign n55272 = n55265 & ~n55271;
  assign n55273 = ~pi299 & ~n49819;
  assign n55274 = ~pi262 & ~n61413;
  assign n55275 = ~n55273 & ~n55274;
  assign n55276 = ~n61240 & n55275;
  assign n55277 = n58992 & ~n55276;
  assign n55278 = ~n55272 & n55277;
  assign n55279 = ~n61240 & ~n55274;
  assign n55280 = n49374 & ~n55255;
  assign n55281 = n55279 & ~n55280;
  assign n55282 = ~n55265 & ~n55281;
  assign n55283 = ~pi207 & n55274;
  assign n55284 = ~pi208 & ~n55283;
  assign n55285 = ~n61240 & ~n55284;
  assign n55286 = ~n55282 & ~n55285;
  assign n55287 = pi299 & ~n55279;
  assign n55288 = ~n51060 & n61413;
  assign n55289 = ~pi299 & ~n55288;
  assign n55290 = ~n55265 & n55289;
  assign n55291 = pi208 & ~n55290;
  assign n55292 = ~n55287 & n55291;
  assign n55293 = n58992 & ~n55292;
  assign n55294 = ~n55286 & n55293;
  assign n55295 = ~n55270 & n55278;
  assign n55296 = ~n51202 & n61413;
  assign n55297 = ~n58992 & ~n55265;
  assign n55298 = ~n55296 & n55297;
  assign n55299 = ~n61415 & ~n55298;
  assign n55300 = ~pi284 & ~n61413;
  assign n55301 = pi1143 & n61413;
  assign n55302 = ~n51492 & n55301;
  assign n55303 = ~n55300 & ~n55302;
  assign n55304 = pi266 & pi992;
  assign n55305 = ~pi280 & n55304;
  assign n55306 = ~pi269 & n55305;
  assign n55307 = ~pi281 & n55306;
  assign n55308 = n45890 & n55307;
  assign n55309 = ~pi264 & n55308;
  assign n55310 = ~pi265 & n55309;
  assign po959 = ~pi274 & n55310;
  assign n55312 = pi274 & ~n55310;
  assign po816 = ~po959 & ~n55312;
  assign n55314 = pi265 & ~n55309;
  assign po976 = ~n55310 & ~n55314;
  assign n55316 = ~pi282 & n55307;
  assign n55317 = ~pi270 & n55316;
  assign n55318 = pi277 & ~n55317;
  assign po977 = ~n55308 & ~n55318;
  assign n55320 = pi270 & ~n55316;
  assign po962 = ~n55317 & ~n55320;
  assign n55322 = pi282 & ~n55307;
  assign po992 = ~n55316 & ~n55322;
  assign n55324 = pi269 & ~n55305;
  assign po974 = ~n55306 & ~n55324;
  assign n55326 = pi280 & ~n55304;
  assign po1070 = ~n55305 & ~n55326;
  assign n55328 = pi311 & ~pi312;
  assign po1080 = n55019 & n55328;
  assign n55330 = ~pi266 & ~pi992;
  assign po1104 = ~n55304 & ~n55330;
  assign n55332 = ~pi949 & pi954;
  assign n55333 = pi313 & ~pi954;
  assign n55334 = ~pi313 & ~pi954;
  assign n55335 = pi949 & pi954;
  assign n55336 = ~n55334 & ~n55335;
  assign n55337 = ~n55332 & ~n55333;
  assign n55338 = n58992 & n44138;
  assign n55339 = n44152 & ~n44774;
  assign n55340 = ~n55338 & ~n55339;
  assign n55341 = ~pi1148 & n55340;
  assign n55342 = ~pi222 & ~pi223;
  assign n55343 = pi937 & ~n55342;
  assign n55344 = pi273 & n26651;
  assign n55345 = ~n55343 & ~n55344;
  assign n55346 = n55338 & n55345;
  assign n55347 = n35591 & ~n44774;
  assign n55348 = ~n55346 & ~n55347;
  assign n55349 = pi237 & ~n55348;
  assign n55350 = ~n6544 & n55346;
  assign n55351 = ~pi215 & n37050;
  assign n55352 = ~pi273 & n55351;
  assign n55353 = pi833 & n3906;
  assign n55354 = ~pi937 & n55353;
  assign n55355 = ~n55352 & ~n55354;
  assign n55356 = ~n44774 & ~n55355;
  assign n55357 = ~n55350 & ~n55356;
  assign n55358 = ~n55349 & n55357;
  assign po459 = ~n55341 & n55358;
  assign n55360 = pi1147 & n55340;
  assign n55361 = ~n6629 & n55339;
  assign n55362 = pi934 & ~n38239;
  assign n55363 = pi271 & n37050;
  assign n55364 = ~n55362 & ~n55363;
  assign n55365 = n55361 & ~n55364;
  assign n55366 = pi222 & ~pi934;
  assign n55367 = ~pi271 & n26651;
  assign n55368 = ~n55366 & ~n55367;
  assign n55369 = n55338 & n55368;
  assign n55370 = ~n55347 & ~n55369;
  assign n55371 = ~n55365 & n55370;
  assign n55372 = ~n55360 & n55371;
  assign n55373 = ~pi233 & ~n55372;
  assign n55374 = n55339 & n55364;
  assign n55375 = n55338 & ~n55368;
  assign n55376 = n35583 & n44774;
  assign n55377 = n58992 & n35582;
  assign n55378 = pi1147 & ~n61417;
  assign n55379 = ~n55375 & n55378;
  assign n55380 = ~n55374 & n55379;
  assign n55381 = ~n6544 & n55338;
  assign n55382 = ~n55361 & ~n55381;
  assign n55383 = ~pi1147 & ~n55382;
  assign n55384 = ~n55371 & n55383;
  assign n55385 = ~n55380 & ~n55384;
  assign n55386 = pi233 & ~n55385;
  assign n55387 = ~n55373 & ~n55386;
  assign n55388 = pi1157 & ~n44152;
  assign n55389 = pi926 & n55353;
  assign n55390 = ~pi243 & n55351;
  assign n55391 = ~n55389 & ~n55390;
  assign n55392 = ~n55388 & n55391;
  assign n55393 = ~n58992 & ~n55392;
  assign n55394 = ~n37051 & ~n37053;
  assign n55395 = ~pi243 & ~n55394;
  assign n55396 = ~n44131 & ~n44138;
  assign n55397 = ~pi1157 & n55396;
  assign n55398 = ~pi926 & ~n55396;
  assign n55399 = ~pi243 & pi1157;
  assign n55400 = ~pi299 & n55342;
  assign n55401 = pi299 & n38239;
  assign n55402 = ~n60434 & ~n55400;
  assign n55403 = ~n55399 & ~n55402;
  assign n55404 = ~n55398 & ~n55403;
  assign n55405 = ~n55397 & n55404;
  assign n55406 = ~n55395 & ~n55405;
  assign n55407 = pi299 & n35591;
  assign n55408 = ~n35582 & ~n60435;
  assign n55409 = pi926 & n55399;
  assign n55410 = ~n55408 & n55409;
  assign n55411 = n58992 & ~n55410;
  assign n55412 = ~n55406 & n55411;
  assign n55413 = pi1157 & n55396;
  assign n55414 = pi926 & ~n55396;
  assign n55415 = ~n55395 & ~n55414;
  assign n55416 = ~n55413 & n55415;
  assign n55417 = ~n55395 & n55403;
  assign n55418 = ~n55410 & ~n55417;
  assign n55419 = ~n55416 & n55418;
  assign n55420 = n58992 & ~n55419;
  assign n55421 = ~n58992 & ~n55390;
  assign n55422 = ~n55388 & ~n55389;
  assign n55423 = n55421 & n55422;
  assign n55424 = ~n55420 & ~n55423;
  assign n55425 = ~n55393 & ~n55412;
  assign n55426 = ~n58992 & ~n55351;
  assign n55427 = n58992 & n55394;
  assign n55428 = n58992 & ~n55394;
  assign n55429 = ~n58992 & n38239;
  assign n55430 = pi216 & n55429;
  assign n55431 = ~n55428 & ~n55430;
  assign n55432 = ~n55426 & ~n55427;
  assign n55433 = ~pi943 & n61419;
  assign n55434 = pi943 & n55382;
  assign n55435 = ~n55433 & ~n55434;
  assign n55436 = ~pi1151 & ~n55435;
  assign n55437 = ~n55340 & n55433;
  assign n55438 = n58992 & ~n55402;
  assign n55439 = ~n55429 & ~n55438;
  assign n55440 = ~pi275 & ~n55439;
  assign n55441 = ~n55347 & ~n61417;
  assign n55442 = pi943 & pi1151;
  assign n55443 = ~n55441 & n55442;
  assign n55444 = ~n55440 & ~n55443;
  assign n55445 = ~n55437 & ~n55440;
  assign n55446 = ~n55443 & n55445;
  assign n55447 = ~n55437 & n55444;
  assign po623 = ~n55436 & n61420;
  assign n55449 = pi1156 & ~n44152;
  assign n55450 = pi942 & n55353;
  assign n55451 = ~pi263 & n55351;
  assign n55452 = ~n55450 & ~n55451;
  assign n55453 = ~n55449 & n55452;
  assign n55454 = ~n58992 & ~n55453;
  assign n55455 = ~pi263 & ~n55394;
  assign n55456 = ~pi1156 & n55396;
  assign n55457 = ~pi942 & ~n55396;
  assign n55458 = ~pi263 & pi1156;
  assign n55459 = ~n55402 & ~n55458;
  assign n55460 = ~n55457 & ~n55459;
  assign n55461 = ~n55456 & n55460;
  assign n55462 = ~n55455 & ~n55461;
  assign n55463 = pi942 & n55458;
  assign n55464 = ~n55408 & n55463;
  assign n55465 = n58992 & ~n55464;
  assign n55466 = ~n55462 & n55465;
  assign n55467 = pi1156 & n55396;
  assign n55468 = pi942 & ~n55396;
  assign n55469 = ~n55455 & ~n55468;
  assign n55470 = ~n55467 & n55469;
  assign n55471 = ~n55455 & n55459;
  assign n55472 = ~n55464 & ~n55471;
  assign n55473 = ~n55470 & n55472;
  assign n55474 = n58992 & ~n55473;
  assign n55475 = ~n58992 & ~n55451;
  assign n55476 = ~n55449 & ~n55450;
  assign n55477 = n55475 & n55476;
  assign n55478 = ~n55474 & ~n55477;
  assign n55479 = ~n55454 & ~n55466;
  assign n55480 = pi1155 & ~n44152;
  assign n55481 = pi925 & n55353;
  assign n55482 = pi267 & n55351;
  assign n55483 = ~n55481 & ~n55482;
  assign n55484 = ~n55480 & n55483;
  assign n55485 = ~n58992 & ~n55484;
  assign n55486 = pi267 & ~n55394;
  assign n55487 = ~pi1155 & n55396;
  assign n55488 = ~pi925 & ~n55396;
  assign n55489 = pi267 & pi1155;
  assign n55490 = ~n55402 & ~n55489;
  assign n55491 = ~n55488 & ~n55490;
  assign n55492 = ~n55487 & n55491;
  assign n55493 = ~n55486 & ~n55492;
  assign n55494 = pi925 & n55489;
  assign n55495 = ~n55408 & n55494;
  assign n55496 = n58992 & ~n55495;
  assign n55497 = ~n55493 & n55496;
  assign n55498 = pi1155 & n55396;
  assign n55499 = pi925 & ~n55396;
  assign n55500 = ~n55486 & ~n55499;
  assign n55501 = ~n55498 & n55500;
  assign n55502 = ~n55486 & n55490;
  assign n55503 = ~n55495 & ~n55502;
  assign n55504 = ~n55501 & n55503;
  assign n55505 = n58992 & ~n55504;
  assign n55506 = ~n58992 & ~n55482;
  assign n55507 = ~n55480 & ~n55481;
  assign n55508 = n55506 & n55507;
  assign n55509 = ~n55505 & ~n55508;
  assign n55510 = ~n55485 & ~n55497;
  assign n55511 = pi1153 & ~n44152;
  assign n55512 = pi941 & n55353;
  assign n55513 = pi253 & n55351;
  assign n55514 = ~n55512 & ~n55513;
  assign n55515 = ~n55511 & n55514;
  assign n55516 = ~n58992 & ~n55515;
  assign n55517 = pi253 & ~n55394;
  assign n55518 = ~pi1153 & n55396;
  assign n55519 = ~pi941 & ~n55396;
  assign n55520 = pi253 & pi1153;
  assign n55521 = ~n55402 & ~n55520;
  assign n55522 = ~n55519 & ~n55521;
  assign n55523 = ~n55518 & n55522;
  assign n55524 = ~n55517 & ~n55523;
  assign n55525 = pi941 & n55520;
  assign n55526 = ~n55408 & n55525;
  assign n55527 = n58992 & ~n55526;
  assign n55528 = ~n55524 & n55527;
  assign n55529 = pi1153 & n55396;
  assign n55530 = pi941 & ~n55396;
  assign n55531 = ~n55517 & ~n55530;
  assign n55532 = ~n55529 & n55531;
  assign n55533 = ~n55517 & n55521;
  assign n55534 = ~n55526 & ~n55533;
  assign n55535 = ~n55532 & n55534;
  assign n55536 = n58992 & ~n55535;
  assign n55537 = ~n58992 & ~n55513;
  assign n55538 = ~n55511 & ~n55512;
  assign n55539 = n55537 & n55538;
  assign n55540 = ~n55536 & ~n55539;
  assign n55541 = ~n55516 & ~n55528;
  assign n55542 = pi1154 & ~n44152;
  assign n55543 = pi923 & n55353;
  assign n55544 = pi254 & n55351;
  assign n55545 = ~n55543 & ~n55544;
  assign n55546 = ~n55542 & n55545;
  assign n55547 = ~n58992 & ~n55546;
  assign n55548 = pi254 & ~n55394;
  assign n55549 = ~pi1154 & n55396;
  assign n55550 = ~pi923 & ~n55396;
  assign n55551 = pi254 & pi1154;
  assign n55552 = ~n55402 & ~n55551;
  assign n55553 = ~n55550 & ~n55552;
  assign n55554 = ~n55549 & n55553;
  assign n55555 = ~n55548 & ~n55554;
  assign n55556 = pi923 & n55551;
  assign n55557 = ~n55408 & n55556;
  assign n55558 = n58992 & ~n55557;
  assign n55559 = ~n55555 & n55558;
  assign n55560 = pi1154 & n55396;
  assign n55561 = pi923 & ~n55396;
  assign n55562 = ~n55548 & ~n55561;
  assign n55563 = ~n55560 & n55562;
  assign n55564 = ~n55548 & n55552;
  assign n55565 = ~n55557 & ~n55564;
  assign n55566 = ~n55563 & n55565;
  assign n55567 = n58992 & ~n55566;
  assign n55568 = ~n58992 & ~n55544;
  assign n55569 = ~n55542 & ~n55543;
  assign n55570 = n55568 & n55569;
  assign n55571 = ~n55567 & ~n55570;
  assign n55572 = ~n55547 & ~n55559;
  assign n55573 = ~pi922 & n61419;
  assign n55574 = pi922 & n55382;
  assign n55575 = ~n55573 & ~n55574;
  assign n55576 = ~pi1152 & ~n55575;
  assign n55577 = ~n55340 & n55573;
  assign n55578 = ~pi268 & ~n55439;
  assign n55579 = pi922 & pi1152;
  assign n55580 = ~n55441 & n55579;
  assign n55581 = ~n55578 & ~n55580;
  assign n55582 = ~n55577 & ~n55578;
  assign n55583 = ~n55580 & n55582;
  assign n55584 = ~n55577 & n55581;
  assign po630 = ~n55576 & n61425;
  assign n55586 = ~pi931 & n61419;
  assign n55587 = pi931 & n55382;
  assign n55588 = ~n55586 & ~n55587;
  assign n55589 = ~pi1150 & ~n55588;
  assign n55590 = ~n55340 & n55586;
  assign n55591 = ~pi272 & ~n55439;
  assign n55592 = pi931 & pi1150;
  assign n55593 = ~n55441 & n55592;
  assign n55594 = ~n55591 & ~n55593;
  assign n55595 = ~n55590 & ~n55591;
  assign n55596 = ~n55593 & n55595;
  assign n55597 = ~n55590 & n55594;
  assign po631 = ~n55589 & n61426;
  assign n55599 = ~pi936 & n61419;
  assign n55600 = pi936 & n55382;
  assign n55601 = ~n55599 & ~n55600;
  assign n55602 = ~pi1149 & ~n55601;
  assign n55603 = ~n55340 & n55599;
  assign n55604 = ~pi283 & ~n55439;
  assign n55605 = pi936 & pi1149;
  assign n55606 = ~n55441 & n55605;
  assign n55607 = ~n55604 & ~n55606;
  assign n55608 = ~n55603 & ~n55604;
  assign n55609 = ~n55606 & n55608;
  assign n55610 = ~n55603 & n55607;
  assign po632 = ~n55602 & n61427;
  assign n55612 = ~pi241 & ~pi506;
  assign n55613 = pi241 & pi506;
  assign n55614 = ~n55612 & ~n55613;
  assign n55615 = pi234 & n45852;
  assign n55616 = pi557 & ~n55615;
  assign n55617 = ~pi557 & ~n55146;
  assign n55618 = ~pi246 & ~pi536;
  assign n55619 = pi246 & pi536;
  assign n55620 = ~n55618 & ~n55619;
  assign n55621 = pi249 & ~pi538;
  assign n55622 = ~pi249 & pi538;
  assign n55623 = ~pi249 & ~pi538;
  assign n55624 = pi249 & pi538;
  assign n55625 = ~n55623 & ~n55624;
  assign n55626 = ~n55621 & ~n55622;
  assign n55627 = pi248 & ~pi537;
  assign n55628 = ~pi248 & pi537;
  assign n55629 = ~n55627 & ~n55628;
  assign n55630 = ~n61428 & n55629;
  assign n55631 = ~n55620 & n55630;
  assign n55632 = ~n55617 & n55631;
  assign n55633 = ~n55617 & ~n55620;
  assign n55634 = ~n55616 & n55633;
  assign n55635 = ~pi538 & n55634;
  assign n55636 = ~pi249 & ~n55635;
  assign n55637 = pi538 & n55634;
  assign n55638 = pi249 & ~n55637;
  assign n55639 = ~n55636 & ~n55638;
  assign n55640 = ~n61428 & n55634;
  assign n55641 = ~pi537 & n61429;
  assign n55642 = ~pi248 & ~n55641;
  assign n55643 = pi537 & n61429;
  assign n55644 = pi248 & ~n55643;
  assign n55645 = ~n55642 & ~n55644;
  assign n55646 = ~n55616 & n55632;
  assign n55647 = ~n55614 & n61430;
  assign n55648 = ~pi240 & ~pi535;
  assign n55649 = pi240 & pi535;
  assign n55650 = ~n55648 & ~n55649;
  assign n55651 = n55647 & ~n55650;
  assign n55652 = pi534 & n55651;
  assign n55653 = ~pi239 & ~n55652;
  assign n55654 = ~pi534 & n55651;
  assign n55655 = pi239 & ~n55654;
  assign n55656 = ~n55653 & ~n55655;
  assign n55657 = pi504 & n55656;
  assign n55658 = pi242 & ~n55657;
  assign n55659 = ~pi504 & n55656;
  assign n55660 = ~pi242 & ~n55659;
  assign n55661 = ~n55658 & ~n55660;
  assign n55662 = pi533 & n55661;
  assign n55663 = pi235 & ~n55662;
  assign n55664 = ~pi533 & n55661;
  assign n55665 = ~pi235 & ~n55664;
  assign n55666 = ~n55663 & ~n55665;
  assign n55667 = pi558 & n55666;
  assign n55668 = pi244 & ~n55667;
  assign n55669 = ~pi558 & n55666;
  assign n55670 = ~pi244 & ~n55669;
  assign n55671 = ~n55668 & ~n55670;
  assign n55672 = pi509 & n55671;
  assign n55673 = pi245 & ~n55672;
  assign n55674 = ~pi509 & n55671;
  assign n55675 = ~pi245 & ~n55674;
  assign n55676 = ~n55673 & ~n55675;
  assign n55677 = pi508 & n55676;
  assign n55678 = pi247 & ~n55677;
  assign n55679 = pi234 & n45855;
  assign n55680 = pi511 & ~n55679;
  assign n55681 = ~pi511 & ~n55168;
  assign n55682 = ~pi248 & ~pi481;
  assign n55683 = pi248 & pi481;
  assign n55684 = ~n55682 & ~n55683;
  assign n55685 = pi249 & ~pi579;
  assign n55686 = ~pi249 & pi579;
  assign n55687 = ~pi249 & ~pi579;
  assign n55688 = pi249 & pi579;
  assign n55689 = ~n55687 & ~n55688;
  assign n55690 = ~n55685 & ~n55686;
  assign n55691 = pi246 & ~pi487;
  assign n55692 = ~pi246 & pi487;
  assign n55693 = pi246 & pi487;
  assign n55694 = ~pi246 & ~pi487;
  assign n55695 = ~n55693 & ~n55694;
  assign n55696 = ~n55691 & ~n55692;
  assign n55697 = ~n61431 & ~n61432;
  assign n55698 = ~n55684 & n55697;
  assign n55699 = ~n55681 & n55698;
  assign n55700 = ~n55681 & ~n61432;
  assign n55701 = ~n55680 & n55700;
  assign n55702 = ~n61431 & n55701;
  assign n55703 = ~n55684 & n55702;
  assign n55704 = ~n55680 & n55699;
  assign n55705 = pi559 & n61433;
  assign n55706 = pi241 & ~n55705;
  assign n55707 = ~pi559 & n61433;
  assign n55708 = ~pi241 & ~n55707;
  assign n55709 = ~n55706 & ~n55708;
  assign n55710 = pi515 & n55709;
  assign n55711 = pi240 & ~n55710;
  assign n55712 = ~pi506 & n61430;
  assign n55713 = n55708 & ~n55712;
  assign n55714 = pi506 & n61430;
  assign n55715 = n55706 & ~n55714;
  assign n55716 = n55623 & n55634;
  assign n55717 = n61431 & ~n55716;
  assign n55718 = ~pi579 & ~n55702;
  assign n55719 = ~n55636 & n55701;
  assign n55720 = pi579 & ~n55719;
  assign n55721 = ~n55718 & ~n55720;
  assign n55722 = n55701 & ~n55717;
  assign n55723 = ~n61429 & ~n61434;
  assign n55724 = ~pi537 & ~n55723;
  assign n55725 = pi537 & n55702;
  assign n55726 = ~pi248 & ~n55725;
  assign n55727 = ~n55724 & n55726;
  assign n55728 = ~n55644 & ~n55727;
  assign n55729 = ~pi481 & ~n55728;
  assign n55730 = pi537 & ~n55723;
  assign n55731 = ~pi537 & n55702;
  assign n55732 = pi248 & ~n55731;
  assign n55733 = ~n55730 & n55732;
  assign n55734 = ~n55642 & ~n55733;
  assign n55735 = pi481 & ~n55734;
  assign n55736 = ~n55729 & ~n55735;
  assign n55737 = ~pi559 & n55736;
  assign n55738 = pi559 & n61430;
  assign n55739 = ~pi241 & ~n55738;
  assign n55740 = ~n55737 & n55739;
  assign n55741 = ~n55706 & ~n55740;
  assign n55742 = ~pi506 & ~n55741;
  assign n55743 = pi559 & n55736;
  assign n55744 = ~pi559 & n61430;
  assign n55745 = pi241 & ~n55744;
  assign n55746 = ~n55743 & n55745;
  assign n55747 = ~n55708 & ~n55746;
  assign n55748 = pi506 & ~n55747;
  assign n55749 = ~n55742 & ~n55748;
  assign n55750 = ~n55713 & ~n55715;
  assign n55751 = ~pi515 & n61435;
  assign n55752 = pi515 & n55647;
  assign n55753 = ~pi240 & ~n55752;
  assign n55754 = ~n55751 & n55753;
  assign n55755 = ~n55711 & ~n55754;
  assign n55756 = ~pi535 & ~n55755;
  assign n55757 = ~pi515 & n55709;
  assign n55758 = ~pi240 & ~n55757;
  assign n55759 = pi515 & n61435;
  assign n55760 = ~pi515 & n55647;
  assign n55761 = pi240 & ~n55760;
  assign n55762 = ~n55759 & n55761;
  assign n55763 = ~n55758 & ~n55762;
  assign n55764 = pi535 & ~n55763;
  assign n55765 = ~n55756 & ~n55764;
  assign n55766 = ~pi534 & n55765;
  assign n55767 = ~n55711 & ~n55758;
  assign n55768 = pi534 & n55767;
  assign n55769 = pi239 & ~n55768;
  assign n55770 = ~n55766 & n55769;
  assign n55771 = ~n55653 & ~n55770;
  assign n55772 = ~pi488 & ~n55771;
  assign n55773 = pi534 & n55765;
  assign n55774 = ~pi534 & n55767;
  assign n55775 = ~pi239 & ~n55774;
  assign n55776 = ~n55773 & n55775;
  assign n55777 = ~n55655 & ~n55776;
  assign n55778 = pi488 & ~n55777;
  assign n55779 = ~n55772 & ~n55778;
  assign n55780 = ~pi504 & n55779;
  assign n55781 = pi239 & ~pi488;
  assign n55782 = ~pi239 & pi488;
  assign n55783 = ~n55781 & ~n55782;
  assign n55784 = n55767 & ~n55783;
  assign n55785 = pi504 & n55784;
  assign n55786 = ~pi242 & ~n55785;
  assign n55787 = ~n55780 & n55786;
  assign n55788 = ~n55658 & ~n55787;
  assign n55789 = ~pi510 & ~n55788;
  assign n55790 = pi504 & n55779;
  assign n55791 = ~pi504 & n55784;
  assign n55792 = pi242 & ~n55791;
  assign n55793 = ~n55790 & n55792;
  assign n55794 = ~n55660 & ~n55793;
  assign n55795 = pi510 & ~n55794;
  assign n55796 = ~n55789 & ~n55795;
  assign n55797 = ~pi533 & n55796;
  assign n55798 = ~pi242 & ~pi510;
  assign n55799 = pi242 & pi510;
  assign n55800 = ~n55798 & ~n55799;
  assign n55801 = n55784 & ~n55800;
  assign n55802 = pi533 & n55801;
  assign n55803 = ~pi235 & ~n55802;
  assign n55804 = ~n55797 & n55803;
  assign n55805 = ~n55663 & ~n55804;
  assign n55806 = ~pi512 & ~n55805;
  assign n55807 = pi533 & n55796;
  assign n55808 = ~pi533 & n55801;
  assign n55809 = pi235 & ~n55808;
  assign n55810 = ~n55807 & n55809;
  assign n55811 = ~n55665 & ~n55810;
  assign n55812 = pi512 & ~n55811;
  assign n55813 = ~n55806 & ~n55812;
  assign n55814 = ~pi558 & n55813;
  assign n55815 = ~pi235 & ~pi512;
  assign n55816 = pi235 & pi512;
  assign n55817 = ~n55815 & ~n55816;
  assign n55818 = n55801 & ~n55817;
  assign n55819 = pi558 & n55818;
  assign n55820 = ~pi244 & ~n55819;
  assign n55821 = ~n55814 & n55820;
  assign n55822 = ~n55668 & ~n55821;
  assign n55823 = ~pi513 & ~n55822;
  assign n55824 = pi558 & n55813;
  assign n55825 = ~pi558 & n55818;
  assign n55826 = pi244 & ~n55825;
  assign n55827 = ~n55824 & n55826;
  assign n55828 = ~n55670 & ~n55827;
  assign n55829 = pi513 & ~n55828;
  assign n55830 = ~n55823 & ~n55829;
  assign n55831 = ~pi509 & n55830;
  assign n55832 = ~pi244 & ~pi513;
  assign n55833 = pi244 & pi513;
  assign n55834 = ~n55832 & ~n55833;
  assign n55835 = n55818 & ~n55834;
  assign n55836 = pi509 & n55835;
  assign n55837 = ~pi245 & ~n55836;
  assign n55838 = ~n55831 & n55837;
  assign n55839 = ~n55673 & ~n55838;
  assign n55840 = ~pi514 & ~n55839;
  assign n55841 = pi509 & n55830;
  assign n55842 = ~pi509 & n55835;
  assign n55843 = pi245 & ~n55842;
  assign n55844 = ~n55841 & n55843;
  assign n55845 = ~n55675 & ~n55844;
  assign n55846 = pi514 & ~n55845;
  assign n55847 = ~n55840 & ~n55846;
  assign n55848 = ~pi508 & n55847;
  assign n55849 = ~pi245 & ~pi514;
  assign n55850 = pi245 & pi514;
  assign n55851 = ~n55849 & ~n55850;
  assign n55852 = n55835 & ~n55851;
  assign n55853 = pi508 & n55852;
  assign n55854 = ~pi247 & ~n55853;
  assign n55855 = ~n55848 & n55854;
  assign n55856 = ~n55678 & ~n55855;
  assign n55857 = ~pi516 & ~n55856;
  assign n55858 = ~pi508 & n55676;
  assign n55859 = ~pi247 & ~n55858;
  assign n55860 = pi508 & n55847;
  assign n55861 = ~pi508 & n55852;
  assign n55862 = pi247 & ~n55861;
  assign n55863 = ~n55860 & n55862;
  assign n55864 = ~n55859 & ~n55863;
  assign n55865 = pi516 & ~n55864;
  assign n55866 = ~n55857 & ~n55865;
  assign n55867 = ~pi238 & n55866;
  assign n55868 = ~pi517 & ~n55867;
  assign n55869 = ~n55678 & ~n55859;
  assign n55870 = ~pi238 & n55869;
  assign n55871 = ~pi247 & ~pi516;
  assign n55872 = pi247 & pi516;
  assign n55873 = ~n55871 & ~n55872;
  assign n55874 = n55852 & ~n55873;
  assign n55875 = pi238 & n55874;
  assign n55876 = pi517 & ~n55875;
  assign n55877 = ~n55870 & n55876;
  assign n55878 = ~pi507 & ~n55877;
  assign n55879 = ~n55868 & n55878;
  assign n55880 = pi238 & n55866;
  assign n55881 = pi517 & ~n55880;
  assign n55882 = pi238 & n55869;
  assign n55883 = ~pi238 & n55874;
  assign n55884 = ~pi517 & ~n55883;
  assign n55885 = ~n55882 & n55884;
  assign n55886 = pi507 & ~n55885;
  assign n55887 = ~n55881 & n55886;
  assign n55888 = ~n55879 & ~n55887;
  assign n55889 = pi233 & ~n55888;
  assign n55890 = ~pi247 & ~pi561;
  assign n55891 = ~pi240 & ~pi542;
  assign n55892 = pi240 & pi542;
  assign n55893 = ~n55891 & ~n55892;
  assign n55894 = pi505 & ~n55615;
  assign n55895 = ~pi505 & ~n55146;
  assign n55896 = ~pi249 & pi496;
  assign n55897 = pi246 & ~pi499;
  assign n55898 = ~n55896 & ~n55897;
  assign n55899 = pi248 & ~pi501;
  assign n55900 = ~pi248 & pi501;
  assign n55901 = ~pi248 & ~pi501;
  assign n55902 = pi248 & pi501;
  assign n55903 = ~n55901 & ~n55902;
  assign n55904 = ~n55899 & ~n55900;
  assign n55905 = n55898 & ~n61436;
  assign n55906 = ~pi241 & ~pi500;
  assign n55907 = pi241 & pi500;
  assign n55908 = ~n55906 & ~n55907;
  assign n55909 = ~pi246 & pi499;
  assign n55910 = pi249 & ~pi496;
  assign n55911 = ~n55909 & ~n55910;
  assign n55912 = ~n55908 & n55911;
  assign n55913 = ~pi246 & ~pi499;
  assign n55914 = pi246 & pi499;
  assign n55915 = ~n55913 & ~n55914;
  assign n55916 = ~n61436 & ~n55915;
  assign n55917 = ~pi249 & ~pi496;
  assign n55918 = pi249 & pi496;
  assign n55919 = ~n55896 & ~n55910;
  assign n55920 = ~n55917 & ~n55918;
  assign n55921 = ~n55908 & n61437;
  assign n55922 = n55916 & n55921;
  assign n55923 = n55905 & n55912;
  assign n55924 = ~n55895 & n61438;
  assign n55925 = ~n61436 & n61437;
  assign n55926 = ~n55915 & n55925;
  assign n55927 = ~n55894 & n55926;
  assign n55928 = ~n55895 & n55927;
  assign n55929 = ~n55908 & n55928;
  assign n55930 = ~n55894 & n55924;
  assign n55931 = ~n55893 & n61439;
  assign n55932 = pi497 & n55931;
  assign n55933 = ~pi239 & ~n55932;
  assign n55934 = ~pi497 & n55931;
  assign n55935 = pi239 & ~n55934;
  assign n55936 = ~n55933 & ~n55935;
  assign n55937 = pi539 & n55936;
  assign n55938 = pi242 & ~n55937;
  assign n55939 = ~pi539 & n55936;
  assign n55940 = ~pi242 & ~n55939;
  assign n55941 = ~n55938 & ~n55940;
  assign n55942 = pi540 & n55941;
  assign n55943 = pi235 & ~n55942;
  assign n55944 = ~pi540 & n55941;
  assign n55945 = ~pi235 & ~n55944;
  assign n55946 = ~n55943 & ~n55945;
  assign n55947 = ~pi244 & ~pi541;
  assign n55948 = pi244 & pi541;
  assign n55949 = ~n55947 & ~n55948;
  assign n55950 = n55946 & ~n55949;
  assign n55951 = ~pi245 & ~pi503;
  assign n55952 = pi245 & pi503;
  assign n55953 = ~n55951 & ~n55952;
  assign n55954 = n55950 & ~n55953;
  assign n55955 = ~pi502 & n55954;
  assign n55956 = ~pi247 & ~n55955;
  assign n55957 = ~n55890 & ~n55956;
  assign n55958 = pi518 & ~n55679;
  assign n55959 = ~pi518 & ~n55168;
  assign n55960 = ~pi246 & pi520;
  assign n55961 = pi248 & ~pi521;
  assign n55962 = ~n55960 & ~n55961;
  assign n55963 = pi249 & ~pi578;
  assign n55964 = ~pi249 & pi578;
  assign n55965 = ~pi249 & ~pi578;
  assign n55966 = pi249 & pi578;
  assign n55967 = ~n55965 & ~n55966;
  assign n55968 = ~n55963 & ~n55964;
  assign n55969 = n55962 & ~n61440;
  assign n55970 = ~pi241 & ~pi574;
  assign n55971 = pi241 & pi574;
  assign n55972 = ~n55970 & ~n55971;
  assign n55973 = ~pi248 & pi521;
  assign n55974 = pi246 & ~pi520;
  assign n55975 = ~n55973 & ~n55974;
  assign n55976 = ~n55972 & n55975;
  assign n55977 = ~pi248 & ~pi521;
  assign n55978 = pi248 & pi521;
  assign n55979 = ~n55961 & ~n55973;
  assign n55980 = ~n55977 & ~n55978;
  assign n55981 = ~n61440 & n61441;
  assign n55982 = ~pi246 & ~pi520;
  assign n55983 = pi246 & pi520;
  assign n55984 = ~n55960 & ~n55974;
  assign n55985 = ~n55982 & ~n55983;
  assign n55986 = ~n55972 & n61442;
  assign n55987 = n55981 & n55986;
  assign n55988 = n55969 & n55976;
  assign n55989 = ~n55959 & n61443;
  assign n55990 = ~n55958 & n61443;
  assign n55991 = ~n55959 & n55990;
  assign n55992 = ~n55958 & n55989;
  assign n55993 = pi582 & n61444;
  assign n55994 = pi240 & ~n55993;
  assign n55995 = ~pi582 & n61444;
  assign n55996 = ~pi240 & ~n55995;
  assign n55997 = ~n55994 & ~n55996;
  assign n55998 = pi239 & ~pi519;
  assign n55999 = ~pi239 & pi519;
  assign n56000 = ~n55998 & ~n55999;
  assign n56001 = n55997 & ~n56000;
  assign n56002 = ~pi242 & ~pi586;
  assign n56003 = pi242 & pi586;
  assign n56004 = ~n56002 & ~n56003;
  assign n56005 = n56001 & ~n56004;
  assign n56006 = ~pi235 & ~pi581;
  assign n56007 = pi235 & pi581;
  assign n56008 = ~n56006 & ~n56007;
  assign n56009 = n56005 & ~n56008;
  assign n56010 = pi585 & n56009;
  assign n56011 = pi244 & ~n56010;
  assign n56012 = ~pi585 & n56009;
  assign n56013 = ~pi244 & ~n56012;
  assign n56014 = ~n56011 & ~n56013;
  assign n56015 = pi584 & n56014;
  assign n56016 = pi245 & ~n56015;
  assign n56017 = ~pi542 & n61439;
  assign n56018 = n55996 & ~n56017;
  assign n56019 = pi542 & n61439;
  assign n56020 = n55994 & ~n56019;
  assign n56021 = ~pi500 & n61439;
  assign n56022 = n55907 & n55928;
  assign n56023 = ~n61444 & ~n56022;
  assign n56024 = ~n56021 & n56023;
  assign n56025 = ~pi582 & ~n56024;
  assign n56026 = pi582 & n61439;
  assign n56027 = ~pi240 & ~n56026;
  assign n56028 = ~n56025 & n56027;
  assign n56029 = ~n55994 & ~n56028;
  assign n56030 = ~pi542 & ~n56029;
  assign n56031 = pi582 & ~n56024;
  assign n56032 = ~pi582 & n61439;
  assign n56033 = pi240 & ~n56032;
  assign n56034 = ~n56031 & n56033;
  assign n56035 = ~n55996 & ~n56034;
  assign n56036 = pi542 & ~n56035;
  assign n56037 = ~n56030 & ~n56036;
  assign n56038 = ~n56018 & ~n56020;
  assign n56039 = ~pi497 & n61445;
  assign n56040 = pi497 & n55997;
  assign n56041 = pi239 & ~n56040;
  assign n56042 = ~n56039 & n56041;
  assign n56043 = ~n55933 & ~n56042;
  assign n56044 = ~pi519 & ~n56043;
  assign n56045 = pi497 & n61445;
  assign n56046 = ~pi497 & n55997;
  assign n56047 = ~pi239 & ~n56046;
  assign n56048 = ~n56045 & n56047;
  assign n56049 = ~n55935 & ~n56048;
  assign n56050 = pi519 & ~n56049;
  assign n56051 = ~n56044 & ~n56050;
  assign n56052 = ~pi539 & n56051;
  assign n56053 = pi539 & n56001;
  assign n56054 = ~pi242 & ~n56053;
  assign n56055 = ~n56052 & n56054;
  assign n56056 = ~n55938 & ~n56055;
  assign n56057 = ~pi586 & ~n56056;
  assign n56058 = pi539 & n56051;
  assign n56059 = ~pi539 & n56001;
  assign n56060 = pi242 & ~n56059;
  assign n56061 = ~n56058 & n56060;
  assign n56062 = ~n55940 & ~n56061;
  assign n56063 = pi586 & ~n56062;
  assign n56064 = ~n56057 & ~n56063;
  assign n56065 = ~pi540 & n56064;
  assign n56066 = pi540 & n56005;
  assign n56067 = ~pi235 & ~n56066;
  assign n56068 = ~n56065 & n56067;
  assign n56069 = ~n55943 & ~n56068;
  assign n56070 = ~pi581 & ~n56069;
  assign n56071 = pi540 & n56064;
  assign n56072 = ~pi540 & n56005;
  assign n56073 = pi235 & ~n56072;
  assign n56074 = ~n56071 & n56073;
  assign n56075 = ~n55945 & ~n56074;
  assign n56076 = pi581 & ~n56075;
  assign n56077 = ~n56070 & ~n56076;
  assign n56078 = ~pi585 & n56077;
  assign n56079 = pi585 & n55946;
  assign n56080 = ~pi244 & ~n56079;
  assign n56081 = ~n56078 & n56080;
  assign n56082 = ~n56011 & ~n56081;
  assign n56083 = ~pi541 & ~n56082;
  assign n56084 = pi585 & n56077;
  assign n56085 = ~pi585 & n55946;
  assign n56086 = pi244 & ~n56085;
  assign n56087 = ~n56084 & n56086;
  assign n56088 = ~n56013 & ~n56087;
  assign n56089 = pi541 & ~n56088;
  assign n56090 = ~n56083 & ~n56089;
  assign n56091 = ~pi584 & n56090;
  assign n56092 = pi584 & n55950;
  assign n56093 = ~pi245 & ~n56092;
  assign n56094 = ~n56091 & n56093;
  assign n56095 = ~n56016 & ~n56094;
  assign n56096 = ~pi503 & ~n56095;
  assign n56097 = ~pi584 & n56014;
  assign n56098 = ~pi245 & ~n56097;
  assign n56099 = pi584 & n56090;
  assign n56100 = ~pi584 & n55950;
  assign n56101 = pi245 & ~n56100;
  assign n56102 = ~n56099 & n56101;
  assign n56103 = ~n56098 & ~n56102;
  assign n56104 = pi503 & ~n56103;
  assign n56105 = ~n56096 & ~n56104;
  assign n56106 = ~pi502 & ~n56105;
  assign n56107 = ~n56016 & ~n56098;
  assign n56108 = pi502 & ~n56107;
  assign n56109 = ~pi561 & ~n56108;
  assign n56110 = ~n56106 & n56109;
  assign n56111 = ~n55957 & ~n56110;
  assign n56112 = pi247 & pi561;
  assign n56113 = pi502 & n55954;
  assign n56114 = pi247 & ~n56113;
  assign n56115 = ~n56112 & ~n56114;
  assign n56116 = pi502 & ~n56105;
  assign n56117 = ~pi502 & ~n56107;
  assign n56118 = pi561 & ~n56117;
  assign n56119 = ~n56116 & n56118;
  assign n56120 = ~n56115 & ~n56119;
  assign n56121 = ~n56111 & ~n56120;
  assign n56122 = ~pi238 & n56121;
  assign n56123 = ~pi522 & ~n56122;
  assign n56124 = ~n55956 & ~n56114;
  assign n56125 = ~pi238 & n56124;
  assign n56126 = ~n55890 & ~n56112;
  assign n56127 = n56107 & ~n56126;
  assign n56128 = pi238 & n56127;
  assign n56129 = pi522 & ~n56128;
  assign n56130 = ~n56125 & n56129;
  assign n56131 = ~pi543 & ~n56130;
  assign n56132 = ~n56123 & n56131;
  assign n56133 = pi238 & n56121;
  assign n56134 = pi522 & ~n56133;
  assign n56135 = pi238 & n56124;
  assign n56136 = ~pi238 & n56127;
  assign n56137 = ~pi522 & ~n56136;
  assign n56138 = ~n56135 & n56137;
  assign n56139 = pi543 & ~n56138;
  assign n56140 = ~n56134 & n56139;
  assign n56141 = ~n56132 & ~n56140;
  assign n56142 = ~pi233 & ~n56141;
  assign n56143 = pi237 & ~n56142;
  assign n56144 = ~n55889 & n56143;
  assign n56145 = ~pi240 & ~pi492;
  assign n56146 = pi240 & pi492;
  assign n56147 = ~n56145 & ~n56146;
  assign n56148 = ~pi241 & ~pi490;
  assign n56149 = pi241 & pi490;
  assign n56150 = ~n56148 & ~n56149;
  assign n56151 = ~pi544 & ~n55146;
  assign n56152 = pi544 & ~n55615;
  assign n56153 = ~pi248 & ~pi548;
  assign n56154 = pi248 & pi548;
  assign n56155 = ~n56153 & ~n56154;
  assign n56156 = pi246 & ~pi546;
  assign n56157 = ~pi246 & pi546;
  assign n56158 = pi246 & pi546;
  assign n56159 = ~pi246 & ~pi546;
  assign n56160 = ~n56158 & ~n56159;
  assign n56161 = ~n56156 & ~n56157;
  assign n56162 = pi249 & ~pi484;
  assign n56163 = ~pi249 & pi484;
  assign n56164 = pi249 & pi484;
  assign n56165 = ~pi249 & ~pi484;
  assign n56166 = ~n56164 & ~n56165;
  assign n56167 = ~n56162 & ~n56163;
  assign n56168 = ~n61446 & ~n61447;
  assign n56169 = ~n56155 & ~n61447;
  assign n56170 = ~n61446 & n56169;
  assign n56171 = ~n56155 & n56168;
  assign n56172 = ~n56152 & n61448;
  assign n56173 = ~n56151 & n61448;
  assign n56174 = ~n56152 & n56173;
  assign n56175 = ~n56151 & n56172;
  assign n56176 = ~n56150 & n61449;
  assign n56177 = ~n56147 & n56176;
  assign n56178 = pi494 & n56177;
  assign n56179 = ~pi239 & ~n56178;
  assign n56180 = ~pi494 & n56177;
  assign n56181 = pi239 & ~n56180;
  assign n56182 = ~n56179 & ~n56181;
  assign n56183 = pi483 & n56182;
  assign n56184 = pi242 & ~n56183;
  assign n56185 = ~pi483 & n56182;
  assign n56186 = ~pi242 & ~n56185;
  assign n56187 = ~n56184 & ~n56186;
  assign n56188 = pi495 & n56187;
  assign n56189 = pi235 & ~n56188;
  assign n56190 = ~pi495 & n56187;
  assign n56191 = ~pi235 & ~n56190;
  assign n56192 = ~n56189 & ~n56191;
  assign n56193 = ~pi244 & ~pi493;
  assign n56194 = pi244 & pi493;
  assign n56195 = ~n56193 & ~n56194;
  assign n56196 = n56192 & ~n56195;
  assign n56197 = pi545 & n56196;
  assign n56198 = pi245 & ~n56197;
  assign n56199 = ~pi545 & n56196;
  assign n56200 = ~pi245 & ~n56199;
  assign n56201 = ~n56198 & ~n56200;
  assign n56202 = pi547 & n56201;
  assign n56203 = pi247 & ~n56202;
  assign n56204 = pi523 & ~n55679;
  assign n56205 = ~pi523 & ~n55168;
  assign n56206 = ~pi248 & ~pi576;
  assign n56207 = pi248 & pi576;
  assign n56208 = ~n56206 & ~n56207;
  assign n56209 = pi246 & ~pi526;
  assign n56210 = ~pi246 & pi526;
  assign n56211 = pi246 & pi526;
  assign n56212 = ~pi246 & ~pi526;
  assign n56213 = ~n56211 & ~n56212;
  assign n56214 = ~n56209 & ~n56210;
  assign n56215 = pi249 & ~pi528;
  assign n56216 = ~pi249 & pi528;
  assign n56217 = pi249 & pi528;
  assign n56218 = ~pi249 & ~pi528;
  assign n56219 = ~n56217 & ~n56218;
  assign n56220 = ~n56215 & ~n56216;
  assign n56221 = ~n61450 & ~n61451;
  assign n56222 = ~n56208 & ~n61451;
  assign n56223 = ~n61450 & n56222;
  assign n56224 = ~n56208 & n56221;
  assign n56225 = ~n56205 & n61452;
  assign n56226 = ~n56204 & n61452;
  assign n56227 = ~n56205 & n56226;
  assign n56228 = ~n56204 & n56225;
  assign n56229 = pi571 & n61453;
  assign n56230 = pi241 & ~n56229;
  assign n56231 = ~pi571 & n61453;
  assign n56232 = ~pi241 & ~n56231;
  assign n56233 = ~n56230 & ~n56232;
  assign n56234 = ~pi530 & n56233;
  assign n56235 = ~pi240 & ~n56234;
  assign n56236 = pi530 & n56233;
  assign n56237 = pi240 & ~n56236;
  assign n56238 = ~n56235 & ~n56237;
  assign n56239 = pi239 & ~pi524;
  assign n56240 = ~pi239 & pi524;
  assign n56241 = ~n56239 & ~n56240;
  assign n56242 = n56238 & ~n56241;
  assign n56243 = ~pi242 & ~pi573;
  assign n56244 = pi242 & pi573;
  assign n56245 = ~n56243 & ~n56244;
  assign n56246 = n56242 & ~n56245;
  assign n56247 = ~pi235 & ~pi575;
  assign n56248 = pi235 & pi575;
  assign n56249 = ~n56247 & ~n56248;
  assign n56250 = n56246 & ~n56249;
  assign n56251 = pi572 & n56250;
  assign n56252 = pi244 & ~n56251;
  assign n56253 = ~n56145 & ~n56235;
  assign n56254 = ~pi490 & n61449;
  assign n56255 = n56232 & ~n56254;
  assign n56256 = pi490 & n61449;
  assign n56257 = n56230 & ~n56256;
  assign n56258 = ~pi241 & ~n61449;
  assign n56259 = ~n56231 & n56258;
  assign n56260 = ~n56230 & ~n56259;
  assign n56261 = ~pi490 & ~n56260;
  assign n56262 = pi241 & ~n61449;
  assign n56263 = ~n56229 & n56262;
  assign n56264 = ~n56232 & ~n56263;
  assign n56265 = pi490 & ~n56264;
  assign n56266 = ~n56261 & ~n56265;
  assign n56267 = ~n56255 & ~n56257;
  assign n56268 = ~pi530 & ~n61454;
  assign n56269 = pi530 & ~n56176;
  assign n56270 = ~pi492 & ~n56269;
  assign n56271 = ~n56268 & n56270;
  assign n56272 = ~n56253 & ~n56271;
  assign n56273 = ~n56146 & ~n56237;
  assign n56274 = pi530 & ~n61454;
  assign n56275 = ~pi530 & ~n56176;
  assign n56276 = pi492 & ~n56275;
  assign n56277 = ~n56274 & n56276;
  assign n56278 = ~n56273 & ~n56277;
  assign n56279 = ~n56272 & ~n56278;
  assign n56280 = ~pi494 & n56279;
  assign n56281 = pi494 & n56238;
  assign n56282 = pi239 & ~n56281;
  assign n56283 = ~n56280 & n56282;
  assign n56284 = ~n56179 & ~n56283;
  assign n56285 = ~pi524 & ~n56284;
  assign n56286 = pi494 & n56279;
  assign n56287 = ~pi494 & n56238;
  assign n56288 = ~pi239 & ~n56287;
  assign n56289 = ~n56286 & n56288;
  assign n56290 = ~n56181 & ~n56289;
  assign n56291 = pi524 & ~n56290;
  assign n56292 = ~n56285 & ~n56291;
  assign n56293 = ~pi483 & n56292;
  assign n56294 = pi483 & n56242;
  assign n56295 = ~pi242 & ~n56294;
  assign n56296 = ~n56293 & n56295;
  assign n56297 = ~n56184 & ~n56296;
  assign n56298 = ~pi573 & ~n56297;
  assign n56299 = pi483 & n56292;
  assign n56300 = ~pi483 & n56242;
  assign n56301 = pi242 & ~n56300;
  assign n56302 = ~n56299 & n56301;
  assign n56303 = ~n56186 & ~n56302;
  assign n56304 = pi573 & ~n56303;
  assign n56305 = ~n56298 & ~n56304;
  assign n56306 = ~pi495 & n56305;
  assign n56307 = pi495 & n56246;
  assign n56308 = ~pi235 & ~n56307;
  assign n56309 = ~n56306 & n56308;
  assign n56310 = ~n56189 & ~n56309;
  assign n56311 = ~pi575 & ~n56310;
  assign n56312 = pi495 & n56305;
  assign n56313 = ~pi495 & n56246;
  assign n56314 = pi235 & ~n56313;
  assign n56315 = ~n56312 & n56314;
  assign n56316 = ~n56191 & ~n56315;
  assign n56317 = pi575 & ~n56316;
  assign n56318 = ~n56311 & ~n56317;
  assign n56319 = ~pi572 & n56318;
  assign n56320 = pi572 & n56192;
  assign n56321 = ~pi244 & ~n56320;
  assign n56322 = ~n56319 & n56321;
  assign n56323 = ~n56252 & ~n56322;
  assign n56324 = ~pi493 & ~n56323;
  assign n56325 = ~pi572 & n56250;
  assign n56326 = ~pi244 & ~n56325;
  assign n56327 = pi572 & n56318;
  assign n56328 = ~pi572 & n56192;
  assign n56329 = pi244 & ~n56328;
  assign n56330 = ~n56327 & n56329;
  assign n56331 = ~n56326 & ~n56330;
  assign n56332 = pi493 & ~n56331;
  assign n56333 = ~n56324 & ~n56332;
  assign n56334 = ~pi545 & n56333;
  assign n56335 = ~n56252 & ~n56326;
  assign n56336 = pi545 & n56335;
  assign n56337 = ~pi245 & ~n56336;
  assign n56338 = ~n56334 & n56337;
  assign n56339 = ~n56198 & ~n56338;
  assign n56340 = ~pi525 & ~n56339;
  assign n56341 = pi545 & n56333;
  assign n56342 = ~pi545 & n56335;
  assign n56343 = pi245 & ~n56342;
  assign n56344 = ~n56341 & n56343;
  assign n56345 = ~n56200 & ~n56344;
  assign n56346 = pi525 & ~n56345;
  assign n56347 = ~n56340 & ~n56346;
  assign n56348 = ~pi547 & n56347;
  assign n56349 = ~pi245 & ~pi525;
  assign n56350 = pi245 & pi525;
  assign n56351 = ~n56349 & ~n56350;
  assign n56352 = n56335 & ~n56351;
  assign n56353 = pi547 & n56352;
  assign n56354 = ~pi247 & ~n56353;
  assign n56355 = ~n56348 & n56354;
  assign n56356 = ~n56203 & ~n56355;
  assign n56357 = ~pi527 & ~n56356;
  assign n56358 = ~pi547 & n56201;
  assign n56359 = ~pi247 & ~n56358;
  assign n56360 = pi547 & n56347;
  assign n56361 = ~pi547 & n56352;
  assign n56362 = pi247 & ~n56361;
  assign n56363 = ~n56360 & n56362;
  assign n56364 = ~n56359 & ~n56363;
  assign n56365 = pi527 & ~n56364;
  assign n56366 = ~n56357 & ~n56365;
  assign n56367 = ~pi238 & n56366;
  assign n56368 = ~pi529 & ~n56367;
  assign n56369 = ~n56203 & ~n56359;
  assign n56370 = ~pi238 & n56369;
  assign n56371 = ~pi247 & ~pi527;
  assign n56372 = pi247 & pi527;
  assign n56373 = ~n56371 & ~n56372;
  assign n56374 = n56352 & ~n56373;
  assign n56375 = pi238 & n56374;
  assign n56376 = pi529 & ~n56375;
  assign n56377 = ~n56370 & n56376;
  assign n56378 = ~pi491 & ~n56377;
  assign n56379 = ~n56368 & n56378;
  assign n56380 = pi238 & n56366;
  assign n56381 = pi529 & ~n56380;
  assign n56382 = pi238 & n56369;
  assign n56383 = ~pi238 & n56374;
  assign n56384 = ~pi529 & ~n56383;
  assign n56385 = ~n56382 & n56384;
  assign n56386 = pi491 & ~n56385;
  assign n56387 = ~n56381 & n56386;
  assign n56388 = ~n56379 & ~n56387;
  assign n56389 = pi233 & ~n56388;
  assign n56390 = pi485 & ~n55615;
  assign n56391 = ~pi485 & ~n55146;
  assign n56392 = ~pi241 & ~pi553;
  assign n56393 = pi241 & pi553;
  assign n56394 = pi241 & ~pi553;
  assign n56395 = ~pi241 & pi553;
  assign n56396 = ~n56394 & ~n56395;
  assign n56397 = ~n56392 & ~n56393;
  assign n56398 = ~pi246 & pi563;
  assign n56399 = pi248 & ~pi554;
  assign n56400 = ~n56398 & ~n56399;
  assign n56401 = pi242 & ~pi489;
  assign n56402 = ~pi242 & pi489;
  assign n56403 = ~n56401 & ~n56402;
  assign n56404 = n56400 & n56403;
  assign n56405 = n61455 & n56404;
  assign n56406 = ~pi240 & pi551;
  assign n56407 = ~pi239 & ~pi550;
  assign n56408 = ~n56406 & ~n56407;
  assign n56409 = pi240 & ~pi551;
  assign n56410 = pi246 & ~pi563;
  assign n56411 = ~n56409 & ~n56410;
  assign n56412 = n56408 & n56411;
  assign n56413 = ~pi248 & pi554;
  assign n56414 = ~pi249 & pi555;
  assign n56415 = ~n56413 & ~n56414;
  assign n56416 = pi249 & ~pi555;
  assign n56417 = pi239 & pi550;
  assign n56418 = ~n56416 & ~n56417;
  assign n56419 = n56415 & n56418;
  assign n56420 = n56412 & n56419;
  assign n56421 = n56405 & n56420;
  assign n56422 = ~n56391 & n56421;
  assign n56423 = ~n56414 & ~n56416;
  assign n56424 = n61455 & n56423;
  assign n56425 = pi240 & pi551;
  assign n56426 = ~pi240 & ~pi551;
  assign n56427 = ~n56425 & ~n56426;
  assign n56428 = ~pi248 & ~pi554;
  assign n56429 = pi248 & pi554;
  assign n56430 = ~n56399 & ~n56413;
  assign n56431 = ~n56428 & ~n56429;
  assign n56432 = ~pi246 & ~pi563;
  assign n56433 = pi246 & pi563;
  assign n56434 = ~n56398 & ~n56410;
  assign n56435 = ~n56432 & ~n56433;
  assign n56436 = n61456 & n61457;
  assign n56437 = ~n56427 & n56436;
  assign n56438 = n56424 & ~n56427;
  assign n56439 = n56436 & n56438;
  assign n56440 = n56424 & n56437;
  assign n56441 = ~n56391 & n61458;
  assign n56442 = ~n56390 & n61458;
  assign n56443 = ~n56391 & n56442;
  assign n56444 = ~n56390 & n56441;
  assign n56445 = pi550 & n61459;
  assign n56446 = ~pi239 & ~n56445;
  assign n56447 = ~pi550 & n61459;
  assign n56448 = pi239 & ~n56447;
  assign n56449 = ~n56446 & ~n56448;
  assign n56450 = ~pi489 & n56449;
  assign n56451 = ~pi242 & ~n56450;
  assign n56452 = pi489 & n56449;
  assign n56453 = pi242 & ~n56452;
  assign n56454 = ~n56451 & ~n56453;
  assign n56455 = ~n56390 & n56422;
  assign n56456 = pi549 & n61460;
  assign n56457 = pi235 & ~n56456;
  assign n56458 = ~pi549 & n61460;
  assign n56459 = ~pi235 & ~n56458;
  assign n56460 = ~n56457 & ~n56459;
  assign n56461 = pi486 & n56460;
  assign n56462 = pi244 & ~n56461;
  assign n56463 = ~pi486 & n56460;
  assign n56464 = ~pi244 & ~n56463;
  assign n56465 = ~n56462 & ~n56464;
  assign n56466 = ~pi245 & ~pi580;
  assign n56467 = pi245 & pi580;
  assign n56468 = ~n56466 & ~n56467;
  assign n56469 = n56465 & ~n56468;
  assign n56470 = pi552 & n56469;
  assign n56471 = pi247 & ~n56470;
  assign n56472 = ~pi235 & ~pi531;
  assign n56473 = pi235 & pi531;
  assign n56474 = ~n56472 & ~n56473;
  assign n56475 = pi570 & ~n55679;
  assign n56476 = ~pi570 & ~n55168;
  assign n56477 = ~pi249 & ~pi482;
  assign n56478 = pi249 & pi482;
  assign n56479 = ~n56477 & ~n56478;
  assign n56480 = ~pi240 & pi560;
  assign n56481 = pi246 & ~pi564;
  assign n56482 = ~n56480 & ~n56481;
  assign n56483 = ~pi239 & ~pi569;
  assign n56484 = pi239 & pi569;
  assign n56485 = ~pi239 & pi569;
  assign n56486 = pi239 & ~pi569;
  assign n56487 = ~n56485 & ~n56486;
  assign n56488 = ~n56483 & ~n56484;
  assign n56489 = n56482 & ~n61461;
  assign n56490 = ~n56479 & n56489;
  assign n56491 = ~pi241 & pi562;
  assign n56492 = pi242 & ~pi556;
  assign n56493 = ~n56491 & ~n56492;
  assign n56494 = pi241 & ~pi562;
  assign n56495 = pi240 & ~pi560;
  assign n56496 = ~n56494 & ~n56495;
  assign n56497 = n56493 & n56496;
  assign n56498 = ~pi246 & pi564;
  assign n56499 = ~pi248 & pi565;
  assign n56500 = ~n56498 & ~n56499;
  assign n56501 = pi248 & ~pi565;
  assign n56502 = ~pi242 & pi556;
  assign n56503 = ~n56501 & ~n56502;
  assign n56504 = n56500 & n56503;
  assign n56505 = n56497 & n56504;
  assign n56506 = n56490 & n56505;
  assign n56507 = ~n56476 & n56506;
  assign n56508 = ~pi242 & ~pi556;
  assign n56509 = pi242 & pi556;
  assign n56510 = ~n56508 & ~n56509;
  assign n56511 = ~n56499 & ~n56501;
  assign n56512 = ~n56479 & n56511;
  assign n56513 = pi241 & pi562;
  assign n56514 = ~pi241 & ~pi562;
  assign n56515 = ~n56513 & ~n56514;
  assign n56516 = ~pi246 & ~pi564;
  assign n56517 = pi246 & pi564;
  assign n56518 = ~n56516 & ~n56517;
  assign n56519 = pi240 & pi560;
  assign n56520 = ~pi240 & ~pi560;
  assign n56521 = ~n56519 & ~n56520;
  assign n56522 = ~n56518 & ~n56521;
  assign n56523 = ~n56515 & n56522;
  assign n56524 = n56512 & n56523;
  assign n56525 = ~n56476 & n56524;
  assign n56526 = ~pi249 & pi482;
  assign n56527 = pi249 & ~pi482;
  assign n56528 = ~n56498 & ~n56527;
  assign n56529 = ~n56526 & n56528;
  assign n56530 = ~n56515 & n56529;
  assign n56531 = ~n56475 & n56530;
  assign n56532 = ~n56476 & n56531;
  assign n56533 = ~n56481 & n56511;
  assign n56534 = ~n56521 & n56533;
  assign n56535 = n56532 & n56534;
  assign n56536 = ~n56475 & n56525;
  assign n56537 = ~n61461 & n61462;
  assign n56538 = ~n56510 & n56537;
  assign n56539 = ~n56475 & n56507;
  assign n56540 = ~n56474 & n61463;
  assign n56541 = ~pi244 & ~pi566;
  assign n56542 = pi244 & pi566;
  assign n56543 = ~n56541 & ~n56542;
  assign n56544 = n56540 & ~n56543;
  assign n56545 = pi568 & n56544;
  assign n56546 = pi245 & ~n56545;
  assign n56547 = ~pi531 & n61463;
  assign n56548 = n56459 & ~n56547;
  assign n56549 = pi531 & n61463;
  assign n56550 = n56457 & ~n56549;
  assign n56551 = ~n56451 & ~n56508;
  assign n56552 = pi569 & n61462;
  assign n56553 = pi569 & ~n56448;
  assign n56554 = n61462 & n56553;
  assign n56555 = ~n56448 & n56552;
  assign n56556 = n56486 & n61462;
  assign n56557 = ~n56449 & ~n56556;
  assign n56558 = ~n61464 & n56557;
  assign n56559 = ~pi489 & n56558;
  assign n56560 = pi489 & ~n56537;
  assign n56561 = ~pi556 & ~n56560;
  assign n56562 = ~n56559 & n56561;
  assign n56563 = ~n56551 & ~n56562;
  assign n56564 = ~n56453 & ~n56509;
  assign n56565 = pi489 & n56558;
  assign n56566 = ~pi489 & ~n56537;
  assign n56567 = pi556 & ~n56566;
  assign n56568 = ~n56565 & n56567;
  assign n56569 = ~n56564 & ~n56568;
  assign n56570 = ~n56563 & ~n56569;
  assign n56571 = ~pi549 & n56570;
  assign n56572 = pi549 & n61463;
  assign n56573 = ~pi235 & ~n56572;
  assign n56574 = ~n56571 & n56573;
  assign n56575 = ~n56457 & ~n56574;
  assign n56576 = ~pi531 & ~n56575;
  assign n56577 = pi549 & n56570;
  assign n56578 = ~pi549 & n61463;
  assign n56579 = pi235 & ~n56578;
  assign n56580 = ~n56577 & n56579;
  assign n56581 = ~n56459 & ~n56580;
  assign n56582 = pi531 & ~n56581;
  assign n56583 = ~n56576 & ~n56582;
  assign n56584 = ~n56548 & ~n56550;
  assign n56585 = ~pi486 & n61465;
  assign n56586 = pi486 & n56540;
  assign n56587 = ~pi244 & ~n56586;
  assign n56588 = ~n56585 & n56587;
  assign n56589 = ~n56462 & ~n56588;
  assign n56590 = ~pi566 & ~n56589;
  assign n56591 = pi486 & n61465;
  assign n56592 = ~pi486 & n56540;
  assign n56593 = pi244 & ~n56592;
  assign n56594 = ~n56591 & n56593;
  assign n56595 = ~n56464 & ~n56594;
  assign n56596 = pi566 & ~n56595;
  assign n56597 = ~n56590 & ~n56596;
  assign n56598 = ~pi568 & n56597;
  assign n56599 = pi568 & n56465;
  assign n56600 = ~pi245 & ~n56599;
  assign n56601 = ~n56598 & n56600;
  assign n56602 = ~n56546 & ~n56601;
  assign n56603 = ~pi580 & ~n56602;
  assign n56604 = ~pi568 & n56544;
  assign n56605 = ~pi245 & ~n56604;
  assign n56606 = pi568 & n56597;
  assign n56607 = ~pi568 & n56465;
  assign n56608 = pi245 & ~n56607;
  assign n56609 = ~n56606 & n56608;
  assign n56610 = ~n56605 & ~n56609;
  assign n56611 = pi580 & ~n56610;
  assign n56612 = ~n56603 & ~n56611;
  assign n56613 = ~pi552 & n56612;
  assign n56614 = ~n56546 & ~n56605;
  assign n56615 = pi552 & n56614;
  assign n56616 = ~pi247 & ~n56615;
  assign n56617 = ~n56613 & n56616;
  assign n56618 = ~n56471 & ~n56617;
  assign n56619 = ~pi532 & ~n56618;
  assign n56620 = ~pi552 & n56469;
  assign n56621 = ~pi247 & ~n56620;
  assign n56622 = pi552 & n56612;
  assign n56623 = ~pi552 & n56614;
  assign n56624 = pi247 & ~n56623;
  assign n56625 = ~n56622 & n56624;
  assign n56626 = ~n56621 & ~n56625;
  assign n56627 = pi532 & ~n56626;
  assign n56628 = ~n56619 & ~n56627;
  assign n56629 = ~pi238 & n56628;
  assign n56630 = ~pi577 & ~n56629;
  assign n56631 = ~n56471 & ~n56621;
  assign n56632 = pi238 & n56631;
  assign n56633 = ~pi247 & ~pi532;
  assign n56634 = pi247 & pi532;
  assign n56635 = ~n56633 & ~n56634;
  assign n56636 = n56614 & ~n56635;
  assign n56637 = ~pi238 & n56636;
  assign n56638 = pi577 & ~n56637;
  assign n56639 = ~n56632 & n56638;
  assign n56640 = ~pi498 & ~n56639;
  assign n56641 = ~n56630 & n56640;
  assign n56642 = pi238 & n56628;
  assign n56643 = pi577 & ~n56642;
  assign n56644 = ~pi238 & n56631;
  assign n56645 = pi238 & n56636;
  assign n56646 = ~pi577 & ~n56645;
  assign n56647 = ~n56644 & n56646;
  assign n56648 = pi498 & ~n56647;
  assign n56649 = ~n56643 & n56648;
  assign n56650 = ~n56641 & ~n56649;
  assign n56651 = ~pi233 & ~n56650;
  assign n56652 = ~pi237 & ~n56651;
  assign n56653 = ~n56389 & n56652;
  assign po750 = ~n56144 & ~n56653;
  assign n56655 = pi534 & ~n44913;
  assign n56656 = ~pi239 & n44913;
  assign po691 = ~n56655 & ~n56656;
  assign n56658 = pi535 & ~n44913;
  assign n56659 = pi240 & n44913;
  assign n56660 = ~n56658 & ~n56659;
  assign n56661 = pi536 & ~n44913;
  assign n56662 = pi246 & n44913;
  assign n56663 = ~n56661 & ~n56662;
  assign n56664 = pi537 & ~n44913;
  assign n56665 = pi248 & n44913;
  assign n56666 = ~n56664 & ~n56665;
  assign n56667 = pi538 & ~n44913;
  assign n56668 = pi249 & n44913;
  assign n56669 = ~n56667 & ~n56668;
  assign n56670 = pi539 & ~n44920;
  assign n56671 = pi242 & n44920;
  assign n56672 = ~n56670 & ~n56671;
  assign n56673 = pi540 & ~n44920;
  assign n56674 = pi235 & n44920;
  assign n56675 = ~n56673 & ~n56674;
  assign n56676 = pi541 & ~n44920;
  assign n56677 = pi244 & n44920;
  assign n56678 = ~n56676 & ~n56677;
  assign n56679 = pi542 & ~n44920;
  assign n56680 = pi240 & n44920;
  assign n56681 = ~n56679 & ~n56680;
  assign n56682 = pi543 & ~n44920;
  assign n56683 = pi238 & n44920;
  assign n56684 = ~n56682 & ~n56683;
  assign n56685 = pi544 & ~n44928;
  assign n56686 = n44923 & n55144;
  assign n56687 = n44928 & n55146;
  assign n56688 = pi544 & ~n56687;
  assign n56689 = ~pi544 & n44923;
  assign n56690 = n55144 & n56689;
  assign n56691 = ~n56688 & ~n56690;
  assign n56692 = ~n56685 & ~n56686;
  assign n56693 = pi545 & ~n44928;
  assign n56694 = pi245 & n44928;
  assign n56695 = ~n56693 & ~n56694;
  assign n56696 = pi546 & ~n44928;
  assign n56697 = pi246 & n44928;
  assign n56698 = ~n56696 & ~n56697;
  assign n56699 = pi547 & ~n44928;
  assign n56700 = pi247 & n44928;
  assign n56701 = ~n56699 & ~n56700;
  assign n56702 = pi548 & ~n44928;
  assign n56703 = pi248 & n44928;
  assign n56704 = ~n56702 & ~n56703;
  assign n56705 = pi549 & ~n44935;
  assign n56706 = pi235 & n44935;
  assign n56707 = ~n56705 & ~n56706;
  assign n56708 = pi550 & ~n44935;
  assign n56709 = ~pi239 & n44935;
  assign po707 = ~n56708 & ~n56709;
  assign n56711 = pi551 & ~n44935;
  assign n56712 = pi240 & n44935;
  assign n56713 = ~n56711 & ~n56712;
  assign n56714 = pi552 & ~n44935;
  assign n56715 = pi247 & n44935;
  assign n56716 = ~n56714 & ~n56715;
  assign n56717 = pi553 & ~n44935;
  assign n56718 = pi241 & n44935;
  assign n56719 = ~n56717 & ~n56718;
  assign n56720 = pi554 & ~n44935;
  assign n56721 = pi248 & n44935;
  assign n56722 = ~n56720 & ~n56721;
  assign n56723 = pi555 & ~n44935;
  assign n56724 = pi249 & n44935;
  assign n56725 = ~n56723 & ~n56724;
  assign n56726 = pi556 & ~n44799;
  assign n56727 = pi242 & n44799;
  assign n56728 = ~n56726 & ~n56727;
  assign n56729 = pi557 & ~n44913;
  assign n56730 = n44556 & n55144;
  assign n56731 = n44913 & n55146;
  assign n56732 = pi557 & ~n56731;
  assign n56733 = ~pi557 & n44556;
  assign n56734 = n55144 & n56733;
  assign n56735 = ~n56732 & ~n56734;
  assign n56736 = ~n56729 & ~n56730;
  assign n56737 = pi558 & ~n44913;
  assign n56738 = pi244 & n44913;
  assign n56739 = ~n56737 & ~n56738;
  assign n56740 = pi559 & ~n44783;
  assign n56741 = pi241 & n44783;
  assign n56742 = ~n56740 & ~n56741;
  assign n56743 = pi560 & ~n44799;
  assign n56744 = pi240 & n44799;
  assign n56745 = ~n56743 & ~n56744;
  assign n56746 = pi561 & ~n44791;
  assign n56747 = pi247 & n44791;
  assign n56748 = ~n56746 & ~n56747;
  assign n56749 = pi562 & ~n44799;
  assign n56750 = pi241 & n44799;
  assign n56751 = ~n56749 & ~n56750;
  assign n56752 = pi563 & ~n44935;
  assign n56753 = pi246 & n44935;
  assign n56754 = ~n56752 & ~n56753;
  assign n56755 = pi564 & ~n44799;
  assign n56756 = pi246 & n44799;
  assign n56757 = ~n56755 & ~n56756;
  assign n56758 = pi565 & ~n44799;
  assign n56759 = pi248 & n44799;
  assign n56760 = ~n56758 & ~n56759;
  assign n56761 = pi566 & ~n44799;
  assign n56762 = pi244 & n44799;
  assign n56763 = ~n56761 & ~n56762;
  assign n56764 = pi568 & ~n44799;
  assign n56765 = pi245 & n44799;
  assign n56766 = ~n56764 & ~n56765;
  assign n56767 = pi569 & ~n44799;
  assign n56768 = ~pi239 & n44799;
  assign po726 = ~n56767 & ~n56768;
  assign n56770 = pi570 & ~n44799;
  assign n56771 = n44794 & n55191;
  assign n56772 = n44799 & n55168;
  assign n56773 = pi570 & ~n56772;
  assign n56774 = ~pi570 & n44794;
  assign n56775 = n55191 & n56774;
  assign n56776 = ~n56773 & ~n56775;
  assign n56777 = ~n56770 & ~n56771;
  assign n56778 = pi571 & ~n44942;
  assign n56779 = pi241 & n44942;
  assign n56780 = ~n56778 & ~n56779;
  assign n56781 = pi572 & ~n44942;
  assign n56782 = pi244 & n44942;
  assign n56783 = ~n56781 & ~n56782;
  assign n56784 = pi573 & ~n44942;
  assign n56785 = pi242 & n44942;
  assign n56786 = ~n56784 & ~n56785;
  assign n56787 = pi574 & ~n44791;
  assign n56788 = pi241 & n44791;
  assign n56789 = ~n56787 & ~n56788;
  assign n56790 = pi575 & ~n44942;
  assign n56791 = pi235 & n44942;
  assign n56792 = ~n56790 & ~n56791;
  assign n56793 = pi576 & ~n44942;
  assign n56794 = pi248 & n44942;
  assign n56795 = ~n56793 & ~n56794;
  assign n56796 = pi577 & ~n44935;
  assign n56797 = pi238 & n44935;
  assign n56798 = ~n56796 & ~n56797;
  assign n56799 = pi578 & ~n44791;
  assign n56800 = pi249 & n44791;
  assign n56801 = ~n56799 & ~n56800;
  assign n56802 = pi579 & ~n44783;
  assign n56803 = pi249 & n44783;
  assign n56804 = ~n56802 & ~n56803;
  assign n56805 = pi580 & ~n44935;
  assign n56806 = pi245 & n44935;
  assign n56807 = ~n56805 & ~n56806;
  assign n56808 = pi581 & ~n44791;
  assign n56809 = pi235 & n44791;
  assign n56810 = ~n56808 & ~n56809;
  assign n56811 = pi582 & ~n44791;
  assign n56812 = pi240 & n44791;
  assign n56813 = ~n56811 & ~n56812;
  assign n56814 = pi584 & ~n44791;
  assign n56815 = pi245 & n44791;
  assign n56816 = ~n56814 & ~n56815;
  assign n56817 = pi585 & ~n44791;
  assign n56818 = pi244 & n44791;
  assign n56819 = ~n56817 & ~n56818;
  assign n56820 = pi586 & ~n44791;
  assign n56821 = pi242 & n44791;
  assign n56822 = ~n56820 & ~n56821;
  assign n56823 = ~pi882 & n58992;
  assign n56824 = pi947 & n56823;
  assign n56825 = pi598 & ~n56824;
  assign n56826 = pi740 & pi780;
  assign n56827 = n2778 & n56826;
  assign n56828 = ~n56825 & ~n56827;
  assign n56829 = pi907 & n56823;
  assign n56830 = ~pi615 & ~n56829;
  assign n56831 = pi779 & pi797;
  assign n56832 = n2781 & n56831;
  assign n56833 = ~n56830 & ~n56832;
  assign n56834 = pi832 & ~pi973;
  assign n56835 = ~pi1054 & pi1066;
  assign n56836 = pi1088 & n56835;
  assign n56837 = n56834 & n56836;
  assign po954 = ~pi953 & n56837;
  assign n56839 = ~pi1116 & po954;
  assign n56840 = ~pi625 & ~po954;
  assign n56841 = ~pi962 & ~n56840;
  assign n56842 = ~pi962 & ~n56839;
  assign n56843 = ~n56840 & n56842;
  assign n56844 = ~n56839 & n56841;
  assign n56845 = ~pi1117 & po954;
  assign n56846 = ~pi627 & ~po954;
  assign n56847 = ~pi962 & ~n56846;
  assign n56848 = ~pi962 & ~n56845;
  assign n56849 = ~n56846 & n56848;
  assign n56850 = ~n56845 & n56847;
  assign n56851 = ~pi1119 & po954;
  assign n56852 = ~pi628 & ~po954;
  assign n56853 = ~pi962 & ~n56852;
  assign n56854 = ~pi962 & ~n56851;
  assign n56855 = ~n56852 & n56854;
  assign n56856 = ~n56851 & n56853;
  assign n56857 = ~pi980 & pi1038;
  assign n56858 = pi1060 & n56857;
  assign n56859 = pi832 & ~pi1061;
  assign n56860 = pi952 & n56859;
  assign n56861 = pi952 & ~pi1061;
  assign n56862 = n56858 & n56861;
  assign n56863 = pi832 & n56862;
  assign n56864 = n56858 & n56860;
  assign n56865 = ~pi1119 & po897;
  assign n56866 = ~pi629 & ~po897;
  assign n56867 = ~pi966 & ~n56866;
  assign n56868 = ~pi966 & ~n56865;
  assign n56869 = ~n56866 & n56868;
  assign n56870 = ~n56865 & n56867;
  assign n56871 = ~pi1120 & po897;
  assign n56872 = ~pi630 & ~po897;
  assign n56873 = ~pi966 & ~n56872;
  assign n56874 = ~pi966 & ~n56871;
  assign n56875 = ~n56872 & n56874;
  assign n56876 = ~n56871 & n56873;
  assign n56877 = pi631 & ~po954;
  assign n56878 = ~pi1113 & po954;
  assign n56879 = ~pi962 & ~n56878;
  assign n56880 = ~pi962 & ~n56877;
  assign n56881 = ~n56878 & n56880;
  assign n56882 = ~n56877 & n56879;
  assign n56883 = pi632 & ~po954;
  assign n56884 = ~pi1115 & po954;
  assign n56885 = ~pi962 & ~n56884;
  assign n56886 = ~pi962 & ~n56883;
  assign n56887 = ~n56884 & n56886;
  assign n56888 = ~n56883 & n56885;
  assign n56889 = ~pi1110 & po897;
  assign n56890 = ~pi633 & ~po897;
  assign n56891 = ~pi966 & ~n56890;
  assign n56892 = ~pi966 & ~n56889;
  assign n56893 = ~n56890 & n56892;
  assign n56894 = ~n56889 & n56891;
  assign n56895 = ~pi1110 & po954;
  assign n56896 = ~pi634 & ~po954;
  assign n56897 = ~pi962 & ~n56896;
  assign n56898 = ~pi962 & ~n56895;
  assign n56899 = ~n56896 & n56898;
  assign n56900 = ~n56895 & n56897;
  assign n56901 = pi635 & ~po954;
  assign n56902 = ~pi1112 & po954;
  assign n56903 = ~pi962 & ~n56902;
  assign n56904 = ~pi962 & ~n56901;
  assign n56905 = ~n56902 & n56904;
  assign n56906 = ~n56901 & n56903;
  assign n56907 = ~pi1127 & po897;
  assign n56908 = ~pi636 & ~po897;
  assign n56909 = ~pi966 & ~n56908;
  assign n56910 = ~pi966 & ~n56907;
  assign n56911 = ~n56908 & n56910;
  assign n56912 = ~n56907 & n56909;
  assign n56913 = ~pi1105 & po954;
  assign n56914 = ~pi637 & ~po954;
  assign n56915 = ~pi962 & ~n56914;
  assign n56916 = ~pi962 & ~n56913;
  assign n56917 = ~n56914 & n56916;
  assign n56918 = ~n56913 & n56915;
  assign n56919 = ~pi1107 & po954;
  assign n56920 = ~pi638 & ~po954;
  assign n56921 = ~pi962 & ~n56920;
  assign n56922 = ~pi962 & ~n56919;
  assign n56923 = ~n56920 & n56922;
  assign n56924 = ~n56919 & n56921;
  assign n56925 = ~pi1109 & po954;
  assign n56926 = ~pi639 & ~po954;
  assign n56927 = ~pi962 & ~n56926;
  assign n56928 = ~pi962 & ~n56925;
  assign n56929 = ~n56926 & n56928;
  assign n56930 = ~n56925 & n56927;
  assign n56931 = ~pi1128 & po897;
  assign n56932 = ~pi640 & ~po897;
  assign n56933 = ~pi966 & ~n56932;
  assign n56934 = ~pi966 & ~n56931;
  assign n56935 = ~n56932 & n56934;
  assign n56936 = ~n56931 & n56933;
  assign n56937 = ~pi1121 & po954;
  assign n56938 = ~pi641 & ~po954;
  assign n56939 = ~pi962 & ~n56938;
  assign n56940 = ~pi962 & ~n56937;
  assign n56941 = ~n56938 & n56940;
  assign n56942 = ~n56937 & n56939;
  assign n56943 = ~pi1104 & po954;
  assign n56944 = ~pi643 & ~po954;
  assign n56945 = ~pi962 & ~n56944;
  assign n56946 = ~pi962 & ~n56943;
  assign n56947 = ~n56944 & n56946;
  assign n56948 = ~n56943 & n56945;
  assign n56949 = ~pi1123 & po897;
  assign n56950 = ~pi644 & ~po897;
  assign n56951 = ~pi966 & ~n56950;
  assign n56952 = ~pi966 & ~n56949;
  assign n56953 = ~n56950 & n56952;
  assign n56954 = ~n56949 & n56951;
  assign n56955 = ~pi1125 & po897;
  assign n56956 = ~pi645 & ~po897;
  assign n56957 = ~pi966 & ~n56956;
  assign n56958 = ~pi966 & ~n56955;
  assign n56959 = ~n56956 & n56958;
  assign n56960 = ~n56955 & n56957;
  assign n56961 = pi646 & ~po954;
  assign n56962 = ~pi1114 & po954;
  assign n56963 = ~pi962 & ~n56962;
  assign n56964 = ~pi962 & ~n56961;
  assign n56965 = ~n56962 & n56964;
  assign n56966 = ~n56961 & n56963;
  assign n56967 = ~pi1120 & po954;
  assign n56968 = ~pi647 & ~po954;
  assign n56969 = ~pi962 & ~n56968;
  assign n56970 = ~pi962 & ~n56967;
  assign n56971 = ~n56968 & n56970;
  assign n56972 = ~n56967 & n56969;
  assign n56973 = ~pi1122 & po954;
  assign n56974 = ~pi648 & ~po954;
  assign n56975 = ~pi962 & ~n56974;
  assign n56976 = ~pi962 & ~n56973;
  assign n56977 = ~n56974 & n56976;
  assign n56978 = ~n56973 & n56975;
  assign n56979 = pi649 & ~po954;
  assign n56980 = ~pi1126 & po954;
  assign n56981 = ~pi962 & ~n56980;
  assign n56982 = ~pi962 & ~n56979;
  assign n56983 = ~n56980 & n56982;
  assign n56984 = ~n56979 & n56981;
  assign n56985 = pi650 & ~po954;
  assign n56986 = ~pi1127 & po954;
  assign n56987 = ~pi962 & ~n56986;
  assign n56988 = ~pi962 & ~n56985;
  assign n56989 = ~n56986 & n56988;
  assign n56990 = ~n56985 & n56987;
  assign n56991 = ~pi1130 & po897;
  assign n56992 = ~pi651 & ~po897;
  assign n56993 = ~pi966 & ~n56992;
  assign n56994 = ~pi966 & ~n56991;
  assign n56995 = ~n56992 & n56994;
  assign n56996 = ~n56991 & n56993;
  assign n56997 = ~pi1131 & po897;
  assign n56998 = ~pi652 & ~po897;
  assign n56999 = ~pi966 & ~n56998;
  assign n57000 = ~pi966 & ~n56997;
  assign n57001 = ~n56998 & n57000;
  assign n57002 = ~n56997 & n56999;
  assign n57003 = ~pi1129 & po897;
  assign n57004 = ~pi653 & ~po897;
  assign n57005 = ~pi966 & ~n57004;
  assign n57006 = ~pi966 & ~n57003;
  assign n57007 = ~n57004 & n57006;
  assign n57008 = ~n57003 & n57005;
  assign n57009 = pi654 & ~po954;
  assign n57010 = ~pi1130 & po954;
  assign n57011 = ~pi962 & ~n57010;
  assign n57012 = ~pi962 & ~n57009;
  assign n57013 = ~n57010 & n57012;
  assign n57014 = ~n57009 & n57011;
  assign n57015 = pi655 & ~po954;
  assign n57016 = ~pi1124 & po954;
  assign n57017 = ~pi962 & ~n57016;
  assign n57018 = ~pi962 & ~n57015;
  assign n57019 = ~n57016 & n57018;
  assign n57020 = ~n57015 & n57017;
  assign n57021 = ~pi1126 & po897;
  assign n57022 = ~pi656 & ~po897;
  assign n57023 = ~pi966 & ~n57022;
  assign n57024 = ~pi966 & ~n57021;
  assign n57025 = ~n57022 & n57024;
  assign n57026 = ~n57021 & n57023;
  assign n57027 = pi657 & ~po954;
  assign n57028 = ~pi1131 & po954;
  assign n57029 = ~pi962 & ~n57028;
  assign n57030 = ~pi962 & ~n57027;
  assign n57031 = ~n57028 & n57030;
  assign n57032 = ~n57027 & n57029;
  assign n57033 = ~pi1124 & po897;
  assign n57034 = ~pi658 & ~po897;
  assign n57035 = ~pi966 & ~n57034;
  assign n57036 = ~pi966 & ~n57033;
  assign n57037 = ~n57034 & n57036;
  assign n57038 = ~n57033 & n57035;
  assign n57039 = ~pi1118 & po954;
  assign n57040 = ~pi660 & ~po954;
  assign n57041 = ~pi962 & ~n57040;
  assign n57042 = ~pi962 & ~n57039;
  assign n57043 = ~n57040 & n57042;
  assign n57044 = ~n57039 & n57041;
  assign n57045 = ~pi1101 & po954;
  assign n57046 = ~pi661 & ~po954;
  assign n57047 = ~pi962 & ~n57046;
  assign n57048 = ~pi962 & ~n57045;
  assign n57049 = ~n57046 & n57048;
  assign n57050 = ~n57045 & n57047;
  assign n57051 = ~pi1102 & po954;
  assign n57052 = ~pi662 & ~po954;
  assign n57053 = ~pi962 & ~n57052;
  assign n57054 = ~pi962 & ~n57051;
  assign n57055 = ~n57052 & n57054;
  assign n57056 = ~n57051 & n57053;
  assign n57057 = ~pi1108 & po954;
  assign n57058 = ~pi665 & ~po954;
  assign n57059 = ~pi962 & ~n57058;
  assign n57060 = ~pi962 & ~n57057;
  assign n57061 = ~n57058 & n57060;
  assign n57062 = ~n57057 & n57059;
  assign n57063 = pi669 & ~po954;
  assign n57064 = ~pi1125 & po954;
  assign n57065 = ~pi962 & ~n57064;
  assign n57066 = ~pi962 & ~n57063;
  assign n57067 = ~n57064 & n57066;
  assign n57068 = ~n57063 & n57065;
  assign n57069 = ~pi1100 & po954;
  assign n57070 = ~pi680 & ~po954;
  assign n57071 = ~pi962 & ~n57070;
  assign n57072 = ~pi962 & ~n57069;
  assign n57073 = ~n57070 & n57072;
  assign n57074 = ~n57069 & n57071;
  assign n57075 = ~pi1103 & po954;
  assign n57076 = ~pi681 & ~po954;
  assign n57077 = ~pi962 & ~n57076;
  assign n57078 = ~pi962 & ~n57075;
  assign n57079 = ~n57076 & n57078;
  assign n57080 = ~n57075 & n57077;
  assign po980 = pi953 & n56837;
  assign n57082 = pi684 & ~po980;
  assign n57083 = ~pi1130 & po980;
  assign n57084 = ~pi962 & ~n57083;
  assign n57085 = ~pi962 & ~n57082;
  assign n57086 = ~n57083 & n57085;
  assign n57087 = ~n57082 & n57084;
  assign n57088 = pi686 & ~po980;
  assign n57089 = ~pi1113 & po980;
  assign n57090 = ~pi962 & ~n57089;
  assign n57091 = ~pi962 & ~n57088;
  assign n57092 = ~n57089 & n57091;
  assign n57093 = ~n57088 & n57090;
  assign n57094 = ~pi1127 & po980;
  assign n57095 = ~pi687 & ~po980;
  assign n57096 = ~pi962 & ~n57095;
  assign n57097 = ~pi962 & ~n57094;
  assign n57098 = ~n57095 & n57097;
  assign n57099 = ~n57094 & n57096;
  assign n57100 = pi688 & ~po980;
  assign n57101 = ~pi1115 & po980;
  assign n57102 = ~pi962 & ~n57101;
  assign n57103 = ~pi962 & ~n57100;
  assign n57104 = ~n57101 & n57103;
  assign n57105 = ~n57100 & n57102;
  assign n57106 = ~pi1108 & po980;
  assign n57107 = ~pi690 & ~po980;
  assign n57108 = ~pi962 & ~n57107;
  assign n57109 = ~pi962 & ~n57106;
  assign n57110 = ~n57107 & n57109;
  assign n57111 = ~n57106 & n57108;
  assign n57112 = ~pi1107 & po980;
  assign n57113 = ~pi691 & ~po980;
  assign n57114 = ~pi962 & ~n57113;
  assign n57115 = ~pi962 & ~n57112;
  assign n57116 = ~n57113 & n57115;
  assign n57117 = ~n57112 & n57114;
  assign n57118 = pi693 & ~po954;
  assign n57119 = ~pi1129 & po954;
  assign n57120 = ~pi962 & ~n57119;
  assign n57121 = ~pi962 & ~n57118;
  assign n57122 = ~n57119 & n57121;
  assign n57123 = ~n57118 & n57120;
  assign n57124 = pi694 & ~po980;
  assign n57125 = ~pi1128 & po980;
  assign n57126 = ~pi962 & ~n57125;
  assign n57127 = ~pi962 & ~n57124;
  assign n57128 = ~n57125 & n57127;
  assign n57129 = ~n57124 & n57126;
  assign n57130 = pi695 & ~po954;
  assign n57131 = ~pi1111 & po954;
  assign n57132 = ~pi962 & ~n57131;
  assign n57133 = ~pi962 & ~n57130;
  assign n57134 = ~n57131 & n57133;
  assign n57135 = ~n57130 & n57132;
  assign n57136 = ~pi1100 & po980;
  assign n57137 = ~pi696 & ~po980;
  assign n57138 = ~pi962 & ~n57137;
  assign n57139 = ~pi962 & ~n57136;
  assign n57140 = ~n57137 & n57139;
  assign n57141 = ~n57136 & n57138;
  assign n57142 = pi697 & ~po980;
  assign n57143 = ~pi1129 & po980;
  assign n57144 = ~pi962 & ~n57143;
  assign n57145 = ~pi962 & ~n57142;
  assign n57146 = ~n57143 & n57145;
  assign n57147 = ~n57142 & n57144;
  assign n57148 = pi698 & ~po980;
  assign n57149 = ~pi1116 & po980;
  assign n57150 = ~pi962 & ~n57149;
  assign n57151 = ~pi962 & ~n57148;
  assign n57152 = ~n57149 & n57151;
  assign n57153 = ~n57148 & n57150;
  assign n57154 = ~pi1103 & po980;
  assign n57155 = ~pi699 & ~po980;
  assign n57156 = ~pi962 & ~n57155;
  assign n57157 = ~pi962 & ~n57154;
  assign n57158 = ~n57155 & n57157;
  assign n57159 = ~n57154 & n57156;
  assign n57160 = ~pi1110 & po980;
  assign n57161 = ~pi700 & ~po980;
  assign n57162 = ~pi962 & ~n57161;
  assign n57163 = ~pi962 & ~n57160;
  assign n57164 = ~n57161 & n57163;
  assign n57165 = ~n57160 & n57162;
  assign n57166 = pi701 & ~po980;
  assign n57167 = ~pi1123 & po980;
  assign n57168 = ~pi962 & ~n57167;
  assign n57169 = ~pi962 & ~n57166;
  assign n57170 = ~n57167 & n57169;
  assign n57171 = ~n57166 & n57168;
  assign n57172 = pi702 & ~po980;
  assign n57173 = ~pi1117 & po980;
  assign n57174 = ~pi962 & ~n57173;
  assign n57175 = ~pi962 & ~n57172;
  assign n57176 = ~n57173 & n57175;
  assign n57177 = ~n57172 & n57174;
  assign n57178 = ~pi1124 & po980;
  assign n57179 = ~pi703 & ~po980;
  assign n57180 = ~pi962 & ~n57179;
  assign n57181 = ~pi962 & ~n57178;
  assign n57182 = ~n57179 & n57181;
  assign n57183 = ~n57178 & n57180;
  assign n57184 = pi704 & ~po980;
  assign n57185 = ~pi1112 & po980;
  assign n57186 = ~pi962 & ~n57185;
  assign n57187 = ~pi962 & ~n57184;
  assign n57188 = ~n57185 & n57187;
  assign n57189 = ~n57184 & n57186;
  assign n57190 = ~pi1125 & po980;
  assign n57191 = ~pi705 & ~po980;
  assign n57192 = ~pi962 & ~n57191;
  assign n57193 = ~pi962 & ~n57190;
  assign n57194 = ~n57191 & n57193;
  assign n57195 = ~n57190 & n57192;
  assign n57196 = ~pi1105 & po980;
  assign n57197 = ~pi706 & ~po980;
  assign n57198 = ~pi962 & ~n57197;
  assign n57199 = ~pi962 & ~n57196;
  assign n57200 = ~n57197 & n57199;
  assign n57201 = ~n57196 & n57198;
  assign n57202 = pi709 & ~po980;
  assign n57203 = ~pi1118 & po980;
  assign n57204 = ~pi962 & ~n57203;
  assign n57205 = ~pi962 & ~n57202;
  assign n57206 = ~n57203 & n57205;
  assign n57207 = ~n57202 & n57204;
  assign n57208 = ~pi1106 & po954;
  assign n57209 = ~pi710 & ~po954;
  assign n57210 = ~pi962 & ~n57209;
  assign n57211 = ~pi962 & ~n57208;
  assign n57212 = ~n57209 & n57211;
  assign n57213 = ~n57208 & n57210;
  assign n57214 = ~pi1123 & po954;
  assign n57215 = ~pi715 & ~po954;
  assign n57216 = ~pi962 & ~n57215;
  assign n57217 = ~pi962 & ~n57214;
  assign n57218 = ~n57215 & n57217;
  assign n57219 = ~n57214 & n57216;
  assign n57220 = pi723 & ~po980;
  assign n57221 = ~pi1111 & po980;
  assign n57222 = ~pi962 & ~n57221;
  assign n57223 = ~pi962 & ~n57220;
  assign n57224 = ~n57221 & n57223;
  assign n57225 = ~n57220 & n57222;
  assign n57226 = pi724 & ~po980;
  assign n57227 = ~pi1114 & po980;
  assign n57228 = ~pi962 & ~n57227;
  assign n57229 = ~pi962 & ~n57226;
  assign n57230 = ~n57227 & n57229;
  assign n57231 = ~n57226 & n57228;
  assign n57232 = pi725 & ~po980;
  assign n57233 = ~pi1120 & po980;
  assign n57234 = ~pi962 & ~n57233;
  assign n57235 = ~pi962 & ~n57232;
  assign n57236 = ~n57233 & n57235;
  assign n57237 = ~n57232 & n57234;
  assign n57238 = ~pi1126 & po980;
  assign n57239 = ~pi726 & ~po980;
  assign n57240 = ~pi962 & ~n57239;
  assign n57241 = ~pi962 & ~n57238;
  assign n57242 = ~n57239 & n57241;
  assign n57243 = ~n57238 & n57240;
  assign n57244 = ~pi1102 & po980;
  assign n57245 = ~pi727 & ~po980;
  assign n57246 = ~pi962 & ~n57245;
  assign n57247 = ~pi962 & ~n57244;
  assign n57248 = ~n57245 & n57247;
  assign n57249 = ~n57244 & n57246;
  assign n57250 = pi728 & ~po980;
  assign n57251 = ~pi1131 & po980;
  assign n57252 = ~pi962 & ~n57251;
  assign n57253 = ~pi962 & ~n57250;
  assign n57254 = ~n57251 & n57253;
  assign n57255 = ~n57250 & n57252;
  assign n57256 = ~pi1104 & po980;
  assign n57257 = ~pi729 & ~po980;
  assign n57258 = ~pi962 & ~n57257;
  assign n57259 = ~pi962 & ~n57256;
  assign n57260 = ~n57257 & n57259;
  assign n57261 = ~n57256 & n57258;
  assign n57262 = ~pi1106 & po980;
  assign n57263 = ~pi730 & ~po980;
  assign n57264 = ~pi962 & ~n57263;
  assign n57265 = ~pi962 & ~n57262;
  assign n57266 = ~n57263 & n57265;
  assign n57267 = ~n57262 & n57264;
  assign n57268 = pi732 & ~po954;
  assign n57269 = ~pi1128 & po954;
  assign n57270 = ~pi962 & ~n57269;
  assign n57271 = ~pi962 & ~n57268;
  assign n57272 = ~n57269 & n57271;
  assign n57273 = ~n57268 & n57270;
  assign n57274 = pi734 & ~po980;
  assign n57275 = ~pi1119 & po980;
  assign n57276 = ~pi962 & ~n57275;
  assign n57277 = ~pi962 & ~n57274;
  assign n57278 = ~n57275 & n57277;
  assign n57279 = ~n57274 & n57276;
  assign n57280 = ~pi1109 & po980;
  assign n57281 = ~pi735 & ~po980;
  assign n57282 = ~pi962 & ~n57281;
  assign n57283 = ~pi962 & ~n57280;
  assign n57284 = ~n57281 & n57283;
  assign n57285 = ~n57280 & n57282;
  assign n57286 = ~pi1101 & po980;
  assign n57287 = ~pi736 & ~po980;
  assign n57288 = ~pi962 & ~n57287;
  assign n57289 = ~pi962 & ~n57286;
  assign n57290 = ~n57287 & n57289;
  assign n57291 = ~n57286 & n57288;
  assign n57292 = pi737 & ~po980;
  assign n57293 = ~pi1122 & po980;
  assign n57294 = ~pi962 & ~n57293;
  assign n57295 = ~pi962 & ~n57292;
  assign n57296 = ~n57293 & n57295;
  assign n57297 = ~n57292 & n57294;
  assign n57298 = pi738 & ~po980;
  assign n57299 = ~pi1121 & po980;
  assign n57300 = ~pi962 & ~n57299;
  assign n57301 = ~pi962 & ~n57298;
  assign n57302 = ~n57299 & n57301;
  assign n57303 = ~n57298 & n57300;
  assign n57304 = ~pi952 & n56859;
  assign n57305 = ~pi952 & ~pi1061;
  assign n57306 = n56858 & n57305;
  assign n57307 = pi832 & n57306;
  assign n57308 = n56858 & n57304;
  assign n57309 = pi739 & ~po988;
  assign n57310 = pi1108 & po988;
  assign n57311 = ~pi966 & ~n57310;
  assign n57312 = ~pi966 & ~n57309;
  assign n57313 = ~n57310 & n57312;
  assign n57314 = ~n57309 & n57311;
  assign n57315 = pi1114 & po988;
  assign n57316 = ~pi741 & ~po988;
  assign n57317 = ~pi966 & ~n57316;
  assign n57318 = ~pi966 & ~n57315;
  assign n57319 = ~n57316 & n57318;
  assign n57320 = ~n57315 & n57317;
  assign n57321 = pi1112 & po988;
  assign n57322 = ~pi742 & ~po988;
  assign n57323 = ~pi966 & ~n57322;
  assign n57324 = ~pi966 & ~n57321;
  assign n57325 = ~n57322 & n57324;
  assign n57326 = ~n57321 & n57323;
  assign n57327 = pi743 & ~po988;
  assign n57328 = pi1109 & po988;
  assign n57329 = ~pi966 & ~n57328;
  assign n57330 = ~pi966 & ~n57327;
  assign n57331 = ~n57328 & n57330;
  assign n57332 = ~n57327 & n57329;
  assign n57333 = pi1131 & po988;
  assign n57334 = ~pi744 & ~po988;
  assign n57335 = ~pi966 & ~n57334;
  assign n57336 = ~pi966 & ~n57333;
  assign n57337 = ~n57334 & n57336;
  assign n57338 = ~n57333 & n57335;
  assign n57339 = pi1111 & po988;
  assign n57340 = ~pi745 & ~po988;
  assign n57341 = ~pi966 & ~n57340;
  assign n57342 = ~pi966 & ~n57339;
  assign n57343 = ~n57340 & n57342;
  assign n57344 = ~n57339 & n57341;
  assign n57345 = pi746 & ~po988;
  assign n57346 = pi1104 & po988;
  assign n57347 = ~pi966 & ~n57346;
  assign n57348 = ~pi966 & ~n57345;
  assign n57349 = ~n57346 & n57348;
  assign n57350 = ~n57345 & n57347;
  assign n57351 = pi748 & ~po988;
  assign n57352 = pi1106 & po988;
  assign n57353 = ~pi966 & ~n57352;
  assign n57354 = ~pi966 & ~n57351;
  assign n57355 = ~n57352 & n57354;
  assign n57356 = ~n57351 & n57353;
  assign n57357 = pi749 & ~po988;
  assign n57358 = pi1105 & po988;
  assign n57359 = ~pi966 & ~n57358;
  assign n57360 = ~pi966 & ~n57357;
  assign n57361 = ~n57358 & n57360;
  assign n57362 = ~n57357 & n57359;
  assign n57363 = pi1130 & po988;
  assign n57364 = ~pi750 & ~po988;
  assign n57365 = ~pi966 & ~n57364;
  assign n57366 = ~pi966 & ~n57363;
  assign n57367 = ~n57364 & n57366;
  assign n57368 = ~n57363 & n57365;
  assign n57369 = pi1123 & po988;
  assign n57370 = ~pi751 & ~po988;
  assign n57371 = ~pi966 & ~n57370;
  assign n57372 = ~pi966 & ~n57369;
  assign n57373 = ~n57370 & n57372;
  assign n57374 = ~n57369 & n57371;
  assign n57375 = pi1124 & po988;
  assign n57376 = ~pi752 & ~po988;
  assign n57377 = ~pi966 & ~n57376;
  assign n57378 = ~pi966 & ~n57375;
  assign n57379 = ~n57376 & n57378;
  assign n57380 = ~n57375 & n57377;
  assign n57381 = pi123 & n35583;
  assign n57382 = pi1131 & ~n57381;
  assign n57383 = pi1127 & ~n57381;
  assign n57384 = ~n57382 & ~n57383;
  assign n57385 = ~pi825 & n57381;
  assign n57386 = n57384 & ~n57385;
  assign n57387 = pi1131 & n57383;
  assign n57388 = ~n57386 & ~n57387;
  assign n57389 = pi1125 & ~pi1126;
  assign n57390 = ~pi1125 & pi1126;
  assign n57391 = ~pi1125 & ~pi1126;
  assign n57392 = pi1125 & pi1126;
  assign n57393 = ~n57391 & ~n57392;
  assign n57394 = ~n57389 & ~n57390;
  assign n57395 = ~pi1128 & ~pi1129;
  assign n57396 = pi1128 & pi1129;
  assign n57397 = pi1128 & ~pi1129;
  assign n57398 = ~pi1128 & pi1129;
  assign n57399 = ~n57397 & ~n57398;
  assign n57400 = ~n57395 & ~n57396;
  assign n57401 = ~pi1124 & ~pi1130;
  assign n57402 = pi1124 & pi1130;
  assign n57403 = pi1124 & ~pi1130;
  assign n57404 = ~pi1124 & pi1130;
  assign n57405 = ~n57403 & ~n57404;
  assign n57406 = ~n57401 & ~n57402;
  assign n57407 = ~n61560 & n61561;
  assign n57408 = n61560 & ~n61561;
  assign n57409 = ~n57407 & ~n57408;
  assign n57410 = ~n61559 & n57409;
  assign n57411 = n61559 & ~n57409;
  assign n57412 = ~n61559 & ~n61560;
  assign n57413 = n61559 & n61560;
  assign n57414 = ~n57412 & ~n57413;
  assign n57415 = n61561 & n57414;
  assign n57416 = ~n61561 & ~n57414;
  assign n57417 = ~n57415 & ~n57416;
  assign n57418 = ~n61559 & ~n61561;
  assign n57419 = n61559 & n61561;
  assign n57420 = ~n57418 & ~n57419;
  assign n57421 = n61560 & n57420;
  assign n57422 = ~n61560 & ~n57420;
  assign n57423 = ~n57421 & ~n57422;
  assign n57424 = ~n57410 & ~n57411;
  assign n57425 = ~n57388 & ~n61562;
  assign n57426 = pi825 & n57381;
  assign n57427 = n57384 & ~n57426;
  assign n57428 = ~n57387 & n61562;
  assign n57429 = ~n57427 & n57428;
  assign po982 = ~n57425 & ~n57429;
  assign n57431 = pi1123 & ~n57381;
  assign n57432 = pi1122 & ~n57381;
  assign n57433 = ~n57431 & ~n57432;
  assign n57434 = ~pi826 & n57381;
  assign n57435 = n57433 & ~n57434;
  assign n57436 = pi1123 & n57432;
  assign n57437 = ~n57435 & ~n57436;
  assign n57438 = pi1116 & ~pi1117;
  assign n57439 = ~pi1116 & pi1117;
  assign n57440 = ~pi1116 & ~pi1117;
  assign n57441 = pi1116 & pi1117;
  assign n57442 = ~n57440 & ~n57441;
  assign n57443 = ~n57438 & ~n57439;
  assign n57444 = ~pi1120 & ~pi1121;
  assign n57445 = pi1120 & pi1121;
  assign n57446 = pi1120 & ~pi1121;
  assign n57447 = ~pi1120 & pi1121;
  assign n57448 = ~n57446 & ~n57447;
  assign n57449 = ~n57444 & ~n57445;
  assign n57450 = ~pi1118 & ~pi1119;
  assign n57451 = pi1118 & pi1119;
  assign n57452 = pi1118 & ~pi1119;
  assign n57453 = ~pi1118 & pi1119;
  assign n57454 = ~n57452 & ~n57453;
  assign n57455 = ~n57450 & ~n57451;
  assign n57456 = ~n61564 & n61565;
  assign n57457 = n61564 & ~n61565;
  assign n57458 = ~n57456 & ~n57457;
  assign n57459 = ~n61563 & n57458;
  assign n57460 = n61563 & ~n57458;
  assign n57461 = ~n61563 & ~n61564;
  assign n57462 = n61563 & n61564;
  assign n57463 = ~n57461 & ~n57462;
  assign n57464 = n61565 & n57463;
  assign n57465 = ~n61565 & ~n57463;
  assign n57466 = ~n57464 & ~n57465;
  assign n57467 = ~n61563 & ~n61565;
  assign n57468 = n61563 & n61565;
  assign n57469 = ~n57467 & ~n57468;
  assign n57470 = n61564 & n57469;
  assign n57471 = ~n61564 & ~n57469;
  assign n57472 = ~n57470 & ~n57471;
  assign n57473 = ~n57459 & ~n57460;
  assign n57474 = ~n57437 & ~n61566;
  assign n57475 = pi826 & n57381;
  assign n57476 = n57433 & ~n57475;
  assign n57477 = ~n57436 & n61566;
  assign n57478 = ~n57476 & n57477;
  assign po983 = ~n57474 & ~n57478;
  assign n57480 = pi1100 & ~n57381;
  assign n57481 = pi1107 & ~n57381;
  assign n57482 = ~n57480 & ~n57481;
  assign n57483 = ~pi827 & n57381;
  assign n57484 = n57482 & ~n57483;
  assign n57485 = pi1100 & n57481;
  assign n57486 = ~n57484 & ~n57485;
  assign n57487 = pi1104 & ~pi1106;
  assign n57488 = ~pi1104 & pi1106;
  assign n57489 = ~pi1104 & ~pi1106;
  assign n57490 = pi1104 & pi1106;
  assign n57491 = ~n57489 & ~n57490;
  assign n57492 = ~n57487 & ~n57488;
  assign n57493 = ~pi1101 & ~pi1102;
  assign n57494 = pi1101 & pi1102;
  assign n57495 = pi1101 & ~pi1102;
  assign n57496 = ~pi1101 & pi1102;
  assign n57497 = ~n57495 & ~n57496;
  assign n57498 = ~n57493 & ~n57494;
  assign n57499 = ~pi1103 & ~pi1105;
  assign n57500 = pi1103 & pi1105;
  assign n57501 = pi1103 & ~pi1105;
  assign n57502 = ~pi1103 & pi1105;
  assign n57503 = ~n57501 & ~n57502;
  assign n57504 = ~n57499 & ~n57500;
  assign n57505 = ~n61568 & n61569;
  assign n57506 = n61568 & ~n61569;
  assign n57507 = ~n57505 & ~n57506;
  assign n57508 = ~n61567 & n57507;
  assign n57509 = n61567 & ~n57507;
  assign n57510 = ~n61567 & ~n61568;
  assign n57511 = n61567 & n61568;
  assign n57512 = ~n57510 & ~n57511;
  assign n57513 = n61569 & n57512;
  assign n57514 = ~n61569 & ~n57512;
  assign n57515 = ~n57513 & ~n57514;
  assign n57516 = ~n61567 & ~n61569;
  assign n57517 = n61567 & n61569;
  assign n57518 = ~n57516 & ~n57517;
  assign n57519 = n61568 & n57518;
  assign n57520 = ~n61568 & ~n57518;
  assign n57521 = ~n57519 & ~n57520;
  assign n57522 = ~n57508 & ~n57509;
  assign n57523 = ~n57486 & ~n61570;
  assign n57524 = pi827 & n57381;
  assign n57525 = n57482 & ~n57524;
  assign n57526 = ~n57485 & n61570;
  assign n57527 = ~n57525 & n57526;
  assign po984 = ~n57523 & ~n57527;
  assign n57529 = pi1115 & ~n57381;
  assign n57530 = pi1114 & ~n57381;
  assign n57531 = ~n57529 & ~n57530;
  assign n57532 = ~pi828 & n57381;
  assign n57533 = n57531 & ~n57532;
  assign n57534 = pi1115 & n57530;
  assign n57535 = ~n57533 & ~n57534;
  assign n57536 = pi1108 & ~pi1109;
  assign n57537 = ~pi1108 & pi1109;
  assign n57538 = ~pi1108 & ~pi1109;
  assign n57539 = pi1108 & pi1109;
  assign n57540 = ~n57538 & ~n57539;
  assign n57541 = ~n57536 & ~n57537;
  assign n57542 = ~pi1112 & ~pi1113;
  assign n57543 = pi1112 & pi1113;
  assign n57544 = pi1112 & ~pi1113;
  assign n57545 = ~pi1112 & pi1113;
  assign n57546 = ~n57544 & ~n57545;
  assign n57547 = ~n57542 & ~n57543;
  assign n57548 = ~pi1110 & ~pi1111;
  assign n57549 = pi1110 & pi1111;
  assign n57550 = pi1110 & ~pi1111;
  assign n57551 = ~pi1110 & pi1111;
  assign n57552 = ~n57550 & ~n57551;
  assign n57553 = ~n57548 & ~n57549;
  assign n57554 = ~n61572 & n61573;
  assign n57555 = n61572 & ~n61573;
  assign n57556 = ~n57554 & ~n57555;
  assign n57557 = ~n61571 & n57556;
  assign n57558 = n61571 & ~n57556;
  assign n57559 = ~n61571 & ~n61572;
  assign n57560 = n61571 & n61572;
  assign n57561 = ~n57559 & ~n57560;
  assign n57562 = n61573 & n57561;
  assign n57563 = ~n61573 & ~n57561;
  assign n57564 = ~n57562 & ~n57563;
  assign n57565 = ~n61571 & ~n61573;
  assign n57566 = n61571 & n61573;
  assign n57567 = ~n57565 & ~n57566;
  assign n57568 = n61572 & n57567;
  assign n57569 = ~n61572 & ~n57567;
  assign n57570 = ~n57568 & ~n57569;
  assign n57571 = ~n57557 & ~n57558;
  assign n57572 = ~n57535 & ~n61574;
  assign n57573 = pi828 & n57381;
  assign n57574 = n57531 & ~n57573;
  assign n57575 = ~n57534 & n61574;
  assign n57576 = ~n57574 & n57575;
  assign po985 = ~n57572 & ~n57576;
  assign n57578 = pi832 & ~pi1100;
  assign n57579 = n56862 & n57578;
  assign n57580 = ~pi1100 & po897;
  assign n57581 = ~pi603 & ~po897;
  assign n57582 = ~pi966 & ~n57581;
  assign n57583 = ~pi966 & ~n61575;
  assign n57584 = ~n57581 & n57583;
  assign n57585 = ~n61575 & n57582;
  assign n57586 = pi871 & pi966;
  assign n57587 = pi872 & pi966;
  assign n57588 = ~n57586 & ~n57587;
  assign n57589 = ~n61576 & n57588;
  assign n57590 = pi606 & ~po897;
  assign n57591 = pi1104 & po897;
  assign n57592 = ~pi606 & ~po897;
  assign n57593 = ~pi1104 & po897;
  assign n57594 = ~n57592 & ~n57593;
  assign n57595 = ~n57590 & ~n57591;
  assign n57596 = ~pi966 & n61577;
  assign n57597 = pi837 & pi966;
  assign n57598 = ~pi966 & ~n61577;
  assign n57599 = ~pi837 & pi966;
  assign n57600 = ~n57598 & ~n57599;
  assign n57601 = ~n57596 & ~n57597;
  assign n57602 = ~pi1102 & po897;
  assign n57603 = ~pi614 & ~po897;
  assign n57604 = ~pi966 & ~n57603;
  assign n57605 = ~pi966 & ~n57602;
  assign n57606 = ~n57603 & n57605;
  assign n57607 = ~n57602 & n57604;
  assign n57608 = ~n57586 & ~n61579;
  assign n57609 = ~pi1101 & po897;
  assign n57610 = ~pi616 & ~po897;
  assign n57611 = ~pi966 & ~n57610;
  assign n57612 = ~pi966 & ~n57609;
  assign n57613 = ~n57610 & n57612;
  assign n57614 = ~n57609 & n57611;
  assign n57615 = ~n57587 & ~n61580;
  assign n57616 = pi617 & ~po897;
  assign n57617 = pi1105 & po897;
  assign n57618 = ~pi617 & ~po897;
  assign n57619 = ~pi1105 & po897;
  assign n57620 = ~n57618 & ~n57619;
  assign n57621 = ~n57616 & ~n57617;
  assign n57622 = ~pi966 & n61581;
  assign n57623 = pi850 & pi966;
  assign n57624 = ~pi966 & ~n61581;
  assign n57625 = ~pi850 & pi966;
  assign n57626 = ~n57624 & ~n57625;
  assign n57627 = ~n57622 & ~n57623;
  assign n57628 = ~pi299 & pi983;
  assign n57629 = ~n37259 & ~n57628;
  assign n57630 = ~n56823 & n57629;
  assign n57631 = pi823 & n6518;
  assign n57632 = ~pi779 & n57631;
  assign n57633 = pi907 & n57628;
  assign n57634 = pi604 & ~n57633;
  assign n57635 = ~n57631 & n57634;
  assign n57636 = ~n57632 & ~n57635;
  assign n57637 = ~pi1107 & po897;
  assign n57638 = ~pi607 & ~po897;
  assign n57639 = ~pi966 & ~n57638;
  assign n57640 = ~pi966 & ~n57637;
  assign n57641 = ~n57638 & n57640;
  assign n57642 = ~n57637 & n57639;
  assign n57643 = ~pi1116 & po897;
  assign n57644 = ~pi608 & ~po897;
  assign n57645 = ~pi966 & ~n57644;
  assign n57646 = ~pi966 & ~n57643;
  assign n57647 = ~n57644 & n57646;
  assign n57648 = ~n57643 & n57645;
  assign n57649 = ~pi1118 & po897;
  assign n57650 = ~pi609 & ~po897;
  assign n57651 = ~pi966 & ~n57650;
  assign n57652 = ~pi966 & ~n57649;
  assign n57653 = ~n57650 & n57652;
  assign n57654 = ~n57649 & n57651;
  assign n57655 = ~pi1113 & po897;
  assign n57656 = ~pi610 & ~po897;
  assign n57657 = ~pi966 & ~n57656;
  assign n57658 = ~pi966 & ~n57655;
  assign n57659 = ~n57656 & n57658;
  assign n57660 = ~n57655 & n57657;
  assign n57661 = ~pi1114 & po897;
  assign n57662 = ~pi611 & ~po897;
  assign n57663 = ~pi966 & ~n57662;
  assign n57664 = ~pi966 & ~n57661;
  assign n57665 = ~n57662 & n57664;
  assign n57666 = ~n57661 & n57663;
  assign n57667 = ~pi1111 & po897;
  assign n57668 = ~pi612 & ~po897;
  assign n57669 = ~pi966 & ~n57668;
  assign n57670 = ~pi966 & ~n57667;
  assign n57671 = ~n57668 & n57670;
  assign n57672 = ~n57667 & n57669;
  assign n57673 = ~pi1115 & po897;
  assign n57674 = ~pi613 & ~po897;
  assign n57675 = ~pi966 & ~n57674;
  assign n57676 = ~pi966 & ~n57673;
  assign n57677 = ~n57674 & n57676;
  assign n57678 = ~n57673 & n57675;
  assign n57679 = ~pi1117 & po897;
  assign n57680 = ~pi618 & ~po897;
  assign n57681 = ~pi966 & ~n57680;
  assign n57682 = ~pi966 & ~n57679;
  assign n57683 = ~n57680 & n57682;
  assign n57684 = ~n57679 & n57681;
  assign n57685 = ~pi1122 & po897;
  assign n57686 = ~pi619 & ~po897;
  assign n57687 = ~pi966 & ~n57686;
  assign n57688 = ~pi966 & ~n57685;
  assign n57689 = ~n57686 & n57688;
  assign n57690 = ~n57685 & n57687;
  assign n57691 = ~pi1112 & po897;
  assign n57692 = ~pi620 & ~po897;
  assign n57693 = ~pi966 & ~n57692;
  assign n57694 = ~pi966 & ~n57691;
  assign n57695 = ~n57692 & n57694;
  assign n57696 = ~n57691 & n57693;
  assign n57697 = ~pi1108 & po897;
  assign n57698 = ~pi621 & ~po897;
  assign n57699 = ~pi966 & ~n57698;
  assign n57700 = ~pi966 & ~n57697;
  assign n57701 = ~n57698 & n57700;
  assign n57702 = ~n57697 & n57699;
  assign n57703 = ~pi1109 & po897;
  assign n57704 = ~pi622 & ~po897;
  assign n57705 = ~pi966 & ~n57704;
  assign n57706 = ~pi966 & ~n57703;
  assign n57707 = ~n57704 & n57706;
  assign n57708 = ~n57703 & n57705;
  assign n57709 = ~pi1106 & po897;
  assign n57710 = ~pi623 & ~po897;
  assign n57711 = ~pi966 & ~n57710;
  assign n57712 = ~pi966 & ~n57709;
  assign n57713 = ~n57710 & n57712;
  assign n57714 = ~n57709 & n57711;
  assign n57715 = pi831 & n6700;
  assign n57716 = ~pi780 & n57715;
  assign n57717 = pi947 & n57628;
  assign n57718 = pi624 & ~n57717;
  assign n57719 = ~n57715 & n57718;
  assign n57720 = ~n57716 & ~n57719;
  assign n57721 = ~pi1121 & po897;
  assign n57722 = ~pi626 & ~po897;
  assign n57723 = ~pi966 & ~n57722;
  assign n57724 = ~pi966 & ~n57721;
  assign n57725 = ~n57722 & n57724;
  assign n57726 = ~n57721 & n57723;
  assign n57727 = ~pi1103 & po897;
  assign n57728 = ~pi642 & ~po897;
  assign n57729 = ~pi966 & ~n57728;
  assign n57730 = ~pi966 & ~n57727;
  assign n57731 = ~n57728 & n57730;
  assign n57732 = ~n57727 & n57729;
  assign n57733 = pi1117 & po988;
  assign n57734 = ~pi753 & ~po988;
  assign n57735 = ~pi966 & ~n57734;
  assign n57736 = ~pi966 & ~n57733;
  assign n57737 = ~n57734 & n57736;
  assign n57738 = ~n57733 & n57735;
  assign n57739 = pi1118 & po988;
  assign n57740 = ~pi754 & ~po988;
  assign n57741 = ~pi966 & ~n57740;
  assign n57742 = ~pi966 & ~n57739;
  assign n57743 = ~n57740 & n57742;
  assign n57744 = ~n57739 & n57741;
  assign n57745 = pi1120 & po988;
  assign n57746 = ~pi755 & ~po988;
  assign n57747 = ~pi966 & ~n57746;
  assign n57748 = ~pi966 & ~n57745;
  assign n57749 = ~n57746 & n57748;
  assign n57750 = ~n57745 & n57747;
  assign n57751 = pi1119 & po988;
  assign n57752 = ~pi756 & ~po988;
  assign n57753 = ~pi966 & ~n57752;
  assign n57754 = ~pi966 & ~n57751;
  assign n57755 = ~n57752 & n57754;
  assign n57756 = ~n57751 & n57753;
  assign n57757 = pi1113 & po988;
  assign n57758 = ~pi757 & ~po988;
  assign n57759 = ~pi966 & ~n57758;
  assign n57760 = ~pi966 & ~n57757;
  assign n57761 = ~n57758 & n57760;
  assign n57762 = ~n57757 & n57759;
  assign n57763 = pi758 & ~po988;
  assign n57764 = pi1101 & po988;
  assign n57765 = ~pi966 & ~n57764;
  assign n57766 = ~pi966 & ~n57763;
  assign n57767 = ~n57764 & n57766;
  assign n57768 = ~n57763 & n57765;
  assign n57769 = pi759 & ~po988;
  assign n57770 = pi1100 & po988;
  assign n57771 = ~pi966 & ~n57770;
  assign n57772 = ~pi759 & ~po988;
  assign n57773 = n57306 & n57578;
  assign n57774 = ~n57772 & ~n57773;
  assign n57775 = ~pi966 & ~n57774;
  assign n57776 = ~n57769 & n57771;
  assign n57777 = pi1115 & po988;
  assign n57778 = ~pi760 & ~po988;
  assign n57779 = ~pi966 & ~n57778;
  assign n57780 = ~pi966 & ~n57777;
  assign n57781 = ~n57778 & n57780;
  assign n57782 = ~n57777 & n57779;
  assign n57783 = pi1121 & po988;
  assign n57784 = ~pi761 & ~po988;
  assign n57785 = ~pi966 & ~n57784;
  assign n57786 = ~pi966 & ~n57783;
  assign n57787 = ~n57784 & n57786;
  assign n57788 = ~n57783 & n57785;
  assign n57789 = pi1129 & po988;
  assign n57790 = ~pi762 & ~po988;
  assign n57791 = ~pi966 & ~n57790;
  assign n57792 = ~pi966 & ~n57789;
  assign n57793 = ~n57790 & n57792;
  assign n57794 = ~n57789 & n57791;
  assign n57795 = pi763 & ~po988;
  assign n57796 = pi1103 & po988;
  assign n57797 = ~pi966 & ~n57796;
  assign n57798 = ~pi966 & ~n57795;
  assign n57799 = ~n57796 & n57798;
  assign n57800 = ~n57795 & n57797;
  assign n57801 = pi764 & ~po988;
  assign n57802 = pi1107 & po988;
  assign n57803 = ~pi966 & ~n57802;
  assign n57804 = ~pi966 & ~n57801;
  assign n57805 = ~n57802 & n57804;
  assign n57806 = ~n57801 & n57803;
  assign n57807 = pi766 & ~po988;
  assign n57808 = pi1110 & po988;
  assign n57809 = ~pi966 & ~n57808;
  assign n57810 = ~pi966 & ~n57807;
  assign n57811 = ~n57808 & n57810;
  assign n57812 = ~n57807 & n57809;
  assign n57813 = pi1116 & po988;
  assign n57814 = ~pi767 & ~po988;
  assign n57815 = ~pi966 & ~n57814;
  assign n57816 = ~pi966 & ~n57813;
  assign n57817 = ~n57814 & n57816;
  assign n57818 = ~n57813 & n57815;
  assign n57819 = pi1125 & po988;
  assign n57820 = ~pi768 & ~po988;
  assign n57821 = ~pi966 & ~n57820;
  assign n57822 = ~pi966 & ~n57819;
  assign n57823 = ~n57820 & n57822;
  assign n57824 = ~n57819 & n57821;
  assign n57825 = pi1126 & po988;
  assign n57826 = ~pi770 & ~po988;
  assign n57827 = ~pi966 & ~n57826;
  assign n57828 = ~pi966 & ~n57825;
  assign n57829 = ~n57826 & n57828;
  assign n57830 = ~n57825 & n57827;
  assign n57831 = pi772 & ~po988;
  assign n57832 = pi1102 & po988;
  assign n57833 = ~pi966 & ~n57832;
  assign n57834 = ~pi966 & ~n57831;
  assign n57835 = ~n57832 & n57834;
  assign n57836 = ~n57831 & n57833;
  assign n57837 = pi1127 & po988;
  assign n57838 = ~pi774 & ~po988;
  assign n57839 = ~pi966 & ~n57838;
  assign n57840 = ~pi966 & ~n57837;
  assign n57841 = ~n57838 & n57840;
  assign n57842 = ~n57837 & n57839;
  assign n57843 = pi1128 & po988;
  assign n57844 = ~pi776 & ~po988;
  assign n57845 = ~pi966 & ~n57844;
  assign n57846 = ~pi966 & ~n57843;
  assign n57847 = ~n57844 & n57846;
  assign n57848 = ~n57843 & n57845;
  assign n57849 = pi1122 & po988;
  assign n57850 = ~pi777 & ~po988;
  assign n57851 = ~pi966 & ~n57850;
  assign n57852 = ~pi966 & ~n57849;
  assign n57853 = ~n57850 & n57852;
  assign n57854 = ~n57849 & n57851;
  assign n57855 = pi779 & ~n56829;
  assign n57856 = pi780 & ~n56824;
  assign n57857 = ~pi604 & ~pi979;
  assign n57858 = pi615 & pi979;
  assign n57859 = ~n57857 & ~n57858;
  assign n57860 = pi604 & ~pi979;
  assign n57861 = ~pi615 & pi979;
  assign n57862 = pi782 & ~n57861;
  assign n57863 = ~n57860 & n57862;
  assign n57864 = pi782 & ~n57859;
  assign n57865 = ~pi782 & ~pi907;
  assign n57866 = ~pi598 & pi979;
  assign n57867 = ~pi624 & ~pi979;
  assign n57868 = pi782 & ~n57867;
  assign n57869 = pi782 & ~n57866;
  assign n57870 = ~n57867 & n57869;
  assign n57871 = ~n57866 & n57868;
  assign n57872 = ~n57865 & ~n61619;
  assign po1063 = ~n61618 & n57872;
  assign n57874 = ~pi782 & pi947;
  assign n57875 = ~n61619 & ~n57874;
  assign n57876 = pi1093 & pi1154;
  assign n57877 = pi923 & ~pi1093;
  assign n57878 = ~pi923 & ~pi1093;
  assign n57879 = pi1093 & ~pi1154;
  assign n57880 = ~n57878 & ~n57879;
  assign n57881 = ~n57876 & ~n57877;
  assign n57882 = pi1093 & pi1155;
  assign n57883 = pi925 & ~pi1093;
  assign n57884 = ~pi925 & ~pi1093;
  assign n57885 = pi1093 & ~pi1155;
  assign n57886 = ~n57884 & ~n57885;
  assign n57887 = ~n57882 & ~n57883;
  assign n57888 = pi1093 & pi1157;
  assign n57889 = pi926 & ~pi1093;
  assign n57890 = ~pi926 & ~pi1093;
  assign n57891 = pi1093 & ~pi1157;
  assign n57892 = ~n57890 & ~n57891;
  assign n57893 = ~n57888 & ~n57889;
  assign n57894 = pi1093 & pi1150;
  assign n57895 = pi931 & ~pi1093;
  assign n57896 = ~pi931 & ~pi1093;
  assign n57897 = pi1093 & ~pi1150;
  assign n57898 = ~n57896 & ~n57897;
  assign n57899 = ~n57894 & ~n57895;
  assign n57900 = pi1093 & pi1147;
  assign n57901 = pi934 & ~pi1093;
  assign n57902 = ~pi934 & ~pi1093;
  assign n57903 = pi1093 & ~pi1147;
  assign n57904 = ~n57902 & ~n57903;
  assign n57905 = ~n57900 & ~n57901;
  assign n57906 = pi1093 & pi1149;
  assign n57907 = pi936 & ~pi1093;
  assign n57908 = ~pi936 & ~pi1093;
  assign n57909 = pi1093 & ~pi1149;
  assign n57910 = ~n57908 & ~n57909;
  assign n57911 = ~n57906 & ~n57907;
  assign n57912 = pi1093 & pi1148;
  assign n57913 = pi937 & ~pi1093;
  assign n57914 = ~pi937 & ~pi1093;
  assign n57915 = pi1093 & ~pi1148;
  assign n57916 = ~n57914 & ~n57915;
  assign n57917 = ~n57912 & ~n57913;
  assign n57918 = pi1093 & pi1153;
  assign n57919 = pi941 & ~pi1093;
  assign n57920 = ~pi941 & ~pi1093;
  assign n57921 = pi1093 & ~pi1153;
  assign n57922 = ~n57920 & ~n57921;
  assign n57923 = ~n57918 & ~n57919;
  assign n57924 = pi1093 & pi1156;
  assign n57925 = pi942 & ~pi1093;
  assign n57926 = ~pi942 & ~pi1093;
  assign n57927 = pi1093 & ~pi1156;
  assign n57928 = ~n57926 & ~n57927;
  assign n57929 = ~n57924 & ~n57925;
  assign n57930 = pi1093 & pi1151;
  assign n57931 = pi943 & ~pi1093;
  assign n57932 = ~pi943 & ~pi1093;
  assign n57933 = pi1093 & ~pi1151;
  assign n57934 = ~n57932 & ~n57933;
  assign n57935 = ~n57930 & ~n57931;
  assign n57936 = ~pi598 & pi615;
  assign n57937 = ~pi604 & ~pi624;
  assign n57938 = pi119 & pi1056;
  assign n57939 = ~pi228 & pi252;
  assign n57940 = ~pi119 & ~n57939;
  assign n57941 = ~pi468 & ~n57940;
  assign n57942 = ~n57938 & n57941;
  assign n57943 = pi119 & pi1077;
  assign n57944 = n57941 & ~n57943;
  assign n57945 = pi119 & pi1073;
  assign n57946 = n57941 & ~n57945;
  assign n57947 = pi119 & pi1041;
  assign n57948 = n57941 & ~n57947;
  assign n57949 = pi119 & pi232;
  assign po236 = ~pi468 & n57949;
  assign n57951 = pi124 & ~pi468;
  assign n57952 = ~pi298 & pi478;
  assign n57953 = ~pi478 & ~pi1044;
  assign n57954 = ~pi478 & pi1044;
  assign n57955 = pi298 & pi478;
  assign n57956 = ~n57954 & ~n57955;
  assign n57957 = ~n57952 & ~n57953;
  assign n57958 = ~pi303 & pi478;
  assign n57959 = ~pi478 & ~pi1049;
  assign n57960 = ~pi478 & pi1049;
  assign n57961 = pi303 & pi478;
  assign n57962 = ~n57960 & ~n57961;
  assign n57963 = ~n57958 & ~n57959;
  assign n57964 = ~pi304 & pi478;
  assign n57965 = ~pi478 & ~pi1048;
  assign n57966 = ~pi478 & pi1048;
  assign n57967 = pi304 & pi478;
  assign n57968 = ~n57966 & ~n57967;
  assign n57969 = ~n57964 & ~n57965;
  assign n57970 = ~pi305 & pi478;
  assign n57971 = ~pi478 & ~pi1084;
  assign n57972 = ~pi478 & pi1084;
  assign n57973 = pi305 & pi478;
  assign n57974 = ~n57972 & ~n57973;
  assign n57975 = ~n57970 & ~n57971;
  assign n57976 = ~pi306 & pi478;
  assign n57977 = ~pi478 & ~pi1059;
  assign n57978 = ~pi478 & pi1059;
  assign n57979 = pi306 & pi478;
  assign n57980 = ~n57978 & ~n57979;
  assign n57981 = ~n57976 & ~n57977;
  assign n57982 = ~pi307 & pi478;
  assign n57983 = ~pi478 & ~pi1053;
  assign n57984 = ~pi478 & pi1053;
  assign n57985 = pi307 & pi478;
  assign n57986 = ~n57984 & ~n57985;
  assign n57987 = ~n57982 & ~n57983;
  assign n57988 = ~pi308 & pi478;
  assign n57989 = ~pi478 & ~pi1037;
  assign n57990 = ~pi478 & pi1037;
  assign n57991 = pi308 & pi478;
  assign n57992 = ~n57990 & ~n57991;
  assign n57993 = ~n57988 & ~n57989;
  assign n57994 = ~pi309 & pi478;
  assign n57995 = ~pi478 & ~pi1072;
  assign n57996 = ~pi478 & pi1072;
  assign n57997 = pi309 & pi478;
  assign n57998 = ~n57996 & ~n57997;
  assign n57999 = ~n57994 & ~n57995;
  assign n58000 = ~pi599 & pi810;
  assign n58001 = pi596 & ~n58000;
  assign n58002 = pi804 & ~n58001;
  assign n58003 = pi815 & ~n58002;
  assign n58004 = pi595 & ~n58003;
  assign n58005 = ~pi804 & ~pi810;
  assign n58006 = ~pi595 & ~n58005;
  assign n58007 = pi594 & pi600;
  assign n58008 = pi597 & n58007;
  assign n58009 = pi601 & n58008;
  assign n58010 = ~n58006 & n58009;
  assign n58011 = ~pi595 & n58005;
  assign n58012 = pi595 & pi815;
  assign n58013 = ~n58002 & n58012;
  assign n58014 = ~n58011 & ~n58013;
  assign n58015 = n58009 & ~n58014;
  assign n58016 = ~n58004 & n58010;
  assign n58017 = ~pi601 & ~n58005;
  assign n58018 = pi600 & ~pi810;
  assign n58019 = pi804 & ~n58018;
  assign n58020 = ~pi815 & ~n58019;
  assign n58021 = ~pi815 & ~n58017;
  assign n58022 = ~n58019 & n58021;
  assign n58023 = ~n58017 & n58020;
  assign n58024 = ~n61638 & ~n61639;
  assign n58025 = pi605 & ~n58024;
  assign n58026 = pi990 & n58007;
  assign n58027 = ~pi815 & n58019;
  assign n58028 = n58026 & n58027;
  assign n58029 = ~n58025 & ~n58028;
  assign po614 = pi821 & ~n58029;
  assign n58031 = ~pi123 & n2872;
  assign n58032 = ~pi591 & n58031;
  assign n58033 = ~pi588 & ~n58031;
  assign n58034 = n45087 & ~n58033;
  assign n58035 = n45087 & ~n58032;
  assign n58036 = ~n58033 & n58035;
  assign n58037 = ~n58032 & n58034;
  assign n58038 = pi590 & ~n58031;
  assign n58039 = pi588 & n58031;
  assign n58040 = n45087 & ~n58039;
  assign n58041 = n45087 & ~n58038;
  assign n58042 = ~n58039 & n58041;
  assign n58043 = ~n58038 & n58040;
  assign n58044 = ~pi592 & n58031;
  assign n58045 = ~pi591 & ~n58031;
  assign n58046 = n45087 & ~n58045;
  assign n58047 = n45087 & ~n58044;
  assign n58048 = ~n58045 & n58047;
  assign n58049 = ~n58044 & n58046;
  assign n58050 = ~pi590 & n58031;
  assign n58051 = ~pi592 & ~n58031;
  assign n58052 = n45087 & ~n58051;
  assign n58053 = n45087 & ~n58050;
  assign n58054 = ~n58051 & n58053;
  assign n58055 = ~n58050 & n58052;
  assign n58056 = ~pi332 & ~pi806;
  assign n58057 = pi990 & n58056;
  assign n58058 = pi595 & n58008;
  assign n58059 = n58057 & n58058;
  assign n58060 = pi596 & n58059;
  assign n58061 = ~pi332 & pi599;
  assign n58062 = ~n58060 & ~n58061;
  assign n58063 = pi599 & n58060;
  assign po756 = ~n58062 & ~n58063;
  assign n58065 = pi605 & ~pi806;
  assign n58066 = n58009 & n58065;
  assign n58067 = pi595 & n58066;
  assign n58068 = ~pi595 & ~n58066;
  assign n58069 = ~pi332 & ~n58068;
  assign po752 = ~n58067 & n58069;
  assign n58071 = ~pi332 & pi596;
  assign n58072 = ~n58059 & ~n58071;
  assign po753 = ~n58060 & ~n58072;
  assign n58074 = ~pi806 & n58026;
  assign n58075 = pi597 & n58074;
  assign n58076 = ~pi597 & ~n58074;
  assign n58077 = ~pi332 & ~n58076;
  assign po754 = ~n58075 & n58077;
  assign n58079 = pi600 & n58057;
  assign n58080 = ~pi332 & pi594;
  assign n58081 = ~n58079 & ~n58080;
  assign po751 = ~n58074 & ~n58081;
  assign n58083 = ~pi332 & pi600;
  assign n58084 = ~n58057 & ~n58083;
  assign po757 = ~n58079 & ~n58084;
  assign n58086 = ~pi601 & pi806;
  assign n58087 = ~pi806 & ~pi989;
  assign n58088 = ~pi332 & ~n58087;
  assign n58089 = ~pi332 & ~n58086;
  assign n58090 = ~n58087 & n58089;
  assign n58091 = ~n58086 & n58088;
  assign n58092 = ~pi287 & pi457;
  assign po444 = ~pi332 & ~n58092;
  assign n58094 = ~pi605 & ~n58056;
  assign n58095 = ~pi332 & ~n58065;
  assign po762 = ~n58094 & n58095;
  assign n58097 = pi721 & pi813;
  assign n58098 = pi765 & ~pi798;
  assign n58099 = ~pi765 & pi798;
  assign n58100 = ~pi765 & ~pi798;
  assign n58101 = pi765 & pi798;
  assign n58102 = ~n58100 & ~n58101;
  assign n58103 = ~n58098 & ~n58099;
  assign n58104 = pi807 & ~n61645;
  assign n58105 = pi747 & n58104;
  assign n58106 = ~pi747 & ~pi807;
  assign n58107 = ~n61645 & n58106;
  assign n58108 = ~n58105 & ~n58107;
  assign n58109 = ~pi771 & ~pi800;
  assign n58110 = pi771 & pi800;
  assign n58111 = ~n58109 & ~n58110;
  assign n58112 = ~pi769 & ~pi794;
  assign n58113 = pi769 & pi794;
  assign n58114 = ~n58112 & ~n58113;
  assign n58115 = ~n58111 & ~n58114;
  assign n58116 = ~n58108 & ~n58114;
  assign n58117 = ~n58111 & n58116;
  assign n58118 = ~n58108 & n58115;
  assign n58119 = pi773 & ~pi801;
  assign n58120 = ~pi773 & pi801;
  assign n58121 = ~pi773 & ~pi801;
  assign n58122 = pi773 & pi801;
  assign n58123 = ~n58121 & ~n58122;
  assign n58124 = ~n58119 & ~n58120;
  assign n58125 = n61646 & ~n61647;
  assign n58126 = n58097 & n58125;
  assign n58127 = ~pi775 & ~pi816;
  assign n58128 = pi775 & pi816;
  assign n58129 = ~n58127 & ~n58128;
  assign n58130 = n58126 & ~n58129;
  assign n58131 = pi731 & ~pi945;
  assign n58132 = pi775 & n58131;
  assign n58133 = pi988 & n58132;
  assign n58134 = ~n58130 & ~n58133;
  assign n58135 = ~pi945 & pi988;
  assign n58136 = pi731 & n58135;
  assign n58137 = ~pi731 & ~pi795;
  assign n58138 = pi731 & pi795;
  assign n58139 = ~n58137 & ~n58138;
  assign n58140 = ~n58136 & n58139;
  assign n58141 = ~n58134 & ~n58140;
  assign n58142 = pi721 & ~pi775;
  assign n58143 = ~n58130 & n58142;
  assign n58144 = n58130 & ~n58139;
  assign n58145 = pi721 & ~n58136;
  assign n58146 = ~n58144 & n58145;
  assign n58147 = ~n58143 & ~n58146;
  assign n58148 = pi721 & ~n58141;
  assign n58149 = ~pi721 & ~pi813;
  assign n58150 = pi794 & pi801;
  assign n58151 = n58149 & n58150;
  assign n58152 = ~n58111 & n58151;
  assign n58153 = n58104 & ~n58111;
  assign n58154 = n58151 & n58153;
  assign n58155 = n58104 & n58152;
  assign n58156 = ~n58126 & ~n61649;
  assign n58157 = pi816 & ~n58156;
  assign n58158 = pi775 & ~n58157;
  assign n58159 = pi795 & ~n58158;
  assign n58160 = pi747 & pi773;
  assign n58161 = pi769 & pi775;
  assign n58162 = n58160 & n58161;
  assign n58163 = pi721 & n58162;
  assign n58164 = ~pi721 & ~n58162;
  assign n58165 = n58136 & ~n58164;
  assign n58166 = pi769 & n58160;
  assign n58167 = ~pi721 & ~n58166;
  assign n58168 = pi721 & n58166;
  assign n58169 = pi775 & ~n58168;
  assign n58170 = ~n58167 & n58169;
  assign n58171 = ~n58142 & ~n58170;
  assign n58172 = n58136 & ~n58171;
  assign n58173 = ~n58163 & n58165;
  assign n58174 = ~n58157 & n58170;
  assign n58175 = pi795 & ~n58174;
  assign n58176 = n61650 & ~n58175;
  assign n58177 = ~n58159 & n61650;
  assign n58178 = n61648 & ~n61651;
  assign n58179 = ~n58097 & ~n58149;
  assign n58180 = n58125 & ~n58179;
  assign n58181 = pi795 & ~n58129;
  assign n58182 = n58180 & n58181;
  assign n58183 = pi731 & n58182;
  assign n58184 = n58135 & n58160;
  assign n58185 = pi731 & n58184;
  assign n58186 = ~n58129 & ~n58179;
  assign n58187 = ~n58111 & n58186;
  assign n58188 = ~pi795 & pi801;
  assign n58189 = ~n58114 & n58188;
  assign n58190 = n58104 & n58189;
  assign n58191 = n58186 & n58189;
  assign n58192 = n58153 & n58191;
  assign n58193 = n58187 & n58190;
  assign n58194 = n58184 & ~n61652;
  assign n58195 = ~pi731 & ~n58194;
  assign n58196 = ~n58185 & ~n58195;
  assign n58197 = ~n58160 & ~n58182;
  assign n58198 = n58136 & ~n58197;
  assign n58199 = pi731 & ~n58182;
  assign n58200 = n58160 & ~n61652;
  assign n58201 = ~pi731 & ~n58200;
  assign n58202 = n58135 & ~n58201;
  assign n58203 = ~n58199 & ~n58202;
  assign n58204 = ~n58198 & ~n58203;
  assign n58205 = ~n58183 & n58196;
  assign n58206 = pi801 & n58107;
  assign n58207 = pi773 & n58135;
  assign n58208 = ~n61647 & ~n58207;
  assign n58209 = n58104 & n58208;
  assign n58210 = ~n58206 & ~n58209;
  assign n58211 = ~n58139 & n58186;
  assign n58212 = n58115 & n58211;
  assign n58213 = ~n58210 & n58212;
  assign n58214 = ~pi747 & ~n58207;
  assign n58215 = ~n58184 & ~n58214;
  assign po904 = ~n58213 & n58215;
  assign n58217 = n58128 & n58180;
  assign n58218 = pi794 & ~n61647;
  assign n58219 = ~n58111 & n58218;
  assign n58220 = n58186 & n58219;
  assign n58221 = n58187 & n58218;
  assign n58222 = ~n58108 & n61654;
  assign n58223 = ~pi775 & n58222;
  assign n58224 = ~n58217 & ~n58223;
  assign n58225 = pi795 & ~n58224;
  assign n58226 = pi775 & n58160;
  assign n58227 = pi769 & ~n58226;
  assign n58228 = ~pi769 & n58226;
  assign n58229 = ~n58227 & ~n58228;
  assign n58230 = n58136 & ~n58229;
  assign n58231 = ~n58225 & n58230;
  assign n58232 = ~n58139 & n58222;
  assign n58233 = pi769 & ~n58136;
  assign n58234 = ~n58232 & n58233;
  assign n58235 = ~n58231 & ~n58234;
  assign n58236 = ~pi765 & ~pi773;
  assign n58237 = ~n58110 & n58236;
  assign n58238 = ~n58113 & n58237;
  assign n58239 = ~n58105 & n58238;
  assign n58240 = ~pi765 & ~n58110;
  assign n58241 = ~n58113 & n58240;
  assign n58242 = ~n58105 & n58241;
  assign n58243 = n58121 & ~n58242;
  assign n58244 = ~n58122 & ~n58243;
  assign n58245 = n61646 & ~n58244;
  assign n58246 = n58125 & ~n58239;
  assign n58247 = ~pi721 & ~n61655;
  assign n58248 = n58127 & ~n58247;
  assign n58249 = ~n58128 & ~n58248;
  assign n58250 = n58137 & ~n58249;
  assign n58251 = ~n58129 & n58138;
  assign n58252 = ~n58250 & ~n58251;
  assign po963 = n58180 & ~n58252;
  assign n58254 = ~pi945 & pi987;
  assign n58255 = ~po963 & n58254;
  assign po978 = n58125 & n58211;
  assign n58257 = pi771 & pi945;
  assign n58258 = ~po978 & n58257;
  assign n58259 = ~n58255 & ~n58258;
  assign n58260 = ~pi801 & n61646;
  assign n58261 = po963 & n58260;
  assign n58262 = n58135 & ~n58261;
  assign n58263 = pi801 & n58211;
  assign n58264 = n61646 & n58263;
  assign n58265 = pi801 & ~n58211;
  assign n58266 = n58125 & ~n58265;
  assign n58267 = pi773 & ~n58266;
  assign n58268 = pi773 & ~n58264;
  assign n58269 = ~n58262 & ~n61656;
  assign po930 = ~n58207 & ~n58269;
  assign n58271 = pi765 & ~po978;
  assign n58272 = pi945 & ~n58271;
  assign n58273 = ~n58126 & ~n58149;
  assign n58274 = n58248 & ~n58273;
  assign n58275 = ~n58217 & ~n58274;
  assign n58276 = n58137 & ~n58275;
  assign n58277 = ~pi765 & ~n58183;
  assign n58278 = ~pi765 & ~n58217;
  assign n58279 = ~n58274 & n58278;
  assign n58280 = ~pi795 & ~n58279;
  assign n58281 = ~pi731 & ~n58280;
  assign n58282 = ~n58199 & ~n58281;
  assign n58283 = ~pi765 & ~n58282;
  assign n58284 = ~n58276 & n58277;
  assign n58285 = ~pi945 & ~n61657;
  assign po922 = ~n58272 & ~n58285;
  assign n58287 = pi765 & pi771;
  assign n58288 = n58160 & n58287;
  assign n58289 = ~n58182 & ~n58288;
  assign n58290 = n58132 & ~n58289;
  assign n58291 = pi775 & ~po978;
  assign n58292 = pi795 & pi800;
  assign n58293 = pi801 & ~pi816;
  assign n58294 = n58292 & n58293;
  assign n58295 = ~n58114 & n58294;
  assign n58296 = ~n58179 & n58295;
  assign n58297 = ~n58179 & n58294;
  assign n58298 = n58116 & n58297;
  assign n58299 = ~n58108 & n58296;
  assign n58300 = n58288 & ~n61658;
  assign n58301 = ~pi775 & ~n58300;
  assign n58302 = n58131 & ~n58301;
  assign n58303 = ~n58131 & po978;
  assign n58304 = pi775 & ~n58303;
  assign n58305 = n58131 & n58288;
  assign n58306 = ~n61658 & n58305;
  assign n58307 = ~n58304 & ~n58306;
  assign n58308 = ~n58291 & ~n58302;
  assign po932 = ~n58290 & ~n61659;
  assign n58310 = pi832 & pi956;
  assign n58311 = ~pi1046 & ~pi1083;
  assign n58312 = pi1085 & n58311;
  assign n58313 = n58310 & n58312;
  assign n58314 = ~pi968 & n58313;
  assign n58315 = pi778 & ~n58314;
  assign n58316 = pi1100 & n58314;
  assign n58317 = ~n58315 & ~n58316;
  assign n58318 = pi781 & ~n58314;
  assign n58319 = pi1101 & n58314;
  assign n58320 = ~n58318 & ~n58319;
  assign n58321 = pi783 & ~n58314;
  assign n58322 = pi1109 & n58314;
  assign n58323 = ~n58321 & ~n58322;
  assign n58324 = pi784 & ~n58314;
  assign n58325 = pi1110 & n58314;
  assign n58326 = ~n58324 & ~n58325;
  assign n58327 = pi785 & ~n58314;
  assign n58328 = pi1102 & n58314;
  assign n58329 = ~n58327 & ~n58328;
  assign n58330 = pi787 & ~n58314;
  assign n58331 = pi1104 & n58314;
  assign n58332 = ~n58330 & ~n58331;
  assign n58333 = pi788 & ~n58314;
  assign n58334 = pi1105 & n58314;
  assign n58335 = ~n58333 & ~n58334;
  assign n58336 = pi789 & ~n58314;
  assign n58337 = pi1106 & n58314;
  assign n58338 = ~n58336 & ~n58337;
  assign n58339 = pi790 & ~n58314;
  assign n58340 = pi1107 & n58314;
  assign n58341 = ~n58339 & ~n58340;
  assign n58342 = pi791 & ~n58314;
  assign n58343 = pi1108 & n58314;
  assign n58344 = ~n58342 & ~n58343;
  assign n58345 = pi792 & ~n58314;
  assign n58346 = pi1103 & n58314;
  assign n58347 = ~n58345 & ~n58346;
  assign n58348 = pi968 & n58313;
  assign n58349 = pi794 & ~n58348;
  assign n58350 = pi1130 & n58348;
  assign n58351 = ~n58349 & ~n58350;
  assign n58352 = pi795 & ~n58348;
  assign n58353 = pi1128 & n58348;
  assign n58354 = ~n58352 & ~n58353;
  assign n58355 = pi798 & ~n58348;
  assign n58356 = pi1124 & n58348;
  assign n58357 = ~n58355 & ~n58356;
  assign n58358 = pi799 & ~n58348;
  assign n58359 = ~pi1107 & n58348;
  assign po956 = ~n58358 & ~n58359;
  assign n58361 = pi800 & ~n58348;
  assign n58362 = pi1125 & n58348;
  assign n58363 = ~n58361 & ~n58362;
  assign n58364 = pi801 & ~n58348;
  assign n58365 = pi1126 & n58348;
  assign n58366 = ~n58364 & ~n58365;
  assign n58367 = pi803 & ~n58348;
  assign n58368 = ~pi1106 & n58348;
  assign po960 = ~n58367 & ~n58368;
  assign n58370 = pi804 & ~n58348;
  assign n58371 = pi1109 & n58348;
  assign n58372 = ~n58370 & ~n58371;
  assign n58373 = pi807 & ~n58348;
  assign n58374 = pi1127 & n58348;
  assign n58375 = ~n58373 & ~n58374;
  assign n58376 = pi808 & ~n58348;
  assign n58377 = pi1101 & n58348;
  assign n58378 = ~n58376 & ~n58377;
  assign n58379 = pi809 & ~n58348;
  assign n58380 = ~pi1103 & n58348;
  assign po966 = ~n58379 & ~n58380;
  assign n58382 = pi810 & ~n58348;
  assign n58383 = pi1108 & n58348;
  assign n58384 = ~n58382 & ~n58383;
  assign n58385 = pi811 & ~n58348;
  assign n58386 = pi1102 & n58348;
  assign n58387 = ~n58385 & ~n58386;
  assign n58388 = pi812 & ~n58348;
  assign n58389 = ~pi1104 & n58348;
  assign po969 = ~n58388 & ~n58389;
  assign n58391 = pi813 & ~n58348;
  assign n58392 = pi1131 & n58348;
  assign n58393 = ~n58391 & ~n58392;
  assign n58394 = pi814 & ~n58348;
  assign n58395 = ~pi1105 & n58348;
  assign po971 = ~n58394 & ~n58395;
  assign n58397 = pi815 & ~n58348;
  assign n58398 = pi1110 & n58348;
  assign n58399 = ~n58397 & ~n58398;
  assign n58400 = pi816 & ~n58348;
  assign n58401 = pi1129 & n58348;
  assign n58402 = ~n58400 & ~n58401;
  assign po979 = ~pi811 & ~pi893;
  assign n58404 = ~pi837 & pi955;
  assign n58405 = ~pi955 & ~pi1049;
  assign n58406 = ~pi955 & pi1049;
  assign n58407 = pi837 & pi955;
  assign n58408 = ~n58406 & ~n58407;
  assign n58409 = ~n58404 & ~n58405;
  assign n58410 = ~pi838 & pi955;
  assign n58411 = ~pi955 & ~pi1047;
  assign n58412 = ~pi955 & pi1047;
  assign n58413 = pi838 & pi955;
  assign n58414 = ~n58412 & ~n58413;
  assign n58415 = ~n58410 & ~n58411;
  assign n58416 = ~pi839 & pi955;
  assign n58417 = ~pi955 & ~pi1074;
  assign n58418 = ~pi955 & pi1074;
  assign n58419 = pi839 & pi955;
  assign n58420 = ~n58418 & ~n58419;
  assign n58421 = ~n58416 & ~n58417;
  assign n58422 = ~pi842 & pi955;
  assign n58423 = ~pi955 & ~pi1035;
  assign n58424 = ~pi955 & pi1035;
  assign n58425 = pi842 & pi955;
  assign n58426 = ~n58424 & ~n58425;
  assign n58427 = ~n58422 & ~n58423;
  assign n58428 = ~pi843 & pi955;
  assign n58429 = ~pi955 & ~pi1079;
  assign n58430 = ~pi955 & pi1079;
  assign n58431 = pi843 & pi955;
  assign n58432 = ~n58430 & ~n58431;
  assign n58433 = ~n58428 & ~n58429;
  assign n58434 = ~pi844 & pi955;
  assign n58435 = ~pi955 & ~pi1078;
  assign n58436 = ~pi955 & pi1078;
  assign n58437 = pi844 & pi955;
  assign n58438 = ~n58436 & ~n58437;
  assign n58439 = ~n58434 & ~n58435;
  assign n58440 = ~pi845 & pi955;
  assign n58441 = ~pi955 & ~pi1043;
  assign n58442 = ~pi955 & pi1043;
  assign n58443 = pi845 & pi955;
  assign n58444 = ~n58442 & ~n58443;
  assign n58445 = ~n58440 & ~n58441;
  assign n58446 = ~pi847 & pi955;
  assign n58447 = ~pi955 & ~pi1055;
  assign n58448 = ~pi955 & pi1055;
  assign n58449 = pi847 & pi955;
  assign n58450 = ~n58448 & ~n58449;
  assign n58451 = ~n58446 & ~n58447;
  assign n58452 = ~pi848 & pi955;
  assign n58453 = ~pi955 & ~pi1039;
  assign n58454 = ~pi955 & pi1039;
  assign n58455 = pi848 & pi955;
  assign n58456 = ~n58454 & ~n58455;
  assign n58457 = ~n58452 & ~n58453;
  assign n58458 = ~pi850 & pi955;
  assign n58459 = ~pi955 & ~pi1048;
  assign n58460 = ~pi955 & pi1048;
  assign n58461 = pi850 & pi955;
  assign n58462 = ~n58460 & ~n58461;
  assign n58463 = ~n58458 & ~n58459;
  assign n58464 = ~pi851 & pi955;
  assign n58465 = ~pi955 & ~pi1045;
  assign n58466 = ~pi955 & pi1045;
  assign n58467 = pi851 & pi955;
  assign n58468 = ~n58466 & ~n58467;
  assign n58469 = ~n58464 & ~n58465;
  assign n58470 = ~pi852 & pi955;
  assign n58471 = ~pi955 & ~pi1062;
  assign n58472 = ~pi955 & pi1062;
  assign n58473 = pi852 & pi955;
  assign n58474 = ~n58472 & ~n58473;
  assign n58475 = ~n58470 & ~n58471;
  assign n58476 = ~pi853 & pi955;
  assign n58477 = ~pi955 & ~pi1080;
  assign n58478 = ~pi955 & pi1080;
  assign n58479 = pi853 & pi955;
  assign n58480 = ~n58478 & ~n58479;
  assign n58481 = ~n58476 & ~n58477;
  assign n58482 = ~pi854 & pi955;
  assign n58483 = ~pi955 & ~pi1051;
  assign n58484 = ~pi955 & pi1051;
  assign n58485 = pi854 & pi955;
  assign n58486 = ~n58484 & ~n58485;
  assign n58487 = ~n58482 & ~n58483;
  assign n58488 = ~pi855 & pi955;
  assign n58489 = ~pi955 & ~pi1065;
  assign n58490 = ~pi955 & pi1065;
  assign n58491 = pi855 & pi955;
  assign n58492 = ~n58490 & ~n58491;
  assign n58493 = ~n58488 & ~n58489;
  assign n58494 = ~pi856 & pi955;
  assign n58495 = ~pi955 & ~pi1067;
  assign n58496 = ~pi955 & pi1067;
  assign n58497 = pi856 & pi955;
  assign n58498 = ~n58496 & ~n58497;
  assign n58499 = ~n58494 & ~n58495;
  assign n58500 = ~pi857 & pi955;
  assign n58501 = ~pi955 & ~pi1058;
  assign n58502 = ~pi955 & pi1058;
  assign n58503 = pi857 & pi955;
  assign n58504 = ~n58502 & ~n58503;
  assign n58505 = ~n58500 & ~n58501;
  assign n58506 = ~pi858 & pi955;
  assign n58507 = ~pi955 & ~pi1087;
  assign n58508 = ~pi955 & pi1087;
  assign n58509 = pi858 & pi955;
  assign n58510 = ~n58508 & ~n58509;
  assign n58511 = ~n58506 & ~n58507;
  assign n58512 = ~pi859 & pi955;
  assign n58513 = ~pi955 & ~pi1070;
  assign n58514 = ~pi955 & pi1070;
  assign n58515 = pi859 & pi955;
  assign n58516 = ~n58514 & ~n58515;
  assign n58517 = ~n58512 & ~n58513;
  assign n58518 = ~pi860 & pi955;
  assign n58519 = ~pi955 & ~pi1076;
  assign n58520 = ~pi955 & pi1076;
  assign n58521 = pi860 & pi955;
  assign n58522 = ~n58520 & ~n58521;
  assign n58523 = ~n58518 & ~n58519;
  assign n58524 = ~pi865 & pi955;
  assign n58525 = ~pi955 & ~pi1040;
  assign n58526 = ~pi955 & pi1040;
  assign n58527 = pi865 & pi955;
  assign n58528 = ~n58526 & ~n58527;
  assign n58529 = ~n58524 & ~n58525;
  assign n58530 = ~pi866 & pi955;
  assign n58531 = ~pi955 & ~pi1053;
  assign n58532 = ~pi955 & pi1053;
  assign n58533 = pi866 & pi955;
  assign n58534 = ~n58532 & ~n58533;
  assign n58535 = ~n58530 & ~n58531;
  assign n58536 = ~pi867 & pi955;
  assign n58537 = ~pi955 & ~pi1057;
  assign n58538 = ~pi955 & pi1057;
  assign n58539 = pi867 & pi955;
  assign n58540 = ~n58538 & ~n58539;
  assign n58541 = ~n58536 & ~n58537;
  assign n58542 = ~pi868 & pi955;
  assign n58543 = ~pi955 & ~pi1063;
  assign n58544 = ~pi955 & pi1063;
  assign n58545 = pi868 & pi955;
  assign n58546 = ~n58544 & ~n58545;
  assign n58547 = ~n58542 & ~n58543;
  assign n58548 = ~pi870 & pi955;
  assign n58549 = ~pi955 & ~pi1069;
  assign n58550 = ~pi955 & pi1069;
  assign n58551 = pi870 & pi955;
  assign n58552 = ~n58550 & ~n58551;
  assign n58553 = ~n58548 & ~n58549;
  assign n58554 = ~pi871 & pi955;
  assign n58555 = ~pi955 & ~pi1072;
  assign n58556 = ~pi955 & pi1072;
  assign n58557 = pi871 & pi955;
  assign n58558 = ~n58556 & ~n58557;
  assign n58559 = ~n58554 & ~n58555;
  assign n58560 = ~pi872 & pi955;
  assign n58561 = ~pi955 & ~pi1084;
  assign n58562 = ~pi955 & pi1084;
  assign n58563 = pi872 & pi955;
  assign n58564 = ~n58562 & ~n58563;
  assign n58565 = ~n58560 & ~n58561;
  assign n58566 = ~pi873 & pi955;
  assign n58567 = ~pi955 & ~pi1044;
  assign n58568 = ~pi955 & pi1044;
  assign n58569 = pi873 & pi955;
  assign n58570 = ~n58568 & ~n58569;
  assign n58571 = ~n58566 & ~n58567;
  assign n58572 = ~pi874 & pi955;
  assign n58573 = ~pi955 & ~pi1036;
  assign n58574 = ~pi955 & pi1036;
  assign n58575 = pi874 & pi955;
  assign n58576 = ~n58574 & ~n58575;
  assign n58577 = ~n58572 & ~n58573;
  assign n58578 = ~pi876 & pi955;
  assign n58579 = ~pi955 & ~pi1037;
  assign n58580 = ~pi955 & pi1037;
  assign n58581 = pi876 & pi955;
  assign n58582 = ~n58580 & ~n58581;
  assign n58583 = ~n58578 & ~n58579;
  assign n58584 = ~pi880 & pi955;
  assign n58585 = ~pi955 & ~pi1081;
  assign n58586 = ~pi955 & pi1081;
  assign n58587 = pi880 & pi955;
  assign n58588 = ~n58586 & ~n58587;
  assign n58589 = ~n58584 & ~n58585;
  assign n58590 = ~pi881 & pi955;
  assign n58591 = ~pi955 & ~pi1059;
  assign n58592 = ~pi955 & pi1059;
  assign n58593 = pi881 & pi955;
  assign n58594 = ~n58592 & ~n58593;
  assign n58595 = ~n58590 & ~n58591;
  assign n58596 = ~pi883 & n57381;
  assign n58597 = ~n57481 & ~n58596;
  assign n58598 = pi1124 & ~n57381;
  assign n58599 = ~pi884 & n57381;
  assign n58600 = ~n58598 & ~n58599;
  assign n58601 = pi1125 & ~n57381;
  assign n58602 = ~pi885 & n57381;
  assign n58603 = ~n58601 & ~n58602;
  assign n58604 = pi1109 & ~n57381;
  assign n58605 = ~pi886 & n57381;
  assign n58606 = ~n58604 & ~n58605;
  assign n58607 = ~pi887 & n57381;
  assign n58608 = ~n57480 & ~n58607;
  assign n58609 = pi1120 & ~n57381;
  assign n58610 = ~pi888 & n57381;
  assign n58611 = ~n58609 & ~n58610;
  assign n58612 = pi1103 & ~n57381;
  assign n58613 = ~pi889 & n57381;
  assign n58614 = ~n58612 & ~n58613;
  assign n58615 = pi1126 & ~n57381;
  assign n58616 = ~pi890 & n57381;
  assign n58617 = ~n58615 & ~n58616;
  assign n58618 = pi1116 & ~n57381;
  assign n58619 = ~pi891 & n57381;
  assign n58620 = ~n58618 & ~n58619;
  assign n58621 = pi1101 & ~n57381;
  assign n58622 = ~pi892 & n57381;
  assign n58623 = ~n58621 & ~n58622;
  assign n58624 = pi1119 & ~n57381;
  assign n58625 = ~pi894 & n57381;
  assign n58626 = ~n58624 & ~n58625;
  assign n58627 = pi1113 & ~n57381;
  assign n58628 = ~pi895 & n57381;
  assign n58629 = ~n58627 & ~n58628;
  assign n58630 = pi1118 & ~n57381;
  assign n58631 = ~pi896 & n57381;
  assign n58632 = ~n58630 & ~n58631;
  assign n58633 = pi1129 & ~n57381;
  assign n58634 = ~pi898 & n57381;
  assign n58635 = ~n58633 & ~n58634;
  assign n58636 = ~pi899 & n57381;
  assign n58637 = ~n57529 & ~n58636;
  assign n58638 = pi1110 & ~n57381;
  assign n58639 = ~pi900 & n57381;
  assign n58640 = ~n58638 & ~n58639;
  assign n58641 = pi1111 & ~n57381;
  assign n58642 = ~pi902 & n57381;
  assign n58643 = ~n58641 & ~n58642;
  assign n58644 = pi1121 & ~n57381;
  assign n58645 = ~pi903 & n57381;
  assign n58646 = ~n58644 & ~n58645;
  assign n58647 = ~pi904 & n57381;
  assign n58648 = ~n57383 & ~n58647;
  assign n58649 = ~pi905 & n57381;
  assign n58650 = ~n57382 & ~n58649;
  assign n58651 = pi1128 & ~n57381;
  assign n58652 = ~pi906 & n57381;
  assign n58653 = ~n58651 & ~n58652;
  assign n58654 = ~pi908 & n57381;
  assign n58655 = ~n57432 & ~n58654;
  assign n58656 = pi1105 & ~n57381;
  assign n58657 = ~pi909 & n57381;
  assign n58658 = ~n58656 & ~n58657;
  assign n58659 = pi1117 & ~n57381;
  assign n58660 = ~pi910 & n57381;
  assign n58661 = ~n58659 & ~n58660;
  assign n58662 = pi1130 & ~n57381;
  assign n58663 = ~pi911 & n57381;
  assign n58664 = ~n58662 & ~n58663;
  assign n58665 = ~pi912 & n57381;
  assign n58666 = ~n57530 & ~n58665;
  assign n58667 = pi1106 & ~n57381;
  assign n58668 = ~pi913 & n57381;
  assign n58669 = ~n58667 & ~n58668;
  assign n58670 = pi1108 & ~n57381;
  assign n58671 = ~pi915 & n57381;
  assign n58672 = ~n58670 & ~n58671;
  assign n58673 = ~pi916 & n57381;
  assign n58674 = ~n57431 & ~n58673;
  assign n58675 = pi1112 & ~n57381;
  assign n58676 = ~pi917 & n57381;
  assign n58677 = ~n58675 & ~n58676;
  assign n58678 = pi1104 & ~n57381;
  assign n58679 = ~pi918 & n57381;
  assign n58680 = ~n58678 & ~n58679;
  assign n58681 = pi1102 & ~n57381;
  assign n58682 = ~pi919 & n57381;
  assign n58683 = ~n58681 & ~n58682;
  assign n58684 = pi1134 & n61413;
  assign n58685 = pi846 & ~n61413;
  assign n58686 = ~n58684 & ~n58685;
  assign n58687 = pi861 & ~pi1093;
  assign n58688 = ~n45960 & ~n58687;
  assign n58689 = ~pi228 & ~n58688;
  assign n58690 = pi123 & ~pi861;
  assign n58691 = ~pi123 & ~pi1141;
  assign n58692 = pi228 & ~n58691;
  assign n58693 = pi228 & ~n58690;
  assign n58694 = ~n58691 & n58693;
  assign n58695 = ~n58690 & n58692;
  assign n58696 = ~n58689 & ~n61692;
  assign n58697 = pi1139 & n61413;
  assign n58698 = pi862 & ~n61413;
  assign n58699 = ~n58697 & ~n58698;
  assign n58700 = pi869 & ~pi1093;
  assign n58701 = ~n45930 & ~n58700;
  assign n58702 = ~pi228 & ~n58701;
  assign n58703 = pi123 & ~pi869;
  assign n58704 = ~pi123 & ~pi1140;
  assign n58705 = pi228 & ~n58704;
  assign n58706 = pi228 & ~n58703;
  assign n58707 = ~n58704 & n58706;
  assign n58708 = ~n58703 & n58705;
  assign n58709 = ~n58702 & ~n61693;
  assign n58710 = ~pi875 & ~pi1093;
  assign n58711 = ~n45939 & ~n58710;
  assign n58712 = ~pi228 & ~n58711;
  assign n58713 = pi123 & pi875;
  assign n58714 = ~pi123 & pi1136;
  assign n58715 = pi228 & ~n58714;
  assign n58716 = pi228 & ~n58713;
  assign n58717 = ~n58714 & n58716;
  assign n58718 = ~n58713 & n58715;
  assign po1031 = ~n58712 & ~n61694;
  assign n58720 = pi877 & ~pi1093;
  assign n58721 = ~n45972 & ~n58720;
  assign n58722 = ~pi228 & ~n58721;
  assign n58723 = pi123 & ~pi877;
  assign n58724 = ~pi123 & ~pi1138;
  assign n58725 = pi228 & ~n58724;
  assign n58726 = pi228 & ~n58723;
  assign n58727 = ~n58724 & n58726;
  assign n58728 = ~n58723 & n58725;
  assign n58729 = ~n58722 & ~n61695;
  assign n58730 = pi878 & ~pi1093;
  assign n58731 = ~n45957 & ~n58730;
  assign n58732 = ~pi228 & ~n58731;
  assign n58733 = pi123 & ~pi878;
  assign n58734 = ~pi123 & ~pi1137;
  assign n58735 = pi228 & ~n58734;
  assign n58736 = pi228 & ~n58733;
  assign n58737 = ~n58734 & n58736;
  assign n58738 = ~n58733 & n58735;
  assign n58739 = ~n58732 & ~n61696;
  assign n58740 = pi879 & ~pi1093;
  assign n58741 = ~n45963 & ~n58740;
  assign n58742 = ~pi228 & ~n58741;
  assign n58743 = pi123 & ~pi879;
  assign n58744 = ~pi123 & ~pi1135;
  assign n58745 = pi228 & ~n58744;
  assign n58746 = pi228 & ~n58743;
  assign n58747 = ~n58744 & n58746;
  assign n58748 = ~n58743 & n58745;
  assign n58749 = ~n58742 & ~n61697;
  assign n58750 = pi840 & ~n2794;
  assign n58751 = pi1196 & n2794;
  assign n58752 = ~n58750 & ~n58751;
  assign n58753 = pi849 & ~n2794;
  assign n58754 = pi1198 & n2794;
  assign n58755 = ~n58753 & ~n58754;
  assign n58756 = pi863 & ~n2794;
  assign n58757 = pi1199 & n2794;
  assign n58758 = ~n58756 & ~n58757;
  assign n58759 = pi864 & ~n2794;
  assign n58760 = pi1197 & n2794;
  assign n58761 = ~n58759 & ~n58760;
  assign po991 = pi946 & n2794;
  assign n58763 = pi1093 & pi1152;
  assign n58764 = pi922 & ~pi1093;
  assign n58765 = ~pi922 & ~pi1093;
  assign n58766 = pi1093 & ~pi1152;
  assign n58767 = ~n58765 & ~n58766;
  assign n58768 = ~n58763 & ~n58764;
  assign po1115 = ~pi782 & pi960;
  assign po1116 = ~pi230 & pi961;
  assign po1118 = ~pi782 & pi963;
  assign po1122 = ~pi230 & pi967;
  assign po1124 = ~pi230 & pi969;
  assign po1125 = ~pi782 & pi970;
  assign po1126 = ~pi230 & pi971;
  assign po1127 = ~pi782 & pi972;
  assign po1128 = ~pi230 & pi974;
  assign po1129 = ~pi782 & pi975;
  assign po1131 = ~pi230 & pi977;
  assign po1132 = ~pi782 & pi978;
  assign n58781 = n2463 | n2464;
  assign n58782 = n2467 | n2468;
  assign n58783 = n2473 | n2474;
  assign n58784 = n2480 | n2481;
  assign n58785 = n2484 | n2485;
  assign n58786 = n2487 | n2488;
  assign n58787 = n2496 | n2497;
  assign n58788 = n2499 | n2500;
  assign n58789 = n2505 | n2506;
  assign n58790 = n2509 | n2510;
  assign n58791 = n2511 | n2512;
  assign n58792 = n2513 | n2514;
  assign n58793 = n2517 | n2518;
  assign n58794 = n2522 | n2523;
  assign n58795 = n2524 | n2525;
  assign n58796 = n2534 | n2535;
  assign n58797 = n2546 | n2536 | n2545;
  assign n58798 = n2537 | n2538 | n2543 | n2544;
  assign n58799 = n2541 | n2542;
  assign n58800 = n2549 | n2550;
  assign n58801 = n2553 | n2551 | n2552;
  assign n58802 = n2563 | n2564;
  assign n58803 = n2566 | n2567;
  assign n58804 = n2570 | n2571;
  assign n58805 = n2576 | n2573 | n2575;
  assign n58806 = n2587 | n2584 | n2586;
  assign n58807 = n2590 | n2591;
  assign n58808 = n2594 | n2595;
  assign n58809 = n2602 | n2603;
  assign n58810 = n2605 | n2606;
  assign n58811 = n2608 | n2609;
  assign n58812 = n2624 | n2619 | n2623;
  assign n58813 = n2626 | n2627;
  assign n58814 = n2629 | n2630;
  assign n58815 = n2637 | n2638;
  assign n58816 = n2639 | n2640;
  assign n58817 = n2644 | n2645;
  assign n58818 = n2646 | n2647;
  assign n58819 = n2652 | n2648 | n2651;
  assign n58820 = n2649 | n2650;
  assign n58821 = n2654 | n2655;
  assign n58822 = n2663 | n2656 | n2662;
  assign n58823 = n2657 | n2658;
  assign n58824 = n2659 | n2660;
  assign n58825 = n2685 | n2686;
  assign n58826 = n2688 | n2689;
  assign n58827 = n2690 | n2691;
  assign n58828 = n2700 | n2701;
  assign n58829 = n2704 | n2705;
  assign n58830 = n2723 | n2724;
  assign n58831 = n2734 | n2735;
  assign n58832 = n2736 | n2737;
  assign n58833 = n2742 | n2738 | n2741;
  assign n58834 = n2739 | n2740;
  assign n58835 = n2748 | n2749;
  assign n58836 = n2759 | n2760;
  assign n58837 = n2762 | n2763;
  assign n58838 = n2799 | n2800;
  assign n58839 = n2809 | n2810;
  assign n58840 = n2812 | n2813;
  assign n58841 = n2814 | n2815;
  assign n58842 = n2818 | n2816 | n2817;
  assign n58843 = n2825 | n2826;
  assign n58844 = n2830 | n2831;
  assign n58845 = n2832 | n2833;
  assign n58846 = n2842 | n2843;
  assign n58847 = n2848 | n2849;
  assign n58848 = n2854 | n2855;
  assign n58849 = n2863 | n2864;
  assign n58850 = n2865 | n2866;
  assign n58851 = n2874 | n2875;
  assign n58852 = n2876 | n2877;
  assign n58853 = n2896 | ~n2897;
  assign n58854 = n2904 | n2905;
  assign n58855 = ~n2929 | n2925 | n2928;
  assign n58856 = n2936 | n2937;
  assign n58857 = n2941 | n2942;
  assign n58858 = n2943 | ~n2944;
  assign n58859 = n2948 | ~n2949;
  assign n58860 = n2955 | ~n2956;
  assign n58861 = n2970 | ~n2971;
  assign n58862 = n2975 | n2976;
  assign n58863 = n2981 | n2982;
  assign n58864 = n2992 | ~n2993;
  assign n58865 = ~n3017 | n3010 | ~n3016;
  assign n58866 = n3022 | ~n3023;
  assign n58867 = n3034 | ~n3035;
  assign n58868 = n3049 | ~n3050;
  assign n58869 = n3058 | ~n3059;
  assign n58870 = n3073 | ~n3074;
  assign n58871 = n3092 | n3088 | ~n3091;
  assign n58872 = n3113 | n3106 | n3112;
  assign n58873 = n3125 | n3121 | ~n3124;
  assign n58874 = n3134 | n3135;
  assign n58875 = n3145 | ~n3146;
  assign n58876 = n3169 | ~n3170;
  assign n58877 = n3178 | ~n3179;
  assign n58878 = n3184 | ~n3185;
  assign n58879 = n3194 | n3195;
  assign n58880 = n3202 | n3203;
  assign n58881 = n3206 | n3207;
  assign n58882 = n3222 | ~n3223;
  assign n58883 = n3234 | ~n3235;
  assign n58884 = n3240 | ~n3241;
  assign n58885 = ~n3256 | n3252 | ~n3255;
  assign n58886 = n3266 | ~n3267;
  assign n58887 = n3278 | ~n3279;
  assign n58888 = n3282 | ~n3283;
  assign n58889 = n3289 | n3290;
  assign n58890 = n3301 | n3302;
  assign n58891 = n3307 | ~n3308;
  assign n58892 = n3319 | ~n3320;
  assign n58893 = n3328 | ~n3329;
  assign n58894 = ~n3362 | n3349 | ~n3361;
  assign n58895 = n3376 | n3377;
  assign n58896 = n3382 | n3383;
  assign n58897 = n3387 | n3388;
  assign n58898 = n3397 | ~n3398;
  assign n58899 = n3406 | ~n3407;
  assign n58900 = n3449 | n3436 | n3448;
  assign n58901 = n3462 | n3463;
  assign n58902 = ~n3474 | n3470 | ~n3473;
  assign n58903 = n3488 | ~n3489;
  assign n58904 = n3497 | ~n3498;
  assign n58905 = n3503 | ~n3504;
  assign n58906 = n3521 | ~n3522;
  assign n58907 = n3527 | ~n3528;
  assign n58908 = n3539 | ~n3540;
  assign n58909 = n3545 | ~n3546;
  assign n58910 = n3581 | n3582;
  assign n58911 = n3583 | n3584;
  assign n58912 = n3589 | ~n3590;
  assign n58913 = n3595 | ~n3596;
  assign n58914 = n3601 | ~n3602;
  assign n58915 = n3607 | ~n3608;
  assign n58916 = n3616 | ~n3617;
  assign n58917 = n3625 | n3626;
  assign n58918 = n3640 | ~n3641;
  assign n58919 = n3642 | n3643;
  assign n58920 = n3652 | ~n3653;
  assign n58921 = n3661 | ~n3662;
  assign n58922 = n3676 | ~n3677;
  assign n58923 = n3695 | n3691 | ~n3694;
  assign n58924 = n3700 | ~n3701;
  assign n58925 = n3736 | n3737;
  assign n58926 = n3738 | n3739;
  assign n58927 = n3747 | n3748;
  assign n58928 = n3762 | ~n3763;
  assign n58929 = n3768 | ~n3769;
  assign n58930 = n3779 | ~n3780;
  assign n58931 = n3786 | ~n3787;
  assign n58932 = n3795 | ~n3796;
  assign n58933 = n3802 | n3803;
  assign n58934 = n3807 | n3808;
  assign n58935 = n3809 | n3810;
  assign n58936 = n3823 | ~n3824;
  assign n58937 = n3828 | ~n3829;
  assign n58938 = n3837 | n3838;
  assign n58939 = n3847 | n3848;
  assign n58940 = n3855 | n3856;
  assign n58941 = n3858 | n3859;
  assign n58942 = n3872 | n3873;
  assign n58943 = n3895 | ~n3896;
  assign n58944 = n3901 | n3902;
  assign n58945 = n3910 | n3911;
  assign n58946 = n3913 | n3914;
  assign n58947 = n3919 | n3920;
  assign n58948 = n3924 | n3925;
  assign n58949 = n3931 | n3932;
  assign n58950 = n4001 | n4002;
  assign n58951 = n4008 | n4009;
  assign n58952 = n4016 | n4017;
  assign n58953 = n4043 | n4044;
  assign n58954 = n4051 | n4052;
  assign n58955 = n4055 | n4056;
  assign n58956 = n4078 | ~n4079;
  assign n58957 = n4085 | ~n4086;
  assign n58958 = n4090 | ~n4091;
  assign n58959 = n4097 | ~n4098;
  assign n58960 = n4102 | ~n4103;
  assign n58961 = n4109 | ~n4110;
  assign n58962 = n4114 | ~n4115;
  assign n58963 = n4131 | n4124 | n4130;
  assign n58964 = n4136 | ~n4137;
  assign n58965 = n4150 | n4151;
  assign n58966 = n4156 | n4157;
  assign n58967 = n4162 | n4159 | n4161;
  assign n58968 = n4170 | n4171;
  assign n58969 = n4175 | n4176;
  assign n58970 = n4177 | n4178;
  assign n58971 = n4179 | n4180;
  assign n58972 = n4181 | n4182;
  assign n58973 = n4192 | n4189 | n4191;
  assign n58974 = n4198 | ~n4199;
  assign n58975 = n4206 | n4207;
  assign n58976 = n4218 | n4219;
  assign n58977 = n4220 | n4221;
  assign n58978 = n4224 | n4225;
  assign n58979 = n4256 | n4257;
  assign n58980 = n4311 | n4308 | n4310;
  assign n58981 = n4337 | n4338;
  assign n58982 = n4343 | n4344;
  assign n58983 = n4350 | n4351;
  assign n58984 = n4354 | n4355;
  assign n58985 = n4388 | ~n4389;
  assign n58986 = n4395 | n4396;
  assign n58987 = n4400 | ~n4401;
  assign n58988 = n4407 | ~n4408;
  assign n58989 = n4417 | n4418;
  assign n58990 = n4425 | n4426;
  assign n58991 = n4429 | n4430;
  assign n58992 = n4442 | n4443;
  assign n58993 = n4451 | ~n4452;
  assign n58994 = n4460 | ~n4461;
  assign n58995 = n4468 | ~n4469;
  assign n58996 = n4472 | n4473;
  assign n58997 = n4481 | ~n4482;
  assign n58998 = n4490 | ~n4491;
  assign n58999 = n4509 | n4502 | ~n4508;
  assign n59000 = n4514 | ~n4515;
  assign n59001 = n4523 | ~n4524;
  assign n59002 = n4542 | ~n4543;
  assign n59003 = n4548 | ~n4549;
  assign n59004 = n4576 | n4566 | n4575;
  assign n59005 = n4587 | ~n4588;
  assign n59006 = n4593 | ~n4594;
  assign n59007 = n4602 | ~n4603;
  assign n59008 = n4611 | ~n4612;
  assign n59009 = n4617 | ~n4618;
  assign n59010 = n4623 | ~n4624;
  assign n59011 = n4659 | n4656 | n4658;
  assign n59012 = n4668 | ~n4669;
  assign n59013 = n4711 | n4712;
  assign n59014 = n4719 | n4720;
  assign n59015 = n4725 | n4726;
  assign n59016 = n4743 | n4744;
  assign n59017 = n4746 | n4747;
  assign n59018 = n4762 | ~n4763;
  assign n59019 = n4767 | ~n4768;
  assign n59020 = n4773 | ~n4774;
  assign n59021 = n4780 | ~n4781;
  assign n59022 = n4803 | ~n4804;
  assign n59023 = n4810 | n4811;
  assign n59024 = n4817 | n4818;
  assign n59025 = n4843 | ~n4844;
  assign n59026 = n4852 | n4853;
  assign n59027 = n4862 | n4863;
  assign n59028 = n4873 | ~n4874;
  assign n59029 = ~n4909 | n4905 | n4908;
  assign n59030 = n4954 | n4955;
  assign n59031 = n4975 | n4976;
  assign n59032 = n4979 | n4980;
  assign n59033 = n4995 | n4996;
  assign n59034 = n5044 | n5045;
  assign n59035 = n5046 | n5047;
  assign n59036 = n5058 | ~n5059;
  assign n59037 = n5067 | n5068;
  assign n59038 = n5080 | ~n5081;
  assign n59039 = n5106 | n5107;
  assign n59040 = n5116 | n5117;
  assign n59041 = n5124 | n5125;
  assign n59042 = n5153 | n5154;
  assign n59043 = n5163 | n5164;
  assign n59044 = n5165 | n5166;
  assign n59045 = n5178 | n5179;
  assign n59046 = n5180 | n5181;
  assign n59047 = n5192 | n5193;
  assign n59048 = n5217 | ~n5218;
  assign n59049 = n5222 | n5223;
  assign n59050 = n5228 | n5229;
  assign n59051 = n5232 | n5233;
  assign n59052 = n5244 | n5245;
  assign n59053 = n5253 | n5254;
  assign n59054 = n5264 | n5265;
  assign n59055 = n5270 | n5271;
  assign n59056 = n5274 | n5275;
  assign n59057 = n5283 | n5284;
  assign n59058 = n5296 | n5297;
  assign n59059 = n5337 | n5333 | ~n5336;
  assign n59060 = n5340 | n5341;
  assign n59061 = n5348 | n5349;
  assign n59062 = n5353 | n5354;
  assign n59063 = n5408 | n5409;
  assign n59064 = n5419 | n5420;
  assign n59065 = n5429 | ~n5430;
  assign n59066 = n5441 | ~n5442;
  assign n59067 = n5469 | ~n5470;
  assign n59068 = n5476 | n5477;
  assign n59069 = n5484 | n5485;
  assign n59070 = n5490 | n5487 | n5489;
  assign n59071 = n5522 | n5523;
  assign n59072 = n5528 | n5529;
  assign n59073 = n5532 | n5533;
  assign n59074 = n5563 | n5564;
  assign n59075 = n5571 | n5572;
  assign n59076 = n5579 | ~n5580;
  assign n59077 = n5584 | n5585;
  assign n59078 = n5591 | n5592;
  assign n59079 = n5596 | n5597;
  assign n59080 = n5623 | n5624;
  assign n59081 = n5629 | n5630;
  assign n59082 = n5641 | n5642;
  assign n59083 = n5647 | n5648;
  assign n59084 = n5653 | n5650 | n5652;
  assign n59085 = n5664 | ~n5665;
  assign n59086 = n5706 | n5707;
  assign n59087 = n5712 | n5709 | n5711;
  assign n59088 = n5719 | n5720;
  assign n59089 = n5752 | n5753;
  assign n59090 = n5758 | n5759;
  assign n59091 = n5760 | ~n5761;
  assign n59092 = n5780 | n5781;
  assign n59093 = n5786 | n5787;
  assign n59094 = n5792 | n5789 | n5791;
  assign n59095 = n5803 | ~n5804;
  assign n59096 = n5841 | n5842;
  assign n59097 = n5847 | n5848;
  assign n59098 = n5850 | n5851;
  assign n59099 = n5878 | n5879;
  assign n59100 = n5886 | n5887;
  assign n59101 = n5917 | n5918;
  assign n59102 = n5925 | n5926;
  assign n59103 = n5933 | ~n5934;
  assign n59104 = n5938 | n5939;
  assign n59105 = n5945 | n5946;
  assign n59106 = n5950 | n5951;
  assign n59107 = n5999 | ~n6000;
  assign n59108 = n6006 | n6007;
  assign n59109 = n6030 | n6031;
  assign n59110 = n6036 | n6033 | n6035;
  assign n59111 = n6051 | n6052;
  assign n59112 = n6085 | n6082 | n6084;
  assign n59113 = n6095 | n6096;
  assign n59114 = n6120 | ~n6121;
  assign n59115 = n6128 | n6129;
  assign n59116 = n6133 | n6134;
  assign n59117 = n6135 | n6136;
  assign n59118 = n6140 | n6141;
  assign n59119 = n6146 | n6147;
  assign n59120 = n6150 | n6151;
  assign n59121 = n6169 | n6170;
  assign n59122 = n6204 | n6205;
  assign n59123 = n6209 | n6210;
  assign n59124 = n6213 | n6214;
  assign n59125 = n6229 | n6230;
  assign n59126 = n6237 | n6238;
  assign n59127 = n6242 | n6243;
  assign n59128 = n6244 | ~n6245;
  assign n59129 = n6249 | ~n6250;
  assign n59130 = n6284 | n6285;
  assign n59131 = n6287 | n6288;
  assign n59132 = n6312 | n6313;
  assign n59133 = n6330 | n6331;
  assign n59134 = n6339 | n6340;
  assign n59135 = n6341 | n6342;
  assign n59136 = n6344 | n6345;
  assign n59137 = n6349 | n6347 | n6348;
  assign n59138 = n6352 | n6350 | n6351;
  assign n59139 = n6363 | n6364;
  assign n59140 = n6367 | n6368;
  assign n59141 = n6387 | n6388;
  assign n59142 = n6397 | n6398;
  assign n59143 = n6413 | n6414;
  assign n59144 = n6417 | n6418;
  assign n59145 = n6432 | n6433;
  assign n59146 = n6441 | n6442;
  assign n59147 = n6457 | ~n6458;
  assign n59148 = n6494 | n6495;
  assign n59149 = n6536 | ~n6537;
  assign n59150 = n6541 | ~n6542;
  assign n59151 = n6573 | ~n6574;
  assign n59152 = n6582 | n6583;
  assign n59153 = n6601 | n6602;
  assign n59154 = n6619 | ~n6620;
  assign n59155 = n6623 | n6624;
  assign n59156 = n6642 | n6643;
  assign n59157 = n6681 | ~n6682;
  assign n59158 = n6717 | n6714 | n6716;
  assign n59159 = n6738 | n6739;
  assign n59160 = n6750 | ~n6751;
  assign n59161 = n6762 | n6759 | n6761;
  assign n59162 = n6776 | ~n6777;
  assign n59163 = n6781 | ~n6782;
  assign n59164 = n6786 | ~n6787;
  assign n59165 = n6807 | ~n6808;
  assign n59166 = n6812 | ~n6813;
  assign n59167 = n6819 | n6820;
  assign n59168 = n6823 | n6824;
  assign n59169 = n6838 | n6839;
  assign n59170 = n6845 | n6846;
  assign n59171 = n6861 | n6862;
  assign n59172 = n6952 | n6953;
  assign n59173 = n6966 | ~n6967;
  assign n59174 = n6974 | ~n6975;
  assign n59175 = n6976 | n6977;
  assign n59176 = n6993 | ~n6994;
  assign n59177 = n6998 | ~n6999;
  assign n59178 = n7003 | ~n7004;
  assign n59179 = n7012 | ~n7013;
  assign n59180 = n7018 | n7019;
  assign n59181 = n7026 | n7027;
  assign n59182 = n7036 | n7037;
  assign n59183 = n7057 | n7058;
  assign n59184 = n7071 | ~n7072;
  assign n59185 = n7074 | n7075;
  assign n59186 = n7084 | n7085;
  assign n59187 = n7098 | n7099;
  assign n59188 = n7102 | n7103;
  assign n59189 = n7125 | n7126;
  assign n59190 = n7141 | n7142;
  assign n59191 = n7150 | n7151;
  assign n59192 = n7152 | n7153;
  assign n59193 = n7200 | n7201;
  assign n59194 = n7207 | n7208;
  assign n59195 = n7218 | ~n7219;
  assign n59196 = n7220 | n7221;
  assign n59197 = n7243 | n7244;
  assign n59198 = n7253 | ~n7254;
  assign n59199 = n7261 | ~n7262;
  assign n59200 = n7263 | n7264;
  assign n59201 = n7272 | n7273;
  assign n59202 = n7282 | ~n7283;
  assign n59203 = n7287 | ~n7288;
  assign n59204 = n7337 | n7338;
  assign n59205 = n7348 | n7349;
  assign n59206 = n7360 | n7361;
  assign n59207 = n7368 | n7365 | n7367;
  assign n59208 = n7373 | n7374;
  assign n59209 = n7386 | n7387;
  assign n59210 = n7390 | n7391;
  assign n59211 = n7396 | n7397;
  assign n59212 = n7414 | n7411 | n7413;
  assign n59213 = n7434 | n7435;
  assign n59214 = n7441 | n7442;
  assign n59215 = n7450 | n7451;
  assign n59216 = n7458 | ~n7459;
  assign n59217 = n7465 | n7466;
  assign n59218 = n7473 | n7474;
  assign n59219 = n7481 | ~n7482;
  assign n59220 = n7486 | ~n7487;
  assign n59221 = n7503 | n7504;
  assign n59222 = n7517 | n7518;
  assign n59223 = n7525 | n7526;
  assign n59224 = n7528 | n7529;
  assign n59225 = n7533 | n7534;
  assign n59226 = n7542 | n7543;
  assign n59227 = n7579 | n7580;
  assign n59228 = n7584 | ~n7585;
  assign n59229 = n7631 | n7628 | n7630;
  assign n59230 = n7636 | ~n7637;
  assign n59231 = n7677 | n7674 | n7676;
  assign n59232 = n7682 | ~n7683;
  assign n59233 = n7721 | ~n7722;
  assign n59234 = n7767 | ~n7768;
  assign n59235 = n7840 | ~n7841;
  assign n59236 = n7860 | n7861;
  assign n59237 = n7924 | ~n7925;
  assign n59238 = n7930 | ~n7931;
  assign n59239 = n7935 | ~n7936;
  assign n59240 = n7966 | n7963 | n7965;
  assign n59241 = n8050 | n8051;
  assign n59242 = n8055 | ~n8056;
  assign n59243 = n8096 | n8097;
  assign n59244 = n8106 | ~n8107;
  assign n59245 = n8119 | n8120;
  assign n59246 = n8132 | ~n8133;
  assign n59247 = n8202 | n8203;
  assign n59248 = n8228 | n8229;
  assign n59249 = n8232 | n8230 | n8231;
  assign n59250 = n8239 | n8240;
  assign n59251 = n8255 | ~n8256;
  assign n59252 = n8291 | ~n8292;
  assign n59253 = n8327 | ~n8328;
  assign n59254 = n8363 | ~n8364;
  assign n59255 = n8398 | ~n8399;
  assign n59256 = n8438 | ~n8439;
  assign n59257 = n8503 | ~n8504;
  assign n59258 = n8523 | n8524;
  assign n59259 = n8574 | ~n8575;
  assign n59260 = n8580 | ~n8581;
  assign n59261 = n8585 | ~n8586;
  assign n59262 = n8681 | n8682;
  assign n59263 = n8719 | n8720;
  assign n59264 = n8732 | n8733;
  assign n59265 = n8745 | ~n8746;
  assign n59266 = n8797 | n8798;
  assign n59267 = n8799 | ~n8800;
  assign n59268 = n8811 | ~n8812;
  assign n59269 = n8816 | ~n8817;
  assign n59270 = n8835 | ~n8836;
  assign n59271 = n8847 | ~n8848;
  assign n59272 = n8854 | n8855;
  assign n59273 = n8885 | ~n8886;
  assign n59274 = n8897 | ~n8898;
  assign n59275 = n8912 | n8913;
  assign n59276 = n8918 | ~n8919;
  assign n59277 = n8929 | ~n8930;
  assign n59278 = n8934 | ~n8935;
  assign n59279 = n8956 | n8957;
  assign n59280 = n8997 | n8998;
  assign n59281 = n9000 | n9001;
  assign n59282 = n9005 | ~n9006;
  assign n59283 = n9028 | n9026 | n9027;
  assign n59284 = n9058 | n9059;
  assign n59285 = n9076 | n9077;
  assign n59286 = n9086 | n9087;
  assign n59287 = n9090 | n9091;
  assign n59288 = n9120 | n9121;
  assign n59289 = n9163 | n9164;
  assign n59290 = n9175 | n9176;
  assign n59291 = n9187 | n9188;
  assign n59292 = n9190 | n9191;
  assign n59293 = n9200 | n9201;
  assign n59294 = n9219 | n9220;
  assign n59295 = n9227 | n9228;
  assign n59296 = n9284 | ~n9285;
  assign n59297 = n9320 | ~n9321;
  assign n59298 = n9355 | ~n9356;
  assign n59299 = n9395 | ~n9396;
  assign n59300 = n9422 | ~n9423;
  assign n59301 = n9463 | ~n9464;
  assign n59302 = n9483 | n9484;
  assign n59303 = n9541 | ~n9542;
  assign n59304 = n9550 | n9551;
  assign n59305 = n9556 | n9557;
  assign n59306 = ~n9605 | n9602 | n9604;
  assign n59307 = n9635 | n9636;
  assign n59308 = n9646 | ~n9647;
  assign n59309 = n9653 | n9654;
  assign n59310 = n9685 | ~n9686;
  assign n59311 = n9691 | ~n9692;
  assign n59312 = n9698 | ~n9699;
  assign n59313 = n9734 | ~n9735;
  assign n59314 = n9740 | ~n9741;
  assign n59315 = n9753 | ~n9754;
  assign n59316 = n9784 | n9785;
  assign n59317 = n9806 | n9807;
  assign n59318 = n9816 | n9817;
  assign n59319 = n9818 | n9819;
  assign n59320 = n9823 | n9824;
  assign n59321 = n9874 | ~n9875;
  assign n59322 = n9910 | ~n9911;
  assign n59323 = n9946 | ~n9947;
  assign n59324 = n9981 | ~n9982;
  assign n59325 = n10021 | ~n10022;
  assign n59326 = n10086 | ~n10087;
  assign n59327 = n10106 | n10107;
  assign n59328 = n10157 | ~n10158;
  assign n59329 = n10163 | ~n10164;
  assign n59330 = n10168 | ~n10169;
  assign n59331 = n10264 | n10265;
  assign n59332 = n10302 | n10303;
  assign n59333 = n10315 | n10316;
  assign n59334 = n10328 | ~n10329;
  assign n59335 = n10399 | n10400;
  assign n59336 = n10415 | n10416;
  assign n59337 = n10445 | ~n10446;
  assign n59338 = n10479 | ~n10480;
  assign n59339 = n10506 | ~n10507;
  assign n59340 = n10540 | ~n10541;
  assign n59341 = n10575 | ~n10576;
  assign n59342 = n10615 | ~n10616;
  assign n59343 = n10680 | ~n10681;
  assign n59344 = n10700 | n10701;
  assign n59345 = n10726 | n10727;
  assign n59346 = n10734 | n10735;
  assign n59347 = n10746 | n10747;
  assign n59348 = n10750 | n10751;
  assign n59349 = n10767 | ~n10768;
  assign n59350 = n10783 | n10784;
  assign n59351 = n10787 | n10788;
  assign n59352 = n10793 | n10794;
  assign n59353 = n10867 | ~n10868;
  assign n59354 = n10892 | n10893;
  assign n59355 = n10900 | n10901;
  assign n59356 = n10903 | n10904;
  assign n59357 = n10910 | n10907 | n10909;
  assign n59358 = n10927 | n10928;
  assign n59359 = n10990 | ~n10991;
  assign n59360 = n10995 | ~n10996;
  assign n59361 = n11001 | ~n11002;
  assign n59362 = n11024 | n11025;
  assign n59363 = n11035 | ~n11036;
  assign n59364 = n11041 | ~n11042;
  assign n59365 = n11060 | ~n11061;
  assign n59366 = n11066 | ~n11067;
  assign n59367 = n11119 | ~n11120;
  assign n59368 = n11125 | ~n11126;
  assign n59369 = n11134 | ~n11135;
  assign n59370 = n11143 | n11144;
  assign n59371 = n11145 | n11146;
  assign n59372 = n11185 | n11186;
  assign n59373 = n11192 | n11193;
  assign n59374 = n11272 | n11273;
  assign n59375 = n11347 | ~n11348;
  assign n59376 = n11353 | ~n11354;
  assign n59377 = n11359 | n11360;
  assign n59378 = n11454 | n11455;
  assign n59379 = n11478 | n11475 | n11477;
  assign n59380 = n11496 | n11497;
  assign n59381 = n11550 | ~n11551;
  assign n59382 = n11555 | ~n11556;
  assign n59383 = n11561 | ~n11562;
  assign n59384 = n11584 | n11585;
  assign n59385 = n11595 | ~n11596;
  assign n59386 = n11601 | ~n11602;
  assign n59387 = n11620 | ~n11621;
  assign n59388 = n11626 | ~n11627;
  assign n59389 = n11679 | ~n11680;
  assign n59390 = n11685 | ~n11686;
  assign n59391 = n11694 | ~n11695;
  assign n59392 = n11703 | n11704;
  assign n59393 = n11705 | n11706;
  assign n59394 = n11740 | n11741;
  assign n59395 = n11747 | n11748;
  assign n59396 = n11827 | n11828;
  assign n59397 = n11901 | ~n11902;
  assign n59398 = n11907 | ~n11908;
  assign n59399 = n11913 | n11914;
  assign n59400 = n12008 | n12009;
  assign n59401 = n12032 | n12029 | n12031;
  assign n59402 = n12049 | n12050;
  assign n59403 = n12101 | ~n12102;
  assign n59404 = n12168 | ~n12169;
  assign n59405 = n12173 | ~n12174;
  assign n59406 = n12179 | ~n12180;
  assign n59407 = n12207 | n12208;
  assign n59408 = n12226 | n12227;
  assign n59409 = n12321 | ~n12322;
  assign n59410 = n12334 | ~n12335;
  assign n59411 = n12399 | ~n12400;
  assign n59412 = n12419 | n12420;
  assign n59413 = n12431 | n12432;
  assign n59414 = n12438 | n12439;
  assign n59415 = n12446 | n12447;
  assign n59416 = n12511 | n12512;
  assign n59417 = n12526 | n12527;
  assign n59418 = n12550 | n12551;
  assign n59419 = n12557 | n12558;
  assign n59420 = n12563 | n12564;
  assign n59421 = n12584 | n12585;
  assign n59422 = n12605 | n12606;
  assign n59423 = n12616 | n12617;
  assign n59424 = n12661 | ~n12662;
  assign n59425 = n12667 | n12668;
  assign n59426 = n12708 | n12709;
  assign n59427 = n12772 | n12773;
  assign n59428 = n12796 | n12793 | n12795;
  assign n59429 = n12813 | n12814;
  assign n59430 = n12868 | ~n12869;
  assign n59431 = n12873 | ~n12874;
  assign n59432 = n12879 | ~n12880;
  assign n59433 = n12901 | n12897 | ~n12900;
  assign n59434 = n12915 | n12916;
  assign n59435 = n12987 | ~n12988;
  assign n59436 = n13009 | n13010;
  assign n59437 = n13013 | n13014;
  assign n59438 = n13016 | n13017;
  assign n59439 = n13020 | n13021;
  assign n59440 = n13025 | n13026;
  assign n59441 = n13028 | n13029;
  assign n59442 = n13048 | n13049;
  assign n59443 = n13067 | n13068;
  assign n59444 = n13083 | n13084;
  assign n59445 = n13148 | n13149;
  assign n59446 = n13164 | n13165;
  assign n59447 = n13215 | ~n13216;
  assign n59448 = n13221 | n13222;
  assign n59449 = n13262 | n13263;
  assign n59450 = n13326 | n13327;
  assign n59451 = n13350 | n13347 | n13349;
  assign n59452 = n13367 | n13368;
  assign n59453 = n13421 | ~n13422;
  assign n59454 = n13426 | ~n13427;
  assign n59455 = n13432 | ~n13433;
  assign n59456 = n13454 | n13450 | ~n13453;
  assign n59457 = n13468 | n13469;
  assign n59458 = n13531 | ~n13532;
  assign n59459 = n13553 | n13554;
  assign n59460 = n13557 | n13558;
  assign n59461 = n13560 | n13561;
  assign n59462 = n13564 | n13565;
  assign n59463 = n13569 | n13570;
  assign n59464 = n13572 | n13573;
  assign n59465 = n13597 | n13598;
  assign n59466 = n13601 | n13602;
  assign n59467 = n13666 | n13667;
  assign n59468 = n13682 | n13683;
  assign n59469 = n13692 | n13693;
  assign n59470 = n13738 | ~n13739;
  assign n59471 = n13744 | n13745;
  assign n59472 = n13785 | n13786;
  assign n59473 = n13849 | n13850;
  assign n59474 = n13873 | n13870 | n13872;
  assign n59475 = n13890 | n13891;
  assign n59476 = n13999 | ~n14000;
  assign n59477 = n14004 | ~n14005;
  assign n59478 = n14010 | ~n14011;
  assign n59479 = n14015 | ~n14016;
  assign n59480 = n14054 | n14055;
  assign n59481 = n14081 | ~n14082;
  assign n59482 = n14133 | n14134;
  assign n59483 = n14181 | n14182;
  assign n59484 = n14194 | ~n14195;
  assign n59485 = n14223 | n14224;
  assign n59486 = n14233 | ~n14234;
  assign n59487 = n14239 | ~n14240;
  assign n59488 = n14253 | ~n14254;
  assign n59489 = n14273 | n14274;
  assign n59490 = n14284 | n14285;
  assign n59491 = n14323 | ~n14324;
  assign n59492 = n14329 | n14330;
  assign n59493 = n14370 | n14371;
  assign n59494 = n14434 | n14435;
  assign n59495 = n14458 | n14455 | n14457;
  assign n59496 = n14475 | n14476;
  assign n59497 = n14528 | ~n14529;
  assign n59498 = n14533 | ~n14534;
  assign n59499 = n14539 | ~n14540;
  assign n59500 = n14560 | ~n14561;
  assign n59501 = n14572 | ~n14573;
  assign n59502 = n14578 | ~n14579;
  assign n59503 = n14597 | n14598;
  assign n59504 = n14652 | ~n14653;
  assign n59505 = n14674 | n14675;
  assign n59506 = n14678 | n14679;
  assign n59507 = n14713 | n14714;
  assign n59508 = n14720 | n14721;
  assign n59509 = n14799 | n14800;
  assign n59510 = n14815 | n14816;
  assign n59511 = n14866 | ~n14867;
  assign n59512 = n14872 | n14873;
  assign n59513 = n14913 | n14914;
  assign n59514 = n14977 | n14978;
  assign n59515 = n15001 | n14998 | n15000;
  assign n59516 = n15018 | n15019;
  assign n59517 = n15072 | ~n15073;
  assign n59518 = n15077 | ~n15078;
  assign n59519 = n15083 | ~n15084;
  assign n59520 = n15088 | ~n15089;
  assign n59521 = n15106 | ~n15107;
  assign n59522 = n15112 | ~n15113;
  assign n59523 = n15127 | n15128;
  assign n59524 = n15222 | n15223;
  assign n59525 = n15225 | n15226;
  assign n59526 = n15257 | ~n15258;
  assign n59527 = n15292 | n15293;
  assign n59528 = n15308 | n15309;
  assign n59529 = n15334 | ~n15335;
  assign n59530 = n15367 | n15368;
  assign n59531 = n15380 | ~n15381;
  assign n59532 = n15394 | ~n15395;
  assign n59533 = n15414 | n15415;
  assign n59534 = n15425 | n15426;
  assign n59535 = n15464 | ~n15465;
  assign n59536 = n15470 | n15471;
  assign n59537 = n15511 | n15512;
  assign n59538 = n15575 | n15576;
  assign n59539 = n15599 | n15596 | n15598;
  assign n59540 = n15616 | n15617;
  assign n59541 = n15669 | ~n15670;
  assign n59542 = n15674 | ~n15675;
  assign n59543 = n15680 | ~n15681;
  assign n59544 = n15701 | ~n15702;
  assign n59545 = n15713 | ~n15714;
  assign n59546 = n15719 | ~n15720;
  assign n59547 = n15794 | ~n15795;
  assign n59548 = n15816 | n15817;
  assign n59549 = n15820 | n15821;
  assign n59550 = n15855 | n15856;
  assign n59551 = n15862 | n15863;
  assign n59552 = n15941 | n15942;
  assign n59553 = n15957 | n15958;
  assign n59554 = n16005 | ~n16006;
  assign n59555 = n16011 | n16012;
  assign n59556 = n16052 | n16053;
  assign n59557 = n16116 | n16117;
  assign n59558 = n16140 | n16137 | n16139;
  assign n59559 = n16157 | n16158;
  assign n59560 = n16210 | ~n16211;
  assign n59561 = n16215 | ~n16216;
  assign n59562 = n16221 | ~n16222;
  assign n59563 = n16242 | ~n16243;
  assign n59564 = n16254 | ~n16255;
  assign n59565 = n16260 | ~n16261;
  assign n59566 = n16335 | ~n16336;
  assign n59567 = n16357 | n16358;
  assign n59568 = n16361 | n16362;
  assign n59569 = n16396 | n16397;
  assign n59570 = n16403 | n16404;
  assign n59571 = n16482 | n16483;
  assign n59572 = n16498 | n16499;
  assign n59573 = n16546 | ~n16547;
  assign n59574 = n16552 | n16553;
  assign n59575 = n16593 | n16594;
  assign n59576 = n16657 | n16658;
  assign n59577 = n16681 | n16678 | n16680;
  assign n59578 = n16698 | n16699;
  assign n59579 = n16751 | ~n16752;
  assign n59580 = n16756 | ~n16757;
  assign n59581 = n16762 | ~n16763;
  assign n59582 = n16783 | ~n16784;
  assign n59583 = n16795 | ~n16796;
  assign n59584 = n16801 | ~n16802;
  assign n59585 = n16820 | n16821;
  assign n59586 = n16875 | ~n16876;
  assign n59587 = n16897 | n16898;
  assign n59588 = n16901 | n16902;
  assign n59589 = n16936 | n16937;
  assign n59590 = n16943 | n16944;
  assign n59591 = n17022 | n17023;
  assign n59592 = n17038 | n17039;
  assign n59593 = n17086 | ~n17087;
  assign n59594 = n17092 | n17093;
  assign n59595 = n17133 | n17134;
  assign n59596 = n17197 | n17198;
  assign n59597 = n17221 | n17218 | n17220;
  assign n59598 = n17238 | n17239;
  assign n59599 = n17291 | ~n17292;
  assign n59600 = n17296 | ~n17297;
  assign n59601 = n17302 | ~n17303;
  assign n59602 = n17323 | ~n17324;
  assign n59603 = n17335 | ~n17336;
  assign n59604 = n17341 | ~n17342;
  assign n59605 = n17360 | n17361;
  assign n59606 = n17415 | ~n17416;
  assign n59607 = n17437 | n17438;
  assign n59608 = n17441 | n17442;
  assign n59609 = n17476 | n17477;
  assign n59610 = n17483 | n17484;
  assign n59611 = n17562 | n17563;
  assign n59612 = n17578 | n17579;
  assign n59613 = n17626 | ~n17627;
  assign n59614 = n17632 | n17633;
  assign n59615 = n17673 | n17674;
  assign n59616 = n17737 | n17738;
  assign n59617 = n17761 | n17758 | n17760;
  assign n59618 = n17778 | n17779;
  assign n59619 = n17831 | ~n17832;
  assign n59620 = n17836 | ~n17837;
  assign n59621 = n17842 | ~n17843;
  assign n59622 = n17863 | ~n17864;
  assign n59623 = n17875 | ~n17876;
  assign n59624 = n17881 | ~n17882;
  assign n59625 = n17900 | n17901;
  assign n59626 = n17955 | ~n17956;
  assign n59627 = n17977 | n17978;
  assign n59628 = n17981 | n17982;
  assign n59629 = n18016 | n18017;
  assign n59630 = n18023 | n18024;
  assign n59631 = n18102 | n18103;
  assign n59632 = n18118 | n18119;
  assign n59633 = n18166 | ~n18167;
  assign n59634 = n18172 | n18173;
  assign n59635 = n18213 | n18214;
  assign n59636 = n18277 | n18278;
  assign n59637 = n18301 | n18298 | n18300;
  assign n59638 = n18318 | n18319;
  assign n59639 = n18371 | ~n18372;
  assign n59640 = n18376 | ~n18377;
  assign n59641 = n18382 | ~n18383;
  assign n59642 = n18403 | ~n18404;
  assign n59643 = n18415 | ~n18416;
  assign n59644 = n18421 | ~n18422;
  assign n59645 = n18496 | ~n18497;
  assign n59646 = n18518 | n18519;
  assign n59647 = n18522 | n18523;
  assign n59648 = n18557 | n18558;
  assign n59649 = n18564 | n18565;
  assign n59650 = n18643 | n18644;
  assign n59651 = n18659 | n18660;
  assign n59652 = n18710 | ~n18711;
  assign n59653 = n18716 | n18717;
  assign n59654 = n18757 | n18758;
  assign n59655 = n18821 | n18822;
  assign n59656 = n18845 | n18842 | n18844;
  assign n59657 = n18862 | n18863;
  assign n59658 = n18970 | ~n18971;
  assign n59659 = n18975 | ~n18976;
  assign n59660 = n18981 | ~n18982;
  assign n59661 = n18986 | ~n18987;
  assign n59662 = n19028 | n19029;
  assign n59663 = n19049 | ~n19050;
  assign n59664 = n19084 | n19085;
  assign n59665 = n19100 | n19101;
  assign n59666 = n19148 | n19149;
  assign n59667 = n19161 | ~n19162;
  assign n59668 = n19190 | n19191;
  assign n59669 = n19200 | ~n19201;
  assign n59670 = n19206 | ~n19207;
  assign n59671 = n19220 | ~n19221;
  assign n59672 = n19240 | n19241;
  assign n59673 = n19251 | n19252;
  assign n59674 = n19293 | ~n19294;
  assign n59675 = n19299 | n19300;
  assign n59676 = n19340 | n19341;
  assign n59677 = n19404 | n19405;
  assign n59678 = n19428 | n19425 | n19427;
  assign n59679 = n19445 | n19446;
  assign n59680 = n19482 | ~n19483;
  assign n59681 = n19561 | ~n19562;
  assign n59682 = n19566 | ~n19567;
  assign n59683 = n19572 | ~n19573;
  assign n59684 = n19577 | ~n19578;
  assign n59685 = n19619 | n19620;
  assign n59686 = n19640 | ~n19641;
  assign n59687 = n19675 | n19676;
  assign n59688 = n19691 | n19692;
  assign n59689 = n19739 | n19740;
  assign n59690 = n19752 | ~n19753;
  assign n59691 = n19781 | n19782;
  assign n59692 = n19791 | ~n19792;
  assign n59693 = n19797 | ~n19798;
  assign n59694 = n19811 | ~n19812;
  assign n59695 = n19831 | n19832;
  assign n59696 = n19842 | n19843;
  assign n59697 = n19884 | ~n19885;
  assign n59698 = n19890 | n19891;
  assign n59699 = n19931 | n19932;
  assign n59700 = n19995 | n19996;
  assign n59701 = n20019 | n20016 | n20018;
  assign n59702 = n20036 | n20037;
  assign n59703 = n20073 | ~n20074;
  assign n59704 = n20152 | ~n20153;
  assign n59705 = n20157 | ~n20158;
  assign n59706 = n20163 | ~n20164;
  assign n59707 = n20168 | ~n20169;
  assign n59708 = n20210 | n20211;
  assign n59709 = n20231 | ~n20232;
  assign n59710 = n20266 | n20267;
  assign n59711 = n20282 | n20283;
  assign n59712 = n20330 | n20331;
  assign n59713 = n20343 | ~n20344;
  assign n59714 = n20372 | n20373;
  assign n59715 = n20382 | ~n20383;
  assign n59716 = n20388 | ~n20389;
  assign n59717 = n20402 | ~n20403;
  assign n59718 = n20422 | n20423;
  assign n59719 = n20433 | n20434;
  assign n59720 = n20440 | n20441;
  assign n59721 = n20447 | n20448;
  assign n59722 = n20455 | n20456;
  assign n59723 = n20527 | n20528;
  assign n59724 = n20551 | n20552;
  assign n59725 = n20558 | n20559;
  assign n59726 = n20564 | n20565;
  assign n59727 = n20590 | n20591;
  assign n59728 = n20650 | ~n20651;
  assign n59729 = n20720 | ~n20721;
  assign n59730 = n20725 | ~n20726;
  assign n59731 = n20731 | ~n20732;
  assign n59732 = n20736 | ~n20737;
  assign n59733 = n20775 | n20776;
  assign n59734 = n20794 | n20795;
  assign n59735 = n20863 | n20864;
  assign n59736 = n20911 | n20912;
  assign n59737 = n20924 | ~n20925;
  assign n59738 = n20958 | n20959;
  assign n59739 = n20965 | ~n20966;
  assign n59740 = n20979 | ~n20980;
  assign n59741 = n20999 | n21000;
  assign n59742 = n21010 | n21011;
  assign n59743 = n21052 | ~n21053;
  assign n59744 = n21058 | n21059;
  assign n59745 = n21099 | n21100;
  assign n59746 = n21163 | n21164;
  assign n59747 = n21187 | n21184 | n21186;
  assign n59748 = n21204 | n21205;
  assign n59749 = n21259 | ~n21260;
  assign n59750 = n21264 | ~n21265;
  assign n59751 = n21270 | ~n21271;
  assign n59752 = n21292 | n21288 | ~n21291;
  assign n59753 = n21306 | n21307;
  assign n59754 = n21378 | ~n21379;
  assign n59755 = n21400 | n21401;
  assign n59756 = n21404 | n21405;
  assign n59757 = n21407 | n21408;
  assign n59758 = n21411 | n21412;
  assign n59759 = n21416 | n21417;
  assign n59760 = n21419 | n21420;
  assign n59761 = n21439 | n21440;
  assign n59762 = n21457 | n21458;
  assign n59763 = n21472 | n21473;
  assign n59764 = n21537 | n21538;
  assign n59765 = n21553 | n21554;
  assign n59766 = n21601 | ~n21602;
  assign n59767 = n21607 | n21608;
  assign n59768 = n21648 | n21649;
  assign n59769 = n21712 | n21713;
  assign n59770 = n21736 | n21733 | n21735;
  assign n59771 = n21753 | n21754;
  assign n59772 = n21808 | ~n21809;
  assign n59773 = n21813 | ~n21814;
  assign n59774 = n21819 | ~n21820;
  assign n59775 = n21841 | n21837 | ~n21840;
  assign n59776 = n21855 | n21856;
  assign n59777 = n21927 | ~n21928;
  assign n59778 = n21949 | n21950;
  assign n59779 = n21953 | n21954;
  assign n59780 = n21956 | n21957;
  assign n59781 = n21960 | n21961;
  assign n59782 = n21965 | n21966;
  assign n59783 = n21968 | n21969;
  assign n59784 = n21988 | n21989;
  assign n59785 = n22006 | n22007;
  assign n59786 = n22021 | n22022;
  assign n59787 = n22086 | n22087;
  assign n59788 = n22102 | n22103;
  assign n59789 = n22150 | ~n22151;
  assign n59790 = n22156 | n22157;
  assign n59791 = n22197 | n22198;
  assign n59792 = n22261 | n22262;
  assign n59793 = n22285 | n22282 | n22284;
  assign n59794 = n22302 | n22303;
  assign n59795 = n22357 | ~n22358;
  assign n59796 = n22362 | ~n22363;
  assign n59797 = n22368 | ~n22369;
  assign n59798 = n22390 | n22386 | ~n22389;
  assign n59799 = n22404 | n22405;
  assign n59800 = n22476 | ~n22477;
  assign n59801 = n22498 | n22499;
  assign n59802 = n22502 | n22503;
  assign n59803 = n22505 | n22506;
  assign n59804 = n22509 | n22510;
  assign n59805 = n22514 | n22515;
  assign n59806 = n22517 | n22518;
  assign n59807 = n22537 | n22538;
  assign n59808 = n22555 | n22556;
  assign n59809 = n22570 | n22571;
  assign n59810 = n22635 | n22636;
  assign n59811 = n22651 | n22652;
  assign n59812 = n22699 | ~n22700;
  assign n59813 = n22705 | n22706;
  assign n59814 = n22746 | n22747;
  assign n59815 = n22810 | n22811;
  assign n59816 = n22834 | n22831 | n22833;
  assign n59817 = n22851 | n22852;
  assign n59818 = n22904 | ~n22905;
  assign n59819 = n22909 | ~n22910;
  assign n59820 = n22915 | ~n22916;
  assign n59821 = n22936 | ~n22937;
  assign n59822 = n22948 | ~n22949;
  assign n59823 = n22954 | ~n22955;
  assign n59824 = n23022 | ~n23023;
  assign n59825 = n23044 | n23045;
  assign n59826 = n23048 | n23049;
  assign n59827 = n23087 | n23088;
  assign n59828 = n23090 | n23091;
  assign n59829 = n23170 | n23171;
  assign n59830 = n23186 | n23187;
  assign n59831 = n23228 | ~n23229;
  assign n59832 = n23233 | ~n23234;
  assign n59833 = n23239 | ~n23240;
  assign n59834 = n23244 | ~n23245;
  assign n59835 = n23262 | ~n23263;
  assign n59836 = n23268 | ~n23269;
  assign n59837 = n23381 | n23382;
  assign n59838 = n23385 | n23386;
  assign n59839 = n23406 | ~n23407;
  assign n59840 = n23441 | n23442;
  assign n59841 = n23457 | n23458;
  assign n59842 = n23483 | ~n23484;
  assign n59843 = n23530 | ~n23531;
  assign n59844 = n23541 | ~n23542;
  assign n59845 = n23554 | ~n23555;
  assign n59846 = n23591 | n23592;
  assign n59847 = n23595 | n23596;
  assign n59848 = n23636 | ~n23637;
  assign n59849 = n23642 | n23643;
  assign n59850 = n23683 | n23684;
  assign n59851 = n23747 | n23748;
  assign n59852 = n23771 | n23768 | n23770;
  assign n59853 = n23788 | n23789;
  assign n59854 = n23850 | ~n23851;
  assign n59855 = n23855 | ~n23856;
  assign n59856 = n23861 | ~n23862;
  assign n59857 = n23866 | ~n23867;
  assign n59858 = n23882 | ~n23883;
  assign n59859 = n23888 | ~n23889;
  assign n59860 = n23915 | ~n23916;
  assign n59861 = n23980 | n23981;
  assign n59862 = n24057 | n24058;
  assign n59863 = n24095 | ~n24096;
  assign n59864 = n24130 | n24131;
  assign n59865 = n24143 | ~n24144;
  assign n59866 = n24157 | ~n24158;
  assign n59867 = n24181 | n24182;
  assign n59868 = n24183 | ~n24184;
  assign n59869 = n24189 | ~n24190;
  assign n59870 = n24211 | n24212;
  assign n59871 = n24237 | ~n24238;
  assign n59872 = n24242 | ~n24243;
  assign n59873 = n24248 | ~n24249;
  assign n59874 = n24294 | ~n24295;
  assign n59875 = n24342 | ~n24343;
  assign n59876 = n24360 | n24361;
  assign n59877 = n24388 | n24389;
  assign n59878 = n24460 | n24461;
  assign n59879 = n24476 | n24477;
  assign n59880 = n24508 | ~n24509;
  assign po357 = n24513 | ~n24514;
  assign n59882 = n24518 | n24519;
  assign n59883 = n24541 | ~n24542;
  assign n59884 = n24546 | ~n24547;
  assign n59885 = n24552 | ~n24553;
  assign n59886 = n24557 | ~n24558;
  assign n59887 = n24563 | ~n24564;
  assign n59888 = n24640 | n24641;
  assign n59889 = n24647 | n24648;
  assign n59890 = n24669 | n24670;
  assign n59891 = n24752 | n24753;
  assign n59892 = n24754 | n24755;
  assign n59893 = n24763 | n24764;
  assign n59894 = n24768 | n24769;
  assign n59895 = n24787 | n24788;
  assign n59896 = n24802 | n24803;
  assign n59897 = n24819 | n24820;
  assign n59898 = n24823 | n24824;
  assign n59899 = n24844 | n24845;
  assign n59900 = n24848 | n24849;
  assign n59901 = n24867 | n24868;
  assign n59902 = n24877 | n24878;
  assign n59903 = n24920 | n24921;
  assign n59904 = n24927 | n24928;
  assign n59905 = n24931 | n24932;
  assign n59906 = n24954 | n24955;
  assign n59907 = n24991 | n24992;
  assign n59908 = n24998 | n24999;
  assign n59909 = n25005 | n25006;
  assign n59910 = n25009 | ~n25010;
  assign n59911 = n25035 | n25036;
  assign n59912 = n25050 | n25051;
  assign n59913 = n25056 | n25057;
  assign n59914 = n25059 | n25060;
  assign n59915 = n25084 | ~n25085;
  assign n59916 = n25104 | n25105;
  assign n59917 = n25109 | ~n25110;
  assign n59918 = n25115 | ~n25116;
  assign n59919 = n25140 | n25141;
  assign n59920 = n25147 | n25148;
  assign n59921 = n25177 | ~n25178;
  assign n59922 = n25197 | n25198;
  assign n59923 = n25202 | ~n25203;
  assign n59924 = n25208 | ~n25209;
  assign n59925 = n25219 | n25220;
  assign n59926 = n25225 | n25226;
  assign n59927 = n25236 | ~n25237;
  assign n59928 = n25258 | n25259;
  assign n59929 = n25260 | n25261;
  assign n59930 = n25278 | ~n25279;
  assign n59931 = n25284 | ~n25285;
  assign n59932 = n25295 | ~n25296;
  assign n59933 = n25310 | n25311;
  assign n59934 = n25350 | n25351;
  assign n59935 = n25360 | n25361;
  assign n59936 = n25370 | n25371;
  assign n59937 = n25397 | n25398;
  assign n59938 = n25401 | n25402;
  assign n59939 = n25410 | n25411;
  assign n59940 = n25417 | n25418;
  assign n59941 = n25480 | n25481;
  assign n59942 = n25484 | n25485;
  assign n59943 = n25575 | n25576;
  assign n59944 = n25584 | ~n25585;
  assign n59945 = n25656 | n25657;
  assign n59946 = n25691 | n25692;
  assign n59947 = n25720 | n25721;
  assign n59948 = n25725 | n25726;
  assign n59949 = n25728 | n25729;
  assign n59950 = n25747 | n25748;
  assign n59951 = n25749 | n25750;
  assign n59952 = n25757 | n25758;
  assign n59953 = n25779 | n25780;
  assign n59954 = n25785 | n25786;
  assign n59955 = n25811 | ~n25812;
  assign n59956 = n25817 | ~n25818;
  assign n59957 = n25827 | n25828;
  assign n59958 = n25849 | n25850;
  assign n59959 = n25868 | n25869;
  assign n59960 = n25879 | n25880;
  assign n59961 = n25895 | n25896;
  assign n59962 = n25917 | n25918;
  assign n59963 = n26000 | ~n26001;
  assign n59964 = n26012 | n26013;
  assign n59965 = n26036 | n26037;
  assign n59966 = n26109 | n26110;
  assign n59967 = n26164 | n26165;
  assign n59968 = n26186 | ~n26187;
  assign n59969 = n26212 | ~n26213;
  assign n59970 = n26227 | n26228;
  assign n59971 = n26238 | n26239;
  assign n59972 = n26241 | n26242;
  assign n59973 = n26292 | n26293;
  assign n59974 = n26299 | n26300;
  assign n59975 = n26306 | n26307;
  assign n59976 = n26315 | ~n26316;
  assign n59977 = n26357 | ~n26358;
  assign n59978 = n26369 | n26370;
  assign n59979 = n26377 | n26378;
  assign n59980 = n26381 | n26382;
  assign n59981 = n26406 | n26407;
  assign n59982 = n26408 | n26409;
  assign n59983 = n26441 | n26442;
  assign n59984 = n26481 | ~n26482;
  assign n59985 = n26487 | ~n26488;
  assign n59986 = n26509 | n26510;
  assign n59987 = n26531 | ~n26532;
  assign n59988 = n26539 | ~n26540;
  assign n59989 = n26550 | n26551;
  assign n59990 = n26553 | n26554;
  assign n59991 = n26585 | n26586;
  assign n59992 = n26616 | n26617;
  assign n59993 = n26622 | n26623;
  assign n59994 = n26628 | n26629;
  assign n59995 = n26656 | ~n26657;
  assign n59996 = n26669 | n26670;
  assign n59997 = n26715 | n26716;
  assign n59998 = n26796 | n26797;
  assign n59999 = n26811 | n26812;
  assign n60000 = n26828 | n26829;
  assign n60001 = n26834 | ~n26835;
  assign n60002 = n26901 | ~n26902;
  assign po379 = n26907 | ~n26908;
  assign n60004 = n26922 | n26923;
  assign n60005 = n27018 | n27019;
  assign n60006 = n27048 | n27049;
  assign n60007 = n27070 | ~n27071;
  assign n60008 = n27112 | ~n27113;
  assign n60009 = n27120 | n27121;
  assign n60010 = n27131 | n27132;
  assign n60011 = n27138 | n27139;
  assign n60012 = n27141 | n27142;
  assign n60013 = n27166 | n27167;
  assign n60014 = n27190 | n27191;
  assign n60015 = n27198 | n27199;
  assign n60016 = n27205 | n27206;
  assign n60017 = n27210 | n27211;
  assign n60018 = n27235 | ~n27236;
  assign n60019 = n27240 | ~n27241;
  assign n60020 = n27249 | ~n27250;
  assign n60021 = n27289 | n27290;
  assign n60022 = n27298 | n27299;
  assign n60023 = n27308 | n27309;
  assign n60024 = n27336 | n27337;
  assign n60025 = n27343 | n27344;
  assign n60026 = n27360 | n27361;
  assign n60027 = n27374 | n27375;
  assign n60028 = n27406 | n27407;
  assign n60029 = n27419 | n27420;
  assign n60030 = n27440 | n27441;
  assign n60031 = n27460 | n27461;
  assign n60032 = n27466 | n27467;
  assign n60033 = n27536 | n27537;
  assign n60034 = n27596 | ~n27597;
  assign po380 = n27602 | ~n27603;
  assign n60036 = n27629 | n27630;
  assign n60037 = n27643 | n27644;
  assign n60038 = n27664 | n27665;
  assign n60039 = n27705 | n27706;
  assign n60040 = n27711 | n27712;
  assign n60041 = n27720 | n27721;
  assign n60042 = n27735 | n27736;
  assign n60043 = n27741 | n27742;
  assign n60044 = n27750 | ~n27751;
  assign n60045 = n27797 | n27798;
  assign n60046 = n27808 | n27809;
  assign n60047 = n27816 | n27817;
  assign n60048 = n27820 | n27821;
  assign n60049 = n27822 | n27823;
  assign n60050 = n27840 | n27841;
  assign n60051 = n27870 | n27871;
  assign n60052 = n27909 | ~n27910;
  assign n60053 = n27915 | ~n27916;
  assign n60054 = n27924 | ~n27925;
  assign n60055 = n28007 | n28008;
  assign n60056 = n28017 | n28014 | n28016;
  assign n60057 = n28048 | n28049;
  assign n60058 = n28062 | n28063;
  assign n60059 = n28079 | n28080;
  assign n60060 = n28083 | ~n28084;
  assign n60061 = n28099 | n28100;
  assign n60062 = n28104 | n28105;
  assign n60063 = n28107 | n28108;
  assign n60064 = n28115 | n28116;
  assign n60065 = n28219 | n28220;
  assign n60066 = n28237 | n28238;
  assign n60067 = n28257 | n28258;
  assign n60068 = n28289 | n28284 | n28285;
  assign n60069 = n28286 | n28287;
  assign n60070 = n28290 | n28291;
  assign n60071 = n28297 | n28298;
  assign n60072 = n28304 | n28305;
  assign n60073 = n28315 | n28316;
  assign n60074 = n28329 | n28330;
  assign n60075 = n28331 | n28332;
  assign n60076 = n28350 | n28351;
  assign n60077 = n28395 | n28396;
  assign n60078 = n28402 | n28403;
  assign n60079 = n28491 | n28492;
  assign n60080 = n28502 | n28503;
  assign n60081 = n28512 | n28513;
  assign n60082 = n28521 | ~n28522;
  assign n60083 = n28530 | ~n28531;
  assign n60084 = n28536 | n28533 | n28535;
  assign n60085 = n28538 | n28539;
  assign n60086 = n28540 | n28541;
  assign n60087 = n28558 | ~n28559;
  assign n60088 = n28572 | ~n28573;
  assign n60089 = n28579 | n28580;
  assign n60090 = n28593 | n28591 | n28592;
  assign n60091 = n28614 | n28615;
  assign n60092 = n28617 | ~n28618;
  assign n60093 = n28658 | n28659;
  assign n60094 = n28671 | n28672;
  assign n60095 = n28680 | n28681;
  assign n60096 = n28687 | n28688;
  assign n60097 = n28731 | n28732;
  assign n60098 = n28771 | n28772;
  assign n60099 = n28781 | n28782;
  assign n60100 = n28783 | n28784;
  assign n60101 = n28817 | n28818;
  assign n60102 = n28826 | n28827;
  assign n60103 = n28830 | n28831;
  assign n60104 = n28836 | n28837;
  assign n60105 = n28856 | n28857;
  assign n60106 = n28912 | n28913;
  assign n60107 = n28915 | n28916;
  assign n60108 = n28922 | n28923;
  assign n60109 = n28925 | n28926;
  assign n60110 = n28930 | n28931;
  assign n60111 = n28982 | n28978 | n28981;
  assign n60112 = n28990 | n28986 | n28989;
  assign n60113 = n28999 | n29000;
  assign n60114 = n29043 | n29044;
  assign n60115 = n29047 | n29048;
  assign n60116 = n29058 | n29059;
  assign n60117 = n29101 | ~n29102;
  assign n60118 = n29133 | n29134;
  assign n60119 = n29137 | n29138;
  assign n60120 = n29144 | n29145;
  assign n60121 = n29148 | n29149;
  assign n60122 = n29186 | ~n29187;
  assign n60123 = n29237 | n29238;
  assign n60124 = n29282 | n29283;
  assign n60125 = n29291 | n29292;
  assign n60126 = n29309 | n29310;
  assign n60127 = n29334 | n29335;
  assign n60128 = n29360 | n29361;
  assign n60129 = n29422 | n29423;
  assign n60130 = n29435 | n29436;
  assign n60131 = n29443 | n29444;
  assign n60132 = n29468 | n29469;
  assign n60133 = n29480 | n29481;
  assign n60134 = n29496 | n29497;
  assign n60135 = n29500 | n29501;
  assign n60136 = n29525 | n29526;
  assign n60137 = n29570 | ~n29571;
  assign n60138 = n29578 | ~n29579;
  assign n60139 = n29596 | n29597;
  assign n60140 = n29603 | n29604;
  assign n60141 = n29618 | n29619;
  assign n60142 = n29620 | n29621;
  assign n60143 = n29639 | n29640;
  assign n60144 = n29646 | n29647;
  assign n60145 = n29648 | n29649;
  assign n60146 = n29663 | n29664;
  assign n60147 = n29667 | ~n29668;
  assign n60148 = n29705 | n29706;
  assign n60149 = n29723 | n29724;
  assign n60150 = n29765 | n29766;
  assign n60151 = n29786 | n29787;
  assign n60152 = n29789 | n29790;
  assign n60153 = n29829 | n29830;
  assign n60154 = n29834 | n29835;
  assign n60155 = n29837 | n29838;
  assign n60156 = n29841 | n29842;
  assign n60157 = n29847 | n29848;
  assign n60158 = n29852 | n29853;
  assign n60159 = n29862 | n29863;
  assign n60160 = n29865 | n29866;
  assign n60161 = n29872 | n29873;
  assign n60162 = n29875 | n29876;
  assign n60163 = n29896 | n29897;
  assign n60164 = n29916 | n29917;
  assign n60165 = n30011 | n30009 | n30010;
  assign n60166 = n30012 | n30013;
  assign n60167 = n30039 | n30040;
  assign n60168 = n30071 | n30068 | n30070;
  assign n60169 = n30081 | n30082;
  assign n60170 = n30095 | n30096;
  assign n60171 = n30101 | n30098 | n30100;
  assign n60172 = n30121 | n30122;
  assign n60173 = n30132 | n30133;
  assign n60174 = n30148 | n30149;
  assign n60175 = n30157 | n30158;
  assign n60176 = n30165 | n30166;
  assign n60177 = n30184 | n30185;
  assign n60178 = n30218 | ~n30219;
  assign n60179 = n30239 | ~n30240;
  assign n60180 = n30270 | n30271;
  assign n60181 = n30434 | n30435;
  assign n60182 = n30473 | n30474;
  assign n60183 = n30494 | n30495;
  assign n60184 = n30553 | n30554;
  assign n60185 = n30640 | n30641;
  assign n60186 = n30650 | n30651;
  assign n60187 = n30675 | n30676;
  assign n60188 = n30683 | n30684;
  assign n60189 = n30690 | n30691;
  assign n60190 = n30711 | n30712;
  assign n60191 = n30722 | n30723;
  assign n60192 = n30764 | n30765;
  assign n60193 = n30766 | n30767;
  assign n60194 = n30790 | n30791;
  assign n60195 = n30792 | n30793;
  assign n60196 = n30809 | n30810;
  assign n60197 = n30814 | n30815;
  assign n60198 = n30816 | n30817;
  assign n60199 = n30819 | n30820;
  assign n60200 = n30826 | n30827;
  assign n60201 = n30846 | n30847;
  assign n60202 = n30859 | n30860;
  assign n60203 = n30906 | n30904 | n30905;
  assign n60204 = n30934 | n30935;
  assign n60205 = n30939 | n30940;
  assign n60206 = n30945 | n30946;
  assign n60207 = n30953 | n30954;
  assign n60208 = n30997 | n30994 | n30996;
  assign n60209 = n31010 | n31011;
  assign n60210 = n31022 | n31023;
  assign n60211 = n31026 | n31027;
  assign n60212 = n31055 | n31052 | n31054;
  assign n60213 = n31062 | n31063;
  assign n60214 = n31070 | n31071;
  assign n60215 = n31079 | n31080;
  assign n60216 = n31082 | n31083;
  assign n60217 = n31089 | n31090;
  assign n60218 = n31095 | n31096;
  assign n60219 = n31104 | n31105;
  assign n60220 = n31110 | n31111;
  assign n60221 = n31124 | n31125;
  assign n60222 = n31136 | n31137;
  assign n60223 = n31147 | n31148;
  assign n60224 = n31149 | ~n31150;
  assign n60225 = n31192 | n31193;
  assign n60226 = n31206 | n31207;
  assign n60227 = n31218 | n31219;
  assign n60228 = n31252 | n31253;
  assign n60229 = n31255 | n31256;
  assign n60230 = n31295 | n31296;
  assign n60231 = n31304 | n31305;
  assign n60232 = n31312 | n31313;
  assign n60233 = n31325 | n31326;
  assign n60234 = n31333 | n31334;
  assign n60235 = n31363 | n31364;
  assign n60236 = n31368 | n31369;
  assign n60237 = n31370 | n31371;
  assign n60238 = n31403 | n31404;
  assign n60239 = n31494 | n31492 | n31493;
  assign n60240 = n31508 | n31509;
  assign n60241 = n31516 | ~n31517;
  assign n60242 = n31526 | n31527;
  assign n60243 = n31538 | n31539;
  assign n60244 = n31546 | n31547;
  assign n60245 = n31554 | n31555;
  assign n60246 = n31568 | n31569;
  assign n60247 = n31589 | n31590;
  assign n60248 = n31597 | n31591 | n31596;
  assign n60249 = n31594 | n31595;
  assign n60250 = n31600 | ~n31601;
  assign n60251 = n31632 | n31633;
  assign n60252 = n31674 | ~n31675;
  assign n60253 = n31761 | n31762;
  assign n60254 = n31777 | n31778;
  assign n60255 = n31795 | ~n31796;
  assign n60256 = n31914 | n31915;
  assign n60257 = n31933 | n31934;
  assign n60258 = n32379 | n32380;
  assign n60259 = n32472 | n32473;
  assign n60260 = n32489 | n32490;
  assign n60261 = n32491 | n32492;
  assign n60262 = n32501 | n32502;
  assign n60263 = n32504 | n32505;
  assign n60264 = n32543 | n32544;
  assign n60265 = n32561 | n32562;
  assign n60266 = n32567 | n32568;
  assign n60267 = n32590 | ~n32591;
  assign n60268 = n32629 | n32630;
  assign n60269 = n32653 | n32654;
  assign n60270 = n32659 | n32660;
  assign n60271 = n32674 | n32675;
  assign n60272 = n32739 | n32740;
  assign n60273 = n32745 | n32746;
  assign n60274 = n32760 | n32761;
  assign n60275 = n32811 | n32812;
  assign n60276 = n32826 | n32827;
  assign n60277 = n32875 | n32876;
  assign n60278 = n32877 | n32878;
  assign n60279 = n32913 | n32909 | n32912;
  assign n60280 = n32910 | n32911;
  assign n60281 = n32915 | n32916;
  assign n60282 = n32937 | n32935 | n32936;
  assign n60283 = n32961 | n32962;
  assign n60284 = n32968 | ~n32969;
  assign n60285 = n32984 | n32985;
  assign n60286 = n32998 | n32999;
  assign n60287 = n33017 | n33018;
  assign n60288 = n33036 | n33037;
  assign n60289 = n33042 | n33039 | n33041;
  assign n60290 = n33047 | n33048;
  assign n60291 = n33051 | n33052;
  assign n60292 = n33083 | n33084;
  assign n60293 = n33132 | n33133;
  assign n60294 = n33142 | n33143;
  assign n60295 = n33147 | n33148;
  assign n60296 = n33156 | n33157;
  assign n60297 = n33158 | ~n33159;
  assign n60298 = n33174 | n33175;
  assign n60299 = n33188 | n33189;
  assign n60300 = n33201 | n33202;
  assign n60301 = n33225 | n33226;
  assign n60302 = n33251 | n33248 | n33250;
  assign n60303 = n33285 | n33286;
  assign n60304 = n33330 | n33331;
  assign n60305 = n33336 | n33337;
  assign n60306 = n33375 | n33376;
  assign n60307 = n33383 | n33384;
  assign n60308 = n33395 | n33396;
  assign n60309 = n33418 | n33419;
  assign n60310 = n33431 | n33429 | n33430;
  assign n60311 = n33434 | n33435;
  assign n60312 = n33480 | n33481;
  assign n60313 = n33507 | n33508;
  assign n60314 = n33514 | n33515;
  assign n60315 = n33522 | n33523;
  assign n60316 = n33532 | n33533;
  assign n60317 = n33583 | n33584;
  assign n60318 = n33610 | n33611;
  assign n60319 = n33617 | n33618;
  assign n60320 = n33663 | n33664;
  assign n60321 = n33672 | n33673;
  assign n60322 = n33679 | n33680;
  assign n60323 = n33723 | n33724;
  assign n60324 = n33730 | n33731;
  assign n60325 = n33735 | n33736;
  assign n60326 = n33745 | n33746;
  assign n60327 = n33756 | n33757;
  assign n60328 = n33821 | n33822;
  assign n60329 = n33832 | n33830 | n33831;
  assign n60330 = n33841 | n33842;
  assign n60331 = n33870 | n33871;
  assign n60332 = n33882 | n33883;
  assign n60333 = n33903 | n33904;
  assign n60334 = n33919 | n33920;
  assign n60335 = n33925 | n33926;
  assign n60336 = n33962 | n33963;
  assign n60337 = n33970 | n33971;
  assign n60338 = n33982 | n33983;
  assign n60339 = n34005 | n34006;
  assign n60340 = n34018 | n34016 | n34017;
  assign n60341 = n34021 | n34022;
  assign n60342 = n34055 | n34056;
  assign n60343 = n34078 | n34079;
  assign n60344 = n34091 | n34089 | n34090;
  assign n60345 = n34094 | n34095;
  assign n60346 = n34147 | n34148;
  assign n60347 = n34153 | n34154;
  assign n60348 = n34191 | n34192;
  assign n60349 = n34199 | n34200;
  assign n60350 = n34231 | n34232;
  assign n60351 = n34254 | n34255;
  assign n60352 = n34261 | n34262;
  assign n60353 = n34310 | n34311;
  assign n60354 = n34333 | n34334;
  assign n60355 = n34339 | n34340;
  assign n60356 = n34362 | n34363;
  assign n60357 = n34371 | n34369 | n34370;
  assign n60358 = n34374 | n34375;
  assign n60359 = n34409 | n34410;
  assign n60360 = n34415 | n34416;
  assign n60361 = n34453 | n34454;
  assign n60362 = n34461 | n34462;
  assign n60363 = n34503 | n34504;
  assign n60364 = n34548 | n34549;
  assign n60365 = n34582 | n34583;
  assign n60366 = n34593 | n34594;
  assign n60367 = n34602 | n34603;
  assign n60368 = n34610 | n34611;
  assign n60369 = n34616 | n34617;
  assign n60370 = n34618 | n34619;
  assign n60371 = n34623 | n34624;
  assign n60372 = n34688 | n34689;
  assign n60373 = n34698 | n34699;
  assign n60374 = n34711 | n34712;
  assign n60375 = n34720 | n34721;
  assign n60376 = n34727 | n34728;
  assign n60377 = n34771 | n34772;
  assign n60378 = n34778 | n34779;
  assign n60379 = n34783 | n34784;
  assign n60380 = n34793 | n34794;
  assign n60381 = n34804 | n34805;
  assign n60382 = n34813 | n34814;
  assign n60383 = n34822 | n34823;
  assign n60384 = n34829 | n34830;
  assign n60385 = n34873 | n34874;
  assign n60386 = n34880 | n34881;
  assign n60387 = n34885 | n34886;
  assign n60388 = n34895 | n34896;
  assign n60389 = n34906 | n34907;
  assign n60390 = n34920 | n34921;
  assign n60391 = n34968 | n34969;
  assign n60392 = n34996 | n34997;
  assign n60393 = n35005 | n35006;
  assign n60394 = n35012 | n35013;
  assign n60395 = n35056 | n35057;
  assign n60396 = n35063 | n35064;
  assign n60397 = n35068 | n35069;
  assign n60398 = n35078 | n35079;
  assign n60399 = n35089 | n35090;
  assign n60400 = n35103 | n35104;
  assign n60401 = n35112 | n35113;
  assign n60402 = n35119 | n35120;
  assign n60403 = n35133 | n35134;
  assign n60404 = n35166 | n35167;
  assign n60405 = n35173 | n35174;
  assign n60406 = n35178 | n35179;
  assign n60407 = n35188 | n35189;
  assign n60408 = n35222 | n35223;
  assign n60409 = n35259 | n35260;
  assign n60410 = n35267 | n35268;
  assign n60411 = n35278 | n35279;
  assign n60412 = n35282 | n35280 | n35281;
  assign n60413 = n35284 | n35285;
  assign n60414 = n35293 | n35294;
  assign n60415 = n35297 | n35298;
  assign n60416 = n35310 | n35311;
  assign n60417 = n35323 | n35324;
  assign n60418 = n35336 | n35337;
  assign n60419 = n35349 | n35350;
  assign n60420 = n35359 | n35360;
  assign n60421 = n35375 | n35376;
  assign n60422 = n35383 | n35384;
  assign n60423 = n35396 | n35397;
  assign n60424 = n35409 | n35410;
  assign n60425 = n35419 | n35420;
  assign n60426 = n35435 | n35436;
  assign n60427 = n35446 | n35447;
  assign n60428 = n35526 | n35527;
  assign n60429 = n35557 | n35558;
  assign n60430 = n35562 | n35563;
  assign n60431 = n35577 | n35578;
  assign n60432 = n35579 | n35580;
  assign n60433 = n35584 | n35585;
  assign n60434 = n35588 | n55401;
  assign n60435 = n55407 | n35589 | n35590;
  assign n60436 = n35592 | n35593;
  assign n60437 = n35614 | n35615;
  assign n60438 = n35631 | n35632;
  assign n60439 = n35675 | n35676;
  assign n60440 = n35679 | n35680;
  assign n60441 = n35692 | n35693;
  assign n60442 = n35695 | n35696;
  assign n60443 = n35738 | n35739;
  assign n60444 = n35781 | n35782;
  assign n60445 = n35787 | n35784 | n35786;
  assign n60446 = n35794 | n35795;
  assign n60447 = n35807 | n35808;
  assign n60448 = n35818 | n35819;
  assign n60449 = n35833 | n35834;
  assign n60450 = n35836 | n35837;
  assign n60451 = n35854 | n35855;
  assign n60452 = n35859 | n35860;
  assign n60453 = n35869 | n35866 | n35868;
  assign n60454 = n35884 | n35885;
  assign n60455 = n35902 | n35903;
  assign n60456 = n35934 | n35935;
  assign n60457 = n35940 | n35937 | n35939;
  assign n60458 = n35956 | n35957;
  assign n60459 = n35962 | n35963;
  assign n60460 = n35974 | n35975;
  assign n60461 = n35980 | n35981;
  assign n60462 = n36030 | n36031;
  assign n60463 = n36047 | n36048;
  assign n60464 = n36066 | n36067;
  assign n60465 = n36072 | n36069 | n36071;
  assign n60466 = n36079 | n36080;
  assign n60467 = n36099 | n36096 | n36098;
  assign n60468 = n36112 | n36113;
  assign n60469 = n36115 | n36116;
  assign n60470 = n36132 | n36133;
  assign n60471 = n36138 | n36139;
  assign n60472 = n36152 | n36153;
  assign n60473 = n36170 | n36171;
  assign n60474 = n36198 | n36199;
  assign n60475 = n36206 | n36207;
  assign n60476 = n36212 | n36213;
  assign n60477 = n36222 | n36223;
  assign n60478 = n36239 | n36240;
  assign po231 = n36275 | n36276;
  assign n60480 = n36282 | n36283;
  assign n60481 = n36299 | n36300;
  assign n60482 = n36335 | n36336;
  assign n60483 = n36356 | n36357;
  assign n60484 = n36407 | n36408;
  assign n60485 = n36411 | n36412;
  assign n60486 = n36444 | n36445;
  assign n60487 = n36456 | n36457;
  assign n60488 = n36458 | n36459;
  assign n60489 = n36463 | n36464;
  assign n60490 = n36465 | n36466;
  assign n60491 = n36467 | n36468;
  assign n60492 = n36504 | n36505;
  assign n60493 = n36529 | n36530;
  assign n60494 = n36531 | n36532;
  assign n60495 = n36536 | n36537;
  assign n60496 = n36541 | n36542;
  assign n60497 = n36550 | n36551;
  assign n60498 = n36562 | n36563;
  assign n60499 = n36589 | n36590;
  assign n60500 = n36591 | n36592;
  assign n60501 = n36593 | n36594;
  assign n60502 = n36610 | n36611;
  assign n60503 = n36622 | n36623;
  assign n60504 = n36671 | n36672;
  assign n60505 = n36687 | n36683 | ~n36686;
  assign n60506 = n36698 | n36699;
  assign n60507 = n36701 | n36702;
  assign n60508 = n36707 | ~n36708;
  assign n60509 = n36764 | n36765;
  assign n60510 = n36788 | n36789;
  assign n60511 = n36872 | n36873;
  assign n60512 = n36879 | n36880;
  assign n60513 = n36884 | n36885;
  assign n60514 = n36911 | n36912;
  assign n60515 = n36940 | n36941;
  assign n60516 = n36945 | n36946;
  assign n60517 = n36974 | n36975;
  assign n60518 = n36983 | n36984;
  assign n60519 = n36988 | n36989;
  assign n60520 = n37031 | n37032;
  assign n60521 = n37077 | n37078;
  assign n60522 = n37104 | n37105;
  assign n60523 = n37131 | n37132;
  assign n60524 = n37137 | n37138;
  assign n60525 = n37163 | n37164;
  assign n60526 = n37170 | ~n37171;
  assign n60527 = n37179 | n37180;
  assign n60528 = n37208 | n37209;
  assign n60529 = n37212 | n37213;
  assign n60530 = n37216 | n37217;
  assign n60531 = n37234 | n37235;
  assign n60532 = n37246 | n37247;
  assign n60533 = n37284 | n37285;
  assign n60534 = n37311 | n37312;
  assign n60535 = n37329 | n37330;
  assign n60536 = n37345 | n37346;
  assign n60537 = n37353 | n37354;
  assign n60538 = n37357 | n37358;
  assign n60539 = n37369 | n37370;
  assign po223 = n37373 | n37374;
  assign n60541 = n37382 | n37383;
  assign n60542 = n37450 | n37451;
  assign n60543 = n37467 | n37468;
  assign n60544 = n37493 | n37494;
  assign n60545 = n37509 | n37510;
  assign n60546 = n37526 | n37527;
  assign n60547 = n37561 | n37562;
  assign n60548 = n37586 | n37587;
  assign n60549 = n37608 | n37609;
  assign n60550 = n37685 | n37686;
  assign n60551 = n37721 | n37722;
  assign n60552 = n37758 | n37759;
  assign n60553 = n37762 | n37763;
  assign n60554 = n37781 | n37782;
  assign n60555 = n37799 | n37800;
  assign n60556 = n37809 | n37810;
  assign n60557 = n37818 | n37816 | n37817;
  assign n60558 = n37872 | n37873;
  assign n60559 = n37887 | n37888;
  assign n60560 = n37897 | n37898;
  assign n60561 = n37903 | n37901 | n37902;
  assign n60562 = n37910 | n37904 | n37909;
  assign n60563 = n54696 | n37906 | n37908;
  assign n60564 = n37914 | n37915;
  assign n60565 = n37933 | n37934;
  assign n60566 = n37963 | n37964;
  assign n60567 = n37977 | n37978;
  assign po234 = n37995 | n37996;
  assign n60569 = n38050 | n38051;
  assign n60570 = n38054 | n38055;
  assign n60571 = n38069 | n38070;
  assign n60572 = n38078 | n38079;
  assign n60573 = n38090 | n38091;
  assign n60574 = n38108 | n38109;
  assign n60575 = n38126 | n38127;
  assign n60576 = n38138 | n38139;
  assign n60577 = n38169 | n38170;
  assign n60578 = n38195 | n38196;
  assign n60579 = n38234 | n38235;
  assign n60580 = n38237 | n38238;
  assign n60581 = n38249 | n38250;
  assign n60582 = n38251 | n38252;
  assign n60583 = n38287 | n38288;
  assign n60584 = n38332 | n38333;
  assign n60585 = n38352 | n38353;
  assign n60586 = n38356 | ~n38357;
  assign n60587 = n38363 | n38364;
  assign n60588 = n38390 | n38391;
  assign n60589 = n38396 | n38397;
  assign n60590 = n38421 | n38422;
  assign n60591 = n38476 | n38477;
  assign n60592 = n38533 | n38534;
  assign n60593 = n38548 | n38549;
  assign n60594 = n38590 | n38591;
  assign n60595 = n38592 | n38593;
  assign n60596 = n38626 | n38627;
  assign n60597 = n38666 | n38667;
  assign n60598 = n38692 | n38693;
  assign n60599 = n38696 | n38697;
  assign n60600 = n38743 | n38744;
  assign n60601 = n38748 | n38749;
  assign n60602 = n38756 | n38757;
  assign n60603 = n38768 | n38769;
  assign n60604 = n38773 | n38774;
  assign n60605 = n38778 | n38779;
  assign n60606 = n38782 | n38783;
  assign n60607 = n38871 | n38872;
  assign n60608 = n38879 | ~n38880;
  assign n60609 = n38893 | n38894;
  assign n60610 = n38908 | n38909;
  assign n60611 = n38927 | n38928;
  assign n60612 = n38948 | n38949;
  assign n60613 = n38959 | n38960;
  assign n60614 = n38975 | n38976;
  assign n60615 = n38980 | n38981;
  assign n60616 = n38983 | n38984;
  assign n60617 = n38989 | n38990;
  assign n60618 = n38996 | n38997;
  assign n60619 = n39026 | n39027;
  assign n60620 = n39037 | n39038;
  assign n60621 = n39048 | n39049;
  assign n60622 = n39091 | n39092;
  assign n60623 = n39093 | n39094;
  assign n60624 = n39095 | n39096;
  assign n60625 = n39098 | n39099;
  assign n60626 = n39103 | n39104;
  assign n60627 = n39116 | n39117;
  assign n60628 = n39129 | n39130;
  assign n60629 = n39145 | n39146;
  assign n60630 = n39153 | n39154;
  assign n60631 = n39170 | n39171;
  assign n60632 = n39198 | n39199;
  assign n60633 = n39208 | n39209;
  assign n60634 = n39231 | n39232;
  assign n60635 = n39340 | n39341;
  assign n60636 = n39353 | n39354;
  assign n60637 = n39362 | n39363;
  assign n60638 = n39367 | n39368;
  assign n60639 = n39440 | n39441;
  assign n60640 = n39466 | n39467;
  assign n60641 = n39476 | n39477;
  assign n60642 = n39503 | n39504;
  assign n60643 = n39532 | n39533;
  assign n60644 = n39538 | n39539;
  assign n60645 = n39553 | ~n39554;
  assign n60646 = n39563 | ~n39564;
  assign n60647 = n39599 | n39600;
  assign n60648 = n39618 | n39615 | n39617;
  assign n60649 = n39642 | n39643;
  assign n60650 = n39646 | n39647;
  assign n60651 = n39701 | n39702;
  assign n60652 = n39714 | n39715;
  assign n60653 = n39749 | n39750;
  assign n60654 = n39837 | n39838;
  assign n60655 = n39866 | n39867;
  assign n60656 = n39880 | n39881;
  assign n60657 = n39891 | n39892;
  assign n60658 = n39893 | n39894;
  assign n60659 = n39944 | n39945;
  assign n60660 = n40021 | n40022;
  assign n60661 = n40027 | n40028;
  assign n60662 = n40037 | n40038;
  assign n60663 = n40042 | n40043;
  assign n60664 = n40056 | n40057;
  assign n60665 = n40078 | n40079;
  assign n60666 = n40090 | n40091;
  assign n60667 = n40142 | n40143;
  assign n60668 = n40147 | n40148;
  assign n60669 = n40158 | n40159;
  assign n60670 = n40169 | n40170;
  assign n60671 = n40187 | n40188;
  assign n60672 = n40191 | n40192;
  assign n60673 = n40223 | n40224;
  assign n60674 = n40237 | n40238;
  assign n60675 = n40270 | ~n40271;
  assign n60676 = n40276 | n40277;
  assign n60677 = n40306 | n40301 | n40305;
  assign n60678 = n40343 | n40344;
  assign n60679 = n40352 | n40353;
  assign n60680 = n40357 | n40358;
  assign n60681 = n40384 | n40385;
  assign n60682 = n40401 | n40402;
  assign n60683 = n40438 | n40439;
  assign n60684 = n40462 | n40463;
  assign n60685 = n40504 | n40505;
  assign n60686 = n40513 | n40514;
  assign n60687 = n40553 | n40554;
  assign n60688 = n40575 | n40576;
  assign n60689 = n40594 | ~n40595;
  assign po252 = n40599 | n40600;
  assign n60691 = n40617 | n40618;
  assign n60692 = n40651 | n40652;
  assign n60693 = n40657 | n40658;
  assign n60694 = n40659 | n40660;
  assign n60695 = n40712 | n40713;
  assign n60696 = n40718 | n40719;
  assign n60697 = n40731 | n40728 | n40730;
  assign n60698 = n40753 | n40754;
  assign n60699 = n40758 | n40759;
  assign n60700 = n40838 | n40839;
  assign n60701 = n40846 | ~n40847;
  assign n60702 = n40908 | n40909;
  assign n60703 = n40944 | n40945;
  assign n60704 = n40974 | n40975;
  assign n60705 = n41023 | n41024;
  assign n60706 = n41088 | n41089;
  assign n60707 = n41092 | n41093;
  assign n60708 = n41101 | n41102;
  assign n60709 = n41149 | n41150;
  assign n60710 = n41188 | n41189;
  assign n60711 = n41213 | n41214;
  assign n60712 = n41222 | n41223;
  assign n60713 = n41261 | n41262;
  assign n60714 = n41307 | n41308;
  assign n60715 = n41326 | n41327;
  assign n60716 = n41354 | n41355;
  assign n60717 = n41376 | n41377;
  assign n60718 = n41488 | n41489;
  assign n60719 = n41577 | n41578;
  assign n60720 = n41597 | n41598;
  assign n60721 = n41616 | n41617;
  assign n60722 = n41642 | n41643;
  assign n60723 = n41654 | n41655;
  assign n60724 = n41685 | n41686;
  assign n60725 = n41730 | n41731;
  assign n60726 = n41747 | n41748;
  assign n60727 = n41755 | n41756;
  assign n60728 = n41826 | n41827;
  assign po158 = n41842 | n41843;
  assign n60730 = n41850 | n41851;
  assign n60731 = n41869 | n41870;
  assign n60732 = n41904 | n41905;
  assign n60733 = n41934 | n41935;
  assign n60734 = n41979 | n41980;
  assign n60735 = n41996 | n41997;
  assign n60736 = n42004 | n42005;
  assign n60737 = n42075 | n42076;
  assign po159 = n42091 | n42092;
  assign n60739 = n42098 | n42099;
  assign n60740 = n42114 | n42115;
  assign n60741 = n42138 | n42139;
  assign n60742 = n42203 | n42204;
  assign n60743 = n42247 | n42248;
  assign n60744 = n42331 | n42332;
  assign n60745 = n42351 | n42352;
  assign n60746 = n42370 | n42371;
  assign n60747 = n42406 | n42407;
  assign n60748 = n42436 | n42437;
  assign n60749 = n42481 | n42482;
  assign n60750 = n42498 | n42499;
  assign n60751 = n42506 | n42507;
  assign n60752 = n42577 | n42578;
  assign po161 = n42593 | n42594;
  assign n60754 = n42601 | n42602;
  assign n60755 = n42620 | n42621;
  assign n60756 = n42656 | n42657;
  assign n60757 = n42686 | n42687;
  assign n60758 = n42731 | n42732;
  assign n60759 = n42748 | n42749;
  assign n60760 = n42756 | n42757;
  assign n60761 = n42827 | n42828;
  assign po162 = n42843 | n42844;
  assign n60763 = n42902 | n42903;
  assign n60764 = n42923 | n42924;
  assign n60765 = n42956 | n42957;
  assign n60766 = n42980 | n42981;
  assign n60767 = n42989 | n42990;
  assign n60768 = n42995 | n42996;
  assign n60769 = n42998 | n42999;
  assign n60770 = n43041 | n43042;
  assign n60771 = n43100 | n43101;
  assign n60772 = n43107 | n43108;
  assign n60773 = n43131 | n43132;
  assign n60774 = n43155 | n43156;
  assign n60775 = n43167 | n43168;
  assign n60776 = n43185 | n43186;
  assign n60777 = n43273 | n43274;
  assign n60778 = n43287 | n43288;
  assign n60779 = n43301 | n43302;
  assign n60780 = n43326 | n43327;
  assign n60781 = n43332 | n43333;
  assign n60782 = n43350 | n43351;
  assign n60783 = n43369 | n43370;
  assign n60784 = n43405 | n43406;
  assign n60785 = n43435 | n43436;
  assign n60786 = n43439 | n43440;
  assign n60787 = n43485 | n43486;
  assign n60788 = n43510 | n43511;
  assign n60789 = n43512 | n43513;
  assign n60790 = n43585 | n43586;
  assign n60791 = n43605 | n43606;
  assign n60792 = n43626 | n43627;
  assign n60793 = n43646 | n43647;
  assign n60794 = n43669 | n43670;
  assign n60795 = n43749 | n43750;
  assign n60796 = n43770 | n43771;
  assign n60797 = n43843 | n43844;
  assign n60798 = n43861 | n43862;
  assign n60799 = n43882 | n43883;
  assign n60800 = n43897 | n43898;
  assign n60801 = n43997 | n43998;
  assign n60802 = n44018 | n44019;
  assign n60803 = n44095 | n44096;
  assign n60804 = n44141 | n44142;
  assign n60805 = n44162 | n44163;
  assign n60806 = n44229 | n44230;
  assign n60807 = n44317 | n44318;
  assign n60808 = n44393 | n44394;
  assign n60809 = n44464 | n44465;
  assign po471 = n44495 | n44496;
  assign po637 = n44535 | n44536;
  assign n60812 = n44591 | n44592;
  assign n60813 = n44669 | n44670;
  assign n60814 = n44681 | n44682;
  assign n60815 = n44690 | n44691;
  assign n60816 = n44699 | n44700;
  assign n60817 = n44702 | n44703;
  assign n60818 = n44743 | ~n44744;
  assign n60819 = n44757 | n44758;
  assign n60820 = n44781 | n44782;
  assign n60821 = n44846 | n44847;
  assign n60822 = n44882 | n44883;
  assign n60823 = n44893 | n44894;
  assign n60824 = n44954 | n44955;
  assign n60825 = n44958 | n44956 | n44957;
  assign n60826 = n44963 | n44964;
  assign n60827 = n44970 | n44971;
  assign n60828 = n44980 | n44981;
  assign n60829 = n45016 | n45017;
  assign n60830 = n45036 | n45033 | n45035;
  assign n60831 = n45044 | ~n45045;
  assign n60832 = n45057 | n45058;
  assign n60833 = n45061 | n45062;
  assign n60834 = n45075 | n45076;
  assign n60835 = n45078 | n45079;
  assign n60836 = n45082 | n45083;
  assign n60837 = n45089 | n45090;
  assign n60838 = n45101 | n45102;
  assign n60839 = n45103 | ~n45104;
  assign n60840 = n45106 | n45107;
  assign n60841 = n45116 | n45117;
  assign n60842 = n45118 | ~n45119;
  assign n60843 = n45122 | n45123;
  assign n60844 = n45125 | ~n45126;
  assign po497 = ~n45135 | n45131 | n45134;
  assign n60846 = n45197 | n45198;
  assign n60847 = n45450 | ~n45451;
  assign n60848 = n45460 | n45461;
  assign po211 = n45471 | n45472;
  assign n60850 = n45506 | n45507;
  assign n60851 = n45539 | n45540;
  assign n60852 = n45563 | n45564;
  assign n60853 = n45565 | n45566;
  assign n60854 = n45593 | n45594;
  assign n60855 = n45598 | n45595 | n45597;
  assign n60856 = n45619 | n45620;
  assign po220 = n45629 | n45630;
  assign po247 = n45642 | n45643;
  assign n60859 = n45647 | n45648;
  assign n60860 = n45649 | n45650;
  assign n60861 = n45653 | n45654;
  assign n60862 = n45692 | n45693;
  assign n60863 = n45695 | n45696;
  assign po206 = n45712 | n45713;
  assign n60865 = n45716 | n45714 | n45715;
  assign po213 = n45728 | n45729;
  assign n60867 = n45732 | n45733;
  assign po222 = n45751 | n45752;
  assign po225 = n45758 | n45759;
  assign n60870 = n45777 | n45778;
  assign n60871 = n45793 | n45794;
  assign n60872 = n45801 | n45802;
  assign n60873 = n45815 | n45816;
  assign n60874 = n45817 | n45818;
  assign po245 = n45820 | n45821;
  assign po261 = n45834 | n45835;
  assign po267 = n45836 | n45837;
  assign po209 = n45848 | n45849;
  assign n60879 = n45859 | n45860;
  assign n60880 = n45865 | n45866;
  assign n60881 = n45873 | n45874;
  assign n60882 = n45879 | n45880;
  assign n60883 = n45885 | n45886;
  assign po943 = n45922 | ~n45923;
  assign n60885 = n45928 | ~n45929;
  assign po1083 = n45937 | ~n45938;
  assign po1085 = n45946 | ~n45947;
  assign po1086 = n45952 | ~n45953;
  assign po1095 = n45970 | ~n45971;
  assign n60890 = n45979 | ~n45980;
  assign n60891 = n46000 | n46001;
  assign n60892 = n46012 | n46013;
  assign n60893 = n46014 | n46015;
  assign n60894 = n46021 | ~n46022;
  assign n60895 = n46039 | n46040;
  assign n60896 = n46044 | n46042 | n46043;
  assign n60897 = n46050 | ~n46051;
  assign n60898 = n46055 | n46056;
  assign n60899 = n46063 | n46064;
  assign n60900 = n46067 | n46068;
  assign n60901 = ~n46077 | n46074 | ~n46076;
  assign n60902 = n46106 | n46107;
  assign n60903 = n46134 | n46135;
  assign n60904 = n46204 | n46205;
  assign n60905 = n46206 | n46207;
  assign n60906 = n46222 | n46223;
  assign n60907 = n46315 | n46316;
  assign n60908 = n46349 | n50485;
  assign n60909 = n46366 | n46367;
  assign n60910 = n46409 | n46410;
  assign n60911 = n46412 | n46413;
  assign n60912 = n46432 | n46433;
  assign n60913 = n46441 | n46442;
  assign n60914 = n46466 | n46467;
  assign n60915 = n46469 | n46470;
  assign n60916 = n46493 | n46494;
  assign n60917 = n46529 | n46519 | n46528;
  assign n60918 = n46526 | n50713;
  assign n60919 = n46546 | n46547;
  assign n60920 = n46586 | n46587;
  assign n60921 = n46595 | n46596;
  assign n60922 = n46599 | n46600;
  assign n60923 = n46616 | n46617;
  assign n60924 = n46662 | n46663;
  assign n60925 = n46670 | n46671;
  assign n60926 = n46689 | n46690;
  assign n60927 = n46691 | n46692;
  assign n60928 = n46697 | n46698;
  assign n60929 = n46719 | n46720;
  assign n60930 = n46729 | n46730;
  assign n60931 = n46739 | n46740;
  assign n60932 = n46749 | n46750;
  assign n60933 = n46829 | n46830;
  assign n60934 = n46854 | n46855;
  assign n60935 = n46863 | n46860 | n46862;
  assign n60936 = n46875 | n46876;
  assign n60937 = n46906 | n46907;
  assign n60938 = n46909 | n46910;
  assign n60939 = n46925 | n46926;
  assign n60940 = n46943 | n46944;
  assign n60941 = n46972 | n46969 | n46971;
  assign n60942 = n46988 | n46989;
  assign n60943 = n47008 | n47009;
  assign n60944 = n47029 | n47030;
  assign n60945 = n47043 | n47044;
  assign n60946 = n47094 | n47095;
  assign n60947 = n47117 | n47118;
  assign n60948 = n47131 | n47132;
  assign n60949 = n47162 | n47163;
  assign n60950 = n47252 | n47253;
  assign n60951 = n47257 | n47258;
  assign n60952 = n47261 | ~n47262;
  assign n60953 = n47264 | n47265;
  assign n60954 = n47278 | n47279;
  assign n60955 = n47288 | n47289;
  assign n60956 = n47312 | n47313;
  assign n60957 = n47325 | n47326;
  assign n60958 = n47355 | n47356;
  assign n60959 = n47370 | n47371;
  assign n60960 = n47382 | n47383;
  assign n60961 = n47400 | n47401;
  assign n60962 = n47408 | n47409;
  assign n60963 = n47411 | n47412;
  assign n60964 = n47439 | ~n47440;
  assign n60965 = n47466 | n47467;
  assign n60966 = n47474 | n47475;
  assign n60967 = n47478 | n47479;
  assign n60968 = n47481 | n47482;
  assign n60969 = n47514 | n47515;
  assign n60970 = n47518 | n47519;
  assign n60971 = n47617 | n47618;
  assign n60972 = n47637 | n47638;
  assign n60973 = n47651 | n47652;
  assign n60974 = n47657 | n47658;
  assign n60975 = n47695 | n47696;
  assign n60976 = n47704 | n47705;
  assign n60977 = n47710 | n47711;
  assign n60978 = n47737 | n47738;
  assign n60979 = n47746 | n47747;
  assign n60980 = n47752 | n47753;
  assign n60981 = n47779 | n47780;
  assign n60982 = n47788 | n47789;
  assign n60983 = n47809 | n47810;
  assign n60984 = n47815 | n47816;
  assign n60985 = n47824 | n47825;
  assign n60986 = n47838 | n47839;
  assign n60987 = n47851 | n47852;
  assign n60988 = n47862 | n47863;
  assign n60989 = n47882 | n47883;
  assign n60990 = n47888 | n47889;
  assign n60991 = n47915 | n47916;
  assign n60992 = n47924 | n47925;
  assign n60993 = n47944 | n47945;
  assign n60994 = n47950 | n47951;
  assign n60995 = n47976 | n47977;
  assign n60996 = n47984 | n47985;
  assign n60997 = n47996 | n47997;
  assign n60998 = n48006 | n48007;
  assign n60999 = n48025 | n48026;
  assign n61000 = n48033 | ~n48034;
  assign n61001 = n48046 | n48047;
  assign n61002 = n48069 | n48070;
  assign n61003 = n48077 | ~n48078;
  assign n61004 = n48089 | n48090;
  assign n61005 = n48098 | n48099;
  assign n61006 = n48117 | n48118;
  assign n61007 = n48137 | n48138;
  assign n61008 = n48153 | ~n48154;
  assign n61009 = n48172 | n48173;
  assign n61010 = n48190 | n48191;
  assign n61011 = n48197 | n48198;
  assign n61012 = n48213 | n48214;
  assign n61013 = n48232 | n48233;
  assign n61014 = n48247 | ~n48248;
  assign n61015 = n48253 | n48254;
  assign n61016 = n48262 | n48263;
  assign n61017 = n48277 | n48278;
  assign n61018 = n48287 | n48288;
  assign n61019 = n48302 | n48303;
  assign n61020 = n48321 | n48322;
  assign n61021 = n48336 | ~n48337;
  assign n61022 = n48348 | n48349;
  assign n61023 = n48356 | n48357;
  assign n61024 = n48368 | n48369;
  assign n61025 = n48376 | n48377;
  assign n61026 = n48400 | n48401;
  assign n61027 = n48416 | n48417;
  assign n61028 = n48423 | n48424;
  assign n61029 = n48441 | ~n48442;
  assign n61030 = n48457 | n48458;
  assign n61031 = n48467 | n48468;
  assign n61032 = n48488 | n48489;
  assign n61033 = n48504 | n48505;
  assign n61034 = n48511 | n48512;
  assign n61035 = n48529 | ~n48530;
  assign n61036 = n48545 | n48546;
  assign n61037 = n48555 | n48556;
  assign n61038 = n48571 | n48572;
  assign n61039 = n48579 | n48580;
  assign n61040 = n48591 | n48592;
  assign n61041 = n48599 | n48600;
  assign n61042 = n48620 | ~n48621;
  assign n61043 = n48635 | n48636;
  assign n61044 = n48641 | n48642;
  assign n61045 = n48675 | n48676;
  assign n61046 = n48681 | n48682;
  assign n61047 = n48709 | n48710;
  assign n61048 = n48717 | n48718;
  assign n61049 = n48723 | n48724;
  assign n61050 = n48731 | n48732;
  assign n61051 = n48743 | n48744;
  assign n61052 = n48749 | n48750;
  assign n61053 = n48776 | n48777;
  assign n61054 = n48796 | n48797;
  assign n61055 = n48804 | n48805;
  assign n61056 = n48810 | n48811;
  assign n61057 = n48818 | n48819;
  assign n61058 = n48830 | n48831;
  assign n61059 = n48850 | n48851;
  assign n61060 = n48866 | n48867;
  assign n61061 = n48886 | n48887;
  assign n61062 = n48902 | n48903;
  assign n61063 = n48922 | n48923;
  assign n61064 = n48938 | n48939;
  assign n61065 = n48958 | n48959;
  assign n61066 = n48974 | n48975;
  assign n61067 = n48994 | n48995;
  assign po412 = n49016 | ~n49017;
  assign po413 = n49022 | ~n49023;
  assign po414 = n49028 | ~n49029;
  assign po415 = n49034 | ~n49035;
  assign po416 = n49040 | ~n49041;
  assign po447 = n49052 | ~n49053;
  assign po448 = n49058 | ~n49059;
  assign po449 = n49064 | ~n49065;
  assign po450 = n49070 | ~n49071;
  assign po451 = n49076 | ~n49077;
  assign po452 = n49082 | ~n49083;
  assign po453 = n49088 | ~n49089;
  assign po454 = n49094 | ~n49095;
  assign n61081 = n49111 | n49112;
  assign n61082 = n49127 | n49128;
  assign n61083 = n49134 | n49135;
  assign n61084 = n49248 | n49249;
  assign n61085 = n49259 | n49260;
  assign n61086 = n49273 | n49274;
  assign n61087 = n49291 | n49292;
  assign n61088 = n49309 | n49310;
  assign n61089 = n49315 | n50173;
  assign n61090 = n49317 | ~n49318;
  assign n61091 = n49331 | n49332;
  assign n61092 = n49353 | ~n49354;
  assign n61093 = n49356 | n49357;
  assign n61094 = n49418 | n49419;
  assign n61095 = n49433 | n49430 | n49432;
  assign n61096 = n49436 | n49437;
  assign n61097 = n49441 | ~n49442;
  assign n61098 = n49443 | n49444;
  assign n61099 = n49470 | n49467 | n49469;
  assign n61100 = n49479 | n49480;
  assign n61101 = n49481 | n49482;
  assign n61102 = n49486 | n49487;
  assign n61103 = n49501 | n49502;
  assign n61104 = n49509 | ~n49510;
  assign n61105 = n49513 | n49514;
  assign n61106 = n49522 | n49523;
  assign n61107 = n49530 | n49531;
  assign n61108 = n49554 | n49555;
  assign n61109 = n49578 | n49579;
  assign n61110 = n49604 | n49605;
  assign n61111 = n49612 | n49613;
  assign n61112 = n49616 | n49617;
  assign n61113 = n49626 | n49627;
  assign n61114 = n49635 | n49636;
  assign n61115 = n49637 | n49638;
  assign n61116 = n49644 | n49645;
  assign n61117 = n49652 | ~n49653;
  assign n61118 = n49698 | n49699;
  assign n61119 = n49710 | n49711;
  assign n61120 = n49734 | n49735;
  assign n61121 = n49741 | n49742;
  assign n61122 = n49755 | n49756;
  assign n61123 = n49757 | n49758;
  assign n61124 = n49764 | n49765;
  assign n61125 = n49777 | n49778;
  assign n61126 = n49782 | n49783;
  assign n61127 = n49786 | n49787;
  assign n61128 = n49804 | n49805;
  assign n61129 = n49827 | n49828;
  assign n61130 = n49830 | n49831;
  assign n61131 = n49843 | n49844;
  assign n61132 = n49850 | n49851;
  assign n61133 = n49862 | n49863;
  assign n61134 = n49864 | n49865;
  assign n61135 = n49880 | n49877 | n49879;
  assign n61136 = n49895 | n49896;
  assign n61137 = n49910 | n49911;
  assign n61138 = n49924 | n49925;
  assign n61139 = n49926 | n49927;
  assign n61140 = n49966 | n49967;
  assign n61141 = n50010 | n50011;
  assign n61142 = n50064 | n50065;
  assign n61143 = n50068 | n50069;
  assign n61144 = n50077 | n50078;
  assign n61145 = n50107 | n50108;
  assign n61146 = n50186 | n50187;
  assign n61147 = n50249 | n50250;
  assign n61148 = n50251 | ~n50252;
  assign n61149 = n50257 | ~n50258;
  assign n61150 = n50273 | ~n50274;
  assign n61151 = n50289 | n50290;
  assign n61152 = n50305 | n50306;
  assign n61153 = n50311 | n50312;
  assign n61154 = n50331 | n50328 | n50330;
  assign n61155 = n50356 | n50357;
  assign n61156 = n50364 | n50365;
  assign n61157 = n50368 | n50369;
  assign n61158 = n50376 | n50377;
  assign n61159 = n50456 | n50457;
  assign n61160 = n50465 | n50466;
  assign n61161 = n50516 | n50517;
  assign n61162 = n50521 | n50522;
  assign n61163 = n50540 | n50541;
  assign n61164 = n50551 | n50552;
  assign n61165 = n50563 | n50564;
  assign n61166 = n50579 | n50580;
  assign n61167 = n50607 | ~n50608;
  assign n61168 = n50654 | n50655;
  assign n61169 = n50689 | n50690;
  assign n61170 = n50756 | n50757;
  assign n61171 = n50777 | n50778;
  assign n61172 = n50814 | n50815;
  assign n61173 = n50829 | n50830;
  assign n61174 = n50863 | n50864;
  assign n61175 = n50886 | n50887;
  assign n61176 = n50892 | n50893;
  assign n61177 = n50906 | n50907;
  assign n61178 = n50911 | n50912;
  assign n61179 = n50917 | n50918;
  assign n61180 = n50924 | n50925;
  assign n61181 = n50930 | n50931;
  assign n61182 = n50980 | n50981;
  assign n61183 = n50991 | n50992;
  assign n61184 = n50995 | n50996;
  assign n61185 = n51112 | n51113;
  assign n61186 = n51136 | n51137;
  assign n61187 = n51142 | n51143;
  assign n61188 = n51187 | n51188;
  assign n61189 = n51199 | n51200;
  assign n61190 = n51204 | n51205;
  assign n61191 = n51209 | n51207 | ~n51208;
  assign n61192 = n51210 | n51211;
  assign n61193 = n51247 | n51248;
  assign n61194 = n51249 | n51250;
  assign n61195 = n51263 | n51264;
  assign n61196 = n51271 | n51269 | n51270;
  assign n61197 = n51273 | n51275 | n51276 | n51277;
  assign n61198 = n51278 | n51279;
  assign n61199 = n51297 | n51294 | n51296;
  assign n61200 = n51366 | ~n51367;
  assign n61201 = n51394 | n51395;
  assign n61202 = n51456 | n51457;
  assign n61203 = n51471 | n51472;
  assign n61204 = n51537 | n51538;
  assign n61205 = n51545 | n51546;
  assign n61206 = n51547 | n51548;
  assign n61207 = n51564 | ~n51565;
  assign n61208 = n51581 | n51582;
  assign n61209 = n51592 | n51593;
  assign n61210 = n51624 | n51625;
  assign n61211 = n51651 | n51652;
  assign n61212 = n51692 | n51693;
  assign n61213 = n51702 | n51703;
  assign n61214 = n51709 | n51710;
  assign n61215 = n51713 | n51714;
  assign n61216 = n51718 | n51719;
  assign n61217 = n51740 | n51741;
  assign n61218 = n51747 | n51748;
  assign n61219 = n51756 | n51757;
  assign n61220 = n51768 | n51769;
  assign n61221 = n51774 | ~n51775;
  assign n61222 = n51828 | n51829;
  assign n61223 = n51839 | n51840;
  assign n61224 = n51842 | n51843;
  assign n61225 = n51875 | n51876;
  assign n61226 = n51909 | n51910;
  assign n61227 = n51939 | n51940;
  assign n61228 = n51956 | ~n51957;
  assign po397 = n51962 | ~n51963;
  assign n61230 = n52039 | n52040;
  assign n61231 = n52045 | n52046;
  assign n61232 = n52068 | n52069;
  assign n61233 = n52083 | n52084;
  assign n61234 = n52107 | n52108;
  assign n61235 = n52117 | ~n52118;
  assign n61236 = n52119 | n52120;
  assign n61237 = n52143 | n52144;
  assign n61238 = n52163 | n52164;
  assign n61239 = n52174 | n52175;
  assign n61240 = n52185 | n52186;
  assign n61241 = n52187 | n52188;
  assign n61242 = n52194 | n52192 | n52193;
  assign n61243 = n52208 | n52209;
  assign n61244 = n52217 | n52218;
  assign n61245 = n52224 | n52225;
  assign n61246 = n52243 | n52244;
  assign n61247 = n52255 | n52256;
  assign n61248 = n52271 | n52272;
  assign n61249 = n52285 | ~n52286;
  assign n61250 = n52300 | n52301;
  assign n61251 = n52311 | n52312;
  assign n61252 = n52321 | ~n52322;
  assign po398 = n52327 | ~n52328;
  assign n61254 = n52352 | n52353;
  assign n61255 = n52363 | n52364;
  assign n61256 = n52373 | n52374;
  assign n61257 = n52376 | ~n52377;
  assign n61258 = n52404 | n52405;
  assign n61259 = n52417 | ~n52418;
  assign n61260 = n52425 | n52426;
  assign n61261 = n52431 | n52432;
  assign n61262 = n52450 | n52451;
  assign n61263 = n52476 | n52477;
  assign n61264 = n52485 | n52486;
  assign n61265 = n52499 | n52500;
  assign n61266 = n52534 | n52535;
  assign n61267 = n52554 | n52555;
  assign n61268 = n52560 | ~n52561;
  assign n61269 = n52585 | n52582 | n52584;
  assign n61270 = n52586 | n52587;
  assign n61271 = n52630 | n52620 | ~n52629;
  assign n61272 = n52661 | n52662;
  assign n61273 = n52663 | n52664;
  assign n61274 = n52695 | n52696;
  assign n61275 = n52709 | n52710;
  assign n61276 = n52724 | n52725;
  assign n61277 = n52760 | n52761;
  assign n61278 = n52778 | ~n52779;
  assign po402 = n52784 | ~n52785;
  assign n61280 = n52813 | n52814;
  assign n61281 = n52828 | n52829;
  assign n61282 = n52865 | n52866;
  assign n61283 = n52904 | n52905;
  assign n61284 = n52919 | n52920;
  assign n61285 = n52927 | n52928;
  assign n61286 = n52931 | n52932;
  assign n61287 = n52943 | ~n52944;
  assign n61288 = n53002 | n53003;
  assign n61289 = n53008 | n53009;
  assign n61290 = n53021 | n53022;
  assign n61291 = n53025 | n53026;
  assign n61292 = n53035 | n53036;
  assign n61293 = n53050 | n53051;
  assign n61294 = n53055 | n53056;
  assign n61295 = n53059 | n53060;
  assign n61296 = n53084 | n53085;
  assign n61297 = n53104 | n53105;
  assign n61298 = n53111 | n53112;
  assign n61299 = n53133 | n53134;
  assign n61300 = n53142 | ~n53143;
  assign po403 = n53148 | ~n53149;
  assign n61302 = n53191 | n53192;
  assign n61303 = n53200 | n53201;
  assign n61304 = n53229 | n53230;
  assign n61305 = n53253 | n53254;
  assign n61306 = n53256 | n53257;
  assign n61307 = n53288 | ~n53289;
  assign n61308 = n53295 | n53296;
  assign n61309 = n53318 | n53319;
  assign n61310 = n53333 | n53334;
  assign n61311 = n53395 | n53396;
  assign n61312 = n53411 | ~n53412;
  assign po404 = n53417 | ~n53418;
  assign n61314 = n53429 | n53430;
  assign n61315 = n53435 | n53436;
  assign n61316 = n53455 | n53456;
  assign n61317 = n53459 | n53460;
  assign n61318 = n53463 | n53464;
  assign n61319 = n53481 | n53482;
  assign n61320 = n53496 | n53497;
  assign n61321 = n53510 | ~n53511;
  assign n61322 = n53520 | n53521;
  assign n61323 = n53531 | ~n53532;
  assign n61324 = n53542 | n53543;
  assign n61325 = n53611 | n53612;
  assign n61326 = n53625 | n53626;
  assign n61327 = n53630 | ~n53631;
  assign po405 = n53636 | ~n53637;
  assign n61329 = n53651 | n53652;
  assign n61330 = n53660 | ~n53661;
  assign n61331 = n53683 | n53684;
  assign n61332 = n53711 | n53708 | n53710;
  assign n61333 = n53714 | n53715;
  assign n61334 = n53731 | n53732;
  assign n61335 = n53799 | n53800;
  assign n61336 = n53834 | ~n53835;
  assign n61337 = n53846 | n53847;
  assign n61338 = n53851 | ~n53852;
  assign po406 = n53857 | ~n53858;
  assign n61340 = n53934 | n53935;
  assign n61341 = n53948 | n53949;
  assign n61342 = n53975 | n53976;
  assign n61343 = n53984 | n53985;
  assign n61344 = n53994 | n53995;
  assign n61345 = n54000 | n54001;
  assign n61346 = n54012 | n54013;
  assign n61347 = n54032 | n54033;
  assign n61348 = n54039 | n54040;
  assign n61349 = n54047 | n54048;
  assign n61350 = n54053 | n54054;
  assign n61351 = n54065 | n54066;
  assign n61352 = n54082 | n54083;
  assign n61353 = n54097 | n54098;
  assign n61354 = n54108 | n54109;
  assign n61355 = n54116 | n54117;
  assign n61356 = n54145 | n54146;
  assign n61357 = n54173 | n54174;
  assign n61358 = n54188 | n54189;
  assign n61359 = n54199 | n54200;
  assign n61360 = n54211 | n54212;
  assign n61361 = n54222 | n54223;
  assign n61362 = n54231 | n54232;
  assign n61363 = n54241 | n54242;
  assign n61364 = n54246 | n54247;
  assign n61365 = n54254 | n54255;
  assign n61366 = n54259 | n54260;
  assign n61367 = n54263 | ~n54264;
  assign n61368 = n54268 | n54269;
  assign n61369 = n54275 | n54276;
  assign n61370 = n54283 | n54284;
  assign n61371 = n54289 | n54290;
  assign n61372 = n54299 | n54300;
  assign n61373 = n54339 | n54340;
  assign n61374 = n54341 | n54342;
  assign n61375 = n54351 | n54352;
  assign n61376 = n54358 | n54359;
  assign n61377 = n54366 | n54367;
  assign n61378 = n54372 | n54373;
  assign n61379 = n54383 | n54384;
  assign n61380 = n54399 | n54400;
  assign n61381 = n54405 | n54406;
  assign n61382 = n54412 | n54413;
  assign n61383 = n54420 | n54421;
  assign n61384 = n54438 | ~n54439;
  assign n61385 = n54488 | n54489;
  assign n61386 = n54497 | n54498;
  assign n61387 = n54552 | n54553;
  assign n61388 = n54560 | n54561;
  assign n61389 = n54585 | n54586;
  assign n61390 = n54587 | ~n54588;
  assign n61391 = n54606 | n54607;
  assign po437 = n54608 | ~n54609;
  assign n61393 = n54622 | n54623;
  assign n61394 = n54634 | n54635;
  assign n61395 = n54665 | n54666;
  assign n61396 = n54678 | n54679;
  assign n61397 = n54698 | n54699;
  assign n61398 = n54708 | n54709;
  assign n61399 = n54819 | n54820;
  assign n61400 = n54879 | n54880;
  assign n61401 = n54965 | n54966;
  assign n61402 = n54997 | n54998;
  assign n61403 = n55023 | n55024;
  assign po468 = n55031 | n55032;
  assign po215 = n55045 | n55046;
  assign po217 = n55053 | n55054;
  assign n61407 = n55058 | n55059;
  assign po221 = n55063 | n55064;
  assign n61409 = n55068 | n55069;
  assign n61410 = n55151 | n55152;
  assign n61411 = n55197 | n55198;
  assign n61412 = n55217 | n55218;
  assign n61413 = n55253 | ~n55254;
  assign n61414 = n55263 | n55264;
  assign n61415 = n55294 | n55295;
  assign n61416 = n55336 | ~n55337;
  assign n61417 = n55376 | n55377;
  assign po622 = n55424 | ~n55425;
  assign n61419 = n55431 | ~n55432;
  assign n61420 = n55446 | n55447;
  assign po626 = n55478 | ~n55479;
  assign po627 = n55509 | ~n55510;
  assign po628 = n55540 | ~n55541;
  assign po629 = n55571 | ~n55572;
  assign n61425 = n55583 | n55584;
  assign n61426 = n55596 | n55597;
  assign n61427 = n55609 | n55610;
  assign n61428 = n55625 | ~n55626;
  assign n61429 = n55639 | n55640;
  assign n61430 = n55645 | n55646;
  assign n61431 = n55689 | ~n55690;
  assign n61432 = n55695 | ~n55696;
  assign n61433 = n55703 | n55704;
  assign n61434 = n55721 | n55722;
  assign n61435 = n55749 | n55750;
  assign n61436 = n55903 | ~n55904;
  assign n61437 = n55919 | ~n55920;
  assign n61438 = n55922 | n55923;
  assign n61439 = n55929 | n55930;
  assign n61440 = n55967 | ~n55968;
  assign n61441 = n55979 | ~n55980;
  assign n61442 = n55984 | ~n55985;
  assign n61443 = n55987 | n55988;
  assign n61444 = n55991 | n55992;
  assign n61445 = n56037 | n56038;
  assign n61446 = n56160 | ~n56161;
  assign n61447 = n56166 | ~n56167;
  assign n61448 = n56170 | n56171;
  assign n61449 = n56174 | n56175;
  assign n61450 = n56213 | ~n56214;
  assign n61451 = n56219 | ~n56220;
  assign n61452 = n56223 | n56224;
  assign n61453 = n56227 | n56228;
  assign n61454 = n56266 | n56267;
  assign n61455 = n56396 | ~n56397;
  assign n61456 = n56430 | ~n56431;
  assign n61457 = n56434 | ~n56435;
  assign n61458 = n56439 | n56440;
  assign n61459 = n56443 | n56444;
  assign n61460 = n56454 | n56455;
  assign n61461 = n56487 | ~n56488;
  assign n61462 = n56535 | n56536;
  assign n61463 = n56538 | n56539;
  assign n61464 = n56554 | n56555;
  assign n61465 = n56583 | n56584;
  assign n61466 = n56691 | n56692;
  assign n61467 = n56735 | n56736;
  assign n61468 = n56776 | n56777;
  assign po782 = n56843 | n56844;
  assign po784 = n56849 | n56850;
  assign po785 = n56855 | n56856;
  assign po897 = n56863 | n56864;
  assign po786 = n56869 | n56870;
  assign po787 = n56875 | n56876;
  assign po788 = n56881 | n56882;
  assign po789 = n56887 | n56888;
  assign po790 = n56893 | n56894;
  assign po791 = n56899 | n56900;
  assign po792 = n56905 | n56906;
  assign po793 = n56911 | n56912;
  assign po794 = n56917 | n56918;
  assign po795 = n56923 | n56924;
  assign po796 = n56929 | n56930;
  assign po797 = n56935 | n56936;
  assign po798 = n56941 | n56942;
  assign po800 = n56947 | n56948;
  assign po801 = n56953 | n56954;
  assign po802 = n56959 | n56960;
  assign po803 = n56965 | n56966;
  assign po804 = n56971 | n56972;
  assign po805 = n56977 | n56978;
  assign po806 = n56983 | n56984;
  assign po807 = n56989 | n56990;
  assign po808 = n56995 | n56996;
  assign po809 = n57001 | n57002;
  assign po810 = n57007 | n57008;
  assign po811 = n57013 | n57014;
  assign po812 = n57019 | n57020;
  assign po813 = n57025 | n57026;
  assign po814 = n57031 | n57032;
  assign po815 = n57037 | n57038;
  assign po817 = n57043 | n57044;
  assign po818 = n57049 | n57050;
  assign po819 = n57055 | n57056;
  assign po822 = n57061 | n57062;
  assign po826 = n57067 | n57068;
  assign po837 = n57073 | n57074;
  assign po838 = n57079 | n57080;
  assign po841 = n57086 | n57087;
  assign po843 = n57092 | n57093;
  assign po844 = n57098 | n57099;
  assign po845 = n57104 | n57105;
  assign po847 = n57110 | n57111;
  assign po848 = n57116 | n57117;
  assign po850 = n57122 | n57123;
  assign po851 = n57128 | n57129;
  assign po852 = n57134 | n57135;
  assign po853 = n57140 | n57141;
  assign po854 = n57146 | n57147;
  assign po855 = n57152 | n57153;
  assign po856 = n57158 | n57159;
  assign po857 = n57164 | n57165;
  assign po858 = n57170 | n57171;
  assign po859 = n57176 | n57177;
  assign po860 = n57182 | n57183;
  assign po861 = n57188 | n57189;
  assign po862 = n57194 | n57195;
  assign po863 = n57200 | n57201;
  assign po866 = n57206 | n57207;
  assign po867 = n57212 | n57213;
  assign po872 = n57218 | n57219;
  assign po880 = n57224 | n57225;
  assign po881 = n57230 | n57231;
  assign po882 = n57236 | n57237;
  assign po883 = n57242 | n57243;
  assign po884 = n57248 | n57249;
  assign po885 = n57254 | n57255;
  assign po886 = n57260 | n57261;
  assign po887 = n57266 | n57267;
  assign po889 = n57272 | n57273;
  assign po891 = n57278 | n57279;
  assign po892 = n57284 | n57285;
  assign po893 = n57290 | n57291;
  assign po894 = n57296 | n57297;
  assign po895 = n57302 | n57303;
  assign po988 = n57307 | n57308;
  assign n61547 = n57313 | n57314;
  assign n61548 = n57319 | n57320;
  assign n61549 = n57325 | n57326;
  assign n61550 = n57331 | n57332;
  assign n61551 = n57337 | n57338;
  assign n61552 = n57343 | n57344;
  assign n61553 = n57349 | n57350;
  assign n61554 = n57355 | n57356;
  assign n61555 = n57361 | n57362;
  assign n61556 = n57367 | n57368;
  assign n61557 = n57373 | n57374;
  assign n61558 = n57379 | n57380;
  assign n61559 = n57393 | ~n57394;
  assign n61560 = n57399 | ~n57400;
  assign n61561 = n57405 | ~n57406;
  assign n61562 = n57424 | n57417 | n57423;
  assign n61563 = n57442 | ~n57443;
  assign n61564 = n57448 | ~n57449;
  assign n61565 = n57454 | ~n57455;
  assign n61566 = n57473 | n57466 | n57472;
  assign n61567 = n57491 | ~n57492;
  assign n61568 = n57497 | ~n57498;
  assign n61569 = n57503 | ~n57504;
  assign n61570 = n57522 | n57515 | n57521;
  assign n61571 = n57540 | ~n57541;
  assign n61572 = n57546 | ~n57547;
  assign n61573 = n57552 | ~n57553;
  assign n61574 = n57571 | n57564 | n57570;
  assign n61575 = n57579 | n57580;
  assign n61576 = n57584 | n57585;
  assign n61577 = n57594 | ~n57595;
  assign po763 = n57600 | ~n57601;
  assign n61579 = n57606 | n57607;
  assign n61580 = n57613 | n57614;
  assign n61581 = n57620 | ~n57621;
  assign po774 = n57626 | ~n57627;
  assign po764 = n57641 | n57642;
  assign po765 = n57647 | n57648;
  assign po766 = n57653 | n57654;
  assign po767 = n57659 | n57660;
  assign po768 = n57665 | n57666;
  assign po769 = n57671 | n57672;
  assign po770 = n57677 | n57678;
  assign po775 = n57683 | n57684;
  assign po776 = n57689 | n57690;
  assign po777 = n57695 | n57696;
  assign po778 = n57701 | n57702;
  assign po779 = n57707 | n57708;
  assign po780 = n57713 | n57714;
  assign po783 = n57725 | n57726;
  assign po799 = n57731 | n57732;
  assign n61598 = n57737 | n57738;
  assign n61599 = n57743 | n57744;
  assign n61600 = n57749 | n57750;
  assign n61601 = n57755 | n57756;
  assign n61602 = n57761 | n57762;
  assign n61603 = n57767 | n57768;
  assign n61604 = n57775 | n57776;
  assign n61605 = n57781 | n57782;
  assign n61606 = n57787 | n57788;
  assign n61607 = n57793 | n57794;
  assign n61608 = n57799 | n57800;
  assign n61609 = n57805 | n57806;
  assign n61610 = n57811 | n57812;
  assign n61611 = n57817 | n57818;
  assign n61612 = n57823 | n57824;
  assign n61613 = n57829 | n57830;
  assign n61614 = n57835 | n57836;
  assign n61615 = n57841 | n57842;
  assign n61616 = n57847 | n57848;
  assign n61617 = n57853 | n57854;
  assign n61618 = n57863 | n57864;
  assign n61619 = n57870 | n57871;
  assign po1079 = n57880 | ~n57881;
  assign po1081 = n57886 | ~n57887;
  assign po1082 = n57892 | ~n57893;
  assign po1087 = n57898 | ~n57899;
  assign po1090 = n57904 | ~n57905;
  assign po1092 = n57910 | ~n57911;
  assign po1093 = n57916 | ~n57917;
  assign po1097 = n57922 | ~n57923;
  assign po1098 = n57928 | ~n57929;
  assign po1099 = n57934 | ~n57935;
  assign n61630 = n57956 | ~n57957;
  assign n61631 = n57962 | ~n57963;
  assign n61632 = n57968 | ~n57969;
  assign n61633 = n57974 | ~n57975;
  assign n61634 = n57980 | ~n57981;
  assign n61635 = n57986 | ~n57987;
  assign n61636 = n57992 | ~n57993;
  assign n61637 = n57998 | ~n57999;
  assign n61638 = n58015 | n58016;
  assign n61639 = n58022 | n58023;
  assign po745 = n58036 | n58037;
  assign n61641 = n58042 | n58043;
  assign po748 = n58048 | n58049;
  assign po749 = n58054 | n58055;
  assign po758 = n58090 | n58091;
  assign n61645 = n58102 | ~n58103;
  assign n61646 = n58117 | n58118;
  assign n61647 = n58123 | ~n58124;
  assign n61648 = n58147 | ~n58148;
  assign n61649 = n58154 | n58155;
  assign n61650 = n58172 | n58173;
  assign n61651 = n58176 | n58177;
  assign n61652 = n58192 | n58193;
  assign po888 = n58204 | n58205;
  assign n61654 = n58220 | n58221;
  assign n61655 = n58245 | n58246;
  assign n61656 = n58267 | n58268;
  assign n61657 = n58283 | n58284;
  assign n61658 = n58298 | n58299;
  assign n61659 = n58307 | n58308;
  assign n61660 = n58408 | ~n58409;
  assign n61661 = n58414 | ~n58415;
  assign n61662 = n58420 | ~n58421;
  assign n61663 = n58426 | ~n58427;
  assign n61664 = n58432 | ~n58433;
  assign n61665 = n58438 | ~n58439;
  assign n61666 = n58444 | ~n58445;
  assign n61667 = n58450 | ~n58451;
  assign n61668 = n58456 | ~n58457;
  assign n61669 = n58462 | ~n58463;
  assign n61670 = n58468 | ~n58469;
  assign n61671 = n58474 | ~n58475;
  assign n61672 = n58480 | ~n58481;
  assign n61673 = n58486 | ~n58487;
  assign n61674 = n58492 | ~n58493;
  assign n61675 = n58498 | ~n58499;
  assign n61676 = n58504 | ~n58505;
  assign n61677 = n58510 | ~n58511;
  assign n61678 = n58516 | ~n58517;
  assign n61679 = n58522 | ~n58523;
  assign n61680 = n58528 | ~n58529;
  assign n61681 = n58534 | ~n58535;
  assign n61682 = n58540 | ~n58541;
  assign n61683 = n58546 | ~n58547;
  assign n61684 = n58552 | ~n58553;
  assign n61685 = n58558 | ~n58559;
  assign n61686 = n58564 | ~n58565;
  assign n61687 = n58570 | ~n58571;
  assign n61688 = n58576 | ~n58577;
  assign n61689 = n58582 | ~n58583;
  assign n61690 = n58588 | ~n58589;
  assign n61691 = n58594 | ~n58595;
  assign n61692 = n58694 | n58695;
  assign n61693 = n58707 | n58708;
  assign n61694 = n58717 | n58718;
  assign n61695 = n58727 | n58728;
  assign n61696 = n58737 | n58738;
  assign n61697 = n58747 | n58748;
  assign po1078 = n58767 | ~n58768;
  assign po0 = pi668;
  assign po1 = pi672;
  assign po2 = pi664;
  assign po3 = pi667;
  assign po4 = pi676;
  assign po5 = pi673;
  assign po6 = pi675;
  assign po7 = pi666;
  assign po8 = pi679;
  assign po9 = pi674;
  assign po10 = pi663;
  assign po11 = pi670;
  assign po12 = pi677;
  assign po13 = pi682;
  assign po14 = pi671;
  assign po15 = pi678;
  assign po16 = pi718;
  assign po17 = pi707;
  assign po18 = pi708;
  assign po19 = pi713;
  assign po20 = pi711;
  assign po21 = pi716;
  assign po22 = pi733;
  assign po23 = pi712;
  assign po24 = pi689;
  assign po25 = pi717;
  assign po26 = pi692;
  assign po27 = pi719;
  assign po28 = pi722;
  assign po29 = pi714;
  assign po30 = pi720;
  assign po31 = pi685;
  assign po32 = pi837;
  assign po33 = pi850;
  assign po34 = pi872;
  assign po35 = pi871;
  assign po36 = pi881;
  assign po37 = pi866;
  assign po38 = pi876;
  assign po39 = pi873;
  assign po40 = pi874;
  assign po41 = pi859;
  assign po42 = pi855;
  assign po43 = pi852;
  assign po44 = pi870;
  assign po45 = pi848;
  assign po46 = pi865;
  assign po47 = pi856;
  assign po48 = pi853;
  assign po49 = pi847;
  assign po50 = pi857;
  assign po51 = pi854;
  assign po52 = pi858;
  assign po53 = pi845;
  assign po54 = pi838;
  assign po55 = pi842;
  assign po56 = pi843;
  assign po57 = pi839;
  assign po58 = pi844;
  assign po59 = pi868;
  assign po60 = pi851;
  assign po61 = pi867;
  assign po62 = pi880;
  assign po63 = pi860;
  assign po64 = pi1030;
  assign po65 = pi1034;
  assign po66 = pi1015;
  assign po67 = pi1020;
  assign po68 = pi1025;
  assign po69 = pi1005;
  assign po70 = pi996;
  assign po71 = pi1012;
  assign po72 = pi993;
  assign po73 = pi1016;
  assign po74 = pi1021;
  assign po75 = pi1010;
  assign po76 = pi1027;
  assign po77 = pi1018;
  assign po78 = pi1017;
  assign po79 = pi1024;
  assign po80 = pi1009;
  assign po81 = pi1032;
  assign po82 = pi1003;
  assign po83 = pi997;
  assign po84 = pi1013;
  assign po85 = pi1011;
  assign po86 = pi1008;
  assign po87 = pi1019;
  assign po88 = pi1031;
  assign po89 = pi1022;
  assign po90 = pi1000;
  assign po91 = pi1023;
  assign po92 = pi1002;
  assign po93 = pi1026;
  assign po94 = pi1006;
  assign po95 = pi998;
  assign po96 = pi31;
  assign po97 = pi80;
  assign po98 = pi893;
  assign po99 = pi467;
  assign po100 = pi78;
  assign po101 = pi112;
  assign po102 = pi13;
  assign po103 = pi25;
  assign po104 = pi226;
  assign po105 = pi127;
  assign po106 = pi822;
  assign po107 = pi808;
  assign po108 = pi227;
  assign po109 = pi477;
  assign po110 = pi834;
  assign po111 = pi229;
  assign po112 = pi12;
  assign po113 = pi11;
  assign po114 = pi10;
  assign po115 = pi9;
  assign po116 = pi8;
  assign po117 = pi7;
  assign po118 = pi6;
  assign po119 = pi5;
  assign po120 = pi4;
  assign po121 = pi3;
  assign po122 = pi0;
  assign po123 = pi2;
  assign po124 = pi1;
  assign po125 = pi310;
  assign po126 = pi302;
  assign po127 = pi475;
  assign po128 = pi474;
  assign po129 = pi466;
  assign po130 = pi473;
  assign po131 = pi471;
  assign po132 = pi472;
  assign po133 = pi470;
  assign po134 = pi469;
  assign po135 = pi465;
  assign po136 = pi1028;
  assign po137 = pi1033;
  assign po138 = pi995;
  assign po139 = pi994;
  assign po140 = pi28;
  assign po141 = pi27;
  assign po142 = pi26;
  assign po143 = pi29;
  assign po144 = pi15;
  assign po145 = pi14;
  assign po146 = pi21;
  assign po147 = pi20;
  assign po148 = pi19;
  assign po149 = pi18;
  assign po150 = pi17;
  assign po151 = pi16;
  assign po152 = pi1096;
  assign po153 = ~n38867;
  assign po154 = ~n43162;
  assign po157 = ~n41590;
  assign po160 = ~n42344;
  assign po163 = ~n43856;
  assign po164 = ~n44108;
  assign po168 = pi228;
  assign po169 = pi22;
  assign po170 = ~pi1090;
  assign po179 = pi1089;
  assign po180 = pi23;
  assign po181 = po167;
  assign po183 = ~n45025;
  assign po184 = ~n57942;
  assign po185 = ~n57944;
  assign po186 = ~n57946;
  assign po187 = ~n57948;
  assign po188 = pi37;
  assign po189 = ~n5145;
  assign po200 = ~n36677;
  assign po201 = ~n36878;
  assign po202 = ~n37623;
  assign po237 = ~n30545;
  assign po257 = ~n37701;
  assign po259 = ~n37796;
  assign po263 = pi117;
  assign po270 = ~n57951;
  assign po276 = ~n30924;
  assign po277 = ~n32942;
  assign po278 = ~n29026;
  assign po279 = ~n39408;
  assign po280 = ~n31396;
  assign po282 = ~n39902;
  assign po283 = ~n60675;
  assign po285 = pi131;
  assign po289 = ~n40562;
  assign po290 = ~n40978;
  assign po291 = ~n41103;
  assign po292 = ~n41226;
  assign po293 = ~n41319;
  assign po294 = ~n44979;
  assign po303 = ~n33061;
  assign po305 = ~n33304;
  assign po309 = ~n33659;
  assign po310 = ~n33761;
  assign po318 = ~n34303;
  assign po323 = ~n34662;
  assign po325 = ~n34809;
  assign po326 = ~n34911;
  assign po327 = ~n34992;
  assign po328 = ~n35094;
  assign po329 = ~n35196;
  assign po352 = ~n32774;
  assign po353 = ~n32858;
  assign po355 = ~n26168;
  assign po356 = ~n59869;
  assign po364 = ~n59918;
  assign po365 = ~n59924;
  assign po366 = ~n25420;
  assign po368 = ~n35318;
  assign po369 = ~n35343;
  assign po370 = ~n35378;
  assign po371 = ~n35403;
  assign po372 = ~n35798;
  assign po374 = ~n25439;
  assign po376 = ~n35438;
  assign po384 = ~n37122;
  assign po385 = ~n36319;
  assign po386 = pi232;
  assign po388 = pi236;
  assign po390 = ~n49796;
  assign po391 = ~n50787;
  assign po394 = ~n50121;
  assign po395 = ~n51373;
  assign po408 = ~n49011;
  assign po417 = ~n49044;
  assign po418 = ~n49047;
  assign po419 = ~n55299;
  assign po421 = ~n54034;
  assign po422 = ~n54084;
  assign po427 = ~n54270;
  assign po430 = ~n53936;
  assign po432 = ~n61149;
  assign po433 = ~n54353;
  assign po434 = ~n54407;
  assign po441 = ~n55303;
  assign po455 = ~n61630;
  assign po457 = ~n55056;
  assign po458 = ~n55035;
  assign po460 = ~n61631;
  assign po461 = ~n61632;
  assign po462 = ~n61633;
  assign po463 = ~n61634;
  assign po464 = ~n61635;
  assign po465 = ~n61636;
  assign po466 = ~n61637;
  assign po467 = ~n55387;
  assign po472 = ~n45205;
  assign po473 = ~n45208;
  assign po474 = ~n45211;
  assign po475 = ~n45214;
  assign po476 = ~n45217;
  assign po477 = ~n45220;
  assign po478 = ~n45223;
  assign po479 = ~n45226;
  assign po480 = ~n45229;
  assign po481 = ~n45232;
  assign po482 = ~n45235;
  assign po483 = ~n45238;
  assign po484 = ~n45241;
  assign po485 = ~n45244;
  assign po486 = ~n45247;
  assign po487 = ~n60839;
  assign po488 = ~n60842;
  assign po490 = ~n45250;
  assign po491 = ~n45253;
  assign po492 = ~n45256;
  assign po493 = ~n54703;
  assign po494 = ~n54706;
  assign po495 = ~n45259;
  assign po496 = ~n45262;
  assign po499 = ~n54712;
  assign po500 = ~n54715;
  assign po501 = ~n45265;
  assign po502 = ~n54718;
  assign po503 = ~n54721;
  assign po504 = ~n54724;
  assign po505 = ~n54727;
  assign po506 = ~n45268;
  assign po507 = ~n54730;
  assign po508 = ~n54733;
  assign po509 = ~n45271;
  assign po510 = ~n45274;
  assign po511 = ~n54736;
  assign po512 = ~n54739;
  assign po513 = ~n54742;
  assign po514 = ~n54745;
  assign po515 = ~n54748;
  assign po516 = ~n54751;
  assign po517 = ~n54754;
  assign po518 = ~n54757;
  assign po519 = ~n54760;
  assign po520 = ~n54763;
  assign po521 = ~n54766;
  assign po522 = ~n45277;
  assign po523 = ~n45280;
  assign po524 = ~n54769;
  assign po525 = ~n54772;
  assign po526 = ~n45283;
  assign po527 = ~n54775;
  assign po528 = ~n45286;
  assign po529 = ~n45289;
  assign po530 = ~n54778;
  assign po531 = ~n54781;
  assign po532 = ~n45292;
  assign po533 = ~n54784;
  assign po534 = ~n45295;
  assign po535 = ~n45298;
  assign po536 = ~n54787;
  assign po537 = ~n54790;
  assign po538 = ~n54793;
  assign po539 = ~n54796;
  assign po540 = ~n54799;
  assign po541 = ~n54802;
  assign po542 = ~n54805;
  assign po543 = ~n54808;
  assign po544 = ~n54811;
  assign po545 = ~n54814;
  assign po546 = ~n54817;
  assign po547 = ~n54823;
  assign po548 = ~n54826;
  assign po549 = ~n54829;
  assign po550 = ~n54832;
  assign po551 = ~n45301;
  assign po552 = ~n54835;
  assign po553 = ~n45304;
  assign po554 = ~n45307;
  assign po555 = ~n54838;
  assign po556 = ~n45310;
  assign po557 = ~n54841;
  assign po558 = ~n54844;
  assign po559 = ~n45313;
  assign po560 = ~n54847;
  assign po561 = ~n54850;
  assign po562 = ~n54853;
  assign po563 = ~n54856;
  assign po564 = ~n54859;
  assign po565 = ~n54862;
  assign po566 = ~n54865;
  assign po567 = ~n54868;
  assign po568 = ~n54871;
  assign po569 = ~n54874;
  assign po570 = ~n54877;
  assign po571 = ~n54883;
  assign po572 = ~n54886;
  assign po573 = ~n45316;
  assign po574 = ~n54889;
  assign po575 = ~n54892;
  assign po576 = ~n45319;
  assign po577 = ~n54895;
  assign po578 = ~n45322;
  assign po579 = ~n45325;
  assign po580 = ~n54898;
  assign po581 = ~n45328;
  assign po582 = ~n54901;
  assign po583 = ~n54904;
  assign po584 = ~n45331;
  assign po585 = ~n54907;
  assign po586 = ~n54910;
  assign po587 = ~n54913;
  assign po588 = ~n54916;
  assign po589 = ~n54919;
  assign po590 = ~n54922;
  assign po591 = ~n54925;
  assign po592 = ~n54928;
  assign po593 = ~n54931;
  assign po594 = ~n54934;
  assign po595 = ~n54937;
  assign po596 = ~n45334;
  assign po597 = ~n45337;
  assign po598 = ~n54940;
  assign po599 = ~n45340;
  assign po600 = ~n54943;
  assign po601 = ~n45343;
  assign po602 = ~n54946;
  assign po603 = ~n45346;
  assign po604 = ~n45349;
  assign po605 = ~n45352;
  assign po606 = ~n45355;
  assign po607 = ~n54949;
  assign po608 = ~n45358;
  assign po609 = ~n54952;
  assign po610 = ~n45361;
  assign po611 = ~n45364;
  assign po612 = ~n54955;
  assign po613 = ~n54958;
  assign po615 = ~n45367;
  assign po616 = ~n45370;
  assign po617 = ~n45373;
  assign po618 = ~n45376;
  assign po619 = ~n45379;
  assign po620 = ~n54961;
  assign po621 = ~n45382;
  assign po625 = ~n45409;
  assign po633 = ~n45517;
  assign po634 = ~n45458;
  assign po636 = pi583;
  assign po638 = ~n55073;
  assign po639 = ~n55076;
  assign po640 = ~n55079;
  assign po641 = ~n55082;
  assign po642 = ~n55085;
  assign po643 = ~n55088;
  assign po644 = ~n55091;
  assign po646 = ~n55097;
  assign po647 = ~n55100;
  assign po648 = ~n55103;
  assign po649 = ~n55106;
  assign po650 = ~n55109;
  assign po652 = ~n55115;
  assign po653 = ~n55118;
  assign po655 = ~n55124;
  assign po656 = ~n55127;
  assign po657 = ~n55130;
  assign po658 = ~n55133;
  assign po659 = ~n55136;
  assign po660 = ~n55139;
  assign po661 = ~n55142;
  assign po662 = ~n61410;
  assign po663 = ~n55155;
  assign po664 = ~n55158;
  assign po665 = ~n55161;
  assign po666 = ~n55164;
  assign po667 = ~n55167;
  assign po668 = ~n55171;
  assign po669 = ~n55174;
  assign po670 = ~n55177;
  assign po671 = ~n55180;
  assign po672 = ~n55183;
  assign po673 = ~n55186;
  assign po674 = ~n55189;
  assign po675 = ~n61411;
  assign po677 = ~n55204;
  assign po678 = ~n55207;
  assign po679 = ~n55210;
  assign po680 = ~n61412;
  assign po682 = ~n55224;
  assign po683 = ~n55227;
  assign po684 = ~n55230;
  assign po685 = ~n55233;
  assign po686 = ~n55236;
  assign po687 = ~n55239;
  assign po688 = ~n55242;
  assign po689 = ~n55245;
  assign po690 = ~n55248;
  assign po692 = ~n56660;
  assign po693 = ~n56663;
  assign po694 = ~n56666;
  assign po695 = ~n56669;
  assign po696 = ~n56672;
  assign po697 = ~n56675;
  assign po698 = ~n56678;
  assign po699 = ~n56681;
  assign po700 = ~n56684;
  assign po701 = ~n61466;
  assign po702 = ~n56695;
  assign po703 = ~n56698;
  assign po704 = ~n56701;
  assign po705 = ~n56704;
  assign po706 = ~n56707;
  assign po708 = ~n56713;
  assign po709 = ~n56716;
  assign po710 = ~n56719;
  assign po711 = ~n56722;
  assign po712 = ~n56725;
  assign po713 = ~n56728;
  assign po714 = ~n61467;
  assign po715 = ~n56739;
  assign po716 = ~n56742;
  assign po717 = ~n56745;
  assign po718 = ~n56748;
  assign po719 = ~n56751;
  assign po720 = ~n56754;
  assign po721 = ~n56757;
  assign po722 = ~n56760;
  assign po723 = ~n56763;
  assign po724 = ~n46140;
  assign po725 = ~n56766;
  assign po727 = ~n61468;
  assign po728 = ~n56780;
  assign po729 = ~n56783;
  assign po730 = ~n56786;
  assign po731 = ~n56789;
  assign po732 = ~n56792;
  assign po733 = ~n56795;
  assign po734 = ~n56798;
  assign po735 = ~n56801;
  assign po736 = ~n56804;
  assign po737 = ~n56807;
  assign po738 = ~n56810;
  assign po739 = ~n56813;
  assign po741 = ~n56816;
  assign po742 = ~n56819;
  assign po743 = ~n56822;
  assign po744 = ~n47396;
  assign po747 = ~n61641;
  assign po755 = ~n56828;
  assign po759 = ~n47413;
  assign po760 = ~n57589;
  assign po761 = ~n57636;
  assign po771 = ~n57608;
  assign po772 = ~n56833;
  assign po773 = ~n57615;
  assign po781 = ~n57720;
  assign po820 = ~n48693;
  assign po821 = ~n48738;
  assign po823 = ~n48780;
  assign po824 = ~n48825;
  assign po825 = ~n47699;
  assign po827 = ~n48861;
  assign po828 = ~n48897;
  assign po829 = ~n47741;
  assign po830 = ~n47783;
  assign po831 = ~n47832;
  assign po832 = ~n47877;
  assign po833 = ~n47919;
  assign po834 = ~n48933;
  assign po835 = ~n48969;
  assign po836 = ~n47962;
  assign po839 = ~n49005;
  assign po840 = ~n35649;
  assign po842 = ~n48014;
  assign po846 = ~n48058;
  assign po849 = ~n48105;
  assign po864 = ~n61008;
  assign po868 = ~n61014;
  assign po869 = ~n48291;
  assign po870 = ~n61021;
  assign po871 = ~n48384;
  assign po874 = ~n48472;
  assign po876 = ~n48560;
  assign po877 = ~n48607;
  assign po878 = ~n58178;
  assign po879 = ~n48652;
  assign po896 = ~n61547;
  assign po898 = ~n61548;
  assign po899 = ~n61549;
  assign po900 = ~n61550;
  assign po901 = ~n61551;
  assign po902 = ~n61552;
  assign po903 = ~n61553;
  assign po905 = ~n61554;
  assign po906 = ~n61555;
  assign po907 = ~n61556;
  assign po908 = ~n61557;
  assign po909 = ~n61558;
  assign po910 = ~n61598;
  assign po911 = ~n61599;
  assign po912 = ~n61600;
  assign po913 = ~n61601;
  assign po914 = ~n61602;
  assign po915 = ~n61603;
  assign po916 = ~n61604;
  assign po917 = ~n61605;
  assign po918 = ~n61606;
  assign po919 = ~n61607;
  assign po920 = ~n61608;
  assign po921 = ~n61609;
  assign po923 = ~n61610;
  assign po924 = ~n61611;
  assign po925 = ~n61612;
  assign po926 = ~n58235;
  assign po927 = ~n61613;
  assign po928 = ~n58259;
  assign po929 = ~n61614;
  assign po931 = ~n61615;
  assign po933 = ~n61616;
  assign po934 = ~n61617;
  assign po935 = ~n58317;
  assign po936 = ~n57855;
  assign po937 = ~n57856;
  assign po938 = ~n58320;
  assign po939 = ~n57630;
  assign po940 = ~n58323;
  assign po941 = ~n58326;
  assign po942 = ~n58329;
  assign po944 = ~n58332;
  assign po945 = ~n58335;
  assign po946 = ~n58338;
  assign po947 = ~n58341;
  assign po948 = ~n58344;
  assign po949 = ~n58347;
  assign po950 = ~n37420;
  assign po951 = ~n58351;
  assign po952 = ~n58354;
  assign po955 = ~n58357;
  assign po957 = ~n58363;
  assign po958 = ~n58366;
  assign po961 = ~n58372;
  assign po964 = ~n58375;
  assign po965 = ~n58378;
  assign po967 = ~n58384;
  assign po968 = ~n58387;
  assign po970 = ~n58393;
  assign po972 = ~n58399;
  assign po973 = ~n58402;
  assign po975 = ~n45901;
  assign po990 = ~n45916;
  assign po993 = ~n61660;
  assign po994 = ~n61661;
  assign po995 = ~n61662;
  assign po996 = ~n58752;
  assign po998 = ~n61663;
  assign po999 = ~n61664;
  assign po1000 = ~n61665;
  assign po1001 = ~n61666;
  assign po1002 = ~n58686;
  assign po1003 = ~n61667;
  assign po1004 = ~n61668;
  assign po1005 = ~n58755;
  assign po1006 = ~n61669;
  assign po1007 = ~n61670;
  assign po1008 = ~n61671;
  assign po1009 = ~n61672;
  assign po1010 = ~n61673;
  assign po1011 = ~n61674;
  assign po1012 = ~n61675;
  assign po1013 = ~n61676;
  assign po1014 = ~n61677;
  assign po1015 = ~n61678;
  assign po1016 = ~n61679;
  assign po1017 = ~n58696;
  assign po1018 = ~n58699;
  assign po1019 = ~n58758;
  assign po1020 = ~n58761;
  assign po1021 = ~n61680;
  assign po1022 = ~n61681;
  assign po1023 = ~n61682;
  assign po1024 = ~n61683;
  assign po1025 = ~n58709;
  assign po1026 = ~n61684;
  assign po1027 = ~n61685;
  assign po1028 = ~n61686;
  assign po1029 = ~n61687;
  assign po1030 = ~n61688;
  assign po1032 = ~n61689;
  assign po1033 = ~n58729;
  assign po1034 = ~n58739;
  assign po1035 = ~n58749;
  assign po1036 = ~n61690;
  assign po1037 = ~n61691;
  assign po1038 = ~n58992;
  assign po1039 = ~n58597;
  assign po1040 = ~n58600;
  assign po1041 = ~n58603;
  assign po1042 = ~n58606;
  assign po1043 = ~n58608;
  assign po1044 = ~n58611;
  assign po1045 = ~n58614;
  assign po1046 = ~n58617;
  assign po1047 = ~n58620;
  assign po1048 = ~n58623;
  assign po1049 = ~n28389;
  assign po1050 = ~n58626;
  assign po1051 = ~n58629;
  assign po1052 = ~n58632;
  assign po1053 = pi67;
  assign po1054 = ~n58635;
  assign po1055 = ~n58637;
  assign po1056 = ~n58640;
  assign po1057 = ~n2707;
  assign po1058 = ~n58643;
  assign po1059 = ~n58646;
  assign po1060 = ~n58648;
  assign po1061 = ~n58650;
  assign po1062 = ~n58653;
  assign po1064 = ~n58655;
  assign po1065 = ~n58658;
  assign po1066 = ~n58661;
  assign po1067 = ~n58664;
  assign po1068 = ~n58666;
  assign po1069 = ~n58669;
  assign po1071 = ~n58672;
  assign po1072 = ~n58674;
  assign po1073 = ~n58677;
  assign po1074 = ~n58680;
  assign po1075 = ~n58683;
  assign po1076 = ~n60885;
  assign po1077 = ~n45932;
  assign po1088 = ~n45956;
  assign po1089 = ~n45959;
  assign po1091 = ~n45962;
  assign po1094 = ~n45965;
  assign po1096 = ~n45974;
  assign po1100 = ~n60890;
  assign po1101 = ~n2782;
  assign po1103 = ~n57875;
  assign po1105 = ~n61416;
  assign po1108 = pi1134;
  assign po1109 = pi964;
  assign po1110 = ~pi954;
  assign po1111 = pi965;
  assign po1112 = ~n45982;
  assign po1113 = pi991;
  assign po1114 = pi985;
  assign po1117 = pi1014;
  assign po1119 = pi1029;
  assign po1120 = pi1004;
  assign po1121 = pi1007;
  assign po1123 = pi1135;
  assign po1130 = ~pi278;
  assign po1133 = ~n57936;
  assign po1134 = pi1064;
  assign po1136 = pi299;
  assign po1137 = ~n57937;
  assign po1138 = pi1075;
  assign po1139 = pi1052;
  assign po1140 = pi771;
  assign po1141 = pi765;
  assign po1142 = pi605;
  assign po1143 = pi601;
  assign po1144 = pi278;
  assign po1145 = pi279;
  assign po1146 = ~pi915;
  assign po1147 = ~pi825;
  assign po1148 = ~pi826;
  assign po1149 = ~pi913;
  assign po1150 = ~pi894;
  assign po1151 = ~pi905;
  assign po1152 = pi1095;
  assign po1153 = ~pi890;
  assign po1154 = pi1094;
  assign po1155 = ~pi906;
  assign po1156 = ~pi896;
  assign po1157 = ~pi909;
  assign po1158 = ~pi911;
  assign po1159 = ~pi908;
  assign po1160 = ~pi891;
  assign po1161 = ~pi902;
  assign po1162 = ~pi903;
  assign po1163 = ~pi883;
  assign po1164 = ~pi888;
  assign po1165 = ~pi919;
  assign po1166 = ~pi886;
  assign po1167 = ~pi912;
  assign po1168 = ~pi895;
  assign po1169 = ~pi916;
  assign po1170 = ~pi889;
  assign po1171 = ~pi900;
  assign po1172 = ~pi885;
  assign po1173 = ~pi904;
  assign po1174 = ~pi899;
  assign po1175 = ~pi918;
  assign po1176 = ~pi898;
  assign po1177 = ~pi917;
  assign po1178 = ~pi827;
  assign po1179 = ~pi887;
  assign po1180 = ~pi884;
  assign po1181 = ~pi910;
  assign po1182 = ~pi828;
  assign po1183 = ~pi892;
  assign po1184 = pi1187;
  assign po1185 = pi1172;
  assign po1186 = pi1170;
  assign po1187 = pi1138;
  assign po1188 = pi1177;
  assign po1189 = pi1178;
  assign po1190 = pi863;
  assign po1191 = pi1203;
  assign po1192 = pi1185;
  assign po1193 = pi1171;
  assign po1194 = pi1192;
  assign po1195 = pi1137;
  assign po1196 = pi1186;
  assign po1197 = pi1165;
  assign po1198 = pi1164;
  assign po1199 = pi1098;
  assign po1200 = pi1183;
  assign po1201 = pi230;
  assign po1202 = pi1169;
  assign po1203 = pi1136;
  assign po1204 = pi1181;
  assign po1205 = pi849;
  assign po1206 = pi1193;
  assign po1207 = pi1182;
  assign po1208 = pi1168;
  assign po1209 = pi1175;
  assign po1210 = pi1191;
  assign po1211 = pi1099;
  assign po1212 = pi1174;
  assign po1213 = pi1179;
  assign po1214 = pi1202;
  assign po1215 = pi1176;
  assign po1216 = pi1173;
  assign po1217 = pi1201;
  assign po1218 = pi1167;
  assign po1219 = pi840;
  assign po1220 = pi1189;
  assign po1221 = pi1195;
  assign po1222 = pi864;
  assign po1223 = pi1190;
  assign po1224 = pi1188;
  assign po1225 = pi1180;
  assign po1226 = pi1194;
  assign po1227 = pi1097;
  assign po1228 = pi1166;
  assign po1229 = pi1200;
  assign po1230 = pi1184;
endmodule
