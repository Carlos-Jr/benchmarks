module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10   );
  input  pi0 , pi1 , pi2 ,
    pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 ;
  output po0 , po1 , po2 ,
    po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 ;
  wire n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379,
    n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414,
    n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463,
    n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568,
    n569, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646,
    n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667,
    n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681,
    n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695,
    n696, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1108;
  assign n22 = ~pi5  & pi7 ;
  assign n23 = pi7  & pi8 ;
  assign n24 = ~pi5  & n23;
  assign n25 = pi8  & n22;
  assign n26 = ~pi0  & ~pi1 ;
  assign n27 = pi2  & ~pi9 ;
  assign n28 = n26 & n27;
  assign n29 = n998 & n28;
  assign n30 = ~pi7  & pi9 ;
  assign n31 = ~n998 & ~n30;
  assign n32 = pi1  & ~n31;
  assign n33 = pi1  & ~pi7 ;
  assign n34 = ~pi5  & ~pi9 ;
  assign n35 = ~n33 & n34;
  assign n36 = ~n32 & ~n35;
  assign n37 = pi0  & ~pi2 ;
  assign n38 = ~n36 & n37;
  assign n39 = ~n29 & ~n38;
  assign n40 = ~pi3  & ~n39;
  assign n41 = ~pi0  & pi9 ;
  assign n42 = pi1  & ~n41;
  assign n43 = ~pi3  & ~pi5 ;
  assign n44 = ~pi1  & pi9 ;
  assign n45 = n43 & ~n44;
  assign n46 = ~n42 & ~n44;
  assign n47 = n43 & n46;
  assign n48 = ~n42 & n45;
  assign n49 = pi0  & ~pi9 ;
  assign n50 = ~pi1  & ~n49;
  assign n51 = pi1  & ~pi9 ;
  assign n52 = ~pi7  & ~n51;
  assign n53 = ~n50 & n52;
  assign n54 = ~n999 & ~n53;
  assign n55 = ~pi2  & ~n54;
  assign n56 = ~pi0  & pi5 ;
  assign n57 = pi0  & ~pi1 ;
  assign n58 = pi2  & ~n57;
  assign n59 = pi1  & pi2 ;
  assign n60 = ~pi2  & ~pi5 ;
  assign n61 = ~pi0  & ~n60;
  assign n62 = ~n59 & ~n61;
  assign n63 = ~n56 & ~n58;
  assign n64 = ~pi9  & ~n1000;
  assign n65 = ~pi2  & ~pi3 ;
  assign n66 = pi9  & ~n65;
  assign n67 = pi0  & pi3 ;
  assign n68 = ~n66 & ~n67;
  assign n69 = ~pi1  & ~n68;
  assign n70 = pi1  & ~pi3 ;
  assign n71 = ~n69 & ~n70;
  assign n72 = ~n64 & n71;
  assign n73 = ~pi7  & ~n72;
  assign n74 = ~n55 & ~n73;
  assign n75 = ~pi8  & ~n74;
  assign n76 = ~n40 & ~n75;
  assign n77 = ~pi6  & ~n76;
  assign n78 = ~pi0  & ~pi2 ;
  assign n79 = n44 & n78;
  assign n80 = ~pi5  & ~n79;
  assign n81 = pi6  & ~n80;
  assign n82 = ~pi0  & ~pi9 ;
  assign n83 = pi0  & pi9 ;
  assign n84 = ~n82 & ~n83;
  assign n85 = ~n41 & ~n49;
  assign n86 = pi1  & pi5 ;
  assign n87 = pi2  & n86;
  assign n88 = pi1  & ~n1001;
  assign n89 = pi2  & n88;
  assign n90 = pi5  & n89;
  assign n91 = ~n1001 & n87;
  assign n92 = ~n81 & ~n1002;
  assign n93 = pi3  & ~n92;
  assign n94 = ~pi2  & ~n49;
  assign n95 = ~pi3  & n42;
  assign n96 = n94 & ~n95;
  assign n97 = ~pi6  & ~n94;
  assign n98 = pi5  & ~n97;
  assign n99 = pi6  & ~n94;
  assign n100 = pi1  & n65;
  assign n101 = n65 & n88;
  assign n102 = ~n1001 & n100;
  assign n103 = ~n99 & ~n1003;
  assign n104 = pi5  & ~n103;
  assign n105 = ~n96 & n98;
  assign n106 = pi2  & pi9 ;
  assign n107 = ~pi2  & n51;
  assign n108 = ~n106 & ~n107;
  assign n109 = ~pi0  & ~pi3 ;
  assign n110 = pi6  & n109;
  assign n111 = ~n108 & n109;
  assign n112 = pi6  & n111;
  assign n113 = ~n108 & n110;
  assign n114 = ~n1004 & ~n1005;
  assign n115 = ~n93 & n114;
  assign n116 = pi8  & ~n115;
  assign n117 = ~pi1  & ~n41;
  assign n118 = ~pi8  & ~n117;
  assign n119 = ~pi1  & pi2 ;
  assign n120 = n49 & n119;
  assign n121 = n27 & n57;
  assign n122 = ~n118 & ~n1006;
  assign n123 = pi3  & ~n122;
  assign n124 = pi1  & ~pi8 ;
  assign n125 = pi2  & ~pi3 ;
  assign n126 = n44 & n125;
  assign n127 = ~n124 & ~n126;
  assign n128 = ~pi0  & ~n127;
  assign n129 = ~pi1  & ~pi9 ;
  assign n130 = ~pi2  & pi6 ;
  assign n131 = pi3  & ~n130;
  assign n132 = n129 & ~n131;
  assign n133 = ~n106 & ~n132;
  assign n134 = ~pi8  & ~n133;
  assign n135 = ~n128 & ~n134;
  assign n136 = ~n123 & n135;
  assign n137 = ~pi5  & ~n136;
  assign n138 = ~pi8  & n129;
  assign n139 = ~pi0  & n65;
  assign n140 = ~pi3  & n78;
  assign n141 = n138 & n1007;
  assign n142 = ~n137 & ~n141;
  assign n143 = pi8  & ~n92;
  assign n144 = ~pi5  & ~n122;
  assign n145 = ~n143 & ~n144;
  assign n146 = pi3  & ~n145;
  assign n147 = ~pi5  & ~n135;
  assign n148 = pi8  & ~n114;
  assign n149 = ~n141 & ~n148;
  assign n150 = ~n141 & ~n147;
  assign n151 = ~n148 & n150;
  assign n152 = ~n147 & n149;
  assign n153 = ~n146 & n1008;
  assign n154 = ~n116 & n142;
  assign n155 = ~pi7  & ~n1009;
  assign n156 = ~n77 & ~n155;
  assign n157 = ~pi4  & ~n156;
  assign n158 = ~pi6  & pi8 ;
  assign n159 = pi5  & ~n158;
  assign n160 = pi4  & pi8 ;
  assign n161 = ~pi6  & ~pi9 ;
  assign n162 = ~n160 & ~n161;
  assign n163 = ~pi8  & ~pi9 ;
  assign n164 = ~pi6  & n163;
  assign n165 = pi6  & n160;
  assign n166 = ~n164 & ~n165;
  assign n167 = pi5  & ~n166;
  assign n168 = n159 & ~n162;
  assign n169 = pi6  & ~pi9 ;
  assign n170 = pi4  & pi9 ;
  assign n171 = ~n169 & ~n170;
  assign n172 = pi5  & pi6 ;
  assign n173 = ~pi8  & ~n172;
  assign n174 = ~n171 & ~n172;
  assign n175 = ~pi8  & n174;
  assign n176 = ~n171 & n173;
  assign n177 = ~n1010 & ~n1011;
  assign n178 = ~pi1  & ~pi3 ;
  assign n179 = ~pi7  & n78;
  assign n180 = n178 & n179;
  assign n181 = ~pi2  & n178;
  assign n182 = ~pi7  & ~n177;
  assign n183 = n181 & n182;
  assign n184 = ~pi0  & n183;
  assign n185 = ~n177 & n180;
  assign n186 = ~n157 & ~n1012;
  assign n187 = ~pi2  & ~pi8 ;
  assign n188 = n82 & n187;
  assign n189 = pi0  & pi8 ;
  assign n190 = pi8  & n83;
  assign n191 = pi9  & n189;
  assign n192 = pi2  & n1013;
  assign n193 = n106 & n189;
  assign n194 = ~n188 & ~n1014;
  assign n195 = pi5  & ~n194;
  assign n196 = ~pi5  & pi8 ;
  assign n197 = pi6  & pi9 ;
  assign n198 = ~n196 & ~n197;
  assign n199 = ~pi0  & ~n198;
  assign n200 = pi8  & pi9 ;
  assign n201 = ~pi8  & pi9 ;
  assign n202 = pi8  & ~pi9 ;
  assign n203 = ~n201 & ~n202;
  assign n204 = ~n163 & ~n200;
  assign n205 = pi5  & ~pi8 ;
  assign n206 = ~pi6  & pi9 ;
  assign n207 = ~n205 & ~n206;
  assign n208 = ~pi8  & n34;
  assign n209 = pi8  & n197;
  assign n210 = ~n208 & ~n209;
  assign n211 = n1015 & n207;
  assign n212 = ~n199 & n1016;
  assign n213 = pi2  & ~n212;
  assign n214 = ~n195 & ~n213;
  assign n215 = ~pi4  & ~n214;
  assign n216 = ~n160 & ~n205;
  assign n217 = ~pi6  & ~n216;
  assign n218 = ~n170 & ~n217;
  assign n219 = n78 & ~n206;
  assign n220 = ~n206 & ~n218;
  assign n221 = n78 & n220;
  assign n222 = ~n218 & n219;
  assign n223 = ~n215 & ~n1017;
  assign n224 = ~pi1  & ~n223;
  assign n225 = n56 & n201;
  assign n226 = pi6  & pi8 ;
  assign n227 = pi0  & ~n226;
  assign n228 = ~n198 & ~n226;
  assign n229 = pi0  & n228;
  assign n230 = ~n198 & n227;
  assign n231 = ~n225 & ~n1018;
  assign n232 = ~pi2  & ~n231;
  assign n233 = ~pi6  & ~pi8 ;
  assign n234 = ~pi0  & pi6 ;
  assign n235 = ~pi2  & ~n234;
  assign n236 = n196 & ~n235;
  assign n237 = ~n233 & ~n236;
  assign n238 = ~pi9  & ~n237;
  assign n239 = ~n232 & ~n238;
  assign n240 = pi1  & ~n239;
  assign n241 = n27 & n158;
  assign n242 = ~n240 & ~n241;
  assign n243 = ~pi4  & ~n242;
  assign n244 = ~pi1  & ~n214;
  assign n245 = ~n241 & ~n244;
  assign n246 = ~n240 & n245;
  assign n247 = ~pi4  & ~n246;
  assign n248 = ~pi1  & ~pi2 ;
  assign n249 = ~pi0  & n248;
  assign n250 = ~pi2  & n26;
  assign n251 = ~pi1  & n78;
  assign n252 = ~n206 & n1019;
  assign n253 = ~n218 & n252;
  assign n254 = ~n247 & ~n253;
  assign n255 = ~n224 & ~n243;
  assign n256 = ~pi3  & ~n1020;
  assign n257 = pi5  & n187;
  assign n258 = ~pi3  & ~pi8 ;
  assign n259 = ~n196 & ~n258;
  assign n260 = pi0  & n259;
  assign n261 = ~n257 & ~n260;
  assign n262 = ~pi1  & ~n261;
  assign n263 = pi3  & pi8 ;
  assign n264 = ~pi2  & ~n263;
  assign n265 = ~pi0  & ~n264;
  assign n266 = ~pi2  & pi8 ;
  assign n267 = pi0  & n266;
  assign n268 = pi0  & ~pi5 ;
  assign n269 = ~n56 & ~n268;
  assign n270 = ~n267 & n269;
  assign n271 = pi1  & ~n270;
  assign n272 = ~n265 & ~n271;
  assign n273 = ~n262 & n272;
  assign n274 = ~pi6  & ~n273;
  assign n275 = ~pi1  & pi6 ;
  assign n276 = pi2  & ~n275;
  assign n277 = ~pi1  & ~pi8 ;
  assign n278 = pi3  & ~n277;
  assign n279 = ~pi2  & ~n277;
  assign n280 = ~pi1  & pi8 ;
  assign n281 = pi6  & n280;
  assign n282 = ~n276 & ~n277;
  assign n283 = ~n279 & ~n281;
  assign n284 = pi3  & n1021;
  assign n285 = ~n276 & n278;
  assign n286 = ~pi0  & pi8 ;
  assign n287 = ~pi2  & ~n286;
  assign n288 = pi0  & pi1 ;
  assign n289 = ~pi1  & ~pi6 ;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~n286 & n290;
  assign n292 = ~pi2  & n291;
  assign n293 = n287 & n290;
  assign n294 = ~n1022 & ~n1023;
  assign n295 = ~pi5  & ~n294;
  assign n296 = ~pi9  & ~n295;
  assign n297 = ~n274 & n296;
  assign n298 = ~pi1  & pi3 ;
  assign n299 = pi3  & ~pi8 ;
  assign n300 = n248 & n299;
  assign n301 = n187 & n298;
  assign n302 = ~n86 & ~n1024;
  assign n303 = pi0  & ~n302;
  assign n304 = pi3  & n59;
  assign n305 = pi5  & ~n65;
  assign n306 = ~pi5  & ~n304;
  assign n307 = ~n65 & ~n306;
  assign n308 = ~n304 & ~n305;
  assign n309 = ~n303 & ~n1025;
  assign n310 = pi6  & ~n309;
  assign n311 = n205 & n304;
  assign n312 = pi9  & ~n311;
  assign n313 = ~n310 & n312;
  assign n314 = ~pi4  & ~n313;
  assign n315 = ~n274 & ~n295;
  assign n316 = ~pi9  & ~n315;
  assign n317 = ~n310 & ~n311;
  assign n318 = pi9  & ~n317;
  assign n319 = ~n316 & ~n318;
  assign n320 = ~pi4  & ~n319;
  assign n321 = ~n297 & n314;
  assign n322 = ~n256 & ~n1026;
  assign n323 = ~pi7  & ~n322;
  assign n324 = n51 & n266;
  assign n325 = n94 & ~n288;
  assign n326 = pi2  & ~n26;
  assign n327 = ~pi8  & ~n326;
  assign n328 = ~n325 & ~n326;
  assign n329 = ~pi8  & n328;
  assign n330 = ~n325 & n327;
  assign n331 = ~n324 & ~n1027;
  assign n332 = pi7  & ~n331;
  assign n333 = ~n28 & ~n332;
  assign n334 = ~pi6  & n43;
  assign n335 = ~pi4  & n334;
  assign n336 = ~pi4  & ~n333;
  assign n337 = ~pi6  & n336;
  assign n338 = n43 & n337;
  assign n339 = ~n333 & n335;
  assign n340 = ~n323 & ~n1028;
  assign n341 = ~n129 & n1015;
  assign n342 = n1015 & ~n277;
  assign n343 = pi2  & ~n1029;
  assign n344 = ~n163 & ~n1013;
  assign n345 = n1015 & ~n286;
  assign n346 = pi5  & n1030;
  assign n347 = ~pi5  & ~n106;
  assign n348 = pi1  & ~n347;
  assign n349 = ~pi5  & n106;
  assign n350 = pi5  & ~n286;
  assign n351 = pi5  & ~n1030;
  assign n352 = n1015 & n350;
  assign n353 = ~n349 & ~n1031;
  assign n354 = pi1  & ~n353;
  assign n355 = ~n346 & n348;
  assign n356 = ~n343 & ~n1032;
  assign n357 = ~pi3  & ~n356;
  assign n358 = n66 & n280;
  assign n359 = pi5  & ~n298;
  assign n360 = ~pi2  & n163;
  assign n361 = ~n359 & n360;
  assign n362 = ~n358 & ~n361;
  assign n363 = pi0  & ~n362;
  assign n364 = ~n357 & ~n363;
  assign n365 = ~pi6  & ~n364;
  assign n366 = pi6  & ~n44;
  assign n367 = ~n51 & ~n366;
  assign n368 = pi8  & ~n367;
  assign n369 = pi1  & pi9 ;
  assign n370 = ~n129 & ~n369;
  assign n371 = n258 & ~n370;
  assign n372 = ~n368 & ~n371;
  assign n373 = ~pi2  & ~n372;
  assign n374 = pi2  & n369;
  assign n375 = ~n280 & ~n374;
  assign n376 = pi6  & ~n375;
  assign n377 = pi8  & ~n27;
  assign n378 = pi2  & n163;
  assign n379 = ~n377 & ~n378;
  assign n380 = ~n376 & n379;
  assign n381 = pi3  & ~n380;
  assign n382 = ~n373 & ~n381;
  assign n383 = n268 & ~n382;
  assign n384 = ~n365 & ~n383;
  assign n385 = ~pi4  & ~n384;
  assign n386 = pi3  & ~n266;
  assign n387 = pi5  & ~n386;
  assign n388 = pi2  & ~pi5 ;
  assign n389 = pi3  & ~n388;
  assign n390 = pi8  & ~n389;
  assign n391 = ~n387 & ~n390;
  assign n392 = pi1  & ~n391;
  assign n393 = ~pi5  & pi6 ;
  assign n394 = ~pi3  & n393;
  assign n395 = ~pi8  & n393;
  assign n396 = n178 & n395;
  assign n397 = n277 & n394;
  assign n398 = ~n392 & ~n1033;
  assign n399 = ~pi9  & ~n398;
  assign n400 = pi1  & pi8 ;
  assign n401 = pi6  & ~n400;
  assign n402 = ~pi9  & ~n401;
  assign n403 = ~pi2  & ~n402;
  assign n404 = ~pi1  & n201;
  assign n405 = ~pi8  & n44;
  assign n406 = ~n403 & ~n1034;
  assign n407 = pi3  & ~n406;
  assign n408 = pi2  & ~n158;
  assign n409 = pi1  & ~n408;
  assign n410 = pi5  & ~n264;
  assign n411 = ~pi1  & ~n264;
  assign n412 = ~n408 & ~n411;
  assign n413 = pi5  & ~n412;
  assign n414 = ~n409 & n410;
  assign n415 = pi6  & ~pi8 ;
  assign n416 = ~pi3  & pi9 ;
  assign n417 = pi1  & n416;
  assign n418 = n415 & n417;
  assign n419 = ~n70 & ~n201;
  assign n420 = ~pi6  & ~n416;
  assign n421 = ~n416 & ~n419;
  assign n422 = ~pi6  & n421;
  assign n423 = ~n419 & n420;
  assign n424 = ~pi4  & ~n1036;
  assign n425 = ~n418 & n424;
  assign n426 = ~n1035 & n425;
  assign n427 = ~n407 & n426;
  assign n428 = ~n399 & n427;
  assign n429 = ~n202 & ~n233;
  assign n430 = ~n200 & ~n415;
  assign n431 = ~pi5  & ~n233;
  assign n432 = ~n202 & n431;
  assign n433 = ~pi5  & n1037;
  assign n434 = n181 & ~n1038;
  assign n435 = pi4  & ~n434;
  assign n436 = ~pi0  & ~n435;
  assign n437 = ~n418 & ~n1036;
  assign n438 = ~n1035 & n437;
  assign n439 = ~n407 & n438;
  assign n440 = ~n407 & ~n418;
  assign n441 = ~n1035 & n440;
  assign n442 = ~n399 & n441;
  assign n443 = ~n1036 & n442;
  assign n444 = ~n399 & n439;
  assign n445 = ~pi4  & ~n1039;
  assign n446 = ~pi3  & pi4 ;
  assign n447 = pi4  & n65;
  assign n448 = ~pi2  & n446;
  assign n449 = ~pi1  & n1040;
  assign n450 = ~pi1  & n446;
  assign n451 = ~n1038 & n450;
  assign n452 = ~pi2  & n451;
  assign n453 = ~n1038 & n449;
  assign n454 = ~n445 & ~n1041;
  assign n455 = ~pi0  & ~n454;
  assign n456 = ~n428 & n436;
  assign n457 = ~n385 & ~n1042;
  assign n458 = ~pi7  & ~n457;
  assign n459 = pi7  & n200;
  assign n460 = pi0  & ~n459;
  assign n461 = n23 & n83;
  assign n462 = ~n82 & ~n461;
  assign n463 = pi1  & ~n462;
  assign n464 = n42 & ~n460;
  assign n465 = n49 & n277;
  assign n466 = ~n1043 & ~n465;
  assign n467 = ~pi5  & ~pi6 ;
  assign n468 = ~pi4  & n65;
  assign n469 = n467 & n468;
  assign n470 = ~pi4  & ~n466;
  assign n471 = n65 & n470;
  assign n472 = n467 & n471;
  assign n473 = ~n466 & n469;
  assign n474 = ~n458 & ~n1044;
  assign n475 = pi2  & ~n259;
  assign n476 = ~pi2  & pi5 ;
  assign n477 = pi5  & pi8 ;
  assign n478 = ~pi2  & n477;
  assign n479 = pi5  & n266;
  assign n480 = pi8  & n476;
  assign n481 = ~n475 & ~n1045;
  assign n482 = ~pi9  & ~n481;
  assign n483 = pi5  & pi9 ;
  assign n484 = ~pi8  & n483;
  assign n485 = pi5  & n201;
  assign n486 = ~pi3  & ~n1046;
  assign n487 = ~pi2  & ~n486;
  assign n488 = ~pi6  & ~n299;
  assign n489 = pi3  & ~pi5 ;
  assign n490 = ~n488 & ~n489;
  assign n491 = ~n487 & ~n490;
  assign n492 = ~n482 & n491;
  assign n493 = pi1  & ~n492;
  assign n494 = n257 & n289;
  assign n495 = ~n394 & ~n494;
  assign n496 = ~pi9  & ~n495;
  assign n497 = ~n493 & ~n496;
  assign n498 = pi0  & ~n497;
  assign n499 = ~n163 & ~n483;
  assign n500 = pi2  & ~n499;
  assign n501 = ~pi3  & ~n415;
  assign n502 = ~n500 & n501;
  assign n503 = pi1  & ~n159;
  assign n504 = n206 & n477;
  assign n505 = ~n208 & ~n504;
  assign n506 = pi2  & ~n505;
  assign n507 = pi3  & ~n159;
  assign n508 = ~n395 & ~n507;
  assign n509 = ~n506 & n508;
  assign n510 = pi1  & ~n509;
  assign n511 = ~n502 & n503;
  assign n512 = pi6  & n388;
  assign n513 = pi2  & n393;
  assign n514 = pi6  & ~n65;
  assign n515 = pi3  & ~pi9 ;
  assign n516 = pi3  & ~n206;
  assign n517 = pi2  & pi6 ;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~n514 & ~n515;
  assign n520 = ~pi1  & ~n1049;
  assign n521 = ~n1048 & ~n520;
  assign n522 = ~n1047 & n521;
  assign n523 = ~pi0  & ~n522;
  assign n524 = pi3  & ~pi6 ;
  assign n525 = pi2  & n524;
  assign n526 = ~n65 & n393;
  assign n527 = ~n525 & ~n526;
  assign n528 = pi9  & ~n527;
  assign n529 = ~pi9  & n393;
  assign n530 = ~n524 & ~n529;
  assign n531 = ~pi8  & ~n530;
  assign n532 = ~n528 & ~n531;
  assign n533 = ~pi1  & ~n532;
  assign n534 = pi1  & n202;
  assign n535 = n393 & n534;
  assign n536 = n400 & n529;
  assign n537 = ~n34 & ~n233;
  assign n538 = ~pi2  & ~n537;
  assign n539 = ~pi6  & ~n483;
  assign n540 = ~n369 & ~n477;
  assign n541 = n539 & ~n540;
  assign n542 = ~n538 & ~n541;
  assign n543 = pi3  & ~n542;
  assign n544 = ~n1050 & ~n543;
  assign n545 = ~n533 & n544;
  assign n546 = ~n523 & n545;
  assign n547 = ~n498 & n546;
  assign n548 = ~pi4  & ~n547;
  assign n549 = ~n172 & ~n467;
  assign n550 = n446 & ~n549;
  assign n551 = ~pi5  & ~n200;
  assign n552 = n1019 & ~n551;
  assign n553 = n550 & n552;
  assign n554 = ~pi4  & ~n1049;
  assign n555 = n1040 & ~n551;
  assign n556 = n200 & n467;
  assign n557 = ~n172 & ~n556;
  assign n558 = n1040 & ~n557;
  assign n559 = ~n549 & n555;
  assign n560 = ~n554 & ~n1051;
  assign n561 = ~pi1  & ~n560;
  assign n562 = ~n1047 & ~n1048;
  assign n563 = ~pi4  & ~n562;
  assign n564 = ~n561 & ~n563;
  assign n565 = ~pi0  & ~n564;
  assign n566 = ~n498 & n545;
  assign n567 = ~pi4  & ~n566;
  assign n568 = ~n565 & ~n567;
  assign n569 = ~n548 & ~n553;
  assign po3  = ~pi7  & ~n1052;
  assign n571 = ~pi1  & pi4 ;
  assign n572 = n1007 & n571;
  assign n573 = n26 & n1040;
  assign n574 = n1019 & n446;
  assign n575 = ~n172 & ~n1053;
  assign n576 = ~pi7  & ~n575;
  assign n577 = ~pi1  & ~pi5 ;
  assign n578 = pi2  & ~n577;
  assign n579 = ~pi9  & ~n578;
  assign n580 = ~pi6  & n579;
  assign n581 = n161 & ~n578;
  assign n582 = pi5  & n369;
  assign n583 = ~n1054 & ~n582;
  assign n584 = pi0  & ~n583;
  assign n585 = ~pi0  & pi2 ;
  assign n586 = ~pi0  & ~n34;
  assign n587 = pi2  & n586;
  assign n588 = ~n34 & n585;
  assign n589 = ~n584 & ~n1055;
  assign n590 = pi8  & ~n589;
  assign n591 = pi2  & n41;
  assign n592 = pi9  & n585;
  assign n593 = ~n138 & ~n1056;
  assign n594 = pi5  & ~n593;
  assign n595 = ~pi2  & ~pi9 ;
  assign n596 = ~pi2  & pi9 ;
  assign n597 = ~n27 & ~n596;
  assign n598 = ~n106 & ~n595;
  assign n599 = pi2  & pi8 ;
  assign n600 = ~n187 & ~n599;
  assign n601 = pi6  & ~n600;
  assign n602 = pi6  & n1015;
  assign n603 = n1057 & n602;
  assign n604 = pi6  & n1057;
  assign n605 = ~n600 & n604;
  assign n606 = n1057 & n601;
  assign n607 = ~n594 & ~n1058;
  assign n608 = ~n590 & ~n594;
  assign n609 = ~n1058 & n608;
  assign n610 = ~n590 & n607;
  assign n611 = ~pi3  & ~n1059;
  assign n612 = ~pi0  & ~pi6 ;
  assign n613 = ~n277 & n612;
  assign n614 = ~n59 & ~n613;
  assign n615 = n370 & ~n614;
  assign n616 = ~pi1  & ~n163;
  assign n617 = pi0  & ~n51;
  assign n618 = ~n138 & ~n369;
  assign n619 = pi0  & ~n618;
  assign n620 = ~n616 & n617;
  assign n621 = pi2  & n51;
  assign n622 = ~n1060 & ~n621;
  assign n623 = ~n277 & n370;
  assign n624 = n612 & n623;
  assign n625 = n622 & ~n624;
  assign n626 = ~n615 & ~n1060;
  assign n627 = ~pi5  & ~n1061;
  assign n628 = pi0  & n226;
  assign n629 = ~pi2  & n628;
  assign n630 = ~n124 & ~n629;
  assign n631 = pi9  & ~n585;
  assign n632 = n124 & ~n585;
  assign n633 = ~pi8  & n288;
  assign n634 = ~n124 & ~n628;
  assign n635 = ~pi2  & ~n634;
  assign n636 = ~n633 & ~n635;
  assign n637 = ~n629 & ~n632;
  assign n638 = pi9  & ~n1062;
  assign n639 = ~n630 & n631;
  assign n640 = ~pi0  & ~pi8 ;
  assign n641 = n51 & ~n268;
  assign n642 = ~n268 & ~n640;
  assign n643 = n51 & n642;
  assign n644 = ~n640 & n641;
  assign n645 = ~n1063 & ~n1064;
  assign n646 = ~n627 & n645;
  assign n647 = pi3  & ~n646;
  assign n648 = ~n1001 & n476;
  assign n649 = ~pi6  & ~n388;
  assign n650 = n41 & ~n649;
  assign n651 = ~n648 & ~n650;
  assign n652 = ~pi8  & ~n651;
  assign n653 = pi2  & ~n163;
  assign n654 = ~n1013 & ~n653;
  assign n655 = pi6  & ~n654;
  assign n656 = ~n652 & ~n655;
  assign n657 = pi1  & ~n656;
  assign n658 = n41 & n599;
  assign n659 = ~pi0  & ~n415;
  assign n660 = ~n477 & n595;
  assign n661 = ~pi8  & ~n612;
  assign n662 = ~n268 & ~n661;
  assign n663 = ~pi9  & ~n662;
  assign n664 = ~pi2  & n663;
  assign n665 = pi8  & ~n268;
  assign n666 = n595 & ~n612;
  assign n667 = ~n665 & n666;
  assign n668 = ~n659 & n660;
  assign n669 = ~n658 & ~n1065;
  assign n670 = ~pi1  & ~n669;
  assign n671 = ~n657 & ~n670;
  assign n672 = ~n647 & n671;
  assign n673 = ~n611 & n672;
  assign n674 = ~pi7  & ~n673;
  assign n675 = pi7  & ~pi9 ;
  assign n676 = pi8  & ~n675;
  assign n677 = n119 & ~n676;
  assign n678 = ~n107 & ~n677;
  assign n679 = ~pi0  & ~n678;
  assign n680 = pi1  & n1013;
  assign n681 = n189 & n369;
  assign n682 = ~n163 & ~n1066;
  assign n683 = ~pi2  & pi7 ;
  assign n684 = pi7  & ~n682;
  assign n685 = ~pi2  & n684;
  assign n686 = ~n682 & n683;
  assign n687 = ~n679 & ~n1067;
  assign n688 = n334 & ~n687;
  assign n689 = ~pi7  & ~n1059;
  assign n690 = n467 & ~n687;
  assign n691 = ~n689 & ~n690;
  assign n692 = ~pi3  & ~n691;
  assign n693 = ~pi7  & ~n672;
  assign n694 = ~n692 & ~n693;
  assign n695 = ~n674 & ~n688;
  assign n696 = ~pi4  & ~n1068;
  assign po6  = ~n576 & ~n696;
  assign n698 = n286 & n524;
  assign n699 = ~n415 & ~n698;
  assign n700 = pi9  & ~n699;
  assign n701 = ~pi3  & pi8 ;
  assign n702 = ~n197 & ~n701;
  assign n703 = pi3  & ~n197;
  assign n704 = pi0  & ~n163;
  assign n705 = ~n233 & n704;
  assign n706 = ~n703 & n705;
  assign n707 = pi0  & ~n702;
  assign n708 = ~pi9  & n226;
  assign n709 = pi6  & n202;
  assign n710 = pi8  & n169;
  assign n711 = ~n1069 & ~n1070;
  assign n712 = ~n700 & ~n1070;
  assign n713 = ~n1069 & n712;
  assign n714 = ~n700 & n711;
  assign n715 = ~pi2  & ~n1071;
  assign n716 = ~pi3  & n164;
  assign n717 = n161 & n258;
  assign n718 = pi3  & ~n200;
  assign n719 = ~n189 & ~n718;
  assign n720 = ~pi6  & ~n719;
  assign n721 = ~pi3  & n200;
  assign n722 = pi8  & n416;
  assign n723 = ~n720 & ~n1073;
  assign n724 = pi2  & ~n723;
  assign n725 = ~n1072 & ~n724;
  assign n726 = ~n715 & ~n1072;
  assign n727 = ~n724 & n726;
  assign n728 = ~n715 & n725;
  assign n729 = pi1  & ~n1074;
  assign n730 = ~pi0  & n602;
  assign n731 = n1015 & n234;
  assign n732 = ~pi6  & ~n200;
  assign n733 = ~n82 & ~n201;
  assign n734 = ~pi6  & ~n733;
  assign n735 = ~pi2  & n734;
  assign n736 = ~pi2  & ~pi6 ;
  assign n737 = ~n733 & n736;
  assign n738 = n94 & n732;
  assign n739 = ~n1075 & ~n1076;
  assign n740 = pi3  & ~n739;
  assign n741 = ~pi0  & n187;
  assign n742 = ~n628 & ~n741;
  assign n743 = ~pi9  & ~n742;
  assign n744 = ~pi6  & ~n258;
  assign n745 = n653 & ~n744;
  assign n746 = ~n743 & ~n745;
  assign n747 = ~n740 & n746;
  assign n748 = ~pi1  & ~n747;
  assign n749 = ~pi2  & n169;
  assign n750 = ~pi2  & pi3 ;
  assign n751 = ~pi9  & n415;
  assign n752 = n750 & n751;
  assign n753 = pi3  & n187;
  assign n754 = n169 & n753;
  assign n755 = n299 & n749;
  assign n756 = ~n748 & ~n1077;
  assign n757 = ~n729 & n756;
  assign n758 = ~pi5  & ~n757;
  assign n759 = pi0  & ~n1057;
  assign n760 = pi5  & ~pi9 ;
  assign n761 = ~pi0  & n760;
  assign n762 = ~pi9  & n56;
  assign n763 = ~n759 & ~n1078;
  assign n764 = pi8  & ~n763;
  assign n765 = pi2  & n1046;
  assign n766 = n106 & n205;
  assign n767 = ~n764 & ~n1079;
  assign n768 = ~pi3  & ~n767;
  assign n769 = pi3  & pi5 ;
  assign n770 = ~n27 & ~n769;
  assign n771 = pi2  & ~n640;
  assign n772 = ~n200 & ~n771;
  assign n773 = pi3  & n476;
  assign n774 = ~pi0  & ~n770;
  assign n775 = ~n773 & ~n774;
  assign n776 = ~pi8  & ~n775;
  assign n777 = n750 & n760;
  assign n778 = ~n776 & ~n777;
  assign n779 = n640 & ~n770;
  assign n780 = ~n773 & ~n779;
  assign n781 = ~n200 & ~n780;
  assign n782 = ~n770 & n772;
  assign n783 = ~n768 & n1080;
  assign n784 = pi1  & ~n783;
  assign n785 = n67 & n378;
  assign n786 = pi2  & pi3 ;
  assign n787 = ~n1015 & ~n786;
  assign n788 = ~pi2  & ~n67;
  assign n789 = pi5  & ~n788;
  assign n790 = n1015 & ~n788;
  assign n791 = ~n786 & ~n790;
  assign n792 = pi5  & ~n791;
  assign n793 = ~n787 & n789;
  assign n794 = ~n785 & ~n1081;
  assign n795 = ~pi1  & ~n794;
  assign n796 = pi8  & n483;
  assign n797 = n786 & n796;
  assign n798 = ~n795 & ~n797;
  assign n799 = ~n784 & n798;
  assign n800 = ~pi6  & ~n799;
  assign n801 = ~n758 & ~n800;
  assign n802 = ~pi7  & ~n801;
  assign n803 = pi2  & ~n1015;
  assign n804 = ~pi0  & n803;
  assign n805 = ~n1015 & n585;
  assign n806 = ~pi9  & n23;
  assign n807 = n37 & n806;
  assign n808 = n267 & n675;
  assign n809 = ~n1082 & ~n1083;
  assign n810 = n43 & n289;
  assign n811 = n178 & n467;
  assign n812 = n289 & ~n809;
  assign n813 = n43 & n812;
  assign n814 = ~n809 & n1084;
  assign n815 = ~n802 & ~n1085;
  assign n816 = ~pi4  & ~n815;
  assign n817 = n60 & n109;
  assign n818 = pi4  & ~pi7 ;
  assign n819 = n289 & n818;
  assign n820 = n43 & n818;
  assign n821 = ~pi5  & ~pi7 ;
  assign n822 = n1053 & n821;
  assign n823 = n1019 & n820;
  assign n824 = ~pi6  & n1086;
  assign n825 = n817 & n819;
  assign po7  = ~n816 & ~n1087;
  assign n827 = n178 & n268;
  assign n828 = n43 & n57;
  assign n829 = ~pi1  & pi5 ;
  assign n830 = ~n43 & ~n829;
  assign n831 = ~n86 & ~n489;
  assign n832 = ~pi2  & ~n109;
  assign n833 = ~n109 & ~n1089;
  assign n834 = ~pi2  & n833;
  assign n835 = ~n1089 & n832;
  assign n836 = ~n1088 & ~n1090;
  assign n837 = pi8  & ~n836;
  assign n838 = ~pi5  & ~n286;
  assign n839 = n59 & ~n769;
  assign n840 = ~n769 & ~n838;
  assign n841 = n59 & n840;
  assign n842 = ~n838 & n839;
  assign n843 = ~n837 & ~n1091;
  assign n844 = ~pi9  & ~n843;
  assign n845 = ~pi2  & ~n129;
  assign n846 = ~n416 & n845;
  assign n847 = ~n129 & ~n416;
  assign n848 = ~n1089 & n847;
  assign n849 = ~pi2  & n848;
  assign n850 = ~n1089 & n846;
  assign n851 = n370 & ~n577;
  assign n852 = n125 & ~n851;
  assign n853 = n248 & n760;
  assign n854 = n129 & n476;
  assign n855 = ~n417 & ~n1093;
  assign n856 = ~pi0  & ~n855;
  assign n857 = ~n852 & ~n856;
  assign n858 = ~n1092 & ~n852;
  assign n859 = ~n856 & n858;
  assign n860 = ~n1092 & n857;
  assign n861 = ~pi8  & ~n1094;
  assign n862 = ~n388 & ~n769;
  assign n863 = pi1  & ~n386;
  assign n864 = ~n386 & ~n862;
  assign n865 = pi1  & n864;
  assign n866 = ~n862 & n863;
  assign n867 = ~n56 & n266;
  assign n868 = ~n56 & n298;
  assign n869 = n266 & n868;
  assign n870 = n298 & n867;
  assign n871 = ~n1095 & ~n1096;
  assign n872 = pi9  & ~n871;
  assign n873 = ~n861 & ~n872;
  assign n874 = ~n844 & ~n872;
  assign n875 = ~n861 & n874;
  assign n876 = ~n844 & n873;
  assign n877 = ~pi6  & ~n1097;
  assign n878 = ~n51 & n286;
  assign n879 = n366 & ~n878;
  assign n880 = ~pi2  & ~n879;
  assign n881 = pi0  & ~n616;
  assign n882 = ~pi6  & ~n124;
  assign n883 = ~n881 & n882;
  assign n884 = n489 & ~n883;
  assign n885 = pi2  & ~n616;
  assign n886 = ~n366 & ~n885;
  assign n887 = pi0  & ~n886;
  assign n888 = pi2  & ~n882;
  assign n889 = pi6  & ~n200;
  assign n890 = pi8  & ~n51;
  assign n891 = n366 & ~n890;
  assign n892 = ~n616 & n889;
  assign n893 = ~n888 & ~n1098;
  assign n894 = ~n887 & n893;
  assign n895 = n489 & ~n894;
  assign n896 = ~n880 & n884;
  assign n897 = ~n877 & ~n1099;
  assign n898 = ~pi7  & ~n897;
  assign n899 = ~pi0  & ~n600;
  assign n900 = ~n267 & ~n899;
  assign n901 = ~pi9  & ~n900;
  assign n902 = ~pi8  & n1056;
  assign n903 = n106 & n640;
  assign n904 = ~n901 & ~n1100;
  assign n905 = ~pi1  & ~n904;
  assign n906 = n369 & n741;
  assign n907 = ~n905 & ~n906;
  assign n908 = n43 & ~n907;
  assign n909 = ~pi6  & n908;
  assign n910 = n334 & ~n907;
  assign n911 = ~n898 & ~n1101;
  assign n912 = ~pi4  & ~n911;
  assign po8  = ~n1086 & ~n912;
  assign n914 = n286 & ~n539;
  assign n915 = n703 & ~n914;
  assign n916 = n446 & ~n467;
  assign n917 = ~pi2  & ~n916;
  assign n918 = ~n197 & ~n914;
  assign n919 = pi3  & ~n918;
  assign n920 = pi4  & ~n467;
  assign n921 = ~pi3  & ~n920;
  assign n922 = ~n919 & ~n921;
  assign n923 = ~pi2  & ~n922;
  assign n924 = ~n915 & n917;
  assign n925 = ~pi3  & ~n551;
  assign n926 = ~pi3  & ~n34;
  assign n927 = ~pi8  & ~n483;
  assign n928 = n926 & ~n927;
  assign n929 = pi2  & n928;
  assign n930 = n653 & n925;
  assign n931 = ~n1102 & ~n1103;
  assign n932 = ~pi1  & ~n931;
  assign n933 = n34 & ~n286;
  assign n934 = ~pi3  & ~n933;
  assign n935 = n41 & n226;
  assign n936 = n286 & ~n703;
  assign n937 = ~n926 & ~n936;
  assign n938 = ~n934 & ~n935;
  assign n939 = ~pi2  & ~n1104;
  assign n940 = ~n200 & n525;
  assign n941 = ~pi5  & n940;
  assign n942 = n525 & n551;
  assign n943 = ~pi6  & ~n796;
  assign n944 = ~pi3  & ~n943;
  assign n945 = ~n1105 & ~n944;
  assign n946 = ~n939 & n945;
  assign n947 = pi1  & ~n946;
  assign n948 = n268 & n525;
  assign n949 = ~pi7  & ~n948;
  assign n950 = ~n616 & ~n949;
  assign n951 = ~pi7  & ~n181;
  assign n952 = pi0  & ~n951;
  assign n953 = ~pi5  & ~n125;
  assign n954 = pi6  & ~n953;
  assign n955 = pi4  & ~n181;
  assign n956 = pi7  & ~n125;
  assign n957 = ~n955 & ~n956;
  assign n958 = ~n954 & ~n956;
  assign n959 = ~n955 & n958;
  assign n960 = ~n954 & n957;
  assign n961 = ~n952 & n1106;
  assign n962 = ~n950 & n961;
  assign n963 = ~n947 & n962;
  assign n964 = ~n932 & ~n954;
  assign n965 = ~n947 & n964;
  assign n966 = ~n956 & n965;
  assign n967 = ~n952 & n966;
  assign n968 = ~n950 & n967;
  assign n969 = ~n955 & n968;
  assign n970 = ~n932 & n963;
  assign n971 = pi8  & ~n42;
  assign n972 = pi3  & ~pi4 ;
  assign n973 = pi2  & n972;
  assign n974 = ~n50 & n973;
  assign n975 = ~pi8  & ~n50;
  assign n976 = ~n42 & ~n975;
  assign n977 = n972 & ~n976;
  assign n978 = pi2  & n977;
  assign n979 = ~n971 & n974;
  assign n980 = ~n1053 & ~n1108;
  assign n981 = ~pi7  & n467;
  assign n982 = ~pi7  & ~n980;
  assign n983 = n467 & n982;
  assign n984 = ~n980 & n981;
  assign n985 = ~pi4  & n326;
  assign n986 = ~n446 & ~n972;
  assign n987 = n1019 & ~n986;
  assign n988 = ~n985 & ~n987;
  assign n989 = ~pi7  & n172;
  assign n990 = ~pi7  & ~n988;
  assign n991 = n172 & n990;
  assign n992 = ~n988 & n989;
  assign n993 = ~n1019 & n972;
  assign n994 = ~n1053 & ~n993;
  assign n995 = ~pi7  & ~n994;
  assign n996 = n172 & n995;
  assign n997 = n989 & ~n994;
  assign n998 = n24 | n25;
  assign n999 = n47 | n48;
  assign n1000 = n62 | n63;
  assign n1001 = n84 | ~n85;
  assign n1002 = n90 | n91;
  assign n1003 = n101 | n102;
  assign n1004 = n104 | n105;
  assign n1005 = n112 | n113;
  assign n1006 = n120 | n121;
  assign n1007 = n139 | n140;
  assign n1008 = n151 | n152;
  assign n1009 = n153 | n154;
  assign n1010 = n167 | n168;
  assign n1011 = n175 | n176;
  assign n1012 = n184 | n185;
  assign n1013 = n190 | n191;
  assign n1014 = n192 | n193;
  assign n1015 = n203 | ~n204;
  assign n1016 = n210 | ~n211;
  assign n1017 = n221 | n222;
  assign n1018 = n229 | n230;
  assign n1019 = n251 | n249 | n250;
  assign n1020 = n254 | n255;
  assign n1021 = n282 | ~n283;
  assign n1022 = n284 | n285;
  assign n1023 = n292 | n293;
  assign n1024 = n300 | n301;
  assign n1025 = n307 | ~n308;
  assign n1026 = n320 | n321;
  assign n1027 = n329 | n330;
  assign n1028 = n338 | n339;
  assign n1029 = n341 | n342;
  assign n1030 = n344 | ~n345;
  assign n1031 = n351 | n352;
  assign n1032 = n354 | n355;
  assign n1033 = n396 | n397;
  assign n1034 = n404 | n405;
  assign n1035 = n413 | n414;
  assign n1036 = n422 | n423;
  assign n1037 = n429 | ~n430;
  assign n1038 = n432 | n433;
  assign n1039 = n443 | n444;
  assign n1040 = n447 | n448;
  assign n1041 = n452 | n453;
  assign n1042 = n455 | n456;
  assign n1043 = n463 | n464;
  assign n1044 = n472 | n473;
  assign n1045 = n480 | n478 | n479;
  assign n1046 = n484 | n485;
  assign n1047 = n510 | n511;
  assign n1048 = n512 | n513;
  assign n1049 = n518 | n519;
  assign n1050 = n535 | n536;
  assign n1051 = n558 | n559;
  assign n1052 = n568 | n569;
  assign n1053 = n574 | n572 | n573;
  assign n1054 = n580 | n581;
  assign n1055 = n587 | n588;
  assign n1056 = n591 | n592;
  assign n1057 = n597 | ~n598;
  assign n1058 = n606 | n603 | n605;
  assign n1059 = n609 | n610;
  assign n1060 = n619 | n620;
  assign n1061 = n625 | n626;
  assign n1062 = n636 | n637;
  assign n1063 = n638 | n639;
  assign n1064 = n643 | n644;
  assign n1065 = n668 | n664 | n667;
  assign n1066 = n680 | n681;
  assign n1067 = n685 | n686;
  assign n1068 = n694 | n695;
  assign n1069 = n706 | n707;
  assign n1070 = n710 | n708 | n709;
  assign n1071 = n713 | n714;
  assign n1072 = n716 | n717;
  assign n1073 = n721 | n722;
  assign n1074 = n727 | n728;
  assign n1075 = n730 | n731;
  assign n1076 = n738 | n735 | n737;
  assign n1077 = n755 | n752 | n754;
  assign n1078 = n761 | n762;
  assign n1079 = n765 | n766;
  assign n1080 = ~n782 | n778 | ~n781;
  assign n1081 = n792 | n793;
  assign n1082 = n804 | n805;
  assign n1083 = n807 | n808;
  assign n1084 = n810 | n811;
  assign n1085 = n813 | n814;
  assign n1086 = n822 | n823;
  assign n1087 = n824 | n825;
  assign n1088 = n827 | n828;
  assign n1089 = n830 | ~n831;
  assign n1090 = n834 | n835;
  assign n1091 = n841 | n842;
  assign n1092 = n849 | n850;
  assign n1093 = n853 | n854;
  assign n1094 = n859 | n860;
  assign n1095 = n865 | n866;
  assign n1096 = n869 | n870;
  assign n1097 = n875 | n876;
  assign n1098 = n891 | n892;
  assign n1099 = n895 | n896;
  assign n1100 = n902 | n903;
  assign n1101 = n909 | n910;
  assign n1102 = n923 | n924;
  assign n1103 = n929 | n930;
  assign n1104 = n937 | n938;
  assign n1105 = n941 | n942;
  assign n1106 = n959 | n960;
  assign po9  = n969 | n970;
  assign n1108 = n978 | n979;
  assign po10  = n983 | n984;
  assign po4  = n991 | n992;
  assign po5  = n996 | n997;
  assign po0  = ~n186;
  assign po1  = ~n340;
  assign po2  = ~n474;
endmodule
