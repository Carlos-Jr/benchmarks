module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29,
    n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n485, n486, n488, n489,
    n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n644, n645,
    n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n674,
    n675, n676;
  assign n23 = pi00 & pi11;
  assign n24 = ~pi08 & ~pi09;
  assign n25 = ~pi10 & ~n24;
  assign n26 = n23 & ~n25;
  assign n27 = pi08 & ~pi10;
  assign n28 = pi04 & n27;
  assign n29 = ~pi00 & pi11;
  assign n30 = n28 & n29;
  assign n31 = ~pi08 & pi10;
  assign n32 = ~pi10 & ~pi11;
  assign n33 = pi08 & n32;
  assign n34 = ~n31 & ~n33;
  assign n35 = pi09 & pi11;
  assign n36 = ~pi10 & ~pi13;
  assign n37 = ~n35 & n36;
  assign n38 = ~pi08 & n37;
  assign n39 = ~pi00 & n38;
  assign n40 = ~pi00 & ~pi04;
  assign n41 = ~pi10 & pi13;
  assign n42 = pi08 & ~pi09;
  assign n43 = ~pi13 & ~n32;
  assign n44 = ~n41 & n42;
  assign n45 = ~n43 & n44;
  assign n46 = ~n40 & n45;
  assign n47 = pi08 & pi09;
  assign n48 = ~n24 & ~n47;
  assign n49 = ~pi10 & pi11;
  assign n50 = ~n48 & n49;
  assign n51 = pi13 & n50;
  assign n52 = ~pi09 & ~pi11;
  assign n53 = n31 & n52;
  assign n54 = ~n51 & ~n53;
  assign n55 = pi00 & pi04;
  assign n56 = ~n54 & n55;
  assign n57 = pi10 & ~pi11;
  assign n58 = ~pi08 & pi09;
  assign n59 = pi13 & n58;
  assign n60 = ~n57 & n59;
  assign n61 = n47 & n57;
  assign n62 = ~pi09 & pi11;
  assign n63 = pi08 & pi10;
  assign n64 = ~pi13 & n62;
  assign n65 = n63 & n64;
  assign n66 = ~n60 & ~n61;
  assign n67 = ~n65 & n66;
  assign n68 = ~pi04 & ~n67;
  assign n69 = ~n40 & ~n55;
  assign n70 = ~pi00 & ~n57;
  assign n71 = n59 & n69;
  assign n72 = ~n70 & n71;
  assign n73 = ~n46 & ~n72;
  assign n74 = ~n56 & n73;
  assign n75 = ~n68 & n74;
  assign n76 = ~n39 & n75;
  assign n77 = ~n34 & n76;
  assign n78 = pi08 & n57;
  assign n79 = ~n23 & ~n78;
  assign n80 = ~pi04 & ~n79;
  assign n81 = ~n30 & ~n80;
  assign n82 = ~n77 & n81;
  assign n83 = ~pi09 & ~n82;
  assign n84 = ~pi08 & pi11;
  assign n85 = pi04 & n84;
  assign n86 = pi00 & ~n75;
  assign n87 = n63 & n86;
  assign n88 = ~pi08 & n57;
  assign n89 = n40 & n88;
  assign n90 = ~pi11 & ~n31;
  assign n91 = n55 & ~n90;
  assign n92 = ~n85 & ~n89;
  assign n93 = ~n91 & n92;
  assign n94 = ~n87 & n93;
  assign n95 = pi09 & ~n94;
  assign n96 = ~pi08 & ~pi10;
  assign n97 = pi04 & n96;
  assign n98 = ~pi09 & ~n27;
  assign n99 = ~n57 & n98;
  assign n100 = ~n97 & ~n99;
  assign n101 = ~n76 & ~n100;
  assign n102 = ~n26 & ~n101;
  assign n103 = ~n83 & n102;
  assign n104 = ~n95 & n103;
  assign n105 = ~pi13 & ~n104;
  assign n106 = ~pi10 & n47;
  assign n107 = ~pi11 & pi13;
  assign n108 = n106 & n107;
  assign n109 = ~pi09 & pi10;
  assign n110 = ~pi13 & n84;
  assign n111 = n109 & n110;
  assign n112 = ~n108 & ~n111;
  assign n113 = pi10 & n47;
  assign n114 = n29 & n113;
  assign n115 = n47 & n49;
  assign n116 = n57 & n58;
  assign n117 = ~n115 & ~n116;
  assign n118 = n23 & ~n47;
  assign n119 = ~pi08 & pi13;
  assign n120 = n35 & n119;
  assign n121 = ~pi10 & n120;
  assign n122 = n55 & n121;
  assign n123 = ~pi00 & n76;
  assign n124 = n120 & ~n123;
  assign n125 = pi13 & n57;
  assign n126 = n24 & n76;
  assign n127 = n47 & n86;
  assign n128 = n42 & n55;
  assign n129 = ~n126 & ~n128;
  assign n130 = ~n127 & n129;
  assign n131 = n125 & ~n130;
  assign n132 = ~n124 & ~n131;
  assign n133 = n42 & n125;
  assign n134 = n132 & n133;
  assign n135 = ~n122 & ~n134;
  assign n136 = pi08 & n52;
  assign n137 = ~n135 & n136;
  assign n138 = ~n118 & ~n137;
  assign n139 = pi10 & ~n138;
  assign n140 = n117 & ~n139;
  assign n141 = n76 & ~n140;
  assign n142 = n49 & n58;
  assign n143 = ~n135 & n142;
  assign n144 = ~n61 & ~n143;
  assign n145 = n132 & ~n144;
  assign n146 = n135 & n142;
  assign n147 = ~pi00 & n53;
  assign n148 = ~n146 & ~n147;
  assign n149 = ~n132 & ~n148;
  assign n150 = n42 & n57;
  assign n151 = n135 & n150;
  assign n152 = ~n25 & n29;
  assign n153 = ~n151 & ~n152;
  assign n154 = ~n76 & ~n153;
  assign n155 = pi00 & ~pi08;
  assign n156 = n132 & n155;
  assign n157 = ~n28 & ~n156;
  assign n158 = n52 & ~n157;
  assign n159 = ~pi09 & n27;
  assign n160 = n69 & n159;
  assign n161 = ~pi09 & n76;
  assign n162 = pi11 & ~n161;
  assign n163 = pi09 & ~n76;
  assign n164 = ~pi00 & ~n163;
  assign n165 = n96 & ~n162;
  assign n166 = ~n164 & n165;
  assign n167 = ~n114 & ~n160;
  assign n168 = ~n166 & n167;
  assign n169 = ~n158 & n168;
  assign n170 = ~n145 & n169;
  assign n171 = ~n149 & ~n154;
  assign n172 = n170 & n171;
  assign n173 = ~n141 & n172;
  assign n174 = ~pi12 & pi13;
  assign n175 = ~n173 & n174;
  assign n176 = pi12 & n173;
  assign n177 = pi13 & ~n175;
  assign n178 = ~n176 & n177;
  assign n179 = ~n105 & n112;
  assign po0 = n178 | ~n179;
  assign n181 = ~pi05 & n78;
  assign n182 = ~pi01 & ~pi05;
  assign n183 = n45 & ~n182;
  assign n184 = pi01 & pi05;
  assign n185 = ~pi09 & n57;
  assign n186 = pi13 & n185;
  assign n187 = n54 & ~n186;
  assign n188 = ~pi00 & pi04;
  assign n189 = ~pi08 & n188;
  assign n190 = n125 & n189;
  assign n191 = n187 & ~n190;
  assign n192 = n184 & ~n191;
  assign n193 = ~pi05 & ~n67;
  assign n194 = ~pi01 & n38;
  assign n195 = n23 & n109;
  assign n196 = ~n182 & n188;
  assign n197 = ~pi01 & pi05;
  assign n198 = n57 & n197;
  assign n199 = pi01 & ~pi05;
  assign n200 = ~n188 & ~n199;
  assign n201 = ~n198 & n200;
  assign n202 = pi09 & ~n196;
  assign n203 = ~n201 & n202;
  assign n204 = ~n195 & ~n203;
  assign n205 = n119 & ~n204;
  assign n206 = ~n183 & ~n194;
  assign n207 = ~n193 & n206;
  assign n208 = ~n205 & n207;
  assign n209 = ~n192 & n208;
  assign n210 = ~n34 & n209;
  assign n211 = pi05 & n27;
  assign n212 = ~pi01 & ~n211;
  assign n213 = pi11 & ~n184;
  assign n214 = ~n212 & n213;
  assign n215 = ~n181 & ~n214;
  assign n216 = ~n210 & n215;
  assign n217 = ~pi09 & ~n216;
  assign n218 = pi11 & ~n25;
  assign n219 = pi09 & ~n209;
  assign n220 = n63 & n219;
  assign n221 = ~n218 & ~n220;
  assign n222 = pi01 & ~n221;
  assign n223 = pi05 & n96;
  assign n224 = ~n99 & ~n223;
  assign n225 = ~n209 & ~n224;
  assign n226 = n88 & n182;
  assign n227 = ~pi01 & ~n84;
  assign n228 = pi05 & ~n90;
  assign n229 = ~n227 & n228;
  assign n230 = ~n226 & ~n229;
  assign n231 = pi09 & ~n230;
  assign n232 = ~n225 & ~n231;
  assign n233 = ~n217 & n232;
  assign n234 = ~n222 & n233;
  assign n235 = ~pi13 & ~n234;
  assign n236 = pi10 & ~n47;
  assign n237 = ~n24 & ~n236;
  assign n238 = pi11 & ~n237;
  assign n239 = n86 & ~n209;
  assign n240 = ~n86 & n209;
  assign n241 = ~n239 & ~n240;
  assign n242 = n238 & n241;
  assign n243 = ~pi01 & n209;
  assign n244 = n120 & ~n243;
  assign n245 = n24 & n209;
  assign n246 = pi05 & ~pi09;
  assign n247 = ~n219 & ~n246;
  assign n248 = pi01 & pi08;
  assign n249 = ~n247 & n248;
  assign n250 = ~n245 & ~n249;
  assign n251 = n125 & ~n250;
  assign n252 = ~n244 & ~n251;
  assign n253 = pi00 & ~n132;
  assign n254 = n252 & ~n253;
  assign n255 = ~n132 & ~n252;
  assign n256 = pi00 & n255;
  assign n257 = ~n254 & ~n256;
  assign n258 = n53 & n257;
  assign n259 = ~n242 & ~n258;
  assign n260 = ~pi01 & ~n259;
  assign n261 = n132 & n252;
  assign n262 = ~n255 & ~n261;
  assign n263 = n113 & ~n262;
  assign n264 = pi09 & n96;
  assign n265 = ~n209 & n264;
  assign n266 = ~n263 & ~n265;
  assign n267 = ~pi11 & ~n266;
  assign n268 = ~pi05 & ~n55;
  assign n269 = n159 & n268;
  assign n270 = ~n57 & ~n237;
  assign n271 = ~n241 & n270;
  assign n272 = n32 & ~n47;
  assign n273 = n23 & n113;
  assign n274 = ~n269 & ~n272;
  assign n275 = ~n273 & n274;
  assign n276 = ~n271 & n275;
  assign n277 = pi01 & ~n276;
  assign n278 = ~pi11 & n58;
  assign n279 = ~n115 & ~n278;
  assign n280 = ~n76 & ~n279;
  assign n281 = ~n209 & n280;
  assign n282 = n76 & n209;
  assign n283 = ~n117 & n282;
  assign n284 = ~pi00 & ~pi01;
  assign n285 = n113 & n284;
  assign n286 = n55 & n182;
  assign n287 = n159 & n286;
  assign n288 = ~n285 & ~n287;
  assign n289 = pi11 & ~n288;
  assign n290 = ~n55 & ~n197;
  assign n291 = n55 & ~n184;
  assign n292 = n159 & ~n290;
  assign n293 = ~n291 & n292;
  assign n294 = n121 & n184;
  assign n295 = n133 & n252;
  assign n296 = ~n294 & ~n295;
  assign n297 = n122 & ~n132;
  assign n298 = ~n296 & n297;
  assign n299 = n296 & ~n297;
  assign n300 = ~n298 & ~n299;
  assign n301 = n252 & ~n300;
  assign n302 = ~n252 & n300;
  assign n303 = n142 & ~n301;
  assign n304 = ~n302 & n303;
  assign n305 = ~n76 & ~n135;
  assign n306 = ~n296 & n305;
  assign n307 = n296 & ~n305;
  assign n308 = ~n306 & ~n307;
  assign n309 = n209 & ~n308;
  assign n310 = ~n209 & n308;
  assign n311 = n63 & ~n309;
  assign n312 = ~n310 & n311;
  assign n313 = pi01 & ~pi08;
  assign n314 = ~n257 & n313;
  assign n315 = ~n211 & ~n314;
  assign n316 = ~n312 & n315;
  assign n317 = n52 & ~n316;
  assign n318 = ~n289 & ~n293;
  assign n319 = ~n281 & n318;
  assign n320 = ~n283 & n319;
  assign n321 = ~n277 & n320;
  assign n322 = ~n267 & n321;
  assign n323 = ~n260 & n322;
  assign n324 = ~n304 & n323;
  assign n325 = ~n317 & n324;
  assign n326 = ~n175 & n325;
  assign n327 = n175 & ~n325;
  assign n328 = pi13 & ~n326;
  assign n329 = ~n327 & n328;
  assign n330 = n112 & ~n235;
  assign po1 = n329 | ~n330;
  assign n332 = ~pi02 & n38;
  assign n333 = ~n188 & ~n197;
  assign n334 = ~n199 & ~n333;
  assign n335 = pi06 & n334;
  assign n336 = n57 & n335;
  assign n337 = ~pi06 & ~n334;
  assign n338 = pi09 & n337;
  assign n339 = ~n336 & ~n338;
  assign n340 = pi02 & ~n339;
  assign n341 = ~n57 & ~n334;
  assign n342 = ~pi02 & pi09;
  assign n343 = ~n335 & n342;
  assign n344 = ~n337 & ~n341;
  assign n345 = n343 & n344;
  assign n346 = pi01 & pi11;
  assign n347 = n109 & n346;
  assign n348 = ~n345 & ~n347;
  assign n349 = ~n340 & n348;
  assign n350 = n119 & ~n349;
  assign n351 = pi02 & pi06;
  assign n352 = ~n187 & n351;
  assign n353 = ~pi02 & ~pi06;
  assign n354 = n45 & ~n353;
  assign n355 = ~pi06 & ~n67;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n352 & n356;
  assign n358 = ~n350 & n357;
  assign n359 = ~n332 & n358;
  assign n360 = ~n34 & n359;
  assign n361 = ~pi06 & n78;
  assign n362 = ~n360 & ~n361;
  assign n363 = ~pi09 & ~n362;
  assign n364 = pi09 & n84;
  assign n365 = ~pi02 & n27;
  assign n366 = n62 & n365;
  assign n367 = ~n364 & ~n366;
  assign n368 = pi06 & ~n367;
  assign n369 = ~n90 & n351;
  assign n370 = n88 & n353;
  assign n371 = ~n369 & ~n370;
  assign n372 = pi09 & ~n371;
  assign n373 = pi02 & pi11;
  assign n374 = ~pi06 & ~pi09;
  assign n375 = n25 & ~n374;
  assign n376 = n373 & ~n375;
  assign n377 = pi06 & n96;
  assign n378 = pi02 & n113;
  assign n379 = ~n99 & ~n377;
  assign n380 = ~n378 & n379;
  assign n381 = ~n359 & ~n380;
  assign n382 = ~n368 & ~n376;
  assign n383 = ~n372 & n382;
  assign n384 = ~n381 & n383;
  assign n385 = ~n363 & n384;
  assign n386 = ~pi13 & ~n385;
  assign n387 = pi06 & n27;
  assign n388 = n121 & n351;
  assign n389 = ~pi02 & n359;
  assign n390 = n120 & ~n389;
  assign n391 = n24 & n359;
  assign n392 = pi09 & n359;
  assign n393 = pi02 & pi08;
  assign n394 = ~n374 & n393;
  assign n395 = ~n392 & n394;
  assign n396 = ~n391 & ~n395;
  assign n397 = n125 & ~n396;
  assign n398 = ~n390 & ~n397;
  assign n399 = n133 & n398;
  assign n400 = ~n388 & ~n399;
  assign n401 = n359 & n400;
  assign n402 = ~n359 & ~n400;
  assign n403 = ~n401 & ~n402;
  assign n404 = ~n209 & ~n307;
  assign n405 = ~n306 & ~n404;
  assign n406 = ~n403 & n405;
  assign n407 = n403 & ~n405;
  assign n408 = n63 & ~n406;
  assign n409 = ~n407 & n408;
  assign n410 = pi01 & ~n254;
  assign n411 = ~n256 & ~n410;
  assign n412 = ~n398 & n411;
  assign n413 = n398 & ~n411;
  assign n414 = ~n412 & ~n413;
  assign n415 = pi02 & ~pi08;
  assign n416 = n414 & n415;
  assign n417 = ~n387 & ~n416;
  assign n418 = ~n409 & n417;
  assign n419 = n52 & ~n418;
  assign n420 = n53 & ~n414;
  assign n421 = pi01 & ~n240;
  assign n422 = ~n239 & ~n421;
  assign n423 = n238 & ~n359;
  assign n424 = n422 & n423;
  assign n425 = ~n420 & ~n424;
  assign n426 = ~pi02 & ~n425;
  assign n427 = ~pi02 & n284;
  assign n428 = pi11 & n427;
  assign n429 = ~n284 & n373;
  assign n430 = n261 & n398;
  assign n431 = ~n261 & ~n398;
  assign n432 = ~n430 & ~n431;
  assign n433 = ~pi11 & ~n432;
  assign n434 = ~n428 & ~n429;
  assign n435 = ~n433 & n434;
  assign n436 = n113 & ~n435;
  assign n437 = n270 & ~n359;
  assign n438 = ~n422 & n437;
  assign n439 = ~n272 & ~n438;
  assign n440 = pi02 & ~n439;
  assign n441 = ~n55 & ~n184;
  assign n442 = ~n182 & ~n441;
  assign n443 = ~n351 & ~n353;
  assign n444 = ~n442 & ~n443;
  assign n445 = pi11 & n353;
  assign n446 = ~n351 & ~n445;
  assign n447 = n442 & n446;
  assign n448 = n159 & ~n444;
  assign n449 = ~n447 & n448;
  assign n450 = n283 & n359;
  assign n451 = ~pi10 & n278;
  assign n452 = n282 & ~n451;
  assign n453 = ~n279 & ~n359;
  assign n454 = ~n452 & n453;
  assign n455 = ~pi02 & n422;
  assign n456 = n270 & n422;
  assign n457 = ~pi02 & n238;
  assign n458 = ~n456 & ~n457;
  assign n459 = n359 & ~n455;
  assign n460 = ~n458 & n459;
  assign n461 = ~n252 & ~n299;
  assign n462 = ~n298 & ~n461;
  assign n463 = n400 & n462;
  assign n464 = ~n400 & ~n462;
  assign n465 = ~n463 & ~n464;
  assign n466 = n398 & ~n465;
  assign n467 = ~n398 & n465;
  assign n468 = n142 & ~n466;
  assign n469 = ~n467 & n468;
  assign n470 = ~n449 & ~n450;
  assign n471 = ~n454 & n470;
  assign n472 = ~n440 & n471;
  assign n473 = ~n460 & n472;
  assign n474 = ~n436 & n473;
  assign n475 = ~n426 & n474;
  assign n476 = ~n419 & n475;
  assign n477 = ~n469 & n476;
  assign n478 = pi13 & n327;
  assign n479 = ~n477 & n478;
  assign n480 = ~n327 & n477;
  assign n481 = pi13 & ~n479;
  assign n482 = ~n480 & n481;
  assign n483 = n112 & ~n386;
  assign po2 = n482 | ~n483;
  assign n485 = ~pi03 & ~pi07;
  assign n486 = n88 & n485;
  assign po5 = pi03 & pi07;
  assign n488 = ~n90 & po5;
  assign n489 = n45 & ~n485;
  assign n490 = pi02 & ~n335;
  assign n491 = ~n337 & ~n490;
  assign n492 = pi07 & pi09;
  assign n493 = n125 & n492;
  assign n494 = ~n491 & n493;
  assign n495 = ~n37 & ~n494;
  assign n496 = ~pi03 & ~n495;
  assign n497 = n109 & n373;
  assign n498 = pi09 & n485;
  assign n499 = n491 & n498;
  assign n500 = ~n497 & ~n499;
  assign n501 = pi13 & ~n500;
  assign n502 = n125 & n491;
  assign n503 = ~n185 & ~n502;
  assign n504 = po5 & ~n503;
  assign n505 = ~n496 & ~n501;
  assign n506 = ~n504 & n505;
  assign n507 = ~pi08 & ~n506;
  assign n508 = pi03 & n59;
  assign n509 = ~n491 & n508;
  assign n510 = n67 & ~n509;
  assign n511 = ~pi07 & ~n510;
  assign n512 = ~n50 & ~n185;
  assign n513 = pi13 & po5;
  assign n514 = ~n512 & n513;
  assign n515 = ~n489 & ~n514;
  assign n516 = ~n511 & n515;
  assign n517 = ~n507 & n516;
  assign n518 = pi03 & ~n517;
  assign n519 = n63 & n518;
  assign n520 = ~n486 & ~n488;
  assign n521 = ~n519 & n520;
  assign n522 = pi09 & ~n521;
  assign n523 = ~n34 & n517;
  assign n524 = ~pi07 & n78;
  assign n525 = ~n523 & ~n524;
  assign n526 = ~pi09 & ~n525;
  assign n527 = pi07 & n96;
  assign n528 = ~n99 & ~n527;
  assign n529 = ~n517 & ~n528;
  assign n530 = pi03 & pi11;
  assign n531 = ~pi07 & ~pi09;
  assign n532 = n25 & ~n531;
  assign n533 = n530 & ~n532;
  assign n534 = ~pi03 & n27;
  assign n535 = n62 & n534;
  assign n536 = ~n364 & ~n535;
  assign n537 = pi07 & ~n536;
  assign n538 = ~n533 & ~n537;
  assign n539 = ~n529 & n538;
  assign n540 = ~n526 & n539;
  assign n541 = ~n522 & n540;
  assign n542 = ~pi13 & ~n541;
  assign n543 = n121 & po5;
  assign n544 = ~pi03 & n517;
  assign n545 = n120 & ~n544;
  assign n546 = n24 & n517;
  assign n547 = n42 & po5;
  assign n548 = n47 & n518;
  assign n549 = ~n546 & ~n547;
  assign n550 = ~n548 & n549;
  assign n551 = n125 & ~n550;
  assign n552 = ~n545 & ~n551;
  assign n553 = n133 & n552;
  assign n554 = ~n543 & ~n553;
  assign n555 = ~n401 & ~n405;
  assign n556 = ~n402 & ~n555;
  assign n557 = n517 & n556;
  assign n558 = ~n517 & ~n556;
  assign n559 = ~n557 & ~n558;
  assign n560 = n554 & ~n559;
  assign n561 = ~n554 & n559;
  assign n562 = pi08 & ~n560;
  assign n563 = ~n561 & n562;
  assign n564 = ~pi02 & n398;
  assign n565 = ~n411 & ~n564;
  assign n566 = pi02 & ~n398;
  assign n567 = ~n565 & ~n566;
  assign n568 = ~n552 & ~n567;
  assign n569 = ~pi03 & ~n568;
  assign n570 = n552 & n567;
  assign n571 = ~pi08 & ~n570;
  assign n572 = n569 & n571;
  assign n573 = ~n563 & ~n572;
  assign n574 = n185 & ~n573;
  assign n575 = pi02 & ~n358;
  assign n576 = n422 & ~n575;
  assign n577 = ~n389 & ~n576;
  assign n578 = ~n517 & ~n577;
  assign n579 = n517 & n577;
  assign n580 = ~n578 & ~n579;
  assign n581 = n238 & ~n580;
  assign n582 = pi07 & n159;
  assign n583 = ~n351 & ~n442;
  assign n584 = ~n353 & ~n583;
  assign n585 = n582 & ~n584;
  assign n586 = ~n581 & ~n585;
  assign n587 = ~pi03 & ~n586;
  assign n588 = n270 & n580;
  assign n589 = ~n272 & ~n588;
  assign n590 = pi03 & ~n589;
  assign n591 = n282 & n359;
  assign n592 = ~n451 & n591;
  assign n593 = ~n279 & ~n517;
  assign n594 = ~n592 & n593;
  assign n595 = n450 & n517;
  assign n596 = n113 & n530;
  assign n597 = ~n427 & n596;
  assign n598 = ~pi07 & n584;
  assign n599 = pi07 & ~n584;
  assign n600 = pi03 & n159;
  assign n601 = ~n598 & n600;
  assign n602 = ~n599 & n601;
  assign n603 = n430 & n552;
  assign n604 = ~n430 & ~n552;
  assign n605 = ~n603 & ~n604;
  assign n606 = n113 & ~n605;
  assign n607 = ~n568 & ~n570;
  assign n608 = pi03 & n24;
  assign n609 = ~n607 & n608;
  assign n610 = ~n582 & ~n606;
  assign n611 = ~n609 & n610;
  assign n612 = ~pi11 & ~n611;
  assign n613 = ~n398 & ~n463;
  assign n614 = ~n464 & ~n613;
  assign n615 = n554 & n614;
  assign n616 = ~n554 & ~n614;
  assign n617 = ~n615 & ~n616;
  assign n618 = n552 & ~n617;
  assign n619 = ~n552 & n617;
  assign n620 = n264 & ~n618;
  assign n621 = ~n619 & n620;
  assign n622 = ~pi03 & n113;
  assign n623 = n427 & n622;
  assign n624 = ~pi03 & n159;
  assign n625 = n598 & n624;
  assign n626 = ~n623 & ~n625;
  assign n627 = ~n621 & n626;
  assign n628 = pi11 & ~n627;
  assign n629 = ~n597 & ~n602;
  assign n630 = ~n595 & n629;
  assign n631 = ~n594 & n630;
  assign n632 = ~n587 & n631;
  assign n633 = ~n590 & n632;
  assign n634 = ~n612 & n633;
  assign n635 = ~n574 & n634;
  assign n636 = ~n628 & n635;
  assign n637 = ~n479 & n636;
  assign n638 = n479 & ~n636;
  assign n639 = pi13 & ~n637;
  assign n640 = ~n638 & n639;
  assign n641 = n112 & ~n542;
  assign po3 = n640 | ~n641;
  assign po4 = n485 | po5;
  assign n644 = ~po5 & ~n584;
  assign n645 = n159 & ~n485;
  assign n646 = ~n644 & n645;
  assign n647 = ~n518 & ~n577;
  assign n648 = ~n237 & ~n544;
  assign n649 = ~n647 & n648;
  assign n650 = n552 & ~n616;
  assign n651 = n264 & ~n615;
  assign n652 = ~n650 & n651;
  assign n653 = ~n623 & ~n646;
  assign n654 = ~n649 & n653;
  assign n655 = ~n652 & n654;
  assign n656 = pi11 & ~n655;
  assign n657 = ~n106 & ~n116;
  assign n658 = n591 & ~n657;
  assign n659 = n517 & n658;
  assign n660 = ~n569 & n571;
  assign n661 = n554 & ~n558;
  assign n662 = pi08 & ~n557;
  assign n663 = ~n661 & n662;
  assign n664 = ~n660 & ~n663;
  assign n665 = n109 & ~n664;
  assign n666 = pi10 & ~n603;
  assign n667 = n47 & ~n666;
  assign n668 = ~n665 & ~n667;
  assign n669 = ~pi11 & ~n668;
  assign n670 = ~n656 & ~n659;
  assign n671 = ~n669 & n670;
  assign n672 = ~n638 & n671;
  assign po6 = pi13 & ~n672;
  assign n674 = ~n182 & ~n184;
  assign n675 = ~n69 & ~n443;
  assign n676 = po4 & ~n674;
  assign po7 = n675 & n676;
endmodule
