module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7;
  wire n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500,
    n501, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n860,
    n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909,
    n910, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931,
    n933, n934, n935, n936, n937, n940, n941,
    n942, n943, n944, n945;
  assign n137 = pi124  & ~pi125 ;
  assign n138 = ~pi126  & ~n137;
  assign n139 = ~pi127  & ~n138;
  assign n140 = ~pi122  & ~n139;
  assign n141 = ~pi123  & pi125 ;
  assign n142 = ~pi126  & n141;
  assign n143 = pi123  & n138;
  assign n144 = ~pi127  & ~n142;
  assign n145 = ~n143 & n144;
  assign n146 = pi122  & ~n145;
  assign n147 = ~n140 & ~n146;
  assign n148 = ~pi120  & ~n147;
  assign n149 = ~pi121  & ~n145;
  assign n150 = pi121  & ~n147;
  assign n151 = ~n149 & ~n150;
  assign n152 = pi120  & ~n151;
  assign n153 = ~n148 & ~n152;
  assign n154 = ~pi118  & ~n153;
  assign n155 = ~pi119  & ~n151;
  assign n156 = pi119  & ~n153;
  assign n157 = ~n155 & ~n156;
  assign n158 = pi118  & ~n157;
  assign n159 = ~n154 & ~n158;
  assign n160 = ~pi116  & ~n159;
  assign n161 = ~pi117  & ~n157;
  assign n162 = pi117  & ~n159;
  assign n163 = ~n161 & ~n162;
  assign n164 = pi116  & ~n163;
  assign n165 = ~n160 & ~n164;
  assign n166 = ~pi114  & ~n165;
  assign n167 = ~pi115  & ~n163;
  assign n168 = pi115  & ~n165;
  assign n169 = ~n167 & ~n168;
  assign n170 = pi114  & ~n169;
  assign n171 = ~n166 & ~n170;
  assign n172 = ~pi112  & ~n171;
  assign n173 = ~pi113  & ~n169;
  assign n174 = pi113  & ~n171;
  assign n175 = ~n173 & ~n174;
  assign n176 = pi112  & ~n175;
  assign n177 = ~n172 & ~n176;
  assign n178 = ~pi110  & ~n177;
  assign n179 = ~pi111  & ~n175;
  assign n180 = pi111  & ~n177;
  assign n181 = ~n179 & ~n180;
  assign n182 = pi110  & ~n181;
  assign n183 = ~n178 & ~n182;
  assign n184 = ~pi108  & ~n183;
  assign n185 = ~pi109  & ~n181;
  assign n186 = pi109  & ~n183;
  assign n187 = ~n185 & ~n186;
  assign n188 = pi108  & ~n187;
  assign n189 = ~n184 & ~n188;
  assign n190 = ~pi106  & ~n189;
  assign n191 = ~pi107  & ~n187;
  assign n192 = pi107  & ~n189;
  assign n193 = ~n191 & ~n192;
  assign n194 = pi106  & ~n193;
  assign n195 = ~n190 & ~n194;
  assign n196 = ~pi104  & ~n195;
  assign n197 = ~pi105  & ~n193;
  assign n198 = pi105  & ~n195;
  assign n199 = ~n197 & ~n198;
  assign n200 = pi104  & ~n199;
  assign n201 = ~n196 & ~n200;
  assign n202 = ~pi102  & ~n201;
  assign n203 = ~pi103  & ~n199;
  assign n204 = pi103  & ~n201;
  assign n205 = ~n203 & ~n204;
  assign n206 = pi102  & ~n205;
  assign n207 = ~n202 & ~n206;
  assign n208 = ~pi100  & ~n207;
  assign n209 = ~pi101  & ~n205;
  assign n210 = pi101  & ~n207;
  assign n211 = ~n209 & ~n210;
  assign n212 = pi100  & ~n211;
  assign n213 = ~n208 & ~n212;
  assign n214 = ~pi98  & ~n213;
  assign n215 = ~pi99  & ~n211;
  assign n216 = pi99  & ~n213;
  assign n217 = ~n215 & ~n216;
  assign n218 = pi98  & ~n217;
  assign n219 = ~n214 & ~n218;
  assign n220 = ~pi96  & ~n219;
  assign n221 = ~pi97  & ~n217;
  assign n222 = pi97  & ~n219;
  assign n223 = ~n221 & ~n222;
  assign n224 = pi96  & ~n223;
  assign n225 = ~n220 & ~n224;
  assign n226 = ~pi94  & ~n225;
  assign n227 = ~pi95  & ~n223;
  assign n228 = pi95  & ~n225;
  assign n229 = ~n227 & ~n228;
  assign n230 = pi94  & ~n229;
  assign n231 = ~n226 & ~n230;
  assign n232 = ~pi92  & ~n231;
  assign n233 = ~pi93  & ~n229;
  assign n234 = pi93  & ~n231;
  assign n235 = ~n233 & ~n234;
  assign n236 = pi92  & ~n235;
  assign n237 = ~n232 & ~n236;
  assign n238 = ~pi90  & ~n237;
  assign n239 = ~pi91  & ~n235;
  assign n240 = pi91  & ~n237;
  assign n241 = ~n239 & ~n240;
  assign n242 = pi90  & ~n241;
  assign n243 = ~n238 & ~n242;
  assign n244 = ~pi88  & ~n243;
  assign n245 = ~pi89  & ~n241;
  assign n246 = pi89  & ~n243;
  assign n247 = ~n245 & ~n246;
  assign n248 = pi88  & ~n247;
  assign n249 = ~n244 & ~n248;
  assign n250 = ~pi86  & ~n249;
  assign n251 = ~pi87  & ~n247;
  assign n252 = pi87  & ~n249;
  assign n253 = ~n251 & ~n252;
  assign n254 = pi86  & ~n253;
  assign n255 = ~n250 & ~n254;
  assign n256 = ~pi84  & ~n255;
  assign n257 = ~pi85  & ~n253;
  assign n258 = pi85  & ~n255;
  assign n259 = ~n257 & ~n258;
  assign n260 = pi84  & ~n259;
  assign n261 = ~n256 & ~n260;
  assign n262 = ~pi82  & ~n261;
  assign n263 = ~pi83  & ~n259;
  assign n264 = pi83  & ~n261;
  assign n265 = ~n263 & ~n264;
  assign n266 = pi82  & ~n265;
  assign n267 = ~n262 & ~n266;
  assign n268 = ~pi80  & ~n267;
  assign n269 = ~pi81  & ~n265;
  assign n270 = pi81  & ~n267;
  assign n271 = ~n269 & ~n270;
  assign n272 = pi80  & ~n271;
  assign n273 = ~n268 & ~n272;
  assign n274 = ~pi78  & ~n273;
  assign n275 = ~pi79  & ~n271;
  assign n276 = pi79  & ~n273;
  assign n277 = ~n275 & ~n276;
  assign n278 = pi78  & ~n277;
  assign n279 = ~n274 & ~n278;
  assign n280 = ~pi76  & ~n279;
  assign n281 = ~pi77  & ~n277;
  assign n282 = pi77  & ~n279;
  assign n283 = ~n281 & ~n282;
  assign n284 = pi76  & ~n283;
  assign n285 = ~n280 & ~n284;
  assign n286 = ~pi74  & ~n285;
  assign n287 = ~pi75  & ~n283;
  assign n288 = pi75  & ~n285;
  assign n289 = ~n287 & ~n288;
  assign n290 = pi74  & ~n289;
  assign n291 = ~n286 & ~n290;
  assign n292 = ~pi72  & ~n291;
  assign n293 = ~pi73  & ~n289;
  assign n294 = pi73  & ~n291;
  assign n295 = ~n293 & ~n294;
  assign n296 = pi72  & ~n295;
  assign n297 = ~n292 & ~n296;
  assign n298 = ~pi70  & ~n297;
  assign n299 = ~pi71  & ~n295;
  assign n300 = pi71  & ~n297;
  assign n301 = ~n299 & ~n300;
  assign n302 = pi70  & ~n301;
  assign n303 = ~n298 & ~n302;
  assign n304 = ~pi68  & ~n303;
  assign n305 = ~pi69  & ~n301;
  assign n306 = pi69  & ~n303;
  assign n307 = ~n305 & ~n306;
  assign n308 = pi68  & ~n307;
  assign n309 = ~n304 & ~n308;
  assign n310 = ~pi66  & ~n309;
  assign n311 = ~pi67  & ~n307;
  assign n312 = pi67  & ~n309;
  assign n313 = ~n311 & ~n312;
  assign n314 = pi66  & ~n313;
  assign n315 = ~n310 & ~n314;
  assign n316 = ~pi64  & ~n315;
  assign n317 = ~pi65  & ~n313;
  assign n318 = pi65  & ~n315;
  assign n319 = ~n317 & ~n318;
  assign n320 = pi64  & ~n319;
  assign n321 = ~n316 & ~n320;
  assign n322 = ~pi62  & ~n321;
  assign n323 = ~pi63  & ~n319;
  assign n324 = pi63  & ~n321;
  assign n325 = ~n323 & ~n324;
  assign n326 = pi62  & ~n325;
  assign n327 = ~n322 & ~n326;
  assign n328 = ~pi60  & ~n327;
  assign n329 = ~pi61  & ~n325;
  assign n330 = pi61  & ~n327;
  assign n331 = ~n329 & ~n330;
  assign n332 = pi60  & ~n331;
  assign n333 = ~n328 & ~n332;
  assign n334 = ~pi58  & ~n333;
  assign n335 = ~pi59  & ~n331;
  assign n336 = pi59  & ~n333;
  assign n337 = ~n335 & ~n336;
  assign n338 = pi58  & ~n337;
  assign n339 = ~n334 & ~n338;
  assign n340 = ~pi56  & ~n339;
  assign n341 = ~pi57  & ~n337;
  assign n342 = pi57  & ~n339;
  assign n343 = ~n341 & ~n342;
  assign n344 = pi56  & ~n343;
  assign n345 = ~n340 & ~n344;
  assign n346 = ~pi54  & ~n345;
  assign n347 = ~pi55  & ~n343;
  assign n348 = pi55  & ~n345;
  assign n349 = ~n347 & ~n348;
  assign n350 = pi54  & ~n349;
  assign n351 = ~n346 & ~n350;
  assign n352 = ~pi52  & ~n351;
  assign n353 = ~pi53  & ~n349;
  assign n354 = pi53  & ~n351;
  assign n355 = ~n353 & ~n354;
  assign n356 = pi52  & ~n355;
  assign n357 = ~n352 & ~n356;
  assign n358 = ~pi50  & ~n357;
  assign n359 = ~pi51  & ~n355;
  assign n360 = pi51  & ~n357;
  assign n361 = ~n359 & ~n360;
  assign n362 = pi50  & ~n361;
  assign n363 = ~n358 & ~n362;
  assign n364 = ~pi48  & ~n363;
  assign n365 = ~pi49  & ~n361;
  assign n366 = pi49  & ~n363;
  assign n367 = ~n365 & ~n366;
  assign n368 = pi48  & ~n367;
  assign n369 = ~n364 & ~n368;
  assign n370 = ~pi46  & ~n369;
  assign n371 = ~pi47  & ~n367;
  assign n372 = pi47  & ~n369;
  assign n373 = ~n371 & ~n372;
  assign n374 = pi46  & ~n373;
  assign n375 = ~n370 & ~n374;
  assign n376 = ~pi44  & ~n375;
  assign n377 = ~pi45  & ~n373;
  assign n378 = pi45  & ~n375;
  assign n379 = ~n377 & ~n378;
  assign n380 = pi44  & ~n379;
  assign n381 = ~n376 & ~n380;
  assign n382 = ~pi42  & ~n381;
  assign n383 = ~pi43  & ~n379;
  assign n384 = pi43  & ~n381;
  assign n385 = ~n383 & ~n384;
  assign n386 = pi42  & ~n385;
  assign n387 = ~n382 & ~n386;
  assign n388 = ~pi40  & ~n387;
  assign n389 = ~pi41  & ~n385;
  assign n390 = pi41  & ~n387;
  assign n391 = ~n389 & ~n390;
  assign n392 = pi40  & ~n391;
  assign n393 = ~n388 & ~n392;
  assign n394 = ~pi38  & ~n393;
  assign n395 = ~pi39  & ~n391;
  assign n396 = pi39  & ~n393;
  assign n397 = ~n395 & ~n396;
  assign n398 = pi38  & ~n397;
  assign n399 = ~n394 & ~n398;
  assign n400 = ~pi36  & ~n399;
  assign n401 = ~pi37  & ~n397;
  assign n402 = pi37  & ~n399;
  assign n403 = ~n401 & ~n402;
  assign n404 = pi36  & ~n403;
  assign n405 = ~n400 & ~n404;
  assign n406 = ~pi34  & ~n405;
  assign n407 = ~pi35  & ~n403;
  assign n408 = pi35  & ~n405;
  assign n409 = ~n407 & ~n408;
  assign n410 = pi34  & ~n409;
  assign n411 = ~n406 & ~n410;
  assign n412 = ~pi32  & ~n411;
  assign n413 = ~pi33  & ~n409;
  assign n414 = pi33  & ~n411;
  assign n415 = ~n413 & ~n414;
  assign n416 = pi32  & ~n415;
  assign n417 = ~n412 & ~n416;
  assign n418 = ~pi30  & ~n417;
  assign n419 = ~pi31  & ~n415;
  assign n420 = pi31  & ~n417;
  assign n421 = ~n419 & ~n420;
  assign n422 = pi30  & ~n421;
  assign n423 = ~n418 & ~n422;
  assign n424 = ~pi28  & ~n423;
  assign n425 = ~pi29  & ~n421;
  assign n426 = pi29  & ~n423;
  assign n427 = ~n425 & ~n426;
  assign n428 = pi28  & ~n427;
  assign n429 = ~n424 & ~n428;
  assign n430 = ~pi26  & ~n429;
  assign n431 = ~pi27  & ~n427;
  assign n432 = pi27  & ~n429;
  assign n433 = ~n431 & ~n432;
  assign n434 = pi26  & ~n433;
  assign n435 = ~n430 & ~n434;
  assign n436 = ~pi24  & ~n435;
  assign n437 = ~pi25  & ~n433;
  assign n438 = pi25  & ~n435;
  assign n439 = ~n437 & ~n438;
  assign n440 = pi24  & ~n439;
  assign n441 = ~n436 & ~n440;
  assign n442 = ~pi22  & ~n441;
  assign n443 = ~pi23  & ~n439;
  assign n444 = pi23  & ~n441;
  assign n445 = ~n443 & ~n444;
  assign n446 = pi22  & ~n445;
  assign n447 = ~n442 & ~n446;
  assign n448 = ~pi20  & ~n447;
  assign n449 = ~pi21  & ~n445;
  assign n450 = pi21  & ~n447;
  assign n451 = ~n449 & ~n450;
  assign n452 = pi20  & ~n451;
  assign n453 = ~n448 & ~n452;
  assign n454 = ~pi18  & ~n453;
  assign n455 = ~pi19  & ~n451;
  assign n456 = pi19  & ~n453;
  assign n457 = ~n455 & ~n456;
  assign n458 = pi18  & ~n457;
  assign n459 = ~n454 & ~n458;
  assign n460 = ~pi16  & ~n459;
  assign n461 = ~pi17  & ~n457;
  assign n462 = pi17  & ~n459;
  assign n463 = ~n461 & ~n462;
  assign n464 = pi16  & ~n463;
  assign n465 = ~n460 & ~n464;
  assign n466 = ~pi14  & ~n465;
  assign n467 = ~pi15  & ~n463;
  assign n468 = pi15  & ~n465;
  assign n469 = ~n467 & ~n468;
  assign n470 = pi14  & ~n469;
  assign n471 = ~n466 & ~n470;
  assign n472 = ~pi12  & ~n471;
  assign n473 = ~pi13  & ~n469;
  assign n474 = pi13  & ~n471;
  assign n475 = ~n473 & ~n474;
  assign n476 = pi12  & ~n475;
  assign n477 = ~n472 & ~n476;
  assign n478 = ~pi10  & ~n477;
  assign n479 = ~pi11  & ~n475;
  assign n480 = pi11  & ~n477;
  assign n481 = ~n479 & ~n480;
  assign n482 = pi10  & ~n481;
  assign n483 = ~n478 & ~n482;
  assign n484 = ~pi8  & ~n483;
  assign n485 = ~pi9  & ~n481;
  assign n486 = pi9  & ~n483;
  assign n487 = ~n485 & ~n486;
  assign n488 = pi8  & ~n487;
  assign n489 = ~n484 & ~n488;
  assign n490 = ~pi6  & ~n489;
  assign n491 = ~pi7  & ~n487;
  assign n492 = pi7  & ~n489;
  assign n493 = ~n491 & ~n492;
  assign n494 = pi6  & ~n493;
  assign n495 = pi1  & ~pi2 ;
  assign n496 = ~pi3  & ~n495;
  assign n497 = ~pi4  & ~n496;
  assign n498 = ~pi5  & ~n497;
  assign n499 = ~n490 & ~n498;
  assign n500 = ~n494 & n499;
  assign n501 = n493 & n498;
  assign po0  = ~n500 & ~n501;
  assign n503 = ~pi10  & ~pi11 ;
  assign n504 = ~pi14  & ~pi15 ;
  assign n505 = ~pi18  & ~pi19 ;
  assign n506 = ~pi22  & ~pi23 ;
  assign n507 = ~pi26  & ~pi27 ;
  assign n508 = ~pi30  & ~pi31 ;
  assign n509 = ~pi34  & ~pi35 ;
  assign n510 = ~pi38  & ~pi39 ;
  assign n511 = ~pi42  & ~pi43 ;
  assign n512 = ~pi46  & ~pi47 ;
  assign n513 = ~pi50  & ~pi51 ;
  assign n514 = ~pi54  & ~pi55 ;
  assign n515 = ~pi58  & ~pi59 ;
  assign n516 = ~pi62  & ~pi63 ;
  assign n517 = ~pi66  & ~pi67 ;
  assign n518 = ~pi70  & ~pi71 ;
  assign n519 = ~pi74  & ~pi75 ;
  assign n520 = ~pi78  & ~pi79 ;
  assign n521 = ~pi82  & ~pi83 ;
  assign n522 = ~pi86  & ~pi87 ;
  assign n523 = ~pi90  & ~pi91 ;
  assign n524 = ~pi94  & ~pi95 ;
  assign n525 = ~pi98  & ~pi99 ;
  assign n526 = ~pi102  & ~pi103 ;
  assign n527 = ~pi106  & ~pi107 ;
  assign n528 = ~pi110  & ~pi111 ;
  assign n529 = ~pi114  & ~pi115 ;
  assign n530 = ~pi116  & ~pi117 ;
  assign n531 = ~pi122  & ~pi123 ;
  assign n532 = pi121  & n531;
  assign n533 = ~pi124  & ~pi125 ;
  assign n534 = ~pi120  & n533;
  assign n535 = ~n532 & n534;
  assign n536 = ~pi126  & pi127 ;
  assign n537 = ~pi126  & ~n536;
  assign n538 = ~n531 & n533;
  assign n539 = pi120  & n538;
  assign n540 = ~n535 & n537;
  assign n541 = ~n539 & n540;
  assign n542 = n530 & ~n541;
  assign n543 = ~pi118  & ~pi119 ;
  assign n544 = n541 & ~n543;
  assign n545 = n537 & n543;
  assign n546 = ~n538 & n545;
  assign n547 = ~n544 & ~n546;
  assign n548 = ~n530 & n547;
  assign n549 = ~n542 & ~n548;
  assign n550 = ~n529 & ~n549;
  assign n551 = n529 & n547;
  assign n552 = ~n550 & ~n551;
  assign n553 = n528 & ~n552;
  assign n554 = ~pi112  & ~pi113 ;
  assign n555 = ~n552 & ~n554;
  assign n556 = ~n549 & n554;
  assign n557 = ~n555 & ~n556;
  assign n558 = ~n528 & ~n557;
  assign n559 = ~n553 & ~n558;
  assign n560 = n527 & ~n559;
  assign n561 = ~pi108  & ~pi109 ;
  assign n562 = ~n559 & ~n561;
  assign n563 = ~n557 & n561;
  assign n564 = ~n562 & ~n563;
  assign n565 = ~n527 & ~n564;
  assign n566 = ~n560 & ~n565;
  assign n567 = n526 & ~n566;
  assign n568 = ~pi104  & ~pi105 ;
  assign n569 = ~n566 & ~n568;
  assign n570 = ~n564 & n568;
  assign n571 = ~n569 & ~n570;
  assign n572 = ~n526 & ~n571;
  assign n573 = ~n567 & ~n572;
  assign n574 = n525 & ~n573;
  assign n575 = ~pi100  & ~pi101 ;
  assign n576 = ~n573 & ~n575;
  assign n577 = ~n571 & n575;
  assign n578 = ~n576 & ~n577;
  assign n579 = ~n525 & ~n578;
  assign n580 = ~n574 & ~n579;
  assign n581 = n524 & ~n580;
  assign n582 = ~pi96  & ~pi97 ;
  assign n583 = ~n580 & ~n582;
  assign n584 = ~n578 & n582;
  assign n585 = ~n583 & ~n584;
  assign n586 = ~n524 & ~n585;
  assign n587 = ~n581 & ~n586;
  assign n588 = n523 & ~n587;
  assign n589 = ~pi92  & ~pi93 ;
  assign n590 = ~n587 & ~n589;
  assign n591 = ~n585 & n589;
  assign n592 = ~n590 & ~n591;
  assign n593 = ~n523 & ~n592;
  assign n594 = ~n588 & ~n593;
  assign n595 = n522 & ~n594;
  assign n596 = ~pi88  & ~pi89 ;
  assign n597 = ~n594 & ~n596;
  assign n598 = ~n592 & n596;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~n522 & ~n599;
  assign n601 = ~n595 & ~n600;
  assign n602 = n521 & ~n601;
  assign n603 = ~pi84  & ~pi85 ;
  assign n604 = ~n601 & ~n603;
  assign n605 = ~n599 & n603;
  assign n606 = ~n604 & ~n605;
  assign n607 = ~n521 & ~n606;
  assign n608 = ~n602 & ~n607;
  assign n609 = n520 & ~n608;
  assign n610 = ~pi80  & ~pi81 ;
  assign n611 = ~n608 & ~n610;
  assign n612 = ~n606 & n610;
  assign n613 = ~n611 & ~n612;
  assign n614 = ~n520 & ~n613;
  assign n615 = ~n609 & ~n614;
  assign n616 = n519 & ~n615;
  assign n617 = ~pi76  & ~pi77 ;
  assign n618 = ~n615 & ~n617;
  assign n619 = ~n613 & n617;
  assign n620 = ~n618 & ~n619;
  assign n621 = ~n519 & ~n620;
  assign n622 = ~n616 & ~n621;
  assign n623 = n518 & ~n622;
  assign n624 = ~pi72  & ~pi73 ;
  assign n625 = ~n622 & ~n624;
  assign n626 = ~n620 & n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = ~n518 & ~n627;
  assign n629 = ~n623 & ~n628;
  assign n630 = n517 & ~n629;
  assign n631 = ~pi68  & ~pi69 ;
  assign n632 = ~n629 & ~n631;
  assign n633 = ~n627 & n631;
  assign n634 = ~n632 & ~n633;
  assign n635 = ~n517 & ~n634;
  assign n636 = ~n630 & ~n635;
  assign n637 = n516 & ~n636;
  assign n638 = ~pi64  & ~pi65 ;
  assign n639 = ~n636 & ~n638;
  assign n640 = ~n634 & n638;
  assign n641 = ~n639 & ~n640;
  assign n642 = ~n516 & ~n641;
  assign n643 = ~n637 & ~n642;
  assign n644 = n515 & ~n643;
  assign n645 = ~pi60  & ~pi61 ;
  assign n646 = ~n643 & ~n645;
  assign n647 = ~n641 & n645;
  assign n648 = ~n646 & ~n647;
  assign n649 = ~n515 & ~n648;
  assign n650 = ~n644 & ~n649;
  assign n651 = n514 & ~n650;
  assign n652 = ~pi56  & ~pi57 ;
  assign n653 = ~n650 & ~n652;
  assign n654 = ~n648 & n652;
  assign n655 = ~n653 & ~n654;
  assign n656 = ~n514 & ~n655;
  assign n657 = ~n651 & ~n656;
  assign n658 = n513 & ~n657;
  assign n659 = ~pi52  & ~pi53 ;
  assign n660 = ~n657 & ~n659;
  assign n661 = ~n655 & n659;
  assign n662 = ~n660 & ~n661;
  assign n663 = ~n513 & ~n662;
  assign n664 = ~n658 & ~n663;
  assign n665 = n512 & ~n664;
  assign n666 = ~pi48  & ~pi49 ;
  assign n667 = ~n664 & ~n666;
  assign n668 = ~n662 & n666;
  assign n669 = ~n667 & ~n668;
  assign n670 = ~n512 & ~n669;
  assign n671 = ~n665 & ~n670;
  assign n672 = n511 & ~n671;
  assign n673 = ~pi44  & ~pi45 ;
  assign n674 = ~n671 & ~n673;
  assign n675 = ~n669 & n673;
  assign n676 = ~n674 & ~n675;
  assign n677 = ~n511 & ~n676;
  assign n678 = ~n672 & ~n677;
  assign n679 = n510 & ~n678;
  assign n680 = ~pi40  & ~pi41 ;
  assign n681 = ~n678 & ~n680;
  assign n682 = ~n676 & n680;
  assign n683 = ~n681 & ~n682;
  assign n684 = ~n510 & ~n683;
  assign n685 = ~n679 & ~n684;
  assign n686 = n509 & ~n685;
  assign n687 = ~pi36  & ~pi37 ;
  assign n688 = ~n685 & ~n687;
  assign n689 = ~n683 & n687;
  assign n690 = ~n688 & ~n689;
  assign n691 = ~n509 & ~n690;
  assign n692 = ~n686 & ~n691;
  assign n693 = n508 & ~n692;
  assign n694 = ~pi32  & ~pi33 ;
  assign n695 = ~n692 & ~n694;
  assign n696 = ~n690 & n694;
  assign n697 = ~n695 & ~n696;
  assign n698 = ~n508 & ~n697;
  assign n699 = ~n693 & ~n698;
  assign n700 = n507 & ~n699;
  assign n701 = ~pi28  & ~pi29 ;
  assign n702 = ~n699 & ~n701;
  assign n703 = ~n697 & n701;
  assign n704 = ~n702 & ~n703;
  assign n705 = ~n507 & ~n704;
  assign n706 = ~n700 & ~n705;
  assign n707 = n506 & ~n706;
  assign n708 = ~pi24  & ~pi25 ;
  assign n709 = ~n706 & ~n708;
  assign n710 = ~n704 & n708;
  assign n711 = ~n709 & ~n710;
  assign n712 = ~n506 & ~n711;
  assign n713 = ~n707 & ~n712;
  assign n714 = n505 & ~n713;
  assign n715 = ~pi20  & ~pi21 ;
  assign n716 = ~n713 & ~n715;
  assign n717 = ~n711 & n715;
  assign n718 = ~n716 & ~n717;
  assign n719 = ~n505 & ~n718;
  assign n720 = ~n714 & ~n719;
  assign n721 = n504 & ~n720;
  assign n722 = ~pi16  & ~pi17 ;
  assign n723 = ~n720 & ~n722;
  assign n724 = ~n718 & n722;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~n504 & ~n725;
  assign n727 = ~n721 & ~n726;
  assign n728 = n503 & ~n727;
  assign n729 = ~pi12  & ~pi13 ;
  assign n730 = ~n727 & ~n729;
  assign n731 = ~n725 & n729;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~n503 & ~n732;
  assign n734 = ~pi8  & ~pi9 ;
  assign n735 = ~pi6  & ~pi7 ;
  assign n736 = ~pi4  & ~pi5 ;
  assign n737 = ~pi2  & ~pi3 ;
  assign n738 = n736 & ~n737;
  assign n739 = n735 & ~n738;
  assign n740 = n734 & ~n739;
  assign n741 = ~n728 & ~n740;
  assign n742 = ~n733 & n741;
  assign n743 = n732 & n740;
  assign po1  = ~n742 & ~n743;
  assign n745 = n506 & n715;
  assign n746 = n508 & n701;
  assign n747 = n510 & n687;
  assign n748 = n512 & n673;
  assign n749 = n514 & n659;
  assign n750 = n516 & n645;
  assign n751 = n518 & n631;
  assign n752 = n521 & n610;
  assign n753 = n523 & n596;
  assign n754 = n525 & n582;
  assign n755 = n527 & n568;
  assign n756 = n533 & n537;
  assign n757 = n530 & n543;
  assign n758 = ~pi120  & ~pi121 ;
  assign n759 = n531 & n758;
  assign n760 = ~n757 & n759;
  assign n761 = n756 & ~n760;
  assign n762 = ~pi114  & n554;
  assign n763 = n761 & ~n762;
  assign n764 = pi115  & n757;
  assign n765 = n759 & ~n764;
  assign n766 = n756 & n762;
  assign n767 = ~n765 & n766;
  assign n768 = ~n763 & ~n767;
  assign n769 = n755 & ~n768;
  assign n770 = n528 & n561;
  assign n771 = ~n761 & n770;
  assign n772 = n768 & ~n770;
  assign n773 = ~n771 & ~n772;
  assign n774 = ~n755 & n773;
  assign n775 = ~n769 & ~n774;
  assign n776 = n754 & ~n775;
  assign n777 = n526 & n575;
  assign n778 = n775 & ~n777;
  assign n779 = ~n773 & n777;
  assign n780 = ~n778 & ~n779;
  assign n781 = ~n754 & n780;
  assign n782 = ~n776 & ~n781;
  assign n783 = n753 & ~n782;
  assign n784 = n524 & n589;
  assign n785 = ~n780 & n784;
  assign n786 = n782 & ~n784;
  assign n787 = ~n785 & ~n786;
  assign n788 = ~n753 & n787;
  assign n789 = ~n783 & ~n788;
  assign n790 = n752 & ~n789;
  assign n791 = n522 & n603;
  assign n792 = ~n787 & n791;
  assign n793 = n789 & ~n791;
  assign n794 = ~n792 & ~n793;
  assign n795 = ~n752 & n794;
  assign n796 = ~n790 & ~n795;
  assign n797 = n520 & n617;
  assign n798 = n796 & ~n797;
  assign n799 = ~n794 & n797;
  assign n800 = ~n798 & ~n799;
  assign n801 = n751 & ~n800;
  assign n802 = n519 & n624;
  assign n803 = ~n796 & n802;
  assign n804 = n800 & ~n802;
  assign n805 = ~n803 & ~n804;
  assign n806 = ~n751 & n805;
  assign n807 = ~n801 & ~n806;
  assign n808 = n750 & ~n807;
  assign n809 = n517 & n638;
  assign n810 = ~n805 & n809;
  assign n811 = n807 & ~n809;
  assign n812 = ~n810 & ~n811;
  assign n813 = ~n750 & n812;
  assign n814 = ~n808 & ~n813;
  assign n815 = n749 & ~n814;
  assign n816 = n515 & n652;
  assign n817 = ~n812 & n816;
  assign n818 = n814 & ~n816;
  assign n819 = ~n817 & ~n818;
  assign n820 = ~n749 & n819;
  assign n821 = ~n815 & ~n820;
  assign n822 = n748 & ~n821;
  assign n823 = n513 & n666;
  assign n824 = ~n819 & n823;
  assign n825 = n821 & ~n823;
  assign n826 = ~n824 & ~n825;
  assign n827 = ~n748 & n826;
  assign n828 = ~n822 & ~n827;
  assign n829 = n747 & ~n828;
  assign n830 = n511 & n680;
  assign n831 = ~n826 & n830;
  assign n832 = n828 & ~n830;
  assign n833 = ~n831 & ~n832;
  assign n834 = ~n747 & n833;
  assign n835 = ~n829 & ~n834;
  assign n836 = n746 & ~n835;
  assign n837 = n509 & n694;
  assign n838 = ~n833 & n837;
  assign n839 = n835 & ~n837;
  assign n840 = ~n838 & ~n839;
  assign n841 = ~n746 & n840;
  assign n842 = ~n836 & ~n841;
  assign n843 = n745 & ~n842;
  assign n844 = n507 & n708;
  assign n845 = ~n840 & n844;
  assign n846 = n842 & ~n844;
  assign n847 = ~n845 & ~n846;
  assign n848 = ~n745 & n847;
  assign n849 = n505 & n722;
  assign n850 = n504 & n729;
  assign n851 = n503 & n734;
  assign n852 = n735 & n736;
  assign n853 = n851 & ~n852;
  assign n854 = n850 & ~n853;
  assign n855 = n849 & ~n854;
  assign n856 = ~n843 & ~n855;
  assign n857 = ~n848 & n856;
  assign n858 = ~n847 & n855;
  assign po2  = ~n857 & ~n858;
  assign n860 = n748 & n830;
  assign n861 = n750 & n816;
  assign n862 = n752 & n791;
  assign n863 = n756 & n759;
  assign n864 = n755 & n770;
  assign n865 = ~pi115  & n757;
  assign n866 = n762 & n865;
  assign n867 = ~n864 & n866;
  assign n868 = n863 & ~n867;
  assign n869 = ~pi102  & n575;
  assign n870 = n754 & n869;
  assign n871 = n868 & ~n870;
  assign n872 = pi103  & n864;
  assign n873 = n866 & ~n872;
  assign n874 = n863 & n870;
  assign n875 = ~n873 & n874;
  assign n876 = ~n871 & ~n875;
  assign n877 = n862 & ~n876;
  assign n878 = n753 & n784;
  assign n879 = ~n868 & n878;
  assign n880 = n876 & ~n878;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n862 & n881;
  assign n883 = ~n877 & ~n882;
  assign n884 = n797 & n802;
  assign n885 = n883 & ~n884;
  assign n886 = ~n881 & n884;
  assign n887 = ~n885 & ~n886;
  assign n888 = n861 & ~n887;
  assign n889 = n751 & n809;
  assign n890 = ~n883 & n889;
  assign n891 = n887 & ~n889;
  assign n892 = ~n890 & ~n891;
  assign n893 = ~n861 & n892;
  assign n894 = ~n888 & ~n893;
  assign n895 = n860 & ~n894;
  assign n896 = n749 & n823;
  assign n897 = ~n892 & n896;
  assign n898 = n894 & ~n896;
  assign n899 = ~n897 & ~n898;
  assign n900 = ~n860 & n899;
  assign n901 = n747 & n837;
  assign n902 = n746 & n844;
  assign n903 = n745 & n849;
  assign n904 = n850 & n851;
  assign n905 = n903 & ~n904;
  assign n906 = n902 & ~n905;
  assign n907 = n901 & ~n906;
  assign n908 = ~n895 & ~n907;
  assign n909 = ~n900 & n908;
  assign n910 = ~n899 & n907;
  assign po3  = ~n909 & ~n910;
  assign n912 = n863 & n866;
  assign n913 = n862 & n878;
  assign n914 = ~pi103  & n864;
  assign n915 = n870 & n914;
  assign n916 = ~n913 & n915;
  assign n917 = n861 & n896;
  assign n918 = n860 & n901;
  assign n919 = n902 & n903;
  assign n920 = n918 & ~n919;
  assign n921 = n917 & ~n920;
  assign n922 = ~pi78  & n617;
  assign n923 = n802 & n922;
  assign n924 = n889 & n923;
  assign n925 = ~n921 & n924;
  assign n926 = n912 & ~n916;
  assign n927 = ~n925 & n926;
  assign n928 = pi79  & n913;
  assign n929 = n915 & ~n928;
  assign n930 = n912 & ~n929;
  assign n931 = n925 & n930;
  assign po4  = ~n927 & ~n931;
  assign n933 = n912 & n915;
  assign n934 = n917 & n918;
  assign n935 = n884 & n889;
  assign n936 = n913 & n935;
  assign n937 = ~n934 & n936;
  assign po5  = ~n933 | n937;
  assign po6  = ~n933 | ~n936;
  assign n940 = ~pi0  & ~pi1 ;
  assign n941 = n737 & n940;
  assign n942 = n852 & n941;
  assign n943 = n904 & n942;
  assign n944 = n919 & n943;
  assign n945 = n934 & n944;
  assign po7 = po6  | ~n945;
endmodule
