module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 ,
    po6 , po7 , po8 , po9 , po10 ,
    po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 ,
    po21 , po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 , po30 ,
    po31 , po32 , po33 , po34 , po35 ,
    po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 ,
    po46 , po47 , po48 , po49 , po50 ,
    po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 ,
    po61 , po62 , po63   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 ;
  wire n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535,
    n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201,
    n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231,
    n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291,
    n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321,
    n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351,
    n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381,
    n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411,
    n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441,
    n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471,
    n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501,
    n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531,
    n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681,
    n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711,
    n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741,
    n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1771,
    n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801,
    n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831,
    n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843,
    n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861,
    n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873,
    n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921,
    n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951,
    n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981,
    n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101,
    n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131,
    n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161,
    n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173,
    n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191,
    n2192, n2193, n2194, n2195, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203,
    n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221,
    n2222, n2223, n2224, n2225, n2226, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233,
    n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281,
    n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311,
    n2312, n2313, n2314, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2323,
    n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341,
    n2342, n2343, n2344, n2345, n2346, n2347,
    n2348, n2349, n2350, n2351, n2352, n2353,
    n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371,
    n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401,
    n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461,
    n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521,
    n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551,
    n2552, n2553, n2554, n2555, n2556, n2557,
    n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581,
    n2582, n2583, n2584, n2585, n2586, n2587,
    n2588, n2589, n2590, n2591, n2592, n2593,
    n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611,
    n2612, n2613, n2614, n2615, n2616, n2617,
    n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641,
    n2642, n2643, n2644, n2645, n2646, n2647,
    n2648, n2649, n2650, n2651, n2652, n2653,
    n2654, n2655, n2656, n2657, n2658, n2659,
    n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671,
    n2672, n2673, n2674, n2675, n2676, n2677,
    n2678, n2679, n2680, n2681, n2682, n2683,
    n2684, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695,
    n2696, n2697, n2698, n2699, n2700, n2701,
    n2702, n2703, n2704, n2705, n2706, n2707,
    n2708, n2709, n2710, n2711, n2712, n2713,
    n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731,
    n2732, n2733, n2734, n2735, n2736, n2737,
    n2738, n2739, n2740, n2741, n2742, n2743,
    n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761,
    n2762, n2763, n2764, n2765, n2766, n2767,
    n2768, n2769, n2770, n2771, n2772, n2773,
    n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791,
    n2792, n2793, n2794, n2795, n2796, n2797,
    n2798, n2799, n2800, n2801, n2802, n2803,
    n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821,
    n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851,
    n2852, n2853, n2854, n2855, n2856, n2857,
    n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2878, n2879, n2880, n2881,
    n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893,
    n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905,
    n2906, n2907, n2908, n2909, n2910, n2911,
    n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2940, n2941,
    n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953,
    n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971,
    n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001,
    n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013,
    n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031,
    n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055,
    n3056, n3057, n3058, n3059, n3060, n3061,
    n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085,
    n3086, n3087, n3088, n3089, n3090, n3091,
    n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109,
    n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3117, n3118, n3119, n3120, n3121,
    n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151,
    n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3174, n3175,
    n3176, n3177, n3178, n3179, n3180, n3181,
    n3182, n3183, n3184, n3185, n3186, n3187,
    n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211,
    n3212, n3213, n3214, n3215, n3216, n3217,
    n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241,
    n3242, n3243, n3244, n3245, n3246, n3247,
    n3248, n3249, n3250, n3251, n3252, n3253,
    n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265,
    n3266, n3267, n3268, n3269, n3270, n3271,
    n3272, n3273, n3274, n3275, n3276, n3277,
    n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535,
    n3536, n3537, n3538, n3539, n3540, n3541,
    n3542, n3543, n3544, n3545, n3546, n3547,
    n3548, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565,
    n3566, n3567, n3568, n3569, n3570, n3571,
    n3572, n3573, n3574, n3575, n3576, n3577,
    n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601,
    n3602, n3603, n3604, n3605, n3606, n3607,
    n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631,
    n3632, n3633, n3634, n3635, n3636, n3637,
    n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661,
    n3662, n3663, n3664, n3665, n3666, n3667,
    n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691,
    n3692, n3693, n3694, n3695, n3696, n3697,
    n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721,
    n3722, n3723, n3724, n3725, n3726, n3727,
    n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751,
    n3752, n3753, n3754, n3755, n3756, n3757,
    n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775,
    n3776, n3777, n3778, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787,
    n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805,
    n3806, n3807, n3808, n3809, n3810, n3811,
    n3812, n3813, n3814, n3815, n3816, n3817,
    n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835,
    n3836, n3837, n3838, n3839, n3840, n3841,
    n3842, n3843, n3844, n3845, n3846, n3847,
    n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865,
    n3866, n3867, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877,
    n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901,
    n3902, n3903, n3904, n3905, n3906, n3907,
    n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931,
    n3932, n3933, n3934, n3935, n3936, n3937,
    n3938, n3939, n3940, n3941, n3942, n3943,
    n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961,
    n3962, n3963, n3964, n3965, n3966, n3967,
    n3968, n3969, n3970, n3971, n3972, n3973,
    n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985,
    n3986, n3987, n3988, n3989, n3990, n3991,
    n3992, n3993, n3994, n3995, n3996, n3997,
    n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027,
    n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057,
    n4058, n4059, n4060, n4061, n4062, n4063,
    n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4083, n4084, n4085, n4086, n4087,
    n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4095, n4096, n4097, n4098, n4099,
    n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117,
    n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141,
    n4142, n4143, n4144, n4145, n4146, n4147,
    n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171,
    n4172, n4173, n4174, n4175, n4176, n4177,
    n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188, n4189,
    n4190, n4191, n4192, n4193, n4194, n4195,
    n4196, n4197, n4198, n4199, n4200, n4201,
    n4202, n4203, n4204, n4205, n4206, n4207,
    n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219,
    n4220, n4221, n4222, n4223, n4224, n4225,
    n4226, n4227, n4228, n4229, n4230, n4231,
    n4232, n4233, n4234, n4235, n4236, n4237,
    n4238, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249,
    n4250, n4251, n4252, n4253, n4254, n4255,
    n4256, n4257, n4258, n4259, n4260, n4261,
    n4262, n4263, n4264, n4265, n4266, n4267,
    n4268, n4269, n4270, n4271, n4272, n4273,
    n4274, n4275, n4276, n4277, n4278, n4279,
    n4280, n4281, n4282, n4283, n4284, n4285,
    n4286, n4287, n4288, n4289, n4290, n4291,
    n4292, n4293, n4294, n4295, n4296, n4297,
    n4298, n4299, n4300, n4301, n4302, n4303,
    n4304, n4305, n4306, n4307, n4308, n4309,
    n4310, n4311, n4312, n4313, n4314, n4315,
    n4316, n4317, n4318, n4319, n4320, n4321,
    n4322, n4323, n4324, n4325, n4326, n4327,
    n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339,
    n4340, n4341, n4342, n4343, n4344, n4345,
    n4346, n4347, n4348, n4349, n4350, n4351,
    n4352, n4353, n4354, n4355, n4356, n4357,
    n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4368, n4369,
    n4370, n4371, n4372, n4373, n4374, n4375,
    n4376, n4377, n4378, n4379, n4380, n4381,
    n4382, n4383, n4384, n4385, n4386, n4387,
    n4388, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4396, n4397, n4398, n4399,
    n4400, n4401, n4402, n4403, n4404, n4405,
    n4406, n4407, n4408, n4409, n4410, n4411,
    n4412, n4413, n4414, n4415, n4416, n4417,
    n4418, n4419, n4420, n4421, n4422, n4423,
    n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4432, n4433, n4434, n4435,
    n4436, n4437, n4438, n4439, n4440, n4441,
    n4442, n4443, n4444, n4445, n4446, n4447,
    n4448, n4449, n4450, n4451, n4452, n4453,
    n4454, n4455, n4456, n4457, n4458, n4459,
    n4460, n4461, n4462, n4463, n4464, n4465,
    n4466, n4467, n4468, n4469, n4470, n4471,
    n4472, n4473, n4474, n4475, n4476, n4477,
    n4478, n4479, n4480, n4481, n4482, n4483,
    n4484, n4485, n4486, n4487, n4488, n4489,
    n4490, n4491, n4492, n4493, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501,
    n4502, n4503, n4504, n4505, n4506, n4507,
    n4508, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525,
    n4526, n4527, n4528, n4529, n4530, n4531,
    n4532, n4533, n4534, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747,
    n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837,
    n4838, n4839, n4840, n4841, n4842, n4843,
    n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861,
    n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873,
    n4874, n4875, n4876, n4877, n4878, n4879,
    n4880, n4881, n4882, n4883, n4884, n4885,
    n4886, n4887, n4888, n4889, n4890, n4891,
    n4892, n4893, n4894, n4895, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101,
    n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5122, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131,
    n5132, n5133, n5134, n5135, n5136, n5137,
    n5138, n5139, n5140, n5141, n5142, n5143,
    n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161,
    n5162, n5163, n5164, n5165, n5166, n5167,
    n5168, n5169, n5170, n5171, n5172, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179,
    n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191,
    n5192, n5193, n5194, n5195, n5196, n5197,
    n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5205, n5206, n5207, n5208, n5209,
    n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221,
    n5222, n5223, n5224, n5225, n5226, n5227,
    n5228, n5229, n5230, n5231, n5232, n5233,
    n5234, n5235, n5236, n5237, n5238, n5239,
    n5240, n5241, n5242, n5243, n5244, n5245,
    n5246, n5247, n5248, n5249, n5250, n5251,
    n5252, n5253, n5254, n5255, n5256, n5257,
    n5258, n5259, n5260, n5261, n5262, n5263,
    n5264, n5265, n5266, n5267, n5268, n5269,
    n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281,
    n5282, n5283, n5284, n5285, n5286, n5287,
    n5288, n5289, n5290, n5291, n5292, n5293,
    n5294, n5295, n5296, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305,
    n5306, n5307, n5308, n5309, n5310, n5311,
    n5312, n5313, n5314, n5315, n5316, n5317,
    n5318, n5319, n5320, n5321, n5322, n5323,
    n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5333, n5334, n5335,
    n5336, n5337, n5338, n5339, n5340, n5341,
    n5342, n5343, n5344, n5345, n5346, n5347,
    n5348, n5349, n5350, n5351, n5352, n5353,
    n5354, n5355, n5356, n5357, n5358, n5359,
    n5360, n5361, n5362, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371,
    n5372, n5373, n5374, n5375, n5376, n5377,
    n5378, n5379, n5380, n5381, n5382, n5383,
    n5384, n5385, n5386, n5387, n5388, n5389,
    n5390, n5391, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401,
    n5402, n5403, n5404, n5405, n5406, n5407,
    n5408, n5409, n5410, n5411, n5412, n5413,
    n5414, n5415, n5416, n5417, n5418, n5419,
    n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431,
    n5432, n5433, n5434, n5435, n5436, n5437,
    n5438, n5439, n5440, n5441, n5442, n5443,
    n5444, n5445, n5446, n5447, n5448, n5449,
    n5450, n5451, n5452, n5453, n5454, n5455,
    n5456, n5457, n5458, n5459, n5460, n5461,
    n5462, n5463, n5464, n5465, n5466, n5467,
    n5468, n5469, n5470, n5471, n5472, n5473,
    n5474, n5475, n5476, n5477, n5478, n5479,
    n5480, n5481, n5482, n5483, n5484, n5485,
    n5486, n5487, n5488, n5489, n5490, n5491,
    n5492, n5493, n5494, n5495, n5496, n5497,
    n5498, n5499, n5500, n5501, n5502, n5503,
    n5504, n5505, n5506, n5507, n5508, n5509,
    n5510, n5511, n5512, n5513, n5514, n5515,
    n5516, n5517, n5518, n5519, n5520, n5521,
    n5522, n5523, n5524, n5525, n5526, n5527,
    n5528, n5529, n5530, n5531, n5532, n5533,
    n5534, n5535, n5536, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551,
    n5552, n5553, n5554, n5555, n5556, n5557,
    n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581,
    n5582, n5583, n5584, n5585, n5586, n5587,
    n5588, n5589, n5590, n5591, n5592, n5593,
    n5594, n5595, n5596, n5597, n5598, n5599,
    n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611,
    n5612, n5613, n5614, n5615, n5616, n5617,
    n5618, n5619, n5620, n5621, n5622, n5623,
    n5624, n5625, n5626, n5627, n5628, n5629,
    n5630, n5631, n5632, n5633, n5634, n5635,
    n5636, n5637, n5638, n5639, n5640, n5641,
    n5642, n5643, n5644, n5645, n5646, n5647,
    n5648, n5649, n5650, n5651, n5652, n5653,
    n5654, n5655, n5656, n5657, n5658, n5659,
    n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5667, n5668, n5669, n5670, n5671,
    n5672, n5673, n5674, n5675, n5676, n5677,
    n5678, n5679, n5680, n5681, n5682, n5683,
    n5684, n5685, n5686, n5687, n5688, n5689,
    n5690, n5691, n5692, n5693, n5694, n5695,
    n5696, n5697, n5698, n5699, n5700, n5701,
    n5702, n5703, n5704, n5705, n5706, n5707,
    n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5715, n5716, n5717, n5718, n5719,
    n5720, n5721, n5722, n5723, n5724, n5725,
    n5726, n5727, n5728, n5729, n5730, n5731,
    n5732, n5733, n5734, n5735, n5736, n5737,
    n5738, n5739, n5740, n5741, n5742, n5743,
    n5744, n5745, n5746, n5747, n5748, n5749,
    n5750, n5751, n5752, n5753, n5754, n5755,
    n5756, n5757, n5758, n5759, n5760, n5761,
    n5762, n5763, n5764, n5765, n5766, n5767,
    n5768, n5769, n5770, n5771, n5772, n5773,
    n5774, n5775, n5776, n5777, n5778, n5779,
    n5780, n5781, n5782, n5783, n5784, n5785,
    n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5794, n5795, n5796, n5797,
    n5798, n5799, n5800, n5801, n5802, n5803,
    n5804, n5805, n5806, n5807, n5808, n5809,
    n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5817, n5818, n5819, n5820, n5821,
    n5822, n5823, n5824, n5825, n5826, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833,
    n5834, n5835, n5836, n5837, n5838, n5839,
    n5840, n5841, n5842, n5843, n5844, n5845,
    n5846, n5847, n5848, n5849, n5850, n5851,
    n5852, n5853, n5854, n5855, n5856, n5857,
    n5858, n5859, n5860, n5861, n5862, n5863,
    n5864, n5865, n5866, n5867, n5868, n5869,
    n5870, n5871, n5872, n5873, n5874, n5875,
    n5876, n5877, n5878, n5879, n5880, n5881,
    n5882, n5883, n5884, n5885, n5886, n5887,
    n5888, n5889, n5890, n5891, n5892, n5893,
    n5894, n5895, n5896, n5897, n5898, n5899,
    n5900, n5901, n5902, n5903, n5904, n5905,
    n5906, n5907, n5908, n5909, n5910, n5911,
    n5912, n5913, n5914, n5915, n5916, n5917,
    n5918, n5919, n5920, n5921, n5922, n5923,
    n5924, n5925, n5926, n5927, n5928, n5929,
    n5930, n5931, n5932, n5933, n5934, n5935,
    n5936, n5937, n5938, n5939, n5940, n5941,
    n5942, n5943, n5944, n5945, n5946, n5947,
    n5948, n5949, n5950, n5951, n5952, n5953,
    n5954, n5955, n5956, n5957, n5958, n5959,
    n5960, n5961, n5962, n5963, n5964, n5965,
    n5966, n5967, n5968, n5969, n5970, n5971,
    n5972, n5973, n5974, n5975, n5976, n5977,
    n5978, n5979, n5980, n5981, n5982, n5983,
    n5984, n5985, n5986, n5987, n5988, n5989,
    n5990, n5991, n5992, n5993, n5994, n5995,
    n5996, n5997, n5998, n5999, n6000, n6001,
    n6002, n6003, n6004, n6005, n6006, n6007,
    n6008, n6009, n6010, n6011, n6012, n6013,
    n6014, n6015, n6016, n6017, n6018, n6019,
    n6020, n6021, n6022, n6023, n6024, n6025,
    n6026, n6027, n6028, n6029, n6030, n6031,
    n6032, n6033, n6034, n6035, n6036, n6037,
    n6038, n6039, n6040, n6041, n6042, n6043,
    n6044, n6045, n6046, n6047, n6048, n6049,
    n6050, n6051, n6052, n6053, n6054, n6055,
    n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067,
    n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079,
    n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097,
    n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6126, n6127,
    n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145,
    n6146, n6147, n6148, n6149, n6150, n6151,
    n6152, n6153, n6154, n6155, n6156, n6157,
    n6158, n6159, n6160, n6161, n6162, n6163,
    n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175,
    n6176, n6177, n6178, n6179, n6180, n6181,
    n6182, n6183, n6184, n6185, n6186, n6187,
    n6188, n6189, n6190, n6191, n6192, n6193,
    n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6202, n6203, n6204, n6205,
    n6206, n6207, n6208, n6209, n6210, n6211,
    n6212, n6213, n6214, n6215, n6216, n6217,
    n6218, n6219, n6220, n6221, n6222, n6223,
    n6224, n6225, n6226, n6227, n6228, n6229,
    n6230, n6231, n6232, n6233, n6234, n6235,
    n6236, n6237, n6238, n6239, n6240, n6241,
    n6242, n6243, n6244, n6245, n6246, n6247,
    n6248, n6249, n6250, n6251, n6252, n6253,
    n6254, n6255, n6256, n6257, n6258, n6259,
    n6260, n6261, n6262, n6263, n6264, n6265,
    n6266, n6267, n6268, n6269, n6270, n6271,
    n6272, n6273, n6274, n6275, n6276, n6277,
    n6278, n6279, n6280, n6281, n6282, n6283,
    n6284, n6285, n6286, n6287, n6288, n6289,
    n6290, n6291, n6292, n6293, n6294, n6295,
    n6296, n6297, n6298, n6299, n6300, n6301,
    n6302, n6303, n6304, n6305, n6306, n6307,
    n6308, n6309, n6310, n6311, n6312, n6313,
    n6314, n6315, n6316, n6317, n6318, n6319,
    n6320, n6321, n6322, n6323, n6324, n6325,
    n6326, n6327, n6328, n6329, n6330, n6331,
    n6332, n6333, n6334, n6335, n6336, n6337,
    n6338, n6339, n6340, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349,
    n6350, n6351, n6352, n6353, n6354, n6355,
    n6356, n6357, n6358, n6359, n6360, n6361,
    n6362, n6363, n6364, n6365, n6366, n6367,
    n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379,
    n6380, n6381, n6382, n6383, n6384, n6385,
    n6386, n6387, n6388, n6389, n6390, n6391,
    n6392, n6393, n6394, n6395, n6396, n6397,
    n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409,
    n6410, n6411, n6412, n6413, n6414, n6415,
    n6416, n6417, n6418, n6419, n6420, n6421,
    n6422, n6423, n6424, n6425, n6426, n6427,
    n6428, n6429, n6430, n6431, n6432, n6433,
    n6434, n6435, n6436, n6437, n6438, n6439,
    n6440, n6441, n6442, n6443, n6444, n6445,
    n6446, n6447, n6448, n6449, n6450, n6451,
    n6452, n6453, n6454, n6455, n6456, n6457,
    n6458, n6459, n6460, n6461, n6462, n6463,
    n6464, n6465, n6466, n6467, n6468, n6469,
    n6470, n6471, n6472, n6473, n6474, n6475,
    n6476, n6477, n6478, n6479, n6480, n6481,
    n6482, n6483, n6484, n6485, n6486, n6487,
    n6488, n6489, n6490, n6491, n6492, n6493,
    n6494, n6495, n6496, n6497, n6498, n6499,
    n6500, n6501, n6502, n6503, n6504, n6505,
    n6506, n6507, n6508, n6509, n6510, n6511,
    n6512, n6513, n6514, n6515, n6516, n6517,
    n6518, n6519, n6520, n6521, n6522, n6523,
    n6524, n6525, n6526, n6527, n6528, n6529,
    n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541,
    n6542, n6543, n6544, n6545, n6546, n6547,
    n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571,
    n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601,
    n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631,
    n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649,
    n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661,
    n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679,
    n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691,
    n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6702, n6703,
    n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721,
    n6722, n6723, n6724, n6725, n6726, n6727,
    n6728, n6729, n6730, n6731, n6732, n6733,
    n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751,
    n6752, n6753, n6754, n6755, n6756, n6757,
    n6758, n6759, n6760, n6761, n6762, n6763,
    n6764, n6765, n6766, n6767, n6768, n6769,
    n6770, n6771, n6772, n6773, n6774, n6775,
    n6776, n6777, n6778, n6779, n6780, n6781,
    n6782, n6783, n6784, n6785, n6786, n6787,
    n6788, n6789, n6790, n6791, n6792, n6793,
    n6794, n6795, n6796, n6797, n6798, n6799,
    n6800, n6801, n6802, n6803, n6804, n6805,
    n6806, n6807, n6808, n6809, n6810, n6811,
    n6812, n6813, n6814, n6815, n6816, n6817,
    n6818, n6819, n6820, n6821, n6822, n6823,
    n6824, n6825, n6826, n6827, n6828, n6829,
    n6830, n6831, n6832, n6833, n6834, n6835,
    n6836, n6837, n6838, n6839, n6840, n6841,
    n6842, n6843, n6844, n6845, n6846, n6847,
    n6848, n6849, n6850, n6851, n6852, n6853,
    n6854, n6855, n6856, n6857, n6858, n6859,
    n6860, n6861, n6862, n6863, n6864, n6865,
    n6866, n6867, n6868, n6869, n6870, n6871,
    n6872, n6873, n6874, n6875, n6876, n6877,
    n6878, n6879, n6880, n6881, n6882, n6883,
    n6884, n6885, n6886, n6887, n6888, n6889,
    n6890, n6891, n6892, n6893, n6894, n6895,
    n6896, n6897, n6898, n6899, n6900, n6901,
    n6902, n6903, n6904, n6905, n6906, n6907,
    n6908, n6909, n6910, n6911, n6912, n6913,
    n6914, n6915, n6916, n6917, n6918, n6919,
    n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931,
    n6932, n6933, n6934, n6935, n6936, n6937,
    n6938, n6939, n6940, n6941, n6942, n6943,
    n6944, n6945, n6946, n6947, n6948, n6949,
    n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961,
    n6962, n6963, n6964, n6965, n6966, n6967,
    n6968, n6969, n6970, n6971, n6972, n6973,
    n6974, n6975, n6976, n6977, n6978, n6979,
    n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991,
    n6992, n6993, n6994, n6995, n6996, n6997,
    n6998, n6999, n7000, n7001, n7002, n7003,
    n7004, n7005, n7006, n7007, n7008, n7009,
    n7010, n7011, n7012, n7013, n7014, n7015,
    n7016, n7017, n7018, n7019, n7020, n7021,
    n7022, n7023, n7024, n7025, n7026, n7027,
    n7028, n7029, n7030, n7031, n7032, n7033,
    n7034, n7035, n7036, n7037, n7038, n7039,
    n7040, n7041, n7042, n7043, n7044, n7045,
    n7046, n7047, n7048, n7049, n7050, n7051,
    n7052, n7053, n7054, n7055, n7056, n7057,
    n7058, n7059, n7060, n7061, n7062, n7063,
    n7064, n7065, n7066, n7067, n7068, n7069,
    n7070, n7071, n7072, n7073, n7074, n7075,
    n7076, n7077, n7078, n7079, n7080, n7081,
    n7082, n7083, n7084, n7085, n7086, n7087,
    n7088, n7089, n7090, n7091, n7092, n7093,
    n7094, n7095, n7096, n7097, n7098, n7099,
    n7100, n7101, n7102, n7103, n7104, n7105,
    n7106, n7107, n7108, n7109, n7110, n7111,
    n7112, n7113, n7114, n7115, n7116, n7117,
    n7118, n7119, n7120, n7121, n7122, n7123,
    n7124, n7125, n7126, n7127, n7128, n7129,
    n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7137, n7138, n7139, n7140, n7141,
    n7142, n7143, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153,
    n7154, n7155, n7156, n7157, n7158, n7159,
    n7160, n7161, n7162, n7163, n7164, n7165,
    n7166, n7167, n7168, n7169, n7170, n7171,
    n7172, n7173, n7174, n7175, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7194, n7195,
    n7196, n7197, n7198, n7199, n7200, n7201,
    n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7227, n7228, n7229, n7230, n7231,
    n7232, n7233, n7234, n7235, n7236, n7237,
    n7238, n7239, n7240, n7241, n7242, n7243,
    n7244, n7245, n7246, n7247, n7248, n7249,
    n7250, n7251, n7252, n7253, n7254, n7255,
    n7256, n7257, n7258, n7259, n7260, n7261,
    n7262, n7263, n7264, n7265, n7266, n7267,
    n7268, n7269, n7270, n7271, n7272, n7273,
    n7274, n7275, n7276, n7277, n7278, n7279,
    n7280, n7281, n7282, n7283, n7284, n7285,
    n7286, n7287, n7288, n7289, n7290, n7291,
    n7292, n7293, n7294, n7295, n7296, n7297,
    n7298, n7299, n7300, n7301, n7302, n7303,
    n7304, n7305, n7306, n7307, n7308, n7309,
    n7310, n7311, n7312, n7313, n7314, n7315,
    n7316, n7317, n7318, n7319, n7320, n7321,
    n7322, n7323, n7324, n7325, n7326, n7327,
    n7328, n7329, n7330, n7331, n7332, n7333,
    n7334, n7335, n7336, n7337, n7338, n7339,
    n7340, n7341, n7342, n7343, n7344, n7345,
    n7346, n7347, n7348, n7349, n7350, n7351,
    n7352, n7353, n7354, n7355, n7356, n7357,
    n7358, n7359, n7360, n7361, n7362, n7363,
    n7364, n7365, n7366, n7367, n7368, n7369,
    n7370, n7371, n7372, n7373, n7374, n7375,
    n7376, n7377, n7378, n7379, n7380, n7381,
    n7382, n7383, n7384, n7385, n7386, n7387,
    n7388, n7389, n7390, n7391, n7392, n7393,
    n7394, n7395, n7396, n7397, n7398, n7399,
    n7400, n7401, n7402, n7403, n7404, n7405,
    n7406, n7407, n7408, n7409, n7410, n7411,
    n7412, n7413, n7414, n7415, n7416, n7417,
    n7418, n7419, n7420, n7421, n7422, n7423,
    n7424, n7425, n7426, n7427, n7428, n7429,
    n7430, n7431, n7432, n7433, n7434, n7435,
    n7436, n7437, n7438, n7439, n7440, n7441,
    n7442, n7443, n7444, n7445, n7446, n7447,
    n7448, n7449, n7450, n7451, n7452, n7453,
    n7454, n7455, n7456, n7457, n7458, n7459,
    n7460, n7461, n7462, n7463, n7464, n7465,
    n7466, n7467, n7468, n7469, n7470, n7471,
    n7472, n7473, n7474, n7475, n7476, n7477,
    n7478, n7479, n7480, n7481, n7482, n7483,
    n7484, n7485, n7486, n7487, n7488, n7489,
    n7490, n7491, n7492, n7493, n7494, n7495,
    n7496, n7497, n7498, n7499, n7500, n7501,
    n7502, n7503, n7504, n7505, n7506, n7507,
    n7508, n7509, n7510, n7511, n7512, n7513,
    n7514, n7515, n7516, n7517, n7518, n7519,
    n7520, n7521, n7522, n7523, n7524, n7525,
    n7526, n7527, n7528, n7529, n7530, n7531,
    n7532, n7533, n7534, n7535, n7536, n7537,
    n7538, n7539, n7540, n7541, n7542, n7543,
    n7544, n7545, n7546, n7547, n7548, n7549,
    n7550, n7551, n7552, n7553, n7554, n7555,
    n7556, n7557, n7558, n7559, n7560, n7561,
    n7562, n7563, n7564, n7565, n7566, n7567,
    n7568, n7569, n7570, n7571, n7572, n7573,
    n7574, n7575, n7576, n7577, n7578, n7579,
    n7580, n7581, n7582, n7583, n7584, n7585,
    n7586, n7587, n7588, n7589, n7590, n7591,
    n7592, n7593, n7594, n7595, n7596, n7597,
    n7598, n7599, n7600, n7601, n7602, n7603,
    n7604, n7605, n7606, n7607, n7608, n7609,
    n7610, n7611, n7612, n7613, n7614, n7615,
    n7616, n7617, n7618, n7619, n7620, n7621,
    n7622, n7623, n7624, n7625, n7626, n7627,
    n7628, n7629, n7630, n7631, n7632, n7633,
    n7634, n7635, n7636, n7637, n7638, n7639,
    n7640, n7641, n7642, n7643, n7644, n7645,
    n7646, n7647, n7648, n7649, n7650, n7651,
    n7652, n7653, n7654, n7655, n7656, n7657,
    n7658, n7659, n7660, n7661, n7662, n7663,
    n7664, n7665, n7666, n7667, n7668, n7669,
    n7670, n7671, n7672, n7673, n7674, n7675,
    n7676, n7677, n7678, n7679, n7680, n7681,
    n7682, n7683, n7684, n7685, n7686, n7687,
    n7688, n7689, n7690, n7691, n7692, n7693,
    n7694, n7695, n7696, n7697, n7698, n7699,
    n7700, n7701, n7702, n7703, n7704, n7705,
    n7706, n7707, n7708, n7709, n7710, n7711,
    n7712, n7713, n7714, n7715, n7716, n7717,
    n7718, n7719, n7720, n7721, n7722, n7723,
    n7724, n7725, n7726, n7727, n7728, n7729,
    n7730, n7731, n7732, n7733, n7734, n7735,
    n7736, n7737, n7738, n7739, n7740, n7741,
    n7742, n7743, n7744, n7745, n7746, n7747,
    n7748, n7749, n7750, n7751, n7752, n7753,
    n7754, n7755, n7756, n7757, n7758, n7759,
    n7760, n7761, n7762, n7763, n7764, n7765,
    n7766, n7767, n7768, n7769, n7770, n7771,
    n7772, n7773, n7774, n7775, n7776, n7777,
    n7778, n7779, n7780, n7781, n7782, n7783,
    n7784, n7785, n7786, n7787, n7788, n7789,
    n7790, n7791, n7792, n7793, n7794, n7795,
    n7796, n7797, n7798, n7799, n7800, n7801,
    n7802, n7803, n7804, n7805, n7806, n7807,
    n7808, n7809, n7810, n7811, n7812, n7813,
    n7814, n7815, n7816, n7817, n7818, n7819,
    n7820, n7821, n7822, n7823, n7824, n7825,
    n7826, n7827, n7828, n7829, n7830, n7831,
    n7832, n7833, n7834, n7835, n7836, n7837,
    n7838, n7839, n7840, n7841, n7842, n7843,
    n7844, n7845, n7846, n7847, n7848, n7849,
    n7850, n7851, n7852, n7853, n7854, n7855,
    n7856, n7857, n7858, n7859, n7860, n7861,
    n7862, n7863, n7864, n7865, n7866, n7867,
    n7868, n7869, n7870, n7871, n7872, n7873,
    n7874, n7875, n7876, n7877, n7878, n7879,
    n7880, n7881, n7882, n7883, n7884, n7885,
    n7886, n7887, n7888, n7889, n7890, n7891,
    n7892, n7893, n7894, n7895, n7896, n7897,
    n7898, n7899, n7900, n7901, n7902, n7903,
    n7904, n7905, n7906, n7907, n7908, n7909,
    n7910, n7911, n7912, n7913, n7914, n7915,
    n7916, n7917, n7918, n7919, n7920, n7921,
    n7922, n7923, n7924, n7925, n7926, n7927,
    n7928, n7929, n7930, n7931, n7932, n7933,
    n7934, n7935, n7936, n7937, n7938, n7939,
    n7940, n7941, n7942, n7943, n7944, n7945,
    n7946, n7947, n7948, n7949, n7950, n7951,
    n7952, n7953, n7954, n7955, n7956, n7957,
    n7958, n7959, n7960, n7961, n7962, n7963,
    n7964, n7965, n7966, n7967, n7968, n7969,
    n7970, n7971, n7972, n7973, n7974, n7975,
    n7976, n7977, n7978, n7979, n7980, n7981,
    n7982, n7983, n7984, n7985, n7986, n7987,
    n7988, n7989, n7990, n7991, n7992, n7993,
    n7994, n7995, n7996, n7997, n7998, n7999,
    n8000, n8001, n8002, n8003, n8004, n8005,
    n8006, n8007, n8008, n8009, n8010, n8011,
    n8012, n8013, n8014, n8015, n8016, n8017,
    n8018, n8019, n8020, n8021, n8022, n8023,
    n8024, n8025, n8026, n8027, n8028, n8029,
    n8030, n8031, n8032, n8033, n8034, n8035,
    n8036, n8037, n8038, n8039, n8040, n8041,
    n8042, n8043, n8044, n8045, n8046, n8047,
    n8048, n8049, n8050, n8051, n8052, n8053,
    n8054, n8055, n8056, n8057, n8058, n8059,
    n8060, n8061, n8062, n8063, n8064, n8065,
    n8066, n8067, n8068, n8069, n8070, n8071,
    n8072, n8073, n8074, n8075, n8076, n8077,
    n8078, n8079, n8080, n8081, n8082, n8083,
    n8084, n8085, n8086, n8087, n8088, n8089,
    n8090, n8091, n8092, n8093, n8094, n8095,
    n8096, n8097, n8098, n8099, n8100, n8101,
    n8102, n8103, n8104, n8105, n8106, n8107,
    n8108, n8109, n8110, n8111, n8112, n8113,
    n8114, n8115, n8116, n8117, n8118, n8119,
    n8120, n8121, n8122, n8123, n8124, n8125,
    n8126, n8127, n8128, n8129, n8130, n8131,
    n8132, n8133, n8134, n8135, n8136, n8137,
    n8138, n8139, n8140, n8141, n8142, n8143,
    n8144, n8145, n8146, n8147, n8148, n8149,
    n8150, n8151, n8152, n8153, n8154, n8155,
    n8156, n8157, n8158, n8159, n8160, n8161,
    n8162, n8163, n8164, n8165, n8166, n8167,
    n8168, n8169, n8170, n8171, n8172, n8173,
    n8174, n8175, n8176, n8177, n8178, n8179,
    n8180, n8181, n8182, n8183, n8184, n8185,
    n8186, n8187, n8188, n8189, n8190, n8191,
    n8192, n8193, n8194, n8195, n8196, n8197,
    n8198, n8199, n8200, n8201, n8202, n8203,
    n8204, n8205, n8206, n8207, n8208, n8209,
    n8210, n8211, n8212, n8213, n8214, n8215,
    n8216, n8217, n8218, n8219, n8220, n8221,
    n8222, n8223, n8224, n8225, n8226, n8227,
    n8228, n8229, n8230, n8231, n8232, n8233,
    n8234, n8235, n8236, n8237, n8238, n8239,
    n8240, n8241, n8242, n8243, n8244, n8245,
    n8246, n8247, n8248, n8249, n8250, n8251,
    n8252, n8253, n8254, n8255, n8256, n8257,
    n8258, n8259, n8260, n8261, n8262, n8263,
    n8264, n8265, n8266, n8267, n8268, n8269,
    n8270, n8271, n8272, n8273, n8274, n8275,
    n8276, n8277, n8278, n8279, n8280, n8281,
    n8282, n8283, n8284, n8285, n8286, n8287,
    n8288, n8289, n8290, n8291, n8292, n8293,
    n8294, n8295, n8296, n8297, n8298, n8299,
    n8300, n8301, n8302, n8303, n8304, n8305,
    n8306, n8307, n8308, n8309, n8310, n8311,
    n8312, n8313, n8314, n8315, n8316, n8317,
    n8318, n8319, n8320, n8321, n8322, n8323,
    n8324, n8325, n8326, n8327, n8328, n8329,
    n8330, n8331, n8332, n8333, n8334, n8335,
    n8336, n8337, n8338, n8339, n8340, n8341,
    n8342, n8343, n8344, n8345, n8346, n8347,
    n8348, n8349, n8350, n8351, n8352, n8353,
    n8354, n8355, n8356, n8357, n8358, n8359,
    n8360, n8361, n8362, n8363, n8364, n8365,
    n8366, n8367, n8368, n8369, n8370, n8371,
    n8372, n8373, n8374, n8375, n8376, n8377,
    n8378, n8379, n8380, n8381, n8382, n8383,
    n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8391, n8392, n8393, n8394, n8395,
    n8396, n8397, n8398, n8399, n8400, n8401,
    n8402, n8403, n8404, n8405, n8406, n8407,
    n8408, n8409, n8410, n8411, n8412, n8413,
    n8414, n8415, n8416, n8417, n8418, n8419,
    n8420, n8421, n8422, n8423, n8424, n8425,
    n8426, n8427, n8428, n8429, n8430, n8431,
    n8432, n8433, n8434, n8435, n8436, n8437,
    n8438, n8439, n8440, n8441, n8442, n8443,
    n8444, n8445, n8446, n8447, n8448, n8449,
    n8450, n8451, n8452, n8453, n8454, n8455,
    n8456, n8457, n8458, n8459, n8460, n8461,
    n8462, n8463, n8464, n8465, n8466, n8467,
    n8468, n8469, n8470, n8471, n8472, n8473,
    n8474, n8475, n8476, n8477, n8478, n8479,
    n8480, n8481, n8482, n8483, n8484, n8485,
    n8486, n8487, n8488, n8489, n8490, n8491,
    n8492, n8493, n8494, n8495, n8496, n8497,
    n8498, n8499, n8500, n8501, n8502, n8503,
    n8504, n8505, n8506, n8507, n8508, n8509,
    n8510, n8511, n8512, n8513, n8514, n8515,
    n8516, n8517, n8518, n8519, n8520, n8521,
    n8522, n8523, n8524, n8525, n8526, n8527,
    n8528, n8529, n8530, n8531, n8532, n8533,
    n8534, n8535, n8536, n8537, n8538, n8539,
    n8540, n8541, n8542, n8543, n8544, n8545,
    n8546, n8547, n8548, n8549, n8550, n8551,
    n8552, n8553, n8554, n8555, n8556, n8557,
    n8558, n8559, n8560, n8561, n8562, n8563,
    n8564, n8565, n8566, n8567, n8568, n8569,
    n8570, n8571, n8572, n8573, n8574, n8575,
    n8576, n8577, n8578, n8579, n8580, n8581,
    n8582, n8583, n8584, n8585, n8586, n8587,
    n8588, n8589, n8590, n8591, n8592, n8593,
    n8594, n8595, n8596, n8597, n8598, n8599,
    n8600, n8601, n8602, n8603, n8604, n8605,
    n8606, n8607, n8608, n8609, n8610, n8611,
    n8612, n8613, n8614, n8615, n8616, n8617,
    n8618, n8619, n8620, n8621, n8622, n8623,
    n8624, n8625, n8626, n8627, n8628, n8629,
    n8630, n8631, n8632, n8633, n8634, n8635,
    n8636, n8637, n8638, n8639, n8640, n8641,
    n8642, n8643, n8644, n8645, n8646, n8647,
    n8648, n8649, n8650, n8651, n8652, n8653,
    n8654, n8655, n8656, n8657, n8658, n8659,
    n8660, n8661, n8662, n8663, n8664, n8665,
    n8666, n8667, n8668, n8669, n8670, n8671,
    n8672, n8673, n8674, n8675, n8676, n8677,
    n8678, n8679, n8680, n8681, n8682, n8683,
    n8684, n8685, n8686, n8687, n8688, n8689,
    n8690, n8691, n8692, n8693, n8694, n8695,
    n8696, n8697, n8698, n8699, n8700, n8701,
    n8702, n8703, n8704, n8705, n8706, n8707,
    n8708, n8709, n8710, n8711, n8712, n8713,
    n8714, n8715, n8716, n8717, n8718, n8719,
    n8720, n8721, n8722, n8723, n8724, n8725,
    n8726, n8727, n8728, n8729, n8730, n8731,
    n8732, n8733, n8734, n8735, n8736, n8737,
    n8738, n8739, n8740, n8741, n8742, n8743,
    n8744, n8745, n8746, n8747, n8748, n8749,
    n8750, n8751, n8752, n8753, n8754, n8755,
    n8756, n8757, n8758, n8759, n8760, n8761,
    n8762, n8763, n8764, n8765, n8766, n8767,
    n8768, n8769, n8770, n8771, n8772, n8773,
    n8774, n8775, n8776, n8777, n8778, n8779,
    n8780, n8781, n8782, n8783, n8784, n8785,
    n8786, n8787, n8788, n8789, n8790, n8791,
    n8792, n8793, n8794, n8795, n8796, n8797,
    n8798, n8799, n8800, n8801, n8802, n8803,
    n8804, n8805, n8806, n8807, n8808, n8809,
    n8810, n8811, n8812, n8813, n8814, n8815,
    n8816, n8817, n8818, n8819, n8820, n8821,
    n8822, n8823, n8824, n8825, n8826, n8827,
    n8828, n8829, n8830, n8831, n8832, n8833,
    n8834, n8835, n8836, n8837, n8838, n8839,
    n8840, n8841, n8842, n8843, n8844, n8845,
    n8846, n8847, n8848, n8849, n8850, n8851,
    n8852, n8853, n8854, n8855, n8856, n8857,
    n8858, n8859, n8860, n8861, n8862, n8863,
    n8864, n8865, n8866, n8867, n8868, n8869,
    n8870, n8871, n8872, n8873, n8874, n8875,
    n8876, n8877, n8878, n8879, n8880, n8881,
    n8882, n8883, n8884, n8885, n8886, n8887,
    n8888, n8889, n8890, n8891, n8892, n8893,
    n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905,
    n8906, n8907, n8908, n8909, n8910, n8911,
    n8912, n8913, n8914, n8915, n8916, n8917,
    n8918, n8919, n8920, n8921, n8922, n8923,
    n8924, n8925, n8926, n8927, n8928, n8929,
    n8930, n8931, n8932, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8940, n8941,
    n8942, n8943, n8944, n8945, n8946, n8947,
    n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8956, n8957, n8958, n8959,
    n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971,
    n8972, n8973, n8974, n8975, n8976, n8977,
    n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989,
    n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001,
    n9002, n9003, n9004, n9005, n9006, n9007,
    n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019,
    n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031,
    n9032, n9033, n9034, n9035, n9036, n9037,
    n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061,
    n9062, n9063, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073,
    n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121,
    n9122, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151,
    n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259,
    n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271,
    n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289,
    n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301,
    n9302, n9303, n9304, n9305, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9313,
    n9314, n9315, n9316, n9317, n9318, n9319,
    n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331,
    n9332, n9333, n9334, n9335, n9336, n9337,
    n9338, n9339, n9340, n9341, n9342, n9343,
    n9344, n9345, n9346, n9347, n9348, n9349,
    n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361,
    n9362, n9363, n9364, n9365, n9366, n9367,
    n9368, n9369, n9370, n9371, n9372, n9373,
    n9374, n9375, n9376, n9377, n9378, n9379,
    n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391,
    n9392, n9393, n9394, n9395, n9396, n9397,
    n9398, n9399, n9400, n9401, n9402, n9403,
    n9404, n9405, n9406, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421,
    n9422, n9423, n9424, n9425, n9426, n9427,
    n9428, n9429, n9430, n9431, n9432, n9433,
    n9434, n9435, n9436, n9437, n9438, n9439,
    n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451,
    n9452, n9453, n9454, n9455, n9456, n9457,
    n9458, n9459, n9460, n9461, n9462, n9463,
    n9464, n9465, n9466, n9467, n9468, n9469,
    n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481,
    n9482, n9483, n9484, n9485, n9486, n9487,
    n9488, n9489, n9490, n9491, n9492, n9493,
    n9494, n9495, n9496, n9497, n9498, n9499,
    n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511,
    n9512, n9513, n9514, n9515, n9516, n9517,
    n9518, n9519, n9520, n9521, n9522, n9523,
    n9524, n9525, n9526, n9527, n9528, n9529,
    n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541,
    n9542, n9543, n9544, n9545, n9546, n9547,
    n9548, n9549, n9550, n9551, n9552, n9553,
    n9554, n9555, n9556, n9557, n9558, n9559,
    n9560, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9570, n9571,
    n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583,
    n9584, n9585, n9586, n9587, n9588, n9589,
    n9590, n9591, n9592, n9593, n9594, n9595,
    n9596, n9597, n9598, n9599, n9600, n9601,
    n9602, n9603, n9604, n9605, n9606, n9607,
    n9608, n9609, n9610, n9611, n9612, n9613,
    n9614, n9615, n9616, n9617, n9618, n9619,
    n9620, n9621, n9622, n9623, n9624, n9625,
    n9626, n9627, n9628, n9629, n9630, n9631,
    n9632, n9633, n9634, n9635, n9636, n9637,
    n9638, n9639, n9640, n9641, n9642, n9643,
    n9644, n9645, n9646, n9647, n9648, n9649,
    n9650, n9651, n9652, n9653, n9654, n9655,
    n9656, n9657, n9658, n9659, n9660, n9661,
    n9662, n9663, n9664, n9665, n9666, n9667,
    n9668, n9669, n9670, n9671, n9672, n9673,
    n9674, n9675, n9676, n9677, n9678, n9679,
    n9680, n9681, n9682, n9683, n9684, n9685,
    n9686, n9687, n9688, n9689, n9690, n9691,
    n9692, n9693, n9694, n9695, n9696, n9697,
    n9698, n9699, n9700, n9701, n9702, n9703,
    n9704, n9705, n9706, n9707, n9708, n9709,
    n9710, n9711, n9712, n9713, n9714, n9715,
    n9716, n9717, n9718, n9719, n9720, n9721,
    n9722, n9723, n9724, n9725, n9726, n9727,
    n9728, n9729, n9730, n9731, n9732, n9733,
    n9734, n9735, n9736, n9737, n9738, n9739,
    n9740, n9741, n9742, n9743, n9744, n9745,
    n9746, n9747, n9748, n9749, n9750, n9751,
    n9752, n9753, n9754, n9755, n9756, n9757,
    n9758, n9759, n9760, n9761, n9762, n9763,
    n9764, n9765, n9766, n9767, n9768, n9769,
    n9770, n9771, n9772, n9773, n9774, n9775,
    n9776, n9777, n9778, n9779, n9780, n9781,
    n9782, n9783, n9784, n9785, n9786, n9787,
    n9788, n9789, n9790, n9791, n9792, n9793,
    n9794, n9795, n9796, n9797, n9798, n9799,
    n9800, n9801, n9802, n9803, n9804, n9805,
    n9806, n9807, n9808, n9809, n9810, n9811,
    n9812, n9813, n9814, n9815, n9816, n9817,
    n9818, n9819, n9820, n9821, n9822, n9823,
    n9824, n9825, n9826, n9827, n9828, n9829,
    n9830, n9831, n9832, n9833, n9834, n9835,
    n9836, n9837, n9838, n9839, n9840, n9841,
    n9842, n9843, n9844, n9845, n9846, n9847,
    n9848, n9849, n9850, n9851, n9852, n9853,
    n9854, n9855, n9856, n9857, n9858, n9859,
    n9860, n9861, n9862, n9863, n9864, n9865,
    n9866, n9867, n9868, n9869, n9870, n9871,
    n9872, n9873, n9874, n9875, n9876, n9877,
    n9878, n9879, n9880, n9881, n9882, n9883,
    n9884, n9885, n9886, n9887, n9888, n9889,
    n9890, n9891, n9892, n9893, n9894, n9895,
    n9896, n9897, n9898, n9899, n9900, n9901,
    n9902, n9903, n9904, n9905, n9906, n9907,
    n9908, n9909, n9910, n9911, n9912, n9913,
    n9914, n9915, n9916, n9917, n9918, n9919,
    n9920, n9921, n9922, n9923, n9924, n9925,
    n9926, n9927, n9928, n9929, n9930, n9931,
    n9932, n9933, n9934, n9935, n9936, n9937,
    n9938, n9939, n9940, n9941, n9942, n9943,
    n9944, n9945, n9946, n9947, n9948, n9949,
    n9950, n9951, n9952, n9953, n9954, n9955,
    n9956, n9957, n9958, n9959, n9960, n9961,
    n9962, n9963, n9964, n9965, n9966, n9967,
    n9968, n9969, n9970, n9971, n9972, n9973,
    n9974, n9975, n9976, n9977, n9978, n9979,
    n9980, n9981, n9982, n9983, n9984, n9985,
    n9986, n9987, n9988, n9989, n9990, n9991,
    n9992, n9993, n9994, n9995, n9996, n9997,
    n9998, n9999, n10000, n10001, n10002, n10003,
    n10004, n10005, n10006, n10007, n10008, n10009,
    n10010, n10011, n10012, n10013, n10014, n10015,
    n10016, n10017, n10018, n10019, n10020, n10021,
    n10022, n10023, n10024, n10025, n10026, n10027,
    n10028, n10029, n10030, n10031, n10032, n10033,
    n10034, n10035, n10036, n10037, n10038, n10039,
    n10040, n10041, n10042, n10043, n10044, n10045,
    n10046, n10047, n10048, n10049, n10050, n10051,
    n10052, n10053, n10054, n10055, n10056, n10057,
    n10058, n10059, n10060, n10061, n10062, n10063,
    n10064, n10065, n10066, n10067, n10068, n10069,
    n10070, n10071, n10072, n10073, n10074, n10075,
    n10076, n10077, n10078, n10079, n10080, n10081,
    n10082, n10083, n10084, n10085, n10086, n10087,
    n10088, n10089, n10090, n10091, n10092, n10093,
    n10094, n10095, n10096, n10097, n10098, n10099,
    n10100, n10101, n10102, n10103, n10104, n10105,
    n10106, n10107, n10108, n10109, n10110, n10111,
    n10112, n10113, n10114, n10115, n10116, n10117,
    n10118, n10119, n10120, n10121, n10122, n10123,
    n10124, n10125, n10126, n10127, n10128, n10129,
    n10130, n10131, n10132, n10133, n10134, n10135,
    n10136, n10137, n10138, n10139, n10140, n10141,
    n10142, n10143, n10144, n10145, n10146, n10147,
    n10148, n10149, n10150, n10151, n10152, n10153,
    n10154, n10155, n10156, n10157, n10158, n10159,
    n10160, n10161, n10162, n10163, n10164, n10165,
    n10166, n10167, n10168, n10169, n10170, n10171,
    n10172, n10173, n10174, n10175, n10176, n10177,
    n10178, n10179, n10180, n10181, n10182, n10183,
    n10184, n10185, n10186, n10187, n10188, n10189,
    n10190, n10191, n10192, n10193, n10194, n10195,
    n10196, n10197, n10198, n10199, n10200, n10201,
    n10202, n10203, n10204, n10205, n10206, n10207,
    n10208, n10209, n10210, n10211, n10212, n10213,
    n10214, n10215, n10216, n10217, n10218, n10219,
    n10220, n10221, n10222, n10223, n10224, n10225,
    n10226, n10227, n10228, n10229, n10230, n10231,
    n10232, n10233, n10234, n10235, n10236, n10237,
    n10238, n10239, n10240, n10241, n10242, n10243,
    n10244, n10245, n10246, n10247, n10248, n10249,
    n10250, n10251, n10252, n10253, n10254, n10255,
    n10256, n10257, n10258, n10259, n10260, n10261,
    n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10269, n10270, n10271, n10272, n10273,
    n10274, n10275, n10276, n10277, n10278, n10279,
    n10280, n10281, n10282, n10283, n10284, n10285,
    n10286, n10287, n10288, n10289, n10290, n10291,
    n10292, n10293, n10294, n10295, n10296, n10297,
    n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309,
    n10310, n10311, n10312, n10313, n10314, n10315,
    n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327,
    n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345,
    n10346, n10347, n10348, n10349, n10350, n10351,
    n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363,
    n10364, n10365, n10366, n10367, n10368, n10369,
    n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381,
    n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10395, n10396, n10397, n10398, n10399,
    n10400, n10401, n10402, n10403, n10404, n10405,
    n10406, n10407, n10408, n10409, n10410, n10411,
    n10412, n10413, n10414, n10415, n10416, n10417,
    n10418, n10419, n10420, n10421, n10422, n10423,
    n10424, n10425, n10426, n10427, n10428, n10429,
    n10430, n10431, n10432, n10433, n10434, n10435,
    n10436, n10437, n10438, n10439, n10440, n10441,
    n10442, n10443, n10444, n10445, n10446, n10447,
    n10448, n10449, n10450, n10451, n10452, n10453,
    n10454, n10455, n10456, n10457, n10458, n10459,
    n10460, n10461, n10462, n10463, n10464, n10465,
    n10466, n10467, n10468, n10469, n10470, n10471,
    n10472, n10473, n10474, n10475, n10476, n10477,
    n10478, n10479, n10480, n10481, n10482, n10483,
    n10484, n10485, n10486, n10487, n10488, n10489,
    n10490, n10491, n10492, n10493, n10494, n10495,
    n10496, n10497, n10498, n10499, n10500, n10501,
    n10502, n10503, n10504, n10505, n10506, n10507,
    n10508, n10509, n10510, n10511, n10512, n10513,
    n10514, n10515, n10516, n10517, n10518, n10519,
    n10520, n10521, n10522, n10523, n10524, n10525,
    n10526, n10527, n10528, n10529, n10530, n10531,
    n10532, n10533, n10534, n10535, n10536, n10537,
    n10538, n10539, n10540, n10541, n10542, n10543,
    n10544, n10545, n10546, n10547, n10548, n10549,
    n10550, n10551, n10552, n10553, n10554, n10555,
    n10556, n10557, n10558, n10559, n10560, n10561,
    n10562, n10563, n10564, n10565, n10566, n10567,
    n10568, n10569, n10570, n10571, n10572, n10573,
    n10574, n10575, n10576, n10577, n10578, n10579,
    n10580, n10581, n10582, n10583, n10584, n10585,
    n10586, n10587, n10588, n10589, n10590, n10591,
    n10592, n10593, n10594, n10595, n10596, n10597,
    n10598, n10599, n10600, n10601, n10602, n10603,
    n10604, n10605, n10606, n10607, n10608, n10609,
    n10610, n10611, n10612, n10613, n10614, n10615,
    n10616, n10617, n10618, n10619, n10620, n10621,
    n10622, n10623, n10624, n10625, n10626, n10627,
    n10628, n10629, n10630, n10631, n10632, n10633,
    n10634, n10635, n10636, n10637, n10638, n10639,
    n10640, n10641, n10642, n10643, n10644, n10645,
    n10646, n10647, n10648, n10649, n10650, n10651,
    n10652, n10653, n10654, n10655, n10656, n10657,
    n10658, n10659, n10660, n10661, n10662, n10663,
    n10664, n10665, n10666, n10667, n10668, n10669,
    n10670, n10671, n10672, n10673, n10674, n10675,
    n10676, n10677, n10678, n10679, n10680, n10681,
    n10682, n10683, n10684, n10685, n10686, n10687,
    n10688, n10689, n10690, n10691, n10692, n10693,
    n10694, n10695, n10696, n10697, n10698, n10699,
    n10700, n10701, n10702, n10703, n10704, n10705,
    n10706, n10707, n10708, n10709, n10710, n10711,
    n10712, n10713, n10714, n10715, n10716, n10717,
    n10718, n10719, n10720, n10721, n10722, n10723,
    n10724, n10725, n10726, n10727, n10728, n10729,
    n10730, n10731, n10732, n10733, n10734, n10735,
    n10736, n10737, n10738, n10739, n10740, n10741,
    n10742, n10743, n10744, n10745, n10746, n10747,
    n10748, n10749, n10750, n10751, n10752, n10753,
    n10754, n10755, n10756, n10757, n10758, n10759,
    n10760, n10761, n10762, n10763, n10764, n10765,
    n10766, n10767, n10768, n10769, n10770, n10771,
    n10772, n10773, n10774, n10775, n10776, n10777,
    n10778, n10779, n10780, n10781, n10782, n10783,
    n10784, n10785, n10786, n10787, n10788, n10789,
    n10790, n10791, n10792, n10793, n10794, n10795,
    n10796, n10797, n10798, n10799, n10800, n10801,
    n10802, n10803, n10804, n10805, n10806, n10807,
    n10808, n10809, n10810, n10811, n10812, n10813,
    n10814, n10815, n10816, n10817, n10818, n10819,
    n10820, n10821, n10822, n10823, n10824, n10825,
    n10826, n10827, n10828, n10829, n10830, n10831,
    n10832, n10833, n10834, n10835, n10836, n10837,
    n10838, n10839, n10840, n10841, n10842, n10843,
    n10844, n10845, n10846, n10847, n10848, n10849,
    n10850, n10851, n10852, n10853, n10854, n10855,
    n10856, n10857, n10858, n10859, n10860, n10861,
    n10862, n10863, n10864, n10865, n10866, n10867,
    n10868, n10869, n10870, n10871, n10872, n10873,
    n10874, n10875, n10876, n10877, n10878, n10879,
    n10880, n10881, n10882, n10883, n10884, n10885,
    n10886, n10887, n10888, n10889, n10890, n10891,
    n10892, n10893, n10894, n10895, n10896, n10897,
    n10898, n10899, n10900, n10901, n10902, n10903,
    n10904, n10905, n10906, n10907, n10908, n10909,
    n10910, n10911, n10912, n10913, n10914, n10915,
    n10916, n10917, n10918, n10919, n10920, n10921,
    n10922, n10923, n10924, n10925, n10926, n10927,
    n10928, n10929, n10930, n10931, n10932, n10933,
    n10934, n10935, n10936, n10937, n10938, n10939,
    n10940, n10941, n10942, n10943, n10944, n10945,
    n10946, n10947, n10948, n10949, n10950, n10951,
    n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10961, n10962, n10963,
    n10964, n10965, n10966, n10967, n10968, n10969,
    n10970, n10971, n10972, n10973, n10974, n10975,
    n10976, n10977, n10978, n10979, n10980, n10981,
    n10982, n10983, n10984, n10985, n10986, n10987,
    n10988, n10989, n10990, n10991, n10992, n10993,
    n10994, n10995, n10996, n10997, n10998, n10999,
    n11000, n11001, n11002, n11003, n11004, n11005,
    n11006, n11007, n11008, n11009, n11010, n11011,
    n11012, n11013, n11014, n11015, n11016, n11017,
    n11018, n11019, n11020, n11021, n11022, n11023,
    n11024, n11025, n11026, n11027, n11028, n11029,
    n11030, n11031, n11032, n11033, n11034, n11035,
    n11036, n11037, n11038, n11039, n11040, n11041,
    n11042, n11043, n11044, n11045, n11046, n11047,
    n11048, n11049, n11050, n11051, n11052, n11053,
    n11054, n11055, n11056, n11057, n11058, n11059,
    n11060, n11061, n11062, n11063, n11064, n11065,
    n11066, n11067, n11068, n11069, n11070, n11071,
    n11072, n11073, n11074, n11075, n11076, n11077,
    n11078, n11079, n11080, n11081, n11082, n11083,
    n11084, n11085, n11086, n11087, n11088, n11089,
    n11090, n11091, n11092, n11093, n11094, n11095,
    n11096, n11097, n11098, n11099, n11100, n11101,
    n11102, n11103, n11104, n11105, n11106, n11107,
    n11108, n11109, n11110, n11111, n11112, n11113,
    n11114, n11115, n11116, n11117, n11118, n11119,
    n11120, n11121, n11122, n11123, n11124, n11125,
    n11126, n11127, n11128, n11129, n11130, n11131,
    n11132, n11133, n11134, n11135, n11136, n11137,
    n11138, n11139, n11140, n11141, n11142, n11143,
    n11144, n11145, n11146, n11147, n11148, n11149,
    n11150, n11151, n11152, n11153, n11154, n11155,
    n11156, n11157, n11158, n11159, n11160, n11161,
    n11162, n11163, n11164, n11165, n11166, n11167,
    n11168, n11169, n11170, n11171, n11172, n11173,
    n11174, n11175, n11176, n11177, n11178, n11179,
    n11180, n11181, n11182, n11183, n11184, n11185,
    n11186, n11187, n11188, n11189, n11190, n11191,
    n11192, n11193, n11194, n11195, n11196, n11197,
    n11198, n11199, n11200, n11201, n11202, n11203,
    n11204, n11205, n11206, n11207, n11208, n11209,
    n11210, n11211, n11212, n11213, n11214, n11215,
    n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227,
    n11228, n11229, n11230, n11231, n11232, n11233,
    n11234, n11235, n11236, n11237, n11238, n11239,
    n11240, n11241, n11242, n11243, n11244, n11245,
    n11246, n11247, n11248, n11249, n11250, n11251,
    n11252, n11253, n11254, n11255, n11256, n11257,
    n11258, n11259, n11260, n11261, n11262, n11263,
    n11264, n11265, n11266, n11267, n11268, n11269,
    n11270, n11271, n11272, n11273, n11274, n11275,
    n11276, n11277, n11278, n11279, n11280, n11281,
    n11282, n11283, n11284, n11285, n11286, n11287,
    n11288, n11289, n11290, n11291, n11292, n11293,
    n11294, n11295, n11296, n11297, n11298, n11299,
    n11300, n11301, n11302, n11303, n11304, n11305,
    n11306, n11307, n11308, n11309, n11310, n11311,
    n11312, n11313, n11314, n11315, n11316, n11317,
    n11318, n11319, n11320, n11321, n11322, n11323,
    n11324, n11325, n11326, n11327, n11328, n11329,
    n11330, n11331, n11332, n11333, n11334, n11335,
    n11336, n11337, n11338, n11339, n11340, n11341,
    n11342, n11343, n11344, n11345, n11346, n11347,
    n11348, n11349, n11350, n11351, n11352, n11353,
    n11354, n11355, n11356, n11357, n11358, n11359,
    n11360, n11361, n11362, n11363, n11364, n11365,
    n11366, n11367, n11368, n11369, n11370, n11371,
    n11372, n11373, n11374, n11375, n11376, n11377,
    n11378, n11379, n11380, n11381, n11382, n11383,
    n11384, n11385, n11386, n11387, n11388, n11389,
    n11390, n11391, n11392, n11393, n11394, n11395,
    n11396, n11397, n11398, n11399, n11400, n11401,
    n11402, n11403, n11404, n11405, n11406, n11407,
    n11408, n11409, n11410, n11411, n11412, n11413,
    n11414, n11415, n11416, n11417, n11418, n11419,
    n11420, n11421, n11422, n11423, n11424, n11425,
    n11426, n11427, n11428, n11429, n11430, n11431,
    n11432, n11433, n11434, n11435, n11436, n11437,
    n11438, n11439, n11440, n11441, n11442, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449,
    n11450, n11451, n11452, n11453, n11454, n11455,
    n11456, n11457, n11458, n11459, n11460, n11461,
    n11462, n11463, n11464, n11465, n11466, n11467,
    n11468, n11469, n11470, n11471, n11472, n11473,
    n11474, n11475, n11476, n11477, n11478, n11479,
    n11480, n11481, n11482, n11483, n11484, n11485,
    n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497,
    n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509,
    n11510, n11511, n11512, n11513, n11514, n11515,
    n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527,
    n11528, n11529, n11530, n11531, n11532, n11533,
    n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545,
    n11546, n11547, n11548, n11549, n11550, n11551,
    n11552, n11553, n11554, n11555, n11556, n11557,
    n11558, n11559, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569,
    n11570, n11571, n11572, n11573, n11574, n11575,
    n11576, n11577, n11578, n11579, n11580, n11581,
    n11582, n11583, n11584, n11585, n11586, n11587,
    n11588, n11589, n11590, n11591, n11592, n11593,
    n11594, n11595, n11596, n11597, n11598, n11599,
    n11600, n11601, n11602, n11603, n11604, n11605,
    n11606, n11607, n11608, n11609, n11610, n11611,
    n11612, n11613, n11614, n11615, n11616, n11617,
    n11618, n11619, n11620, n11621, n11622, n11623,
    n11624, n11625, n11626, n11627, n11628, n11629,
    n11630, n11631, n11632, n11633, n11634, n11635,
    n11636, n11637, n11638, n11639, n11640, n11641,
    n11642, n11643, n11644, n11645, n11646, n11647,
    n11648, n11649, n11650, n11651, n11652, n11653,
    n11654, n11655, n11656, n11657, n11658, n11659,
    n11660, n11661, n11662, n11663, n11664, n11665,
    n11666, n11667, n11668, n11669, n11670, n11671,
    n11672, n11673, n11674, n11675, n11676, n11677,
    n11678, n11679, n11680, n11681, n11682, n11683,
    n11684, n11685, n11686, n11687, n11688, n11689,
    n11690, n11691, n11692, n11693, n11694, n11695,
    n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11704, n11705, n11706, n11707,
    n11708, n11709, n11710, n11711, n11712, n11713,
    n11714, n11715, n11716, n11717, n11718, n11719,
    n11720, n11721, n11722, n11723, n11724, n11725,
    n11726, n11727, n11728, n11729, n11730, n11731,
    n11732, n11733, n11734, n11735, n11736, n11737,
    n11738, n11739, n11740, n11741, n11742, n11743,
    n11744, n11745, n11746, n11747, n11748, n11749,
    n11750, n11751, n11752, n11753, n11754, n11755,
    n11756, n11757, n11758, n11759, n11760, n11761,
    n11762, n11763, n11764, n11765, n11766, n11767,
    n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779,
    n11780, n11781, n11782, n11783, n11784, n11785,
    n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797,
    n11798, n11799, n11800, n11801, n11802, n11803,
    n11804, n11805, n11806, n11807, n11808, n11809,
    n11810, n11811, n11812, n11813, n11814, n11815,
    n11816, n11817, n11818, n11819, n11820, n11821,
    n11822, n11823, n11824, n11825, n11826, n11827,
    n11828, n11829, n11830, n11831, n11832, n11833,
    n11834, n11835, n11836, n11837, n11838, n11839,
    n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11849, n11850, n11851,
    n11852, n11853, n11854, n11855, n11856, n11857,
    n11858, n11859, n11860, n11861, n11862, n11863,
    n11864, n11865, n11866, n11867, n11868, n11869,
    n11870, n11871, n11872, n11873, n11874, n11875,
    n11876, n11877, n11878, n11879, n11880, n11881,
    n11882, n11883, n11884, n11885, n11886, n11887,
    n11888, n11889, n11890, n11891, n11892, n11893,
    n11894, n11895, n11896, n11897, n11898, n11899,
    n11900, n11901, n11902, n11903, n11904, n11905,
    n11906, n11907, n11908, n11909, n11910, n11911,
    n11912, n11913, n11914, n11915, n11916, n11917,
    n11918, n11919, n11920, n11921, n11922, n11923,
    n11924, n11925, n11926, n11927, n11928, n11929,
    n11930, n11931, n11932, n11933, n11934, n11935,
    n11936, n11937, n11938, n11939, n11940, n11941,
    n11942, n11943, n11944, n11945, n11946, n11947,
    n11948, n11949, n11950, n11951, n11952, n11953,
    n11954, n11955, n11956, n11957, n11958, n11959,
    n11960, n11961, n11962, n11963, n11964, n11965,
    n11966, n11967, n11968, n11969, n11970, n11971,
    n11972, n11973, n11974, n11975, n11976, n11977,
    n11978, n11979, n11980, n11981, n11982, n11983,
    n11984, n11985, n11986, n11987, n11988, n11989,
    n11990, n11991, n11992, n11993, n11994, n11995,
    n11996, n11997, n11998, n11999, n12000, n12001,
    n12002, n12003, n12004, n12005, n12006, n12007,
    n12008, n12009, n12010, n12011, n12012, n12013,
    n12014, n12015, n12016, n12017, n12018, n12019,
    n12020, n12021, n12022, n12023, n12024, n12025,
    n12026, n12027, n12028, n12029, n12030, n12031,
    n12032, n12033, n12034, n12035, n12036, n12037,
    n12038, n12039, n12040, n12041, n12042, n12043,
    n12044, n12045, n12046, n12047, n12048, n12049,
    n12050, n12051, n12052, n12053, n12054, n12055,
    n12056, n12057, n12058, n12059, n12060, n12061,
    n12062, n12063, n12064, n12065, n12066, n12067,
    n12068, n12069, n12070, n12071, n12072, n12073,
    n12074, n12075, n12076, n12077, n12078, n12079,
    n12080, n12081, n12082, n12083, n12084, n12085,
    n12086, n12087, n12088, n12089, n12090, n12091,
    n12092, n12093, n12094, n12095, n12096, n12097,
    n12098, n12099, n12100, n12101, n12102, n12103,
    n12104, n12105, n12106, n12107, n12108, n12109,
    n12110, n12111, n12112, n12113, n12114, n12115,
    n12116, n12117, n12118, n12119, n12120, n12121,
    n12122, n12123, n12124, n12125, n12126, n12127,
    n12128, n12129, n12130, n12131, n12132, n12133,
    n12134, n12135, n12136, n12137, n12138, n12139,
    n12140, n12141, n12142, n12143, n12144, n12145,
    n12146, n12147, n12148, n12149, n12150, n12151,
    n12152, n12153, n12154, n12155, n12156, n12157,
    n12158, n12159, n12160, n12161, n12162, n12163,
    n12164, n12165, n12166, n12167, n12168, n12169,
    n12170, n12171, n12172, n12173, n12174, n12175,
    n12176, n12177, n12178, n12179, n12180, n12181,
    n12182, n12183, n12184, n12185, n12186, n12187,
    n12188, n12189, n12190, n12191, n12192, n12193,
    n12194, n12195, n12196, n12197, n12198, n12199,
    n12200, n12201, n12202, n12203, n12204, n12205,
    n12206, n12207, n12208, n12209, n12210, n12211,
    n12212, n12213, n12214, n12215, n12216, n12217,
    n12218, n12219, n12220, n12221, n12222, n12223,
    n12224, n12225, n12226, n12227, n12228, n12229,
    n12230, n12231, n12232, n12233, n12234, n12235,
    n12236, n12237, n12238, n12239, n12240, n12241,
    n12242, n12243, n12244, n12245, n12246, n12247,
    n12248, n12249, n12250, n12251, n12252, n12253,
    n12254, n12255, n12256, n12257, n12258, n12259,
    n12260, n12261, n12262, n12263, n12264, n12265,
    n12266, n12267, n12268, n12269, n12270, n12271,
    n12272, n12273, n12274, n12275, n12276, n12277,
    n12278, n12279, n12280, n12281, n12282, n12283,
    n12284, n12285, n12286, n12287, n12288, n12289,
    n12290, n12291, n12292, n12293, n12294, n12295,
    n12296, n12297, n12298, n12299, n12300, n12301,
    n12302, n12303, n12304, n12305, n12306, n12307,
    n12308, n12309, n12310, n12311, n12312, n12313,
    n12314, n12315, n12316, n12317, n12318, n12319,
    n12320, n12321, n12322, n12323, n12324, n12325,
    n12326, n12327, n12328, n12329, n12330, n12331,
    n12332, n12333, n12334, n12335, n12336, n12337,
    n12338, n12339, n12340, n12341, n12342, n12343,
    n12344, n12345, n12346, n12347, n12348, n12349,
    n12350, n12351, n12352, n12353, n12354, n12355,
    n12356, n12357, n12358, n12359, n12360, n12361,
    n12362, n12363, n12364, n12365, n12366, n12367,
    n12368, n12369, n12370, n12371, n12372, n12373,
    n12374, n12375, n12376, n12377, n12378, n12379,
    n12380, n12381, n12382, n12383, n12384, n12385,
    n12386, n12387, n12388, n12389, n12390, n12391,
    n12392, n12393, n12394, n12395, n12396, n12397,
    n12398, n12399, n12400, n12401, n12402, n12403,
    n12404, n12405, n12406, n12407, n12408, n12409,
    n12410, n12411, n12412, n12413, n12414, n12415,
    n12416, n12417, n12418, n12419, n12420, n12421,
    n12422, n12423, n12424, n12425, n12426, n12427,
    n12428, n12429, n12430, n12431, n12432, n12433,
    n12434, n12435, n12436, n12437, n12438, n12439,
    n12440, n12441, n12442, n12443, n12444, n12445,
    n12446, n12447, n12448, n12449, n12450, n12451,
    n12452, n12453, n12454, n12455, n12456, n12457,
    n12458, n12459, n12460, n12461, n12462, n12463,
    n12464, n12465, n12466, n12467, n12468, n12469,
    n12470, n12471, n12472, n12473, n12474, n12475,
    n12476, n12477, n12478, n12479, n12480, n12481,
    n12482, n12483, n12484, n12485, n12486, n12487,
    n12488, n12489, n12490, n12491, n12492, n12493,
    n12494, n12495, n12496, n12497, n12498, n12499,
    n12500, n12501, n12502, n12503, n12504, n12505,
    n12506, n12507, n12508, n12509, n12510, n12511,
    n12512, n12513, n12514, n12515, n12516, n12517,
    n12518, n12519, n12520, n12521, n12522, n12523,
    n12524, n12525, n12526, n12527, n12528, n12529,
    n12530, n12531, n12532, n12533, n12534, n12535,
    n12536, n12537, n12538, n12539, n12540, n12541,
    n12542, n12543, n12544, n12545, n12546, n12547,
    n12548, n12549, n12550, n12551, n12552, n12553,
    n12554, n12555, n12556, n12557, n12558, n12559,
    n12560, n12561, n12562, n12563, n12564, n12565,
    n12566, n12567, n12568, n12569, n12570, n12571,
    n12572, n12573, n12574, n12575, n12576, n12577,
    n12578, n12579, n12580, n12581, n12582, n12583,
    n12584, n12585, n12586, n12587, n12588, n12589,
    n12590, n12591, n12592, n12593, n12594, n12595,
    n12596, n12597, n12598, n12599, n12600, n12601,
    n12602, n12603, n12604, n12605, n12606, n12607,
    n12608, n12609, n12610, n12611, n12612, n12613,
    n12614, n12615, n12616, n12617, n12618, n12619,
    n12620, n12621, n12622, n12623, n12624, n12625,
    n12626, n12627, n12628, n12629, n12630, n12631,
    n12632, n12633, n12634, n12635, n12636, n12637,
    n12638, n12639, n12640, n12641, n12642, n12643,
    n12644, n12645, n12646, n12647, n12648, n12649,
    n12650, n12651, n12652, n12653, n12654, n12655,
    n12656, n12657, n12658, n12659, n12660, n12661,
    n12662, n12663, n12664, n12665, n12666, n12667,
    n12668, n12669, n12670, n12671, n12672, n12673,
    n12674, n12675, n12676, n12677, n12678, n12679,
    n12680, n12681, n12682, n12683, n12684, n12685,
    n12686, n12687, n12688, n12689, n12690, n12691,
    n12692, n12693, n12694, n12695, n12696, n12697,
    n12698, n12699, n12700, n12701, n12702, n12703,
    n12704, n12705, n12706, n12707, n12708, n12709,
    n12710, n12711, n12712, n12713, n12714, n12715,
    n12716, n12717, n12718, n12719, n12720, n12721,
    n12722, n12723, n12724, n12725, n12726, n12727,
    n12728, n12729, n12730, n12731, n12732, n12733,
    n12734, n12735, n12736, n12737, n12738, n12739,
    n12740, n12741, n12742, n12743, n12744, n12745,
    n12746, n12747, n12748, n12749, n12750, n12751,
    n12752, n12753, n12754, n12755, n12756, n12757,
    n12758, n12759, n12760, n12761, n12762, n12763,
    n12764, n12765, n12766, n12767, n12768, n12769,
    n12770, n12771, n12772, n12773, n12774, n12775,
    n12776, n12777, n12778, n12779, n12780, n12781,
    n12782, n12783, n12784, n12785, n12786, n12787,
    n12788, n12789, n12790, n12791, n12792, n12793,
    n12794, n12795, n12796, n12797, n12798, n12799,
    n12800, n12801, n12802, n12803, n12804, n12805,
    n12806, n12807, n12808, n12809, n12810, n12811,
    n12812, n12813, n12814, n12815, n12816, n12817,
    n12818, n12819, n12820, n12821, n12822, n12823,
    n12824, n12825, n12826, n12827, n12828, n12829,
    n12830, n12831, n12832, n12833, n12834, n12835,
    n12836, n12837, n12838, n12839, n12840, n12841,
    n12842, n12843, n12844, n12845, n12846, n12847,
    n12848, n12849, n12850, n12851, n12852, n12853,
    n12854, n12855, n12856, n12857, n12858, n12859,
    n12860, n12861, n12862, n12863, n12864, n12865,
    n12866, n12867, n12868, n12869, n12870, n12871,
    n12872, n12873, n12874, n12875, n12876, n12877,
    n12878, n12879, n12880, n12881, n12882, n12883,
    n12884, n12885, n12886, n12887, n12888, n12889,
    n12890, n12891, n12892, n12893, n12894, n12895,
    n12896, n12897, n12898, n12899, n12900, n12901,
    n12902, n12903, n12904, n12905, n12906, n12907,
    n12908, n12909, n12910, n12911, n12912, n12913,
    n12914, n12915, n12916, n12917, n12918, n12919,
    n12920, n12921, n12922, n12923, n12924, n12925,
    n12926, n12927, n12928, n12929, n12930, n12931,
    n12932, n12933, n12934, n12935, n12936, n12937,
    n12938, n12939, n12940, n12941, n12942, n12943,
    n12944, n12945, n12946, n12947, n12948, n12949,
    n12950, n12951, n12952, n12953, n12954, n12955,
    n12956, n12957, n12958, n12959, n12960, n12961,
    n12962, n12963, n12964, n12965, n12966, n12967,
    n12968, n12969, n12970, n12971, n12972, n12973,
    n12974, n12975, n12976, n12977, n12978, n12979,
    n12980, n12981, n12982, n12983, n12984, n12985,
    n12986, n12987, n12988, n12989, n12990, n12991,
    n12992, n12993, n12994, n12995, n12996, n12997,
    n12998, n12999, n13000, n13001, n13002, n13003,
    n13004, n13005, n13006, n13007, n13008, n13009,
    n13010, n13011, n13012, n13013, n13014, n13015,
    n13016, n13017, n13018, n13019, n13020, n13021,
    n13022, n13023, n13024, n13025, n13026, n13027,
    n13028, n13029, n13030, n13031, n13032, n13033,
    n13034, n13035, n13036, n13037, n13038, n13039,
    n13040, n13041, n13042, n13043, n13044, n13045,
    n13046, n13047, n13048, n13049, n13050, n13051,
    n13052, n13053, n13054, n13055, n13056, n13057,
    n13058, n13059, n13060, n13061, n13062, n13063,
    n13064, n13065, n13066, n13067, n13068, n13069,
    n13070, n13071, n13072, n13073, n13074, n13075,
    n13076, n13077, n13078, n13079, n13080, n13081,
    n13082, n13083, n13084, n13085, n13086, n13087,
    n13088, n13089, n13090, n13091, n13092, n13093,
    n13094, n13095, n13096, n13097, n13098, n13099,
    n13100, n13101, n13102, n13103, n13104, n13105,
    n13106, n13107, n13108, n13109, n13110, n13111,
    n13112, n13113, n13114, n13115, n13116, n13117,
    n13118, n13119, n13120, n13121, n13122, n13123,
    n13124, n13125, n13126, n13127, n13128, n13129,
    n13130, n13131, n13132, n13133, n13134, n13135,
    n13136, n13137, n13138, n13139, n13140, n13141,
    n13142, n13143, n13144, n13145, n13146, n13147,
    n13148, n13149, n13150, n13151, n13152, n13153,
    n13154, n13155, n13156, n13157, n13158, n13159,
    n13160, n13161, n13162, n13163, n13164, n13165,
    n13166, n13167, n13168, n13169, n13170, n13171,
    n13172, n13173, n13174, n13175, n13176, n13177,
    n13178, n13179, n13180, n13181, n13182, n13183,
    n13184, n13185, n13186, n13187, n13188, n13189,
    n13190, n13191, n13192, n13193, n13194, n13195,
    n13196, n13197, n13198, n13199, n13200, n13201,
    n13202, n13203, n13204, n13205, n13206, n13207,
    n13208, n13209, n13210, n13211, n13212, n13213,
    n13214, n13215, n13216, n13217, n13218, n13219,
    n13220, n13221, n13222, n13223, n13224, n13225,
    n13226, n13227, n13228, n13229, n13230, n13231,
    n13232, n13233, n13234, n13235, n13236, n13237,
    n13238, n13239, n13240, n13241, n13242, n13243,
    n13244, n13245, n13246, n13247, n13248, n13249,
    n13250, n13251, n13252, n13253, n13254, n13255,
    n13256, n13257, n13258, n13259, n13260, n13261,
    n13262, n13263, n13264, n13265, n13266, n13267,
    n13268, n13269, n13270, n13271, n13272, n13273,
    n13274, n13275, n13276, n13277, n13278, n13279,
    n13280, n13281, n13282, n13283, n13284, n13285,
    n13286, n13287, n13288, n13289, n13290, n13291,
    n13292, n13293, n13294, n13295, n13296, n13297,
    n13298, n13299, n13300, n13301, n13302, n13303,
    n13304, n13305, n13306, n13307, n13308, n13309,
    n13310, n13311, n13312, n13313, n13314, n13315,
    n13316, n13317, n13318, n13319, n13320, n13321,
    n13322, n13323, n13324, n13325, n13326, n13327,
    n13328, n13329, n13330, n13331, n13332, n13333,
    n13334, n13335, n13336, n13337, n13338, n13339,
    n13340, n13341, n13342, n13343, n13344, n13345,
    n13346, n13347, n13348, n13349, n13350, n13351,
    n13352, n13353, n13354, n13355, n13356, n13357,
    n13358, n13359, n13360, n13361, n13362, n13363,
    n13364, n13365, n13366, n13367, n13368, n13369,
    n13370, n13371, n13372, n13373, n13374, n13375,
    n13376, n13377, n13378, n13379, n13380, n13381,
    n13382, n13383, n13384, n13385, n13386, n13387,
    n13388, n13389, n13390, n13391, n13392, n13393,
    n13394, n13395, n13396, n13397, n13398, n13399,
    n13400, n13401, n13402, n13403, n13404, n13405,
    n13406, n13407, n13408, n13409, n13410, n13411,
    n13412, n13413, n13414, n13415, n13416, n13417,
    n13418, n13419, n13420, n13421, n13422, n13423,
    n13424, n13425, n13426, n13427, n13428, n13429,
    n13430, n13431, n13432, n13433, n13434, n13435,
    n13436, n13437, n13438, n13439, n13440, n13441,
    n13442, n13443, n13444, n13445, n13446, n13447,
    n13448, n13449, n13450, n13451, n13452, n13453,
    n13454, n13455, n13456, n13457, n13458, n13459,
    n13460, n13461, n13462, n13463, n13464, n13465,
    n13466, n13467, n13468, n13469, n13470, n13471,
    n13472, n13473, n13474, n13475, n13476, n13477,
    n13478, n13479, n13480, n13481, n13482, n13483,
    n13484, n13485, n13486, n13487, n13488, n13489,
    n13490, n13491, n13492, n13493, n13494, n13495,
    n13496, n13497, n13498, n13499, n13500, n13501,
    n13502, n13503, n13504, n13505, n13506, n13507,
    n13508, n13509, n13510, n13511, n13512, n13513,
    n13514, n13515, n13516, n13517, n13518, n13519,
    n13520, n13521, n13522, n13523, n13524, n13525,
    n13526, n13527, n13528, n13529, n13530, n13531,
    n13532, n13533, n13534, n13535, n13536, n13537,
    n13538, n13539, n13540, n13541, n13542, n13543,
    n13544, n13545, n13546, n13547, n13548, n13549,
    n13550, n13551, n13552, n13553, n13554, n13555,
    n13556, n13557, n13558, n13559, n13560, n13561,
    n13562, n13563, n13564, n13565, n13566, n13567,
    n13568, n13569, n13570, n13571, n13572, n13573,
    n13574, n13575, n13576, n13577, n13578, n13579,
    n13580, n13581, n13582, n13583, n13584, n13585,
    n13586, n13587, n13588, n13589, n13590, n13591,
    n13592, n13593, n13594, n13595, n13596, n13597,
    n13598, n13599, n13600, n13601, n13602, n13603,
    n13604, n13605, n13606, n13607, n13608, n13609,
    n13610, n13611, n13612, n13613, n13614, n13615,
    n13616, n13617, n13618, n13619, n13620, n13621,
    n13622, n13623, n13624, n13625, n13626, n13627,
    n13628, n13629, n13630, n13631, n13632, n13633,
    n13634, n13635, n13636, n13637, n13638, n13639,
    n13640, n13641, n13642, n13643, n13644, n13645,
    n13646, n13647, n13648, n13649, n13650, n13651,
    n13652, n13653, n13654, n13655, n13656, n13657,
    n13658, n13659, n13660, n13661, n13662, n13663,
    n13664, n13665, n13666, n13667, n13668, n13669,
    n13670, n13671, n13672, n13673, n13674, n13675,
    n13676, n13677, n13678, n13679, n13680, n13681,
    n13682, n13683, n13684, n13685, n13686, n13687,
    n13688, n13689, n13690, n13691, n13692, n13693,
    n13694, n13695, n13696, n13697, n13698, n13699,
    n13700, n13701, n13702, n13703, n13704, n13705,
    n13706, n13707, n13708, n13709, n13710, n13711,
    n13712, n13713, n13714, n13715, n13716, n13717,
    n13718, n13719, n13720, n13721, n13722, n13723,
    n13724, n13725, n13726, n13727, n13728, n13729,
    n13730, n13731, n13732, n13733, n13734, n13735,
    n13736, n13737, n13738, n13739, n13740, n13741,
    n13742, n13743, n13744, n13745, n13746, n13747,
    n13748, n13749, n13750, n13751, n13752, n13753,
    n13754, n13755, n13756, n13757, n13758, n13759,
    n13760, n13761, n13762, n13763, n13764, n13765,
    n13766, n13767, n13768, n13769, n13770, n13771,
    n13772, n13773, n13774, n13775, n13776, n13777,
    n13778, n13779, n13780, n13781, n13782, n13783,
    n13784, n13785, n13786, n13787, n13788, n13789,
    n13790, n13791, n13792, n13793, n13794, n13795,
    n13796, n13797, n13798, n13799, n13800, n13801,
    n13802, n13803, n13804, n13805, n13806, n13807,
    n13808, n13809, n13810, n13811, n13812, n13813,
    n13814, n13815, n13816, n13817, n13818, n13819,
    n13820, n13821, n13822, n13823, n13824, n13825,
    n13826, n13827, n13828, n13829, n13830, n13831,
    n13832, n13833, n13834, n13835, n13836, n13837,
    n13838, n13839, n13840, n13841, n13842, n13843,
    n13844, n13845, n13846, n13847, n13848, n13849,
    n13850, n13851, n13852, n13853, n13854, n13855,
    n13856, n13857, n13858, n13859, n13860, n13861,
    n13862, n13863, n13864, n13865, n13866, n13867,
    n13868, n13869, n13870, n13871, n13872, n13873,
    n13874, n13875, n13876, n13877, n13878, n13879,
    n13880, n13881, n13882, n13883, n13884, n13885,
    n13886, n13887, n13888, n13889, n13890, n13891,
    n13892, n13893, n13894, n13895, n13896, n13897,
    n13898, n13899, n13900, n13901, n13902, n13903,
    n13904, n13905, n13906, n13907, n13908, n13909,
    n13910, n13911, n13912, n13913, n13914, n13915,
    n13916, n13917, n13918, n13919, n13920, n13921,
    n13922, n13923, n13924, n13925, n13926, n13927,
    n13928, n13929, n13930, n13931, n13932, n13933,
    n13934, n13935, n13936, n13937, n13938, n13939,
    n13940, n13941, n13942, n13943, n13944, n13945,
    n13946, n13947, n13948, n13949, n13950, n13951,
    n13952, n13953, n13954, n13955, n13956, n13957,
    n13958, n13959, n13960, n13961, n13962, n13963,
    n13964, n13965, n13966, n13967, n13968, n13969,
    n13970, n13971, n13972, n13973, n13974, n13975,
    n13976, n13977, n13978, n13979, n13980, n13981,
    n13982, n13983, n13984, n13985, n13986, n13987,
    n13988, n13989, n13990, n13991, n13992, n13993,
    n13994, n13995, n13996, n13997, n13998, n13999,
    n14000, n14001, n14002, n14003, n14004, n14005,
    n14006, n14007, n14008, n14009, n14010, n14011,
    n14012, n14013, n14014, n14015, n14016, n14017,
    n14018, n14019, n14020, n14021, n14022, n14023,
    n14024, n14025, n14026, n14027, n14028, n14029,
    n14030, n14031, n14032, n14033, n14034, n14035,
    n14036, n14037, n14038, n14039, n14040, n14041,
    n14042, n14043, n14044, n14045, n14046, n14047,
    n14048, n14049, n14050, n14051, n14052, n14053,
    n14054, n14055, n14056, n14057, n14058, n14059,
    n14060, n14061, n14062, n14063, n14064, n14065,
    n14066, n14067, n14068, n14069, n14070, n14071,
    n14072, n14073, n14074, n14075, n14076, n14077,
    n14078, n14079, n14080, n14081, n14082, n14083,
    n14084, n14085, n14086, n14087, n14088, n14089,
    n14090, n14091, n14092, n14093, n14094, n14095,
    n14096, n14097, n14098, n14099, n14100, n14101,
    n14102, n14103, n14104, n14105, n14106, n14107,
    n14108, n14109, n14110, n14111, n14112, n14113,
    n14114, n14115, n14116, n14117, n14118, n14119,
    n14120, n14121, n14122, n14123, n14124, n14125,
    n14126, n14127, n14128, n14129, n14130, n14131,
    n14132, n14133, n14134, n14135, n14136, n14137,
    n14138, n14139, n14140, n14141, n14142, n14143,
    n14144, n14145, n14146, n14147, n14148, n14149,
    n14150, n14151, n14152, n14153, n14154, n14155,
    n14156, n14157, n14158, n14159, n14160, n14161,
    n14162, n14163, n14164, n14165, n14166, n14167,
    n14168, n14169, n14170, n14171, n14172, n14173,
    n14174, n14175, n14176, n14177, n14178, n14179,
    n14180, n14181, n14182, n14183, n14184, n14185,
    n14186, n14187, n14188, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197,
    n14198, n14199, n14200, n14201, n14202, n14203,
    n14204, n14205, n14206, n14207, n14208, n14209,
    n14210, n14211, n14212, n14213, n14214, n14215,
    n14216, n14217, n14218, n14219, n14220, n14221,
    n14222, n14223, n14224, n14225, n14226, n14227,
    n14228, n14229, n14230, n14231, n14232, n14233,
    n14234, n14235, n14236, n14237, n14238, n14239,
    n14240, n14241, n14242, n14243, n14244, n14245,
    n14246, n14247, n14248, n14249, n14250, n14251,
    n14252, n14253, n14254, n14255, n14256, n14257,
    n14258, n14259, n14260, n14261, n14262, n14263,
    n14264, n14265, n14266, n14267, n14268, n14269,
    n14270, n14271, n14272, n14273, n14274, n14275,
    n14276, n14277, n14278, n14279, n14280, n14281,
    n14282, n14283, n14284, n14285, n14286, n14287,
    n14288, n14289, n14290, n14291, n14292, n14293,
    n14294, n14295, n14296, n14297, n14298, n14299,
    n14300, n14301, n14302, n14303, n14304, n14305,
    n14306, n14307, n14308, n14309, n14310, n14311,
    n14312, n14313, n14314, n14315, n14316, n14317,
    n14318, n14319, n14320, n14321, n14322, n14323,
    n14324, n14325, n14326, n14327, n14328, n14329,
    n14330, n14331, n14332, n14333, n14334, n14335,
    n14336, n14337, n14338, n14339, n14340, n14341,
    n14342, n14343, n14344, n14345, n14346, n14347,
    n14348, n14349, n14350, n14351, n14352, n14353,
    n14354, n14355, n14356, n14357, n14358, n14359,
    n14360, n14361, n14362, n14363, n14364, n14365,
    n14366, n14367, n14368, n14369, n14370, n14371,
    n14372, n14373, n14374, n14375, n14376, n14377,
    n14378, n14379, n14380, n14381, n14382, n14383,
    n14384, n14385, n14386, n14387, n14388, n14389,
    n14390, n14391, n14392, n14393, n14394, n14395,
    n14396, n14397, n14398, n14399, n14400, n14401,
    n14402, n14403, n14404, n14405, n14406, n14407,
    n14408, n14409, n14410, n14411, n14412, n14413,
    n14414, n14415, n14416, n14417, n14418, n14419,
    n14420, n14421, n14422, n14423, n14424, n14425,
    n14426, n14427, n14428, n14429, n14430, n14431,
    n14432, n14433, n14434, n14435, n14436, n14437,
    n14438, n14439, n14440, n14441, n14442, n14443,
    n14444, n14445, n14446, n14447, n14448, n14449,
    n14450, n14451, n14452, n14453, n14454, n14455,
    n14456, n14457, n14458, n14459, n14460, n14461,
    n14462, n14463, n14464, n14465, n14466, n14467,
    n14468, n14469, n14470, n14471, n14472, n14473,
    n14474, n14475, n14476, n14477, n14478, n14479,
    n14480, n14481, n14482, n14483, n14484, n14485,
    n14486, n14487, n14488, n14489, n14490, n14491,
    n14492, n14493, n14494, n14495, n14496, n14497,
    n14498, n14499, n14500, n14501, n14502, n14503,
    n14504, n14505, n14506, n14507, n14508, n14509,
    n14510, n14511, n14512, n14513, n14514, n14515,
    n14516, n14517, n14518, n14519, n14520, n14521,
    n14522, n14523, n14524, n14525, n14526, n14527,
    n14528, n14529, n14530, n14531, n14532, n14533,
    n14534, n14535, n14536, n14537, n14538, n14539,
    n14540, n14541, n14542, n14543, n14544, n14545,
    n14546, n14547, n14548, n14549, n14550, n14551,
    n14552, n14553, n14554, n14555, n14556, n14557,
    n14558, n14559, n14560, n14561, n14562, n14563,
    n14564, n14565, n14566, n14567, n14568, n14569,
    n14570, n14571, n14572, n14573, n14574, n14575,
    n14576, n14577, n14578, n14579, n14580, n14581,
    n14582, n14583, n14584, n14585, n14586, n14587,
    n14588, n14589, n14590, n14591, n14592, n14593,
    n14594, n14595, n14596, n14597, n14598, n14599,
    n14600, n14601, n14602, n14603, n14604, n14605,
    n14606, n14607, n14608, n14609, n14610, n14611,
    n14612, n14613, n14614, n14615, n14616, n14617,
    n14618, n14619, n14620, n14621, n14622, n14623,
    n14624, n14625, n14626, n14627, n14628, n14629,
    n14630, n14631, n14632, n14633, n14634, n14635,
    n14636, n14637, n14638, n14639, n14640, n14641,
    n14642, n14643, n14644, n14645, n14646, n14647,
    n14648, n14649, n14650, n14651, n14652, n14653,
    n14654, n14655, n14656, n14657, n14658, n14659,
    n14660, n14661, n14662, n14663, n14664, n14665,
    n14666, n14667, n14668, n14669, n14670, n14671,
    n14672, n14673, n14674, n14675, n14676, n14677,
    n14678, n14679, n14680, n14681, n14682, n14683,
    n14684, n14685, n14686, n14687, n14688, n14689,
    n14690, n14691, n14692, n14693, n14694, n14695,
    n14696, n14697, n14698, n14699, n14700, n14701,
    n14702, n14703, n14704, n14705, n14706, n14707,
    n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14715, n14716, n14717, n14718, n14719,
    n14720, n14721, n14722, n14723, n14724, n14725,
    n14726, n14727, n14728, n14729, n14730, n14731,
    n14732, n14733, n14734, n14735, n14736, n14737,
    n14738, n14739, n14740, n14741, n14742, n14743,
    n14744, n14745, n14746, n14747, n14748, n14749,
    n14750, n14751, n14752, n14753, n14754, n14755,
    n14756, n14757, n14758, n14759, n14760, n14761,
    n14762, n14763, n14764, n14765, n14766, n14767,
    n14768, n14769, n14770, n14771, n14772, n14773,
    n14774, n14775, n14776, n14777, n14778, n14779,
    n14780, n14781, n14782, n14783, n14784, n14785,
    n14786, n14787, n14788, n14789, n14790, n14791,
    n14792, n14793, n14794, n14795, n14796, n14797,
    n14798, n14799, n14800, n14801, n14802, n14803,
    n14804, n14805, n14806, n14807, n14808, n14809,
    n14810, n14811, n14812, n14813, n14814, n14815,
    n14816, n14817, n14818, n14819, n14820, n14821,
    n14822, n14823, n14824, n14825, n14826, n14827,
    n14828, n14829, n14830, n14831, n14832, n14833,
    n14834, n14835, n14836, n14837, n14838, n14839,
    n14840, n14841, n14842, n14843, n14844, n14845,
    n14846, n14847, n14848, n14849, n14850, n14851,
    n14852, n14853, n14854, n14855, n14856, n14857,
    n14858, n14859, n14860, n14861, n14862, n14863,
    n14864, n14865, n14866, n14867, n14868, n14869,
    n14870, n14871, n14872, n14873, n14874, n14875,
    n14876, n14877, n14878, n14879, n14880, n14881,
    n14882, n14883, n14884, n14885, n14886, n14887,
    n14888, n14889, n14890, n14891, n14892, n14893,
    n14894, n14895, n14896, n14897, n14898, n14899,
    n14900, n14901, n14902, n14903, n14904, n14905,
    n14906, n14907, n14908, n14909, n14910, n14911,
    n14912, n14913, n14914, n14915, n14916, n14917,
    n14918, n14919, n14920, n14921, n14922, n14923,
    n14924, n14925, n14926, n14927, n14928, n14929,
    n14930, n14931, n14932, n14933, n14934, n14935,
    n14936, n14937, n14938, n14939, n14940, n14941,
    n14942, n14943, n14944, n14945, n14946, n14947,
    n14948, n14949, n14950, n14951, n14952, n14953,
    n14954, n14955, n14956, n14957, n14958, n14959,
    n14960, n14961, n14962, n14963, n14964, n14965,
    n14966, n14967, n14968, n14969, n14970, n14971,
    n14972, n14973, n14974, n14975, n14976, n14977,
    n14978, n14979, n14980, n14981, n14982, n14983,
    n14984, n14985, n14986, n14987, n14988, n14989,
    n14990, n14991, n14992, n14993, n14994, n14995,
    n14996, n14997, n14998, n14999, n15000, n15001,
    n15002, n15003, n15004, n15005, n15006, n15007,
    n15008, n15009, n15010, n15011, n15012, n15013,
    n15014, n15015, n15016, n15017, n15018, n15019,
    n15020, n15021, n15022, n15023, n15024, n15025,
    n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037,
    n15038, n15039, n15040, n15041, n15042, n15043,
    n15044, n15045, n15046, n15047, n15048, n15049,
    n15050, n15051, n15052, n15053, n15054, n15055,
    n15056, n15057, n15058, n15059, n15060, n15061,
    n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073,
    n15074, n15075, n15076, n15077, n15078, n15079,
    n15080, n15081, n15082, n15083, n15084, n15085,
    n15086, n15087, n15088, n15089, n15090, n15091,
    n15092, n15093, n15094, n15095, n15096, n15097,
    n15098, n15099, n15100, n15101, n15102, n15103,
    n15104, n15105, n15106, n15107, n15108, n15109,
    n15110, n15111, n15112, n15113, n15114, n15115,
    n15116, n15117, n15118, n15119, n15120, n15121,
    n15122, n15123, n15124, n15125, n15126, n15127,
    n15128, n15129, n15130, n15131, n15132, n15133,
    n15134, n15135, n15136, n15137, n15138, n15139,
    n15140, n15141, n15142, n15143, n15144, n15145,
    n15146, n15147, n15148, n15149, n15150, n15151,
    n15152, n15153, n15154, n15155, n15156, n15157,
    n15158, n15159, n15160, n15161, n15162, n15163,
    n15164, n15165, n15166, n15167, n15168, n15169,
    n15170, n15171, n15172, n15173, n15174, n15175,
    n15176, n15177, n15178, n15179, n15180, n15181,
    n15182, n15183, n15184, n15185, n15186, n15187,
    n15188, n15189, n15190, n15191, n15192, n15193,
    n15194, n15195, n15196, n15197, n15198, n15199,
    n15200, n15201, n15202, n15203, n15204, n15205,
    n15206, n15207, n15208, n15209, n15210, n15211,
    n15212, n15213, n15214, n15215, n15216, n15217,
    n15218, n15219, n15220, n15221, n15222, n15223,
    n15224, n15225, n15226, n15227, n15228, n15229,
    n15230, n15231, n15232, n15233, n15234, n15235,
    n15236, n15237, n15238, n15239, n15240, n15241,
    n15242, n15243, n15244, n15245, n15246, n15247,
    n15248, n15249, n15250, n15251, n15252, n15253,
    n15254, n15255, n15256, n15257, n15258, n15259,
    n15260, n15261, n15262, n15263, n15264, n15265,
    n15266, n15267, n15268, n15269, n15270, n15271,
    n15272, n15273, n15274, n15275, n15276, n15277,
    n15278, n15279, n15280, n15281, n15282, n15283,
    n15284, n15285, n15286, n15287, n15288, n15289,
    n15290, n15291, n15292, n15293, n15294, n15295,
    n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307,
    n15308, n15309, n15310, n15311, n15312, n15313,
    n15314, n15315, n15316, n15317, n15318, n15319,
    n15320, n15321, n15322, n15323, n15324, n15325,
    n15326, n15327, n15328, n15329, n15330, n15331,
    n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343,
    n15344, n15345, n15346, n15347, n15348, n15349,
    n15350, n15351, n15352, n15353, n15354, n15355,
    n15356, n15357, n15358, n15359, n15360, n15361,
    n15362, n15363, n15364, n15365, n15366, n15367,
    n15368, n15369, n15370, n15371, n15372, n15373,
    n15374, n15375, n15376, n15377, n15378, n15379,
    n15380, n15381, n15382, n15383, n15384, n15385,
    n15386, n15387, n15388, n15389, n15390, n15391,
    n15392, n15393, n15394, n15395, n15396, n15397,
    n15398, n15399, n15400, n15401, n15402, n15403,
    n15404, n15405, n15406, n15407, n15408, n15409,
    n15410, n15411, n15412, n15413, n15414, n15415,
    n15416, n15417, n15418, n15419, n15420, n15421,
    n15422, n15423, n15424, n15425, n15426, n15427,
    n15428, n15429, n15430, n15431, n15432, n15433,
    n15434, n15435, n15436, n15437, n15438, n15439,
    n15440, n15441, n15442, n15443, n15444, n15445,
    n15446, n15447, n15448, n15449, n15450, n15451,
    n15452, n15453, n15454, n15455, n15456, n15457,
    n15458, n15459, n15460, n15461, n15462, n15463,
    n15464, n15465, n15466, n15467, n15468, n15469,
    n15470, n15471, n15472, n15473, n15474, n15475,
    n15476, n15477, n15478, n15479, n15480, n15481,
    n15482, n15483, n15484, n15485, n15486, n15487,
    n15488, n15489, n15490, n15491, n15492, n15493,
    n15494, n15495, n15496, n15497, n15498, n15499,
    n15500, n15501, n15502, n15503, n15504, n15505,
    n15506, n15507, n15508, n15509, n15510, n15511,
    n15512, n15513, n15514, n15515, n15516, n15517,
    n15518, n15519, n15520, n15521, n15522, n15523,
    n15524, n15525, n15526, n15527, n15528, n15529,
    n15530, n15531, n15532, n15533, n15534, n15535,
    n15536, n15537, n15538, n15539, n15540, n15541,
    n15542, n15543, n15544, n15545, n15546, n15547,
    n15548, n15549, n15550, n15551, n15552, n15553,
    n15554, n15555, n15556, n15557, n15558, n15559,
    n15560, n15561, n15562, n15563, n15564, n15565,
    n15566, n15567, n15568, n15569, n15570, n15571,
    n15572, n15573, n15574, n15575, n15576, n15577,
    n15578, n15579, n15580, n15581, n15582, n15583,
    n15584, n15585, n15586, n15587, n15588, n15589,
    n15590, n15591, n15592, n15593, n15594, n15595,
    n15596, n15597, n15598, n15599, n15600, n15601,
    n15602, n15603, n15604, n15605, n15606, n15607,
    n15608, n15609, n15610, n15611, n15612, n15613,
    n15614, n15615, n15616, n15617, n15618, n15619,
    n15620, n15621, n15622, n15623, n15624, n15625,
    n15626, n15627, n15628, n15629, n15630, n15631,
    n15632, n15633, n15634, n15635, n15636, n15637,
    n15638, n15639, n15640, n15641, n15642, n15643,
    n15644, n15645, n15646, n15647, n15648, n15649,
    n15650, n15651, n15652, n15653, n15654, n15655,
    n15656, n15657, n15658, n15659, n15660, n15661,
    n15662, n15663, n15664, n15665, n15666, n15667,
    n15668, n15669, n15670, n15671, n15672, n15673,
    n15674, n15675, n15676, n15677, n15678, n15679,
    n15680, n15681, n15682, n15683, n15684, n15685,
    n15686, n15687, n15688, n15689, n15690, n15691,
    n15692, n15693, n15694, n15695, n15696, n15697,
    n15698, n15699, n15700, n15701, n15702, n15703,
    n15704, n15705, n15706, n15707, n15708, n15709,
    n15710, n15711, n15712, n15713, n15714, n15715,
    n15716, n15717, n15718, n15719, n15720, n15721,
    n15722, n15723, n15724, n15725, n15726, n15727,
    n15728, n15729, n15730, n15731, n15732, n15733,
    n15734, n15735, n15736, n15737, n15738, n15739,
    n15740, n15741, n15742, n15743, n15744, n15745,
    n15746, n15747, n15748, n15749, n15750, n15751,
    n15752, n15753, n15754, n15755, n15756, n15757,
    n15758, n15759, n15760, n15761, n15762, n15763,
    n15764, n15765, n15766, n15767, n15768, n15769,
    n15770, n15771, n15772, n15773, n15774, n15775,
    n15776, n15777, n15778, n15779, n15780, n15781,
    n15782, n15783, n15784, n15785, n15786, n15787,
    n15788, n15789, n15790, n15791, n15792, n15793,
    n15794, n15795, n15796, n15797, n15798, n15799,
    n15800, n15801, n15802, n15803, n15804, n15805,
    n15806, n15807, n15808, n15809, n15810, n15811,
    n15812, n15813, n15814, n15815, n15816, n15817,
    n15818, n15819, n15820, n15821, n15822, n15823,
    n15824, n15825, n15826, n15827, n15828, n15829,
    n15830, n15831, n15832, n15833, n15834, n15835,
    n15836, n15837, n15838, n15839, n15840, n15841,
    n15842, n15843, n15844, n15845, n15846, n15847,
    n15848, n15849, n15850, n15851, n15852, n15853,
    n15854, n15855, n15856, n15857, n15858, n15859,
    n15860, n15861, n15862, n15863, n15864, n15865,
    n15866, n15867, n15868, n15869, n15870, n15871,
    n15872, n15873, n15874, n15875, n15876, n15877,
    n15878, n15879, n15880, n15881, n15882, n15883,
    n15884, n15885, n15886, n15887, n15888, n15889,
    n15890, n15891, n15892, n15893, n15894, n15895,
    n15896, n15897, n15898, n15899, n15900, n15901,
    n15902, n15903, n15904, n15905, n15906, n15907,
    n15908, n15909, n15910, n15911, n15912, n15913,
    n15914, n15915, n15916, n15917, n15918, n15919,
    n15920, n15921, n15922, n15923, n15924, n15925,
    n15926, n15927, n15928, n15929, n15930, n15931,
    n15932, n15933, n15934, n15935, n15936, n15937,
    n15938, n15939, n15940, n15941, n15942, n15943,
    n15944, n15945, n15946, n15947, n15948, n15949,
    n15950, n15951, n15952, n15953, n15954, n15955,
    n15956, n15957, n15958, n15959, n15960, n15961,
    n15962, n15963, n15964, n15965, n15966, n15967,
    n15968, n15969, n15970, n15971, n15972, n15973,
    n15974, n15975, n15976, n15977, n15978, n15979,
    n15980, n15981, n15982, n15983, n15984, n15985,
    n15986, n15987, n15988, n15989, n15990, n15991,
    n15992, n15993, n15994, n15995, n15996, n15997,
    n15998, n15999, n16000, n16001, n16002, n16003,
    n16004, n16005, n16006, n16007, n16008, n16009,
    n16010, n16011, n16012, n16013, n16014, n16015,
    n16016, n16017, n16018, n16019, n16020, n16021,
    n16022, n16023, n16024, n16025, n16026, n16027,
    n16028, n16029, n16030, n16031, n16032, n16033,
    n16034, n16035, n16036, n16037, n16038, n16039,
    n16040, n16041, n16042, n16043, n16044, n16045,
    n16046, n16047, n16048, n16049, n16050, n16051,
    n16052, n16053, n16054, n16055, n16056, n16057,
    n16058, n16059, n16060, n16061, n16062, n16063,
    n16064, n16065, n16066, n16067, n16068, n16069,
    n16070, n16071, n16072, n16073, n16074, n16075,
    n16076, n16077, n16078, n16079, n16080, n16081,
    n16082, n16083, n16084, n16085, n16086, n16087,
    n16088, n16089, n16090, n16091, n16092, n16093,
    n16094, n16095, n16096, n16097, n16098, n16099,
    n16100, n16101, n16102, n16103, n16104, n16105,
    n16106, n16107, n16108, n16109, n16110, n16111,
    n16112, n16113, n16114, n16115, n16116, n16117,
    n16118, n16119, n16120, n16121, n16122, n16123,
    n16124, n16125, n16126, n16127, n16128, n16129,
    n16130, n16131, n16132, n16133, n16134, n16135,
    n16136, n16137, n16138, n16139, n16140, n16141,
    n16142, n16143, n16144, n16145, n16146, n16147,
    n16148, n16149, n16150, n16151, n16152, n16153,
    n16154, n16155, n16156, n16157, n16158, n16159,
    n16160, n16161, n16162, n16163, n16164, n16165,
    n16166, n16167, n16168, n16169, n16170, n16171,
    n16172, n16173, n16174, n16175, n16176, n16177,
    n16178, n16179, n16180, n16181, n16182, n16183,
    n16184, n16185, n16186, n16187, n16188, n16189,
    n16190, n16191, n16192, n16193, n16194, n16195,
    n16196, n16197, n16198, n16199, n16200, n16201,
    n16202, n16203, n16204, n16205, n16206, n16207,
    n16208, n16209, n16210, n16211, n16212, n16213,
    n16214, n16215, n16216, n16217, n16218, n16219,
    n16220, n16221, n16222, n16223, n16224, n16225,
    n16226, n16227, n16228, n16229, n16230, n16231,
    n16232, n16233, n16234, n16235, n16236, n16237,
    n16238, n16239, n16240, n16241, n16242, n16243,
    n16244, n16245, n16246, n16247, n16248, n16249,
    n16250, n16251, n16252, n16253, n16254, n16255,
    n16256, n16257, n16258, n16259, n16260, n16261,
    n16262, n16263, n16264, n16265, n16266, n16267,
    n16268, n16269, n16270, n16271, n16272, n16273,
    n16274, n16275, n16276, n16277, n16278, n16279,
    n16280, n16281, n16282, n16283, n16284, n16285,
    n16286, n16287, n16288, n16289, n16290, n16291,
    n16292, n16293, n16294, n16295, n16296, n16297,
    n16298, n16299, n16300, n16301, n16302, n16303,
    n16304, n16305, n16306, n16307, n16308, n16309,
    n16310, n16311, n16312, n16313, n16314, n16315,
    n16316, n16317, n16318, n16319, n16320, n16321,
    n16322, n16323, n16324, n16325, n16326, n16327,
    n16328, n16329, n16330, n16331, n16332, n16333,
    n16334, n16335, n16336, n16337, n16338, n16339,
    n16340, n16341, n16342, n16343, n16344, n16345,
    n16346, n16347, n16348, n16349, n16350, n16351,
    n16352, n16353, n16354, n16355, n16356, n16357,
    n16358, n16359, n16360, n16361, n16362, n16363,
    n16364, n16365, n16366, n16367, n16368, n16369,
    n16370, n16371, n16372, n16373, n16374, n16375,
    n16376, n16377, n16378, n16379, n16380, n16381,
    n16382, n16383, n16384, n16385, n16386, n16387,
    n16388, n16389, n16390, n16391, n16392, n16393,
    n16394, n16395, n16396, n16397, n16398, n16399,
    n16400, n16401, n16402, n16403, n16404, n16405,
    n16406, n16407, n16408, n16409, n16410, n16411,
    n16412, n16413, n16414, n16415, n16416, n16417,
    n16418, n16419, n16420, n16421, n16422, n16423,
    n16424, n16425, n16426, n16427, n16428, n16429,
    n16430, n16431, n16432, n16433, n16434, n16435,
    n16436, n16437, n16438, n16439, n16440, n16441,
    n16442, n16443, n16444, n16445, n16446, n16447,
    n16448, n16449, n16450, n16451, n16452, n16453,
    n16454, n16455, n16456, n16457, n16458, n16459,
    n16460, n16461, n16462, n16463, n16464, n16465,
    n16466, n16467, n16468, n16469, n16470, n16471,
    n16472, n16473, n16474, n16475, n16476, n16477,
    n16478, n16479, n16480, n16481, n16482, n16483,
    n16484, n16485, n16486, n16487, n16488, n16489,
    n16490, n16491, n16492, n16493, n16494, n16495,
    n16496, n16497, n16498, n16499, n16500, n16501,
    n16502, n16503, n16504, n16505, n16506, n16507,
    n16508, n16509, n16510, n16511, n16512, n16513,
    n16514, n16515, n16516, n16517, n16518, n16519,
    n16520, n16521, n16522, n16523, n16524, n16525,
    n16526, n16527, n16528, n16529, n16530, n16531,
    n16532, n16533, n16534, n16535, n16536, n16537,
    n16538, n16539, n16540, n16541, n16542, n16543,
    n16544, n16545, n16546, n16547, n16548, n16549,
    n16550, n16551, n16552, n16553, n16554, n16555,
    n16556, n16557, n16558, n16559, n16560, n16561,
    n16562, n16563, n16564, n16565, n16566, n16567,
    n16568, n16569, n16570, n16571, n16572, n16573,
    n16574, n16575, n16576, n16577, n16578, n16579,
    n16580, n16581, n16582, n16583, n16584, n16585,
    n16586, n16587, n16588, n16589, n16590, n16591,
    n16592, n16593, n16594, n16595, n16596, n16597,
    n16598, n16599, n16600, n16601, n16602, n16603,
    n16604, n16605, n16606, n16607, n16608, n16609,
    n16610, n16611, n16612, n16613, n16614, n16615,
    n16616, n16617, n16618, n16619, n16620, n16621,
    n16622, n16623, n16624, n16625, n16626, n16627,
    n16628, n16629, n16630, n16631, n16632, n16633,
    n16634, n16635, n16636, n16637, n16638, n16639,
    n16640, n16641, n16642, n16643, n16644, n16645,
    n16646, n16647, n16648, n16649, n16650, n16651,
    n16652, n16653, n16654, n16655, n16656, n16657,
    n16658, n16659, n16660, n16661, n16662, n16663,
    n16664, n16665, n16666, n16667, n16668, n16669,
    n16670, n16671, n16672, n16673, n16674, n16675,
    n16676, n16677, n16678, n16679, n16680, n16681,
    n16682, n16683, n16684, n16685, n16686, n16687,
    n16688, n16689, n16690, n16691, n16692, n16693,
    n16694, n16695, n16696, n16697, n16698, n16699,
    n16700, n16701, n16702, n16703, n16704, n16705,
    n16706, n16707, n16708, n16709, n16710, n16711,
    n16712, n16713, n16714, n16715, n16716, n16717,
    n16718, n16719, n16720, n16721, n16722, n16723,
    n16724, n16725, n16726, n16727, n16728, n16729,
    n16730, n16731, n16732, n16733, n16734, n16735,
    n16736, n16737, n16738, n16739, n16740, n16741,
    n16742, n16743, n16744, n16745, n16746, n16747,
    n16748, n16749, n16750, n16751, n16752, n16753,
    n16754, n16755, n16756, n16757, n16758, n16759,
    n16760, n16761, n16762, n16763, n16764, n16765,
    n16766, n16767, n16768, n16769, n16770, n16771,
    n16772, n16773, n16774, n16775, n16776, n16777,
    n16778, n16779, n16780, n16781, n16782, n16783,
    n16784, n16785, n16786, n16787, n16788, n16789,
    n16790, n16791, n16792, n16793, n16794, n16795,
    n16796, n16797, n16798, n16799, n16800, n16801,
    n16802, n16803, n16804, n16805, n16806, n16807,
    n16808, n16809, n16810, n16811, n16812, n16813,
    n16814, n16815, n16816, n16817, n16818, n16819,
    n16820, n16821, n16822, n16823, n16824, n16825,
    n16826, n16827, n16828, n16829, n16830, n16831,
    n16832, n16833, n16834, n16835, n16836, n16837,
    n16838, n16839, n16840, n16841, n16842, n16843,
    n16844, n16845, n16846, n16847, n16848, n16849,
    n16850, n16851, n16852, n16853, n16854, n16855,
    n16856, n16857, n16858, n16859, n16860, n16861,
    n16862, n16863, n16864, n16865, n16866, n16867,
    n16868, n16869, n16870, n16871, n16872, n16873,
    n16874, n16875, n16876, n16877, n16878, n16879,
    n16880, n16881, n16882, n16883, n16884, n16885,
    n16886, n16887, n16888, n16889, n16890, n16891,
    n16892, n16893, n16894, n16895, n16896, n16897,
    n16898, n16899, n16900, n16901, n16902, n16903,
    n16904, n16905, n16906, n16907, n16908, n16909,
    n16910, n16911, n16912, n16913, n16914, n16915,
    n16916, n16917, n16918, n16919, n16920, n16921,
    n16922, n16923, n16924, n16925, n16926, n16927,
    n16928, n16929, n16930, n16931, n16932, n16933,
    n16934, n16935, n16936, n16937, n16938, n16939,
    n16940, n16941, n16942, n16943, n16944, n16945,
    n16946, n16947, n16948, n16949, n16950, n16951,
    n16952, n16953, n16954, n16955, n16956, n16957,
    n16958, n16959, n16960, n16961, n16962, n16963,
    n16964, n16965, n16966, n16967, n16968, n16969,
    n16970, n16971, n16972, n16973, n16974, n16975,
    n16976, n16977, n16978, n16979, n16980, n16981,
    n16982, n16983, n16984, n16985, n16986, n16987,
    n16988, n16989, n16990, n16991, n16992, n16993,
    n16994, n16995, n16996, n16997, n16998, n16999,
    n17000, n17001, n17002, n17003, n17004, n17005,
    n17006, n17007, n17008, n17009, n17010, n17011,
    n17012, n17013, n17014, n17015, n17016, n17017,
    n17018, n17019, n17020, n17021, n17022, n17023,
    n17024, n17025, n17026, n17027, n17028, n17029,
    n17030, n17031, n17032, n17033, n17034, n17035,
    n17036, n17037, n17038, n17039, n17040, n17041,
    n17042, n17043, n17044, n17045, n17046, n17047,
    n17048, n17049, n17050, n17051, n17052, n17053,
    n17054, n17055, n17056, n17057, n17058, n17059,
    n17060, n17061, n17062, n17063, n17064, n17065,
    n17066, n17067, n17068, n17069, n17070, n17071,
    n17072, n17073, n17074, n17075, n17076, n17077,
    n17078, n17079, n17080, n17081, n17082, n17083,
    n17084, n17085, n17086, n17087, n17088, n17089,
    n17090, n17091, n17092, n17093, n17094, n17095,
    n17096, n17097, n17098, n17099, n17100, n17101,
    n17102, n17103, n17104, n17105, n17106, n17107,
    n17108, n17109, n17110, n17111, n17112, n17113,
    n17114, n17115, n17116, n17117, n17118, n17119,
    n17120, n17121, n17122, n17123, n17124, n17125,
    n17126, n17127, n17128, n17129, n17130, n17131,
    n17132, n17133, n17134, n17135, n17136, n17137,
    n17138, n17139, n17140, n17141, n17142, n17143,
    n17144, n17145, n17146, n17147, n17148, n17149,
    n17150, n17151, n17152, n17153, n17154, n17155,
    n17156, n17157, n17158, n17159, n17160, n17161,
    n17162, n17163, n17164, n17165, n17166, n17167,
    n17168, n17169, n17170, n17171, n17172, n17173,
    n17174, n17175, n17176, n17177, n17178, n17179,
    n17180, n17181, n17182, n17183, n17184, n17185,
    n17186, n17187, n17188, n17189, n17190, n17191,
    n17192, n17193, n17194, n17195, n17196, n17197,
    n17198, n17199, n17200, n17201, n17202, n17203,
    n17204, n17205, n17206, n17207, n17208, n17209,
    n17210, n17211, n17212, n17213, n17214, n17215,
    n17216, n17217, n17218, n17219, n17220, n17221,
    n17222, n17223, n17224, n17225, n17226, n17227,
    n17228, n17229, n17230, n17231, n17232, n17233,
    n17234, n17235, n17236, n17237, n17238, n17239,
    n17240, n17241, n17242, n17243, n17244, n17245,
    n17246, n17247, n17248, n17249, n17250, n17251,
    n17252, n17253, n17254, n17255, n17256, n17257,
    n17258, n17259, n17260, n17261, n17262, n17263,
    n17264, n17265, n17266, n17267, n17268, n17269,
    n17270, n17271, n17272, n17273, n17274, n17275,
    n17276, n17277, n17278, n17279, n17280, n17281,
    n17282, n17283, n17284, n17285, n17286, n17287,
    n17288, n17289, n17290, n17291, n17292, n17293,
    n17294, n17295, n17296, n17297, n17298, n17299,
    n17300, n17301, n17302, n17303, n17304, n17305,
    n17306, n17307, n17308, n17309, n17310, n17311,
    n17312, n17313, n17314, n17315, n17316, n17317,
    n17318, n17319, n17320, n17321, n17322, n17323,
    n17324, n17325, n17326, n17327, n17328, n17329,
    n17330, n17331, n17332, n17333, n17334, n17335,
    n17336, n17337, n17338, n17339, n17340, n17341,
    n17342, n17343, n17344, n17345, n17346, n17347,
    n17348, n17349, n17350, n17351, n17352, n17353,
    n17354, n17355, n17356, n17357, n17358, n17359,
    n17360, n17361, n17362, n17363, n17364, n17365,
    n17366, n17367, n17368, n17369, n17370, n17371,
    n17372, n17373, n17374, n17375, n17376, n17377,
    n17378, n17379, n17380, n17381, n17382, n17383,
    n17384, n17385, n17386, n17387, n17388, n17389,
    n17390, n17391, n17392, n17393, n17394, n17395,
    n17396, n17397, n17398, n17399, n17400, n17401,
    n17402, n17403, n17404, n17405, n17406, n17407,
    n17408, n17409, n17410, n17411, n17412, n17413,
    n17414, n17415, n17416, n17417, n17418, n17419,
    n17420, n17421, n17422, n17423, n17424, n17425,
    n17426, n17427, n17428, n17429, n17430, n17431,
    n17432, n17433, n17434, n17435, n17436, n17437,
    n17438, n17439, n17440, n17441, n17442, n17443,
    n17444, n17445, n17446, n17447, n17448, n17449,
    n17450, n17451, n17452, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461,
    n17462, n17463, n17464, n17465, n17466, n17467,
    n17468, n17469, n17470, n17471, n17472, n17473,
    n17474, n17475, n17476, n17477, n17478, n17479,
    n17480, n17481, n17482, n17483, n17484, n17485,
    n17486, n17487, n17488, n17489, n17490, n17491,
    n17492, n17493, n17494, n17495, n17496, n17497,
    n17498, n17499, n17500, n17501, n17502, n17503,
    n17504, n17505, n17506, n17507, n17508, n17509,
    n17510, n17511, n17512, n17513, n17514, n17515,
    n17516, n17517, n17518, n17519, n17520, n17521,
    n17522, n17523, n17524, n17525, n17526, n17527,
    n17528, n17529, n17530, n17531, n17532, n17533,
    n17534, n17535, n17536, n17537, n17538, n17539,
    n17540, n17541, n17542, n17543, n17544, n17545,
    n17546, n17547, n17548, n17549, n17550, n17551,
    n17552, n17553, n17554, n17555, n17556, n17557,
    n17558, n17559, n17560, n17561, n17562, n17563,
    n17564, n17565, n17566, n17567, n17568, n17569,
    n17570, n17571, n17572, n17573, n17574, n17575,
    n17576, n17577, n17578, n17579, n17580, n17581,
    n17582, n17583, n17584, n17585, n17586, n17587,
    n17588, n17589, n17590, n17591, n17592, n17593,
    n17594, n17595, n17596, n17597, n17598, n17599,
    n17600, n17601, n17602, n17603, n17604, n17605,
    n17606, n17607, n17608, n17609, n17610, n17611,
    n17612, n17613, n17614, n17615, n17616, n17617,
    n17618, n17619, n17620, n17621, n17622, n17623,
    n17624, n17625, n17626, n17627, n17628, n17629,
    n17630, n17631, n17632, n17633, n17634, n17635,
    n17636, n17637, n17638, n17639, n17640, n17641,
    n17642, n17643, n17644, n17645, n17646, n17647,
    n17648, n17649, n17650, n17651, n17652, n17653,
    n17654, n17655, n17656, n17657, n17658, n17659,
    n17660, n17661, n17662, n17663, n17664, n17665,
    n17666, n17667, n17668, n17669, n17670, n17671,
    n17672, n17673, n17674, n17675, n17676, n17677,
    n17678, n17679, n17680, n17681, n17682, n17683,
    n17684, n17685, n17686, n17687, n17688, n17689,
    n17690, n17691, n17692, n17693, n17694, n17695,
    n17696, n17697, n17698, n17699, n17700, n17701,
    n17702, n17703, n17704, n17705, n17706, n17707,
    n17708, n17709, n17710, n17711, n17712, n17713,
    n17714, n17715, n17716, n17717, n17718, n17719,
    n17720, n17721, n17722, n17723, n17724, n17725,
    n17726, n17727, n17728, n17729, n17730, n17731,
    n17732, n17733, n17734, n17735, n17736, n17737,
    n17738, n17739, n17740, n17741, n17742, n17743,
    n17744, n17745, n17746, n17747, n17748, n17749,
    n17750, n17751, n17752, n17753, n17754, n17755,
    n17756, n17757, n17758, n17759, n17760, n17761,
    n17762, n17763, n17764, n17765, n17766, n17767,
    n17768, n17769, n17770, n17771, n17772, n17773,
    n17774, n17775, n17776, n17777, n17778, n17779,
    n17780, n17781, n17782, n17783, n17784, n17785,
    n17786, n17787, n17788, n17789, n17790, n17791,
    n17792, n17793, n17794, n17795, n17796, n17797,
    n17798, n17799, n17800, n17801, n17802, n17803,
    n17804, n17805, n17806, n17807, n17808, n17809,
    n17810, n17811, n17812, n17813, n17814, n17815,
    n17816, n17817, n17818, n17819, n17820, n17821,
    n17822, n17823, n17824, n17825, n17826, n17827,
    n17828, n17829, n17830, n17831, n17832, n17833,
    n17834, n17835, n17836, n17837, n17838, n17839,
    n17840, n17841, n17842, n17843, n17844, n17845,
    n17846, n17847, n17848, n17849, n17850, n17851,
    n17852, n17853, n17854, n17855, n17856, n17857,
    n17858, n17859, n17860, n17861, n17862, n17863,
    n17864, n17865, n17866, n17867, n17868, n17869,
    n17870, n17871, n17872, n17873, n17874, n17875,
    n17876, n17877, n17878, n17879, n17880, n17881,
    n17882, n17883, n17884, n17885, n17886, n17887,
    n17888, n17889, n17890, n17891, n17892, n17893,
    n17894, n17895, n17896, n17897, n17898, n17899,
    n17900, n17901, n17902, n17903, n17904, n17905,
    n17906, n17907, n17908, n17909, n17910, n17911,
    n17912, n17913, n17914, n17915, n17916, n17917,
    n17918, n17919, n17920, n17921, n17922, n17923,
    n17924, n17925, n17926, n17927, n17928, n17929,
    n17930, n17931, n17932, n17933, n17934, n17935,
    n17936, n17937, n17938, n17939, n17940, n17941,
    n17942, n17943, n17944, n17945, n17946, n17947,
    n17948, n17949, n17950, n17951, n17952, n17953,
    n17954, n17955, n17956, n17957, n17958, n17959,
    n17960, n17961, n17962, n17963, n17964, n17965,
    n17966, n17967, n17968, n17969, n17970, n17971,
    n17972, n17973, n17974, n17975, n17976, n17977,
    n17978, n17979, n17980, n17981, n17982, n17983,
    n17984, n17985, n17986, n17987, n17988, n17989,
    n17990, n17991, n17992, n17993, n17994, n17995,
    n17996, n17997, n17998, n17999, n18000, n18001,
    n18002, n18003, n18004, n18005, n18006, n18007,
    n18008, n18009, n18010, n18011, n18012, n18013,
    n18014, n18015, n18016, n18017, n18018, n18019,
    n18020, n18021, n18022, n18023, n18024, n18025,
    n18026, n18027, n18028, n18029, n18030, n18031,
    n18032, n18033, n18034, n18035, n18036, n18037,
    n18038, n18039, n18040, n18041, n18042, n18043,
    n18044, n18045, n18046, n18047, n18048, n18049,
    n18050, n18051, n18052, n18053, n18054, n18055,
    n18056, n18057, n18058, n18059, n18060, n18061,
    n18062, n18063, n18064, n18065, n18066, n18067,
    n18068, n18069, n18070, n18071, n18072, n18073,
    n18074, n18075, n18076, n18077, n18078, n18079,
    n18080, n18081, n18082, n18083, n18084, n18085,
    n18086, n18087, n18088, n18089, n18090, n18091,
    n18092, n18093, n18094, n18095, n18096, n18097,
    n18098, n18099, n18100, n18101, n18102, n18103,
    n18104, n18105, n18106, n18107, n18108, n18109,
    n18110, n18111, n18112, n18113, n18114, n18115,
    n18116, n18117, n18118, n18119, n18120, n18121,
    n18122, n18123, n18124, n18125, n18126, n18127,
    n18128, n18129, n18130, n18131, n18132, n18133,
    n18134, n18135, n18136, n18137, n18138, n18139,
    n18140, n18141, n18142, n18143, n18144, n18145,
    n18146, n18147, n18148, n18149, n18150, n18151,
    n18152, n18153, n18154, n18155, n18156, n18157,
    n18158, n18159, n18160, n18161, n18162, n18163,
    n18164, n18165, n18166, n18167, n18168, n18169,
    n18170, n18171, n18172, n18173, n18174, n18175,
    n18176, n18177, n18178, n18179, n18180, n18181,
    n18182, n18183, n18184, n18185, n18186, n18187,
    n18188, n18189, n18190, n18191, n18192, n18193,
    n18194, n18195, n18196, n18197, n18198, n18199,
    n18200, n18201, n18202, n18203, n18204, n18205,
    n18206, n18207, n18208, n18209, n18210, n18211,
    n18212, n18213, n18214, n18215, n18216, n18217,
    n18218, n18219, n18220, n18221, n18222, n18223,
    n18224, n18225, n18226, n18227, n18228, n18229,
    n18230, n18231, n18232, n18233, n18234, n18235,
    n18236, n18237, n18238, n18239, n18240, n18241,
    n18242, n18243, n18244, n18245, n18246, n18247,
    n18248, n18249, n18250, n18251, n18252, n18253,
    n18254, n18255, n18256, n18257, n18258, n18259,
    n18260, n18261, n18262, n18263, n18264, n18265,
    n18266, n18267, n18268, n18269, n18270, n18271,
    n18272, n18273, n18274, n18275, n18276, n18277,
    n18278, n18279, n18280, n18281, n18282, n18283,
    n18284, n18285, n18286, n18287, n18288, n18289,
    n18290, n18291, n18292, n18293, n18294, n18295,
    n18296, n18297, n18298, n18299, n18300, n18301,
    n18302, n18303, n18304, n18305, n18306, n18307,
    n18308, n18309, n18310, n18311, n18312, n18313,
    n18314, n18315, n18316, n18317, n18318, n18319,
    n18320, n18321, n18322, n18323, n18324, n18325,
    n18326, n18327, n18328, n18329, n18330, n18331,
    n18332, n18333, n18334, n18335, n18336, n18337,
    n18338, n18339, n18340, n18341, n18342, n18343,
    n18344, n18345, n18346, n18347, n18348, n18349,
    n18350, n18351, n18352, n18353, n18354, n18355,
    n18356, n18357, n18358, n18359, n18360, n18361,
    n18362, n18363, n18364, n18365, n18366, n18367,
    n18368, n18369, n18370, n18371, n18372, n18373,
    n18374, n18375, n18376, n18377, n18378, n18379,
    n18380, n18381, n18382, n18383, n18384, n18385,
    n18386, n18387, n18388, n18389, n18390, n18391,
    n18392, n18393, n18394, n18395, n18396, n18397,
    n18398, n18399, n18400, n18401, n18402, n18403,
    n18404, n18405, n18406, n18407, n18408, n18409,
    n18410, n18411, n18412, n18413, n18414, n18415,
    n18416, n18417, n18418, n18419, n18420, n18421,
    n18422, n18423, n18424, n18425, n18426, n18427,
    n18428, n18429, n18430, n18431, n18432, n18433,
    n18434, n18435, n18436, n18437, n18438, n18439,
    n18440, n18441, n18442, n18443, n18444, n18445,
    n18446, n18447, n18448, n18449, n18450, n18451,
    n18452, n18453, n18454, n18455, n18456, n18457,
    n18458, n18459, n18460, n18461, n18462, n18463,
    n18464, n18465, n18466, n18467, n18468, n18469,
    n18470, n18471, n18472, n18473, n18474, n18475,
    n18476, n18477, n18478, n18479, n18480, n18481,
    n18482, n18483, n18484, n18485, n18486, n18487,
    n18488, n18489, n18490, n18491, n18492, n18493,
    n18494, n18495, n18496, n18497, n18498, n18499,
    n18500, n18501, n18502, n18503, n18504, n18505,
    n18506, n18507, n18508, n18509, n18510, n18511,
    n18512, n18513, n18514, n18515, n18516, n18517,
    n18518, n18519, n18520, n18521, n18522, n18523,
    n18524, n18525, n18526, n18527, n18528, n18529,
    n18530, n18531, n18532, n18533, n18534, n18535,
    n18536, n18537, n18538, n18539, n18540, n18541,
    n18542, n18543, n18544, n18545, n18546, n18547,
    n18548, n18549, n18550, n18551, n18552, n18553,
    n18554, n18555, n18556, n18557, n18558, n18559,
    n18560, n18561, n18562, n18563, n18564, n18565,
    n18566, n18567, n18568, n18569, n18570, n18571,
    n18572, n18573, n18574, n18575, n18576, n18577,
    n18578, n18579, n18580, n18581, n18582, n18583,
    n18584, n18585, n18586, n18587, n18588, n18589,
    n18590, n18591, n18592, n18593, n18594, n18595,
    n18596, n18597, n18598, n18599, n18600, n18601,
    n18602, n18603, n18604, n18605, n18606, n18607,
    n18608, n18609, n18610, n18611, n18612, n18613,
    n18614, n18615, n18616, n18617, n18618, n18619,
    n18620, n18621, n18622, n18623, n18624, n18625,
    n18626, n18627, n18628, n18629, n18630, n18631,
    n18632, n18633, n18634, n18635, n18636, n18637,
    n18638, n18639, n18640, n18641, n18642, n18643,
    n18644, n18645, n18646, n18647, n18648, n18649,
    n18650, n18651, n18652, n18653, n18654, n18655,
    n18656, n18657, n18658, n18659, n18660, n18661,
    n18662, n18663, n18664, n18665, n18666, n18667,
    n18668, n18669, n18670, n18671, n18672, n18673,
    n18674, n18675, n18676, n18677, n18678, n18679,
    n18680, n18681, n18682, n18683, n18684, n18685,
    n18686, n18687, n18688, n18689, n18690, n18691,
    n18692, n18693, n18694, n18695, n18696, n18697,
    n18698, n18699, n18700, n18701, n18702, n18703,
    n18704, n18705, n18706, n18707, n18708, n18709,
    n18710, n18711, n18712, n18713, n18714, n18715,
    n18716, n18717, n18718, n18719, n18720, n18721,
    n18722, n18723, n18724, n18725, n18726, n18727,
    n18728, n18729, n18730, n18731, n18732, n18733,
    n18734, n18735, n18736, n18737, n18738, n18739,
    n18740, n18741, n18742, n18743, n18744, n18745,
    n18746, n18747, n18748, n18749, n18750, n18751,
    n18752, n18753, n18754, n18755, n18756, n18757,
    n18758, n18759, n18760, n18761, n18762, n18763,
    n18764, n18765, n18766, n18767, n18768, n18769,
    n18770, n18771, n18772, n18773, n18774, n18775,
    n18776, n18777, n18778, n18779, n18780, n18781,
    n18782, n18783, n18784, n18785, n18786, n18787,
    n18788, n18789, n18790, n18791, n18792, n18793,
    n18794, n18795, n18796, n18797, n18798, n18799,
    n18800, n18801, n18802, n18803, n18804, n18805,
    n18806, n18807, n18808, n18809, n18810, n18811,
    n18812, n18813, n18814, n18815, n18816, n18817,
    n18818, n18819, n18820, n18821, n18822, n18823,
    n18824, n18825, n18826, n18827, n18828, n18829,
    n18830, n18831, n18832, n18833, n18834, n18835,
    n18836, n18837, n18838, n18839, n18840, n18841,
    n18842, n18843, n18844, n18845, n18846, n18847,
    n18848, n18849, n18850, n18851, n18852, n18853,
    n18854, n18855, n18856, n18857, n18858, n18859,
    n18860, n18861, n18862, n18863, n18864, n18865,
    n18866, n18867, n18868, n18869, n18870, n18871,
    n18872, n18873, n18874, n18875, n18876, n18877,
    n18878, n18879, n18880, n18881, n18882, n18883,
    n18884, n18885, n18886, n18887, n18888, n18889,
    n18890, n18891, n18892, n18893, n18894, n18895,
    n18896, n18897, n18898, n18899, n18900, n18901,
    n18902, n18903, n18904, n18905, n18906, n18907,
    n18908, n18909, n18910, n18911, n18912, n18913,
    n18914, n18915, n18916, n18917, n18918, n18919,
    n18920, n18921, n18922, n18923, n18924, n18925,
    n18926, n18927, n18928, n18929, n18930, n18931,
    n18932, n18933, n18934, n18935, n18936, n18937,
    n18938, n18939, n18940, n18941, n18942, n18943,
    n18944, n18945, n18946, n18947, n18948, n18949,
    n18950, n18951, n18952, n18953, n18954, n18955,
    n18956, n18957, n18958, n18959, n18960, n18961,
    n18962, n18963, n18964, n18965, n18966, n18967,
    n18968, n18969, n18970, n18971, n18972, n18973,
    n18974, n18975, n18976, n18977, n18978, n18979,
    n18980, n18981, n18982, n18983, n18984, n18985,
    n18986, n18987, n18988, n18989, n18990, n18991,
    n18992, n18993, n18994, n18995, n18996, n18997,
    n18998, n18999, n19000, n19001, n19002, n19003,
    n19004, n19005, n19006, n19007, n19008, n19009,
    n19010, n19011, n19012, n19013, n19014, n19015,
    n19016, n19017, n19018, n19019, n19020, n19021,
    n19022, n19023, n19024, n19025, n19026, n19027,
    n19028, n19029, n19030, n19031, n19032, n19033,
    n19034, n19035, n19036, n19037, n19038, n19039,
    n19040, n19041, n19042, n19043, n19044, n19045,
    n19046, n19047, n19048, n19049, n19050, n19051,
    n19052, n19053, n19054, n19055, n19056, n19057,
    n19058, n19059, n19060, n19061, n19062, n19063,
    n19064, n19065, n19066, n19067, n19068, n19069,
    n19070, n19071, n19072, n19073, n19074, n19075,
    n19076, n19077, n19078, n19079, n19080, n19081,
    n19082, n19083, n19084, n19085, n19086, n19087,
    n19088, n19089, n19090, n19091, n19092, n19093,
    n19094, n19095, n19096, n19097, n19098, n19099,
    n19100, n19101, n19102, n19103, n19104, n19105,
    n19106, n19107, n19108, n19109, n19110, n19111,
    n19112, n19113, n19114, n19115, n19116, n19117,
    n19118, n19119, n19120, n19121, n19122, n19123,
    n19124, n19125, n19126, n19127, n19128, n19129,
    n19130, n19131, n19132, n19133, n19134, n19135,
    n19136, n19137, n19138, n19139, n19140, n19141,
    n19142, n19143, n19144, n19145, n19146, n19147,
    n19148, n19149, n19150, n19151, n19152, n19153,
    n19154, n19155, n19156, n19157, n19158, n19159,
    n19160, n19161, n19162, n19163, n19164, n19165,
    n19166, n19167, n19168, n19169, n19170, n19171,
    n19172, n19173, n19174, n19175, n19176, n19177,
    n19178, n19179, n19180, n19181, n19182, n19183,
    n19184, n19185, n19186, n19187, n19188, n19189,
    n19190, n19191, n19192, n19193, n19194, n19195,
    n19196, n19197, n19198, n19199, n19200, n19201,
    n19202, n19203, n19204, n19205, n19206, n19207,
    n19208, n19209, n19210, n19211, n19212, n19213,
    n19214, n19215, n19216, n19217, n19218, n19219,
    n19220, n19221, n19222, n19223, n19224, n19225,
    n19226, n19227, n19228, n19229, n19230, n19231,
    n19232, n19233, n19234, n19235, n19236, n19237,
    n19238, n19239, n19240, n19241, n19242, n19243,
    n19244, n19245, n19246, n19247, n19248, n19249,
    n19250, n19251, n19252, n19253, n19254, n19255,
    n19256, n19257, n19258, n19259, n19260, n19261,
    n19262, n19263, n19264, n19265, n19266, n19267,
    n19268, n19269, n19270, n19271, n19272, n19273,
    n19274, n19275, n19276, n19277, n19278, n19279,
    n19280, n19281, n19282, n19283, n19284, n19285,
    n19286, n19287, n19288, n19289, n19290, n19291,
    n19292, n19293, n19294, n19295, n19296, n19297,
    n19298, n19299, n19300, n19301, n19302, n19303,
    n19304, n19305, n19306, n19307, n19308, n19309,
    n19310, n19311, n19312, n19313, n19314, n19315,
    n19316, n19317, n19318, n19319, n19320, n19321,
    n19322, n19323, n19324, n19325, n19326, n19327,
    n19328, n19329, n19330, n19331, n19332, n19333,
    n19334, n19335, n19336, n19337, n19338, n19339,
    n19340, n19341, n19342, n19343, n19344, n19345,
    n19346, n19347, n19348, n19349, n19350, n19351,
    n19352, n19353, n19354, n19355, n19356, n19357,
    n19358, n19359, n19360, n19361, n19362, n19363,
    n19364, n19365, n19366, n19367, n19368, n19369,
    n19370, n19371, n19372, n19373, n19374, n19375,
    n19376, n19377, n19378, n19379, n19380, n19381,
    n19382, n19383, n19384, n19385, n19386, n19387,
    n19388, n19389, n19390, n19391, n19392, n19393,
    n19394, n19395, n19396, n19397, n19398, n19399,
    n19400, n19401, n19402, n19403, n19404, n19405,
    n19406, n19407, n19408, n19409, n19410, n19411,
    n19412, n19413, n19414, n19415, n19416, n19417,
    n19418, n19419, n19420, n19421, n19422, n19423,
    n19424, n19425, n19426, n19427, n19428, n19429,
    n19430, n19431, n19432, n19433, n19434, n19435,
    n19436, n19437, n19438, n19439, n19440, n19441,
    n19442, n19443, n19444, n19445, n19446, n19447,
    n19448, n19449, n19450, n19451, n19452, n19453,
    n19454, n19455, n19456, n19457, n19458, n19459,
    n19460, n19461, n19462, n19463, n19464, n19465,
    n19466, n19467, n19468, n19469, n19470, n19471,
    n19472, n19473, n19474, n19475, n19476, n19477,
    n19478, n19479, n19480, n19481, n19482, n19483,
    n19484, n19485, n19486, n19487, n19488, n19489,
    n19490, n19491, n19492, n19493, n19494, n19495,
    n19496, n19497, n19498, n19499, n19500, n19501,
    n19502, n19503, n19504, n19505, n19506, n19507,
    n19508, n19509, n19510, n19511, n19512, n19513,
    n19514, n19515, n19516, n19517, n19518, n19519,
    n19520, n19521, n19522, n19523, n19524, n19525,
    n19526, n19527, n19528, n19529, n19530, n19531,
    n19532, n19533, n19534, n19535, n19536, n19537,
    n19538, n19539, n19540, n19541, n19542, n19543,
    n19544, n19545, n19546, n19547, n19548, n19549,
    n19550, n19551, n19552, n19553, n19554, n19555,
    n19556, n19557, n19558, n19559, n19560, n19561,
    n19562, n19563, n19564, n19565, n19566, n19567,
    n19568, n19569, n19570, n19571, n19572, n19573,
    n19574, n19575, n19576, n19577, n19578, n19579,
    n19580, n19581, n19582, n19583, n19584, n19585,
    n19586, n19587, n19588, n19589, n19590, n19591,
    n19592, n19593, n19594, n19595, n19596, n19597,
    n19598, n19599, n19600, n19601, n19602, n19603,
    n19604, n19605, n19606, n19607, n19608, n19609,
    n19610, n19611, n19612, n19613, n19614, n19615,
    n19616, n19617, n19618, n19619, n19620, n19621,
    n19622, n19623, n19624, n19625, n19626, n19627,
    n19628, n19629, n19630, n19631, n19632, n19633,
    n19634, n19635, n19636, n19637, n19638, n19639,
    n19640, n19641, n19642, n19643, n19644, n19645,
    n19646, n19647, n19648, n19649, n19650, n19651,
    n19652, n19653, n19654, n19655, n19656, n19657,
    n19658, n19659, n19660, n19661, n19662, n19663,
    n19664, n19665, n19666, n19667, n19668, n19669,
    n19670, n19671, n19672, n19673, n19674, n19675,
    n19676, n19677, n19678, n19679, n19680, n19681,
    n19682, n19683, n19684, n19685, n19686, n19687,
    n19688, n19689, n19690, n19691, n19692, n19693,
    n19694, n19695, n19696, n19697, n19698, n19699,
    n19700, n19701, n19702, n19703, n19704, n19705,
    n19706, n19707, n19708, n19709, n19710, n19711,
    n19712, n19713, n19714, n19715, n19716, n19717,
    n19718, n19719, n19720, n19721, n19722, n19723,
    n19724, n19725, n19726, n19727, n19728, n19729,
    n19730, n19731, n19732, n19733, n19734, n19735,
    n19736, n19737, n19738, n19739, n19740, n19741,
    n19742, n19743, n19744, n19745, n19746, n19747,
    n19748, n19749, n19750, n19751, n19752, n19753,
    n19754, n19755, n19756, n19757, n19758, n19759,
    n19760, n19761, n19762, n19763, n19764, n19765,
    n19766, n19767, n19768, n19769, n19770, n19771,
    n19772, n19773, n19774, n19775, n19776, n19777,
    n19778, n19779, n19780, n19781, n19782, n19783,
    n19784, n19785, n19786, n19787, n19788, n19789,
    n19790, n19791, n19792, n19793, n19794, n19795,
    n19796, n19797, n19798, n19799, n19800, n19801,
    n19802, n19803, n19804, n19805, n19806, n19807,
    n19808, n19809, n19810, n19811, n19812, n19813,
    n19814, n19815, n19816, n19817, n19818, n19819,
    n19820, n19821, n19822, n19823, n19824, n19825,
    n19826, n19827, n19828, n19829, n19830, n19831,
    n19832, n19833, n19834, n19835, n19836, n19837,
    n19838, n19839, n19840, n19841, n19842, n19843,
    n19844, n19845, n19846, n19847, n19848, n19849,
    n19850, n19851, n19852, n19853, n19854, n19855,
    n19856, n19857, n19858, n19859, n19860, n19861,
    n19862, n19863, n19864, n19865, n19866, n19867,
    n19868, n19869, n19870, n19871, n19872, n19873,
    n19874, n19875, n19876, n19877, n19878, n19879,
    n19880, n19881, n19882, n19883, n19884, n19885,
    n19886, n19887, n19888, n19889, n19890, n19891,
    n19892, n19893, n19894, n19895, n19896, n19897,
    n19898, n19899, n19900, n19901, n19902, n19903,
    n19904, n19905, n19906, n19907, n19908, n19909,
    n19910, n19911, n19912, n19913, n19914, n19915,
    n19916, n19917, n19918, n19919, n19920, n19921,
    n19922, n19923, n19924, n19925, n19926, n19927,
    n19928, n19929, n19930, n19931, n19932, n19933,
    n19934, n19935, n19936, n19937, n19938, n19939,
    n19940, n19941, n19942, n19943, n19944, n19945,
    n19946, n19947, n19948, n19949, n19950, n19951,
    n19952, n19953, n19954, n19955, n19956, n19957,
    n19958, n19959, n19960, n19961, n19962, n19963,
    n19964, n19965, n19966, n19967, n19968, n19969,
    n19970, n19971, n19972, n19973, n19974, n19975,
    n19976, n19977, n19978, n19979, n19980, n19981,
    n19982, n19983, n19984, n19985, n19986, n19987,
    n19988, n19989, n19990, n19991, n19992, n19993,
    n19994, n19995, n19996, n19997, n19998, n19999,
    n20000, n20001, n20002, n20003, n20004, n20005,
    n20006, n20007, n20008, n20009, n20010, n20011,
    n20012, n20013, n20014, n20015, n20016, n20017,
    n20018, n20019, n20020, n20021, n20022, n20023,
    n20024, n20025, n20026, n20027, n20028, n20029,
    n20030, n20031, n20032, n20033, n20034, n20035,
    n20036, n20037, n20038, n20039, n20040, n20041,
    n20042, n20043, n20044, n20045, n20046, n20047,
    n20048, n20049, n20050, n20051, n20052, n20053,
    n20054, n20055, n20056, n20057, n20058, n20059,
    n20060, n20061, n20062, n20063, n20064, n20065,
    n20066, n20067, n20068, n20069, n20070, n20071,
    n20072, n20073, n20074, n20075, n20076, n20077,
    n20078, n20079, n20080, n20081, n20082, n20083,
    n20084, n20085, n20086, n20087, n20088, n20089,
    n20090, n20091, n20092, n20093, n20094, n20095,
    n20096, n20097, n20098, n20099, n20100, n20101,
    n20102, n20103, n20104, n20105, n20106, n20107,
    n20108, n20109, n20110, n20111, n20112, n20113,
    n20114, n20115, n20116, n20117, n20118, n20119,
    n20120, n20121, n20122, n20123, n20124, n20125,
    n20126, n20127, n20128, n20129, n20130, n20131,
    n20132, n20133, n20134, n20135, n20136, n20137,
    n20138, n20139, n20140, n20141, n20142, n20143,
    n20144, n20145, n20146, n20147, n20148, n20149,
    n20150, n20151, n20152, n20153, n20154, n20155,
    n20156, n20157, n20158, n20159, n20160, n20161,
    n20162, n20163, n20164, n20165, n20166, n20167,
    n20168, n20169, n20170, n20171, n20172, n20173,
    n20174, n20175, n20176, n20177, n20178, n20179,
    n20180, n20181, n20182, n20183, n20184, n20185,
    n20186, n20187, n20188, n20189, n20190, n20191,
    n20192, n20193, n20194, n20195, n20196, n20197,
    n20198, n20199, n20200, n20201, n20202, n20203,
    n20204, n20205, n20206, n20207, n20208, n20209,
    n20210, n20211, n20212, n20213, n20214, n20215,
    n20216, n20217, n20218, n20219, n20220, n20221,
    n20222, n20223, n20224, n20225, n20226, n20227,
    n20228, n20229, n20230, n20231, n20232, n20233,
    n20234, n20235, n20236, n20237, n20238, n20239,
    n20240, n20241, n20242, n20243, n20244, n20245,
    n20246, n20247, n20248, n20249, n20250, n20251,
    n20252, n20253, n20254, n20255, n20256, n20257,
    n20258, n20259, n20260, n20261, n20262, n20263,
    n20264, n20265, n20266, n20267, n20268, n20269,
    n20270, n20271, n20272, n20273, n20274, n20275,
    n20276, n20277, n20278, n20279, n20280, n20281,
    n20282, n20283, n20284, n20285, n20286, n20287,
    n20288, n20289, n20290, n20291, n20292, n20293,
    n20294, n20295, n20296, n20297, n20298, n20299,
    n20300, n20301, n20302, n20303, n20304, n20305,
    n20306, n20307, n20308, n20309, n20310, n20311,
    n20312, n20313, n20314, n20315, n20316, n20317,
    n20318, n20319, n20320, n20321, n20322, n20323,
    n20324, n20325, n20326, n20327, n20328, n20329,
    n20330, n20331, n20332, n20333, n20334, n20335,
    n20336, n20337, n20338, n20339, n20340, n20341,
    n20342, n20343, n20344, n20345, n20346, n20347,
    n20348, n20349, n20350, n20351, n20352, n20353,
    n20354, n20355, n20356, n20357, n20358, n20359,
    n20360, n20361, n20362, n20363, n20364, n20365,
    n20366, n20367, n20368, n20369, n20370, n20371,
    n20372, n20373, n20374, n20375, n20376, n20377,
    n20378, n20379, n20380, n20381, n20382, n20383,
    n20384, n20385, n20386, n20387, n20388, n20389,
    n20390, n20391, n20392, n20393, n20394, n20395,
    n20396, n20397, n20398, n20399, n20400, n20401,
    n20402, n20403, n20404, n20405, n20406, n20407,
    n20408, n20409, n20410, n20411, n20412, n20413,
    n20414, n20415, n20416, n20417, n20418, n20419,
    n20420, n20421, n20422, n20423, n20424, n20425,
    n20426, n20427, n20428, n20429, n20430, n20431,
    n20432, n20433, n20434, n20435, n20436, n20437,
    n20438, n20439, n20440, n20441, n20442, n20443,
    n20444, n20445, n20446, n20447, n20448, n20449,
    n20450, n20451, n20452, n20453, n20454, n20455,
    n20456, n20457, n20458, n20459, n20460, n20461,
    n20462, n20463, n20464, n20465, n20466, n20467,
    n20468, n20469, n20470, n20471, n20472, n20473,
    n20474, n20475, n20476, n20477, n20478, n20479,
    n20480, n20481, n20482, n20483, n20484, n20485,
    n20486, n20487, n20488, n20489, n20490, n20491,
    n20492, n20493, n20494, n20495, n20496, n20497,
    n20498, n20499, n20500, n20501, n20502, n20503,
    n20504, n20505, n20506, n20507, n20508, n20509,
    n20510, n20511, n20512, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521,
    n20522, n20523, n20524, n20525, n20526, n20527,
    n20528, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539,
    n20540, n20541, n20542, n20543, n20544, n20545,
    n20546, n20547, n20548, n20549, n20550, n20551,
    n20552, n20553, n20554, n20555, n20556, n20557,
    n20558, n20559, n20560, n20561, n20562, n20563,
    n20564, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581,
    n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599,
    n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617,
    n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20631, n20632, n20633, n20634, n20635,
    n20636, n20637, n20638, n20639, n20640, n20641,
    n20642, n20643, n20644, n20645, n20646, n20647,
    n20648, n20649, n20650, n20651, n20652, n20653,
    n20654, n20655, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665,
    n20666, n20667, n20668, n20669, n20670, n20671,
    n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683,
    n20684, n20685, n20686, n20687, n20688, n20689,
    n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701,
    n20702, n20703, n20704, n20705, n20706, n20707,
    n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719,
    n20720, n20721, n20722, n20723, n20724, n20725,
    n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737,
    n20738, n20739, n20740, n20741, n20742, n20743,
    n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755,
    n20756, n20757, n20758, n20759, n20760, n20761,
    n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773,
    n20774, n20775, n20776, n20777, n20778, n20779,
    n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20789, n20790, n20791,
    n20792, n20793, n20794, n20795, n20796, n20797,
    n20798, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809,
    n20810, n20811, n20812, n20813, n20814, n20815,
    n20816, n20817, n20818, n20819, n20820, n20821,
    n20822, n20823, n20824, n20825, n20826, n20827,
    n20828, n20829, n20830, n20831, n20832, n20833,
    n20834, n20835, n20836, n20837, n20838, n20839,
    n20840, n20841, n20842, n20843, n20844, n20845,
    n20846, n20847, n20848, n20849, n20850, n20851,
    n20852, n20853, n20854, n20855, n20856, n20857,
    n20858, n20859, n20860, n20861, n20862, n20863,
    n20864, n20865, n20866, n20867, n20868, n20869,
    n20870, n20871, n20872, n20873, n20874, n20875,
    n20876, n20877, n20878, n20879, n20880, n20881,
    n20882, n20883, n20884, n20885, n20886, n20887,
    n20888, n20889, n20890, n20891, n20892, n20893,
    n20894, n20895, n20896, n20897, n20898, n20899,
    n20900, n20901, n20902, n20903, n20904, n20905,
    n20906, n20907, n20908, n20909, n20910, n20911,
    n20912, n20913, n20914, n20915, n20916, n20917,
    n20918, n20919, n20920, n20921, n20922, n20923,
    n20924, n20925, n20926, n20927, n20928, n20929,
    n20930, n20931, n20932, n20933, n20934, n20935,
    n20936, n20937, n20938, n20939, n20940, n20941,
    n20942, n20943, n20944, n20945, n20946, n20947,
    n20948, n20949, n20950, n20951, n20952, n20953,
    n20954, n20955, n20956, n20957, n20958, n20959,
    n20960, n20961, n20962, n20963, n20964, n20965,
    n20966, n20967, n20968, n20969, n20970, n20971,
    n20972, n20973, n20974, n20975, n20976, n20977,
    n20978, n20979, n20980, n20981, n20982, n20983,
    n20984, n20985, n20986, n20987, n20988, n20989,
    n20990, n20991, n20992, n20993, n20994, n20995,
    n20996, n20997, n20998, n20999, n21000, n21001,
    n21002, n21003, n21004, n21005, n21006, n21007,
    n21008, n21009, n21010, n21011, n21012, n21013,
    n21014, n21015, n21016, n21017, n21018, n21019,
    n21020, n21021, n21022, n21023, n21024, n21025,
    n21026, n21027, n21028, n21029, n21030, n21031,
    n21032, n21033, n21034, n21035, n21036, n21037,
    n21038, n21039, n21040, n21041, n21042, n21043,
    n21044, n21045, n21046, n21047, n21048, n21049,
    n21050, n21051, n21052, n21053, n21054, n21055,
    n21056, n21057, n21058, n21059, n21060, n21061,
    n21062, n21063, n21064, n21065, n21066, n21067,
    n21068, n21069, n21070, n21071, n21072, n21073,
    n21074, n21075, n21076, n21077, n21078, n21079,
    n21080, n21081, n21082, n21083, n21084, n21085,
    n21086, n21087, n21088, n21089, n21090, n21091,
    n21092, n21093, n21094, n21095, n21096, n21097,
    n21098, n21099, n21100, n21101, n21102, n21103,
    n21104, n21105, n21106, n21107, n21108, n21109,
    n21110, n21111, n21112, n21113, n21114, n21115,
    n21116, n21117, n21118, n21119, n21120, n21121,
    n21122, n21123, n21124, n21125, n21126, n21127,
    n21128, n21129, n21130, n21131, n21132, n21133,
    n21134, n21135, n21136, n21137, n21138, n21139,
    n21140, n21141, n21142, n21143, n21144, n21145,
    n21146, n21147, n21148, n21149, n21150, n21151,
    n21152, n21153, n21154, n21155, n21156, n21157,
    n21158, n21159, n21160, n21161, n21162, n21163,
    n21164, n21165, n21166, n21167, n21168, n21169,
    n21170, n21171, n21172, n21173, n21174, n21175,
    n21176, n21177, n21178, n21179, n21180, n21181,
    n21182, n21183, n21184, n21185, n21186, n21187,
    n21188, n21189, n21190, n21191, n21192, n21193,
    n21194, n21195, n21196, n21197, n21198, n21199,
    n21200, n21201, n21202, n21203, n21204, n21205,
    n21206, n21207, n21208, n21209, n21210, n21211,
    n21212, n21213, n21214, n21215, n21216, n21217,
    n21218, n21219, n21220, n21221, n21222, n21223,
    n21224, n21225, n21226, n21227, n21228, n21229,
    n21230, n21231, n21232, n21233, n21234, n21235,
    n21236, n21237, n21238, n21239, n21240, n21241,
    n21242, n21243, n21244, n21245, n21246, n21247,
    n21248, n21249, n21250, n21251, n21252, n21253,
    n21254, n21255, n21256, n21257, n21258, n21259,
    n21260, n21261, n21262, n21263, n21264, n21265,
    n21266, n21267, n21268, n21269, n21270, n21271,
    n21272, n21273, n21274, n21275, n21276, n21277,
    n21278, n21279, n21280, n21281, n21282, n21283,
    n21284, n21285, n21286, n21287, n21288, n21289,
    n21290, n21291, n21292, n21293, n21294, n21295,
    n21296, n21297, n21298, n21299, n21300, n21301,
    n21302, n21303, n21304, n21305, n21306, n21307,
    n21308, n21309, n21310, n21311, n21312, n21313,
    n21314, n21315, n21316, n21317, n21318, n21319,
    n21320, n21321, n21322, n21323, n21324, n21325,
    n21326, n21327, n21328, n21329, n21330, n21331,
    n21332, n21333, n21334, n21335, n21336, n21337,
    n21338, n21339, n21340, n21341, n21342, n21343,
    n21344, n21345, n21346, n21347, n21348, n21349,
    n21350, n21351, n21352, n21353, n21354, n21355,
    n21356, n21357, n21358, n21359, n21360, n21361,
    n21362, n21363, n21364, n21365, n21366, n21367,
    n21368, n21369, n21370, n21371, n21372, n21373,
    n21374, n21375, n21376, n21377, n21378, n21379,
    n21380, n21381, n21382, n21383, n21384, n21385,
    n21386, n21387, n21388, n21389, n21390, n21391,
    n21392, n21393, n21394, n21395, n21396, n21397,
    n21398, n21399, n21400, n21401, n21402, n21403,
    n21404, n21405, n21406, n21407, n21408, n21409,
    n21410, n21411, n21412, n21413, n21414, n21415,
    n21416, n21417, n21418, n21419, n21420, n21421,
    n21422, n21423, n21424, n21425, n21426, n21427,
    n21428, n21429, n21430, n21431, n21432, n21433,
    n21434, n21435, n21436, n21437, n21438, n21439,
    n21440, n21441, n21442, n21443, n21444, n21445,
    n21446, n21447, n21448, n21449, n21450, n21451,
    n21452, n21453, n21454, n21455, n21456, n21457,
    n21458, n21459, n21460, n21461, n21462, n21463,
    n21464, n21465, n21466, n21467, n21468, n21469,
    n21470, n21471, n21472, n21473, n21474, n21475,
    n21476, n21477, n21478, n21479, n21480, n21481,
    n21482, n21483, n21484, n21485, n21486, n21487,
    n21488, n21489, n21490, n21491, n21492, n21493,
    n21494, n21495, n21496, n21497, n21498, n21499,
    n21500, n21501, n21502, n21503, n21504, n21505,
    n21506, n21507, n21508, n21509, n21510, n21511,
    n21512, n21513, n21514, n21515, n21516, n21517,
    n21518, n21519, n21520, n21521, n21522, n21523,
    n21524, n21525, n21526, n21527, n21528, n21529,
    n21530, n21531, n21532, n21533, n21534, n21535,
    n21536, n21537, n21538, n21539, n21540, n21541,
    n21542, n21543, n21544, n21545, n21546, n21547,
    n21548, n21549, n21550, n21551, n21552, n21553,
    n21554, n21555, n21556, n21557, n21558, n21559,
    n21560, n21561, n21562, n21563, n21564, n21565,
    n21566, n21567, n21568, n21569, n21570, n21571,
    n21572, n21573, n21574, n21575, n21576, n21577,
    n21578, n21579, n21580, n21581, n21582, n21583,
    n21584, n21585, n21586, n21587, n21588, n21589,
    n21590, n21591, n21592, n21593, n21594, n21595,
    n21596, n21597, n21598, n21599, n21600, n21601,
    n21602, n21603, n21604, n21605, n21606, n21607,
    n21608, n21609, n21610, n21611, n21612, n21613,
    n21614, n21615, n21616, n21617, n21618, n21619,
    n21620, n21621, n21622, n21623, n21624, n21625,
    n21626, n21627, n21628, n21629, n21630, n21631,
    n21632, n21633, n21634, n21635, n21636, n21637,
    n21638, n21639, n21640, n21641, n21642, n21643,
    n21644, n21645, n21646, n21647, n21648, n21649,
    n21650, n21651, n21652, n21653, n21654, n21655,
    n21656, n21657, n21658, n21659, n21660, n21661,
    n21662, n21663, n21664, n21665, n21666, n21667,
    n21668, n21669, n21670, n21671, n21672, n21673,
    n21674, n21675, n21676, n21677, n21678, n21679,
    n21680, n21681, n21682, n21683, n21684, n21685,
    n21686, n21687, n21688, n21689, n21690, n21691,
    n21692, n21693, n21694, n21695, n21696, n21697,
    n21698, n21699, n21700, n21701, n21702, n21703,
    n21704, n21705, n21706, n21707, n21708, n21709,
    n21710, n21711, n21712, n21713, n21714, n21715,
    n21716, n21717, n21718, n21719, n21720, n21721,
    n21722, n21723, n21724, n21725, n21726, n21727,
    n21728, n21729, n21730, n21731, n21732, n21733,
    n21734, n21735, n21736, n21737, n21738, n21739,
    n21740, n21741, n21742, n21743, n21744, n21745,
    n21746, n21747, n21748, n21749, n21750, n21751,
    n21752, n21753, n21754, n21755, n21756, n21757,
    n21758, n21759, n21760, n21761, n21762, n21763,
    n21764, n21765, n21766, n21767, n21768, n21769,
    n21770, n21771, n21772, n21773, n21774, n21775,
    n21776, n21777, n21778, n21779, n21780, n21781,
    n21782, n21783, n21784, n21785, n21786, n21787,
    n21788, n21789, n21790, n21791, n21792, n21793,
    n21794, n21795, n21796, n21797, n21798, n21799,
    n21800, n21801, n21802, n21803, n21804, n21805,
    n21806, n21807, n21808, n21809, n21810, n21811,
    n21812, n21813, n21814, n21815, n21816, n21817,
    n21818, n21819, n21820, n21821, n21822, n21823,
    n21824, n21825, n21826, n21827, n21828, n21829,
    n21830, n21831, n21832, n21833, n21834, n21835,
    n21836, n21837, n21838, n21839, n21840, n21841,
    n21842, n21843, n21844, n21845, n21846, n21847,
    n21848, n21849, n21850, n21851, n21852, n21853,
    n21854, n21855, n21856, n21857, n21858, n21859,
    n21860, n21861, n21862, n21863, n21864, n21865,
    n21866, n21867, n21868, n21869, n21870, n21871,
    n21872, n21873, n21874, n21875, n21876, n21877,
    n21878, n21879, n21880, n21881, n21882, n21883,
    n21884, n21885, n21886, n21887, n21888, n21889,
    n21890, n21891, n21892, n21893, n21894, n21895,
    n21896, n21897, n21898, n21899, n21900, n21901,
    n21902, n21903, n21904, n21905, n21906, n21907,
    n21908, n21909, n21910, n21911, n21912, n21913,
    n21914, n21915, n21916, n21917, n21918, n21919,
    n21920, n21921, n21922, n21923, n21924, n21925,
    n21926, n21927, n21928, n21929, n21930, n21931,
    n21932, n21933, n21934, n21935, n21936, n21937,
    n21938, n21939, n21940, n21941, n21942, n21943,
    n21944, n21945, n21946, n21947, n21948, n21949,
    n21950, n21951, n21952, n21953, n21954, n21955,
    n21956, n21957, n21958, n21959, n21960, n21961,
    n21962, n21963, n21964, n21965, n21966, n21967,
    n21968, n21969, n21970, n21971, n21972, n21973,
    n21974, n21975, n21976, n21977, n21978, n21979,
    n21980, n21981, n21982, n21983, n21984, n21985,
    n21986, n21987, n21988, n21989, n21990, n21991,
    n21992, n21993, n21994, n21995, n21996, n21997,
    n21998, n21999, n22000, n22001, n22002, n22003,
    n22004, n22005, n22006, n22007, n22008, n22009,
    n22010, n22011, n22012, n22013, n22014, n22015,
    n22016, n22017, n22018, n22019, n22020, n22021,
    n22022, n22023, n22024, n22025, n22026, n22027,
    n22028, n22029, n22030, n22031, n22032, n22033,
    n22034, n22035, n22036, n22037, n22038, n22039,
    n22040, n22041, n22042, n22043, n22044, n22045,
    n22046, n22047, n22048, n22049, n22050, n22051,
    n22052, n22053, n22054, n22055, n22056, n22057,
    n22058, n22059, n22060, n22061, n22062, n22063,
    n22064, n22065, n22066, n22067, n22068, n22069,
    n22070, n22071, n22072, n22073, n22074, n22075,
    n22076, n22077, n22078, n22079, n22080, n22081,
    n22082, n22083, n22084, n22085, n22086, n22087,
    n22088, n22089, n22090, n22091, n22092, n22093,
    n22094, n22095, n22096, n22097, n22098, n22099,
    n22100, n22101, n22102, n22103, n22104, n22105,
    n22106, n22107, n22108, n22109, n22110, n22111,
    n22112, n22113, n22114, n22115, n22116, n22117,
    n22118, n22119, n22120, n22121, n22122, n22123,
    n22124, n22125, n22126, n22127, n22128, n22129,
    n22130, n22131, n22132, n22133, n22134, n22135,
    n22136, n22137, n22138, n22139, n22140, n22141,
    n22142, n22143, n22144, n22145, n22146, n22147,
    n22148, n22149, n22150, n22151, n22152, n22153,
    n22154, n22155, n22156, n22157, n22158, n22159,
    n22160, n22161, n22162, n22163, n22164, n22165,
    n22166, n22167, n22168, n22169, n22170, n22171,
    n22172, n22173, n22174, n22175, n22176, n22177,
    n22178, n22179, n22180, n22181, n22182, n22183,
    n22184, n22185, n22186, n22187, n22188, n22189,
    n22190, n22191, n22192, n22193, n22194, n22195,
    n22196, n22197, n22198, n22199, n22200, n22201,
    n22202, n22203, n22204, n22205, n22206, n22207,
    n22208, n22209, n22210, n22211, n22212, n22213,
    n22214, n22215, n22216, n22217, n22218, n22219,
    n22220, n22221, n22222, n22223, n22224, n22225,
    n22226, n22227, n22228, n22229, n22230, n22231,
    n22232, n22233, n22234, n22235, n22236, n22237,
    n22238, n22239, n22240, n22241, n22242, n22243,
    n22244, n22245, n22246, n22247, n22248, n22249,
    n22250, n22251, n22252, n22253, n22254, n22255,
    n22256, n22257, n22258, n22259, n22260, n22261,
    n22262, n22263, n22264, n22265, n22266, n22267,
    n22268, n22269, n22270, n22271, n22272, n22273,
    n22274, n22275, n22276, n22277, n22278, n22279,
    n22280, n22281, n22282, n22283, n22284, n22285,
    n22286, n22287, n22288, n22289, n22290, n22291,
    n22292, n22293, n22294, n22295, n22296, n22297,
    n22298, n22299, n22300, n22301, n22302, n22303,
    n22304, n22305, n22306, n22307, n22308, n22309,
    n22310, n22311, n22312, n22313, n22314, n22315,
    n22316, n22317, n22318, n22319, n22320, n22321,
    n22322, n22323, n22324, n22325, n22326, n22327,
    n22328, n22329, n22330, n22331, n22332, n22333,
    n22334, n22335, n22336, n22337, n22338, n22339,
    n22340, n22341, n22342, n22343, n22344, n22345,
    n22346, n22347, n22348, n22349, n22350, n22351,
    n22352, n22353, n22354, n22355, n22356, n22357,
    n22358, n22359, n22360, n22361, n22362, n22363,
    n22364, n22365, n22366, n22367, n22368, n22369,
    n22370, n22371, n22372, n22373, n22374, n22375,
    n22376, n22377, n22378, n22379, n22380, n22381,
    n22382, n22383, n22384, n22385, n22386, n22387,
    n22388, n22389, n22390, n22391, n22392, n22393,
    n22394, n22395, n22396, n22397, n22398, n22399,
    n22400, n22401, n22402, n22403, n22404, n22405,
    n22406, n22407, n22408, n22409, n22410, n22411,
    n22412, n22413, n22414, n22415, n22416, n22417,
    n22418, n22419, n22420, n22421, n22422, n22423,
    n22424, n22425, n22426, n22427, n22428, n22429,
    n22430, n22431, n22432, n22433, n22434, n22435,
    n22436, n22437, n22438, n22439, n22440, n22441,
    n22442, n22443, n22444, n22445, n22446, n22447,
    n22448, n22449, n22450, n22451, n22452, n22453,
    n22454, n22455, n22456, n22457, n22458, n22459,
    n22460, n22461, n22462, n22463, n22464, n22465,
    n22466, n22467, n22468, n22469, n22470, n22471,
    n22472, n22473, n22474, n22475, n22476, n22477,
    n22478, n22479, n22480, n22481, n22482, n22483,
    n22484, n22485, n22486, n22487, n22488, n22489,
    n22490, n22491, n22492, n22493, n22494, n22495,
    n22496, n22497, n22498, n22499, n22500, n22501,
    n22502, n22503, n22504, n22505, n22506, n22507,
    n22508, n22509, n22510, n22511, n22512, n22513,
    n22514, n22515, n22516, n22517, n22518, n22519,
    n22520, n22521, n22522, n22523, n22524, n22525,
    n22526, n22527, n22528, n22529, n22530, n22531,
    n22532, n22533, n22534, n22535, n22536, n22537,
    n22538, n22539, n22540, n22541, n22542, n22543,
    n22544, n22545, n22546, n22547, n22548, n22549,
    n22550, n22551, n22552, n22553, n22554, n22555,
    n22556, n22557, n22558, n22559, n22560, n22561,
    n22562, n22563, n22564, n22565, n22566, n22567,
    n22568, n22569, n22570, n22571, n22572, n22573,
    n22574, n22575, n22576, n22577, n22578, n22579,
    n22580, n22581, n22582, n22583, n22584, n22585,
    n22586, n22587, n22588, n22589, n22590, n22591,
    n22592, n22593, n22594, n22595, n22596, n22597,
    n22598, n22599, n22600, n22601, n22602, n22603,
    n22604, n22605, n22606, n22607, n22608, n22609,
    n22610, n22611, n22612, n22613, n22614, n22615,
    n22616, n22617, n22618, n22619, n22620, n22621,
    n22622, n22623, n22624, n22625, n22626, n22627,
    n22628, n22629, n22630, n22631, n22632, n22633,
    n22634, n22635, n22636, n22637, n22638, n22639,
    n22640, n22641, n22642, n22643, n22644, n22645,
    n22646, n22647, n22648, n22649, n22650, n22651,
    n22652, n22653, n22654, n22655, n22656, n22657,
    n22658, n22659, n22660, n22661, n22662, n22663,
    n22664, n22665, n22666, n22667, n22668, n22669,
    n22670, n22671, n22672, n22673, n22674, n22675,
    n22676, n22677, n22678, n22679, n22680, n22681,
    n22682, n22683, n22684, n22685, n22686, n22687,
    n22688, n22689, n22690, n22691, n22692, n22693,
    n22694, n22695, n22696, n22697, n22698, n22699,
    n22700, n22701, n22702, n22703, n22704, n22705,
    n22706, n22707, n22708, n22709, n22710, n22711,
    n22712, n22713, n22714, n22715, n22716, n22717,
    n22718, n22719, n22720, n22721, n22722, n22723,
    n22724, n22725, n22726, n22727, n22728, n22729,
    n22730, n22731, n22732, n22733, n22734, n22735,
    n22736, n22737, n22738, n22739, n22740, n22741,
    n22742, n22743, n22744, n22745, n22746, n22747,
    n22748, n22749, n22750, n22751, n22752, n22753,
    n22754, n22755, n22756, n22757, n22758, n22759,
    n22760, n22761, n22762, n22763, n22764, n22765,
    n22766, n22767, n22768, n22769, n22770, n22771,
    n22772, n22773, n22774, n22775, n22776, n22777,
    n22778, n22779, n22780, n22781, n22782, n22783,
    n22784, n22785, n22786, n22787, n22788, n22789,
    n22790, n22791, n22792, n22793, n22794, n22795,
    n22796, n22797, n22798, n22799, n22800, n22801,
    n22802, n22803, n22804, n22805, n22806, n22807,
    n22808, n22809, n22810, n22811, n22812, n22813,
    n22814, n22815, n22816, n22817, n22818, n22819,
    n22820, n22821, n22822, n22823, n22824, n22825,
    n22826, n22827, n22828, n22829, n22830, n22831,
    n22832, n22833, n22834, n22835, n22836, n22837,
    n22838, n22839, n22840, n22841, n22842, n22843,
    n22844, n22845, n22846, n22847, n22848, n22849,
    n22850, n22851, n22852, n22853, n22854, n22855,
    n22856, n22857, n22858, n22859, n22860, n22861,
    n22862, n22863, n22864, n22865, n22866, n22867,
    n22868, n22869, n22870, n22871, n22872, n22873,
    n22874, n22875, n22876, n22877, n22878, n22879,
    n22880, n22881, n22882, n22883, n22884, n22885,
    n22886, n22887, n22888, n22889, n22890, n22891,
    n22892, n22893, n22894, n22895, n22896, n22897,
    n22898, n22899, n22900, n22901, n22902, n22903,
    n22904, n22905, n22906, n22907, n22908, n22909,
    n22910, n22911, n22912, n22913, n22914, n22915,
    n22916, n22917, n22918, n22919, n22920, n22921,
    n22922, n22923, n22924, n22925, n22926, n22927,
    n22928, n22929, n22930, n22931, n22932, n22933,
    n22934, n22935, n22936, n22937, n22938, n22939,
    n22940, n22941, n22942, n22943, n22944, n22945,
    n22946, n22947, n22948, n22949, n22950, n22951,
    n22952, n22953, n22954, n22955, n22956, n22957,
    n22958, n22959, n22960, n22961, n22962, n22963,
    n22964, n22965, n22966, n22967, n22968, n22969,
    n22970, n22971, n22972, n22973, n22974, n22975,
    n22976, n22977, n22978, n22979, n22980, n22981,
    n22982, n22983, n22984, n22985, n22986, n22987,
    n22988, n22989, n22990, n22991, n22992, n22993,
    n22994, n22995, n22996, n22997, n22998, n22999,
    n23000, n23001, n23002, n23003, n23004, n23005,
    n23006, n23007, n23008, n23009, n23010, n23011,
    n23012, n23013, n23014, n23015, n23016, n23017,
    n23018, n23019, n23020, n23021, n23022, n23023,
    n23024, n23025, n23026, n23027, n23028, n23029,
    n23030, n23031, n23032, n23033, n23034, n23035,
    n23036, n23037, n23038, n23039, n23040, n23041,
    n23042, n23043, n23044, n23045, n23046, n23047,
    n23048, n23049, n23050, n23051, n23052, n23053,
    n23054, n23055, n23056, n23057, n23058, n23059,
    n23060, n23061, n23062, n23063, n23064, n23065,
    n23066, n23067, n23068, n23069, n23070, n23071,
    n23072, n23073, n23074, n23075, n23076, n23077,
    n23078, n23079, n23080, n23081, n23082, n23083,
    n23084, n23085, n23086, n23087, n23088, n23089,
    n23090, n23091, n23092, n23093, n23094, n23095,
    n23096, n23097, n23098, n23099, n23100, n23101,
    n23102, n23103, n23104, n23105, n23106, n23107,
    n23108, n23109, n23110, n23111, n23112, n23113,
    n23114, n23115, n23116, n23117, n23118, n23119,
    n23120, n23121, n23122, n23123, n23124, n23125,
    n23126, n23127, n23128, n23129, n23130, n23131,
    n23132, n23133, n23134, n23135, n23136, n23137,
    n23138, n23139, n23140, n23141, n23142, n23143,
    n23144, n23145, n23146, n23147, n23148, n23149,
    n23150, n23151, n23152, n23153, n23154, n23155,
    n23156, n23157, n23158, n23159, n23160, n23161,
    n23162, n23163, n23164, n23165, n23166, n23167,
    n23168, n23169, n23170, n23171, n23172, n23173,
    n23174, n23175, n23176, n23177, n23178, n23179,
    n23180, n23181, n23182, n23183, n23184, n23185,
    n23186, n23187, n23188, n23189, n23190, n23191,
    n23192, n23193, n23194, n23195, n23196, n23197,
    n23198, n23199, n23200, n23201, n23202, n23203,
    n23204, n23205, n23206, n23207, n23208, n23209,
    n23210, n23211, n23212, n23213, n23214, n23215,
    n23216, n23217, n23218, n23219, n23220, n23221,
    n23222, n23223, n23224, n23225, n23226, n23227,
    n23228, n23229, n23230, n23231, n23232, n23233,
    n23234, n23235, n23236, n23237, n23238, n23239,
    n23240, n23241, n23242, n23243, n23244, n23245,
    n23246, n23247, n23248, n23249, n23250, n23251,
    n23252, n23253, n23254, n23255, n23256, n23257,
    n23258, n23259, n23260, n23261, n23262, n23263,
    n23264, n23265, n23266, n23267, n23268, n23269,
    n23270, n23271, n23272, n23273, n23274, n23275,
    n23276, n23277, n23278, n23279, n23280, n23281,
    n23282, n23283, n23284, n23285, n23286, n23287,
    n23288, n23289, n23290, n23291, n23292, n23293,
    n23294, n23295, n23296, n23297, n23298, n23299,
    n23300, n23301, n23302, n23303, n23304, n23305,
    n23306, n23307, n23308, n23309, n23310, n23311,
    n23312, n23313, n23314, n23315, n23316, n23317,
    n23318, n23319, n23320, n23321, n23322, n23323,
    n23324, n23325, n23326, n23327, n23328, n23329,
    n23330, n23331, n23332, n23333, n23334, n23335,
    n23336, n23337, n23338, n23339, n23340, n23341,
    n23342, n23343, n23344, n23345, n23346, n23347,
    n23348, n23349, n23350, n23351, n23352, n23353,
    n23354, n23355, n23356, n23357, n23358, n23359,
    n23360, n23361, n23362, n23363, n23364, n23365,
    n23366, n23367, n23368, n23369, n23370, n23371,
    n23372, n23373, n23374, n23375, n23376, n23377,
    n23378, n23379, n23380, n23381, n23382, n23383,
    n23384, n23385, n23386, n23387, n23388, n23389,
    n23390, n23391, n23392, n23393, n23394, n23395,
    n23396, n23397, n23398, n23399, n23400, n23401,
    n23402, n23403, n23404, n23405, n23406, n23407,
    n23408, n23409, n23410, n23411, n23412, n23413,
    n23414, n23415, n23416, n23417, n23418, n23419,
    n23420, n23421, n23422, n23423, n23424, n23425,
    n23426, n23427, n23428, n23429, n23430, n23431,
    n23432, n23433, n23434, n23435, n23436, n23437,
    n23438, n23439, n23440, n23441, n23442, n23443,
    n23444, n23445, n23446, n23447, n23448, n23449,
    n23450, n23451, n23452, n23453, n23454, n23455,
    n23456, n23457, n23458, n23459, n23460, n23461,
    n23462, n23463, n23464, n23465, n23466, n23467,
    n23468, n23469, n23470, n23471, n23472, n23473,
    n23474, n23475, n23476, n23477, n23478, n23479,
    n23480, n23481, n23482, n23483, n23484, n23485,
    n23486, n23487, n23488, n23489, n23490, n23491,
    n23492, n23493, n23494, n23495, n23496, n23497,
    n23498, n23499, n23500, n23501, n23502, n23503,
    n23504, n23505, n23506, n23507, n23508, n23509,
    n23510, n23511, n23512, n23513, n23514, n23515,
    n23516, n23517, n23518, n23519, n23520, n23521,
    n23522, n23523, n23524, n23525, n23526, n23527,
    n23528, n23529, n23530, n23531, n23532, n23533,
    n23534, n23535, n23536, n23537, n23538, n23539,
    n23540, n23541, n23542, n23543, n23544, n23545,
    n23546, n23547, n23548, n23549, n23550, n23551,
    n23552, n23553, n23554, n23555, n23556, n23557,
    n23558, n23559, n23560, n23561, n23562, n23563,
    n23564, n23565, n23566, n23567, n23568, n23569,
    n23570, n23571, n23572, n23573, n23574, n23575,
    n23576, n23577, n23578, n23579, n23580, n23581,
    n23582, n23583, n23584, n23585, n23586, n23587,
    n23588, n23589, n23590, n23591, n23592, n23593,
    n23594, n23595, n23596, n23597, n23598, n23599,
    n23600, n23601, n23602, n23603, n23604, n23605,
    n23606, n23607, n23608, n23609, n23610, n23611,
    n23612, n23613, n23614, n23615, n23616, n23617,
    n23618, n23619, n23620, n23621, n23622, n23623,
    n23624, n23625, n23626, n23627, n23628, n23629,
    n23630, n23631, n23632, n23633, n23634, n23635,
    n23636, n23637, n23638, n23639, n23640, n23641,
    n23642, n23643, n23644, n23645, n23646, n23647,
    n23648, n23649, n23650, n23651, n23652, n23653,
    n23654, n23655, n23656, n23657, n23658, n23659,
    n23660, n23661, n23662, n23663, n23664, n23665,
    n23666, n23667, n23668, n23669, n23670, n23671,
    n23672, n23673, n23674, n23675, n23676, n23677,
    n23678, n23679, n23680, n23681, n23682, n23683,
    n23684, n23685, n23686, n23687, n23688, n23689,
    n23690, n23691, n23692, n23693, n23694, n23695,
    n23696, n23697, n23698, n23699, n23700, n23701,
    n23702, n23703, n23704, n23705, n23706, n23707,
    n23708, n23709, n23710, n23711, n23712, n23713,
    n23714, n23715, n23716, n23717, n23718, n23719,
    n23720, n23721, n23722, n23723, n23724, n23725,
    n23726, n23727, n23728, n23729, n23730, n23731,
    n23732, n23733, n23734, n23735, n23736, n23737,
    n23738, n23739, n23740, n23741, n23742, n23743,
    n23744, n23745, n23746, n23747, n23748, n23749,
    n23750, n23751, n23752, n23753, n23754, n23755,
    n23756, n23757, n23758, n23759, n23760, n23761,
    n23762, n23763, n23764, n23765, n23766, n23767,
    n23768, n23769, n23770, n23771, n23772, n23773,
    n23774, n23775, n23776, n23777, n23778, n23779,
    n23780, n23781, n23782, n23783, n23784, n23785,
    n23786, n23787, n23788, n23789, n23790, n23791,
    n23792, n23793, n23794, n23795, n23796, n23797,
    n23798, n23799, n23800, n23801, n23802, n23803,
    n23804, n23805, n23806, n23807, n23808, n23809,
    n23810, n23811, n23812, n23813, n23814, n23815,
    n23816, n23817, n23818, n23819, n23820, n23821,
    n23822, n23823, n23824, n23825, n23826, n23827,
    n23828, n23829, n23830, n23831, n23832, n23833,
    n23834, n23835, n23836, n23837, n23838, n23839,
    n23840, n23841, n23842, n23843, n23844, n23845,
    n23846, n23847, n23848, n23849, n23850, n23851,
    n23852, n23853, n23854, n23855, n23856, n23857,
    n23858, n23859, n23860, n23861, n23862, n23863,
    n23864, n23865, n23866, n23867, n23868, n23869,
    n23870, n23871, n23872, n23873, n23874, n23875,
    n23876, n23877, n23878, n23879, n23880, n23881,
    n23882, n23883, n23884, n23885, n23886, n23887,
    n23888, n23889, n23890, n23891, n23892, n23893,
    n23894, n23895, n23896, n23897, n23898, n23899,
    n23900, n23901, n23902, n23903, n23904, n23905,
    n23906, n23907, n23908, n23909, n23910, n23911,
    n23912, n23913, n23914, n23915, n23916, n23917,
    n23918, n23919, n23920, n23921, n23922, n23923,
    n23924, n23925, n23926, n23927, n23928, n23929,
    n23930, n23931, n23932, n23933, n23934, n23935,
    n23936, n23937, n23938, n23939, n23940, n23941,
    n23942, n23943, n23944, n23945, n23946, n23947,
    n23948, n23949, n23950, n23951, n23952, n23953,
    n23954, n23955, n23956, n23957, n23958, n23959,
    n23960, n23961, n23962, n23963, n23964, n23965,
    n23966, n23967, n23968, n23969, n23970, n23971,
    n23972, n23973, n23974, n23975, n23976, n23977,
    n23978, n23979, n23980, n23981, n23982, n23983,
    n23984, n23985, n23986, n23987, n23988, n23989,
    n23990, n23991, n23992, n23993, n23994, n23995,
    n23996, n23997, n23998, n23999, n24000, n24001,
    n24002, n24003, n24004, n24005, n24006, n24007,
    n24008, n24009, n24010, n24011, n24012, n24013,
    n24014, n24015, n24016, n24017, n24018, n24019,
    n24020, n24021, n24022, n24023, n24024, n24025,
    n24026, n24027, n24028, n24029, n24030, n24031,
    n24032, n24033, n24034, n24035, n24036, n24037,
    n24038, n24039, n24040, n24041, n24042, n24043,
    n24044, n24045, n24046, n24047, n24048, n24049,
    n24050, n24051, n24052, n24053, n24054, n24055,
    n24056, n24057, n24058, n24059, n24060, n24061,
    n24062, n24063, n24064, n24065, n24066, n24067,
    n24068, n24069, n24070, n24071, n24072, n24073,
    n24074, n24075, n24076, n24077, n24078, n24079,
    n24080, n24081, n24082, n24083, n24084, n24085,
    n24086, n24087, n24088, n24089, n24090, n24091,
    n24092, n24093, n24094, n24095, n24096, n24097,
    n24098, n24099, n24100, n24101, n24102, n24103,
    n24104, n24105, n24106, n24107, n24108, n24109,
    n24110, n24111, n24112, n24113, n24114, n24115,
    n24116, n24117, n24118, n24119, n24120, n24121,
    n24122, n24123, n24124, n24125, n24126, n24127,
    n24128, n24129, n24130, n24131, n24132, n24133,
    n24134, n24135, n24136, n24137, n24138, n24139,
    n24140, n24141, n24142, n24143, n24144, n24145,
    n24146, n24147, n24148, n24149, n24150, n24151,
    n24152, n24153, n24154, n24155, n24156, n24157,
    n24158, n24159, n24160, n24161, n24162, n24163,
    n24164, n24165, n24166, n24167, n24168, n24169,
    n24170, n24171, n24172, n24173, n24174, n24175,
    n24176, n24177, n24178, n24179, n24180, n24181,
    n24182, n24183, n24184, n24185, n24186, n24187,
    n24188, n24189, n24190, n24191, n24192, n24193,
    n24194, n24195, n24196, n24197, n24198, n24199,
    n24200, n24201, n24202, n24203, n24204, n24205,
    n24206, n24207, n24208, n24209, n24210, n24211,
    n24212, n24213, n24214, n24215, n24216, n24217,
    n24218, n24219, n24220, n24221, n24222, n24223,
    n24224, n24225, n24226, n24227, n24228, n24229,
    n24230, n24231, n24232, n24233, n24234, n24235,
    n24236, n24237, n24238, n24239, n24240, n24241,
    n24242, n24243, n24244, n24245, n24246, n24247,
    n24248, n24249, n24250, n24251, n24252, n24253,
    n24254, n24255, n24256, n24257, n24258, n24259,
    n24260, n24261, n24262, n24263, n24264, n24265,
    n24266, n24267, n24268, n24269, n24270, n24271,
    n24272, n24273, n24274, n24275, n24276, n24277,
    n24278, n24279, n24280, n24281, n24282, n24283,
    n24284, n24285, n24286, n24287, n24288, n24289,
    n24290, n24291, n24292, n24293, n24294, n24295,
    n24296, n24297, n24298, n24299, n24300, n24301,
    n24302, n24303, n24304, n24305, n24306, n24307,
    n24308, n24309, n24310, n24311, n24312, n24313,
    n24314, n24315, n24316, n24317, n24318, n24319,
    n24320, n24321, n24322, n24323, n24324, n24325,
    n24326, n24327, n24328, n24329, n24330, n24331,
    n24332, n24333, n24334, n24335, n24336, n24337,
    n24338, n24339, n24340, n24341, n24342, n24343,
    n24344, n24345, n24346, n24347, n24348, n24349,
    n24350, n24351, n24352, n24353, n24354, n24355,
    n24356, n24357, n24358, n24359, n24360, n24361,
    n24362, n24363, n24364, n24365, n24366, n24367,
    n24368, n24369, n24370, n24371, n24372, n24373,
    n24374, n24375, n24376, n24377, n24378, n24379,
    n24380, n24381, n24382, n24383, n24384, n24385,
    n24386, n24387, n24388, n24389, n24390, n24391,
    n24392, n24393, n24394, n24395, n24396, n24397,
    n24398, n24399, n24400, n24401, n24402, n24403,
    n24404, n24405, n24406, n24407, n24408, n24409,
    n24410, n24411, n24412, n24413, n24414, n24415,
    n24416, n24417, n24418, n24419, n24420, n24421,
    n24422, n24423, n24424, n24425, n24426, n24427,
    n24428, n24429, n24430, n24431, n24432, n24433,
    n24434, n24435, n24436, n24437, n24438, n24439,
    n24440, n24441, n24442, n24443, n24444, n24445,
    n24446, n24447, n24448, n24449, n24450, n24451,
    n24452, n24453, n24454, n24455, n24456, n24457,
    n24458, n24459, n24460, n24461, n24462, n24463,
    n24464, n24465, n24466, n24467, n24468, n24469,
    n24470, n24471, n24472, n24473, n24474, n24475,
    n24476, n24477, n24478, n24479, n24480, n24481,
    n24482, n24483, n24484, n24485, n24486, n24487,
    n24488, n24489, n24490, n24491, n24492, n24493,
    n24494, n24495, n24496, n24497, n24498, n24499,
    n24500, n24501, n24502, n24503, n24504, n24505,
    n24506, n24507, n24508, n24509, n24510, n24511,
    n24512, n24513, n24514, n24515, n24516, n24517,
    n24518, n24519, n24520, n24521, n24522, n24523,
    n24524, n24525, n24526, n24527, n24528, n24529,
    n24530, n24531, n24532, n24533, n24534, n24535,
    n24536, n24537, n24538, n24539, n24540, n24541,
    n24542, n24543, n24544, n24545, n24546, n24547,
    n24548, n24549, n24550, n24551, n24552, n24553,
    n24554, n24555, n24556, n24557, n24558, n24559,
    n24560, n24561, n24562, n24563, n24564, n24565,
    n24566, n24567, n24568, n24569, n24570, n24571,
    n24572, n24573, n24574, n24575, n24576, n24577,
    n24578, n24579, n24580, n24581, n24582, n24583,
    n24584, n24585, n24586, n24587, n24588, n24589,
    n24590, n24591, n24592, n24593, n24594, n24595,
    n24596, n24597, n24598, n24599, n24600, n24601,
    n24602, n24603, n24604, n24605, n24606, n24607,
    n24608, n24609, n24610, n24611, n24612, n24613,
    n24614, n24615, n24616, n24617, n24618, n24619,
    n24620, n24621, n24622, n24623, n24624, n24625,
    n24626, n24627, n24628, n24629, n24630, n24631,
    n24632, n24633, n24634, n24635, n24636, n24637,
    n24638, n24639, n24640, n24641, n24642, n24643,
    n24644, n24645, n24646, n24647, n24648, n24649,
    n24650, n24651, n24652, n24653, n24654, n24655,
    n24656, n24657, n24658, n24659, n24660, n24661,
    n24662, n24663, n24664, n24665, n24666, n24667,
    n24668, n24669, n24670, n24671, n24672, n24673,
    n24674, n24675, n24676, n24677, n24678, n24679,
    n24680, n24681, n24682, n24683, n24684, n24685,
    n24686, n24687, n24688, n24689, n24690, n24691,
    n24692, n24693, n24694, n24695, n24696, n24697,
    n24698, n24699, n24700, n24701, n24702, n24703,
    n24704, n24705, n24706, n24707, n24708, n24709,
    n24710, n24711, n24712, n24713, n24714, n24715,
    n24716, n24717, n24718, n24719, n24720, n24721,
    n24722, n24723, n24724, n24725, n24726, n24727,
    n24728, n24729, n24730, n24731, n24732, n24733,
    n24734, n24735, n24736, n24737, n24738, n24739,
    n24740, n24741, n24742, n24743, n24744, n24745,
    n24746, n24747, n24748, n24749, n24750, n24751,
    n24752, n24753, n24754, n24755, n24756, n24757,
    n24758, n24759, n24760, n24761, n24762, n24763,
    n24764, n24765, n24766, n24767, n24768, n24769,
    n24770, n24771, n24772, n24773, n24774, n24775,
    n24776, n24777, n24778, n24779, n24780, n24781,
    n24782, n24783, n24784, n24785, n24786, n24787,
    n24788, n24789, n24790, n24791, n24792, n24793,
    n24794, n24795, n24796, n24797, n24798, n24799,
    n24800, n24801, n24802, n24803, n24804, n24805,
    n24806, n24807, n24808, n24809, n24810, n24811,
    n24812, n24813, n24814, n24815, n24816, n24817,
    n24818, n24819, n24820, n24821, n24822, n24823,
    n24824, n24825, n24826, n24827, n24828, n24829,
    n24830, n24831, n24832, n24833, n24834, n24835,
    n24836, n24837, n24838, n24839, n24840, n24841,
    n24842, n24843, n24844, n24845, n24846, n24847,
    n24848, n24849, n24850, n24851, n24852, n24853,
    n24854, n24855, n24856, n24857, n24858, n24859,
    n24860, n24861, n24862, n24863, n24864, n24865,
    n24866, n24867, n24868, n24869, n24870, n24871,
    n24872, n24873, n24874, n24875, n24876, n24877,
    n24878, n24879, n24880, n24881, n24882, n24883,
    n24884, n24885, n24886, n24887, n24888, n24889,
    n24890, n24891, n24892, n24893, n24894, n24895,
    n24896, n24897, n24898, n24899, n24900, n24901,
    n24902, n24903, n24904, n24905, n24906, n24907,
    n24908, n24909, n24910, n24911, n24912, n24913,
    n24914, n24915, n24916, n24917, n24918, n24919,
    n24920, n24921, n24922, n24923, n24924, n24925,
    n24926, n24927, n24928, n24929, n24930, n24931,
    n24932, n24933, n24934, n24935, n24936, n24937,
    n24938, n24939, n24940, n24941, n24942, n24943,
    n24944, n24945, n24946, n24947, n24948, n24949,
    n24950, n24951, n24952, n24953, n24954, n24955,
    n24956, n24957, n24958, n24959, n24960, n24961,
    n24962, n24963, n24964, n24965, n24966, n24967,
    n24968, n24969, n24970, n24971, n24972, n24973,
    n24974, n24975, n24976, n24977, n24978, n24979,
    n24980, n24981, n24982, n24983, n24984, n24985,
    n24986, n24987, n24988, n24989, n24990, n24991,
    n24992, n24993, n24994, n24995, n24996, n24997,
    n24998, n24999, n25000, n25001, n25002, n25003,
    n25004, n25005, n25006, n25007, n25008, n25009,
    n25010, n25011, n25012, n25013, n25014, n25015,
    n25016, n25017, n25018, n25019, n25020, n25021,
    n25022, n25023, n25024, n25025, n25026, n25027,
    n25028, n25029, n25030, n25031, n25032, n25033,
    n25034, n25035, n25036, n25037, n25038, n25039,
    n25040, n25041, n25042, n25043, n25044, n25045,
    n25046, n25047, n25048, n25049, n25050, n25051,
    n25052, n25053, n25054, n25055, n25056, n25057,
    n25058, n25059, n25060, n25061, n25062, n25063,
    n25064, n25065, n25066, n25067, n25068, n25069,
    n25070, n25071, n25072, n25073, n25074, n25075,
    n25076, n25077, n25078, n25079, n25080, n25081,
    n25082, n25083, n25084, n25085, n25086, n25087,
    n25088, n25089, n25090, n25091, n25092, n25093,
    n25094, n25095, n25096, n25097, n25098, n25099,
    n25100, n25101, n25102, n25103, n25104, n25105,
    n25106, n25107, n25108, n25109, n25110, n25111,
    n25112, n25113, n25114, n25115, n25116, n25117,
    n25118, n25119, n25120, n25121, n25122, n25123,
    n25124, n25125, n25126, n25127, n25128, n25129,
    n25130, n25131, n25132, n25133, n25134, n25135,
    n25136, n25137, n25138, n25139, n25140, n25141,
    n25142, n25143, n25144, n25145, n25146, n25147,
    n25148, n25149, n25150, n25151, n25152, n25153,
    n25154, n25155, n25156, n25157, n25158, n25159,
    n25160, n25161, n25162, n25163, n25164, n25165,
    n25166, n25167, n25168, n25169, n25170, n25171,
    n25172, n25173, n25174, n25175, n25176, n25177,
    n25178, n25179, n25180, n25181, n25182, n25183,
    n25184, n25185, n25186, n25187, n25188, n25189,
    n25190, n25191, n25192, n25193, n25194, n25195,
    n25196, n25197, n25198, n25199, n25200, n25201,
    n25202, n25203, n25204, n25205, n25206, n25207,
    n25208, n25209, n25210, n25211, n25212, n25213,
    n25214, n25215, n25216, n25217, n25218, n25219,
    n25220, n25221, n25222, n25223, n25224, n25225,
    n25226, n25227, n25228, n25229, n25230, n25231,
    n25232, n25233, n25234, n25235, n25236, n25237,
    n25238, n25239, n25240, n25241, n25242, n25243,
    n25244, n25245, n25246, n25247, n25248, n25249,
    n25250, n25251, n25252, n25253, n25254, n25255,
    n25256, n25257, n25258, n25259, n25260, n25261,
    n25262, n25263, n25264, n25265, n25266, n25267,
    n25268, n25269, n25270, n25271, n25272, n25273,
    n25274, n25275, n25276, n25277, n25278, n25279,
    n25280, n25281, n25282, n25283, n25284, n25285,
    n25286, n25287, n25288, n25289, n25290, n25291,
    n25292, n25293, n25294, n25295, n25296, n25297,
    n25298, n25299, n25300, n25301, n25302, n25303,
    n25304, n25305, n25306, n25307, n25308, n25309,
    n25310, n25311, n25312, n25313, n25314, n25315,
    n25316, n25317, n25318, n25319, n25320, n25321,
    n25322, n25323, n25324, n25325, n25326, n25327,
    n25328, n25329, n25330, n25331, n25332, n25333,
    n25334, n25335, n25336, n25337, n25338, n25339,
    n25340, n25341, n25342, n25343, n25344, n25345,
    n25346, n25347, n25348, n25349, n25350, n25351,
    n25352, n25353, n25354, n25355, n25356, n25357,
    n25358, n25359, n25360, n25361, n25362, n25363,
    n25364, n25365, n25366, n25367, n25368, n25369,
    n25370, n25371, n25372, n25373, n25374, n25375,
    n25376, n25377, n25378, n25379, n25380, n25381,
    n25382, n25383, n25384, n25385, n25386, n25387,
    n25388, n25389, n25390, n25391, n25392, n25393,
    n25394, n25395, n25396, n25397, n25398, n25399,
    n25400, n25401, n25402, n25403, n25404, n25405,
    n25406, n25407, n25408, n25409, n25410, n25411,
    n25412, n25413, n25414, n25415, n25416, n25417,
    n25418, n25419, n25420, n25421, n25422, n25423,
    n25424, n25425, n25426, n25427, n25428, n25429,
    n25430, n25431, n25432, n25433, n25434, n25435,
    n25436, n25437, n25438, n25439, n25440, n25441,
    n25442, n25443, n25444, n25445, n25446, n25447,
    n25448, n25449, n25450, n25451, n25452, n25453,
    n25454, n25455, n25456, n25457, n25458, n25459,
    n25460, n25461, n25462, n25463, n25464, n25465,
    n25466, n25467, n25468, n25469, n25470, n25471,
    n25472, n25473, n25474, n25475, n25476, n25477,
    n25478, n25479, n25480, n25481, n25482, n25483,
    n25484, n25485, n25486, n25487, n25488, n25489,
    n25490, n25491, n25492, n25493, n25494, n25495,
    n25496, n25497, n25498, n25499, n25500, n25501,
    n25502, n25503, n25504, n25505, n25506, n25507,
    n25508, n25509, n25510, n25511, n25512, n25513,
    n25514, n25515, n25516, n25517, n25518, n25519,
    n25520, n25521, n25522, n25523, n25524, n25525,
    n25526, n25527, n25528, n25529, n25530, n25531,
    n25532, n25533, n25534, n25535, n25536, n25537,
    n25538, n25539, n25540, n25541, n25542, n25543,
    n25544, n25545, n25546, n25547, n25548, n25549,
    n25550, n25551, n25552, n25553, n25554, n25555,
    n25556, n25557, n25558, n25559, n25560, n25561,
    n25562, n25563, n25564, n25565, n25566, n25567,
    n25568, n25569, n25570, n25571, n25572, n25573,
    n25574, n25575, n25576, n25577, n25578, n25579,
    n25580, n25581, n25582, n25583, n25584, n25585,
    n25586, n25587, n25588, n25589, n25590, n25591,
    n25592, n25593, n25594, n25595, n25596, n25597,
    n25598, n25599, n25600, n25601, n25602, n25603,
    n25604, n25605, n25606, n25607, n25608, n25609,
    n25610, n25611, n25612, n25613, n25614, n25615,
    n25616, n25617, n25618, n25619, n25620, n25621,
    n25622, n25623, n25624, n25625, n25626, n25627,
    n25628, n25629, n25630, n25631, n25632, n25633,
    n25634, n25635, n25636, n25637, n25638, n25639,
    n25640, n25641, n25642, n25643, n25644, n25645,
    n25646, n25647, n25648, n25649, n25650, n25651,
    n25652, n25653, n25654, n25655, n25656, n25657,
    n25658, n25659, n25660, n25661, n25662, n25663,
    n25664, n25665, n25666, n25667, n25668, n25669,
    n25670, n25671, n25672, n25673, n25674, n25675,
    n25676, n25677, n25678, n25679, n25680, n25681,
    n25682, n25683, n25684, n25685, n25686, n25687,
    n25688, n25689, n25690, n25691, n25692, n25693,
    n25694, n25695, n25696, n25697, n25698, n25699,
    n25700, n25701, n25702, n25703, n25704, n25705,
    n25706, n25707, n25708, n25709, n25710, n25711,
    n25712, n25713, n25714, n25715, n25716, n25717,
    n25718, n25719, n25720, n25721, n25722, n25723,
    n25724, n25725, n25726, n25727, n25728, n25729,
    n25730, n25731, n25732, n25733, n25734, n25735,
    n25736, n25737, n25738, n25739, n25740, n25741,
    n25742, n25743, n25744, n25745, n25746, n25747,
    n25748, n25749, n25750, n25751, n25752, n25753,
    n25754, n25755, n25756, n25757, n25758, n25759,
    n25760, n25761, n25762, n25763, n25764, n25765,
    n25766, n25767, n25768, n25769, n25770, n25771,
    n25772, n25773, n25774, n25775, n25776, n25777,
    n25778, n25779, n25780, n25781, n25782, n25783,
    n25784, n25785, n25786, n25787, n25788, n25789,
    n25790, n25791, n25792, n25793, n25794, n25795,
    n25796, n25797, n25798, n25799, n25800, n25801,
    n25802, n25803, n25804, n25805, n25806, n25807,
    n25808, n25809, n25810, n25811, n25812, n25813,
    n25814, n25815, n25816, n25817, n25818, n25819,
    n25820, n25821, n25822, n25823, n25824, n25825,
    n25826, n25827, n25828, n25829, n25830, n25831,
    n25832, n25833, n25834, n25835, n25836, n25837,
    n25838, n25839, n25840, n25841, n25842, n25843,
    n25844, n25845, n25846, n25847, n25848, n25849,
    n25850, n25851, n25852, n25853, n25854, n25855,
    n25856, n25857, n25858, n25859, n25860, n25861,
    n25862, n25863, n25864, n25865, n25866, n25867,
    n25868, n25869, n25870, n25871, n25872, n25873,
    n25874, n25875, n25876, n25877, n25878, n25879,
    n25880, n25881, n25882, n25883, n25884, n25885,
    n25886, n25887, n25888, n25889, n25890, n25891,
    n25892, n25893, n25894, n25895, n25896, n25897,
    n25898, n25899, n25900, n25901, n25902, n25903,
    n25904, n25905, n25906, n25907, n25908, n25909,
    n25910, n25911, n25912, n25913, n25914, n25915,
    n25916, n25917, n25918, n25919, n25920, n25921,
    n25922, n25923, n25924, n25925, n25926, n25927,
    n25928, n25929, n25930, n25931, n25932, n25933,
    n25934, n25935, n25936, n25937, n25938, n25939,
    n25940, n25941, n25942, n25943, n25944, n25945,
    n25946, n25947, n25948, n25949, n25950, n25951,
    n25952, n25953, n25954, n25955, n25956, n25957,
    n25958, n25959, n25960, n25961, n25962, n25963,
    n25964, n25965, n25966, n25967, n25968, n25969,
    n25970, n25971, n25972, n25973, n25974, n25975,
    n25976, n25977, n25978, n25979, n25980, n25981,
    n25982, n25983, n25984, n25985, n25986, n25987,
    n25988, n25989, n25990, n25991, n25992, n25993,
    n25994, n25995, n25996, n25997, n25998, n25999,
    n26000, n26001, n26002, n26003, n26004, n26005,
    n26006, n26007, n26008, n26009, n26010, n26011,
    n26012, n26013, n26014, n26015, n26016, n26017,
    n26018, n26019, n26020, n26021, n26022, n26023,
    n26024, n26025, n26026, n26027, n26028, n26029,
    n26030, n26031, n26032, n26033, n26034, n26035,
    n26036, n26037, n26038, n26039, n26040, n26041,
    n26042, n26043, n26044, n26045, n26046, n26047,
    n26048, n26049, n26050, n26051, n26052, n26053,
    n26054, n26055, n26056, n26057, n26058, n26059,
    n26060, n26061, n26062, n26063, n26064, n26065,
    n26066, n26067, n26068, n26069, n26070, n26071,
    n26072, n26073, n26074, n26075, n26076, n26077,
    n26078, n26079, n26080, n26081, n26082, n26083,
    n26084, n26085, n26086, n26087, n26088, n26089,
    n26090, n26091, n26092, n26093, n26094, n26095,
    n26096, n26097, n26098, n26099, n26100, n26101,
    n26102, n26103, n26104, n26105, n26106, n26107,
    n26108, n26109, n26110, n26111, n26112, n26113,
    n26114, n26115, n26116, n26117, n26118, n26119,
    n26120, n26121, n26122, n26123, n26124, n26125,
    n26126, n26127, n26128, n26129, n26130, n26131,
    n26132, n26133, n26134, n26135, n26136, n26137,
    n26138, n26139, n26140, n26141, n26142, n26143,
    n26144, n26145, n26146, n26147, n26148, n26149,
    n26150, n26151, n26152, n26153, n26154, n26155,
    n26156, n26157, n26158, n26159, n26160, n26161,
    n26162, n26163, n26164, n26165, n26166, n26167,
    n26168, n26169, n26170, n26171, n26172, n26173,
    n26174, n26175, n26176, n26177, n26178, n26179,
    n26180, n26181, n26182, n26183, n26184, n26185,
    n26186, n26187, n26188, n26189, n26190, n26191,
    n26192, n26193, n26194, n26195, n26196, n26197,
    n26198, n26199, n26200, n26201, n26202, n26203,
    n26204, n26205, n26206, n26207, n26208, n26209,
    n26210, n26211, n26212, n26213, n26214, n26215,
    n26216, n26217, n26218, n26219, n26220, n26221,
    n26222, n26223, n26224, n26225, n26226, n26227,
    n26228, n26229, n26230, n26231, n26232, n26233,
    n26234, n26235, n26236, n26237, n26238, n26239,
    n26240, n26241, n26242, n26243, n26244, n26245,
    n26246, n26247, n26248, n26249, n26250, n26251,
    n26252, n26253, n26254, n26255, n26256, n26257,
    n26258, n26259, n26260, n26261, n26262, n26263,
    n26264, n26265, n26266, n26267, n26268, n26269,
    n26270, n26271, n26272, n26273, n26274, n26275,
    n26276, n26277, n26278, n26279, n26280, n26281,
    n26282, n26283, n26284, n26285, n26286, n26287,
    n26288, n26289, n26290, n26291, n26292, n26293,
    n26294, n26295, n26296, n26297, n26298, n26299,
    n26300, n26301, n26302, n26303, n26304, n26305,
    n26306, n26307, n26308, n26309, n26310, n26311,
    n26312, n26313, n26314, n26315, n26316, n26317,
    n26318, n26319, n26320, n26321, n26322, n26323,
    n26324, n26325, n26326, n26327, n26328, n26329,
    n26330, n26331, n26332, n26333, n26334, n26335,
    n26336, n26337, n26338, n26339, n26340, n26341,
    n26342, n26343, n26344, n26345, n26346, n26347,
    n26348, n26349, n26350, n26351, n26352, n26353,
    n26354, n26355, n26356, n26357, n26358, n26359,
    n26360, n26361, n26362, n26363, n26364, n26365,
    n26366, n26367, n26368, n26369, n26370, n26371,
    n26372, n26373, n26374, n26375, n26376, n26377,
    n26378, n26379, n26380, n26381, n26382, n26383,
    n26384, n26385, n26386, n26387, n26388, n26389,
    n26390, n26391, n26392, n26393, n26394, n26395,
    n26396, n26397, n26398, n26399, n26400, n26401,
    n26402, n26403, n26404, n26405, n26406, n26407,
    n26408, n26409, n26410, n26411, n26412, n26413,
    n26414, n26415, n26416, n26417, n26418, n26419,
    n26420, n26421, n26422, n26423, n26424, n26425,
    n26426, n26427, n26428, n26429, n26430, n26431,
    n26432, n26433, n26434, n26435, n26436, n26437,
    n26438, n26439, n26440, n26441, n26442, n26443,
    n26444, n26445, n26446, n26447, n26448, n26449,
    n26450, n26451, n26452, n26453, n26454, n26455,
    n26456, n26457, n26458, n26459, n26460, n26461,
    n26462, n26463, n26464, n26465, n26466, n26467,
    n26468, n26469, n26470, n26471, n26472, n26473,
    n26474, n26475, n26476, n26477, n26478, n26479,
    n26480, n26481, n26482, n26483, n26484, n26485,
    n26486, n26487, n26488, n26489, n26490, n26491,
    n26492, n26493, n26494, n26495, n26496, n26497,
    n26498, n26499, n26500, n26501, n26502, n26503,
    n26504, n26505, n26506, n26507, n26508, n26509,
    n26510, n26511, n26512, n26513, n26514, n26515,
    n26516, n26517, n26518, n26519, n26520, n26521,
    n26522, n26523, n26524, n26525, n26526, n26527,
    n26528, n26529, n26530, n26531, n26532, n26533,
    n26534, n26535, n26536, n26537, n26538, n26539,
    n26540, n26541, n26542, n26543, n26544, n26545,
    n26546, n26547, n26548, n26549, n26550, n26551,
    n26552, n26553, n26554, n26555, n26556, n26557,
    n26558, n26559, n26560, n26561, n26562, n26563,
    n26564, n26565, n26566, n26567, n26568, n26569,
    n26570, n26571, n26572, n26573, n26574, n26575,
    n26576, n26577, n26578, n26579, n26580, n26581,
    n26582, n26583, n26584, n26585, n26586, n26587,
    n26588, n26589, n26590, n26591, n26592, n26593,
    n26594, n26595, n26596, n26597, n26598, n26599,
    n26600, n26601, n26602, n26603, n26604, n26605,
    n26606, n26607, n26608, n26609, n26610, n26611,
    n26612, n26613, n26614, n26615, n26616, n26617,
    n26618, n26619, n26620, n26621, n26622, n26623,
    n26624, n26625, n26626, n26627, n26628, n26629,
    n26630, n26631, n26632, n26633, n26634, n26635,
    n26636, n26637, n26638, n26639, n26640, n26641,
    n26642, n26643, n26644, n26645, n26646, n26647,
    n26648, n26649, n26650, n26651, n26652, n26653,
    n26654, n26655, n26656, n26657, n26658, n26659,
    n26660, n26661, n26662, n26663, n26664, n26665,
    n26666, n26667, n26668, n26669, n26670, n26671,
    n26672, n26673, n26674, n26675, n26676, n26677,
    n26678, n26679, n26680, n26681, n26682, n26683,
    n26684, n26685, n26686, n26687, n26688, n26689,
    n26690, n26691, n26692, n26693, n26694, n26695,
    n26696, n26697, n26698, n26699, n26700, n26701,
    n26702, n26703, n26704, n26705, n26706, n26707,
    n26708, n26709, n26710, n26711, n26712, n26713,
    n26714, n26715, n26716, n26717, n26718, n26719,
    n26720, n26721, n26722, n26723, n26724, n26725,
    n26726, n26727, n26728, n26729, n26730, n26731,
    n26732, n26733, n26734, n26735, n26736, n26737,
    n26738, n26739, n26740, n26741, n26742, n26743,
    n26744, n26745, n26746, n26747, n26748, n26749,
    n26750, n26751, n26752, n26753, n26754, n26755,
    n26756, n26757, n26758, n26759, n26760, n26761,
    n26762, n26763, n26764, n26765, n26766, n26767,
    n26768, n26769, n26770, n26771, n26772, n26773,
    n26774, n26775, n26776, n26777, n26778, n26779,
    n26780, n26781, n26782, n26783, n26784, n26785,
    n26786, n26787, n26788, n26789, n26790, n26791,
    n26792, n26793, n26794, n26795, n26796, n26797,
    n26798, n26799, n26800, n26801, n26802, n26803,
    n26804, n26805, n26806, n26807, n26808, n26809,
    n26810, n26811, n26812, n26813, n26814, n26815,
    n26816, n26817, n26818, n26819, n26820, n26821,
    n26822, n26823, n26824, n26825, n26826, n26827,
    n26828, n26829, n26830, n26831, n26832, n26833,
    n26834, n26835, n26836, n26837, n26838, n26839,
    n26840, n26841, n26842, n26843, n26844, n26845,
    n26846, n26847, n26848, n26849, n26850, n26851,
    n26852, n26853, n26854, n26855, n26856, n26857,
    n26858, n26859, n26860, n26861, n26862, n26863,
    n26864, n26865, n26866, n26867, n26868, n26869,
    n26870, n26871, n26872, n26873, n26874, n26875,
    n26876, n26877, n26878, n26879, n26880, n26881,
    n26882, n26883, n26884, n26885, n26886, n26887,
    n26888, n26889, n26890, n26891, n26892, n26893,
    n26894, n26895, n26896, n26897, n26898, n26899,
    n26900, n26901, n26902, n26903, n26904, n26905,
    n26906, n26907, n26908, n26909, n26910, n26911,
    n26912, n26913, n26914, n26915, n26916, n26917,
    n26918, n26919, n26920, n26921, n26922, n26923,
    n26924, n26925, n26926, n26927, n26928, n26929,
    n26930, n26931, n26932, n26933, n26934, n26935,
    n26936, n26937, n26938, n26939, n26940, n26941,
    n26942, n26943, n26944, n26945, n26946, n26947,
    n26948, n26949, n26950, n26951, n26952, n26953,
    n26954, n26955, n26956, n26957, n26958, n26959,
    n26960, n26961, n26962, n26963, n26964, n26965,
    n26966, n26967, n26968, n26969, n26970, n26971,
    n26972, n26973, n26974, n26975, n26976, n26977,
    n26978, n26979, n26980, n26981, n26982, n26983,
    n26984, n26985, n26986, n26987, n26988, n26989,
    n26990, n26991, n26992, n26993, n26994, n26995,
    n26996, n26997, n26998, n26999, n27000, n27001,
    n27002, n27003, n27004, n27005, n27006, n27007,
    n27008, n27009, n27010, n27011, n27012, n27013,
    n27014, n27015, n27016, n27017, n27018, n27019,
    n27020, n27021, n27022, n27023, n27024, n27025,
    n27026, n27027, n27028, n27029, n27030, n27031,
    n27032, n27033, n27034, n27035, n27036, n27037,
    n27038, n27039, n27040, n27041, n27042, n27043,
    n27044, n27045, n27046, n27047, n27048, n27049,
    n27050, n27051, n27052, n27053, n27054, n27055,
    n27056, n27057, n27058, n27059, n27060, n27061,
    n27062, n27063, n27064, n27065, n27066, n27067,
    n27068, n27069, n27070, n27071, n27072, n27073,
    n27074, n27075, n27076, n27077, n27078, n27079,
    n27080, n27081, n27082, n27083, n27084, n27085,
    n27086, n27087, n27088, n27089, n27090, n27091,
    n27092, n27093, n27094, n27095, n27096, n27097,
    n27098, n27099, n27100, n27101, n27102, n27103,
    n27104, n27105, n27106, n27107, n27108, n27109,
    n27110, n27111, n27112, n27113, n27114, n27115,
    n27116, n27117, n27118, n27119, n27120, n27121,
    n27122, n27123, n27124, n27125, n27126, n27127,
    n27128, n27129, n27130, n27131, n27132, n27133,
    n27134, n27135, n27136, n27137, n27138, n27139,
    n27140, n27141, n27142, n27143, n27144, n27145,
    n27146, n27147, n27148, n27149, n27150, n27151,
    n27152, n27153, n27154, n27155, n27156, n27157,
    n27158, n27159, n27160, n27161, n27162, n27163,
    n27164, n27165, n27166, n27167, n27168, n27169,
    n27170, n27171, n27172, n27173, n27174, n27175,
    n27176, n27177, n27178, n27179, n27180, n27181,
    n27182, n27183, n27184, n27185, n27186, n27187,
    n27188, n27189, n27190, n27191, n27192, n27193,
    n27194, n27195, n27196, n27197, n27198, n27199,
    n27200, n27201, n27202, n27203, n27204, n27205,
    n27206, n27207, n27208, n27209, n27210, n27211,
    n27212, n27213, n27214, n27215, n27216, n27217,
    n27218, n27219, n27220, n27221, n27222, n27223,
    n27224, n27225, n27226, n27227, n27228, n27229,
    n27230, n27231, n27232, n27233, n27234, n27235,
    n27236, n27237, n27238, n27239, n27240, n27241,
    n27242, n27243, n27244, n27245, n27246, n27247,
    n27248, n27249, n27250, n27251, n27252, n27253,
    n27254, n27255, n27256, n27257, n27258, n27259,
    n27260, n27261, n27262, n27263, n27264, n27265,
    n27266, n27267, n27268, n27269, n27270, n27271,
    n27272, n27273, n27274, n27275, n27276, n27277,
    n27278, n27279, n27280, n27281, n27282, n27283,
    n27284, n27285, n27286, n27287, n27288, n27289,
    n27290, n27291, n27292, n27293, n27294, n27295,
    n27296, n27297, n27298, n27299, n27300, n27301,
    n27302, n27303, n27304, n27305, n27306, n27307,
    n27308, n27309, n27310, n27311, n27312, n27313,
    n27314, n27315, n27316, n27317, n27318, n27319,
    n27320, n27321, n27322, n27323, n27324, n27325,
    n27326, n27327, n27328, n27329, n27330, n27331,
    n27332, n27333, n27334, n27335, n27336, n27337,
    n27338, n27339, n27340, n27341, n27342, n27343,
    n27344, n27345, n27346, n27347, n27348, n27349,
    n27350, n27351, n27352, n27353, n27354, n27355,
    n27356, n27357, n27358, n27359, n27360, n27361,
    n27362, n27363, n27364, n27365, n27366, n27367,
    n27368, n27369, n27370, n27371, n27372, n27373,
    n27374, n27375, n27376, n27377, n27378, n27379,
    n27380, n27381, n27382, n27383, n27384, n27385,
    n27386, n27387, n27388, n27389, n27390, n27391,
    n27392, n27393, n27394, n27395, n27396, n27397,
    n27398, n27399, n27400, n27401, n27402, n27403,
    n27404, n27405, n27406, n27407, n27408, n27409,
    n27410, n27411, n27412, n27413, n27414, n27415,
    n27416, n27417, n27418, n27419, n27420, n27421,
    n27422, n27423, n27424, n27425, n27426, n27427,
    n27428, n27429, n27430, n27431, n27432, n27433,
    n27434, n27435, n27436, n27437, n27438, n27439,
    n27440, n27441, n27442, n27443, n27444, n27445,
    n27446, n27447, n27448, n27449, n27450, n27451,
    n27452, n27453, n27454, n27455, n27456, n27457,
    n27458, n27459, n27460, n27461, n27462, n27463,
    n27464, n27465, n27466, n27467, n27468, n27469,
    n27470, n27471, n27472, n27473, n27474, n27475,
    n27476, n27477, n27478, n27479, n27480, n27481,
    n27482, n27483, n27484, n27485, n27486, n27487,
    n27488, n27489, n27490, n27491, n27492, n27493,
    n27494, n27495, n27496, n27497, n27498, n27499,
    n27500, n27501, n27502, n27503, n27504, n27505,
    n27506, n27507, n27508, n27509, n27510, n27511,
    n27512, n27513, n27514, n27515, n27516, n27517,
    n27518, n27519, n27520, n27521, n27522, n27523,
    n27524, n27525, n27526, n27527, n27528, n27529,
    n27530, n27531, n27532, n27533, n27534, n27535,
    n27536, n27537, n27538, n27539, n27540, n27541,
    n27542, n27543, n27544, n27545, n27546, n27547,
    n27548, n27549, n27550, n27551, n27552, n27553,
    n27554, n27555, n27556, n27557, n27558, n27559,
    n27560, n27561, n27562, n27563, n27564, n27565,
    n27566, n27567, n27568, n27569, n27570, n27571,
    n27572, n27573, n27574, n27575, n27576, n27577,
    n27578, n27579, n27580, n27581, n27582, n27583,
    n27584, n27585, n27586, n27587, n27588, n27589,
    n27590, n27591, n27592, n27593, n27594, n27595,
    n27596, n27597, n27598, n27599, n27600, n27601,
    n27602, n27603, n27604, n27605, n27606, n27607,
    n27608, n27609, n27610, n27611, n27612, n27613,
    n27614, n27615, n27616, n27617, n27618, n27619,
    n27620, n27621, n27622, n27623, n27624, n27625,
    n27626, n27627, n27628, n27629, n27630, n27631,
    n27632, n27633, n27634, n27635, n27636, n27637,
    n27638, n27639, n27640, n27641, n27642, n27643,
    n27644, n27645, n27646, n27647, n27648, n27649,
    n27650, n27651, n27652, n27653, n27654, n27655,
    n27656, n27657, n27658, n27659, n27660, n27661,
    n27662, n27663, n27664, n27665, n27666, n27667,
    n27668, n27669, n27670, n27671, n27672, n27673,
    n27674, n27675, n27676, n27677, n27678, n27679,
    n27680, n27681, n27682, n27683, n27684, n27685,
    n27686, n27687, n27688, n27689, n27690, n27691,
    n27692, n27693, n27694, n27695, n27696, n27697,
    n27698, n27699, n27700, n27701, n27702, n27703,
    n27704, n27705, n27706, n27707, n27708, n27709,
    n27710, n27711, n27712, n27713, n27714, n27715,
    n27716, n27717, n27718, n27719, n27720, n27721,
    n27722, n27723, n27724, n27725, n27726, n27727,
    n27728, n27729, n27730, n27731, n27732, n27733,
    n27734, n27735, n27736, n27737, n27738, n27739,
    n27740, n27741, n27742, n27743, n27744, n27745,
    n27746, n27747, n27748, n27749, n27750, n27751,
    n27752, n27753, n27754, n27755, n27756, n27757,
    n27758, n27759, n27760, n27761, n27762, n27763,
    n27764, n27765, n27766, n27767, n27768, n27769,
    n27770, n27771, n27772, n27773, n27774, n27775,
    n27776, n27777, n27778, n27779, n27780, n27781,
    n27782, n27783, n27784, n27785, n27786, n27787,
    n27788, n27789, n27790, n27791, n27792, n27793,
    n27794, n27795, n27796, n27797, n27798, n27799,
    n27800, n27801, n27802, n27803, n27804, n27805,
    n27806, n27807, n27808, n27809, n27810, n27811,
    n27812, n27813, n27814, n27815, n27816, n27817,
    n27818, n27819, n27820, n27821, n27822, n27823,
    n27824, n27825, n27826, n27827, n27828, n27829,
    n27830, n27831, n27832, n27833, n27834, n27835,
    n27836, n27837, n27838, n27839, n27840, n27841,
    n27842, n27843, n27844, n27845, n27846, n27847,
    n27848, n27849, n27850, n27851, n27852, n27853,
    n27854, n27855, n27856, n27857, n27858, n27859,
    n27860, n27861, n27862, n27863, n27864, n27865,
    n27866, n27867, n27868, n27869, n27870, n27871,
    n27872, n27873, n27874, n27875, n27876, n27877,
    n27878, n27879, n27880, n27881, n27882, n27883,
    n27884, n27885, n27886, n27887, n27888, n27889,
    n27890, n27891, n27892, n27893, n27894, n27895,
    n27896, n27897, n27898, n27899, n27900, n27901,
    n27902, n27903, n27904, n27905, n27906, n27907,
    n27908, n27909, n27910, n27911, n27912, n27913,
    n27914, n27915, n27916, n27917, n27918, n27919,
    n27920, n27921, n27922, n27923, n27924, n27925,
    n27926, n27927, n27928, n27929, n27930, n27931,
    n27932, n27933, n27934, n27935, n27936, n27937,
    n27938, n27939, n27940, n27941, n27942, n27943,
    n27944, n27945, n27946, n27947, n27948, n27949,
    n27950, n27951, n27952, n27953, n27954, n27955,
    n27956, n27957, n27958, n27959, n27960, n27961,
    n27962, n27963, n27964, n27965, n27966, n27967,
    n27968, n27969, n27970, n27971, n27972, n27973,
    n27974, n27975, n27976, n27977, n27978, n27979,
    n27980, n27981, n27982, n27983, n27984, n27985,
    n27986, n27987, n27988, n27989, n27990, n27991,
    n27992, n27993, n27994, n27995, n27996, n27997,
    n27998, n27999, n28000, n28001, n28002, n28003,
    n28004, n28005, n28006, n28007, n28008, n28009,
    n28010, n28011, n28012, n28013, n28014, n28015,
    n28016, n28017, n28018, n28019, n28020, n28021,
    n28022, n28023, n28024, n28025, n28026, n28027,
    n28028, n28029, n28030, n28031, n28032, n28033,
    n28034, n28035, n28036, n28037, n28038, n28039,
    n28040, n28041, n28042, n28043, n28044, n28045,
    n28046, n28047, n28048, n28049, n28050, n28051,
    n28052, n28053, n28054, n28055, n28056, n28057,
    n28058, n28059, n28060, n28061, n28062, n28063,
    n28064, n28065, n28066, n28067, n28068, n28069,
    n28070, n28071, n28072, n28073, n28074, n28075,
    n28076, n28077, n28078, n28079, n28080, n28081,
    n28082, n28083, n28084, n28085, n28086, n28087,
    n28088, n28089, n28090, n28091, n28092, n28093,
    n28094, n28095, n28096, n28097, n28098, n28099,
    n28100, n28101, n28102, n28103, n28104, n28105,
    n28106, n28107, n28108, n28109, n28110, n28111,
    n28112, n28113, n28114, n28115, n28116, n28117,
    n28118, n28119, n28120, n28121, n28122, n28123,
    n28124, n28125, n28126, n28127, n28128, n28129,
    n28130, n28131, n28132, n28133, n28134, n28135,
    n28136, n28137, n28138, n28139, n28140, n28141,
    n28142, n28143, n28144, n28145, n28146, n28147,
    n28148, n28149, n28150, n28151, n28152, n28153,
    n28154, n28155, n28156, n28157, n28158, n28159,
    n28160, n28161, n28162, n28163, n28164, n28165,
    n28166, n28167, n28168, n28169, n28170, n28171,
    n28172, n28173, n28174, n28175, n28176, n28177,
    n28178, n28179, n28180, n28181, n28182, n28183,
    n28184, n28185, n28186, n28187, n28188, n28189,
    n28190, n28191, n28192, n28193, n28194, n28195,
    n28196, n28197, n28198, n28199, n28200, n28201,
    n28202, n28203, n28204, n28205, n28206, n28207,
    n28208, n28209, n28210, n28211, n28212, n28213,
    n28214, n28215, n28216, n28217, n28218, n28219,
    n28220, n28221, n28222, n28223, n28224, n28225,
    n28226, n28227, n28228, n28229, n28230, n28231,
    n28232, n28233, n28234, n28235, n28236, n28237,
    n28238, n28239, n28240, n28241, n28242, n28243,
    n28244, n28245, n28246, n28247, n28248, n28249,
    n28250, n28251, n28252, n28253, n28254, n28255,
    n28256, n28257, n28258, n28259, n28260, n28261,
    n28262, n28263, n28264, n28265, n28266, n28267,
    n28268, n28269, n28270, n28271, n28272, n28273,
    n28274, n28275, n28276, n28277, n28278, n28279,
    n28280, n28281, n28282, n28283, n28284, n28285,
    n28286, n28287, n28288, n28289, n28290, n28291,
    n28292, n28293, n28294, n28295, n28296, n28297,
    n28298, n28299, n28300, n28301, n28302, n28303,
    n28304, n28305, n28306, n28307, n28308, n28309,
    n28310, n28311, n28312, n28313, n28314, n28315,
    n28316, n28317, n28318, n28319, n28320, n28321,
    n28322, n28323, n28324, n28325, n28326, n28327,
    n28328, n28329, n28330, n28331, n28332, n28333,
    n28334, n28335, n28336, n28337, n28338, n28339,
    n28340, n28341, n28342, n28343, n28344, n28345,
    n28346, n28347, n28348, n28349, n28350, n28351,
    n28352, n28353, n28354, n28355, n28356, n28357,
    n28358, n28359, n28360, n28361, n28362, n28363,
    n28364, n28365, n28366, n28367, n28368, n28369,
    n28370, n28371, n28372, n28373, n28374, n28375,
    n28376, n28377, n28378, n28379, n28380, n28381,
    n28382, n28383, n28384, n28385, n28386, n28387,
    n28388, n28389, n28390, n28391, n28392, n28393,
    n28394, n28395, n28396, n28397, n28398, n28399,
    n28400, n28401, n28402, n28403, n28404, n28405,
    n28406, n28407, n28408, n28409, n28410, n28411,
    n28412, n28413, n28414, n28415, n28416, n28417,
    n28418, n28419, n28420, n28421, n28422, n28423,
    n28424, n28425, n28426, n28427, n28428, n28429,
    n28430, n28431, n28432, n28433, n28434, n28435,
    n28436, n28437, n28438, n28439, n28440, n28441,
    n28442, n28443, n28444, n28445, n28446, n28447,
    n28448, n28449, n28450, n28451, n28452, n28453,
    n28454, n28455, n28456, n28457, n28458, n28459,
    n28460, n28461, n28462, n28463, n28464, n28465,
    n28466, n28467, n28468, n28469, n28470, n28471,
    n28472, n28473, n28474, n28475, n28476, n28477,
    n28478, n28479, n28480, n28481, n28482, n28483,
    n28484, n28485, n28486, n28487, n28488, n28489,
    n28490, n28491, n28492, n28493, n28494, n28495,
    n28496, n28497, n28498, n28499, n28500, n28501,
    n28502, n28503, n28504, n28505, n28506, n28507,
    n28508, n28509, n28510, n28511, n28512, n28513,
    n28514, n28515, n28516, n28517, n28518, n28519,
    n28520, n28521, n28522, n28523, n28524, n28525,
    n28526, n28527, n28528, n28529, n28530, n28531,
    n28532, n28533, n28534, n28535, n28536, n28537,
    n28538, n28539, n28540, n28541, n28542, n28543,
    n28544, n28545, n28546, n28547, n28548, n28549,
    n28550, n28551, n28552, n28553, n28554, n28555,
    n28556, n28557, n28558, n28559, n28560, n28561,
    n28562, n28563, n28564, n28565, n28566, n28567,
    n28568, n28569, n28570, n28571, n28572, n28573,
    n28574, n28575, n28576, n28577, n28578, n28579,
    n28580, n28581, n28582, n28583, n28584, n28585,
    n28586, n28587, n28588, n28589, n28590, n28591,
    n28592, n28593, n28594, n28595, n28596, n28597,
    n28598, n28599, n28600, n28601, n28602, n28603,
    n28604, n28605, n28606, n28607, n28608, n28609,
    n28610, n28611, n28612, n28613, n28614, n28615,
    n28616, n28617, n28618, n28619, n28620, n28621,
    n28622, n28623, n28624, n28625, n28626, n28627,
    n28628, n28629, n28630, n28631, n28632, n28633,
    n28634, n28635, n28636, n28637, n28638, n28639,
    n28640, n28641, n28642, n28643, n28644, n28645,
    n28646, n28647, n28648, n28649, n28650, n28651,
    n28652, n28653, n28654, n28655, n28656, n28657,
    n28658, n28659, n28660, n28661, n28662, n28663,
    n28664, n28665, n28666, n28667, n28668, n28669,
    n28670, n28671, n28672, n28673, n28674, n28675,
    n28676, n28677, n28678, n28679, n28680, n28681,
    n28682, n28683, n28684, n28685, n28686, n28687,
    n28688, n28689, n28690, n28691, n28692, n28693,
    n28694, n28695, n28696, n28697, n28698, n28699,
    n28700, n28701, n28702, n28703, n28704, n28705,
    n28706, n28707, n28708, n28709, n28710, n28711,
    n28712, n28713, n28714, n28715, n28716, n28717,
    n28718, n28719, n28720, n28721, n28722, n28723,
    n28724, n28725, n28726, n28727, n28728, n28729,
    n28730, n28731, n28732, n28733, n28734, n28735,
    n28736, n28737, n28738, n28739, n28740, n28741,
    n28742, n28743, n28744, n28745, n28746, n28747,
    n28748, n28749, n28750, n28751, n28752, n28753,
    n28754, n28755, n28756, n28757, n28758, n28759,
    n28760, n28761, n28762, n28763, n28764, n28765,
    n28766, n28767, n28768, n28769, n28770, n28771,
    n28772, n28773, n28774, n28775, n28776, n28777,
    n28778, n28779, n28780, n28781, n28782, n28783,
    n28784, n28785, n28786, n28787, n28788, n28789,
    n28790, n28791, n28792, n28793, n28794, n28795,
    n28796, n28797, n28798, n28799, n28800, n28801,
    n28802, n28803, n28804, n28805, n28806, n28807,
    n28808, n28809, n28810, n28811, n28812, n28813,
    n28814, n28815, n28816, n28817, n28818, n28819,
    n28820, n28821, n28822, n28823, n28824, n28825,
    n28826, n28827, n28828, n28829, n28830, n28831,
    n28832, n28833, n28834, n28835, n28836, n28837,
    n28838, n28839, n28840, n28841, n28842, n28843,
    n28844, n28845, n28846, n28847, n28848, n28849,
    n28850, n28851, n28852, n28853, n28854, n28855,
    n28856, n28857, n28858, n28859, n28860, n28861,
    n28862, n28863, n28864, n28865, n28866, n28867,
    n28868, n28869, n28870, n28871, n28872, n28873,
    n28874, n28875, n28876, n28877, n28878, n28879,
    n28880, n28881, n28882, n28883, n28884, n28885,
    n28886, n28887, n28888, n28889, n28890, n28891,
    n28892, n28893, n28894, n28895, n28896, n28897,
    n28898, n28899, n28900, n28901, n28902, n28903,
    n28904, n28905, n28906, n28907, n28908, n28909,
    n28910, n28911, n28912, n28913, n28914, n28915,
    n28916, n28917, n28918, n28919, n28920, n28921,
    n28922, n28923, n28924, n28925, n28926, n28927,
    n28928, n28929, n28930, n28931, n28932, n28933,
    n28934, n28935, n28936, n28937, n28938, n28939,
    n28940, n28941, n28942, n28943, n28944, n28945,
    n28946, n28947, n28948, n28949, n28950, n28951,
    n28952, n28953, n28954, n28955, n28956, n28957,
    n28958, n28959, n28960, n28961, n28962, n28963,
    n28964, n28965, n28966, n28967, n28968, n28969,
    n28970, n28971, n28972, n28973, n28974, n28975,
    n28976, n28977, n28978, n28979, n28980, n28981,
    n28982, n28983, n28984, n28985, n28986, n28987,
    n28988, n28989, n28990, n28991, n28992, n28993,
    n28994, n28995, n28996, n28997, n28998, n28999,
    n29000, n29001, n29002, n29003, n29004, n29005,
    n29006, n29007, n29008, n29009, n29010, n29011,
    n29012, n29013, n29014, n29015, n29016, n29017,
    n29018, n29019, n29020, n29021, n29022, n29023,
    n29024, n29025, n29026, n29027, n29028, n29029,
    n29030, n29031, n29032, n29033, n29034, n29035,
    n29036, n29037, n29038, n29039, n29040, n29041,
    n29042, n29043, n29044, n29045, n29046, n29047,
    n29048, n29049, n29050, n29051, n29052, n29053,
    n29054, n29055, n29056, n29057, n29058, n29059,
    n29060, n29061, n29062, n29063, n29064, n29065,
    n29066, n29067, n29068, n29069, n29070, n29071,
    n29072, n29073, n29074, n29075, n29076, n29077,
    n29078, n29079, n29080, n29081, n29082, n29083,
    n29084, n29085, n29086, n29087, n29088, n29089,
    n29090, n29091, n29092, n29093, n29094, n29095,
    n29096, n29097, n29098, n29099, n29100, n29101,
    n29102, n29103, n29104, n29105, n29106, n29107,
    n29108, n29109, n29110, n29111, n29112, n29113,
    n29114, n29115, n29116, n29117, n29118, n29119,
    n29120, n29121, n29122, n29123, n29124, n29125,
    n29126, n29127, n29128, n29129, n29130, n29131,
    n29132, n29133, n29134, n29135, n29136, n29137,
    n29138, n29139, n29140, n29141, n29142, n29143,
    n29144, n29145, n29146, n29147, n29148, n29149,
    n29150, n29151, n29152, n29153, n29154, n29155,
    n29156, n29157, n29158, n29159, n29160, n29161,
    n29162, n29163, n29164, n29165, n29166, n29167,
    n29168, n29169, n29170, n29171, n29172, n29173,
    n29174, n29175, n29176, n29177, n29178, n29179,
    n29180, n29181, n29182, n29183, n29184, n29185,
    n29186, n29187, n29188, n29189, n29190, n29191,
    n29192, n29193, n29194, n29195, n29196, n29197,
    n29198, n29199, n29200, n29201, n29202, n29203,
    n29204, n29205, n29206, n29207, n29208, n29209,
    n29210, n29211, n29212, n29213, n29214, n29215,
    n29216, n29217, n29218, n29219, n29220, n29221,
    n29222, n29223, n29224, n29225, n29226, n29227,
    n29228, n29229, n29230, n29231, n29232, n29233,
    n29234, n29235, n29236, n29237, n29238, n29239,
    n29240, n29241, n29242, n29243, n29244, n29245,
    n29246, n29247, n29248, n29249, n29250, n29251,
    n29252, n29253, n29254, n29255, n29256, n29257,
    n29258, n29259, n29260, n29261, n29262, n29263,
    n29264, n29265, n29266, n29267, n29268, n29269,
    n29270, n29271, n29272, n29273, n29274, n29275,
    n29276, n29277, n29278, n29279, n29280, n29281,
    n29282, n29283, n29284, n29285, n29286, n29287,
    n29288, n29289, n29290, n29291, n29292, n29293,
    n29294, n29295, n29296, n29297, n29298, n29299,
    n29300, n29301, n29302, n29303, n29304, n29305,
    n29306, n29307, n29308, n29309, n29310, n29311,
    n29312, n29313, n29314, n29315, n29316, n29317,
    n29318, n29319, n29320, n29321, n29322, n29323,
    n29324, n29325, n29326, n29327, n29328, n29329,
    n29330, n29331, n29332, n29333, n29334, n29335,
    n29336, n29337, n29338, n29339, n29340, n29341,
    n29342, n29343, n29344, n29345, n29346, n29347,
    n29348, n29349, n29350, n29351, n29352, n29353,
    n29354, n29355, n29356, n29357, n29358, n29359,
    n29360, n29361, n29362, n29363, n29364, n29365,
    n29366, n29367, n29368, n29369, n29370, n29371,
    n29372, n29373, n29374, n29375, n29376, n29377,
    n29378, n29379, n29380, n29381, n29382, n29383,
    n29384, n29385, n29386, n29387, n29388, n29389,
    n29390, n29391, n29392, n29393, n29394, n29395,
    n29396, n29397, n29398, n29399, n29400, n29401,
    n29402, n29403, n29404, n29405, n29406, n29407,
    n29408, n29409, n29410, n29411, n29412, n29413,
    n29414, n29415, n29416, n29417, n29418, n29419,
    n29420, n29421, n29422, n29423, n29424, n29425,
    n29426, n29427, n29428, n29429, n29430, n29431,
    n29432, n29433, n29434, n29435, n29436, n29437,
    n29438, n29439, n29440, n29441, n29442, n29443,
    n29444, n29445, n29446, n29447, n29448, n29449,
    n29450, n29451, n29452, n29453, n29454, n29455,
    n29456, n29457, n29458, n29459, n29460, n29461,
    n29462, n29463, n29464, n29465, n29466, n29467,
    n29468, n29469, n29470, n29471, n29472, n29473,
    n29474, n29475, n29476, n29477, n29478, n29479,
    n29480, n29481, n29482, n29483, n29484, n29485,
    n29486, n29487, n29488, n29489, n29490, n29491,
    n29492, n29493, n29494, n29495, n29496, n29497,
    n29498, n29499, n29500, n29501, n29502, n29503,
    n29504, n29505, n29506, n29507, n29508, n29509,
    n29510, n29511, n29512, n29513, n29514, n29515,
    n29516, n29517, n29518, n29519, n29520, n29521,
    n29522, n29523, n29524, n29525, n29526, n29527,
    n29528, n29529, n29530, n29531, n29532, n29533,
    n29534, n29535, n29536, n29537, n29538, n29539,
    n29540, n29541, n29542, n29543, n29544, n29545,
    n29546, n29547, n29548, n29549, n29550, n29551,
    n29552, n29553, n29554, n29555, n29556, n29557,
    n29558, n29559, n29560, n29561, n29562, n29563,
    n29564, n29565, n29566, n29567, n29568, n29569,
    n29570, n29571, n29572, n29573, n29574, n29575,
    n29576, n29577, n29578, n29579, n29580, n29581,
    n29582, n29583, n29584, n29585, n29586, n29587,
    n29588, n29589, n29590, n29591, n29592, n29593,
    n29594, n29595, n29596, n29597, n29598, n29599,
    n29600, n29601, n29602, n29603, n29604, n29605,
    n29606, n29607, n29608, n29609, n29610, n29611,
    n29612, n29613, n29614, n29615, n29616, n29617,
    n29618, n29619, n29620, n29621, n29622, n29623,
    n29624, n29625, n29626, n29627, n29628, n29629,
    n29630, n29631, n29632, n29633, n29634, n29635,
    n29636, n29637, n29638, n29639, n29640, n29641,
    n29642, n29643, n29644, n29645, n29646, n29647,
    n29648, n29649, n29650, n29651, n29652, n29653,
    n29654, n29655, n29656, n29657, n29658, n29659,
    n29660, n29661, n29662, n29663, n29664, n29665,
    n29666, n29667, n29668, n29669, n29670, n29671,
    n29672, n29673, n29674, n29675, n29676, n29677,
    n29678, n29679, n29680, n29681, n29682, n29683,
    n29684, n29685, n29686, n29687, n29688, n29689,
    n29690, n29691, n29692, n29693, n29694, n29695,
    n29696, n29697, n29698, n29699, n29700, n29701,
    n29702, n29703, n29704, n29705, n29706, n29707,
    n29708, n29709, n29710, n29711, n29712, n29713,
    n29714, n29715, n29716, n29717, n29718, n29719,
    n29720, n29721, n29722, n29723, n29724, n29725,
    n29726, n29727, n29728, n29729, n29730, n29731,
    n29732, n29733, n29734, n29735, n29736, n29737,
    n29738, n29739, n29740, n29741, n29742, n29743,
    n29744, n29745, n29746, n29747, n29748, n29749,
    n29750, n29751, n29752, n29753, n29754, n29755,
    n29756, n29757, n29758, n29759, n29760, n29761,
    n29762, n29763, n29764, n29765, n29766, n29767,
    n29768, n29769, n29770, n29771, n29772, n29773,
    n29774, n29775, n29776, n29777, n29778, n29779,
    n29780, n29781, n29782, n29783, n29784, n29785,
    n29786, n29787, n29788, n29789, n29790, n29791,
    n29792, n29793, n29794, n29795, n29796, n29797,
    n29798, n29799, n29800, n29801, n29802, n29803,
    n29804, n29805, n29806, n29807, n29808, n29809,
    n29810, n29811, n29812, n29813, n29814, n29815,
    n29816, n29817, n29818, n29819, n29820, n29821,
    n29822, n29823, n29824, n29825, n29826, n29827,
    n29828, n29829, n29830, n29831, n29832, n29833,
    n29834, n29835, n29836, n29837, n29838, n29839,
    n29840, n29841, n29842, n29843, n29844, n29845,
    n29846, n29847, n29848, n29849, n29850, n29851,
    n29852, n29853, n29854, n29855, n29856, n29857,
    n29858, n29859, n29860, n29861, n29862, n29863,
    n29864, n29865, n29866, n29867, n29868, n29869,
    n29870, n29871, n29872, n29873, n29874, n29875,
    n29876, n29877, n29878, n29879, n29880, n29881,
    n29882, n29883, n29884, n29885, n29886, n29887,
    n29888, n29889, n29890, n29891, n29892, n29893,
    n29894, n29895, n29896, n29897, n29898, n29899,
    n29900, n29901, n29902, n29903, n29904, n29905,
    n29906, n29907, n29908, n29909, n29910, n29911,
    n29912, n29913, n29914, n29915, n29916, n29917,
    n29918, n29919, n29920, n29921, n29922, n29923,
    n29924, n29925, n29926, n29927, n29928, n29929,
    n29930, n29931, n29932, n29933, n29934, n29935,
    n29936, n29937, n29938, n29939, n29940, n29941,
    n29942, n29943, n29944, n29945, n29946, n29947,
    n29948, n29949, n29950, n29951, n29952, n29953,
    n29954, n29955, n29956, n29957, n29958, n29959,
    n29960, n29961, n29962, n29963, n29964, n29965,
    n29966, n29967, n29968, n29969, n29970, n29971,
    n29972, n29973, n29974, n29975, n29976, n29977,
    n29978, n29979, n29980, n29981, n29982, n29983,
    n29984, n29985, n29986, n29987, n29988, n29989,
    n29990, n29991, n29992, n29993, n29994, n29995,
    n29996, n29997, n29998, n29999, n30000, n30001,
    n30002, n30003, n30004, n30005, n30006, n30007,
    n30008, n30009, n30010, n30011, n30012, n30013,
    n30014, n30015, n30016, n30017, n30018, n30019,
    n30020, n30021, n30022, n30023, n30024, n30025,
    n30026, n30027, n30028, n30029, n30030, n30031,
    n30032, n30033, n30034, n30035, n30036, n30037,
    n30038, n30039, n30040, n30041, n30042, n30043,
    n30044, n30045, n30046, n30047, n30048, n30049,
    n30050, n30051, n30052, n30053, n30054, n30055,
    n30056, n30057, n30058, n30059, n30060, n30061,
    n30062, n30063, n30064, n30065, n30066, n30067,
    n30068, n30069, n30070, n30071, n30072, n30073,
    n30074, n30075, n30076, n30077, n30078, n30079,
    n30080, n30081, n30082, n30083, n30084, n30085,
    n30086, n30087, n30088, n30089, n30090, n30091,
    n30092, n30093, n30094, n30095, n30096, n30097,
    n30098, n30099, n30100, n30101, n30102, n30103,
    n30104, n30105, n30106, n30107, n30108, n30109,
    n30110, n30111, n30112, n30113, n30114, n30115,
    n30116, n30117, n30118, n30119, n30120, n30121,
    n30122, n30123, n30124, n30125, n30126, n30127,
    n30128, n30129, n30130, n30131, n30132, n30133,
    n30134, n30135, n30136, n30137, n30138, n30139,
    n30140, n30141, n30142, n30143, n30144, n30145,
    n30146, n30147, n30148, n30149, n30150, n30151,
    n30152, n30153, n30154, n30155, n30156, n30157,
    n30158, n30159, n30160, n30161, n30162, n30163,
    n30164, n30165, n30166, n30167, n30168, n30169,
    n30170, n30171, n30172, n30173, n30174, n30175,
    n30176, n30177, n30178, n30179, n30180, n30181,
    n30182, n30183, n30184, n30185, n30186, n30187,
    n30188, n30189, n30190, n30191, n30192, n30193,
    n30194, n30195, n30196, n30197, n30198, n30199,
    n30200, n30201, n30202, n30203, n30204, n30205,
    n30206, n30207, n30208, n30209, n30210, n30211,
    n30212, n30213, n30214, n30215, n30216, n30217,
    n30218, n30219, n30220, n30221, n30222, n30223,
    n30224, n30225, n30226, n30227, n30228, n30229,
    n30230, n30231, n30232, n30233, n30234, n30235,
    n30236, n30237, n30238, n30239, n30240, n30241,
    n30242, n30243, n30244, n30245, n30246, n30247,
    n30248, n30249, n30250, n30251, n30252, n30253,
    n30254, n30255, n30256, n30257, n30258, n30259,
    n30260, n30261, n30262, n30263, n30264, n30265,
    n30266, n30267, n30268, n30269, n30270, n30271,
    n30272, n30273, n30274, n30275, n30276, n30277,
    n30278, n30279, n30280, n30281, n30282, n30283,
    n30284, n30285, n30286, n30287, n30288, n30289,
    n30290, n30291, n30292, n30293, n30294, n30295,
    n30296, n30297, n30298, n30299, n30300, n30301,
    n30302, n30303, n30304, n30305, n30306, n30307,
    n30308, n30309, n30310, n30311, n30312, n30313,
    n30314, n30315, n30316, n30317, n30318, n30319,
    n30320, n30321, n30322, n30323, n30324, n30325,
    n30326, n30327, n30328, n30329, n30330, n30331,
    n30332, n30333, n30334, n30335, n30336, n30337,
    n30338, n30339, n30340, n30341, n30342, n30343,
    n30344, n30345, n30346, n30347, n30348, n30349,
    n30350, n30351, n30352, n30353, n30354, n30355,
    n30356, n30357, n30358, n30359, n30360, n30361,
    n30362, n30363, n30364, n30365, n30366, n30367,
    n30368, n30369, n30370, n30371, n30372, n30373,
    n30374, n30375, n30376, n30377, n30378, n30379,
    n30380, n30381, n30382, n30383, n30384, n30385,
    n30386, n30387, n30388, n30389, n30390, n30391,
    n30392, n30393, n30394, n30395, n30396, n30397,
    n30398, n30399, n30400, n30401, n30402, n30403,
    n30404, n30405, n30406, n30407, n30408, n30409,
    n30410, n30411, n30412, n30413, n30414, n30415,
    n30416, n30417, n30418, n30419, n30420, n30421,
    n30422, n30423, n30424, n30425, n30426, n30427,
    n30428, n30429, n30430, n30431, n30432, n30433,
    n30434, n30435, n30436, n30437, n30438, n30439,
    n30440, n30441, n30442, n30443, n30444, n30445,
    n30446, n30447, n30448, n30449, n30450, n30451,
    n30452, n30453, n30454, n30455, n30456, n30457,
    n30458, n30459, n30460, n30461, n30462, n30463,
    n30464, n30465, n30466, n30467, n30468, n30469,
    n30470, n30471, n30472, n30473, n30474, n30475,
    n30476, n30477, n30478, n30479, n30480, n30481,
    n30482, n30483, n30484, n30485, n30486, n30487,
    n30488, n30489, n30490, n30491, n30492, n30493,
    n30494, n30495, n30496, n30497, n30498, n30499,
    n30500, n30501, n30502, n30503, n30504, n30505,
    n30506, n30507, n30508, n30509, n30510, n30511,
    n30512, n30513, n30514, n30515, n30516, n30517,
    n30518, n30519, n30520, n30521, n30522, n30523,
    n30524, n30525, n30526, n30527, n30528, n30529,
    n30530, n30531, n30532, n30533, n30534, n30535,
    n30536, n30537, n30538, n30539, n30540, n30541,
    n30542, n30543, n30544, n30545, n30546, n30547,
    n30548, n30549, n30550, n30551, n30552, n30553,
    n30554, n30555, n30556, n30557, n30558, n30559,
    n30560, n30561, n30562, n30563, n30564, n30565,
    n30566, n30567, n30568, n30569, n30570, n30571,
    n30572, n30573, n30574, n30575, n30576, n30577,
    n30578, n30579, n30580, n30581, n30582, n30583,
    n30584, n30585, n30586, n30587, n30588, n30589,
    n30590, n30591, n30592, n30593, n30594, n30595,
    n30596, n30597, n30598, n30599, n30600, n30601,
    n30602, n30603, n30604, n30605, n30606, n30607,
    n30608, n30609, n30610, n30611, n30612, n30613,
    n30614, n30615, n30616, n30617, n30618, n30619,
    n30620, n30621, n30622, n30623, n30624, n30625,
    n30626, n30627, n30628, n30629, n30630, n30631,
    n30632, n30633, n30634, n30635, n30636, n30637,
    n30638, n30639, n30640, n30641, n30642, n30643,
    n30644, n30645, n30646, n30647, n30648, n30649,
    n30650, n30651, n30652, n30653, n30654, n30655,
    n30656, n30657, n30658, n30659, n30660, n30661,
    n30662, n30663, n30664, n30665, n30666, n30667,
    n30668, n30669, n30670, n30671, n30672, n30673,
    n30674, n30675, n30676, n30677, n30678, n30679,
    n30680, n30681, n30682, n30683, n30684, n30685,
    n30686, n30687, n30688, n30689, n30690, n30691,
    n30692, n30693, n30694, n30695, n30696, n30697,
    n30698, n30699, n30700, n30701, n30702, n30703,
    n30704, n30705, n30706, n30707, n30708, n30709,
    n30710, n30711, n30712, n30713, n30714, n30715,
    n30716, n30717, n30718, n30719, n30720, n30721,
    n30722, n30723, n30724, n30725, n30726, n30727,
    n30728, n30729, n30730, n30731, n30732, n30733,
    n30734, n30735, n30736, n30737, n30738, n30739,
    n30740, n30741, n30742, n30743, n30744, n30745,
    n30746, n30747, n30748, n30749, n30750, n30751,
    n30752, n30753, n30754, n30755, n30756, n30757,
    n30758, n30759, n30760, n30761, n30762, n30763,
    n30764, n30765, n30766, n30767, n30768, n30769,
    n30770, n30771, n30772, n30773, n30774, n30775,
    n30776, n30777, n30778, n30779, n30780, n30781,
    n30782, n30783, n30784, n30785, n30786, n30787,
    n30788, n30789, n30790, n30791, n30792, n30793,
    n30794, n30795, n30796, n30797, n30798, n30799,
    n30800, n30801, n30802, n30803, n30804, n30805,
    n30806, n30807, n30808, n30809, n30810, n30811,
    n30812, n30813, n30814, n30815, n30816, n30817,
    n30818, n30819, n30820, n30821, n30822, n30823,
    n30824, n30825, n30826, n30827, n30828, n30829,
    n30830, n30831, n30832, n30833, n30834, n30835,
    n30836, n30837, n30838, n30839, n30840, n30841,
    n30842, n30843, n30844, n30845, n30846, n30847,
    n30848, n30849, n30850, n30851, n30852, n30853,
    n30854, n30855, n30856, n30857, n30858, n30859,
    n30860, n30861, n30862, n30863, n30864, n30865,
    n30866, n30867, n30868, n30869, n30870, n30871,
    n30872, n30873, n30874, n30875, n30876, n30877,
    n30878, n30879, n30880, n30881, n30882, n30883,
    n30884, n30885, n30886, n30887, n30888, n30889,
    n30890, n30891, n30892, n30893, n30894, n30895,
    n30896, n30897, n30898, n30899, n30900, n30901,
    n30902, n30903, n30904, n30905, n30906, n30907,
    n30908, n30909, n30910, n30911, n30912, n30913,
    n30914, n30915, n30916, n30917, n30918, n30919,
    n30920, n30921, n30922, n30923, n30924, n30925,
    n30926, n30927, n30928, n30929, n30930, n30931,
    n30932, n30933, n30934, n30935, n30936, n30937,
    n30938, n30939, n30940, n30941, n30942, n30943,
    n30944, n30945, n30946, n30947, n30948, n30949,
    n30950, n30951, n30952, n30953, n30954, n30955,
    n30956, n30957, n30958, n30959, n30960, n30961,
    n30962, n30963, n30964, n30965, n30966, n30967,
    n30968, n30969, n30970, n30971, n30972, n30973,
    n30974, n30975, n30976, n30977, n30978, n30979,
    n30980, n30981, n30982, n30983, n30984, n30985,
    n30986, n30987, n30988, n30989, n30990, n30991,
    n30992, n30993, n30994, n30995, n30996, n30997,
    n30998, n30999, n31000, n31001, n31002, n31003,
    n31004, n31005, n31006, n31007, n31008, n31009,
    n31010, n31011, n31012, n31013, n31014, n31015,
    n31016, n31017, n31018, n31019, n31020, n31021,
    n31022, n31023, n31024, n31025, n31026, n31027,
    n31028, n31029, n31030, n31031, n31032, n31033,
    n31034, n31035, n31036, n31037, n31038, n31039,
    n31040, n31041, n31042, n31043, n31044, n31045,
    n31046, n31047, n31048, n31049, n31050, n31051,
    n31052, n31053, n31054, n31055, n31056, n31057,
    n31058, n31059, n31060, n31061, n31062, n31063,
    n31064, n31065, n31066, n31067, n31068, n31069,
    n31070, n31071, n31072, n31073, n31074, n31075,
    n31076, n31077, n31078, n31079, n31080, n31081,
    n31082, n31083, n31084, n31085, n31086, n31087,
    n31088, n31089, n31090, n31091, n31092, n31093,
    n31094, n31095, n31096, n31097, n31098, n31099,
    n31100, n31101, n31102, n31103, n31104, n31105,
    n31106, n31107, n31108, n31109, n31110, n31111,
    n31112, n31113, n31114, n31115, n31116, n31117,
    n31118, n31119, n31120, n31121, n31122, n31123,
    n31124, n31125, n31126, n31127, n31128, n31129,
    n31130, n31131, n31132, n31133, n31134, n31135,
    n31136, n31137, n31138, n31139, n31140, n31141,
    n31142, n31143, n31144, n31145, n31146, n31147,
    n31148, n31149, n31150, n31151, n31152, n31153,
    n31154, n31155, n31156, n31157, n31158, n31159,
    n31160, n31161, n31162, n31163, n31164, n31165,
    n31166, n31167, n31168, n31169, n31170, n31171,
    n31172, n31173, n31174, n31175, n31176, n31177,
    n31178, n31179, n31180, n31181, n31182, n31183,
    n31184, n31185, n31186, n31187, n31188, n31189,
    n31190, n31191, n31192, n31193, n31194, n31195,
    n31196, n31197, n31198, n31199, n31200, n31201,
    n31202, n31203, n31204, n31205, n31206, n31207,
    n31208, n31209, n31210, n31211, n31212, n31213,
    n31214, n31215, n31216, n31217, n31218, n31219,
    n31220, n31221, n31222, n31223, n31224, n31225,
    n31226, n31227, n31228, n31229, n31230, n31231,
    n31232, n31233, n31234, n31235, n31236, n31237,
    n31238, n31239, n31240, n31241, n31242, n31243,
    n31244, n31245, n31246, n31247, n31248, n31249,
    n31250, n31251, n31252, n31253, n31254, n31255,
    n31256, n31257, n31258, n31259, n31260, n31261,
    n31262, n31263, n31264, n31265, n31266, n31267,
    n31268, n31269, n31270, n31271, n31272, n31273,
    n31274, n31275, n31276, n31277, n31278, n31279,
    n31280, n31281, n31282, n31283, n31284, n31285,
    n31286, n31287, n31288, n31289, n31290, n31291,
    n31292, n31293, n31294, n31295, n31296, n31297,
    n31298, n31299, n31300, n31301, n31302, n31303,
    n31304, n31305, n31306, n31307, n31308, n31309,
    n31310, n31311, n31312, n31313, n31314, n31315,
    n31316, n31317, n31318, n31319, n31320, n31321,
    n31322, n31323, n31324, n31325, n31326, n31327,
    n31328, n31329, n31330, n31331, n31332, n31333,
    n31334, n31335, n31336, n31337, n31338, n31339,
    n31340, n31341, n31342, n31343, n31344, n31345,
    n31346, n31347, n31348, n31349, n31350, n31351,
    n31352, n31353, n31354, n31355, n31356, n31357,
    n31358, n31359, n31360, n31361, n31362, n31363,
    n31364, n31365, n31366, n31367, n31368, n31369,
    n31370, n31371, n31372, n31373, n31374, n31375,
    n31376, n31377, n31378, n31379, n31380, n31381,
    n31382, n31383, n31384, n31385, n31386, n31387,
    n31388, n31389, n31390, n31391, n31392, n31393,
    n31394, n31395, n31396, n31397, n31398, n31399,
    n31400, n31401, n31402, n31403, n31404, n31405,
    n31406, n31407, n31408, n31409, n31410, n31411,
    n31412, n31413, n31414, n31415, n31416, n31417,
    n31418, n31419, n31420, n31421, n31422, n31423,
    n31424, n31425, n31426, n31427, n31428, n31429,
    n31430, n31431, n31432, n31433, n31434, n31435,
    n31436, n31437, n31438, n31439, n31440, n31441,
    n31442, n31443, n31444, n31445, n31446, n31447,
    n31448, n31449, n31450, n31451, n31452, n31453,
    n31454, n31455, n31456, n31457, n31458, n31459,
    n31460, n31461, n31462, n31463, n31464, n31465,
    n31466, n31467, n31468, n31469, n31470, n31471,
    n31472, n31473, n31474, n31475, n31476, n31477,
    n31478, n31479, n31480, n31481, n31482, n31483,
    n31484, n31485, n31486, n31487, n31488, n31489,
    n31490, n31491, n31492, n31493, n31494, n31495,
    n31496, n31497, n31498, n31499, n31500, n31501,
    n31502, n31503, n31504, n31505, n31506, n31507,
    n31508, n31509, n31510, n31511, n31512, n31513,
    n31514, n31515, n31516, n31517, n31518, n31519,
    n31520, n31521, n31522, n31523, n31524, n31525,
    n31526, n31527, n31528, n31529, n31530, n31531,
    n31532, n31533, n31534, n31535, n31536, n31537,
    n31538, n31539, n31540, n31541, n31542, n31543,
    n31544, n31545, n31546, n31547, n31548, n31549,
    n31550, n31551, n31552, n31553, n31554, n31555,
    n31556, n31557, n31558, n31559, n31560, n31561,
    n31562, n31563, n31564, n31565, n31566, n31567,
    n31568, n31569, n31570, n31571, n31572, n31573,
    n31574, n31575, n31576, n31577, n31578, n31579,
    n31580, n31581, n31582, n31583, n31584, n31585,
    n31586, n31587, n31588, n31589, n31590, n31591,
    n31592, n31593, n31594, n31595, n31596, n31597,
    n31598, n31599, n31600, n31601, n31602, n31603,
    n31604, n31605, n31606, n31607, n31608, n31609,
    n31610, n31611, n31612, n31613, n31614, n31615,
    n31616, n31617, n31618, n31619, n31620, n31621,
    n31622, n31623, n31624, n31625, n31626, n31627,
    n31628, n31629, n31630, n31631, n31632, n31633,
    n31634, n31635, n31636, n31637, n31638, n31639,
    n31640, n31641, n31642, n31643, n31644, n31645,
    n31646, n31647, n31648, n31649, n31650, n31651,
    n31652, n31653, n31654, n31655, n31656, n31657,
    n31658, n31659, n31660, n31661, n31662, n31663,
    n31664, n31665, n31666, n31667, n31668, n31669,
    n31670, n31671, n31672, n31673, n31674, n31675,
    n31676, n31677, n31678, n31679, n31680, n31681,
    n31682, n31683, n31684, n31685, n31686, n31687,
    n31688, n31689, n31690, n31691, n31692, n31693,
    n31694, n31695, n31696, n31697, n31698, n31699,
    n31700, n31701, n31702, n31703, n31704, n31705,
    n31706, n31707, n31708, n31709, n31710, n31711,
    n31712, n31713, n31714, n31715, n31716, n31717,
    n31718, n31719, n31720, n31721, n31722, n31723,
    n31724, n31725, n31726, n31727, n31728, n31729,
    n31730, n31731, n31732, n31733, n31734, n31735,
    n31736, n31737, n31738, n31739, n31740, n31741,
    n31742, n31743, n31744, n31745, n31746, n31747,
    n31748, n31749, n31750, n31751, n31752, n31753,
    n31754, n31755, n31756, n31757, n31758, n31759,
    n31760, n31761, n31762, n31763, n31764, n31765,
    n31766, n31767, n31768, n31769, n31770, n31771,
    n31772, n31773, n31774, n31775, n31776, n31777,
    n31778, n31779, n31780, n31781, n31782, n31783,
    n31784, n31785, n31786, n31787, n31788, n31789,
    n31790, n31791, n31792, n31793, n31794, n31795,
    n31796, n31797, n31798, n31799, n31800, n31801,
    n31802, n31803, n31804, n31805, n31806, n31807,
    n31808, n31809, n31810, n31811, n31812, n31813,
    n31814, n31815, n31816, n31817, n31818, n31819,
    n31820, n31821, n31822, n31823, n31824, n31825,
    n31826, n31827, n31828, n31829, n31830, n31831,
    n31832, n31833, n31834, n31835, n31836, n31837,
    n31838, n31839, n31840, n31841, n31842, n31843,
    n31844, n31845, n31846, n31847, n31848, n31849,
    n31850, n31851, n31852, n31853, n31854, n31855,
    n31856, n31857, n31858, n31859, n31860, n31861,
    n31862, n31863, n31864, n31865, n31866, n31867,
    n31868, n31869, n31870, n31871, n31872, n31873,
    n31874, n31875, n31876, n31877, n31878, n31879,
    n31880, n31881, n31882, n31883, n31884, n31885,
    n31886, n31887, n31888, n31889, n31890, n31891,
    n31892, n31893, n31894, n31895, n31896, n31897,
    n31898, n31899, n31900, n31901, n31902, n31903,
    n31904, n31905, n31906, n31907, n31908, n31909,
    n31910, n31911, n31912, n31913, n31914, n31915,
    n31916, n31917, n31918, n31919, n31920, n31921,
    n31922, n31923, n31924, n31925, n31926, n31927,
    n31928, n31929, n31930, n31931, n31932, n31933,
    n31934, n31935, n31936, n31937, n31938, n31939,
    n31940, n31941, n31942, n31943, n31944, n31945,
    n31946, n31947, n31948, n31949, n31950, n31951,
    n31952, n31953, n31954, n31955, n31956, n31957,
    n31958, n31959, n31960, n31961, n31962, n31963,
    n31964, n31965, n31966, n31967, n31968, n31969,
    n31970, n31971, n31972, n31973, n31974, n31975,
    n31976, n31977, n31978, n31979, n31980, n31981,
    n31982, n31983, n31984, n31985, n31986, n31987,
    n31988, n31989, n31990, n31991, n31992, n31993,
    n31994, n31995, n31996, n31997, n31998, n31999,
    n32000, n32001, n32002, n32003, n32004, n32005,
    n32006, n32007, n32008, n32009, n32010, n32011,
    n32012, n32013, n32014, n32015, n32016, n32017,
    n32018, n32019, n32020, n32021, n32022, n32023,
    n32024, n32025, n32026, n32027, n32028, n32029,
    n32030, n32031, n32032, n32033, n32034, n32035,
    n32036, n32037, n32038, n32039, n32040, n32041,
    n32042, n32043, n32044, n32045, n32046, n32047,
    n32048, n32049, n32050, n32051, n32052, n32053,
    n32054, n32055, n32056, n32057, n32058, n32059,
    n32060, n32061, n32062, n32063, n32064, n32065,
    n32066, n32067, n32068, n32069, n32070, n32071,
    n32072, n32073, n32074, n32075, n32076, n32077,
    n32078, n32079, n32080, n32081, n32082, n32083,
    n32084, n32085, n32086, n32087, n32088, n32089,
    n32090, n32091, n32092, n32093, n32094, n32095,
    n32096, n32097, n32098, n32099, n32100, n32101,
    n32102, n32103, n32104, n32105, n32106, n32107,
    n32108, n32109, n32110, n32111, n32112, n32113,
    n32114, n32115, n32116, n32117, n32118, n32119,
    n32120, n32121, n32122, n32123, n32124, n32125,
    n32126, n32127, n32128, n32129, n32130, n32131,
    n32132, n32133, n32134, n32135, n32136, n32137,
    n32138, n32139, n32140, n32141, n32142, n32143,
    n32144, n32145, n32146, n32147, n32148, n32149,
    n32150, n32151, n32152, n32153, n32154, n32155,
    n32156, n32157, n32158, n32159, n32160, n32161,
    n32162, n32163, n32164, n32165, n32166, n32167,
    n32168, n32169, n32170, n32171, n32172, n32173,
    n32174, n32175, n32176, n32177, n32178, n32179,
    n32180, n32181, n32182, n32183, n32184, n32185,
    n32186, n32187, n32188, n32189, n32190, n32191,
    n32192, n32193, n32194, n32195, n32196, n32197,
    n32198, n32199, n32200, n32201, n32202, n32203,
    n32204, n32205, n32206, n32207, n32208, n32209,
    n32210, n32211, n32212, n32213, n32214, n32215,
    n32216, n32217, n32218, n32219, n32220, n32221,
    n32222, n32223, n32224, n32225, n32226, n32227,
    n32228, n32229, n32230, n32231, n32232, n32233,
    n32234, n32235, n32236, n32237, n32238, n32239,
    n32240, n32241, n32242, n32243, n32244, n32245,
    n32246, n32247, n32248, n32249, n32250, n32251,
    n32252, n32253, n32254, n32255, n32256, n32257,
    n32258, n32259, n32260, n32261, n32262, n32263,
    n32264, n32265, n32266, n32267, n32268, n32269,
    n32270, n32271, n32272, n32273, n32274, n32275,
    n32276, n32277, n32278, n32279, n32280, n32281,
    n32282, n32283, n32284, n32285, n32286, n32287,
    n32288, n32289, n32290, n32291, n32292, n32293,
    n32294, n32295, n32296, n32297, n32298, n32299,
    n32300, n32301, n32302, n32303, n32304, n32305,
    n32306, n32307, n32308, n32309, n32310, n32311,
    n32312, n32313, n32314, n32315, n32316, n32317,
    n32318, n32319, n32320, n32321, n32322, n32323,
    n32324, n32325, n32326, n32327, n32328, n32329,
    n32330, n32331, n32332, n32333, n32334, n32335,
    n32336, n32337, n32338, n32339, n32340, n32341,
    n32342, n32343, n32344, n32345, n32346, n32347,
    n32348, n32349, n32350, n32351, n32352, n32353,
    n32354, n32355, n32356, n32357, n32358, n32359,
    n32360, n32361, n32362, n32363, n32364, n32365,
    n32366, n32367, n32368, n32369, n32370, n32371,
    n32372, n32373, n32374, n32375, n32376, n32377,
    n32378, n32379, n32380, n32381, n32382, n32383,
    n32384, n32385, n32386, n32387, n32388, n32389,
    n32390, n32391, n32392, n32393, n32394, n32395,
    n32396, n32397, n32398, n32399, n32400, n32401,
    n32402, n32403, n32404, n32405, n32406, n32407,
    n32408, n32409, n32410, n32411, n32412, n32413,
    n32414, n32415, n32416, n32417, n32418, n32419,
    n32420, n32421, n32422, n32423, n32424, n32425,
    n32426, n32427, n32428, n32429, n32430, n32431,
    n32432, n32433, n32434, n32435, n32436, n32437,
    n32438, n32439, n32440, n32441, n32442, n32443,
    n32444, n32445, n32446, n32447, n32448, n32449,
    n32450, n32451, n32452, n32453, n32454, n32455,
    n32456, n32457, n32458, n32459, n32460, n32461,
    n32462, n32463, n32464, n32465, n32466, n32467,
    n32468, n32469, n32470, n32471, n32472, n32473,
    n32474, n32475, n32476, n32477, n32478, n32479,
    n32480, n32481, n32482, n32483, n32484, n32485,
    n32486, n32487, n32488, n32489, n32490, n32491,
    n32492, n32493, n32494, n32495, n32496, n32497,
    n32498, n32499, n32500, n32501, n32502, n32503,
    n32504, n32505, n32506, n32507, n32508, n32509,
    n32510, n32511, n32512, n32513, n32514, n32515,
    n32516, n32517, n32518, n32519, n32520, n32521,
    n32522, n32523, n32524, n32525, n32526, n32527,
    n32528, n32529, n32530, n32531, n32532, n32533,
    n32534, n32535, n32536, n32537, n32538, n32539,
    n32540, n32541, n32542, n32543, n32544, n32545,
    n32546, n32547, n32548, n32549, n32550, n32551,
    n32552, n32553, n32554, n32555, n32556, n32557,
    n32558, n32559, n32560, n32561, n32562, n32563,
    n32564, n32565, n32566, n32567, n32568, n32569,
    n32570, n32571, n32572, n32573, n32574, n32575,
    n32576, n32577, n32578, n32579, n32580, n32581,
    n32582, n32583, n32584, n32585, n32586, n32587,
    n32588, n32589, n32590, n32591, n32592, n32593,
    n32594, n32595, n32596, n32597, n32598, n32599,
    n32600, n32601, n32602, n32603, n32604, n32605,
    n32606, n32607, n32608, n32609, n32610, n32611,
    n32612, n32613, n32614, n32615, n32616, n32617,
    n32618, n32619, n32620, n32621, n32622, n32623,
    n32624, n32625, n32626, n32627, n32628, n32629,
    n32630, n32631, n32632, n32633, n32634, n32635,
    n32636, n32637, n32638, n32639, n32640, n32641,
    n32642, n32643, n32644, n32645, n32646, n32647,
    n32648, n32649, n32650, n32651, n32652, n32653,
    n32654, n32655, n32656, n32657, n32658, n32659,
    n32660, n32661, n32662, n32663, n32664, n32665,
    n32666, n32667, n32668, n32669, n32670, n32671,
    n32672, n32673, n32674, n32675, n32676, n32677,
    n32678, n32679, n32680, n32681, n32682, n32683,
    n32684, n32685, n32686, n32687, n32688, n32689,
    n32690, n32691, n32692, n32693, n32694, n32695,
    n32696, n32697, n32698, n32699, n32700, n32701,
    n32702, n32703, n32704, n32705, n32706, n32707,
    n32708, n32709, n32710, n32711, n32712, n32713,
    n32714, n32715, n32716, n32717, n32718, n32719,
    n32720, n32721, n32722, n32723, n32724, n32725,
    n32726, n32727, n32728, n32729, n32730, n32731,
    n32732, n32733, n32734, n32735, n32736, n32737,
    n32738, n32739, n32740, n32741, n32742, n32743,
    n32744, n32745, n32746, n32747, n32748, n32749,
    n32750, n32751, n32752, n32753, n32754, n32755,
    n32756, n32757, n32758, n32759, n32760, n32761,
    n32762, n32763, n32764, n32765, n32766, n32767,
    n32768, n32769, n32770, n32771, n32772, n32773,
    n32774, n32775, n32776, n32777, n32778, n32779,
    n32780, n32781, n32782, n32783, n32784, n32785,
    n32786, n32787, n32788, n32789, n32790, n32791,
    n32792, n32793, n32794, n32795, n32796, n32797,
    n32798, n32799, n32800, n32801, n32802, n32803,
    n32804, n32805, n32806, n32807, n32808, n32809,
    n32810, n32811, n32812, n32813, n32814, n32815,
    n32816, n32817, n32818, n32819, n32820, n32821,
    n32822, n32823, n32824, n32825, n32826, n32827,
    n32828, n32829, n32830, n32831, n32832, n32833,
    n32834, n32835, n32836, n32837, n32838, n32839,
    n32840, n32841, n32842, n32843, n32844, n32845,
    n32846, n32847, n32848, n32849, n32850, n32851,
    n32852, n32853, n32854, n32855, n32856, n32857,
    n32858, n32859, n32860, n32861, n32862, n32863,
    n32864, n32865, n32866, n32867, n32868, n32869,
    n32870, n32871, n32872, n32873, n32874, n32875,
    n32876, n32877, n32878, n32879, n32880, n32881,
    n32882, n32883, n32884, n32885, n32886, n32887,
    n32888, n32889, n32890, n32891, n32892, n32893,
    n32894, n32895, n32896, n32897, n32898, n32899,
    n32900, n32901, n32902, n32903, n32904, n32905,
    n32906, n32907, n32908, n32909, n32910, n32911,
    n32912, n32913, n32914, n32915, n32916, n32917,
    n32918, n32919, n32920, n32921, n32922, n32923,
    n32924, n32925, n32926, n32927, n32928, n32929,
    n32930, n32931, n32932, n32933, n32934, n32935,
    n32936, n32937, n32938, n32939, n32940, n32941,
    n32942, n32943, n32944, n32945, n32946, n32947,
    n32948, n32949, n32950, n32951, n32952, n32953,
    n32954, n32955, n32956, n32957, n32958, n32959,
    n32960, n32961, n32962, n32963, n32964, n32965,
    n32966, n32967, n32968, n32969, n32970, n32971,
    n32972, n32973, n32974, n32975, n32976, n32977,
    n32978, n32979, n32980, n32981, n32982, n32983,
    n32984, n32985, n32986, n32987, n32988, n32989,
    n32990, n32991, n32992, n32993, n32994, n32995,
    n32996, n32997, n32998, n32999, n33000, n33001,
    n33002, n33003, n33004, n33005, n33006, n33007,
    n33008, n33009, n33010, n33011, n33012, n33013,
    n33014, n33015, n33016, n33017, n33018, n33019,
    n33020, n33021, n33022, n33023, n33024, n33025,
    n33026, n33027, n33028, n33029, n33030, n33031,
    n33032, n33033, n33034, n33035, n33036, n33037,
    n33038, n33039, n33040, n33041, n33042, n33043,
    n33044, n33045, n33046, n33047, n33048, n33049,
    n33050, n33051, n33052, n33053, n33054, n33055,
    n33056, n33057, n33058, n33059, n33060, n33061,
    n33062, n33063, n33064, n33065, n33066, n33067,
    n33068, n33069, n33070, n33071, n33072, n33073,
    n33074, n33075, n33076, n33077, n33078, n33079,
    n33080, n33081, n33082, n33083, n33084, n33085,
    n33086, n33087, n33088, n33089, n33090, n33091,
    n33092, n33093, n33094, n33095, n33096, n33097,
    n33098, n33099, n33100, n33101, n33102, n33103,
    n33104, n33105, n33106, n33107, n33108, n33109,
    n33110, n33111, n33112, n33113, n33114, n33115,
    n33116, n33117, n33118, n33119, n33120, n33121,
    n33122, n33123, n33124, n33125, n33126, n33127,
    n33128, n33129, n33130, n33131, n33132, n33133,
    n33134, n33135, n33136, n33137, n33138, n33139,
    n33140, n33141, n33142, n33143, n33144, n33145,
    n33146, n33147, n33148, n33149, n33150, n33151,
    n33152, n33153, n33154, n33155, n33156, n33157,
    n33158, n33159, n33160, n33161, n33162, n33163,
    n33164, n33165, n33166, n33167, n33168, n33169,
    n33170, n33171, n33172, n33173, n33174, n33175,
    n33176, n33177, n33178, n33179, n33180, n33181,
    n33182, n33183, n33184, n33185, n33186, n33187,
    n33188, n33189, n33190, n33191, n33192, n33193,
    n33194, n33195, n33196, n33197, n33198, n33199,
    n33200, n33201, n33202, n33203, n33204, n33205,
    n33206, n33207, n33208, n33209, n33210, n33211,
    n33212, n33213, n33214, n33215, n33216, n33217,
    n33218, n33219, n33220, n33221, n33222, n33223,
    n33224, n33225, n33226, n33227, n33228, n33229,
    n33230, n33231, n33232, n33233, n33234, n33235,
    n33236, n33237, n33238, n33239, n33240, n33241,
    n33242, n33243, n33244, n33245, n33246, n33247,
    n33248, n33249, n33250, n33251, n33252, n33253,
    n33254, n33255, n33256, n33257, n33258, n33259,
    n33260, n33261, n33262, n33263, n33264, n33265,
    n33266, n33267, n33268, n33269, n33270, n33271,
    n33272, n33273, n33274, n33275, n33276, n33277,
    n33278, n33279, n33280, n33281, n33282, n33283,
    n33284, n33285, n33286, n33287, n33288, n33289,
    n33290, n33291, n33292, n33293, n33294, n33295,
    n33296, n33297, n33298, n33299, n33300, n33301,
    n33302, n33303, n33304, n33305, n33306, n33307,
    n33308, n33309, n33310, n33311, n33312, n33313,
    n33314, n33315, n33316, n33317, n33318, n33319,
    n33320, n33321, n33322, n33323, n33324, n33325,
    n33326, n33327, n33328, n33329, n33330, n33331,
    n33332, n33333, n33334, n33335, n33336, n33337,
    n33338, n33339, n33340, n33341, n33342, n33343,
    n33344, n33345, n33346, n33347, n33348, n33349,
    n33350, n33351, n33352, n33353, n33354, n33355,
    n33356, n33357, n33358, n33359, n33360, n33361,
    n33362, n33363, n33364, n33365, n33366, n33367,
    n33368, n33369, n33370, n33371, n33372, n33373,
    n33374, n33375, n33376, n33377, n33378, n33379,
    n33380, n33381, n33382, n33383, n33384, n33385,
    n33386, n33387, n33388, n33389, n33390, n33391,
    n33392, n33393, n33394, n33395, n33396, n33397,
    n33398, n33399, n33400, n33401, n33402, n33403,
    n33404, n33405, n33406, n33407, n33408, n33409,
    n33410, n33411, n33412, n33413, n33414, n33415,
    n33416, n33417, n33418, n33419, n33420, n33421,
    n33422, n33423, n33424, n33425, n33426, n33427,
    n33428, n33429, n33430, n33431, n33432, n33433,
    n33434, n33435, n33436, n33437, n33438, n33439,
    n33440, n33441, n33442, n33443, n33444, n33445,
    n33446, n33447, n33448, n33449, n33450, n33451,
    n33452, n33453, n33454, n33455, n33456, n33457,
    n33458, n33459, n33460, n33461, n33462, n33463,
    n33464, n33465, n33466, n33467, n33468, n33469,
    n33470, n33471, n33472, n33473, n33474, n33475,
    n33476, n33477, n33478, n33479, n33480, n33481,
    n33482, n33483, n33484, n33485, n33486, n33487,
    n33488, n33489, n33490, n33491, n33492, n33493,
    n33494, n33495, n33496, n33497, n33498, n33499,
    n33500, n33501, n33502, n33503, n33504, n33505,
    n33506, n33507, n33508, n33509, n33510, n33511,
    n33512, n33513, n33514, n33515, n33516, n33517,
    n33518, n33519, n33520, n33521, n33522, n33523,
    n33524, n33525, n33526, n33527, n33528, n33529,
    n33530, n33531, n33532, n33533, n33534, n33535,
    n33536, n33537, n33538, n33539, n33540, n33541,
    n33542, n33543, n33544, n33545, n33546, n33547,
    n33548, n33549, n33550, n33551, n33552, n33553,
    n33554, n33555, n33556, n33557, n33558, n33559,
    n33560, n33561, n33562, n33563, n33564, n33565,
    n33566, n33567, n33568, n33569, n33570, n33571,
    n33572, n33573, n33574, n33575, n33576, n33577,
    n33578, n33579, n33580, n33581, n33582, n33583,
    n33584, n33585, n33586, n33587, n33588, n33589,
    n33590, n33591, n33592, n33593, n33594, n33595,
    n33596, n33597, n33598, n33599, n33600, n33601,
    n33602, n33603, n33604, n33605, n33606, n33607,
    n33608, n33609, n33610, n33611, n33612, n33613,
    n33614, n33615, n33616, n33617, n33618, n33619,
    n33620, n33621, n33622, n33623, n33624, n33625,
    n33626, n33627, n33628, n33629, n33630, n33631,
    n33632, n33633, n33634, n33635, n33636, n33637,
    n33638, n33639, n33640, n33641, n33642, n33643,
    n33644, n33645, n33646, n33647, n33648, n33649,
    n33650, n33651, n33652, n33653, n33654, n33655,
    n33656, n33657, n33658, n33659, n33660, n33661,
    n33662, n33663, n33664, n33665, n33666, n33667,
    n33668, n33669, n33670, n33671, n33672, n33673,
    n33674, n33675, n33676, n33677, n33678, n33679,
    n33680, n33681, n33682, n33683, n33684, n33685,
    n33686, n33687, n33688, n33689, n33690, n33691,
    n33692, n33693, n33694, n33695, n33696, n33697,
    n33698, n33699, n33700, n33701, n33702, n33703,
    n33704, n33705, n33706, n33707, n33708, n33709,
    n33710, n33711, n33712, n33713, n33714, n33715,
    n33716, n33717, n33718, n33719, n33720, n33721,
    n33722, n33723, n33724, n33725, n33726, n33727,
    n33728, n33729, n33730, n33731, n33732, n33733,
    n33734, n33735, n33736, n33737, n33738, n33739,
    n33740, n33741, n33742, n33743, n33744, n33745,
    n33746, n33747, n33748, n33749, n33750, n33751,
    n33752, n33753, n33754, n33755, n33756, n33757,
    n33758, n33759, n33760, n33761, n33762, n33763,
    n33764, n33765, n33766, n33767, n33768, n33769,
    n33770, n33771, n33772, n33773, n33774, n33775,
    n33776, n33777, n33778, n33779, n33780, n33781,
    n33782, n33783, n33784, n33785, n33786, n33787,
    n33788, n33789, n33790, n33791, n33792, n33793,
    n33794, n33795, n33796, n33797, n33798, n33799,
    n33800, n33801, n33802, n33803, n33804, n33805,
    n33806, n33807, n33808, n33809, n33810, n33811,
    n33812, n33813, n33814, n33815, n33816, n33817,
    n33818, n33819, n33820, n33821, n33822, n33823,
    n33824, n33825, n33826, n33827, n33828, n33829,
    n33830, n33831, n33832, n33833, n33834, n33835,
    n33836, n33837, n33838, n33839, n33840, n33841,
    n33842, n33843, n33844, n33845, n33846, n33847,
    n33848, n33849, n33850, n33851, n33852, n33853,
    n33854, n33855, n33856, n33857, n33858, n33859,
    n33860, n33861, n33862, n33863, n33864, n33865,
    n33866, n33867, n33868, n33869, n33870, n33871,
    n33872, n33873, n33874, n33875, n33876, n33877,
    n33878, n33879, n33880, n33881, n33882, n33883,
    n33884, n33885, n33886, n33887, n33888, n33889,
    n33890, n33891, n33892, n33893, n33894, n33895,
    n33896, n33897, n33898, n33899, n33900, n33901,
    n33902, n33903, n33904, n33905, n33906, n33907,
    n33908, n33909, n33910, n33911, n33912, n33913,
    n33914, n33915, n33916, n33917, n33918, n33919,
    n33920, n33921, n33922, n33923, n33924, n33925,
    n33926, n33927, n33928, n33929, n33930, n33931,
    n33932, n33933, n33934, n33935, n33936, n33937,
    n33938, n33939, n33940, n33941, n33942, n33943,
    n33944, n33945, n33946, n33947, n33948, n33949,
    n33950, n33951, n33952, n33953, n33954, n33955,
    n33956, n33957, n33958, n33959, n33960, n33961,
    n33962, n33963, n33964, n33965, n33966, n33967,
    n33968, n33969, n33970, n33971, n33972, n33973,
    n33974, n33975, n33976, n33977, n33978, n33979,
    n33980, n33981, n33982, n33983, n33984, n33985,
    n33986, n33987, n33988, n33989, n33990, n33991,
    n33992, n33993, n33994, n33995, n33996, n33997,
    n33998, n33999, n34000, n34001, n34002, n34003,
    n34004, n34005, n34006, n34007, n34008, n34009,
    n34010, n34011, n34012, n34013, n34014, n34015,
    n34016, n34017, n34018, n34019, n34020, n34021,
    n34022, n34023, n34024, n34025, n34026, n34027,
    n34028, n34029, n34030, n34031, n34032, n34033,
    n34034, n34035, n34036, n34037, n34038, n34039,
    n34040, n34041, n34042, n34043, n34044, n34045,
    n34046, n34047, n34048, n34049, n34050, n34051,
    n34052, n34053, n34054, n34055, n34056, n34057,
    n34058, n34059, n34060, n34061, n34062, n34063,
    n34064, n34065, n34066, n34067, n34068, n34069,
    n34070, n34071, n34072, n34073, n34074, n34075,
    n34076, n34077, n34078, n34079, n34080, n34081,
    n34082, n34083, n34084, n34085, n34086, n34087,
    n34088, n34089, n34090, n34091, n34092, n34093,
    n34094, n34095, n34096, n34097, n34098, n34099,
    n34100, n34101, n34102, n34103, n34104, n34105,
    n34106, n34107, n34108, n34109, n34110, n34111,
    n34112, n34113, n34114, n34115, n34116, n34117,
    n34118, n34119, n34120, n34121, n34122, n34123,
    n34124, n34125, n34126, n34127, n34128, n34129,
    n34130, n34131, n34132, n34133, n34134, n34135,
    n34136, n34137, n34138, n34139, n34140, n34141,
    n34142, n34143, n34144, n34145, n34146, n34147,
    n34148, n34149, n34150, n34151, n34152, n34153,
    n34154, n34155, n34156, n34157, n34158, n34159,
    n34160, n34161, n34162, n34163, n34164, n34165,
    n34166, n34167, n34168, n34169, n34170, n34171,
    n34172, n34173, n34174, n34175, n34176, n34177,
    n34178, n34179, n34180, n34181, n34182, n34183,
    n34184, n34185, n34186, n34187, n34188, n34189,
    n34190, n34191, n34192, n34193, n34194, n34195,
    n34196, n34197, n34198, n34199, n34200, n34201,
    n34202, n34203, n34204, n34205, n34206, n34207,
    n34208, n34209, n34210, n34211, n34212, n34213,
    n34214, n34215, n34216, n34217, n34218, n34219,
    n34220, n34221, n34222, n34223, n34224, n34225,
    n34226, n34227, n34228, n34229, n34230, n34231,
    n34232, n34233, n34234, n34235, n34236, n34237,
    n34238, n34239, n34240, n34241, n34242, n34243,
    n34244, n34245, n34246, n34247, n34248, n34249,
    n34250, n34251, n34252, n34253, n34254, n34255,
    n34256, n34257, n34258, n34259, n34260, n34261,
    n34262, n34263, n34264, n34265, n34266, n34267,
    n34268, n34269, n34270, n34271, n34272, n34273,
    n34274, n34275, n34276, n34277, n34278, n34279,
    n34280, n34281, n34282, n34283, n34284, n34285,
    n34286, n34287, n34288, n34289, n34290, n34291,
    n34292, n34293, n34294, n34295, n34296, n34297,
    n34298, n34299, n34300, n34301, n34302, n34303,
    n34304, n34305, n34306, n34307, n34308, n34309,
    n34310, n34311, n34312, n34313, n34314, n34315,
    n34316, n34317, n34318, n34319, n34320, n34321,
    n34322, n34323, n34324, n34325, n34326, n34327,
    n34328, n34329, n34330, n34331, n34332, n34333,
    n34334, n34335, n34336, n34337, n34338, n34339,
    n34340, n34341, n34342, n34343, n34344, n34345,
    n34346, n34347, n34348, n34349, n34350, n34351,
    n34352, n34353, n34354, n34355, n34356, n34357,
    n34358, n34359, n34360, n34361, n34362, n34363,
    n34364, n34365, n34366, n34367, n34368, n34369,
    n34370, n34371, n34372, n34373, n34374, n34375,
    n34376, n34377, n34378, n34379, n34380, n34381,
    n34382, n34383, n34384, n34385, n34386, n34387,
    n34388, n34389, n34390, n34391, n34392, n34393,
    n34394, n34395, n34396, n34397, n34398, n34399,
    n34400, n34401, n34402, n34403, n34404, n34405,
    n34406, n34407, n34408, n34409, n34410, n34411,
    n34412, n34413, n34414, n34415, n34416, n34417,
    n34418, n34419, n34420, n34421, n34422, n34423,
    n34424, n34425, n34426, n34427, n34428, n34429,
    n34430, n34431, n34432, n34433, n34434, n34435,
    n34436, n34437, n34438, n34439, n34440, n34441,
    n34442, n34443, n34444, n34445, n34446, n34447,
    n34448, n34449, n34450, n34451, n34452, n34453,
    n34454, n34455, n34456, n34457, n34458, n34459,
    n34460, n34461, n34462, n34463, n34464, n34465,
    n34466, n34467, n34468, n34469, n34470, n34471,
    n34472, n34473, n34474, n34475, n34476, n34477,
    n34478, n34479, n34480, n34481, n34482, n34483,
    n34484, n34485, n34486, n34487, n34488, n34489,
    n34490, n34491, n34492, n34493, n34494, n34495,
    n34496, n34497, n34498, n34499, n34500, n34501,
    n34502, n34503, n34504, n34505, n34506, n34507,
    n34508, n34509, n34510, n34511, n34512, n34513,
    n34514, n34515, n34516, n34517, n34518, n34519,
    n34520, n34521, n34522, n34523, n34524, n34525,
    n34526, n34527, n34528, n34529, n34530, n34531,
    n34532, n34533, n34534, n34535, n34536, n34537,
    n34538, n34539, n34540, n34541, n34542, n34543,
    n34544, n34545, n34546, n34547, n34548, n34549,
    n34550, n34551, n34552, n34553, n34554, n34555,
    n34556, n34557, n34558, n34559, n34560, n34561,
    n34562, n34563, n34564, n34565, n34566, n34567,
    n34568, n34569, n34570, n34571, n34572, n34573,
    n34574, n34575, n34576, n34577, n34578, n34579,
    n34580, n34581, n34582, n34583, n34584, n34585,
    n34586, n34587, n34588, n34589, n34590, n34591,
    n34592, n34593, n34594, n34595, n34596, n34597,
    n34598, n34599, n34600, n34601, n34602, n34603,
    n34604, n34605, n34606, n34607, n34608, n34609,
    n34610, n34611, n34612, n34613, n34614, n34615,
    n34616, n34617, n34618, n34619, n34620, n34621,
    n34622, n34623, n34624, n34625, n34626, n34627,
    n34628, n34629, n34630, n34631, n34632, n34633,
    n34634, n34635, n34636, n34637, n34638, n34639,
    n34640, n34641, n34642, n34643, n34644, n34645,
    n34646, n34647, n34648, n34649, n34650, n34651,
    n34652, n34653, n34654, n34655, n34656, n34657,
    n34658, n34659, n34660, n34661, n34662, n34663,
    n34664, n34665, n34666, n34667, n34668, n34669,
    n34670, n34671, n34672, n34673, n34674, n34675,
    n34676, n34677, n34678, n34679, n34680, n34681,
    n34682, n34683, n34684, n34685, n34686, n34687,
    n34688, n34689, n34690, n34691, n34692, n34693,
    n34694, n34695, n34696, n34697, n34698, n34699,
    n34700, n34701, n34702, n34703, n34704, n34705,
    n34706, n34707, n34708, n34709, n34710, n34711,
    n34712, n34713, n34714, n34715, n34716, n34717,
    n34718, n34719, n34720, n34721, n34722, n34723,
    n34724, n34725, n34726, n34727, n34728, n34729,
    n34730, n34731, n34732, n34733, n34734, n34735,
    n34736, n34737, n34738, n34739, n34740, n34741,
    n34742, n34743, n34744, n34745, n34746, n34747,
    n34748, n34749, n34750, n34751, n34752, n34753,
    n34754, n34755, n34756, n34757, n34758, n34759,
    n34760, n34761, n34762, n34763, n34764, n34765,
    n34766, n34767, n34768, n34769, n34770, n34771,
    n34772, n34773, n34774, n34775, n34776, n34777,
    n34778, n34779, n34780, n34781, n34782, n34783,
    n34784, n34785, n34786, n34787, n34788, n34789,
    n34790, n34791, n34792, n34793, n34794, n34795,
    n34796, n34797, n34798, n34799, n34800, n34801,
    n34802, n34803, n34804, n34805, n34806, n34807,
    n34808, n34809, n34810, n34811, n34812, n34813,
    n34814, n34815, n34816, n34817, n34818, n34819,
    n34820, n34821, n34822, n34823, n34824, n34825,
    n34826, n34827, n34828, n34829, n34830, n34831,
    n34832, n34833, n34834, n34835, n34836, n34837,
    n34838, n34839, n34840, n34841, n34842, n34843,
    n34844, n34845, n34846, n34847, n34848, n34849,
    n34850, n34851, n34852, n34853, n34854, n34855,
    n34856, n34857, n34858, n34859, n34860, n34861,
    n34862, n34863, n34864, n34865, n34866, n34867,
    n34868, n34869, n34870, n34871, n34872, n34873,
    n34874, n34875, n34876, n34877, n34878, n34879,
    n34880, n34881, n34882, n34883, n34884, n34885,
    n34886, n34887, n34888, n34889, n34890, n34891,
    n34892, n34893, n34894, n34895, n34896, n34897,
    n34898, n34899, n34900, n34901, n34902, n34903,
    n34904, n34905, n34906, n34907, n34908, n34909,
    n34910, n34911, n34912, n34913, n34914, n34915,
    n34916, n34917, n34918, n34919, n34920, n34921,
    n34922, n34923, n34924, n34925, n34926, n34927,
    n34928, n34929, n34930, n34931, n34932, n34933,
    n34934, n34935, n34936, n34937, n34938, n34939,
    n34940, n34941, n34942, n34943, n34944, n34945,
    n34946, n34947, n34948, n34949, n34950, n34951,
    n34952, n34953, n34954, n34955, n34956, n34957,
    n34958, n34959, n34960, n34961, n34962, n34963,
    n34964, n34965, n34966, n34967, n34968, n34969,
    n34970, n34971, n34972, n34973, n34974, n34975,
    n34976, n34977, n34978, n34979, n34980, n34981,
    n34982, n34983, n34984, n34985, n34986, n34987,
    n34988, n34989, n34990, n34991, n34992, n34993,
    n34994, n34995, n34996, n34997, n34998, n34999,
    n35000, n35001, n35002, n35003, n35004, n35005,
    n35006, n35007, n35008, n35009, n35010, n35011,
    n35012, n35013, n35014, n35015, n35016, n35017,
    n35018, n35019, n35020, n35021, n35022, n35023,
    n35024, n35025, n35026, n35027, n35028, n35029,
    n35030, n35031, n35032, n35033, n35034, n35035,
    n35036, n35037, n35038, n35039, n35040, n35041,
    n35042, n35043, n35044, n35045, n35046, n35047,
    n35048, n35049, n35050, n35051, n35052, n35053,
    n35054, n35055, n35056, n35057, n35058, n35059,
    n35060, n35061, n35062, n35063, n35064, n35065,
    n35066, n35067, n35068, n35069, n35070, n35071,
    n35072, n35073, n35074, n35075, n35076, n35077,
    n35078, n35079, n35080, n35081, n35082, n35083,
    n35084, n35085, n35086, n35087, n35088, n35089,
    n35090, n35091, n35092, n35093, n35094, n35095,
    n35096, n35097, n35098, n35099, n35100, n35101,
    n35102, n35103, n35104, n35105, n35106, n35107,
    n35108, n35109, n35110, n35111, n35112, n35113,
    n35114, n35115, n35116, n35117, n35118, n35119,
    n35120, n35121, n35122, n35123, n35124, n35125,
    n35126, n35127, n35128, n35129, n35130, n35131,
    n35132, n35133, n35134, n35135, n35136, n35137,
    n35138, n35139, n35140, n35141, n35142, n35143,
    n35144, n35145, n35146, n35147, n35148, n35149,
    n35150, n35151, n35152, n35153, n35154, n35155,
    n35156, n35157, n35158, n35159, n35160, n35161,
    n35162, n35163, n35164, n35165, n35166, n35167,
    n35168, n35169, n35170, n35171, n35172, n35173,
    n35174, n35175, n35176, n35177, n35178, n35179,
    n35180, n35181, n35182, n35183, n35184, n35185,
    n35186, n35187, n35188, n35189, n35190, n35191,
    n35192, n35193, n35194, n35195, n35196, n35197,
    n35198, n35199, n35200, n35201, n35202, n35203,
    n35204, n35205, n35206, n35207, n35208, n35209,
    n35210, n35211, n35212, n35213, n35214, n35215,
    n35216, n35217, n35218, n35219, n35220, n35221,
    n35222, n35223, n35224, n35225, n35226, n35227,
    n35228, n35229, n35230, n35231, n35232, n35233,
    n35234, n35235, n35236, n35237, n35238, n35239,
    n35240, n35241, n35242, n35243, n35244, n35245,
    n35246, n35247, n35248, n35249, n35250, n35251,
    n35252, n35253, n35254, n35255, n35256, n35257,
    n35258, n35259, n35260, n35261, n35262, n35263,
    n35264, n35265, n35266, n35267, n35268, n35269,
    n35270, n35271, n35272, n35273, n35274, n35275,
    n35276, n35277, n35278, n35279, n35280, n35281,
    n35282, n35283, n35284, n35285, n35286, n35287,
    n35288, n35289, n35290, n35291, n35292, n35293,
    n35294, n35295, n35296, n35297, n35298, n35299,
    n35300, n35301, n35302, n35303, n35304, n35305,
    n35306, n35307, n35308, n35309, n35310, n35311,
    n35312, n35313, n35314, n35315, n35316, n35317,
    n35318, n35319, n35320, n35321, n35322, n35323,
    n35324, n35325, n35326, n35327, n35328, n35329,
    n35330, n35331, n35332, n35333, n35334, n35335,
    n35336, n35337, n35338, n35339, n35340, n35341,
    n35342, n35343, n35344, n35345, n35346, n35347,
    n35348, n35349, n35350, n35351, n35352, n35353,
    n35354, n35355, n35356, n35357, n35358, n35359,
    n35360, n35361, n35362, n35363, n35364, n35365,
    n35366, n35367, n35368, n35369, n35370, n35371,
    n35372, n35373, n35374, n35375, n35376, n35377,
    n35378, n35379, n35380, n35381, n35382, n35383,
    n35384, n35385, n35386, n35387, n35388, n35389,
    n35390, n35391, n35392, n35393, n35394, n35395,
    n35396, n35397, n35398, n35399, n35400, n35401,
    n35402, n35403, n35404, n35405, n35406, n35407,
    n35408, n35409, n35410, n35411, n35412, n35413,
    n35414, n35415, n35416, n35417, n35418, n35419,
    n35420, n35421, n35422, n35423, n35424, n35425,
    n35426, n35427, n35428, n35429, n35430, n35431,
    n35432, n35433, n35434, n35435, n35436, n35437,
    n35438, n35439, n35440, n35441, n35442, n35443,
    n35444, n35445, n35446, n35447, n35448, n35449,
    n35450, n35451, n35452, n35453, n35454, n35455,
    n35456, n35457, n35458, n35459, n35460, n35461,
    n35462, n35463, n35464, n35465, n35466, n35467,
    n35468, n35469, n35470, n35471, n35472, n35473,
    n35474, n35475, n35476, n35477, n35478, n35479,
    n35480, n35481, n35482, n35483, n35484, n35485,
    n35486, n35487, n35488, n35489, n35490, n35491,
    n35492, n35493, n35494, n35495, n35496, n35497,
    n35498, n35499, n35500, n35501, n35502, n35503,
    n35504, n35505, n35506, n35507, n35508, n35509,
    n35510, n35511, n35512, n35513, n35514, n35515,
    n35516, n35517, n35518, n35519, n35520, n35521,
    n35522, n35523, n35524, n35525, n35526, n35527,
    n35528, n35529, n35530, n35531, n35532, n35533,
    n35534, n35535, n35536, n35537, n35538, n35539,
    n35540, n35541, n35542, n35543, n35544, n35545,
    n35546, n35547, n35548, n35549, n35550, n35551,
    n35552, n35553, n35554, n35555, n35556, n35557,
    n35558, n35559, n35560, n35561, n35562, n35563,
    n35564, n35565, n35566, n35567, n35568, n35569,
    n35570, n35571, n35572, n35573, n35574, n35575,
    n35576, n35577, n35578, n35579, n35580, n35581,
    n35582, n35583, n35584, n35585, n35586, n35587,
    n35588, n35589, n35590, n35591, n35592, n35593,
    n35594, n35595, n35596, n35597, n35598, n35599,
    n35600, n35601, n35602, n35603, n35604, n35605,
    n35606, n35607, n35608, n35609, n35610, n35611,
    n35612, n35613, n35614, n35615, n35616, n35617,
    n35618, n35619, n35620, n35621, n35622, n35623,
    n35624, n35625, n35626, n35627, n35628, n35629,
    n35630, n35631, n35632, n35633, n35634, n35635,
    n35636, n35637, n35638, n35639, n35640, n35641,
    n35642, n35643, n35644, n35645, n35646, n35647,
    n35648, n35649, n35650, n35651, n35652, n35653,
    n35654, n35655, n35656, n35657, n35658, n35659,
    n35660, n35661, n35662, n35663, n35664, n35665,
    n35666, n35667, n35668, n35669, n35670, n35671,
    n35672, n35673, n35674, n35675, n35676, n35677,
    n35678, n35679, n35680, n35681, n35682, n35683,
    n35684, n35685, n35686, n35687, n35688, n35689,
    n35690, n35691, n35692, n35693, n35694, n35695,
    n35696, n35697, n35698, n35699, n35700, n35701,
    n35702, n35703, n35704, n35705, n35706, n35707,
    n35708, n35709, n35710, n35711, n35712, n35713,
    n35714, n35715, n35716, n35717, n35718, n35719,
    n35720, n35721, n35722, n35723, n35724, n35725,
    n35726, n35727, n35728, n35729, n35730, n35731,
    n35732, n35733, n35734, n35735, n35736, n35737,
    n35738, n35739, n35740, n35741, n35742, n35743,
    n35744, n35745, n35746, n35747, n35748, n35749,
    n35750, n35751, n35752, n35753, n35754, n35755,
    n35756, n35757, n35758, n35759, n35760, n35761,
    n35762, n35763, n35764, n35765, n35766, n35767,
    n35768, n35769, n35770, n35771, n35772, n35773,
    n35774, n35775, n35776, n35777, n35778, n35779,
    n35780, n35781, n35782, n35783, n35784, n35785,
    n35786, n35787, n35788, n35789, n35790, n35791,
    n35792, n35793, n35794, n35795, n35796, n35797,
    n35798, n35799, n35800, n35801, n35802, n35803,
    n35804, n35805, n35806, n35807, n35808, n35809,
    n35810, n35811, n35812, n35813, n35814, n35815,
    n35816, n35817, n35818, n35819, n35820, n35821,
    n35822, n35823, n35824, n35825, n35826, n35827,
    n35828, n35829, n35830, n35831, n35832, n35833,
    n35834, n35835, n35836, n35837, n35838, n35839,
    n35840, n35841, n35842, n35843, n35844, n35845,
    n35846, n35847, n35848, n35849, n35850, n35851,
    n35852, n35853, n35854, n35855, n35856, n35857,
    n35858, n35859, n35860, n35861, n35862, n35863,
    n35864, n35865, n35866, n35867, n35868, n35869,
    n35870, n35871, n35872, n35873, n35874, n35875,
    n35876, n35877, n35878, n35879, n35880, n35881,
    n35882, n35883, n35884, n35885, n35886, n35887,
    n35888, n35889, n35890, n35891, n35892, n35893,
    n35894, n35895, n35896, n35897, n35898, n35899,
    n35900, n35901, n35902, n35903, n35904, n35905,
    n35906, n35907, n35908, n35909, n35910, n35911,
    n35912, n35913, n35914, n35915, n35916, n35917,
    n35918, n35919, n35920, n35921, n35922, n35923,
    n35924, n35925, n35926, n35927, n35928, n35929,
    n35930, n35931, n35932, n35933, n35934, n35935,
    n35936, n35937, n35938, n35939, n35940, n35941,
    n35942, n35943, n35944, n35945, n35946, n35947,
    n35948, n35949, n35950, n35951, n35952, n35953,
    n35954, n35955, n35956, n35957, n35958, n35959,
    n35960, n35961, n35962, n35963, n35964, n35965,
    n35966, n35967, n35968, n35969, n35970, n35971,
    n35972, n35973, n35974, n35975, n35976, n35977,
    n35978, n35979, n35980, n35981, n35982, n35983,
    n35984, n35985, n35986, n35987, n35988, n35989,
    n35990, n35991, n35992, n35993, n35994, n35995,
    n35996, n35997, n35998, n35999, n36000, n36001,
    n36002, n36003, n36004, n36005, n36006, n36007,
    n36008, n36009, n36010, n36011, n36012, n36013,
    n36014, n36015, n36016, n36017, n36018, n36019,
    n36020, n36021, n36022, n36023, n36024, n36025,
    n36026, n36027, n36028, n36029, n36030, n36031,
    n36032, n36033, n36034, n36035, n36036, n36037,
    n36038, n36039, n36040, n36041, n36042, n36043,
    n36044, n36045, n36046, n36047, n36048, n36049,
    n36050, n36051, n36052, n36053, n36054, n36055,
    n36056, n36057, n36058, n36059, n36060, n36061,
    n36062, n36063, n36064, n36065, n36066, n36067,
    n36068, n36069, n36070, n36071, n36072, n36073,
    n36074, n36075, n36076, n36077, n36078, n36079,
    n36080, n36081, n36082, n36083, n36084, n36085,
    n36086, n36087, n36088, n36089, n36090, n36091,
    n36092, n36093, n36094, n36095, n36096, n36097,
    n36098, n36099, n36100, n36101, n36102, n36103,
    n36104, n36105, n36106, n36107, n36108, n36109,
    n36110, n36111, n36112, n36113, n36114, n36115,
    n36116, n36117, n36118, n36119, n36120, n36121,
    n36122, n36123, n36124, n36125, n36126, n36127,
    n36128, n36129, n36130, n36131, n36132, n36133,
    n36134, n36135, n36136, n36137, n36138, n36139,
    n36140, n36141, n36142, n36143, n36144, n36145,
    n36146, n36147, n36148, n36149, n36150, n36151,
    n36152, n36153, n36154, n36155, n36156, n36157,
    n36158, n36159, n36160, n36161, n36162, n36163,
    n36164, n36165, n36166, n36167, n36168, n36169,
    n36170, n36171, n36172, n36173, n36174, n36175,
    n36176, n36177, n36178, n36179, n36180, n36181,
    n36182, n36183, n36184, n36185, n36186, n36187,
    n36188, n36189, n36190, n36191, n36192, n36193,
    n36194, n36195, n36196, n36197, n36198, n36199,
    n36200, n36201, n36202, n36203, n36204, n36205,
    n36206, n36207, n36208, n36209, n36210, n36211,
    n36212, n36213, n36214, n36215, n36216, n36217,
    n36218, n36219, n36220, n36221, n36222, n36223,
    n36224, n36225, n36226, n36227, n36228, n36229,
    n36230, n36231, n36232, n36233, n36234, n36235,
    n36236, n36237, n36238, n36239, n36240, n36241,
    n36242, n36243, n36244, n36245, n36246, n36247,
    n36248, n36249, n36250, n36251, n36252, n36253,
    n36254, n36255, n36256, n36257, n36258, n36259,
    n36260, n36261, n36262, n36263, n36264, n36265,
    n36266, n36267, n36268, n36269, n36270, n36271,
    n36272, n36273, n36274, n36275, n36276, n36277,
    n36278, n36279, n36280, n36281, n36282, n36283,
    n36284, n36285, n36286, n36287, n36288, n36289,
    n36290, n36291, n36292, n36293, n36294, n36295,
    n36296, n36297, n36298, n36299, n36300, n36301,
    n36302, n36303, n36304, n36305, n36306, n36307,
    n36308, n36309, n36310, n36311, n36312, n36313,
    n36314, n36315, n36316, n36317, n36318, n36319,
    n36320, n36321, n36322, n36323, n36324, n36325,
    n36326, n36327, n36328, n36329, n36330, n36331,
    n36332, n36333, n36334, n36335, n36336, n36337,
    n36338, n36339, n36340, n36341, n36342, n36343,
    n36344, n36345, n36346, n36347, n36348, n36349,
    n36350, n36351, n36352, n36353, n36354, n36355,
    n36356, n36357, n36358, n36359, n36360, n36361,
    n36362, n36363, n36364, n36365, n36366, n36367,
    n36368, n36369, n36370, n36371, n36372, n36373,
    n36374, n36375, n36376, n36377, n36378, n36379,
    n36380, n36381, n36382, n36383, n36384, n36385,
    n36386, n36387, n36388, n36389, n36390, n36391,
    n36392, n36393, n36394, n36395, n36396, n36397,
    n36398, n36399, n36400, n36401, n36402, n36403,
    n36404, n36405, n36406, n36407, n36408, n36409,
    n36410, n36411, n36412, n36413, n36414, n36415,
    n36416, n36417, n36418, n36419, n36420, n36421,
    n36422, n36423, n36424, n36425, n36426, n36427,
    n36428, n36429, n36430, n36431, n36432, n36433,
    n36434, n36435, n36436, n36437, n36438, n36439,
    n36440, n36441, n36442, n36443, n36444, n36445,
    n36446, n36447, n36448, n36449, n36450, n36451,
    n36452, n36453, n36454, n36455, n36456, n36457,
    n36458, n36459, n36460, n36461, n36462, n36463,
    n36464, n36465, n36466, n36467, n36468, n36469,
    n36470, n36471, n36472, n36473, n36474, n36475,
    n36476, n36477, n36478, n36479, n36480, n36481,
    n36482, n36483, n36484, n36485, n36486, n36487,
    n36488, n36489, n36490, n36491, n36492, n36493,
    n36494, n36495, n36496, n36497, n36498, n36499,
    n36500, n36501, n36502, n36503, n36504, n36505,
    n36506, n36507, n36508, n36509, n36510, n36511;
  assign n193 = ~pi126  & ~pi127 ;
  assign n194 = ~pi62  & ~pi63 ;
  assign n195 = pi126  & pi127 ;
  assign n196 = ~pi124  & ~pi125 ;
  assign n197 = ~pi126  & ~n196;
  assign n198 = ~n195 & ~n197;
  assign n199 = ~pi124  & ~n198;
  assign n200 = pi125  & ~n199;
  assign n201 = n196 & ~n198;
  assign n202 = n195 & n196;
  assign n203 = ~n200 & ~n32240;
  assign n204 = pi124  & ~n198;
  assign n205 = ~pi122  & ~pi123 ;
  assign n206 = ~pi124  & n205;
  assign n207 = ~n204 & ~n206;
  assign n208 = n203 & ~n207;
  assign n209 = n193 & ~n208;
  assign n210 = ~n203 & n207;
  assign n211 = pi126  & n196;
  assign n212 = pi127  & ~n197;
  assign n213 = pi127  & ~n211;
  assign n214 = ~n197 & n213;
  assign n215 = ~n211 & n212;
  assign n216 = ~n210 & ~n32241;
  assign n217 = ~n209 & n216;
  assign n218 = pi122  & ~n217;
  assign n219 = ~pi120  & ~pi121 ;
  assign n220 = ~pi122  & n219;
  assign n221 = ~n195 & ~n220;
  assign n222 = ~n197 & n221;
  assign n223 = ~pi122  & ~n219;
  assign n224 = pi122  & n217;
  assign n225 = ~n223 & ~n224;
  assign n226 = ~n218 & ~n220;
  assign n227 = n198 & ~n32242;
  assign n228 = ~n218 & n222;
  assign n229 = ~n198 & n32242;
  assign n230 = ~pi122  & ~n217;
  assign n231 = ~pi123  & n230;
  assign n232 = n205 & ~n217;
  assign n233 = pi123  & ~n230;
  assign n234 = ~n32244 & ~n233;
  assign n235 = ~n229 & ~n234;
  assign n236 = ~n32243 & n234;
  assign n237 = ~n229 & ~n236;
  assign n238 = ~n32243 & ~n235;
  assign n239 = ~n198 & ~n32241;
  assign n240 = ~n210 & n239;
  assign n241 = ~n198 & n217;
  assign n242 = ~n209 & n240;
  assign n243 = ~n32244 & ~n32246;
  assign n244 = pi124  & ~n243;
  assign n245 = ~pi124  & ~n32246;
  assign n246 = ~pi124  & n243;
  assign n247 = ~n32244 & n245;
  assign n248 = ~n244 & ~n32247;
  assign n249 = n203 & ~n32241;
  assign n250 = ~n208 & ~n210;
  assign n251 = n208 & ~n217;
  assign n252 = n208 & n32241;
  assign n253 = ~n210 & ~n32248;
  assign n254 = ~n249 & ~n250;
  assign n255 = ~n248 & n32249;
  assign n256 = ~n32245 & ~n248;
  assign n257 = n32249 & n256;
  assign n258 = ~n32245 & n255;
  assign n259 = n193 & ~n32250;
  assign n260 = n32245 & n248;
  assign n261 = ~n193 & ~n249;
  assign n262 = ~n193 & ~n208;
  assign n263 = ~n210 & n262;
  assign n264 = n207 & ~n32241;
  assign n265 = n263 & ~n264;
  assign n266 = n203 & ~n217;
  assign n267 = n207 & ~n266;
  assign n268 = n262 & ~n267;
  assign n269 = n250 & n261;
  assign n270 = ~n260 & ~n32251;
  assign n271 = ~n259 & n270;
  assign n272 = pi120  & ~n271;
  assign n273 = ~pi118  & ~pi119 ;
  assign n274 = ~pi120  & n273;
  assign n275 = ~n272 & ~n274;
  assign n276 = ~n217 & ~n275;
  assign n277 = ~pi120  & ~n271;
  assign n278 = pi121  & ~n277;
  assign n279 = ~pi121  & n277;
  assign n280 = n219 & ~n271;
  assign n281 = ~n278 & ~n32252;
  assign n282 = ~n32241 & ~n274;
  assign n283 = ~n210 & n282;
  assign n284 = ~n209 & n283;
  assign n285 = n217 & n275;
  assign n286 = ~n272 & n284;
  assign n287 = n281 & ~n32253;
  assign n288 = ~n276 & ~n287;
  assign n289 = ~n198 & ~n288;
  assign n290 = n198 & ~n276;
  assign n291 = ~n287 & n290;
  assign n292 = ~n217 & ~n263;
  assign n293 = ~n217 & ~n32251;
  assign n294 = ~n209 & n32249;
  assign n295 = ~n260 & n32254;
  assign n296 = ~n259 & n295;
  assign n297 = ~n32252 & ~n296;
  assign n298 = pi122  & ~n297;
  assign n299 = ~pi122  & ~n296;
  assign n300 = ~pi122  & n297;
  assign n301 = ~n32252 & n299;
  assign n302 = ~n298 & ~n32255;
  assign n303 = ~n291 & ~n302;
  assign n304 = ~n289 & ~n303;
  assign n305 = ~n32243 & ~n229;
  assign n306 = ~n271 & n305;
  assign n307 = n234 & ~n306;
  assign n308 = ~n234 & n305;
  assign n309 = ~n234 & n306;
  assign n310 = ~n271 & n308;
  assign n311 = ~n307 & ~n32256;
  assign n312 = n256 & ~n271;
  assign n313 = ~n260 & ~n312;
  assign n314 = ~n311 & n313;
  assign n315 = ~n304 & n314;
  assign n316 = n193 & ~n315;
  assign n317 = ~n289 & n311;
  assign n318 = ~n303 & n317;
  assign n319 = n304 & n311;
  assign n320 = ~n248 & n271;
  assign n321 = ~n193 & ~n256;
  assign n322 = ~n260 & n321;
  assign n323 = ~n271 & ~n322;
  assign n324 = n32245 & ~n271;
  assign n325 = ~n248 & ~n324;
  assign n326 = ~n193 & ~n260;
  assign n327 = ~n325 & n326;
  assign n328 = ~n320 & ~n323;
  assign n329 = ~n32257 & ~n32258;
  assign n330 = ~n316 & n329;
  assign n331 = pi118  & ~n330;
  assign n332 = ~pi116  & ~pi117 ;
  assign n333 = ~pi118  & n332;
  assign n334 = ~n331 & ~n333;
  assign n335 = ~n271 & ~n334;
  assign n336 = ~n203 & ~n32241;
  assign n337 = ~n210 & n336;
  assign n338 = ~n203 & n217;
  assign n339 = ~n209 & n337;
  assign n340 = ~n333 & ~n32259;
  assign n341 = ~n32251 & n340;
  assign n342 = ~n260 & n341;
  assign n343 = ~n259 & n342;
  assign n344 = n271 & n334;
  assign n345 = ~n331 & n343;
  assign n346 = ~pi118  & ~n330;
  assign n347 = pi119  & ~n346;
  assign n348 = ~pi119  & n346;
  assign n349 = n273 & ~n330;
  assign n350 = ~n347 & ~n32261;
  assign n351 = ~n32260 & n350;
  assign n352 = ~n335 & ~n351;
  assign n353 = ~n217 & ~n352;
  assign n354 = ~n32257 & n323;
  assign n355 = ~n316 & n354;
  assign n356 = ~n32261 & ~n355;
  assign n357 = pi120  & ~n356;
  assign n358 = ~pi120  & ~n355;
  assign n359 = ~pi120  & n356;
  assign n360 = ~n32261 & n358;
  assign n361 = ~n357 & ~n32262;
  assign n362 = n217 & ~n335;
  assign n363 = n217 & n352;
  assign n364 = ~n351 & n362;
  assign n365 = ~n361 & ~n32263;
  assign n366 = ~n353 & ~n365;
  assign n367 = ~n198 & ~n366;
  assign n368 = n198 & ~n353;
  assign n369 = ~n365 & n368;
  assign n370 = ~n276 & ~n32253;
  assign n371 = ~n330 & n370;
  assign n372 = n281 & ~n371;
  assign n373 = ~n281 & ~n32253;
  assign n374 = ~n276 & n373;
  assign n375 = ~n281 & n370;
  assign n376 = ~n281 & n371;
  assign n377 = ~n330 & n32264;
  assign n378 = ~n372 & ~n32265;
  assign n379 = ~n369 & ~n378;
  assign n380 = ~n367 & ~n379;
  assign n381 = ~n289 & ~n291;
  assign n382 = ~n330 & n381;
  assign n383 = ~n302 & ~n382;
  assign n384 = ~n291 & n302;
  assign n385 = ~n289 & n384;
  assign n386 = n302 & n382;
  assign n387 = ~n330 & n385;
  assign n388 = ~n383 & ~n32266;
  assign n389 = ~n304 & ~n311;
  assign n390 = ~n330 & n389;
  assign n391 = ~n32257 & ~n390;
  assign n392 = ~n388 & n391;
  assign n393 = ~n380 & n392;
  assign n394 = n193 & ~n393;
  assign n395 = ~n367 & n388;
  assign n396 = n380 & n388;
  assign n397 = ~n379 & n395;
  assign n398 = n304 & ~n330;
  assign n399 = ~n311 & ~n398;
  assign n400 = ~n193 & ~n32257;
  assign n401 = ~n399 & n400;
  assign n402 = ~n32267 & ~n401;
  assign n403 = ~n394 & n402;
  assign n404 = pi116  & ~n403;
  assign n405 = ~pi114  & ~pi115 ;
  assign n406 = ~pi116  & n405;
  assign n407 = ~n404 & ~n406;
  assign n408 = ~n330 & ~n407;
  assign n409 = ~pi116  & ~n403;
  assign n410 = pi117  & ~n409;
  assign n411 = ~pi117  & n409;
  assign n412 = n332 & ~n403;
  assign n413 = ~n410 & ~n32268;
  assign n414 = ~n32247 & ~n32259;
  assign n415 = ~n244 & n414;
  assign n416 = ~n32251 & n415;
  assign n417 = ~n260 & n416;
  assign n418 = ~n259 & n417;
  assign n419 = ~n406 & ~n418;
  assign n420 = ~n32258 & n419;
  assign n421 = ~n32257 & n420;
  assign n422 = ~n316 & n421;
  assign n423 = n330 & n407;
  assign n424 = ~n404 & n422;
  assign n425 = n413 & ~n32269;
  assign n426 = ~n408 & ~n425;
  assign n427 = ~n271 & ~n426;
  assign n428 = n271 & ~n408;
  assign n429 = ~n425 & n428;
  assign n430 = ~n330 & ~n401;
  assign n431 = ~n32267 & n430;
  assign n432 = ~n394 & n431;
  assign n433 = ~n32268 & ~n432;
  assign n434 = pi118  & ~n433;
  assign n435 = ~pi118  & ~n432;
  assign n436 = ~pi118  & n433;
  assign n437 = ~n32268 & n435;
  assign n438 = ~n434 & ~n32270;
  assign n439 = ~n429 & ~n438;
  assign n440 = ~n427 & ~n439;
  assign n441 = ~n217 & ~n440;
  assign n442 = n217 & ~n427;
  assign n443 = ~n439 & n442;
  assign n444 = n217 & n440;
  assign n445 = ~n335 & ~n32260;
  assign n446 = ~n403 & n445;
  assign n447 = n350 & ~n446;
  assign n448 = ~n350 & n445;
  assign n449 = ~n350 & n446;
  assign n450 = ~n403 & n448;
  assign n451 = ~n447 & ~n32272;
  assign n452 = ~n32271 & ~n451;
  assign n453 = ~n441 & ~n452;
  assign n454 = ~n198 & ~n453;
  assign n455 = n198 & ~n441;
  assign n456 = ~n452 & n455;
  assign n457 = ~n353 & ~n32263;
  assign n458 = ~n353 & ~n403;
  assign n459 = ~n32263 & n458;
  assign n460 = ~n403 & n457;
  assign n461 = n361 & ~n32273;
  assign n462 = n365 & n458;
  assign n463 = n361 & ~n32263;
  assign n464 = ~n353 & n463;
  assign n465 = ~n403 & n464;
  assign n466 = ~n361 & ~n32273;
  assign n467 = ~n465 & ~n466;
  assign n468 = ~n461 & ~n462;
  assign n469 = ~n456 & ~n32274;
  assign n470 = ~n454 & ~n469;
  assign n471 = ~n367 & ~n369;
  assign n472 = ~n403 & n471;
  assign n473 = n378 & ~n472;
  assign n474 = ~n378 & n472;
  assign n475 = ~n367 & n378;
  assign n476 = ~n369 & n475;
  assign n477 = n378 & n472;
  assign n478 = ~n403 & n476;
  assign n479 = ~n378 & ~n472;
  assign n480 = ~n32275 & ~n479;
  assign n481 = ~n473 & ~n474;
  assign n482 = ~n380 & ~n388;
  assign n483 = ~n388 & ~n403;
  assign n484 = ~n380 & n483;
  assign n485 = ~n403 & n482;
  assign n486 = ~n32267 & ~n32277;
  assign n487 = ~n32276 & n486;
  assign n488 = ~n470 & n487;
  assign n489 = n193 & ~n488;
  assign n490 = ~n454 & n32276;
  assign n491 = ~n469 & n490;
  assign n492 = n470 & n32276;
  assign n493 = n380 & ~n483;
  assign n494 = ~n193 & ~n482;
  assign n495 = ~n493 & n494;
  assign n496 = ~n32278 & ~n495;
  assign n497 = ~n489 & n496;
  assign n498 = pi114  & ~n497;
  assign n499 = ~pi112  & ~pi113 ;
  assign n500 = ~pi114  & n499;
  assign n501 = ~n498 & ~n500;
  assign n502 = ~n403 & ~n501;
  assign n503 = ~n32256 & ~n418;
  assign n504 = ~n307 & n503;
  assign n505 = ~n32258 & n504;
  assign n506 = ~n32257 & n505;
  assign n507 = n311 & n330;
  assign n508 = ~n316 & n506;
  assign n509 = ~n500 & ~n32279;
  assign n510 = ~n401 & n509;
  assign n511 = ~n32267 & n510;
  assign n512 = ~n394 & n511;
  assign n513 = n403 & n501;
  assign n514 = ~n498 & n512;
  assign n515 = ~pi114  & ~n497;
  assign n516 = pi115  & ~n515;
  assign n517 = ~pi115  & n515;
  assign n518 = n405 & ~n497;
  assign n519 = ~n516 & ~n32281;
  assign n520 = ~n32280 & n519;
  assign n521 = ~n502 & ~n520;
  assign n522 = ~n330 & ~n521;
  assign n523 = ~n403 & ~n495;
  assign n524 = ~n32278 & n523;
  assign n525 = ~n489 & n524;
  assign n526 = ~n32281 & ~n525;
  assign n527 = pi116  & ~n526;
  assign n528 = ~pi116  & ~n525;
  assign n529 = ~pi116  & n526;
  assign n530 = ~n32281 & n528;
  assign n531 = ~n527 & ~n32282;
  assign n532 = n330 & ~n502;
  assign n533 = n330 & n521;
  assign n534 = ~n520 & n532;
  assign n535 = ~n531 & ~n32283;
  assign n536 = ~n522 & ~n535;
  assign n537 = ~n271 & ~n536;
  assign n538 = n271 & ~n522;
  assign n539 = ~n535 & n538;
  assign n540 = ~n408 & ~n32269;
  assign n541 = ~n497 & n540;
  assign n542 = n413 & ~n541;
  assign n543 = ~n413 & n540;
  assign n544 = ~n413 & n541;
  assign n545 = ~n497 & n543;
  assign n546 = ~n542 & ~n32284;
  assign n547 = ~n539 & ~n546;
  assign n548 = ~n537 & ~n547;
  assign n549 = ~n217 & ~n548;
  assign n550 = ~n427 & ~n429;
  assign n551 = ~n497 & n550;
  assign n552 = ~n438 & ~n551;
  assign n553 = ~n429 & n438;
  assign n554 = ~n427 & n553;
  assign n555 = n438 & n551;
  assign n556 = ~n497 & n554;
  assign n557 = ~n552 & ~n32285;
  assign n558 = n217 & ~n537;
  assign n559 = n217 & n548;
  assign n560 = ~n547 & n558;
  assign n561 = ~n557 & ~n32286;
  assign n562 = ~n549 & ~n561;
  assign n563 = ~n198 & ~n562;
  assign n564 = n198 & ~n549;
  assign n565 = ~n561 & n564;
  assign n566 = ~n441 & ~n32271;
  assign n567 = ~n497 & n566;
  assign n568 = n451 & ~n567;
  assign n569 = ~n451 & n567;
  assign n570 = ~n441 & n451;
  assign n571 = ~n32271 & n570;
  assign n572 = n451 & n567;
  assign n573 = ~n497 & n571;
  assign n574 = ~n451 & ~n567;
  assign n575 = ~n32287 & ~n574;
  assign n576 = ~n568 & ~n569;
  assign n577 = ~n565 & ~n32288;
  assign n578 = ~n563 & ~n577;
  assign n579 = ~n454 & ~n456;
  assign n580 = ~n497 & n579;
  assign n581 = ~n32274 & ~n580;
  assign n582 = ~n456 & n32274;
  assign n583 = ~n454 & n582;
  assign n584 = n32274 & n580;
  assign n585 = ~n497 & n583;
  assign n586 = ~n581 & ~n32289;
  assign n587 = ~n470 & ~n32276;
  assign n588 = ~n32276 & ~n497;
  assign n589 = ~n470 & n588;
  assign n590 = ~n497 & n587;
  assign n591 = ~n32278 & ~n32290;
  assign n592 = ~n586 & n591;
  assign n593 = ~n578 & n592;
  assign n594 = n193 & ~n593;
  assign n595 = ~n563 & n586;
  assign n596 = n578 & n586;
  assign n597 = ~n577 & n595;
  assign n598 = n470 & ~n588;
  assign n599 = ~n193 & ~n587;
  assign n600 = ~n598 & n599;
  assign n601 = ~n32291 & ~n600;
  assign n602 = ~n594 & n601;
  assign n603 = pi112  & ~n602;
  assign n604 = ~pi110  & ~pi111 ;
  assign n605 = ~pi112  & n604;
  assign n606 = ~n603 & ~n605;
  assign n607 = ~n497 & ~n606;
  assign n608 = ~pi112  & ~n602;
  assign n609 = pi113  & ~n608;
  assign n610 = ~pi113  & n608;
  assign n611 = n499 & ~n602;
  assign n612 = ~n609 & ~n32292;
  assign n613 = ~n32266 & ~n32279;
  assign n614 = ~n383 & n613;
  assign n615 = ~n401 & n614;
  assign n616 = ~n32267 & n615;
  assign n617 = n388 & n403;
  assign n618 = ~n394 & n616;
  assign n619 = ~n605 & ~n32293;
  assign n620 = ~n495 & n619;
  assign n621 = ~n32278 & n620;
  assign n622 = ~n489 & n621;
  assign n623 = n497 & n606;
  assign n624 = ~n603 & n622;
  assign n625 = n612 & ~n32294;
  assign n626 = ~n607 & ~n625;
  assign n627 = ~n403 & ~n626;
  assign n628 = n403 & ~n607;
  assign n629 = ~n625 & n628;
  assign n630 = ~n497 & ~n600;
  assign n631 = ~n32291 & n630;
  assign n632 = ~n594 & n631;
  assign n633 = ~n32292 & ~n632;
  assign n634 = pi114  & ~n633;
  assign n635 = ~pi114  & ~n632;
  assign n636 = ~pi114  & n633;
  assign n637 = ~n32292 & n635;
  assign n638 = ~n634 & ~n32295;
  assign n639 = ~n629 & ~n638;
  assign n640 = ~n627 & ~n639;
  assign n641 = ~n330 & ~n640;
  assign n642 = n330 & ~n627;
  assign n643 = ~n639 & n642;
  assign n644 = n330 & n640;
  assign n645 = ~n502 & ~n32280;
  assign n646 = ~n602 & n645;
  assign n647 = n519 & ~n646;
  assign n648 = ~n519 & n645;
  assign n649 = ~n519 & n646;
  assign n650 = ~n602 & n648;
  assign n651 = ~n647 & ~n32297;
  assign n652 = ~n32296 & ~n651;
  assign n653 = ~n641 & ~n652;
  assign n654 = ~n271 & ~n653;
  assign n655 = n271 & ~n641;
  assign n656 = ~n652 & n655;
  assign n657 = ~n522 & ~n32283;
  assign n658 = ~n522 & ~n602;
  assign n659 = ~n32283 & n658;
  assign n660 = ~n602 & n657;
  assign n661 = n531 & ~n32298;
  assign n662 = n535 & n658;
  assign n663 = n531 & ~n32283;
  assign n664 = ~n522 & n663;
  assign n665 = ~n602 & n664;
  assign n666 = ~n531 & ~n32298;
  assign n667 = ~n665 & ~n666;
  assign n668 = ~n661 & ~n662;
  assign n669 = ~n656 & ~n32299;
  assign n670 = ~n654 & ~n669;
  assign n671 = ~n217 & ~n670;
  assign n672 = n217 & ~n654;
  assign n673 = ~n669 & n672;
  assign n674 = n217 & n670;
  assign n675 = ~n537 & ~n539;
  assign n676 = ~n602 & n675;
  assign n677 = n546 & ~n676;
  assign n678 = ~n546 & n676;
  assign n679 = ~n537 & n546;
  assign n680 = ~n539 & n679;
  assign n681 = n546 & n676;
  assign n682 = ~n602 & n680;
  assign n683 = ~n546 & ~n676;
  assign n684 = ~n32301 & ~n683;
  assign n685 = ~n677 & ~n678;
  assign n686 = ~n32300 & ~n32302;
  assign n687 = ~n671 & ~n686;
  assign n688 = ~n198 & ~n687;
  assign n689 = n198 & ~n671;
  assign n690 = ~n686 & n689;
  assign n691 = ~n549 & ~n32286;
  assign n692 = ~n549 & ~n602;
  assign n693 = ~n32286 & n692;
  assign n694 = ~n602 & n691;
  assign n695 = n557 & ~n32303;
  assign n696 = n561 & n692;
  assign n697 = n557 & ~n32286;
  assign n698 = ~n549 & n697;
  assign n699 = ~n602 & n698;
  assign n700 = ~n557 & ~n32303;
  assign n701 = ~n699 & ~n700;
  assign n702 = ~n695 & ~n696;
  assign n703 = ~n690 & ~n32304;
  assign n704 = ~n688 & ~n703;
  assign n705 = ~n563 & ~n565;
  assign n706 = ~n602 & n705;
  assign n707 = ~n32288 & n706;
  assign n708 = n32288 & ~n706;
  assign n709 = ~n563 & n32288;
  assign n710 = ~n565 & n709;
  assign n711 = ~n602 & n710;
  assign n712 = ~n32288 & ~n706;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~n707 & ~n708;
  assign n715 = ~n578 & ~n586;
  assign n716 = ~n586 & ~n602;
  assign n717 = ~n578 & n716;
  assign n718 = ~n602 & n715;
  assign n719 = ~n32291 & ~n32306;
  assign n720 = ~n32305 & n719;
  assign n721 = ~n704 & n720;
  assign n722 = n193 & ~n721;
  assign n723 = ~n688 & n32305;
  assign n724 = ~n703 & n723;
  assign n725 = n704 & n32305;
  assign n726 = n578 & ~n716;
  assign n727 = ~n193 & ~n715;
  assign n728 = ~n726 & n727;
  assign n729 = ~n32307 & ~n728;
  assign n730 = ~n722 & n729;
  assign n731 = pi110  & ~n730;
  assign n732 = ~pi108  & ~pi109 ;
  assign n733 = ~pi110  & n732;
  assign n734 = ~n731 & ~n733;
  assign n735 = ~n602 & ~n734;
  assign n736 = ~n32275 & ~n32293;
  assign n737 = ~n479 & n736;
  assign n738 = ~n495 & n737;
  assign n739 = ~n32278 & n738;
  assign n740 = n32276 & n497;
  assign n741 = ~n489 & n739;
  assign n742 = ~n733 & ~n32308;
  assign n743 = ~n600 & n742;
  assign n744 = ~n32291 & n743;
  assign n745 = ~n594 & n744;
  assign n746 = n602 & n734;
  assign n747 = ~n731 & n745;
  assign n748 = ~pi110  & ~n730;
  assign n749 = pi111  & ~n748;
  assign n750 = ~pi111  & n748;
  assign n751 = n604 & ~n730;
  assign n752 = ~n749 & ~n32310;
  assign n753 = ~n32309 & n752;
  assign n754 = ~n735 & ~n753;
  assign n755 = ~n497 & ~n754;
  assign n756 = ~n602 & ~n728;
  assign n757 = ~n32307 & n756;
  assign n758 = ~n722 & n757;
  assign n759 = ~n32310 & ~n758;
  assign n760 = pi112  & ~n759;
  assign n761 = ~pi112  & ~n758;
  assign n762 = ~pi112  & n759;
  assign n763 = ~n32310 & n761;
  assign n764 = ~n760 & ~n32311;
  assign n765 = n497 & ~n735;
  assign n766 = n497 & n754;
  assign n767 = ~n753 & n765;
  assign n768 = ~n764 & ~n32312;
  assign n769 = ~n755 & ~n768;
  assign n770 = ~n403 & ~n769;
  assign n771 = n403 & ~n755;
  assign n772 = ~n768 & n771;
  assign n773 = ~n607 & ~n32294;
  assign n774 = ~n730 & n773;
  assign n775 = n612 & ~n774;
  assign n776 = ~n612 & ~n32294;
  assign n777 = ~n607 & n776;
  assign n778 = ~n612 & n773;
  assign n779 = ~n612 & n774;
  assign n780 = ~n730 & n32313;
  assign n781 = ~n775 & ~n32314;
  assign n782 = ~n772 & ~n781;
  assign n783 = ~n770 & ~n782;
  assign n784 = ~n330 & ~n783;
  assign n785 = ~n627 & ~n629;
  assign n786 = ~n730 & n785;
  assign n787 = ~n638 & ~n786;
  assign n788 = ~n629 & n638;
  assign n789 = ~n627 & n788;
  assign n790 = n638 & n786;
  assign n791 = ~n730 & n789;
  assign n792 = ~n787 & ~n32315;
  assign n793 = n330 & ~n770;
  assign n794 = n330 & n783;
  assign n795 = ~n782 & n793;
  assign n796 = ~n792 & ~n32316;
  assign n797 = ~n784 & ~n796;
  assign n798 = ~n271 & ~n797;
  assign n799 = n271 & ~n784;
  assign n800 = ~n796 & n799;
  assign n801 = ~n641 & ~n32296;
  assign n802 = ~n730 & n801;
  assign n803 = n651 & ~n802;
  assign n804 = ~n651 & n802;
  assign n805 = ~n641 & n651;
  assign n806 = ~n32296 & n805;
  assign n807 = n651 & n802;
  assign n808 = ~n730 & n806;
  assign n809 = ~n651 & ~n802;
  assign n810 = ~n32317 & ~n809;
  assign n811 = ~n803 & ~n804;
  assign n812 = ~n800 & ~n32318;
  assign n813 = ~n798 & ~n812;
  assign n814 = ~n217 & ~n813;
  assign n815 = ~n654 & ~n656;
  assign n816 = ~n730 & n815;
  assign n817 = ~n32299 & ~n816;
  assign n818 = ~n656 & n32299;
  assign n819 = ~n654 & n818;
  assign n820 = n32299 & n816;
  assign n821 = ~n730 & n819;
  assign n822 = ~n817 & ~n32319;
  assign n823 = n217 & ~n798;
  assign n824 = n217 & n813;
  assign n825 = ~n812 & n823;
  assign n826 = ~n822 & ~n32320;
  assign n827 = ~n814 & ~n826;
  assign n828 = ~n198 & ~n827;
  assign n829 = n198 & ~n814;
  assign n830 = ~n826 & n829;
  assign n831 = ~n671 & ~n32300;
  assign n832 = ~n730 & n831;
  assign n833 = ~n32302 & n832;
  assign n834 = n32302 & ~n832;
  assign n835 = ~n671 & n32302;
  assign n836 = ~n32300 & n835;
  assign n837 = ~n730 & n836;
  assign n838 = ~n32302 & ~n832;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~n833 & ~n834;
  assign n841 = ~n830 & ~n32321;
  assign n842 = ~n828 & ~n841;
  assign n843 = ~n688 & ~n690;
  assign n844 = ~n730 & n843;
  assign n845 = ~n32304 & ~n844;
  assign n846 = ~n690 & n32304;
  assign n847 = ~n688 & n846;
  assign n848 = n32304 & n844;
  assign n849 = ~n730 & n847;
  assign n850 = ~n845 & ~n32322;
  assign n851 = ~n704 & ~n32305;
  assign n852 = ~n32305 & ~n730;
  assign n853 = ~n704 & n852;
  assign n854 = ~n730 & n851;
  assign n855 = ~n32307 & ~n32323;
  assign n856 = ~n850 & n855;
  assign n857 = ~n842 & n856;
  assign n858 = n193 & ~n857;
  assign n859 = ~n828 & n850;
  assign n860 = n842 & n850;
  assign n861 = ~n841 & n859;
  assign n862 = n704 & ~n852;
  assign n863 = ~n193 & ~n851;
  assign n864 = ~n862 & n863;
  assign n865 = ~n32324 & ~n864;
  assign n866 = ~n858 & n865;
  assign n867 = pi108  & ~n866;
  assign n868 = ~pi106  & ~pi107 ;
  assign n869 = ~pi108  & n868;
  assign n870 = ~n867 & ~n869;
  assign n871 = ~n730 & ~n870;
  assign n872 = ~pi108  & ~n866;
  assign n873 = pi109  & ~n872;
  assign n874 = ~pi109  & n872;
  assign n875 = n732 & ~n866;
  assign n876 = ~n873 & ~n32325;
  assign n877 = ~n32289 & ~n32308;
  assign n878 = ~n581 & n877;
  assign n879 = ~n600 & n878;
  assign n880 = ~n32291 & n879;
  assign n881 = n586 & n602;
  assign n882 = ~n594 & n880;
  assign n883 = ~n869 & ~n32326;
  assign n884 = ~n728 & n883;
  assign n885 = ~n32307 & n884;
  assign n886 = ~n722 & n885;
  assign n887 = n730 & n870;
  assign n888 = ~n867 & n886;
  assign n889 = n876 & ~n32327;
  assign n890 = ~n871 & ~n889;
  assign n891 = ~n602 & ~n890;
  assign n892 = n602 & ~n871;
  assign n893 = ~n889 & n892;
  assign n894 = ~n730 & ~n864;
  assign n895 = ~n32324 & n894;
  assign n896 = ~n858 & n895;
  assign n897 = ~n32325 & ~n896;
  assign n898 = pi110  & ~n897;
  assign n899 = ~pi110  & ~n896;
  assign n900 = ~pi110  & n897;
  assign n901 = ~n32325 & n899;
  assign n902 = ~n898 & ~n32328;
  assign n903 = ~n893 & ~n902;
  assign n904 = ~n891 & ~n903;
  assign n905 = ~n497 & ~n904;
  assign n906 = n497 & ~n891;
  assign n907 = ~n903 & n906;
  assign n908 = n497 & n904;
  assign n909 = ~n735 & ~n32309;
  assign n910 = ~n866 & n909;
  assign n911 = n752 & ~n910;
  assign n912 = ~n752 & n909;
  assign n913 = ~n752 & n910;
  assign n914 = ~n866 & n912;
  assign n915 = ~n911 & ~n32330;
  assign n916 = ~n32329 & ~n915;
  assign n917 = ~n905 & ~n916;
  assign n918 = ~n403 & ~n917;
  assign n919 = n403 & ~n905;
  assign n920 = ~n916 & n919;
  assign n921 = ~n755 & ~n32312;
  assign n922 = ~n755 & ~n866;
  assign n923 = ~n32312 & n922;
  assign n924 = ~n866 & n921;
  assign n925 = n764 & ~n32331;
  assign n926 = n768 & n922;
  assign n927 = n764 & ~n32312;
  assign n928 = ~n755 & n927;
  assign n929 = ~n866 & n928;
  assign n930 = ~n764 & ~n32331;
  assign n931 = ~n929 & ~n930;
  assign n932 = ~n925 & ~n926;
  assign n933 = ~n920 & ~n32332;
  assign n934 = ~n918 & ~n933;
  assign n935 = ~n330 & ~n934;
  assign n936 = n330 & ~n918;
  assign n937 = ~n933 & n936;
  assign n938 = n330 & n934;
  assign n939 = ~n770 & ~n772;
  assign n940 = ~n866 & n939;
  assign n941 = n781 & ~n940;
  assign n942 = ~n781 & n940;
  assign n943 = ~n770 & n781;
  assign n944 = ~n772 & n943;
  assign n945 = n781 & n940;
  assign n946 = ~n866 & n944;
  assign n947 = ~n781 & ~n940;
  assign n948 = ~n32334 & ~n947;
  assign n949 = ~n941 & ~n942;
  assign n950 = ~n32333 & ~n32335;
  assign n951 = ~n935 & ~n950;
  assign n952 = ~n271 & ~n951;
  assign n953 = n271 & ~n935;
  assign n954 = ~n950 & n953;
  assign n955 = ~n784 & ~n32316;
  assign n956 = ~n784 & ~n866;
  assign n957 = ~n32316 & n956;
  assign n958 = ~n866 & n955;
  assign n959 = n792 & ~n32336;
  assign n960 = n796 & n956;
  assign n961 = n792 & ~n32316;
  assign n962 = ~n784 & n961;
  assign n963 = ~n866 & n962;
  assign n964 = ~n792 & ~n32336;
  assign n965 = ~n963 & ~n964;
  assign n966 = ~n959 & ~n960;
  assign n967 = ~n954 & ~n32337;
  assign n968 = ~n952 & ~n967;
  assign n969 = ~n217 & ~n968;
  assign n970 = n217 & ~n952;
  assign n971 = ~n967 & n970;
  assign n972 = n217 & n968;
  assign n973 = ~n798 & ~n800;
  assign n974 = ~n866 & n973;
  assign n975 = ~n32318 & n974;
  assign n976 = n32318 & ~n974;
  assign n977 = ~n798 & n32318;
  assign n978 = ~n800 & n977;
  assign n979 = ~n866 & n978;
  assign n980 = ~n32318 & ~n974;
  assign n981 = ~n979 & ~n980;
  assign n982 = ~n975 & ~n976;
  assign n983 = ~n32338 & ~n32339;
  assign n984 = ~n969 & ~n983;
  assign n985 = ~n198 & ~n984;
  assign n986 = n198 & ~n969;
  assign n987 = ~n983 & n986;
  assign n988 = ~n814 & ~n32320;
  assign n989 = ~n814 & ~n866;
  assign n990 = ~n32320 & n989;
  assign n991 = ~n866 & n988;
  assign n992 = n822 & ~n32340;
  assign n993 = n826 & n989;
  assign n994 = n822 & ~n32320;
  assign n995 = ~n814 & n994;
  assign n996 = ~n866 & n995;
  assign n997 = ~n822 & ~n32340;
  assign n998 = ~n996 & ~n997;
  assign n999 = ~n992 & ~n993;
  assign n1000 = ~n987 & ~n32341;
  assign n1001 = ~n985 & ~n1000;
  assign n1002 = ~n828 & ~n830;
  assign n1003 = ~n866 & n1002;
  assign n1004 = ~n32321 & ~n1003;
  assign n1005 = ~n828 & n32321;
  assign n1006 = ~n830 & n1005;
  assign n1007 = n32321 & n1003;
  assign n1008 = ~n866 & n1006;
  assign n1009 = n32321 & ~n1003;
  assign n1010 = ~n32321 & n1003;
  assign n1011 = ~n1009 & ~n1010;
  assign n1012 = ~n1004 & ~n32342;
  assign n1013 = ~n842 & ~n850;
  assign n1014 = ~n850 & ~n866;
  assign n1015 = ~n842 & n1014;
  assign n1016 = ~n866 & n1013;
  assign n1017 = ~n32324 & ~n32344;
  assign n1018 = n32343 & n1017;
  assign n1019 = ~n1001 & n1018;
  assign n1020 = n193 & ~n1019;
  assign n1021 = ~n985 & ~n32343;
  assign n1022 = ~n1000 & n1021;
  assign n1023 = n1001 & ~n32343;
  assign n1024 = n842 & ~n1014;
  assign n1025 = ~n193 & ~n1013;
  assign n1026 = ~n1024 & n1025;
  assign n1027 = ~n32345 & ~n1026;
  assign n1028 = ~n1020 & n1027;
  assign n1029 = pi106  & ~n1028;
  assign n1030 = ~pi104  & ~pi105 ;
  assign n1031 = ~pi106  & n1030;
  assign n1032 = ~n1029 & ~n1031;
  assign n1033 = ~n866 & ~n1032;
  assign n1034 = ~n711 & ~n32326;
  assign n1035 = ~n712 & n1034;
  assign n1036 = ~n728 & n1035;
  assign n1037 = ~n32307 & n1036;
  assign n1038 = n32305 & n730;
  assign n1039 = ~n722 & n1037;
  assign n1040 = ~n1031 & ~n32346;
  assign n1041 = ~n864 & n1040;
  assign n1042 = ~n32324 & n1041;
  assign n1043 = ~n858 & n1042;
  assign n1044 = n866 & n1032;
  assign n1045 = ~n1029 & n1043;
  assign n1046 = ~pi106  & ~n1028;
  assign n1047 = pi107  & ~n1046;
  assign n1048 = ~pi107  & n1046;
  assign n1049 = n868 & ~n1028;
  assign n1050 = ~n1047 & ~n32348;
  assign n1051 = ~n32347 & n1050;
  assign n1052 = ~n1033 & ~n1051;
  assign n1053 = ~n730 & ~n1052;
  assign n1054 = ~n866 & ~n1026;
  assign n1055 = ~n32345 & n1054;
  assign n1056 = ~n1020 & n1055;
  assign n1057 = ~n32348 & ~n1056;
  assign n1058 = pi108  & ~n1057;
  assign n1059 = ~pi108  & ~n1056;
  assign n1060 = ~pi108  & n1057;
  assign n1061 = ~n32348 & n1059;
  assign n1062 = ~n1058 & ~n32349;
  assign n1063 = n730 & ~n1033;
  assign n1064 = n730 & n1052;
  assign n1065 = ~n1051 & n1063;
  assign n1066 = ~n1062 & ~n32350;
  assign n1067 = ~n1053 & ~n1066;
  assign n1068 = ~n602 & ~n1067;
  assign n1069 = n602 & ~n1053;
  assign n1070 = ~n1066 & n1069;
  assign n1071 = ~n871 & ~n32327;
  assign n1072 = ~n1028 & n1071;
  assign n1073 = n876 & ~n1072;
  assign n1074 = ~n876 & n1071;
  assign n1075 = ~n876 & n1072;
  assign n1076 = ~n1028 & n1074;
  assign n1077 = ~n1073 & ~n32351;
  assign n1078 = ~n1070 & ~n1077;
  assign n1079 = ~n1068 & ~n1078;
  assign n1080 = ~n497 & ~n1079;
  assign n1081 = ~n891 & ~n893;
  assign n1082 = ~n1028 & n1081;
  assign n1083 = ~n902 & ~n1082;
  assign n1084 = ~n893 & n902;
  assign n1085 = ~n891 & n1084;
  assign n1086 = n902 & n1082;
  assign n1087 = ~n1028 & n1085;
  assign n1088 = ~n1083 & ~n32352;
  assign n1089 = n497 & ~n1068;
  assign n1090 = n497 & n1079;
  assign n1091 = ~n1078 & n1089;
  assign n1092 = ~n1088 & ~n32353;
  assign n1093 = ~n1080 & ~n1092;
  assign n1094 = ~n403 & ~n1093;
  assign n1095 = n403 & ~n1080;
  assign n1096 = ~n1092 & n1095;
  assign n1097 = ~n905 & ~n32329;
  assign n1098 = ~n1028 & n1097;
  assign n1099 = n915 & ~n1098;
  assign n1100 = ~n915 & n1098;
  assign n1101 = ~n905 & n915;
  assign n1102 = ~n32329 & n1101;
  assign n1103 = n915 & n1098;
  assign n1104 = ~n1028 & n1102;
  assign n1105 = ~n915 & ~n1098;
  assign n1106 = ~n32354 & ~n1105;
  assign n1107 = ~n1099 & ~n1100;
  assign n1108 = ~n1096 & ~n32355;
  assign n1109 = ~n1094 & ~n1108;
  assign n1110 = ~n330 & ~n1109;
  assign n1111 = ~n918 & ~n920;
  assign n1112 = ~n1028 & n1111;
  assign n1113 = ~n32332 & ~n1112;
  assign n1114 = ~n920 & n32332;
  assign n1115 = ~n918 & n1114;
  assign n1116 = n32332 & n1112;
  assign n1117 = ~n1028 & n1115;
  assign n1118 = ~n1113 & ~n32356;
  assign n1119 = n330 & ~n1094;
  assign n1120 = n330 & n1109;
  assign n1121 = ~n1108 & n1119;
  assign n1122 = ~n1118 & ~n32357;
  assign n1123 = ~n1110 & ~n1122;
  assign n1124 = ~n271 & ~n1123;
  assign n1125 = n271 & ~n1110;
  assign n1126 = ~n1122 & n1125;
  assign n1127 = ~n935 & ~n32333;
  assign n1128 = ~n1028 & n1127;
  assign n1129 = ~n32335 & n1128;
  assign n1130 = n32335 & ~n1128;
  assign n1131 = ~n935 & n32335;
  assign n1132 = ~n32333 & n1131;
  assign n1133 = ~n1028 & n1132;
  assign n1134 = ~n32335 & ~n1128;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = ~n1129 & ~n1130;
  assign n1137 = ~n1126 & ~n32358;
  assign n1138 = ~n1124 & ~n1137;
  assign n1139 = ~n217 & ~n1138;
  assign n1140 = ~n952 & ~n954;
  assign n1141 = ~n1028 & n1140;
  assign n1142 = ~n32337 & ~n1141;
  assign n1143 = ~n954 & n32337;
  assign n1144 = ~n952 & n1143;
  assign n1145 = n32337 & n1141;
  assign n1146 = ~n1028 & n1144;
  assign n1147 = ~n1142 & ~n32359;
  assign n1148 = n217 & ~n1124;
  assign n1149 = n217 & n1138;
  assign n1150 = ~n1137 & n1148;
  assign n1151 = ~n1147 & ~n32360;
  assign n1152 = ~n1139 & ~n1151;
  assign n1153 = ~n198 & ~n1152;
  assign n1154 = n198 & ~n1139;
  assign n1155 = ~n1151 & n1154;
  assign n1156 = ~n969 & ~n32338;
  assign n1157 = ~n1028 & n1156;
  assign n1158 = ~n32339 & ~n1157;
  assign n1159 = ~n969 & n32339;
  assign n1160 = ~n32338 & n1159;
  assign n1161 = n32339 & n1157;
  assign n1162 = ~n1028 & n1160;
  assign n1163 = n32339 & ~n1157;
  assign n1164 = ~n32339 & n1157;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = ~n1158 & ~n32361;
  assign n1167 = ~n1155 & n32362;
  assign n1168 = ~n1153 & ~n1167;
  assign n1169 = ~n985 & ~n987;
  assign n1170 = ~n1028 & n1169;
  assign n1171 = ~n32341 & ~n1170;
  assign n1172 = ~n987 & n32341;
  assign n1173 = ~n985 & n1172;
  assign n1174 = n32341 & n1170;
  assign n1175 = ~n1028 & n1173;
  assign n1176 = ~n1171 & ~n32363;
  assign n1177 = ~n1001 & n32343;
  assign n1178 = n32343 & ~n1028;
  assign n1179 = ~n1001 & n1178;
  assign n1180 = ~n1028 & n1177;
  assign n1181 = ~n32345 & ~n32364;
  assign n1182 = ~n1176 & n1181;
  assign n1183 = ~n1168 & n1182;
  assign n1184 = n193 & ~n1183;
  assign n1185 = ~n1153 & n1176;
  assign n1186 = n1168 & n1176;
  assign n1187 = ~n1167 & n1185;
  assign n1188 = n1001 & ~n1178;
  assign n1189 = ~n193 & ~n1177;
  assign n1190 = ~n1188 & n1189;
  assign n1191 = ~n32365 & ~n1190;
  assign n1192 = ~n1184 & n1191;
  assign n1193 = pi104  & ~n1192;
  assign n1194 = ~pi102  & ~pi103 ;
  assign n1195 = ~pi104  & n1194;
  assign n1196 = ~n1193 & ~n1195;
  assign n1197 = ~n1028 & ~n1196;
  assign n1198 = ~pi104  & ~n1192;
  assign n1199 = pi105  & ~n1198;
  assign n1200 = ~pi105  & n1198;
  assign n1201 = n1030 & ~n1192;
  assign n1202 = ~n1199 & ~n32366;
  assign n1203 = ~n32322 & ~n32346;
  assign n1204 = ~n845 & n1203;
  assign n1205 = ~n864 & n1204;
  assign n1206 = ~n32324 & n1205;
  assign n1207 = n850 & n866;
  assign n1208 = ~n858 & n1206;
  assign n1209 = ~n1195 & ~n32367;
  assign n1210 = ~n1026 & n1209;
  assign n1211 = ~n32345 & n1210;
  assign n1212 = ~n1020 & n1211;
  assign n1213 = n1028 & n1196;
  assign n1214 = ~n1193 & n1212;
  assign n1215 = n1202 & ~n32368;
  assign n1216 = ~n1197 & ~n1215;
  assign n1217 = ~n866 & ~n1216;
  assign n1218 = n866 & ~n1197;
  assign n1219 = ~n1215 & n1218;
  assign n1220 = ~n1028 & ~n1190;
  assign n1221 = ~n32365 & n1220;
  assign n1222 = ~n1184 & n1221;
  assign n1223 = ~n32366 & ~n1222;
  assign n1224 = pi106  & ~n1223;
  assign n1225 = ~pi106  & ~n1222;
  assign n1226 = ~pi106  & n1223;
  assign n1227 = ~n32366 & n1225;
  assign n1228 = ~n1224 & ~n32369;
  assign n1229 = ~n1219 & ~n1228;
  assign n1230 = ~n1217 & ~n1229;
  assign n1231 = ~n730 & ~n1230;
  assign n1232 = n730 & ~n1217;
  assign n1233 = ~n1229 & n1232;
  assign n1234 = n730 & n1230;
  assign n1235 = ~n1033 & ~n32347;
  assign n1236 = ~n1192 & n1235;
  assign n1237 = n1050 & ~n1236;
  assign n1238 = ~n1050 & n1235;
  assign n1239 = ~n1050 & n1236;
  assign n1240 = ~n1192 & n1238;
  assign n1241 = ~n1237 & ~n32371;
  assign n1242 = ~n32370 & ~n1241;
  assign n1243 = ~n1231 & ~n1242;
  assign n1244 = ~n602 & ~n1243;
  assign n1245 = n602 & ~n1231;
  assign n1246 = ~n1242 & n1245;
  assign n1247 = ~n1053 & ~n32350;
  assign n1248 = ~n1053 & ~n1192;
  assign n1249 = ~n32350 & n1248;
  assign n1250 = ~n1192 & n1247;
  assign n1251 = n1062 & ~n32372;
  assign n1252 = n1066 & n1248;
  assign n1253 = n1062 & ~n32350;
  assign n1254 = ~n1053 & n1253;
  assign n1255 = ~n1192 & n1254;
  assign n1256 = ~n1062 & ~n32372;
  assign n1257 = ~n1255 & ~n1256;
  assign n1258 = ~n1251 & ~n1252;
  assign n1259 = ~n1246 & ~n32373;
  assign n1260 = ~n1244 & ~n1259;
  assign n1261 = ~n497 & ~n1260;
  assign n1262 = n497 & ~n1244;
  assign n1263 = ~n1259 & n1262;
  assign n1264 = n497 & n1260;
  assign n1265 = ~n1068 & ~n1070;
  assign n1266 = ~n1192 & n1265;
  assign n1267 = n1077 & ~n1266;
  assign n1268 = ~n1077 & n1266;
  assign n1269 = ~n1068 & n1077;
  assign n1270 = ~n1070 & n1269;
  assign n1271 = n1077 & n1266;
  assign n1272 = ~n1192 & n1270;
  assign n1273 = ~n1077 & ~n1266;
  assign n1274 = ~n32375 & ~n1273;
  assign n1275 = ~n1267 & ~n1268;
  assign n1276 = ~n32374 & ~n32376;
  assign n1277 = ~n1261 & ~n1276;
  assign n1278 = ~n403 & ~n1277;
  assign n1279 = n403 & ~n1261;
  assign n1280 = ~n1276 & n1279;
  assign n1281 = ~n1080 & ~n32353;
  assign n1282 = ~n1080 & ~n1192;
  assign n1283 = ~n32353 & n1282;
  assign n1284 = ~n1192 & n1281;
  assign n1285 = n1088 & ~n32377;
  assign n1286 = n1092 & n1282;
  assign n1287 = n1088 & ~n32353;
  assign n1288 = ~n1080 & n1287;
  assign n1289 = ~n1192 & n1288;
  assign n1290 = ~n1088 & ~n32377;
  assign n1291 = ~n1289 & ~n1290;
  assign n1292 = ~n1285 & ~n1286;
  assign n1293 = ~n1280 & ~n32378;
  assign n1294 = ~n1278 & ~n1293;
  assign n1295 = ~n330 & ~n1294;
  assign n1296 = n330 & ~n1278;
  assign n1297 = ~n1293 & n1296;
  assign n1298 = n330 & n1294;
  assign n1299 = ~n1094 & ~n1096;
  assign n1300 = ~n1192 & n1299;
  assign n1301 = ~n32355 & n1300;
  assign n1302 = n32355 & ~n1300;
  assign n1303 = ~n1094 & n32355;
  assign n1304 = ~n1096 & n1303;
  assign n1305 = ~n1192 & n1304;
  assign n1306 = ~n32355 & ~n1300;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n1301 & ~n1302;
  assign n1309 = ~n32379 & ~n32380;
  assign n1310 = ~n1295 & ~n1309;
  assign n1311 = ~n271 & ~n1310;
  assign n1312 = n271 & ~n1295;
  assign n1313 = ~n1309 & n1312;
  assign n1314 = ~n1110 & ~n32357;
  assign n1315 = ~n1110 & ~n1192;
  assign n1316 = ~n32357 & n1315;
  assign n1317 = ~n1192 & n1314;
  assign n1318 = n1118 & ~n32381;
  assign n1319 = n1122 & n1315;
  assign n1320 = n1118 & ~n32357;
  assign n1321 = ~n1110 & n1320;
  assign n1322 = ~n1192 & n1321;
  assign n1323 = ~n1118 & ~n32381;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = ~n1318 & ~n1319;
  assign n1326 = ~n1313 & ~n32382;
  assign n1327 = ~n1311 & ~n1326;
  assign n1328 = ~n217 & ~n1327;
  assign n1329 = n217 & ~n1311;
  assign n1330 = ~n1326 & n1329;
  assign n1331 = n217 & n1327;
  assign n1332 = ~n1124 & ~n1126;
  assign n1333 = ~n1192 & n1332;
  assign n1334 = ~n32358 & ~n1333;
  assign n1335 = ~n1124 & n32358;
  assign n1336 = ~n1126 & n1335;
  assign n1337 = n32358 & n1333;
  assign n1338 = ~n1192 & n1336;
  assign n1339 = ~n32358 & n1333;
  assign n1340 = n32358 & ~n1333;
  assign n1341 = ~n1339 & ~n1340;
  assign n1342 = ~n1334 & ~n32384;
  assign n1343 = ~n32383 & n32385;
  assign n1344 = ~n1328 & ~n1343;
  assign n1345 = ~n198 & ~n1344;
  assign n1346 = n198 & ~n1328;
  assign n1347 = ~n1343 & n1346;
  assign n1348 = ~n1139 & ~n32360;
  assign n1349 = ~n1139 & ~n1192;
  assign n1350 = ~n32360 & n1349;
  assign n1351 = ~n1192 & n1348;
  assign n1352 = n1147 & ~n32386;
  assign n1353 = n1151 & n1349;
  assign n1354 = n1147 & ~n32360;
  assign n1355 = ~n1139 & n1354;
  assign n1356 = ~n1192 & n1355;
  assign n1357 = ~n1147 & ~n32386;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = ~n1352 & ~n1353;
  assign n1360 = ~n1347 & ~n32387;
  assign n1361 = ~n1345 & ~n1360;
  assign n1362 = ~n1153 & ~n1155;
  assign n1363 = ~n1192 & n1362;
  assign n1364 = n32362 & ~n1363;
  assign n1365 = ~n1153 & ~n32362;
  assign n1366 = ~n1155 & n1365;
  assign n1367 = ~n32362 & n1363;
  assign n1368 = ~n1192 & n1366;
  assign n1369 = n32362 & n1363;
  assign n1370 = ~n32362 & ~n1363;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = ~n1364 & ~n32388;
  assign n1373 = ~n1168 & ~n1176;
  assign n1374 = ~n1176 & ~n1192;
  assign n1375 = ~n1168 & n1374;
  assign n1376 = ~n1192 & n1373;
  assign n1377 = ~n32365 & ~n32390;
  assign n1378 = n32389 & n1377;
  assign n1379 = ~n1361 & n1378;
  assign n1380 = n193 & ~n1379;
  assign n1381 = ~n1345 & ~n32389;
  assign n1382 = ~n1360 & n1381;
  assign n1383 = n1361 & ~n32389;
  assign n1384 = n1168 & ~n1374;
  assign n1385 = ~n193 & ~n1373;
  assign n1386 = ~n1384 & n1385;
  assign n1387 = ~n32391 & ~n1386;
  assign n1388 = ~n1380 & n1387;
  assign n1389 = pi102  & ~n1388;
  assign n1390 = ~pi100  & ~pi101 ;
  assign n1391 = ~pi102  & n1390;
  assign n1392 = ~n1389 & ~n1391;
  assign n1393 = ~n1192 & ~n1392;
  assign n1394 = ~n32342 & ~n32367;
  assign n1395 = ~n1004 & n1394;
  assign n1396 = ~n1026 & n1395;
  assign n1397 = ~n32345 & n1396;
  assign n1398 = ~n32343 & n1028;
  assign n1399 = ~n1020 & n1397;
  assign n1400 = ~n1391 & ~n32392;
  assign n1401 = ~n1190 & n1400;
  assign n1402 = ~n32365 & n1401;
  assign n1403 = ~n1184 & n1402;
  assign n1404 = n1192 & n1392;
  assign n1405 = ~n1389 & n1403;
  assign n1406 = ~pi102  & ~n1388;
  assign n1407 = pi103  & ~n1406;
  assign n1408 = ~pi103  & n1406;
  assign n1409 = n1194 & ~n1388;
  assign n1410 = ~n1407 & ~n32394;
  assign n1411 = ~n32393 & n1410;
  assign n1412 = ~n1393 & ~n1411;
  assign n1413 = ~n1028 & ~n1412;
  assign n1414 = ~n1192 & ~n1386;
  assign n1415 = ~n32391 & n1414;
  assign n1416 = ~n1380 & n1415;
  assign n1417 = ~n32394 & ~n1416;
  assign n1418 = pi104  & ~n1417;
  assign n1419 = ~pi104  & ~n1416;
  assign n1420 = ~pi104  & n1417;
  assign n1421 = ~n32394 & n1419;
  assign n1422 = ~n1418 & ~n32395;
  assign n1423 = n1028 & ~n1393;
  assign n1424 = n1028 & n1412;
  assign n1425 = ~n1411 & n1423;
  assign n1426 = ~n1422 & ~n32396;
  assign n1427 = ~n1413 & ~n1426;
  assign n1428 = ~n866 & ~n1427;
  assign n1429 = n866 & ~n1413;
  assign n1430 = ~n1426 & n1429;
  assign n1431 = ~n1197 & ~n32368;
  assign n1432 = ~n1388 & n1431;
  assign n1433 = n1202 & ~n1432;
  assign n1434 = ~n1202 & n1431;
  assign n1435 = ~n1202 & n1432;
  assign n1436 = ~n1388 & n1434;
  assign n1437 = ~n1433 & ~n32397;
  assign n1438 = ~n1430 & ~n1437;
  assign n1439 = ~n1428 & ~n1438;
  assign n1440 = ~n730 & ~n1439;
  assign n1441 = ~n1217 & ~n1219;
  assign n1442 = ~n1388 & n1441;
  assign n1443 = ~n1228 & ~n1442;
  assign n1444 = ~n1219 & n1228;
  assign n1445 = ~n1217 & n1444;
  assign n1446 = n1228 & n1442;
  assign n1447 = ~n1388 & n1445;
  assign n1448 = ~n1443 & ~n32398;
  assign n1449 = n730 & ~n1428;
  assign n1450 = n730 & n1439;
  assign n1451 = ~n1438 & n1449;
  assign n1452 = ~n1448 & ~n32399;
  assign n1453 = ~n1440 & ~n1452;
  assign n1454 = ~n602 & ~n1453;
  assign n1455 = n602 & ~n1440;
  assign n1456 = ~n1452 & n1455;
  assign n1457 = ~n1231 & ~n32370;
  assign n1458 = ~n1388 & n1457;
  assign n1459 = n1241 & ~n1458;
  assign n1460 = ~n1241 & n1458;
  assign n1461 = ~n1231 & n1241;
  assign n1462 = ~n32370 & n1461;
  assign n1463 = n1241 & n1458;
  assign n1464 = ~n1388 & n1462;
  assign n1465 = ~n1241 & ~n1458;
  assign n1466 = ~n32400 & ~n1465;
  assign n1467 = ~n1459 & ~n1460;
  assign n1468 = ~n1456 & ~n32401;
  assign n1469 = ~n1454 & ~n1468;
  assign n1470 = ~n497 & ~n1469;
  assign n1471 = ~n1244 & ~n1246;
  assign n1472 = ~n1388 & n1471;
  assign n1473 = ~n32373 & ~n1472;
  assign n1474 = ~n1246 & n32373;
  assign n1475 = ~n1244 & n1474;
  assign n1476 = n32373 & n1472;
  assign n1477 = ~n1388 & n1475;
  assign n1478 = ~n1473 & ~n32402;
  assign n1479 = n497 & ~n1454;
  assign n1480 = n497 & n1469;
  assign n1481 = ~n1468 & n1479;
  assign n1482 = ~n1478 & ~n32403;
  assign n1483 = ~n1470 & ~n1482;
  assign n1484 = ~n403 & ~n1483;
  assign n1485 = n403 & ~n1470;
  assign n1486 = ~n1482 & n1485;
  assign n1487 = ~n1261 & ~n32374;
  assign n1488 = ~n1388 & n1487;
  assign n1489 = ~n32376 & n1488;
  assign n1490 = n32376 & ~n1488;
  assign n1491 = ~n1261 & n32376;
  assign n1492 = ~n32374 & n1491;
  assign n1493 = ~n1388 & n1492;
  assign n1494 = ~n32376 & ~n1488;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = ~n1489 & ~n1490;
  assign n1497 = ~n1486 & ~n32404;
  assign n1498 = ~n1484 & ~n1497;
  assign n1499 = ~n330 & ~n1498;
  assign n1500 = ~n1278 & ~n1280;
  assign n1501 = ~n1388 & n1500;
  assign n1502 = ~n32378 & ~n1501;
  assign n1503 = ~n1280 & n32378;
  assign n1504 = ~n1278 & n1503;
  assign n1505 = n32378 & n1501;
  assign n1506 = ~n1388 & n1504;
  assign n1507 = ~n1502 & ~n32405;
  assign n1508 = n330 & ~n1484;
  assign n1509 = n330 & n1498;
  assign n1510 = ~n1497 & n1508;
  assign n1511 = ~n1507 & ~n32406;
  assign n1512 = ~n1499 & ~n1511;
  assign n1513 = ~n271 & ~n1512;
  assign n1514 = n271 & ~n1499;
  assign n1515 = ~n1511 & n1514;
  assign n1516 = ~n1295 & ~n32379;
  assign n1517 = ~n1388 & n1516;
  assign n1518 = ~n32380 & ~n1517;
  assign n1519 = ~n1295 & n32380;
  assign n1520 = ~n32379 & n1519;
  assign n1521 = n32380 & n1517;
  assign n1522 = ~n1388 & n1520;
  assign n1523 = n32380 & ~n1517;
  assign n1524 = ~n32380 & n1517;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = ~n1518 & ~n32407;
  assign n1527 = ~n1515 & n32408;
  assign n1528 = ~n1513 & ~n1527;
  assign n1529 = ~n217 & ~n1528;
  assign n1530 = ~n1311 & ~n1313;
  assign n1531 = ~n1388 & n1530;
  assign n1532 = ~n32382 & ~n1531;
  assign n1533 = ~n1313 & n32382;
  assign n1534 = ~n1311 & n1533;
  assign n1535 = n32382 & n1531;
  assign n1536 = ~n1388 & n1534;
  assign n1537 = ~n1532 & ~n32409;
  assign n1538 = n217 & ~n1513;
  assign n1539 = n217 & n1528;
  assign n1540 = ~n1527 & n1538;
  assign n1541 = ~n1537 & ~n32410;
  assign n1542 = ~n1529 & ~n1541;
  assign n1543 = ~n198 & ~n1542;
  assign n1544 = n198 & ~n1529;
  assign n1545 = ~n1541 & n1544;
  assign n1546 = ~n1328 & ~n32383;
  assign n1547 = ~n1388 & n1546;
  assign n1548 = ~n32385 & ~n1547;
  assign n1549 = n32385 & n1547;
  assign n1550 = ~n1328 & ~n32385;
  assign n1551 = ~n32383 & n1550;
  assign n1552 = ~n32385 & n1547;
  assign n1553 = ~n1388 & n1551;
  assign n1554 = n32385 & ~n1547;
  assign n1555 = ~n32411 & ~n1554;
  assign n1556 = ~n1548 & ~n1549;
  assign n1557 = ~n1545 & ~n32412;
  assign n1558 = ~n1543 & ~n1557;
  assign n1559 = ~n1345 & ~n1347;
  assign n1560 = ~n1388 & n1559;
  assign n1561 = ~n32387 & ~n1560;
  assign n1562 = ~n1347 & n32387;
  assign n1563 = ~n1345 & n1562;
  assign n1564 = n32387 & n1560;
  assign n1565 = ~n1388 & n1563;
  assign n1566 = ~n1561 & ~n32413;
  assign n1567 = ~n1361 & n32389;
  assign n1568 = n32389 & ~n1388;
  assign n1569 = ~n1361 & n1568;
  assign n1570 = ~n1388 & n1567;
  assign n1571 = ~n32391 & ~n32414;
  assign n1572 = ~n1566 & n1571;
  assign n1573 = ~n1558 & n1572;
  assign n1574 = n193 & ~n1573;
  assign n1575 = ~n1543 & n1566;
  assign n1576 = n1558 & n1566;
  assign n1577 = ~n1557 & n1575;
  assign n1578 = n1361 & ~n1568;
  assign n1579 = ~n193 & ~n1567;
  assign n1580 = ~n1578 & n1579;
  assign n1581 = ~n32415 & ~n1580;
  assign n1582 = ~n1574 & n1581;
  assign n1583 = pi100  & ~n1582;
  assign n1584 = ~pi98  & ~pi99 ;
  assign n1585 = ~pi100  & n1584;
  assign n1586 = ~n1583 & ~n1585;
  assign n1587 = ~n1388 & ~n1586;
  assign n1588 = ~pi100  & ~n1582;
  assign n1589 = pi101  & ~n1588;
  assign n1590 = ~pi101  & n1588;
  assign n1591 = n1390 & ~n1582;
  assign n1592 = ~n1589 & ~n32416;
  assign n1593 = ~n32363 & ~n32392;
  assign n1594 = ~n1171 & n1593;
  assign n1595 = ~n1190 & n1594;
  assign n1596 = ~n32365 & n1595;
  assign n1597 = n1176 & n1192;
  assign n1598 = ~n1184 & n1596;
  assign n1599 = ~n1585 & ~n32417;
  assign n1600 = ~n1386 & n1599;
  assign n1601 = ~n32391 & n1600;
  assign n1602 = ~n1380 & n1601;
  assign n1603 = n1388 & n1586;
  assign n1604 = ~n1583 & n1602;
  assign n1605 = n1592 & ~n32418;
  assign n1606 = ~n1587 & ~n1605;
  assign n1607 = ~n1192 & ~n1606;
  assign n1608 = n1192 & ~n1587;
  assign n1609 = ~n1605 & n1608;
  assign n1610 = ~n1388 & ~n1580;
  assign n1611 = ~n32415 & n1610;
  assign n1612 = ~n1574 & n1611;
  assign n1613 = ~n32416 & ~n1612;
  assign n1614 = pi102  & ~n1613;
  assign n1615 = ~pi102  & ~n1612;
  assign n1616 = ~pi102  & n1613;
  assign n1617 = ~n32416 & n1615;
  assign n1618 = ~n1614 & ~n32419;
  assign n1619 = ~n1609 & ~n1618;
  assign n1620 = ~n1607 & ~n1619;
  assign n1621 = ~n1028 & ~n1620;
  assign n1622 = n1028 & ~n1607;
  assign n1623 = ~n1619 & n1622;
  assign n1624 = n1028 & n1620;
  assign n1625 = ~n1393 & ~n32393;
  assign n1626 = ~n1582 & n1625;
  assign n1627 = n1410 & ~n1626;
  assign n1628 = ~n1410 & n1625;
  assign n1629 = ~n1410 & n1626;
  assign n1630 = ~n1582 & n1628;
  assign n1631 = ~n1627 & ~n32421;
  assign n1632 = ~n32420 & ~n1631;
  assign n1633 = ~n1621 & ~n1632;
  assign n1634 = ~n866 & ~n1633;
  assign n1635 = n866 & ~n1621;
  assign n1636 = ~n1632 & n1635;
  assign n1637 = ~n1413 & ~n32396;
  assign n1638 = ~n1413 & ~n1582;
  assign n1639 = ~n32396 & n1638;
  assign n1640 = ~n1582 & n1637;
  assign n1641 = n1422 & ~n32422;
  assign n1642 = n1426 & n1638;
  assign n1643 = n1422 & ~n32396;
  assign n1644 = ~n1413 & n1643;
  assign n1645 = ~n1582 & n1644;
  assign n1646 = ~n1422 & ~n32422;
  assign n1647 = ~n1645 & ~n1646;
  assign n1648 = ~n1641 & ~n1642;
  assign n1649 = ~n1636 & ~n32423;
  assign n1650 = ~n1634 & ~n1649;
  assign n1651 = ~n730 & ~n1650;
  assign n1652 = n730 & ~n1634;
  assign n1653 = ~n1649 & n1652;
  assign n1654 = n730 & n1650;
  assign n1655 = ~n1428 & ~n1430;
  assign n1656 = ~n1582 & n1655;
  assign n1657 = n1437 & ~n1656;
  assign n1658 = ~n1437 & n1656;
  assign n1659 = ~n1428 & n1437;
  assign n1660 = ~n1430 & n1659;
  assign n1661 = n1437 & n1656;
  assign n1662 = ~n1582 & n1660;
  assign n1663 = ~n1437 & ~n1656;
  assign n1664 = ~n32425 & ~n1663;
  assign n1665 = ~n1657 & ~n1658;
  assign n1666 = ~n32424 & ~n32426;
  assign n1667 = ~n1651 & ~n1666;
  assign n1668 = ~n602 & ~n1667;
  assign n1669 = n602 & ~n1651;
  assign n1670 = ~n1666 & n1669;
  assign n1671 = ~n1440 & ~n32399;
  assign n1672 = ~n1440 & ~n1582;
  assign n1673 = ~n32399 & n1672;
  assign n1674 = ~n1582 & n1671;
  assign n1675 = n1448 & ~n32427;
  assign n1676 = n1452 & n1672;
  assign n1677 = n1448 & ~n32399;
  assign n1678 = ~n1440 & n1677;
  assign n1679 = ~n1582 & n1678;
  assign n1680 = ~n1448 & ~n32427;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = ~n1675 & ~n1676;
  assign n1683 = ~n1670 & ~n32428;
  assign n1684 = ~n1668 & ~n1683;
  assign n1685 = ~n497 & ~n1684;
  assign n1686 = n497 & ~n1668;
  assign n1687 = ~n1683 & n1686;
  assign n1688 = n497 & n1684;
  assign n1689 = ~n1454 & ~n1456;
  assign n1690 = ~n1582 & n1689;
  assign n1691 = ~n32401 & n1690;
  assign n1692 = n32401 & ~n1690;
  assign n1693 = ~n1454 & n32401;
  assign n1694 = ~n1456 & n1693;
  assign n1695 = ~n1582 & n1694;
  assign n1696 = ~n32401 & ~n1690;
  assign n1697 = ~n1695 & ~n1696;
  assign n1698 = ~n1691 & ~n1692;
  assign n1699 = ~n32429 & ~n32430;
  assign n1700 = ~n1685 & ~n1699;
  assign n1701 = ~n403 & ~n1700;
  assign n1702 = n403 & ~n1685;
  assign n1703 = ~n1699 & n1702;
  assign n1704 = ~n1470 & ~n32403;
  assign n1705 = ~n1470 & ~n1582;
  assign n1706 = ~n32403 & n1705;
  assign n1707 = ~n1582 & n1704;
  assign n1708 = n1478 & ~n32431;
  assign n1709 = n1482 & n1705;
  assign n1710 = n1478 & ~n32403;
  assign n1711 = ~n1470 & n1710;
  assign n1712 = ~n1582 & n1711;
  assign n1713 = ~n1478 & ~n32431;
  assign n1714 = ~n1712 & ~n1713;
  assign n1715 = ~n1708 & ~n1709;
  assign n1716 = ~n1703 & ~n32432;
  assign n1717 = ~n1701 & ~n1716;
  assign n1718 = ~n330 & ~n1717;
  assign n1719 = n330 & ~n1701;
  assign n1720 = ~n1716 & n1719;
  assign n1721 = n330 & n1717;
  assign n1722 = ~n1484 & ~n1486;
  assign n1723 = ~n1582 & n1722;
  assign n1724 = ~n32404 & ~n1723;
  assign n1725 = ~n1484 & n32404;
  assign n1726 = ~n1486 & n1725;
  assign n1727 = n32404 & n1723;
  assign n1728 = ~n1582 & n1726;
  assign n1729 = n32404 & ~n1723;
  assign n1730 = ~n32404 & n1723;
  assign n1731 = ~n1729 & ~n1730;
  assign n1732 = ~n1724 & ~n32434;
  assign n1733 = ~n32433 & n32435;
  assign n1734 = ~n1718 & ~n1733;
  assign n1735 = ~n271 & ~n1734;
  assign n1736 = n271 & ~n1718;
  assign n1737 = ~n1733 & n1736;
  assign n1738 = ~n1499 & ~n32406;
  assign n1739 = ~n1499 & ~n1582;
  assign n1740 = ~n32406 & n1739;
  assign n1741 = ~n1582 & n1738;
  assign n1742 = n1507 & ~n32436;
  assign n1743 = n1511 & n1739;
  assign n1744 = n1507 & ~n32406;
  assign n1745 = ~n1499 & n1744;
  assign n1746 = ~n1582 & n1745;
  assign n1747 = ~n1507 & ~n32436;
  assign n1748 = ~n1746 & ~n1747;
  assign n1749 = ~n1742 & ~n1743;
  assign n1750 = ~n1737 & ~n32437;
  assign n1751 = ~n1735 & ~n1750;
  assign n1752 = ~n217 & ~n1751;
  assign n1753 = n217 & ~n1735;
  assign n1754 = ~n1750 & n1753;
  assign n1755 = n217 & n1751;
  assign n1756 = ~n1513 & ~n1515;
  assign n1757 = ~n1582 & n1756;
  assign n1758 = n32408 & ~n1757;
  assign n1759 = ~n1513 & ~n32408;
  assign n1760 = ~n1515 & n1759;
  assign n1761 = ~n32408 & n1757;
  assign n1762 = ~n1582 & n1760;
  assign n1763 = n32408 & n1757;
  assign n1764 = ~n32408 & ~n1757;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = ~n1758 & ~n32439;
  assign n1767 = ~n32438 & n32440;
  assign n1768 = ~n1752 & ~n1767;
  assign n1769 = ~n198 & ~n1768;
  assign n1770 = n198 & ~n1752;
  assign n1771 = ~n1767 & n1770;
  assign n1772 = ~n1529 & ~n32410;
  assign n1773 = ~n1529 & ~n1582;
  assign n1774 = ~n32410 & n1773;
  assign n1775 = ~n1582 & n1772;
  assign n1776 = n1537 & ~n32441;
  assign n1777 = n1541 & n1773;
  assign n1778 = n1537 & ~n32410;
  assign n1779 = ~n1529 & n1778;
  assign n1780 = ~n1582 & n1779;
  assign n1781 = ~n1537 & ~n32441;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = ~n1776 & ~n1777;
  assign n1784 = ~n1771 & ~n32442;
  assign n1785 = ~n1769 & ~n1784;
  assign n1786 = ~n1543 & ~n1545;
  assign n1787 = ~n1582 & n1786;
  assign n1788 = ~n32412 & n1787;
  assign n1789 = n32412 & ~n1787;
  assign n1790 = ~n1543 & n32412;
  assign n1791 = ~n1545 & n1790;
  assign n1792 = n32412 & n1787;
  assign n1793 = ~n1582 & n1791;
  assign n1794 = ~n32412 & ~n1787;
  assign n1795 = ~n32443 & ~n1794;
  assign n1796 = ~n1788 & ~n1789;
  assign n1797 = ~n1558 & ~n1566;
  assign n1798 = ~n1566 & ~n1582;
  assign n1799 = ~n1558 & n1798;
  assign n1800 = ~n1582 & n1797;
  assign n1801 = ~n32415 & ~n32445;
  assign n1802 = ~n32444 & n1801;
  assign n1803 = ~n1785 & n1802;
  assign n1804 = n193 & ~n1803;
  assign n1805 = ~n1769 & n32444;
  assign n1806 = ~n1784 & n1805;
  assign n1807 = n1785 & n32444;
  assign n1808 = n1558 & ~n1798;
  assign n1809 = ~n193 & ~n1797;
  assign n1810 = ~n1808 & n1809;
  assign n1811 = ~n32446 & ~n1810;
  assign n1812 = ~n1804 & n1811;
  assign n1813 = pi98  & ~n1812;
  assign n1814 = ~pi96  & ~pi97 ;
  assign n1815 = ~pi98  & n1814;
  assign n1816 = ~n1813 & ~n1815;
  assign n1817 = ~n1582 & ~n1816;
  assign n1818 = ~n32388 & ~n32417;
  assign n1819 = ~n1364 & n1818;
  assign n1820 = ~n1386 & n1819;
  assign n1821 = ~n32391 & n1820;
  assign n1822 = ~n32389 & n1388;
  assign n1823 = ~n1380 & n1821;
  assign n1824 = ~n1815 & ~n32447;
  assign n1825 = ~n1580 & n1824;
  assign n1826 = ~n32415 & n1825;
  assign n1827 = ~n1574 & n1826;
  assign n1828 = n1582 & n1816;
  assign n1829 = ~n1813 & n1827;
  assign n1830 = ~pi98  & ~n1812;
  assign n1831 = pi99  & ~n1830;
  assign n1832 = ~pi99  & n1830;
  assign n1833 = n1584 & ~n1812;
  assign n1834 = ~n1831 & ~n32449;
  assign n1835 = ~n32448 & n1834;
  assign n1836 = ~n1817 & ~n1835;
  assign n1837 = ~n1388 & ~n1836;
  assign n1838 = ~n1582 & ~n1810;
  assign n1839 = ~n32446 & n1838;
  assign n1840 = ~n1804 & n1839;
  assign n1841 = ~n32449 & ~n1840;
  assign n1842 = pi100  & ~n1841;
  assign n1843 = ~pi100  & ~n1840;
  assign n1844 = ~pi100  & n1841;
  assign n1845 = ~n32449 & n1843;
  assign n1846 = ~n1842 & ~n32450;
  assign n1847 = n1388 & ~n1817;
  assign n1848 = n1388 & n1836;
  assign n1849 = ~n1835 & n1847;
  assign n1850 = ~n1846 & ~n32451;
  assign n1851 = ~n1837 & ~n1850;
  assign n1852 = ~n1192 & ~n1851;
  assign n1853 = n1192 & ~n1837;
  assign n1854 = ~n1850 & n1853;
  assign n1855 = ~n1587 & ~n32418;
  assign n1856 = ~n1812 & n1855;
  assign n1857 = n1592 & ~n1856;
  assign n1858 = ~n1592 & n1855;
  assign n1859 = ~n1592 & n1856;
  assign n1860 = ~n1812 & n1858;
  assign n1861 = ~n1857 & ~n32452;
  assign n1862 = ~n1854 & ~n1861;
  assign n1863 = ~n1852 & ~n1862;
  assign n1864 = ~n1028 & ~n1863;
  assign n1865 = ~n1607 & ~n1609;
  assign n1866 = ~n1812 & n1865;
  assign n1867 = ~n1618 & ~n1866;
  assign n1868 = ~n1609 & n1618;
  assign n1869 = ~n1607 & n1868;
  assign n1870 = n1618 & n1866;
  assign n1871 = ~n1812 & n1869;
  assign n1872 = ~n1867 & ~n32453;
  assign n1873 = n1028 & ~n1852;
  assign n1874 = n1028 & n1863;
  assign n1875 = ~n1862 & n1873;
  assign n1876 = ~n1872 & ~n32454;
  assign n1877 = ~n1864 & ~n1876;
  assign n1878 = ~n866 & ~n1877;
  assign n1879 = n866 & ~n1864;
  assign n1880 = ~n1876 & n1879;
  assign n1881 = ~n1621 & ~n32420;
  assign n1882 = ~n1812 & n1881;
  assign n1883 = n1631 & ~n1882;
  assign n1884 = ~n1631 & n1882;
  assign n1885 = ~n1621 & n1631;
  assign n1886 = ~n32420 & n1885;
  assign n1887 = n1631 & n1882;
  assign n1888 = ~n1812 & n1886;
  assign n1889 = ~n1631 & ~n1882;
  assign n1890 = ~n32455 & ~n1889;
  assign n1891 = ~n1883 & ~n1884;
  assign n1892 = ~n1880 & ~n32456;
  assign n1893 = ~n1878 & ~n1892;
  assign n1894 = ~n730 & ~n1893;
  assign n1895 = ~n1634 & ~n1636;
  assign n1896 = ~n1812 & n1895;
  assign n1897 = ~n32423 & ~n1896;
  assign n1898 = ~n1636 & n32423;
  assign n1899 = ~n1634 & n1898;
  assign n1900 = n32423 & n1896;
  assign n1901 = ~n1812 & n1899;
  assign n1902 = ~n1897 & ~n32457;
  assign n1903 = n730 & ~n1878;
  assign n1904 = n730 & n1893;
  assign n1905 = ~n1892 & n1903;
  assign n1906 = ~n1902 & ~n32458;
  assign n1907 = ~n1894 & ~n1906;
  assign n1908 = ~n602 & ~n1907;
  assign n1909 = n602 & ~n1894;
  assign n1910 = ~n1906 & n1909;
  assign n1911 = ~n1651 & ~n32424;
  assign n1912 = ~n1812 & n1911;
  assign n1913 = ~n32426 & n1912;
  assign n1914 = n32426 & ~n1912;
  assign n1915 = ~n1651 & n32426;
  assign n1916 = ~n32424 & n1915;
  assign n1917 = ~n1812 & n1916;
  assign n1918 = ~n32426 & ~n1912;
  assign n1919 = ~n1917 & ~n1918;
  assign n1920 = ~n1913 & ~n1914;
  assign n1921 = ~n1910 & ~n32459;
  assign n1922 = ~n1908 & ~n1921;
  assign n1923 = ~n497 & ~n1922;
  assign n1924 = ~n1668 & ~n1670;
  assign n1925 = ~n1812 & n1924;
  assign n1926 = ~n32428 & ~n1925;
  assign n1927 = ~n1670 & n32428;
  assign n1928 = ~n1668 & n1927;
  assign n1929 = n32428 & n1925;
  assign n1930 = ~n1812 & n1928;
  assign n1931 = ~n1926 & ~n32460;
  assign n1932 = n497 & ~n1908;
  assign n1933 = n497 & n1922;
  assign n1934 = ~n1921 & n1932;
  assign n1935 = ~n1931 & ~n32461;
  assign n1936 = ~n1923 & ~n1935;
  assign n1937 = ~n403 & ~n1936;
  assign n1938 = n403 & ~n1923;
  assign n1939 = ~n1935 & n1938;
  assign n1940 = ~n1685 & ~n32429;
  assign n1941 = ~n1812 & n1940;
  assign n1942 = ~n32430 & ~n1941;
  assign n1943 = ~n1685 & n32430;
  assign n1944 = ~n32429 & n1943;
  assign n1945 = n32430 & n1941;
  assign n1946 = ~n1812 & n1944;
  assign n1947 = n32430 & ~n1941;
  assign n1948 = ~n32430 & n1941;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = ~n1942 & ~n32462;
  assign n1951 = ~n1939 & n32463;
  assign n1952 = ~n1937 & ~n1951;
  assign n1953 = ~n330 & ~n1952;
  assign n1954 = ~n1701 & ~n1703;
  assign n1955 = ~n1812 & n1954;
  assign n1956 = ~n32432 & ~n1955;
  assign n1957 = ~n1703 & n32432;
  assign n1958 = ~n1701 & n1957;
  assign n1959 = n32432 & n1955;
  assign n1960 = ~n1812 & n1958;
  assign n1961 = ~n1956 & ~n32464;
  assign n1962 = n330 & ~n1937;
  assign n1963 = n330 & n1952;
  assign n1964 = ~n1951 & n1962;
  assign n1965 = ~n1961 & ~n32465;
  assign n1966 = ~n1953 & ~n1965;
  assign n1967 = ~n271 & ~n1966;
  assign n1968 = n271 & ~n1953;
  assign n1969 = ~n1965 & n1968;
  assign n1970 = ~n1718 & ~n32433;
  assign n1971 = ~n1812 & n1970;
  assign n1972 = n32435 & ~n1971;
  assign n1973 = ~n1718 & ~n32435;
  assign n1974 = ~n32433 & n1973;
  assign n1975 = ~n32435 & n1971;
  assign n1976 = ~n1812 & n1974;
  assign n1977 = n32435 & n1971;
  assign n1978 = ~n32435 & ~n1971;
  assign n1979 = ~n1977 & ~n1978;
  assign n1980 = ~n1972 & ~n32466;
  assign n1981 = ~n1969 & n32467;
  assign n1982 = ~n1967 & ~n1981;
  assign n1983 = ~n217 & ~n1982;
  assign n1984 = ~n1735 & ~n1737;
  assign n1985 = ~n1812 & n1984;
  assign n1986 = ~n32437 & ~n1985;
  assign n1987 = ~n1737 & n32437;
  assign n1988 = ~n1735 & n1987;
  assign n1989 = n32437 & n1985;
  assign n1990 = ~n1812 & n1988;
  assign n1991 = ~n1986 & ~n32468;
  assign n1992 = n217 & ~n1967;
  assign n1993 = n217 & n1982;
  assign n1994 = ~n1981 & n1992;
  assign n1995 = ~n1991 & ~n32469;
  assign n1996 = ~n1983 & ~n1995;
  assign n1997 = ~n198 & ~n1996;
  assign n1998 = n198 & ~n1983;
  assign n1999 = ~n1995 & n1998;
  assign n2000 = ~n1752 & ~n32438;
  assign n2001 = ~n1752 & ~n1812;
  assign n2002 = ~n32438 & n2001;
  assign n2003 = ~n1812 & n2000;
  assign n2004 = ~n32440 & ~n32470;
  assign n2005 = n1767 & n2001;
  assign n2006 = n32440 & n32470;
  assign n2007 = ~n1752 & ~n32440;
  assign n2008 = ~n32438 & n2007;
  assign n2009 = ~n1812 & n2008;
  assign n2010 = n32440 & ~n32470;
  assign n2011 = ~n2009 & ~n2010;
  assign n2012 = ~n2004 & ~n32471;
  assign n2013 = ~n1999 & ~n32472;
  assign n2014 = ~n1997 & ~n2013;
  assign n2015 = ~n1769 & ~n1771;
  assign n2016 = ~n1812 & n2015;
  assign n2017 = ~n32442 & ~n2016;
  assign n2018 = ~n1771 & n32442;
  assign n2019 = ~n1769 & n2018;
  assign n2020 = n32442 & n2016;
  assign n2021 = ~n1812 & n2019;
  assign n2022 = ~n2017 & ~n32473;
  assign n2023 = ~n1785 & ~n32444;
  assign n2024 = ~n32444 & ~n1812;
  assign n2025 = ~n1785 & n2024;
  assign n2026 = ~n1812 & n2023;
  assign n2027 = ~n32446 & ~n32474;
  assign n2028 = ~n2022 & n2027;
  assign n2029 = ~n2014 & n2028;
  assign n2030 = n193 & ~n2029;
  assign n2031 = ~n1997 & n2022;
  assign n2032 = n2014 & n2022;
  assign n2033 = ~n2013 & n2031;
  assign n2034 = n1785 & ~n2024;
  assign n2035 = ~n193 & ~n2023;
  assign n2036 = ~n2034 & n2035;
  assign n2037 = ~n32475 & ~n2036;
  assign n2038 = ~n2030 & n2037;
  assign n2039 = pi96  & ~n2038;
  assign n2040 = ~pi94  & ~pi95 ;
  assign n2041 = ~pi96  & n2040;
  assign n2042 = ~n2039 & ~n2041;
  assign n2043 = ~n1812 & ~n2042;
  assign n2044 = ~pi96  & ~n2038;
  assign n2045 = pi97  & ~n2044;
  assign n2046 = ~pi97  & n2044;
  assign n2047 = n1814 & ~n2038;
  assign n2048 = ~n2045 & ~n32476;
  assign n2049 = ~n32413 & ~n32447;
  assign n2050 = ~n1561 & n2049;
  assign n2051 = ~n1580 & n2050;
  assign n2052 = ~n32415 & n2051;
  assign n2053 = n1566 & n1582;
  assign n2054 = ~n1574 & n2052;
  assign n2055 = ~n2041 & ~n32477;
  assign n2056 = ~n1810 & n2055;
  assign n2057 = ~n32446 & n2056;
  assign n2058 = ~n1804 & n2057;
  assign n2059 = n1812 & n2042;
  assign n2060 = ~n2039 & n2058;
  assign n2061 = n2048 & ~n32478;
  assign n2062 = ~n2043 & ~n2061;
  assign n2063 = ~n1582 & ~n2062;
  assign n2064 = n1582 & ~n2043;
  assign n2065 = ~n2061 & n2064;
  assign n2066 = ~n1812 & ~n2036;
  assign n2067 = ~n32475 & n2066;
  assign n2068 = ~n2030 & n2067;
  assign n2069 = ~n32476 & ~n2068;
  assign n2070 = pi98  & ~n2069;
  assign n2071 = ~pi98  & ~n2068;
  assign n2072 = ~pi98  & n2069;
  assign n2073 = ~n32476 & n2071;
  assign n2074 = ~n2070 & ~n32479;
  assign n2075 = ~n2065 & ~n2074;
  assign n2076 = ~n2063 & ~n2075;
  assign n2077 = ~n1388 & ~n2076;
  assign n2078 = n1388 & ~n2063;
  assign n2079 = ~n2075 & n2078;
  assign n2080 = n1388 & n2076;
  assign n2081 = ~n1817 & ~n32448;
  assign n2082 = ~n2038 & n2081;
  assign n2083 = n1834 & ~n2082;
  assign n2084 = ~n1834 & n2081;
  assign n2085 = ~n1834 & n2082;
  assign n2086 = ~n2038 & n2084;
  assign n2087 = ~n2083 & ~n32481;
  assign n2088 = ~n32480 & ~n2087;
  assign n2089 = ~n2077 & ~n2088;
  assign n2090 = ~n1192 & ~n2089;
  assign n2091 = n1192 & ~n2077;
  assign n2092 = ~n2088 & n2091;
  assign n2093 = ~n1837 & ~n32451;
  assign n2094 = ~n1837 & ~n2038;
  assign n2095 = ~n32451 & n2094;
  assign n2096 = ~n2038 & n2093;
  assign n2097 = n1846 & ~n32482;
  assign n2098 = n1850 & n2094;
  assign n2099 = n1846 & ~n32451;
  assign n2100 = ~n1837 & n2099;
  assign n2101 = ~n2038 & n2100;
  assign n2102 = ~n1846 & ~n32482;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = ~n2097 & ~n2098;
  assign n2105 = ~n2092 & ~n32483;
  assign n2106 = ~n2090 & ~n2105;
  assign n2107 = ~n1028 & ~n2106;
  assign n2108 = n1028 & ~n2090;
  assign n2109 = ~n2105 & n2108;
  assign n2110 = n1028 & n2106;
  assign n2111 = ~n1852 & ~n1854;
  assign n2112 = ~n2038 & n2111;
  assign n2113 = n1861 & ~n2112;
  assign n2114 = ~n1861 & n2112;
  assign n2115 = ~n1852 & n1861;
  assign n2116 = ~n1854 & n2115;
  assign n2117 = n1861 & n2112;
  assign n2118 = ~n2038 & n2116;
  assign n2119 = ~n1861 & ~n2112;
  assign n2120 = ~n32485 & ~n2119;
  assign n2121 = ~n2113 & ~n2114;
  assign n2122 = ~n32484 & ~n32486;
  assign n2123 = ~n2107 & ~n2122;
  assign n2124 = ~n866 & ~n2123;
  assign n2125 = n866 & ~n2107;
  assign n2126 = ~n2122 & n2125;
  assign n2127 = ~n1864 & ~n32454;
  assign n2128 = ~n1864 & ~n2038;
  assign n2129 = ~n32454 & n2128;
  assign n2130 = ~n2038 & n2127;
  assign n2131 = n1872 & ~n32487;
  assign n2132 = n1876 & n2128;
  assign n2133 = n1872 & ~n32454;
  assign n2134 = ~n1864 & n2133;
  assign n2135 = ~n2038 & n2134;
  assign n2136 = ~n1872 & ~n32487;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = ~n2131 & ~n2132;
  assign n2139 = ~n2126 & ~n32488;
  assign n2140 = ~n2124 & ~n2139;
  assign n2141 = ~n730 & ~n2140;
  assign n2142 = n730 & ~n2124;
  assign n2143 = ~n2139 & n2142;
  assign n2144 = n730 & n2140;
  assign n2145 = ~n1878 & ~n1880;
  assign n2146 = ~n2038 & n2145;
  assign n2147 = ~n32456 & n2146;
  assign n2148 = n32456 & ~n2146;
  assign n2149 = ~n1878 & n32456;
  assign n2150 = ~n1880 & n2149;
  assign n2151 = ~n2038 & n2150;
  assign n2152 = ~n32456 & ~n2146;
  assign n2153 = ~n2151 & ~n2152;
  assign n2154 = ~n2147 & ~n2148;
  assign n2155 = ~n32489 & ~n32490;
  assign n2156 = ~n2141 & ~n2155;
  assign n2157 = ~n602 & ~n2156;
  assign n2158 = n602 & ~n2141;
  assign n2159 = ~n2155 & n2158;
  assign n2160 = ~n1894 & ~n32458;
  assign n2161 = ~n1894 & ~n2038;
  assign n2162 = ~n32458 & n2161;
  assign n2163 = ~n2038 & n2160;
  assign n2164 = n1902 & ~n32491;
  assign n2165 = n1906 & n2161;
  assign n2166 = n1902 & ~n32458;
  assign n2167 = ~n1894 & n2166;
  assign n2168 = ~n2038 & n2167;
  assign n2169 = ~n1902 & ~n32491;
  assign n2170 = ~n2168 & ~n2169;
  assign n2171 = ~n2164 & ~n2165;
  assign n2172 = ~n2159 & ~n32492;
  assign n2173 = ~n2157 & ~n2172;
  assign n2174 = ~n497 & ~n2173;
  assign n2175 = n497 & ~n2157;
  assign n2176 = ~n2172 & n2175;
  assign n2177 = n497 & n2173;
  assign n2178 = ~n1908 & ~n1910;
  assign n2179 = ~n2038 & n2178;
  assign n2180 = ~n32459 & ~n2179;
  assign n2181 = ~n1908 & n32459;
  assign n2182 = ~n1910 & n2181;
  assign n2183 = n32459 & n2179;
  assign n2184 = ~n2038 & n2182;
  assign n2185 = n32459 & ~n2179;
  assign n2186 = ~n32459 & n2179;
  assign n2187 = ~n2185 & ~n2186;
  assign n2188 = ~n2180 & ~n32494;
  assign n2189 = ~n32493 & n32495;
  assign n2190 = ~n2174 & ~n2189;
  assign n2191 = ~n403 & ~n2190;
  assign n2192 = n403 & ~n2174;
  assign n2193 = ~n2189 & n2192;
  assign n2194 = ~n1923 & ~n32461;
  assign n2195 = ~n1923 & ~n2038;
  assign n2196 = ~n32461 & n2195;
  assign n2197 = ~n2038 & n2194;
  assign n2198 = n1931 & ~n32496;
  assign n2199 = n1935 & n2195;
  assign n2200 = n1931 & ~n32461;
  assign n2201 = ~n1923 & n2200;
  assign n2202 = ~n2038 & n2201;
  assign n2203 = ~n1931 & ~n32496;
  assign n2204 = ~n2202 & ~n2203;
  assign n2205 = ~n2198 & ~n2199;
  assign n2206 = ~n2193 & ~n32497;
  assign n2207 = ~n2191 & ~n2206;
  assign n2208 = ~n330 & ~n2207;
  assign n2209 = n330 & ~n2191;
  assign n2210 = ~n2206 & n2209;
  assign n2211 = n330 & n2207;
  assign n2212 = ~n1937 & ~n1939;
  assign n2213 = ~n2038 & n2212;
  assign n2214 = n32463 & ~n2213;
  assign n2215 = ~n1937 & ~n32463;
  assign n2216 = ~n1939 & n2215;
  assign n2217 = ~n32463 & n2213;
  assign n2218 = ~n2038 & n2216;
  assign n2219 = n32463 & n2213;
  assign n2220 = ~n32463 & ~n2213;
  assign n2221 = ~n2219 & ~n2220;
  assign n2222 = ~n2214 & ~n32499;
  assign n2223 = ~n32498 & n32500;
  assign n2224 = ~n2208 & ~n2223;
  assign n2225 = ~n271 & ~n2224;
  assign n2226 = n271 & ~n2208;
  assign n2227 = ~n2223 & n2226;
  assign n2228 = ~n1953 & ~n32465;
  assign n2229 = ~n1953 & ~n2038;
  assign n2230 = ~n32465 & n2229;
  assign n2231 = ~n2038 & n2228;
  assign n2232 = n1961 & ~n32501;
  assign n2233 = n1965 & n2229;
  assign n2234 = n1961 & ~n32465;
  assign n2235 = ~n1953 & n2234;
  assign n2236 = ~n2038 & n2235;
  assign n2237 = ~n1961 & ~n32501;
  assign n2238 = ~n2236 & ~n2237;
  assign n2239 = ~n2232 & ~n2233;
  assign n2240 = ~n2227 & ~n32502;
  assign n2241 = ~n2225 & ~n2240;
  assign n2242 = ~n217 & ~n2241;
  assign n2243 = n217 & ~n2225;
  assign n2244 = ~n2240 & n2243;
  assign n2245 = n217 & n2241;
  assign n2246 = ~n1967 & ~n1969;
  assign n2247 = ~n1967 & ~n2038;
  assign n2248 = ~n1969 & n2247;
  assign n2249 = ~n2038 & n2246;
  assign n2250 = ~n32467 & ~n32504;
  assign n2251 = n1981 & n2247;
  assign n2252 = n32467 & n32504;
  assign n2253 = ~n1967 & ~n32467;
  assign n2254 = ~n1969 & n2253;
  assign n2255 = ~n2038 & n2254;
  assign n2256 = n32467 & ~n32504;
  assign n2257 = ~n2255 & ~n2256;
  assign n2258 = ~n2250 & ~n32505;
  assign n2259 = ~n32503 & ~n32506;
  assign n2260 = ~n2242 & ~n2259;
  assign n2261 = ~n198 & ~n2260;
  assign n2262 = n198 & ~n2242;
  assign n2263 = ~n2259 & n2262;
  assign n2264 = ~n1983 & ~n32469;
  assign n2265 = ~n1983 & ~n2038;
  assign n2266 = ~n32469 & n2265;
  assign n2267 = ~n2038 & n2264;
  assign n2268 = n1991 & ~n32507;
  assign n2269 = n1995 & n2265;
  assign n2270 = n1991 & ~n32469;
  assign n2271 = ~n1983 & n2270;
  assign n2272 = ~n2038 & n2271;
  assign n2273 = ~n1991 & ~n32507;
  assign n2274 = ~n2272 & ~n2273;
  assign n2275 = ~n2268 & ~n2269;
  assign n2276 = ~n2263 & ~n32508;
  assign n2277 = ~n2261 & ~n2276;
  assign n2278 = ~n1997 & ~n1999;
  assign n2279 = ~n2038 & n2278;
  assign n2280 = ~n32472 & ~n2279;
  assign n2281 = ~n1997 & n32472;
  assign n2282 = ~n1999 & n2281;
  assign n2283 = n32472 & n2279;
  assign n2284 = ~n2038 & n2282;
  assign n2285 = ~n2280 & ~n32509;
  assign n2286 = ~n2014 & ~n2022;
  assign n2287 = ~n2022 & ~n2038;
  assign n2288 = ~n2014 & n2287;
  assign n2289 = ~n2038 & n2286;
  assign n2290 = ~n32475 & ~n32510;
  assign n2291 = ~n2285 & n2290;
  assign n2292 = ~n2277 & n2291;
  assign n2293 = n193 & ~n2292;
  assign n2294 = ~n2261 & n2285;
  assign n2295 = ~n2276 & n2294;
  assign n2296 = n2277 & n2285;
  assign n2297 = n2014 & ~n2287;
  assign n2298 = ~n193 & ~n2286;
  assign n2299 = ~n2297 & n2298;
  assign n2300 = ~n32511 & ~n2299;
  assign n2301 = ~n2293 & n2300;
  assign n2302 = pi94  & ~n2301;
  assign n2303 = ~pi92  & ~pi93 ;
  assign n2304 = ~pi94  & n2303;
  assign n2305 = ~n2302 & ~n2304;
  assign n2306 = ~n2038 & ~n2305;
  assign n2307 = ~n32443 & ~n32477;
  assign n2308 = ~n1794 & n2307;
  assign n2309 = ~n1810 & n2308;
  assign n2310 = ~n32446 & n2309;
  assign n2311 = n32444 & n1812;
  assign n2312 = ~n1804 & n2310;
  assign n2313 = ~n2304 & ~n32512;
  assign n2314 = ~n2036 & n2313;
  assign n2315 = ~n32475 & n2314;
  assign n2316 = ~n2030 & n2315;
  assign n2317 = n2038 & n2305;
  assign n2318 = ~n2302 & n2316;
  assign n2319 = ~pi94  & ~n2301;
  assign n2320 = pi95  & ~n2319;
  assign n2321 = ~pi95  & n2319;
  assign n2322 = n2040 & ~n2301;
  assign n2323 = ~n2320 & ~n32514;
  assign n2324 = ~n32513 & n2323;
  assign n2325 = ~n2306 & ~n2324;
  assign n2326 = ~n1812 & ~n2325;
  assign n2327 = ~n2038 & ~n2299;
  assign n2328 = ~n32511 & n2327;
  assign n2329 = ~n2293 & n2328;
  assign n2330 = ~n32514 & ~n2329;
  assign n2331 = pi96  & ~n2330;
  assign n2332 = ~pi96  & ~n2329;
  assign n2333 = ~pi96  & n2330;
  assign n2334 = ~n32514 & n2332;
  assign n2335 = ~n2331 & ~n32515;
  assign n2336 = n1812 & ~n2306;
  assign n2337 = n1812 & n2325;
  assign n2338 = ~n2324 & n2336;
  assign n2339 = ~n2335 & ~n32516;
  assign n2340 = ~n2326 & ~n2339;
  assign n2341 = ~n1582 & ~n2340;
  assign n2342 = n1582 & ~n2326;
  assign n2343 = ~n2339 & n2342;
  assign n2344 = ~n2043 & ~n32478;
  assign n2345 = ~n2301 & n2344;
  assign n2346 = n2048 & ~n2345;
  assign n2347 = ~n2048 & ~n32478;
  assign n2348 = ~n2043 & n2347;
  assign n2349 = ~n2048 & n2344;
  assign n2350 = ~n2048 & n2345;
  assign n2351 = ~n2301 & n32517;
  assign n2352 = ~n2346 & ~n32518;
  assign n2353 = ~n2343 & ~n2352;
  assign n2354 = ~n2341 & ~n2353;
  assign n2355 = ~n1388 & ~n2354;
  assign n2356 = ~n2063 & ~n2065;
  assign n2357 = ~n2301 & n2356;
  assign n2358 = ~n2074 & ~n2357;
  assign n2359 = ~n2065 & n2074;
  assign n2360 = ~n2063 & n2359;
  assign n2361 = n2074 & n2357;
  assign n2362 = ~n2301 & n2360;
  assign n2363 = ~n2358 & ~n32519;
  assign n2364 = n1388 & ~n2341;
  assign n2365 = n1388 & n2354;
  assign n2366 = ~n2353 & n2364;
  assign n2367 = ~n2363 & ~n32520;
  assign n2368 = ~n2355 & ~n2367;
  assign n2369 = ~n1192 & ~n2368;
  assign n2370 = n1192 & ~n2355;
  assign n2371 = ~n2367 & n2370;
  assign n2372 = ~n2077 & ~n32480;
  assign n2373 = ~n2301 & n2372;
  assign n2374 = n2087 & ~n2373;
  assign n2375 = ~n2087 & n2373;
  assign n2376 = ~n2077 & n2087;
  assign n2377 = ~n32480 & n2376;
  assign n2378 = n2087 & n2373;
  assign n2379 = ~n2301 & n2377;
  assign n2380 = ~n2087 & ~n2373;
  assign n2381 = ~n32521 & ~n2380;
  assign n2382 = ~n2374 & ~n2375;
  assign n2383 = ~n2371 & ~n32522;
  assign n2384 = ~n2369 & ~n2383;
  assign n2385 = ~n1028 & ~n2384;
  assign n2386 = ~n2090 & ~n2092;
  assign n2387 = ~n2301 & n2386;
  assign n2388 = ~n32483 & ~n2387;
  assign n2389 = ~n2092 & n32483;
  assign n2390 = ~n2090 & n2389;
  assign n2391 = n32483 & n2387;
  assign n2392 = ~n2301 & n2390;
  assign n2393 = ~n2388 & ~n32523;
  assign n2394 = n1028 & ~n2369;
  assign n2395 = n1028 & n2384;
  assign n2396 = ~n2383 & n2394;
  assign n2397 = ~n2393 & ~n32524;
  assign n2398 = ~n2385 & ~n2397;
  assign n2399 = ~n866 & ~n2398;
  assign n2400 = n866 & ~n2385;
  assign n2401 = ~n2397 & n2400;
  assign n2402 = ~n2107 & ~n32484;
  assign n2403 = ~n2301 & n2402;
  assign n2404 = ~n32486 & n2403;
  assign n2405 = n32486 & ~n2403;
  assign n2406 = ~n2107 & n32486;
  assign n2407 = ~n32484 & n2406;
  assign n2408 = ~n2301 & n2407;
  assign n2409 = ~n32486 & ~n2403;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = ~n2404 & ~n2405;
  assign n2412 = ~n2401 & ~n32525;
  assign n2413 = ~n2399 & ~n2412;
  assign n2414 = ~n730 & ~n2413;
  assign n2415 = ~n2124 & ~n2126;
  assign n2416 = ~n2301 & n2415;
  assign n2417 = ~n32488 & ~n2416;
  assign n2418 = ~n2126 & n32488;
  assign n2419 = ~n2124 & n2418;
  assign n2420 = n32488 & n2416;
  assign n2421 = ~n2301 & n2419;
  assign n2422 = ~n2417 & ~n32526;
  assign n2423 = n730 & ~n2399;
  assign n2424 = n730 & n2413;
  assign n2425 = ~n2412 & n2423;
  assign n2426 = ~n2422 & ~n32527;
  assign n2427 = ~n2414 & ~n2426;
  assign n2428 = ~n602 & ~n2427;
  assign n2429 = n602 & ~n2414;
  assign n2430 = ~n2426 & n2429;
  assign n2431 = ~n2141 & ~n32489;
  assign n2432 = ~n2301 & n2431;
  assign n2433 = ~n32490 & ~n2432;
  assign n2434 = ~n2141 & n32490;
  assign n2435 = ~n32489 & n2434;
  assign n2436 = n32490 & n2432;
  assign n2437 = ~n2301 & n2435;
  assign n2438 = n32490 & ~n2432;
  assign n2439 = ~n32490 & n2432;
  assign n2440 = ~n2438 & ~n2439;
  assign n2441 = ~n2433 & ~n32528;
  assign n2442 = ~n2430 & n32529;
  assign n2443 = ~n2428 & ~n2442;
  assign n2444 = ~n497 & ~n2443;
  assign n2445 = ~n2157 & ~n2159;
  assign n2446 = ~n2301 & n2445;
  assign n2447 = ~n32492 & ~n2446;
  assign n2448 = ~n2159 & n32492;
  assign n2449 = ~n2157 & n2448;
  assign n2450 = n32492 & n2446;
  assign n2451 = ~n2301 & n2449;
  assign n2452 = ~n2447 & ~n32530;
  assign n2453 = n497 & ~n2428;
  assign n2454 = n497 & n2443;
  assign n2455 = ~n2442 & n2453;
  assign n2456 = ~n2452 & ~n32531;
  assign n2457 = ~n2444 & ~n2456;
  assign n2458 = ~n403 & ~n2457;
  assign n2459 = n403 & ~n2444;
  assign n2460 = ~n2456 & n2459;
  assign n2461 = ~n2174 & ~n32493;
  assign n2462 = ~n2301 & n2461;
  assign n2463 = n32495 & ~n2462;
  assign n2464 = ~n2174 & ~n32495;
  assign n2465 = ~n32493 & n2464;
  assign n2466 = ~n32495 & n2462;
  assign n2467 = ~n2301 & n2465;
  assign n2468 = n32495 & n2462;
  assign n2469 = ~n32495 & ~n2462;
  assign n2470 = ~n2468 & ~n2469;
  assign n2471 = ~n2463 & ~n32532;
  assign n2472 = ~n2460 & n32533;
  assign n2473 = ~n2458 & ~n2472;
  assign n2474 = ~n330 & ~n2473;
  assign n2475 = ~n2191 & ~n2193;
  assign n2476 = ~n2301 & n2475;
  assign n2477 = ~n32497 & ~n2476;
  assign n2478 = ~n2193 & n32497;
  assign n2479 = ~n2191 & n2478;
  assign n2480 = n32497 & n2476;
  assign n2481 = ~n2301 & n2479;
  assign n2482 = ~n2477 & ~n32534;
  assign n2483 = n330 & ~n2458;
  assign n2484 = n330 & n2473;
  assign n2485 = ~n2472 & n2483;
  assign n2486 = ~n2482 & ~n32535;
  assign n2487 = ~n2474 & ~n2486;
  assign n2488 = ~n271 & ~n2487;
  assign n2489 = n271 & ~n2474;
  assign n2490 = ~n2486 & n2489;
  assign n2491 = ~n2208 & ~n32498;
  assign n2492 = ~n2208 & ~n2301;
  assign n2493 = ~n32498 & n2492;
  assign n2494 = ~n2301 & n2491;
  assign n2495 = ~n32500 & ~n32536;
  assign n2496 = n2223 & n2492;
  assign n2497 = n32500 & n32536;
  assign n2498 = ~n2208 & ~n32500;
  assign n2499 = ~n32498 & n2498;
  assign n2500 = ~n2301 & n2499;
  assign n2501 = n32500 & ~n32536;
  assign n2502 = ~n2500 & ~n2501;
  assign n2503 = ~n2495 & ~n32537;
  assign n2504 = ~n2490 & ~n32538;
  assign n2505 = ~n2488 & ~n2504;
  assign n2506 = ~n217 & ~n2505;
  assign n2507 = ~n2225 & ~n2227;
  assign n2508 = ~n2301 & n2507;
  assign n2509 = ~n32502 & ~n2508;
  assign n2510 = ~n2227 & n32502;
  assign n2511 = ~n2225 & n2510;
  assign n2512 = n32502 & n2508;
  assign n2513 = ~n2301 & n2511;
  assign n2514 = ~n2509 & ~n32539;
  assign n2515 = n217 & ~n2488;
  assign n2516 = n217 & n2505;
  assign n2517 = ~n2504 & n2515;
  assign n2518 = ~n2514 & ~n32540;
  assign n2519 = ~n2506 & ~n2518;
  assign n2520 = ~n198 & ~n2519;
  assign n2521 = n198 & ~n2506;
  assign n2522 = ~n2518 & n2521;
  assign n2523 = ~n2242 & ~n32503;
  assign n2524 = ~n2301 & n2523;
  assign n2525 = ~n32506 & ~n2524;
  assign n2526 = ~n2242 & n32506;
  assign n2527 = ~n32503 & n2526;
  assign n2528 = n32506 & n2524;
  assign n2529 = ~n2301 & n2527;
  assign n2530 = ~n2525 & ~n32541;
  assign n2531 = ~n2522 & ~n2530;
  assign n2532 = ~n2520 & ~n2531;
  assign n2533 = ~n2261 & ~n2263;
  assign n2534 = ~n2301 & n2533;
  assign n2535 = ~n32508 & ~n2534;
  assign n2536 = ~n2263 & n32508;
  assign n2537 = ~n2261 & n2536;
  assign n2538 = n32508 & n2534;
  assign n2539 = ~n2301 & n2537;
  assign n2540 = ~n2535 & ~n32542;
  assign n2541 = ~n2277 & ~n2285;
  assign n2542 = ~n2285 & ~n2301;
  assign n2543 = ~n2277 & n2542;
  assign n2544 = ~n2301 & n2541;
  assign n2545 = ~n32511 & ~n32543;
  assign n2546 = ~n2540 & n2545;
  assign n2547 = ~n2532 & n2546;
  assign n2548 = n193 & ~n2547;
  assign n2549 = ~n2520 & n2540;
  assign n2550 = n2532 & n2540;
  assign n2551 = ~n2531 & n2549;
  assign n2552 = n2277 & ~n2542;
  assign n2553 = ~n193 & ~n2541;
  assign n2554 = ~n2552 & n2553;
  assign n2555 = ~n32544 & ~n2554;
  assign n2556 = ~n2548 & n2555;
  assign n2557 = pi92  & ~n2556;
  assign n2558 = ~pi90  & ~pi91 ;
  assign n2559 = ~pi92  & n2558;
  assign n2560 = ~n2557 & ~n2559;
  assign n2561 = ~n2301 & ~n2560;
  assign n2562 = ~pi92  & ~n2556;
  assign n2563 = pi93  & ~n2562;
  assign n2564 = ~pi93  & n2562;
  assign n2565 = n2303 & ~n2556;
  assign n2566 = ~n2563 & ~n32545;
  assign n2567 = ~n32473 & ~n32512;
  assign n2568 = ~n2017 & n2567;
  assign n2569 = ~n2036 & n2568;
  assign n2570 = ~n32475 & n2569;
  assign n2571 = n2022 & n2038;
  assign n2572 = ~n2030 & n2570;
  assign n2573 = ~n2559 & ~n32546;
  assign n2574 = ~n2299 & n2573;
  assign n2575 = ~n32511 & n2574;
  assign n2576 = ~n2293 & n2575;
  assign n2577 = n2301 & n2560;
  assign n2578 = ~n2557 & n2576;
  assign n2579 = n2566 & ~n32547;
  assign n2580 = ~n2561 & ~n2579;
  assign n2581 = ~n2038 & ~n2580;
  assign n2582 = n2038 & ~n2561;
  assign n2583 = ~n2579 & n2582;
  assign n2584 = ~n2301 & ~n2554;
  assign n2585 = ~n32544 & n2584;
  assign n2586 = ~n2548 & n2585;
  assign n2587 = ~n32545 & ~n2586;
  assign n2588 = pi94  & ~n2587;
  assign n2589 = ~pi94  & ~n2586;
  assign n2590 = ~pi94  & n2587;
  assign n2591 = ~n32545 & n2589;
  assign n2592 = ~n2588 & ~n32548;
  assign n2593 = ~n2583 & ~n2592;
  assign n2594 = ~n2581 & ~n2593;
  assign n2595 = ~n1812 & ~n2594;
  assign n2596 = n1812 & ~n2581;
  assign n2597 = ~n2593 & n2596;
  assign n2598 = n1812 & n2594;
  assign n2599 = ~n2306 & ~n32513;
  assign n2600 = ~n2556 & n2599;
  assign n2601 = n2323 & ~n2600;
  assign n2602 = ~n2323 & n2599;
  assign n2603 = ~n2323 & n2600;
  assign n2604 = ~n2556 & n2602;
  assign n2605 = ~n2601 & ~n32550;
  assign n2606 = ~n32549 & ~n2605;
  assign n2607 = ~n2595 & ~n2606;
  assign n2608 = ~n1582 & ~n2607;
  assign n2609 = n1582 & ~n2595;
  assign n2610 = ~n2606 & n2609;
  assign n2611 = ~n2326 & ~n32516;
  assign n2612 = ~n2326 & ~n2556;
  assign n2613 = ~n32516 & n2612;
  assign n2614 = ~n2556 & n2611;
  assign n2615 = n2335 & ~n32551;
  assign n2616 = n2339 & n2612;
  assign n2617 = n2335 & ~n32516;
  assign n2618 = ~n2326 & n2617;
  assign n2619 = ~n2556 & n2618;
  assign n2620 = ~n2335 & ~n32551;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = ~n2615 & ~n2616;
  assign n2623 = ~n2610 & ~n32552;
  assign n2624 = ~n2608 & ~n2623;
  assign n2625 = ~n1388 & ~n2624;
  assign n2626 = n1388 & ~n2608;
  assign n2627 = ~n2623 & n2626;
  assign n2628 = n1388 & n2624;
  assign n2629 = ~n2341 & ~n2343;
  assign n2630 = ~n2556 & n2629;
  assign n2631 = n2352 & ~n2630;
  assign n2632 = ~n2352 & n2630;
  assign n2633 = ~n2341 & n2352;
  assign n2634 = ~n2343 & n2633;
  assign n2635 = n2352 & n2630;
  assign n2636 = ~n2556 & n2634;
  assign n2637 = ~n2352 & ~n2630;
  assign n2638 = ~n32554 & ~n2637;
  assign n2639 = ~n2631 & ~n2632;
  assign n2640 = ~n32553 & ~n32555;
  assign n2641 = ~n2625 & ~n2640;
  assign n2642 = ~n1192 & ~n2641;
  assign n2643 = n1192 & ~n2625;
  assign n2644 = ~n2640 & n2643;
  assign n2645 = ~n2355 & ~n32520;
  assign n2646 = ~n2355 & ~n2556;
  assign n2647 = ~n32520 & n2646;
  assign n2648 = ~n2556 & n2645;
  assign n2649 = n2363 & ~n32556;
  assign n2650 = n2367 & n2646;
  assign n2651 = n2363 & ~n32520;
  assign n2652 = ~n2355 & n2651;
  assign n2653 = ~n2556 & n2652;
  assign n2654 = ~n2363 & ~n32556;
  assign n2655 = ~n2653 & ~n2654;
  assign n2656 = ~n2649 & ~n2650;
  assign n2657 = ~n2644 & ~n32557;
  assign n2658 = ~n2642 & ~n2657;
  assign n2659 = ~n1028 & ~n2658;
  assign n2660 = n1028 & ~n2642;
  assign n2661 = ~n2657 & n2660;
  assign n2662 = n1028 & n2658;
  assign n2663 = ~n2369 & ~n2371;
  assign n2664 = ~n2556 & n2663;
  assign n2665 = ~n32522 & n2664;
  assign n2666 = n32522 & ~n2664;
  assign n2667 = ~n2369 & n32522;
  assign n2668 = ~n2371 & n2667;
  assign n2669 = ~n2556 & n2668;
  assign n2670 = ~n32522 & ~n2664;
  assign n2671 = ~n2669 & ~n2670;
  assign n2672 = ~n2665 & ~n2666;
  assign n2673 = ~n32558 & ~n32559;
  assign n2674 = ~n2659 & ~n2673;
  assign n2675 = ~n866 & ~n2674;
  assign n2676 = n866 & ~n2659;
  assign n2677 = ~n2673 & n2676;
  assign n2678 = ~n2385 & ~n32524;
  assign n2679 = ~n2385 & ~n2556;
  assign n2680 = ~n32524 & n2679;
  assign n2681 = ~n2556 & n2678;
  assign n2682 = n2393 & ~n32560;
  assign n2683 = n2397 & n2679;
  assign n2684 = n2393 & ~n32524;
  assign n2685 = ~n2385 & n2684;
  assign n2686 = ~n2556 & n2685;
  assign n2687 = ~n2393 & ~n32560;
  assign n2688 = ~n2686 & ~n2687;
  assign n2689 = ~n2682 & ~n2683;
  assign n2690 = ~n2677 & ~n32561;
  assign n2691 = ~n2675 & ~n2690;
  assign n2692 = ~n730 & ~n2691;
  assign n2693 = n730 & ~n2675;
  assign n2694 = ~n2690 & n2693;
  assign n2695 = n730 & n2691;
  assign n2696 = ~n2399 & ~n2401;
  assign n2697 = ~n2556 & n2696;
  assign n2698 = ~n32525 & ~n2697;
  assign n2699 = ~n2399 & n32525;
  assign n2700 = ~n2401 & n2699;
  assign n2701 = n32525 & n2697;
  assign n2702 = ~n2556 & n2700;
  assign n2703 = n32525 & ~n2697;
  assign n2704 = ~n32525 & n2697;
  assign n2705 = ~n2703 & ~n2704;
  assign n2706 = ~n2698 & ~n32563;
  assign n2707 = ~n32562 & n32564;
  assign n2708 = ~n2692 & ~n2707;
  assign n2709 = ~n602 & ~n2708;
  assign n2710 = n602 & ~n2692;
  assign n2711 = ~n2707 & n2710;
  assign n2712 = ~n2414 & ~n32527;
  assign n2713 = ~n2414 & ~n2556;
  assign n2714 = ~n32527 & n2713;
  assign n2715 = ~n2556 & n2712;
  assign n2716 = n2422 & ~n32565;
  assign n2717 = n2426 & n2713;
  assign n2718 = n2422 & ~n32527;
  assign n2719 = ~n2414 & n2718;
  assign n2720 = ~n2556 & n2719;
  assign n2721 = ~n2422 & ~n32565;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = ~n2716 & ~n2717;
  assign n2724 = ~n2711 & ~n32566;
  assign n2725 = ~n2709 & ~n2724;
  assign n2726 = ~n497 & ~n2725;
  assign n2727 = n497 & ~n2709;
  assign n2728 = ~n2724 & n2727;
  assign n2729 = n497 & n2725;
  assign n2730 = ~n2428 & ~n2430;
  assign n2731 = ~n2556 & n2730;
  assign n2732 = n32529 & ~n2731;
  assign n2733 = ~n2428 & ~n32529;
  assign n2734 = ~n2430 & n2733;
  assign n2735 = ~n32529 & n2731;
  assign n2736 = ~n2556 & n2734;
  assign n2737 = n32529 & n2731;
  assign n2738 = ~n32529 & ~n2731;
  assign n2739 = ~n2737 & ~n2738;
  assign n2740 = ~n2732 & ~n32568;
  assign n2741 = ~n32567 & n32569;
  assign n2742 = ~n2726 & ~n2741;
  assign n2743 = ~n403 & ~n2742;
  assign n2744 = n403 & ~n2726;
  assign n2745 = ~n2741 & n2744;
  assign n2746 = ~n2444 & ~n32531;
  assign n2747 = ~n2444 & ~n2556;
  assign n2748 = ~n32531 & n2747;
  assign n2749 = ~n2556 & n2746;
  assign n2750 = n2452 & ~n32570;
  assign n2751 = n2456 & n2747;
  assign n2752 = n2452 & ~n32531;
  assign n2753 = ~n2444 & n2752;
  assign n2754 = ~n2556 & n2753;
  assign n2755 = ~n2452 & ~n32570;
  assign n2756 = ~n2754 & ~n2755;
  assign n2757 = ~n2750 & ~n2751;
  assign n2758 = ~n2745 & ~n32571;
  assign n2759 = ~n2743 & ~n2758;
  assign n2760 = ~n330 & ~n2759;
  assign n2761 = n330 & ~n2743;
  assign n2762 = ~n2758 & n2761;
  assign n2763 = n330 & n2759;
  assign n2764 = ~n2458 & ~n2460;
  assign n2765 = ~n2458 & ~n2556;
  assign n2766 = ~n2460 & n2765;
  assign n2767 = ~n2556 & n2764;
  assign n2768 = ~n32533 & ~n32573;
  assign n2769 = n2472 & n2765;
  assign n2770 = n32533 & n32573;
  assign n2771 = ~n2458 & ~n32533;
  assign n2772 = ~n2460 & n2771;
  assign n2773 = ~n2556 & n2772;
  assign n2774 = n32533 & ~n32573;
  assign n2775 = ~n2773 & ~n2774;
  assign n2776 = ~n2768 & ~n32574;
  assign n2777 = ~n32572 & ~n32575;
  assign n2778 = ~n2760 & ~n2777;
  assign n2779 = ~n271 & ~n2778;
  assign n2780 = n271 & ~n2760;
  assign n2781 = ~n2777 & n2780;
  assign n2782 = ~n2474 & ~n32535;
  assign n2783 = ~n2474 & ~n2556;
  assign n2784 = ~n32535 & n2783;
  assign n2785 = ~n2556 & n2782;
  assign n2786 = n2482 & ~n32576;
  assign n2787 = n2486 & n2783;
  assign n2788 = n2482 & ~n32535;
  assign n2789 = ~n2474 & n2788;
  assign n2790 = ~n2556 & n2789;
  assign n2791 = ~n2482 & ~n32576;
  assign n2792 = ~n2790 & ~n2791;
  assign n2793 = ~n2786 & ~n2787;
  assign n2794 = ~n2781 & ~n32577;
  assign n2795 = ~n2779 & ~n2794;
  assign n2796 = ~n217 & ~n2795;
  assign n2797 = n217 & ~n2779;
  assign n2798 = ~n2794 & n2797;
  assign n2799 = n217 & n2795;
  assign n2800 = ~n2488 & ~n2490;
  assign n2801 = ~n2556 & n2800;
  assign n2802 = ~n32538 & ~n2801;
  assign n2803 = ~n2488 & n32538;
  assign n2804 = ~n2490 & n2803;
  assign n2805 = n32538 & n2801;
  assign n2806 = ~n2556 & n2804;
  assign n2807 = ~n2802 & ~n32579;
  assign n2808 = ~n32578 & ~n2807;
  assign n2809 = ~n2796 & ~n2808;
  assign n2810 = ~n198 & ~n2809;
  assign n2811 = n198 & ~n2796;
  assign n2812 = ~n2808 & n2811;
  assign n2813 = ~n2506 & ~n32540;
  assign n2814 = ~n2506 & ~n2556;
  assign n2815 = ~n32540 & n2814;
  assign n2816 = ~n2556 & n2813;
  assign n2817 = n2514 & ~n32580;
  assign n2818 = n2518 & n2814;
  assign n2819 = n2514 & ~n32540;
  assign n2820 = ~n2506 & n2819;
  assign n2821 = ~n2556 & n2820;
  assign n2822 = ~n2514 & ~n32580;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = ~n2817 & ~n2818;
  assign n2825 = ~n2812 & ~n32581;
  assign n2826 = ~n2810 & ~n2825;
  assign n2827 = ~n2520 & ~n2522;
  assign n2828 = ~n2520 & ~n2556;
  assign n2829 = ~n2522 & n2828;
  assign n2830 = ~n2556 & n2827;
  assign n2831 = n2530 & ~n32582;
  assign n2832 = n2531 & n2828;
  assign n2833 = ~n2530 & n32582;
  assign n2834 = ~n2520 & n2530;
  assign n2835 = ~n2522 & n2834;
  assign n2836 = ~n2556 & n2835;
  assign n2837 = ~n2530 & ~n32582;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = ~n2831 & ~n32583;
  assign n2840 = ~n2532 & ~n2540;
  assign n2841 = ~n2540 & ~n2556;
  assign n2842 = ~n2532 & n2841;
  assign n2843 = ~n2556 & n2840;
  assign n2844 = ~n32544 & ~n32585;
  assign n2845 = ~n32584 & n2844;
  assign n2846 = ~n2826 & n2845;
  assign n2847 = n193 & ~n2846;
  assign n2848 = ~n2810 & n32584;
  assign n2849 = ~n2825 & n2848;
  assign n2850 = n2826 & n32584;
  assign n2851 = n2532 & ~n2841;
  assign n2852 = ~n193 & ~n2840;
  assign n2853 = ~n2851 & n2852;
  assign n2854 = ~n32586 & ~n2853;
  assign n2855 = ~n2847 & n2854;
  assign n2856 = pi90  & ~n2855;
  assign n2857 = ~pi88  & ~pi89 ;
  assign n2858 = ~pi90  & n2857;
  assign n2859 = ~n2856 & ~n2858;
  assign n2860 = ~n2556 & ~n2859;
  assign n2861 = ~n32509 & ~n32546;
  assign n2862 = ~n2280 & n2861;
  assign n2863 = ~n2299 & n2862;
  assign n2864 = ~n32511 & n2863;
  assign n2865 = n2285 & n2301;
  assign n2866 = ~n2293 & n2864;
  assign n2867 = ~n2858 & ~n32587;
  assign n2868 = ~n2554 & n2867;
  assign n2869 = ~n32544 & n2868;
  assign n2870 = ~n2548 & n2869;
  assign n2871 = n2556 & n2859;
  assign n2872 = ~n2856 & n2870;
  assign n2873 = ~pi90  & ~n2855;
  assign n2874 = pi91  & ~n2873;
  assign n2875 = ~pi91  & n2873;
  assign n2876 = n2558 & ~n2855;
  assign n2877 = ~n2874 & ~n32589;
  assign n2878 = ~n32588 & n2877;
  assign n2879 = ~n2860 & ~n2878;
  assign n2880 = ~n2301 & ~n2879;
  assign n2881 = ~n2556 & ~n2853;
  assign n2882 = ~n32586 & n2881;
  assign n2883 = ~n2847 & n2882;
  assign n2884 = ~n32589 & ~n2883;
  assign n2885 = pi92  & ~n2884;
  assign n2886 = ~pi92  & ~n2883;
  assign n2887 = ~pi92  & n2884;
  assign n2888 = ~n32589 & n2886;
  assign n2889 = ~n2885 & ~n32590;
  assign n2890 = n2301 & ~n2860;
  assign n2891 = n2301 & n2879;
  assign n2892 = ~n2878 & n2890;
  assign n2893 = ~n2889 & ~n32591;
  assign n2894 = ~n2880 & ~n2893;
  assign n2895 = ~n2038 & ~n2894;
  assign n2896 = n2038 & ~n2880;
  assign n2897 = ~n2893 & n2896;
  assign n2898 = ~n2561 & ~n32547;
  assign n2899 = ~n2855 & n2898;
  assign n2900 = n2566 & ~n2899;
  assign n2901 = ~n2566 & n2898;
  assign n2902 = ~n2566 & n2899;
  assign n2903 = ~n2855 & n2901;
  assign n2904 = ~n2900 & ~n32592;
  assign n2905 = ~n2897 & ~n2904;
  assign n2906 = ~n2895 & ~n2905;
  assign n2907 = ~n1812 & ~n2906;
  assign n2908 = ~n2581 & ~n2583;
  assign n2909 = ~n2855 & n2908;
  assign n2910 = ~n2592 & ~n2909;
  assign n2911 = ~n2583 & n2592;
  assign n2912 = ~n2581 & n2911;
  assign n2913 = n2592 & n2909;
  assign n2914 = ~n2855 & n2912;
  assign n2915 = ~n2910 & ~n32593;
  assign n2916 = n1812 & ~n2895;
  assign n2917 = n1812 & n2906;
  assign n2918 = ~n2905 & n2916;
  assign n2919 = ~n2915 & ~n32594;
  assign n2920 = ~n2907 & ~n2919;
  assign n2921 = ~n1582 & ~n2920;
  assign n2922 = n1582 & ~n2907;
  assign n2923 = ~n2919 & n2922;
  assign n2924 = ~n2595 & ~n32549;
  assign n2925 = ~n2855 & n2924;
  assign n2926 = n2605 & ~n2925;
  assign n2927 = ~n2605 & n2925;
  assign n2928 = ~n2595 & n2605;
  assign n2929 = ~n32549 & n2928;
  assign n2930 = n2605 & n2925;
  assign n2931 = ~n2855 & n2929;
  assign n2932 = ~n2605 & ~n2925;
  assign n2933 = ~n32595 & ~n2932;
  assign n2934 = ~n2926 & ~n2927;
  assign n2935 = ~n2923 & ~n32596;
  assign n2936 = ~n2921 & ~n2935;
  assign n2937 = ~n1388 & ~n2936;
  assign n2938 = ~n2608 & ~n2610;
  assign n2939 = ~n2855 & n2938;
  assign n2940 = ~n32552 & ~n2939;
  assign n2941 = ~n2610 & n32552;
  assign n2942 = ~n2608 & n2941;
  assign n2943 = n32552 & n2939;
  assign n2944 = ~n2855 & n2942;
  assign n2945 = ~n2940 & ~n32597;
  assign n2946 = n1388 & ~n2921;
  assign n2947 = n1388 & n2936;
  assign n2948 = ~n2935 & n2946;
  assign n2949 = ~n2945 & ~n32598;
  assign n2950 = ~n2937 & ~n2949;
  assign n2951 = ~n1192 & ~n2950;
  assign n2952 = n1192 & ~n2937;
  assign n2953 = ~n2949 & n2952;
  assign n2954 = ~n2625 & ~n32553;
  assign n2955 = ~n2855 & n2954;
  assign n2956 = ~n32555 & n2955;
  assign n2957 = n32555 & ~n2955;
  assign n2958 = ~n2625 & n32555;
  assign n2959 = ~n32553 & n2958;
  assign n2960 = ~n2855 & n2959;
  assign n2961 = ~n32555 & ~n2955;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = ~n2956 & ~n2957;
  assign n2964 = ~n2953 & ~n32599;
  assign n2965 = ~n2951 & ~n2964;
  assign n2966 = ~n1028 & ~n2965;
  assign n2967 = ~n2642 & ~n2644;
  assign n2968 = ~n2855 & n2967;
  assign n2969 = ~n32557 & ~n2968;
  assign n2970 = ~n2644 & n32557;
  assign n2971 = ~n2642 & n2970;
  assign n2972 = n32557 & n2968;
  assign n2973 = ~n2855 & n2971;
  assign n2974 = ~n2969 & ~n32600;
  assign n2975 = n1028 & ~n2951;
  assign n2976 = n1028 & n2965;
  assign n2977 = ~n2964 & n2975;
  assign n2978 = ~n2974 & ~n32601;
  assign n2979 = ~n2966 & ~n2978;
  assign n2980 = ~n866 & ~n2979;
  assign n2981 = n866 & ~n2966;
  assign n2982 = ~n2978 & n2981;
  assign n2983 = ~n2659 & ~n32558;
  assign n2984 = ~n2855 & n2983;
  assign n2985 = ~n32559 & ~n2984;
  assign n2986 = ~n2659 & n32559;
  assign n2987 = ~n32558 & n2986;
  assign n2988 = n32559 & n2984;
  assign n2989 = ~n2855 & n2987;
  assign n2990 = n32559 & ~n2984;
  assign n2991 = ~n32559 & n2984;
  assign n2992 = ~n2990 & ~n2991;
  assign n2993 = ~n2985 & ~n32602;
  assign n2994 = ~n2982 & n32603;
  assign n2995 = ~n2980 & ~n2994;
  assign n2996 = ~n730 & ~n2995;
  assign n2997 = ~n2675 & ~n2677;
  assign n2998 = ~n2855 & n2997;
  assign n2999 = ~n32561 & ~n2998;
  assign n3000 = ~n2677 & n32561;
  assign n3001 = ~n2675 & n3000;
  assign n3002 = n32561 & n2998;
  assign n3003 = ~n2855 & n3001;
  assign n3004 = ~n2999 & ~n32604;
  assign n3005 = n730 & ~n2980;
  assign n3006 = n730 & n2995;
  assign n3007 = ~n2994 & n3005;
  assign n3008 = ~n3004 & ~n32605;
  assign n3009 = ~n2996 & ~n3008;
  assign n3010 = ~n602 & ~n3009;
  assign n3011 = n602 & ~n2996;
  assign n3012 = ~n3008 & n3011;
  assign n3013 = ~n2692 & ~n32562;
  assign n3014 = ~n2855 & n3013;
  assign n3015 = n32564 & ~n3014;
  assign n3016 = ~n2692 & ~n32564;
  assign n3017 = ~n32562 & n3016;
  assign n3018 = ~n32564 & n3014;
  assign n3019 = ~n2855 & n3017;
  assign n3020 = n32564 & n3014;
  assign n3021 = ~n32564 & ~n3014;
  assign n3022 = ~n3020 & ~n3021;
  assign n3023 = ~n3015 & ~n32606;
  assign n3024 = ~n3012 & n32607;
  assign n3025 = ~n3010 & ~n3024;
  assign n3026 = ~n497 & ~n3025;
  assign n3027 = ~n2709 & ~n2711;
  assign n3028 = ~n2855 & n3027;
  assign n3029 = ~n32566 & ~n3028;
  assign n3030 = ~n2711 & n32566;
  assign n3031 = ~n2709 & n3030;
  assign n3032 = n32566 & n3028;
  assign n3033 = ~n2855 & n3031;
  assign n3034 = ~n3029 & ~n32608;
  assign n3035 = n497 & ~n3010;
  assign n3036 = n497 & n3025;
  assign n3037 = ~n3024 & n3035;
  assign n3038 = ~n3034 & ~n32609;
  assign n3039 = ~n3026 & ~n3038;
  assign n3040 = ~n403 & ~n3039;
  assign n3041 = n403 & ~n3026;
  assign n3042 = ~n3038 & n3041;
  assign n3043 = ~n2726 & ~n32567;
  assign n3044 = ~n2726 & ~n2855;
  assign n3045 = ~n32567 & n3044;
  assign n3046 = ~n2855 & n3043;
  assign n3047 = ~n32569 & ~n32610;
  assign n3048 = n2741 & n3044;
  assign n3049 = n32569 & n32610;
  assign n3050 = ~n2726 & ~n32569;
  assign n3051 = ~n32567 & n3050;
  assign n3052 = ~n2855 & n3051;
  assign n3053 = n32569 & ~n32610;
  assign n3054 = ~n3052 & ~n3053;
  assign n3055 = ~n3047 & ~n32611;
  assign n3056 = ~n3042 & ~n32612;
  assign n3057 = ~n3040 & ~n3056;
  assign n3058 = ~n330 & ~n3057;
  assign n3059 = ~n2743 & ~n2745;
  assign n3060 = ~n2855 & n3059;
  assign n3061 = ~n32571 & ~n3060;
  assign n3062 = ~n2745 & n32571;
  assign n3063 = ~n2743 & n3062;
  assign n3064 = n32571 & n3060;
  assign n3065 = ~n2855 & n3063;
  assign n3066 = ~n3061 & ~n32613;
  assign n3067 = n330 & ~n3040;
  assign n3068 = n330 & n3057;
  assign n3069 = ~n3056 & n3067;
  assign n3070 = ~n3066 & ~n32614;
  assign n3071 = ~n3058 & ~n3070;
  assign n3072 = ~n271 & ~n3071;
  assign n3073 = n271 & ~n3058;
  assign n3074 = ~n3070 & n3073;
  assign n3075 = ~n2760 & ~n32572;
  assign n3076 = ~n2855 & n3075;
  assign n3077 = ~n32575 & ~n3076;
  assign n3078 = ~n2760 & n32575;
  assign n3079 = ~n32572 & n3078;
  assign n3080 = n32575 & n3076;
  assign n3081 = ~n2855 & n3079;
  assign n3082 = ~n3077 & ~n32615;
  assign n3083 = ~n3074 & ~n3082;
  assign n3084 = ~n3072 & ~n3083;
  assign n3085 = ~n217 & ~n3084;
  assign n3086 = ~n2779 & ~n2781;
  assign n3087 = ~n2855 & n3086;
  assign n3088 = ~n32577 & ~n3087;
  assign n3089 = ~n2781 & n32577;
  assign n3090 = ~n2779 & n3089;
  assign n3091 = n32577 & n3087;
  assign n3092 = ~n2855 & n3090;
  assign n3093 = ~n3088 & ~n32616;
  assign n3094 = n217 & ~n3072;
  assign n3095 = n217 & n3084;
  assign n3096 = ~n3083 & n3094;
  assign n3097 = ~n3093 & ~n32617;
  assign n3098 = ~n3085 & ~n3097;
  assign n3099 = ~n198 & ~n3098;
  assign n3100 = n198 & ~n3085;
  assign n3101 = ~n3097 & n3100;
  assign n3102 = ~n2796 & ~n32578;
  assign n3103 = ~n2796 & ~n2855;
  assign n3104 = ~n32578 & n3103;
  assign n3105 = ~n2855 & n3102;
  assign n3106 = n2807 & ~n32618;
  assign n3107 = n2808 & n3103;
  assign n3108 = ~n2807 & n32618;
  assign n3109 = ~n2796 & n2807;
  assign n3110 = ~n32578 & n3109;
  assign n3111 = ~n2855 & n3110;
  assign n3112 = ~n2807 & ~n32618;
  assign n3113 = ~n3111 & ~n3112;
  assign n3114 = ~n3106 & ~n32619;
  assign n3115 = ~n3101 & ~n32620;
  assign n3116 = ~n3099 & ~n3115;
  assign n3117 = ~n2810 & ~n2812;
  assign n3118 = ~n2855 & n3117;
  assign n3119 = ~n32581 & ~n3118;
  assign n3120 = ~n2812 & n32581;
  assign n3121 = ~n2810 & n3120;
  assign n3122 = n32581 & n3118;
  assign n3123 = ~n2855 & n3121;
  assign n3124 = ~n3119 & ~n32621;
  assign n3125 = ~n2826 & ~n32584;
  assign n3126 = ~n32584 & ~n2855;
  assign n3127 = ~n2826 & n3126;
  assign n3128 = ~n2855 & n3125;
  assign n3129 = ~n32586 & ~n32622;
  assign n3130 = ~n3124 & n3129;
  assign n3131 = ~n3116 & n3130;
  assign n3132 = n193 & ~n3131;
  assign n3133 = ~n3099 & n3124;
  assign n3134 = n3116 & n3124;
  assign n3135 = ~n3115 & n3133;
  assign n3136 = n2826 & ~n3126;
  assign n3137 = ~n193 & ~n3125;
  assign n3138 = ~n3136 & n3137;
  assign n3139 = ~n32623 & ~n3138;
  assign n3140 = ~n3132 & n3139;
  assign n3141 = pi88  & ~n3140;
  assign n3142 = ~pi86  & ~pi87 ;
  assign n3143 = ~pi88  & n3142;
  assign n3144 = ~n3141 & ~n3143;
  assign n3145 = ~n2855 & ~n3144;
  assign n3146 = ~pi88  & ~n3140;
  assign n3147 = pi89  & ~n3146;
  assign n3148 = ~pi89  & n3146;
  assign n3149 = n2857 & ~n3140;
  assign n3150 = ~n3147 & ~n32624;
  assign n3151 = ~n32542 & ~n32587;
  assign n3152 = ~n2535 & n3151;
  assign n3153 = ~n2554 & n3152;
  assign n3154 = ~n32544 & n3153;
  assign n3155 = n2540 & n2556;
  assign n3156 = ~n2548 & n3154;
  assign n3157 = ~n3143 & ~n32625;
  assign n3158 = ~n2853 & n3157;
  assign n3159 = ~n32586 & n3158;
  assign n3160 = ~n2847 & n3159;
  assign n3161 = n2855 & n3144;
  assign n3162 = ~n3141 & n3160;
  assign n3163 = n3150 & ~n32626;
  assign n3164 = ~n3145 & ~n3163;
  assign n3165 = ~n2556 & ~n3164;
  assign n3166 = n2556 & ~n3145;
  assign n3167 = ~n3163 & n3166;
  assign n3168 = ~n2855 & ~n3138;
  assign n3169 = ~n32623 & n3168;
  assign n3170 = ~n3132 & n3169;
  assign n3171 = ~n32624 & ~n3170;
  assign n3172 = pi90  & ~n3171;
  assign n3173 = ~pi90  & ~n3170;
  assign n3174 = ~pi90  & n3171;
  assign n3175 = ~n32624 & n3173;
  assign n3176 = ~n3172 & ~n32627;
  assign n3177 = ~n3167 & ~n3176;
  assign n3178 = ~n3165 & ~n3177;
  assign n3179 = ~n2301 & ~n3178;
  assign n3180 = n2301 & ~n3165;
  assign n3181 = ~n3177 & n3180;
  assign n3182 = n2301 & n3178;
  assign n3183 = ~n2860 & ~n32588;
  assign n3184 = ~n3140 & n3183;
  assign n3185 = n2877 & ~n3184;
  assign n3186 = ~n2877 & n3183;
  assign n3187 = ~n2877 & n3184;
  assign n3188 = ~n3140 & n3186;
  assign n3189 = ~n3185 & ~n32629;
  assign n3190 = ~n32628 & ~n3189;
  assign n3191 = ~n3179 & ~n3190;
  assign n3192 = ~n2038 & ~n3191;
  assign n3193 = n2038 & ~n3179;
  assign n3194 = ~n3190 & n3193;
  assign n3195 = ~n2880 & ~n32591;
  assign n3196 = ~n2880 & ~n3140;
  assign n3197 = ~n32591 & n3196;
  assign n3198 = ~n3140 & n3195;
  assign n3199 = n2889 & ~n32630;
  assign n3200 = n2893 & n3196;
  assign n3201 = n2889 & ~n32591;
  assign n3202 = ~n2880 & n3201;
  assign n3203 = ~n3140 & n3202;
  assign n3204 = ~n2889 & ~n32630;
  assign n3205 = ~n3203 & ~n3204;
  assign n3206 = ~n3199 & ~n3200;
  assign n3207 = ~n3194 & ~n32631;
  assign n3208 = ~n3192 & ~n3207;
  assign n3209 = ~n1812 & ~n3208;
  assign n3210 = n1812 & ~n3192;
  assign n3211 = ~n3207 & n3210;
  assign n3212 = n1812 & n3208;
  assign n3213 = ~n2895 & ~n2897;
  assign n3214 = ~n3140 & n3213;
  assign n3215 = n2904 & ~n3214;
  assign n3216 = ~n2904 & n3214;
  assign n3217 = ~n2895 & n2904;
  assign n3218 = ~n2897 & n3217;
  assign n3219 = n2904 & n3214;
  assign n3220 = ~n3140 & n3218;
  assign n3221 = ~n2904 & ~n3214;
  assign n3222 = ~n32633 & ~n3221;
  assign n3223 = ~n3215 & ~n3216;
  assign n3224 = ~n32632 & ~n32634;
  assign n3225 = ~n3209 & ~n3224;
  assign n3226 = ~n1582 & ~n3225;
  assign n3227 = n1582 & ~n3209;
  assign n3228 = ~n3224 & n3227;
  assign n3229 = ~n2907 & ~n32594;
  assign n3230 = ~n2907 & ~n3140;
  assign n3231 = ~n32594 & n3230;
  assign n3232 = ~n3140 & n3229;
  assign n3233 = n2915 & ~n32635;
  assign n3234 = n2919 & n3230;
  assign n3235 = n2915 & ~n32594;
  assign n3236 = ~n2907 & n3235;
  assign n3237 = ~n3140 & n3236;
  assign n3238 = ~n2915 & ~n32635;
  assign n3239 = ~n3237 & ~n3238;
  assign n3240 = ~n3233 & ~n3234;
  assign n3241 = ~n3228 & ~n32636;
  assign n3242 = ~n3226 & ~n3241;
  assign n3243 = ~n1388 & ~n3242;
  assign n3244 = n1388 & ~n3226;
  assign n3245 = ~n3241 & n3244;
  assign n3246 = n1388 & n3242;
  assign n3247 = ~n2921 & ~n2923;
  assign n3248 = ~n3140 & n3247;
  assign n3249 = ~n32596 & n3248;
  assign n3250 = n32596 & ~n3248;
  assign n3251 = ~n2921 & n32596;
  assign n3252 = ~n2923 & n3251;
  assign n3253 = ~n3140 & n3252;
  assign n3254 = ~n32596 & ~n3248;
  assign n3255 = ~n3253 & ~n3254;
  assign n3256 = ~n3249 & ~n3250;
  assign n3257 = ~n32637 & ~n32638;
  assign n3258 = ~n3243 & ~n3257;
  assign n3259 = ~n1192 & ~n3258;
  assign n3260 = n1192 & ~n3243;
  assign n3261 = ~n3257 & n3260;
  assign n3262 = ~n2937 & ~n32598;
  assign n3263 = ~n2937 & ~n3140;
  assign n3264 = ~n32598 & n3263;
  assign n3265 = ~n3140 & n3262;
  assign n3266 = n2945 & ~n32639;
  assign n3267 = n2949 & n3263;
  assign n3268 = n2945 & ~n32598;
  assign n3269 = ~n2937 & n3268;
  assign n3270 = ~n3140 & n3269;
  assign n3271 = ~n2945 & ~n32639;
  assign n3272 = ~n3270 & ~n3271;
  assign n3273 = ~n3266 & ~n3267;
  assign n3274 = ~n3261 & ~n32640;
  assign n3275 = ~n3259 & ~n3274;
  assign n3276 = ~n1028 & ~n3275;
  assign n3277 = n1028 & ~n3259;
  assign n3278 = ~n3274 & n3277;
  assign n3279 = n1028 & n3275;
  assign n3280 = ~n2951 & ~n2953;
  assign n3281 = ~n3140 & n3280;
  assign n3282 = ~n32599 & ~n3281;
  assign n3283 = ~n2951 & n32599;
  assign n3284 = ~n2953 & n3283;
  assign n3285 = n32599 & n3281;
  assign n3286 = ~n3140 & n3284;
  assign n3287 = ~n32599 & n3281;
  assign n3288 = n32599 & ~n3281;
  assign n3289 = ~n3287 & ~n3288;
  assign n3290 = ~n3282 & ~n32642;
  assign n3291 = ~n32641 & n32643;
  assign n3292 = ~n3276 & ~n3291;
  assign n3293 = ~n866 & ~n3292;
  assign n3294 = n866 & ~n3276;
  assign n3295 = ~n3291 & n3294;
  assign n3296 = ~n2966 & ~n32601;
  assign n3297 = ~n2966 & ~n3140;
  assign n3298 = ~n32601 & n3297;
  assign n3299 = ~n3140 & n3296;
  assign n3300 = n2974 & ~n32644;
  assign n3301 = n2978 & n3297;
  assign n3302 = n2974 & ~n32601;
  assign n3303 = ~n2966 & n3302;
  assign n3304 = ~n3140 & n3303;
  assign n3305 = ~n2974 & ~n32644;
  assign n3306 = ~n3304 & ~n3305;
  assign n3307 = ~n3300 & ~n3301;
  assign n3308 = ~n3295 & ~n32645;
  assign n3309 = ~n3293 & ~n3308;
  assign n3310 = ~n730 & ~n3309;
  assign n3311 = n730 & ~n3293;
  assign n3312 = ~n3308 & n3311;
  assign n3313 = n730 & n3309;
  assign n3314 = ~n2980 & ~n2982;
  assign n3315 = ~n3140 & n3314;
  assign n3316 = n32603 & ~n3315;
  assign n3317 = ~n2980 & ~n32603;
  assign n3318 = ~n2982 & n3317;
  assign n3319 = ~n32603 & n3315;
  assign n3320 = ~n3140 & n3318;
  assign n3321 = n32603 & n3315;
  assign n3322 = ~n32603 & ~n3315;
  assign n3323 = ~n3321 & ~n3322;
  assign n3324 = ~n3316 & ~n32647;
  assign n3325 = ~n32646 & n32648;
  assign n3326 = ~n3310 & ~n3325;
  assign n3327 = ~n602 & ~n3326;
  assign n3328 = n602 & ~n3310;
  assign n3329 = ~n3325 & n3328;
  assign n3330 = ~n2996 & ~n32605;
  assign n3331 = ~n2996 & ~n3140;
  assign n3332 = ~n32605 & n3331;
  assign n3333 = ~n3140 & n3330;
  assign n3334 = n3004 & ~n32649;
  assign n3335 = n3008 & n3331;
  assign n3336 = n3004 & ~n32605;
  assign n3337 = ~n2996 & n3336;
  assign n3338 = ~n3140 & n3337;
  assign n3339 = ~n3004 & ~n32649;
  assign n3340 = ~n3338 & ~n3339;
  assign n3341 = ~n3334 & ~n3335;
  assign n3342 = ~n3329 & ~n32650;
  assign n3343 = ~n3327 & ~n3342;
  assign n3344 = ~n497 & ~n3343;
  assign n3345 = n497 & ~n3327;
  assign n3346 = ~n3342 & n3345;
  assign n3347 = n497 & n3343;
  assign n3348 = ~n3010 & ~n3012;
  assign n3349 = ~n3010 & ~n3140;
  assign n3350 = ~n3012 & n3349;
  assign n3351 = ~n3140 & n3348;
  assign n3352 = ~n32607 & ~n32652;
  assign n3353 = n3024 & n3349;
  assign n3354 = n32607 & n32652;
  assign n3355 = ~n3010 & ~n32607;
  assign n3356 = ~n3012 & n3355;
  assign n3357 = ~n3140 & n3356;
  assign n3358 = n32607 & ~n32652;
  assign n3359 = ~n3357 & ~n3358;
  assign n3360 = ~n3352 & ~n32653;
  assign n3361 = ~n32651 & ~n32654;
  assign n3362 = ~n3344 & ~n3361;
  assign n3363 = ~n403 & ~n3362;
  assign n3364 = n403 & ~n3344;
  assign n3365 = ~n3361 & n3364;
  assign n3366 = ~n3026 & ~n32609;
  assign n3367 = ~n3026 & ~n3140;
  assign n3368 = ~n32609 & n3367;
  assign n3369 = ~n3140 & n3366;
  assign n3370 = n3034 & ~n32655;
  assign n3371 = n3038 & n3367;
  assign n3372 = n3034 & ~n32609;
  assign n3373 = ~n3026 & n3372;
  assign n3374 = ~n3140 & n3373;
  assign n3375 = ~n3034 & ~n32655;
  assign n3376 = ~n3374 & ~n3375;
  assign n3377 = ~n3370 & ~n3371;
  assign n3378 = ~n3365 & ~n32656;
  assign n3379 = ~n3363 & ~n3378;
  assign n3380 = ~n330 & ~n3379;
  assign n3381 = n330 & ~n3363;
  assign n3382 = ~n3378 & n3381;
  assign n3383 = n330 & n3379;
  assign n3384 = ~n3040 & ~n3042;
  assign n3385 = ~n3140 & n3384;
  assign n3386 = ~n32612 & ~n3385;
  assign n3387 = ~n3040 & n32612;
  assign n3388 = ~n3042 & n3387;
  assign n3389 = n32612 & n3385;
  assign n3390 = ~n3140 & n3388;
  assign n3391 = ~n3386 & ~n32658;
  assign n3392 = ~n32657 & ~n3391;
  assign n3393 = ~n3380 & ~n3392;
  assign n3394 = ~n271 & ~n3393;
  assign n3395 = n271 & ~n3380;
  assign n3396 = ~n3392 & n3395;
  assign n3397 = ~n3058 & ~n32614;
  assign n3398 = ~n3058 & ~n3140;
  assign n3399 = ~n32614 & n3398;
  assign n3400 = ~n3140 & n3397;
  assign n3401 = n3066 & ~n32659;
  assign n3402 = n3070 & n3398;
  assign n3403 = n3066 & ~n32614;
  assign n3404 = ~n3058 & n3403;
  assign n3405 = ~n3140 & n3404;
  assign n3406 = ~n3066 & ~n32659;
  assign n3407 = ~n3405 & ~n3406;
  assign n3408 = ~n3401 & ~n3402;
  assign n3409 = ~n3396 & ~n32660;
  assign n3410 = ~n3394 & ~n3409;
  assign n3411 = ~n217 & ~n3410;
  assign n3412 = n217 & ~n3394;
  assign n3413 = ~n3409 & n3412;
  assign n3414 = n217 & n3410;
  assign n3415 = ~n3072 & ~n3074;
  assign n3416 = ~n3072 & ~n3140;
  assign n3417 = ~n3074 & n3416;
  assign n3418 = ~n3140 & n3415;
  assign n3419 = n3082 & ~n32662;
  assign n3420 = n3083 & n3416;
  assign n3421 = ~n3082 & n32662;
  assign n3422 = ~n3072 & n3082;
  assign n3423 = ~n3074 & n3422;
  assign n3424 = ~n3140 & n3423;
  assign n3425 = ~n3082 & ~n32662;
  assign n3426 = ~n3424 & ~n3425;
  assign n3427 = ~n3419 & ~n32663;
  assign n3428 = ~n32661 & ~n32664;
  assign n3429 = ~n3411 & ~n3428;
  assign n3430 = ~n198 & ~n3429;
  assign n3431 = n198 & ~n3411;
  assign n3432 = ~n3428 & n3431;
  assign n3433 = ~n3085 & ~n32617;
  assign n3434 = ~n3085 & ~n3140;
  assign n3435 = ~n32617 & n3434;
  assign n3436 = ~n3140 & n3433;
  assign n3437 = n3093 & ~n32665;
  assign n3438 = n3097 & n3434;
  assign n3439 = n3093 & ~n32617;
  assign n3440 = ~n3085 & n3439;
  assign n3441 = ~n3140 & n3440;
  assign n3442 = ~n3093 & ~n32665;
  assign n3443 = ~n3441 & ~n3442;
  assign n3444 = ~n3437 & ~n3438;
  assign n3445 = ~n3432 & ~n32666;
  assign n3446 = ~n3430 & ~n3445;
  assign n3447 = ~n3099 & ~n3101;
  assign n3448 = ~n3140 & n3447;
  assign n3449 = ~n32620 & n3448;
  assign n3450 = n32620 & ~n3448;
  assign n3451 = ~n3099 & n32620;
  assign n3452 = ~n3101 & n3451;
  assign n3453 = n32620 & n3448;
  assign n3454 = ~n3140 & n3452;
  assign n3455 = ~n32620 & ~n3448;
  assign n3456 = ~n32667 & ~n3455;
  assign n3457 = ~n3449 & ~n3450;
  assign n3458 = ~n3116 & ~n3124;
  assign n3459 = ~n3124 & ~n3140;
  assign n3460 = ~n3116 & n3459;
  assign n3461 = ~n3140 & n3458;
  assign n3462 = ~n32623 & ~n32669;
  assign n3463 = ~n32668 & n3462;
  assign n3464 = ~n3446 & n3463;
  assign n3465 = n193 & ~n3464;
  assign n3466 = ~n3430 & n32668;
  assign n3467 = ~n3445 & n3466;
  assign n3468 = n3446 & n32668;
  assign n3469 = n3116 & ~n3459;
  assign n3470 = ~n193 & ~n3458;
  assign n3471 = ~n3469 & n3470;
  assign n3472 = ~n32670 & ~n3471;
  assign n3473 = ~n3465 & n3472;
  assign n3474 = pi86  & ~n3473;
  assign n3475 = ~pi84  & ~pi85 ;
  assign n3476 = ~pi86  & n3475;
  assign n3477 = ~n3474 & ~n3476;
  assign n3478 = ~n3140 & ~n3477;
  assign n3479 = ~n2836 & ~n32625;
  assign n3480 = ~n2837 & n3479;
  assign n3481 = ~n2853 & n3480;
  assign n3482 = ~n32586 & n3481;
  assign n3483 = n32584 & n2855;
  assign n3484 = ~n2847 & n3482;
  assign n3485 = ~n3476 & ~n32671;
  assign n3486 = ~n3138 & n3485;
  assign n3487 = ~n32623 & n3486;
  assign n3488 = ~n3132 & n3487;
  assign n3489 = n3140 & n3477;
  assign n3490 = ~n3474 & n3488;
  assign n3491 = ~pi86  & ~n3473;
  assign n3492 = pi87  & ~n3491;
  assign n3493 = ~pi87  & n3491;
  assign n3494 = n3142 & ~n3473;
  assign n3495 = ~n3492 & ~n32673;
  assign n3496 = ~n32672 & n3495;
  assign n3497 = ~n3478 & ~n3496;
  assign n3498 = ~n2855 & ~n3497;
  assign n3499 = ~n3140 & ~n3471;
  assign n3500 = ~n32670 & n3499;
  assign n3501 = ~n3465 & n3500;
  assign n3502 = ~n32673 & ~n3501;
  assign n3503 = pi88  & ~n3502;
  assign n3504 = ~pi88  & ~n3501;
  assign n3505 = ~pi88  & n3502;
  assign n3506 = ~n32673 & n3504;
  assign n3507 = ~n3503 & ~n32674;
  assign n3508 = n2855 & ~n3478;
  assign n3509 = n2855 & n3497;
  assign n3510 = ~n3496 & n3508;
  assign n3511 = ~n3507 & ~n32675;
  assign n3512 = ~n3498 & ~n3511;
  assign n3513 = ~n2556 & ~n3512;
  assign n3514 = n2556 & ~n3498;
  assign n3515 = ~n3511 & n3514;
  assign n3516 = ~n3145 & ~n32626;
  assign n3517 = ~n3473 & n3516;
  assign n3518 = n3150 & ~n3517;
  assign n3519 = ~n3150 & n3516;
  assign n3520 = ~n3150 & n3517;
  assign n3521 = ~n3473 & n3519;
  assign n3522 = ~n3518 & ~n32676;
  assign n3523 = ~n3515 & ~n3522;
  assign n3524 = ~n3513 & ~n3523;
  assign n3525 = ~n2301 & ~n3524;
  assign n3526 = ~n3165 & ~n3167;
  assign n3527 = ~n3473 & n3526;
  assign n3528 = ~n3176 & ~n3527;
  assign n3529 = ~n3167 & n3176;
  assign n3530 = ~n3165 & n3529;
  assign n3531 = n3176 & n3527;
  assign n3532 = ~n3473 & n3530;
  assign n3533 = ~n3528 & ~n32677;
  assign n3534 = n2301 & ~n3513;
  assign n3535 = n2301 & n3524;
  assign n3536 = ~n3523 & n3534;
  assign n3537 = ~n3533 & ~n32678;
  assign n3538 = ~n3525 & ~n3537;
  assign n3539 = ~n2038 & ~n3538;
  assign n3540 = n2038 & ~n3525;
  assign n3541 = ~n3537 & n3540;
  assign n3542 = ~n3179 & ~n32628;
  assign n3543 = ~n3473 & n3542;
  assign n3544 = n3189 & ~n3543;
  assign n3545 = ~n3189 & n3543;
  assign n3546 = ~n3179 & n3189;
  assign n3547 = ~n32628 & n3546;
  assign n3548 = n3189 & n3543;
  assign n3549 = ~n3473 & n3547;
  assign n3550 = ~n3189 & ~n3543;
  assign n3551 = ~n32679 & ~n3550;
  assign n3552 = ~n3544 & ~n3545;
  assign n3553 = ~n3541 & ~n32680;
  assign n3554 = ~n3539 & ~n3553;
  assign n3555 = ~n1812 & ~n3554;
  assign n3556 = ~n3192 & ~n3194;
  assign n3557 = ~n3473 & n3556;
  assign n3558 = ~n32631 & ~n3557;
  assign n3559 = ~n3194 & n32631;
  assign n3560 = ~n3192 & n3559;
  assign n3561 = n32631 & n3557;
  assign n3562 = ~n3473 & n3560;
  assign n3563 = ~n3558 & ~n32681;
  assign n3564 = n1812 & ~n3539;
  assign n3565 = n1812 & n3554;
  assign n3566 = ~n3553 & n3564;
  assign n3567 = ~n3563 & ~n32682;
  assign n3568 = ~n3555 & ~n3567;
  assign n3569 = ~n1582 & ~n3568;
  assign n3570 = n1582 & ~n3555;
  assign n3571 = ~n3567 & n3570;
  assign n3572 = ~n3209 & ~n32632;
  assign n3573 = ~n3473 & n3572;
  assign n3574 = ~n32634 & n3573;
  assign n3575 = n32634 & ~n3573;
  assign n3576 = ~n3209 & n32634;
  assign n3577 = ~n32632 & n3576;
  assign n3578 = ~n3473 & n3577;
  assign n3579 = ~n32634 & ~n3573;
  assign n3580 = ~n3578 & ~n3579;
  assign n3581 = ~n3574 & ~n3575;
  assign n3582 = ~n3571 & ~n32683;
  assign n3583 = ~n3569 & ~n3582;
  assign n3584 = ~n1388 & ~n3583;
  assign n3585 = ~n3226 & ~n3228;
  assign n3586 = ~n3473 & n3585;
  assign n3587 = ~n32636 & ~n3586;
  assign n3588 = ~n3228 & n32636;
  assign n3589 = ~n3226 & n3588;
  assign n3590 = n32636 & n3586;
  assign n3591 = ~n3473 & n3589;
  assign n3592 = ~n3587 & ~n32684;
  assign n3593 = n1388 & ~n3569;
  assign n3594 = n1388 & n3583;
  assign n3595 = ~n3582 & n3593;
  assign n3596 = ~n3592 & ~n32685;
  assign n3597 = ~n3584 & ~n3596;
  assign n3598 = ~n1192 & ~n3597;
  assign n3599 = n1192 & ~n3584;
  assign n3600 = ~n3596 & n3599;
  assign n3601 = ~n3243 & ~n32637;
  assign n3602 = ~n3473 & n3601;
  assign n3603 = ~n32638 & ~n3602;
  assign n3604 = ~n3243 & n32638;
  assign n3605 = ~n32637 & n3604;
  assign n3606 = n32638 & n3602;
  assign n3607 = ~n3473 & n3605;
  assign n3608 = n32638 & ~n3602;
  assign n3609 = ~n32638 & n3602;
  assign n3610 = ~n3608 & ~n3609;
  assign n3611 = ~n3603 & ~n32686;
  assign n3612 = ~n3600 & n32687;
  assign n3613 = ~n3598 & ~n3612;
  assign n3614 = ~n1028 & ~n3613;
  assign n3615 = ~n3259 & ~n3261;
  assign n3616 = ~n3473 & n3615;
  assign n3617 = ~n32640 & ~n3616;
  assign n3618 = ~n3261 & n32640;
  assign n3619 = ~n3259 & n3618;
  assign n3620 = n32640 & n3616;
  assign n3621 = ~n3473 & n3619;
  assign n3622 = ~n3617 & ~n32688;
  assign n3623 = n1028 & ~n3598;
  assign n3624 = n1028 & n3613;
  assign n3625 = ~n3612 & n3623;
  assign n3626 = ~n3622 & ~n32689;
  assign n3627 = ~n3614 & ~n3626;
  assign n3628 = ~n866 & ~n3627;
  assign n3629 = n866 & ~n3614;
  assign n3630 = ~n3626 & n3629;
  assign n3631 = ~n3276 & ~n32641;
  assign n3632 = ~n3473 & n3631;
  assign n3633 = ~n32643 & ~n3632;
  assign n3634 = n32643 & n3632;
  assign n3635 = ~n3276 & ~n32643;
  assign n3636 = ~n32641 & n3635;
  assign n3637 = ~n32643 & n3632;
  assign n3638 = ~n3473 & n3636;
  assign n3639 = n32643 & ~n3632;
  assign n3640 = ~n32690 & ~n3639;
  assign n3641 = ~n3633 & ~n3634;
  assign n3642 = ~n3630 & ~n32691;
  assign n3643 = ~n3628 & ~n3642;
  assign n3644 = ~n730 & ~n3643;
  assign n3645 = ~n3293 & ~n3295;
  assign n3646 = ~n3473 & n3645;
  assign n3647 = ~n32645 & ~n3646;
  assign n3648 = ~n3295 & n32645;
  assign n3649 = ~n3293 & n3648;
  assign n3650 = n32645 & n3646;
  assign n3651 = ~n3473 & n3649;
  assign n3652 = ~n3647 & ~n32692;
  assign n3653 = n730 & ~n3628;
  assign n3654 = n730 & n3643;
  assign n3655 = ~n3642 & n3653;
  assign n3656 = ~n3652 & ~n32693;
  assign n3657 = ~n3644 & ~n3656;
  assign n3658 = ~n602 & ~n3657;
  assign n3659 = n602 & ~n3644;
  assign n3660 = ~n3656 & n3659;
  assign n3661 = ~n3310 & ~n32646;
  assign n3662 = ~n3310 & ~n3473;
  assign n3663 = ~n32646 & n3662;
  assign n3664 = ~n3473 & n3661;
  assign n3665 = ~n32648 & ~n32694;
  assign n3666 = n3325 & n3662;
  assign n3667 = n32648 & n32694;
  assign n3668 = ~n3310 & ~n32648;
  assign n3669 = ~n32646 & n3668;
  assign n3670 = ~n3473 & n3669;
  assign n3671 = n32648 & ~n32694;
  assign n3672 = ~n3670 & ~n3671;
  assign n3673 = ~n3665 & ~n32695;
  assign n3674 = ~n3660 & ~n32696;
  assign n3675 = ~n3658 & ~n3674;
  assign n3676 = ~n497 & ~n3675;
  assign n3677 = ~n3327 & ~n3329;
  assign n3678 = ~n3473 & n3677;
  assign n3679 = ~n32650 & ~n3678;
  assign n3680 = ~n3329 & n32650;
  assign n3681 = ~n3327 & n3680;
  assign n3682 = n32650 & n3678;
  assign n3683 = ~n3473 & n3681;
  assign n3684 = ~n3679 & ~n32697;
  assign n3685 = n497 & ~n3658;
  assign n3686 = n497 & n3675;
  assign n3687 = ~n3674 & n3685;
  assign n3688 = ~n3684 & ~n32698;
  assign n3689 = ~n3676 & ~n3688;
  assign n3690 = ~n403 & ~n3689;
  assign n3691 = n403 & ~n3676;
  assign n3692 = ~n3688 & n3691;
  assign n3693 = ~n3344 & ~n32651;
  assign n3694 = ~n3473 & n3693;
  assign n3695 = ~n32654 & ~n3694;
  assign n3696 = ~n3344 & n32654;
  assign n3697 = ~n32651 & n3696;
  assign n3698 = n32654 & n3694;
  assign n3699 = ~n3473 & n3697;
  assign n3700 = ~n3695 & ~n32699;
  assign n3701 = ~n3692 & ~n3700;
  assign n3702 = ~n3690 & ~n3701;
  assign n3703 = ~n330 & ~n3702;
  assign n3704 = ~n3363 & ~n3365;
  assign n3705 = ~n3473 & n3704;
  assign n3706 = ~n32656 & ~n3705;
  assign n3707 = ~n3365 & n32656;
  assign n3708 = ~n3363 & n3707;
  assign n3709 = n32656 & n3705;
  assign n3710 = ~n3473 & n3708;
  assign n3711 = ~n3706 & ~n32700;
  assign n3712 = n330 & ~n3690;
  assign n3713 = n330 & n3702;
  assign n3714 = ~n3701 & n3712;
  assign n3715 = ~n3711 & ~n32701;
  assign n3716 = ~n3703 & ~n3715;
  assign n3717 = ~n271 & ~n3716;
  assign n3718 = n271 & ~n3703;
  assign n3719 = ~n3715 & n3718;
  assign n3720 = ~n3380 & ~n32657;
  assign n3721 = ~n3380 & ~n3473;
  assign n3722 = ~n32657 & n3721;
  assign n3723 = ~n3473 & n3720;
  assign n3724 = n3391 & ~n32702;
  assign n3725 = n3392 & n3721;
  assign n3726 = ~n3391 & n32702;
  assign n3727 = ~n3380 & n3391;
  assign n3728 = ~n32657 & n3727;
  assign n3729 = ~n3473 & n3728;
  assign n3730 = ~n3391 & ~n32702;
  assign n3731 = ~n3729 & ~n3730;
  assign n3732 = ~n3724 & ~n32703;
  assign n3733 = ~n3719 & ~n32704;
  assign n3734 = ~n3717 & ~n3733;
  assign n3735 = ~n217 & ~n3734;
  assign n3736 = ~n3394 & ~n3396;
  assign n3737 = ~n3473 & n3736;
  assign n3738 = ~n32660 & ~n3737;
  assign n3739 = ~n3396 & n32660;
  assign n3740 = ~n3394 & n3739;
  assign n3741 = n32660 & n3737;
  assign n3742 = ~n3473 & n3740;
  assign n3743 = ~n3738 & ~n32705;
  assign n3744 = n217 & ~n3717;
  assign n3745 = n217 & n3734;
  assign n3746 = ~n3733 & n3744;
  assign n3747 = ~n3743 & ~n32706;
  assign n3748 = ~n3735 & ~n3747;
  assign n3749 = ~n198 & ~n3748;
  assign n3750 = n198 & ~n3735;
  assign n3751 = ~n3747 & n3750;
  assign n3752 = ~n3411 & ~n32661;
  assign n3753 = ~n3473 & n3752;
  assign n3754 = ~n32664 & n3753;
  assign n3755 = n32664 & ~n3753;
  assign n3756 = ~n3411 & n32664;
  assign n3757 = ~n32661 & n3756;
  assign n3758 = n32664 & n3753;
  assign n3759 = ~n3473 & n3757;
  assign n3760 = ~n32664 & ~n3753;
  assign n3761 = ~n32707 & ~n3760;
  assign n3762 = ~n3754 & ~n3755;
  assign n3763 = ~n3751 & ~n32708;
  assign n3764 = ~n3749 & ~n3763;
  assign n3765 = ~n3430 & ~n3432;
  assign n3766 = ~n3473 & n3765;
  assign n3767 = ~n32666 & ~n3766;
  assign n3768 = ~n3432 & n32666;
  assign n3769 = ~n3430 & n3768;
  assign n3770 = n32666 & n3766;
  assign n3771 = ~n3473 & n3769;
  assign n3772 = ~n3767 & ~n32709;
  assign n3773 = ~n3446 & ~n32668;
  assign n3774 = ~n32668 & ~n3473;
  assign n3775 = ~n3446 & n3774;
  assign n3776 = ~n3473 & n3773;
  assign n3777 = ~n32670 & ~n32710;
  assign n3778 = ~n3772 & n3777;
  assign n3779 = ~n3764 & n3778;
  assign n3780 = n193 & ~n3779;
  assign n3781 = ~n3749 & n3772;
  assign n3782 = n3764 & n3772;
  assign n3783 = ~n3763 & n3781;
  assign n3784 = n3446 & ~n3774;
  assign n3785 = ~n193 & ~n3773;
  assign n3786 = ~n3784 & n3785;
  assign n3787 = ~n32711 & ~n3786;
  assign n3788 = ~n3780 & n3787;
  assign n3789 = pi84  & ~n3788;
  assign n3790 = ~pi82  & ~pi83 ;
  assign n3791 = ~pi84  & n3790;
  assign n3792 = ~n3789 & ~n3791;
  assign n3793 = ~n3473 & ~n3792;
  assign n3794 = ~pi84  & ~n3788;
  assign n3795 = pi85  & ~n3794;
  assign n3796 = ~pi85  & n3794;
  assign n3797 = n3475 & ~n3788;
  assign n3798 = ~n3795 & ~n32712;
  assign n3799 = ~n32621 & ~n32671;
  assign n3800 = ~n3119 & n3799;
  assign n3801 = ~n3138 & n3800;
  assign n3802 = ~n32623 & n3801;
  assign n3803 = n3124 & n3140;
  assign n3804 = ~n3132 & n3802;
  assign n3805 = ~n3791 & ~n32713;
  assign n3806 = ~n3471 & n3805;
  assign n3807 = ~n32670 & n3806;
  assign n3808 = ~n3465 & n3807;
  assign n3809 = n3473 & n3792;
  assign n3810 = ~n3789 & n3808;
  assign n3811 = n3798 & ~n32714;
  assign n3812 = ~n3793 & ~n3811;
  assign n3813 = ~n3140 & ~n3812;
  assign n3814 = n3140 & ~n3793;
  assign n3815 = ~n3811 & n3814;
  assign n3816 = ~n3473 & ~n3786;
  assign n3817 = ~n32711 & n3816;
  assign n3818 = ~n3780 & n3817;
  assign n3819 = ~n32712 & ~n3818;
  assign n3820 = pi86  & ~n3819;
  assign n3821 = ~pi86  & ~n3818;
  assign n3822 = ~pi86  & n3819;
  assign n3823 = ~n32712 & n3821;
  assign n3824 = ~n3820 & ~n32715;
  assign n3825 = ~n3815 & ~n3824;
  assign n3826 = ~n3813 & ~n3825;
  assign n3827 = ~n2855 & ~n3826;
  assign n3828 = n2855 & ~n3813;
  assign n3829 = ~n3825 & n3828;
  assign n3830 = n2855 & n3826;
  assign n3831 = ~n3478 & ~n32672;
  assign n3832 = ~n3788 & n3831;
  assign n3833 = n3495 & ~n3832;
  assign n3834 = ~n3495 & n3831;
  assign n3835 = ~n3495 & n3832;
  assign n3836 = ~n3788 & n3834;
  assign n3837 = ~n3833 & ~n32717;
  assign n3838 = ~n32716 & ~n3837;
  assign n3839 = ~n3827 & ~n3838;
  assign n3840 = ~n2556 & ~n3839;
  assign n3841 = n2556 & ~n3827;
  assign n3842 = ~n3838 & n3841;
  assign n3843 = ~n3498 & ~n32675;
  assign n3844 = ~n3498 & ~n3788;
  assign n3845 = ~n32675 & n3844;
  assign n3846 = ~n3788 & n3843;
  assign n3847 = n3507 & ~n32718;
  assign n3848 = n3511 & n3844;
  assign n3849 = n3507 & ~n32675;
  assign n3850 = ~n3498 & n3849;
  assign n3851 = ~n3788 & n3850;
  assign n3852 = ~n3507 & ~n32718;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = ~n3847 & ~n3848;
  assign n3855 = ~n3842 & ~n32719;
  assign n3856 = ~n3840 & ~n3855;
  assign n3857 = ~n2301 & ~n3856;
  assign n3858 = n2301 & ~n3840;
  assign n3859 = ~n3855 & n3858;
  assign n3860 = n2301 & n3856;
  assign n3861 = ~n3513 & ~n3515;
  assign n3862 = ~n3788 & n3861;
  assign n3863 = n3522 & ~n3862;
  assign n3864 = ~n3522 & n3862;
  assign n3865 = ~n3513 & n3522;
  assign n3866 = ~n3515 & n3865;
  assign n3867 = n3522 & n3862;
  assign n3868 = ~n3788 & n3866;
  assign n3869 = ~n3522 & ~n3862;
  assign n3870 = ~n32721 & ~n3869;
  assign n3871 = ~n3863 & ~n3864;
  assign n3872 = ~n32720 & ~n32722;
  assign n3873 = ~n3857 & ~n3872;
  assign n3874 = ~n2038 & ~n3873;
  assign n3875 = n2038 & ~n3857;
  assign n3876 = ~n3872 & n3875;
  assign n3877 = ~n3525 & ~n32678;
  assign n3878 = ~n3525 & ~n3788;
  assign n3879 = ~n32678 & n3878;
  assign n3880 = ~n3788 & n3877;
  assign n3881 = n3533 & ~n32723;
  assign n3882 = n3537 & n3878;
  assign n3883 = n3533 & ~n32678;
  assign n3884 = ~n3525 & n3883;
  assign n3885 = ~n3788 & n3884;
  assign n3886 = ~n3533 & ~n32723;
  assign n3887 = ~n3885 & ~n3886;
  assign n3888 = ~n3881 & ~n3882;
  assign n3889 = ~n3876 & ~n32724;
  assign n3890 = ~n3874 & ~n3889;
  assign n3891 = ~n1812 & ~n3890;
  assign n3892 = n1812 & ~n3874;
  assign n3893 = ~n3889 & n3892;
  assign n3894 = n1812 & n3890;
  assign n3895 = ~n3539 & ~n3541;
  assign n3896 = ~n3788 & n3895;
  assign n3897 = ~n32680 & n3896;
  assign n3898 = n32680 & ~n3896;
  assign n3899 = ~n3539 & n32680;
  assign n3900 = ~n3541 & n3899;
  assign n3901 = ~n3788 & n3900;
  assign n3902 = ~n32680 & ~n3896;
  assign n3903 = ~n3901 & ~n3902;
  assign n3904 = ~n3897 & ~n3898;
  assign n3905 = ~n32725 & ~n32726;
  assign n3906 = ~n3891 & ~n3905;
  assign n3907 = ~n1582 & ~n3906;
  assign n3908 = n1582 & ~n3891;
  assign n3909 = ~n3905 & n3908;
  assign n3910 = ~n3555 & ~n32682;
  assign n3911 = ~n3555 & ~n3788;
  assign n3912 = ~n32682 & n3911;
  assign n3913 = ~n3788 & n3910;
  assign n3914 = n3563 & ~n32727;
  assign n3915 = n3567 & n3911;
  assign n3916 = n3563 & ~n32682;
  assign n3917 = ~n3555 & n3916;
  assign n3918 = ~n3788 & n3917;
  assign n3919 = ~n3563 & ~n32727;
  assign n3920 = ~n3918 & ~n3919;
  assign n3921 = ~n3914 & ~n3915;
  assign n3922 = ~n3909 & ~n32728;
  assign n3923 = ~n3907 & ~n3922;
  assign n3924 = ~n1388 & ~n3923;
  assign n3925 = n1388 & ~n3907;
  assign n3926 = ~n3922 & n3925;
  assign n3927 = n1388 & n3923;
  assign n3928 = ~n3569 & ~n3571;
  assign n3929 = ~n3788 & n3928;
  assign n3930 = ~n32683 & ~n3929;
  assign n3931 = ~n3569 & n32683;
  assign n3932 = ~n3571 & n3931;
  assign n3933 = n32683 & n3929;
  assign n3934 = ~n3788 & n3932;
  assign n3935 = n32683 & ~n3929;
  assign n3936 = ~n32683 & n3929;
  assign n3937 = ~n3935 & ~n3936;
  assign n3938 = ~n3930 & ~n32730;
  assign n3939 = ~n32729 & n32731;
  assign n3940 = ~n3924 & ~n3939;
  assign n3941 = ~n1192 & ~n3940;
  assign n3942 = n1192 & ~n3924;
  assign n3943 = ~n3939 & n3942;
  assign n3944 = ~n3584 & ~n32685;
  assign n3945 = ~n3584 & ~n3788;
  assign n3946 = ~n32685 & n3945;
  assign n3947 = ~n3788 & n3944;
  assign n3948 = n3592 & ~n32732;
  assign n3949 = n3596 & n3945;
  assign n3950 = n3592 & ~n32685;
  assign n3951 = ~n3584 & n3950;
  assign n3952 = ~n3788 & n3951;
  assign n3953 = ~n3592 & ~n32732;
  assign n3954 = ~n3952 & ~n3953;
  assign n3955 = ~n3948 & ~n3949;
  assign n3956 = ~n3943 & ~n32733;
  assign n3957 = ~n3941 & ~n3956;
  assign n3958 = ~n1028 & ~n3957;
  assign n3959 = n1028 & ~n3941;
  assign n3960 = ~n3956 & n3959;
  assign n3961 = n1028 & n3957;
  assign n3962 = ~n3598 & ~n3600;
  assign n3963 = ~n3788 & n3962;
  assign n3964 = n32687 & ~n3963;
  assign n3965 = ~n3598 & ~n32687;
  assign n3966 = ~n3600 & n3965;
  assign n3967 = ~n32687 & n3963;
  assign n3968 = ~n3788 & n3966;
  assign n3969 = n32687 & n3963;
  assign n3970 = ~n32687 & ~n3963;
  assign n3971 = ~n3969 & ~n3970;
  assign n3972 = ~n3964 & ~n32735;
  assign n3973 = ~n32734 & n32736;
  assign n3974 = ~n3958 & ~n3973;
  assign n3975 = ~n866 & ~n3974;
  assign n3976 = n866 & ~n3958;
  assign n3977 = ~n3973 & n3976;
  assign n3978 = ~n3614 & ~n32689;
  assign n3979 = ~n3614 & ~n3788;
  assign n3980 = ~n32689 & n3979;
  assign n3981 = ~n3788 & n3978;
  assign n3982 = n3622 & ~n32737;
  assign n3983 = n3626 & n3979;
  assign n3984 = n3622 & ~n32689;
  assign n3985 = ~n3614 & n3984;
  assign n3986 = ~n3788 & n3985;
  assign n3987 = ~n3622 & ~n32737;
  assign n3988 = ~n3986 & ~n3987;
  assign n3989 = ~n3982 & ~n3983;
  assign n3990 = ~n3977 & ~n32738;
  assign n3991 = ~n3975 & ~n3990;
  assign n3992 = ~n730 & ~n3991;
  assign n3993 = n730 & ~n3975;
  assign n3994 = ~n3990 & n3993;
  assign n3995 = n730 & n3991;
  assign n3996 = ~n3628 & ~n3630;
  assign n3997 = ~n3788 & n3996;
  assign n3998 = ~n32691 & n3997;
  assign n3999 = n32691 & ~n3997;
  assign n4000 = ~n3628 & n32691;
  assign n4001 = ~n3630 & n4000;
  assign n4002 = n32691 & n3997;
  assign n4003 = ~n3788 & n4001;
  assign n4004 = ~n32691 & ~n3997;
  assign n4005 = ~n32740 & ~n4004;
  assign n4006 = ~n3998 & ~n3999;
  assign n4007 = ~n32739 & ~n32741;
  assign n4008 = ~n3992 & ~n4007;
  assign n4009 = ~n602 & ~n4008;
  assign n4010 = n602 & ~n3992;
  assign n4011 = ~n4007 & n4010;
  assign n4012 = ~n3644 & ~n32693;
  assign n4013 = ~n3644 & ~n3788;
  assign n4014 = ~n32693 & n4013;
  assign n4015 = ~n3788 & n4012;
  assign n4016 = n3652 & ~n32742;
  assign n4017 = n3656 & n4013;
  assign n4018 = n3652 & ~n32693;
  assign n4019 = ~n3644 & n4018;
  assign n4020 = ~n3788 & n4019;
  assign n4021 = ~n3652 & ~n32742;
  assign n4022 = ~n4020 & ~n4021;
  assign n4023 = ~n4016 & ~n4017;
  assign n4024 = ~n4011 & ~n32743;
  assign n4025 = ~n4009 & ~n4024;
  assign n4026 = ~n497 & ~n4025;
  assign n4027 = n497 & ~n4009;
  assign n4028 = ~n4024 & n4027;
  assign n4029 = n497 & n4025;
  assign n4030 = ~n3658 & ~n3660;
  assign n4031 = ~n3788 & n4030;
  assign n4032 = ~n32696 & ~n4031;
  assign n4033 = ~n3658 & n32696;
  assign n4034 = ~n3660 & n4033;
  assign n4035 = n32696 & n4031;
  assign n4036 = ~n3788 & n4034;
  assign n4037 = ~n4032 & ~n32745;
  assign n4038 = ~n32744 & ~n4037;
  assign n4039 = ~n4026 & ~n4038;
  assign n4040 = ~n403 & ~n4039;
  assign n4041 = n403 & ~n4026;
  assign n4042 = ~n4038 & n4041;
  assign n4043 = ~n3676 & ~n32698;
  assign n4044 = ~n3676 & ~n3788;
  assign n4045 = ~n32698 & n4044;
  assign n4046 = ~n3788 & n4043;
  assign n4047 = n3684 & ~n32746;
  assign n4048 = n3688 & n4044;
  assign n4049 = n3684 & ~n32698;
  assign n4050 = ~n3676 & n4049;
  assign n4051 = ~n3788 & n4050;
  assign n4052 = ~n3684 & ~n32746;
  assign n4053 = ~n4051 & ~n4052;
  assign n4054 = ~n4047 & ~n4048;
  assign n4055 = ~n4042 & ~n32747;
  assign n4056 = ~n4040 & ~n4055;
  assign n4057 = ~n330 & ~n4056;
  assign n4058 = n330 & ~n4040;
  assign n4059 = ~n4055 & n4058;
  assign n4060 = n330 & n4056;
  assign n4061 = ~n3690 & ~n3692;
  assign n4062 = ~n3690 & ~n3788;
  assign n4063 = ~n3692 & n4062;
  assign n4064 = ~n3788 & n4061;
  assign n4065 = n3700 & ~n32749;
  assign n4066 = n3701 & n4062;
  assign n4067 = ~n3700 & n32749;
  assign n4068 = ~n3690 & n3700;
  assign n4069 = ~n3692 & n4068;
  assign n4070 = ~n3788 & n4069;
  assign n4071 = ~n3700 & ~n32749;
  assign n4072 = ~n4070 & ~n4071;
  assign n4073 = ~n4065 & ~n32750;
  assign n4074 = ~n32748 & ~n32751;
  assign n4075 = ~n4057 & ~n4074;
  assign n4076 = ~n271 & ~n4075;
  assign n4077 = n271 & ~n4057;
  assign n4078 = ~n4074 & n4077;
  assign n4079 = ~n3703 & ~n32701;
  assign n4080 = ~n3703 & ~n3788;
  assign n4081 = ~n32701 & n4080;
  assign n4082 = ~n3788 & n4079;
  assign n4083 = n3711 & ~n32752;
  assign n4084 = n3715 & n4080;
  assign n4085 = n3711 & ~n32701;
  assign n4086 = ~n3703 & n4085;
  assign n4087 = ~n3788 & n4086;
  assign n4088 = ~n3711 & ~n32752;
  assign n4089 = ~n4087 & ~n4088;
  assign n4090 = ~n4083 & ~n4084;
  assign n4091 = ~n4078 & ~n32753;
  assign n4092 = ~n4076 & ~n4091;
  assign n4093 = ~n217 & ~n4092;
  assign n4094 = n217 & ~n4076;
  assign n4095 = ~n4091 & n4094;
  assign n4096 = n217 & n4092;
  assign n4097 = ~n3717 & ~n3719;
  assign n4098 = ~n3788 & n4097;
  assign n4099 = ~n32704 & n4098;
  assign n4100 = n32704 & ~n4098;
  assign n4101 = ~n3717 & n32704;
  assign n4102 = ~n3719 & n4101;
  assign n4103 = n32704 & n4098;
  assign n4104 = ~n3788 & n4102;
  assign n4105 = ~n32704 & ~n4098;
  assign n4106 = ~n32755 & ~n4105;
  assign n4107 = ~n4099 & ~n4100;
  assign n4108 = ~n32754 & ~n32756;
  assign n4109 = ~n4093 & ~n4108;
  assign n4110 = ~n198 & ~n4109;
  assign n4111 = n198 & ~n4093;
  assign n4112 = ~n4108 & n4111;
  assign n4113 = ~n3735 & ~n32706;
  assign n4114 = ~n3735 & ~n3788;
  assign n4115 = ~n32706 & n4114;
  assign n4116 = ~n3788 & n4113;
  assign n4117 = n3743 & ~n32757;
  assign n4118 = n3747 & n4114;
  assign n4119 = n3743 & ~n32706;
  assign n4120 = ~n3735 & n4119;
  assign n4121 = ~n3788 & n4120;
  assign n4122 = ~n3743 & ~n32757;
  assign n4123 = ~n4121 & ~n4122;
  assign n4124 = ~n4117 & ~n4118;
  assign n4125 = ~n4112 & ~n32758;
  assign n4126 = ~n4110 & ~n4125;
  assign n4127 = ~n3749 & ~n3751;
  assign n4128 = ~n3749 & ~n3788;
  assign n4129 = ~n3751 & n4128;
  assign n4130 = ~n3788 & n4127;
  assign n4131 = n32708 & ~n32759;
  assign n4132 = n3763 & n4128;
  assign n4133 = ~n32708 & n32759;
  assign n4134 = ~n3749 & n32708;
  assign n4135 = ~n3751 & n4134;
  assign n4136 = ~n3788 & n4135;
  assign n4137 = ~n32708 & ~n32759;
  assign n4138 = ~n4136 & ~n4137;
  assign n4139 = ~n4131 & ~n32760;
  assign n4140 = ~n3764 & ~n3772;
  assign n4141 = ~n3772 & ~n3788;
  assign n4142 = ~n3764 & n4141;
  assign n4143 = ~n3788 & n4140;
  assign n4144 = ~n32711 & ~n32762;
  assign n4145 = ~n32761 & n4144;
  assign n4146 = ~n4126 & n4145;
  assign n4147 = n193 & ~n4146;
  assign n4148 = ~n4110 & n32761;
  assign n4149 = ~n4125 & n4148;
  assign n4150 = n4126 & n32761;
  assign n4151 = n3764 & ~n4141;
  assign n4152 = ~n193 & ~n4140;
  assign n4153 = ~n4151 & n4152;
  assign n4154 = ~n32763 & ~n4153;
  assign n4155 = ~n4147 & n4154;
  assign n4156 = pi82  & ~n4155;
  assign n4157 = ~pi80  & ~pi81 ;
  assign n4158 = ~pi82  & n4157;
  assign n4159 = ~n4156 & ~n4158;
  assign n4160 = ~n3788 & ~n4159;
  assign n4161 = ~n32667 & ~n32713;
  assign n4162 = ~n3455 & n4161;
  assign n4163 = ~n3471 & n4162;
  assign n4164 = ~n32670 & n4163;
  assign n4165 = n32668 & n3473;
  assign n4166 = ~n3465 & n4164;
  assign n4167 = ~n4158 & ~n32764;
  assign n4168 = ~n3786 & n4167;
  assign n4169 = ~n32711 & n4168;
  assign n4170 = ~n3780 & n4169;
  assign n4171 = n3788 & n4159;
  assign n4172 = ~n4156 & n4170;
  assign n4173 = ~pi82  & ~n4155;
  assign n4174 = pi83  & ~n4173;
  assign n4175 = ~pi83  & n4173;
  assign n4176 = n3790 & ~n4155;
  assign n4177 = ~n4174 & ~n32766;
  assign n4178 = ~n32765 & n4177;
  assign n4179 = ~n4160 & ~n4178;
  assign n4180 = ~n3473 & ~n4179;
  assign n4181 = ~n3788 & ~n4153;
  assign n4182 = ~n32763 & n4181;
  assign n4183 = ~n4147 & n4182;
  assign n4184 = ~n32766 & ~n4183;
  assign n4185 = pi84  & ~n4184;
  assign n4186 = ~pi84  & ~n4183;
  assign n4187 = ~pi84  & n4184;
  assign n4188 = ~n32766 & n4186;
  assign n4189 = ~n4185 & ~n32767;
  assign n4190 = n3473 & ~n4160;
  assign n4191 = n3473 & n4179;
  assign n4192 = ~n4178 & n4190;
  assign n4193 = ~n4189 & ~n32768;
  assign n4194 = ~n4180 & ~n4193;
  assign n4195 = ~n3140 & ~n4194;
  assign n4196 = n3140 & ~n4180;
  assign n4197 = ~n4193 & n4196;
  assign n4198 = ~n3793 & ~n32714;
  assign n4199 = ~n4155 & n4198;
  assign n4200 = n3798 & ~n4199;
  assign n4201 = ~n3798 & n4198;
  assign n4202 = ~n3798 & n4199;
  assign n4203 = ~n4155 & n4201;
  assign n4204 = ~n4200 & ~n32769;
  assign n4205 = ~n4197 & ~n4204;
  assign n4206 = ~n4195 & ~n4205;
  assign n4207 = ~n2855 & ~n4206;
  assign n4208 = ~n3813 & ~n3815;
  assign n4209 = ~n4155 & n4208;
  assign n4210 = ~n3824 & ~n4209;
  assign n4211 = ~n3815 & n3824;
  assign n4212 = ~n3813 & n4211;
  assign n4213 = n3824 & n4209;
  assign n4214 = ~n4155 & n4212;
  assign n4215 = ~n4210 & ~n32770;
  assign n4216 = n2855 & ~n4195;
  assign n4217 = n2855 & n4206;
  assign n4218 = ~n4205 & n4216;
  assign n4219 = ~n4215 & ~n32771;
  assign n4220 = ~n4207 & ~n4219;
  assign n4221 = ~n2556 & ~n4220;
  assign n4222 = n2556 & ~n4207;
  assign n4223 = ~n4219 & n4222;
  assign n4224 = ~n3827 & ~n32716;
  assign n4225 = ~n4155 & n4224;
  assign n4226 = n3837 & ~n4225;
  assign n4227 = ~n3837 & n4225;
  assign n4228 = ~n3827 & n3837;
  assign n4229 = ~n32716 & n4228;
  assign n4230 = n3837 & n4225;
  assign n4231 = ~n4155 & n4229;
  assign n4232 = ~n3837 & ~n4225;
  assign n4233 = ~n32772 & ~n4232;
  assign n4234 = ~n4226 & ~n4227;
  assign n4235 = ~n4223 & ~n32773;
  assign n4236 = ~n4221 & ~n4235;
  assign n4237 = ~n2301 & ~n4236;
  assign n4238 = ~n3840 & ~n3842;
  assign n4239 = ~n4155 & n4238;
  assign n4240 = ~n32719 & ~n4239;
  assign n4241 = ~n3842 & n32719;
  assign n4242 = ~n3840 & n4241;
  assign n4243 = n32719 & n4239;
  assign n4244 = ~n4155 & n4242;
  assign n4245 = ~n4240 & ~n32774;
  assign n4246 = n2301 & ~n4221;
  assign n4247 = n2301 & n4236;
  assign n4248 = ~n4235 & n4246;
  assign n4249 = ~n4245 & ~n32775;
  assign n4250 = ~n4237 & ~n4249;
  assign n4251 = ~n2038 & ~n4250;
  assign n4252 = n2038 & ~n4237;
  assign n4253 = ~n4249 & n4252;
  assign n4254 = ~n3857 & ~n32720;
  assign n4255 = ~n4155 & n4254;
  assign n4256 = ~n32722 & n4255;
  assign n4257 = n32722 & ~n4255;
  assign n4258 = ~n3857 & n32722;
  assign n4259 = ~n32720 & n4258;
  assign n4260 = ~n4155 & n4259;
  assign n4261 = ~n32722 & ~n4255;
  assign n4262 = ~n4260 & ~n4261;
  assign n4263 = ~n4256 & ~n4257;
  assign n4264 = ~n4253 & ~n32776;
  assign n4265 = ~n4251 & ~n4264;
  assign n4266 = ~n1812 & ~n4265;
  assign n4267 = ~n3874 & ~n3876;
  assign n4268 = ~n4155 & n4267;
  assign n4269 = ~n32724 & ~n4268;
  assign n4270 = ~n3876 & n32724;
  assign n4271 = ~n3874 & n4270;
  assign n4272 = n32724 & n4268;
  assign n4273 = ~n4155 & n4271;
  assign n4274 = ~n4269 & ~n32777;
  assign n4275 = n1812 & ~n4251;
  assign n4276 = n1812 & n4265;
  assign n4277 = ~n4264 & n4275;
  assign n4278 = ~n4274 & ~n32778;
  assign n4279 = ~n4266 & ~n4278;
  assign n4280 = ~n1582 & ~n4279;
  assign n4281 = n1582 & ~n4266;
  assign n4282 = ~n4278 & n4281;
  assign n4283 = ~n3891 & ~n32725;
  assign n4284 = ~n4155 & n4283;
  assign n4285 = ~n32726 & ~n4284;
  assign n4286 = ~n3891 & n32726;
  assign n4287 = ~n32725 & n4286;
  assign n4288 = n32726 & n4284;
  assign n4289 = ~n4155 & n4287;
  assign n4290 = n32726 & ~n4284;
  assign n4291 = ~n32726 & n4284;
  assign n4292 = ~n4290 & ~n4291;
  assign n4293 = ~n4285 & ~n32779;
  assign n4294 = ~n4282 & n32780;
  assign n4295 = ~n4280 & ~n4294;
  assign n4296 = ~n1388 & ~n4295;
  assign n4297 = ~n3907 & ~n3909;
  assign n4298 = ~n4155 & n4297;
  assign n4299 = ~n32728 & ~n4298;
  assign n4300 = ~n3909 & n32728;
  assign n4301 = ~n3907 & n4300;
  assign n4302 = n32728 & n4298;
  assign n4303 = ~n4155 & n4301;
  assign n4304 = ~n4299 & ~n32781;
  assign n4305 = n1388 & ~n4280;
  assign n4306 = n1388 & n4295;
  assign n4307 = ~n4294 & n4305;
  assign n4308 = ~n4304 & ~n32782;
  assign n4309 = ~n4296 & ~n4308;
  assign n4310 = ~n1192 & ~n4309;
  assign n4311 = n1192 & ~n4296;
  assign n4312 = ~n4308 & n4311;
  assign n4313 = ~n3924 & ~n32729;
  assign n4314 = ~n4155 & n4313;
  assign n4315 = n32731 & ~n4314;
  assign n4316 = ~n3924 & ~n32731;
  assign n4317 = ~n32729 & n4316;
  assign n4318 = ~n32731 & n4314;
  assign n4319 = ~n4155 & n4317;
  assign n4320 = n32731 & n4314;
  assign n4321 = ~n32731 & ~n4314;
  assign n4322 = ~n4320 & ~n4321;
  assign n4323 = ~n4315 & ~n32783;
  assign n4324 = ~n4312 & n32784;
  assign n4325 = ~n4310 & ~n4324;
  assign n4326 = ~n1028 & ~n4325;
  assign n4327 = ~n3941 & ~n3943;
  assign n4328 = ~n4155 & n4327;
  assign n4329 = ~n32733 & ~n4328;
  assign n4330 = ~n3943 & n32733;
  assign n4331 = ~n3941 & n4330;
  assign n4332 = n32733 & n4328;
  assign n4333 = ~n4155 & n4331;
  assign n4334 = ~n4329 & ~n32785;
  assign n4335 = n1028 & ~n4310;
  assign n4336 = n1028 & n4325;
  assign n4337 = ~n4324 & n4335;
  assign n4338 = ~n4334 & ~n32786;
  assign n4339 = ~n4326 & ~n4338;
  assign n4340 = ~n866 & ~n4339;
  assign n4341 = n866 & ~n4326;
  assign n4342 = ~n4338 & n4341;
  assign n4343 = ~n3958 & ~n32734;
  assign n4344 = ~n3958 & ~n4155;
  assign n4345 = ~n32734 & n4344;
  assign n4346 = ~n4155 & n4343;
  assign n4347 = ~n32736 & ~n32787;
  assign n4348 = n3973 & n4344;
  assign n4349 = n32736 & n32787;
  assign n4350 = ~n3958 & ~n32736;
  assign n4351 = ~n32734 & n4350;
  assign n4352 = ~n4155 & n4351;
  assign n4353 = n32736 & ~n32787;
  assign n4354 = ~n4352 & ~n4353;
  assign n4355 = ~n4347 & ~n32788;
  assign n4356 = ~n4342 & ~n32789;
  assign n4357 = ~n4340 & ~n4356;
  assign n4358 = ~n730 & ~n4357;
  assign n4359 = ~n3975 & ~n3977;
  assign n4360 = ~n4155 & n4359;
  assign n4361 = ~n32738 & ~n4360;
  assign n4362 = ~n3977 & n32738;
  assign n4363 = ~n3975 & n4362;
  assign n4364 = n32738 & n4360;
  assign n4365 = ~n4155 & n4363;
  assign n4366 = ~n4361 & ~n32790;
  assign n4367 = n730 & ~n4340;
  assign n4368 = n730 & n4357;
  assign n4369 = ~n4356 & n4367;
  assign n4370 = ~n4366 & ~n32791;
  assign n4371 = ~n4358 & ~n4370;
  assign n4372 = ~n602 & ~n4371;
  assign n4373 = n602 & ~n4358;
  assign n4374 = ~n4370 & n4373;
  assign n4375 = ~n3992 & ~n32739;
  assign n4376 = ~n3992 & ~n4155;
  assign n4377 = ~n32739 & n4376;
  assign n4378 = ~n4155 & n4375;
  assign n4379 = n4007 & n4376;
  assign n4380 = ~n32741 & n32792;
  assign n4381 = n32741 & ~n32792;
  assign n4382 = ~n3992 & n32741;
  assign n4383 = ~n32739 & n4382;
  assign n4384 = n32741 & n32792;
  assign n4385 = ~n4155 & n4383;
  assign n4386 = ~n32741 & ~n32792;
  assign n4387 = ~n32794 & ~n4386;
  assign n4388 = ~n32793 & ~n4381;
  assign n4389 = ~n4374 & ~n32795;
  assign n4390 = ~n4372 & ~n4389;
  assign n4391 = ~n497 & ~n4390;
  assign n4392 = ~n4009 & ~n4011;
  assign n4393 = ~n4155 & n4392;
  assign n4394 = ~n32743 & ~n4393;
  assign n4395 = ~n4011 & n32743;
  assign n4396 = ~n4009 & n4395;
  assign n4397 = n32743 & n4393;
  assign n4398 = ~n4155 & n4396;
  assign n4399 = ~n4394 & ~n32796;
  assign n4400 = n497 & ~n4372;
  assign n4401 = n497 & n4390;
  assign n4402 = ~n4389 & n4400;
  assign n4403 = ~n4399 & ~n32797;
  assign n4404 = ~n4391 & ~n4403;
  assign n4405 = ~n403 & ~n4404;
  assign n4406 = n403 & ~n4391;
  assign n4407 = ~n4403 & n4406;
  assign n4408 = ~n4026 & ~n32744;
  assign n4409 = ~n4026 & ~n4155;
  assign n4410 = ~n32744 & n4409;
  assign n4411 = ~n4155 & n4408;
  assign n4412 = n4037 & ~n32798;
  assign n4413 = n4038 & n4409;
  assign n4414 = ~n4037 & n32798;
  assign n4415 = ~n4026 & n4037;
  assign n4416 = ~n32744 & n4415;
  assign n4417 = ~n4155 & n4416;
  assign n4418 = ~n4037 & ~n32798;
  assign n4419 = ~n4417 & ~n4418;
  assign n4420 = ~n4412 & ~n32799;
  assign n4421 = ~n4407 & ~n32800;
  assign n4422 = ~n4405 & ~n4421;
  assign n4423 = ~n330 & ~n4422;
  assign n4424 = ~n4040 & ~n4042;
  assign n4425 = ~n4155 & n4424;
  assign n4426 = ~n32747 & ~n4425;
  assign n4427 = ~n4042 & n32747;
  assign n4428 = ~n4040 & n4427;
  assign n4429 = n32747 & n4425;
  assign n4430 = ~n4155 & n4428;
  assign n4431 = ~n4426 & ~n32801;
  assign n4432 = n330 & ~n4405;
  assign n4433 = n330 & n4422;
  assign n4434 = ~n4421 & n4432;
  assign n4435 = ~n4431 & ~n32802;
  assign n4436 = ~n4423 & ~n4435;
  assign n4437 = ~n271 & ~n4436;
  assign n4438 = n271 & ~n4423;
  assign n4439 = ~n4435 & n4438;
  assign n4440 = ~n4057 & ~n32748;
  assign n4441 = ~n4155 & n4440;
  assign n4442 = ~n32751 & n4441;
  assign n4443 = n32751 & ~n4441;
  assign n4444 = ~n4057 & n32751;
  assign n4445 = ~n32748 & n4444;
  assign n4446 = n32751 & n4441;
  assign n4447 = ~n4155 & n4445;
  assign n4448 = ~n32751 & ~n4441;
  assign n4449 = ~n32803 & ~n4448;
  assign n4450 = ~n4442 & ~n4443;
  assign n4451 = ~n4439 & ~n32804;
  assign n4452 = ~n4437 & ~n4451;
  assign n4453 = ~n217 & ~n4452;
  assign n4454 = ~n4076 & ~n4078;
  assign n4455 = ~n4155 & n4454;
  assign n4456 = ~n32753 & ~n4455;
  assign n4457 = ~n4078 & n32753;
  assign n4458 = ~n4076 & n4457;
  assign n4459 = n32753 & n4455;
  assign n4460 = ~n4155 & n4458;
  assign n4461 = ~n4456 & ~n32805;
  assign n4462 = n217 & ~n4437;
  assign n4463 = n217 & n4452;
  assign n4464 = ~n4451 & n4462;
  assign n4465 = ~n4461 & ~n32806;
  assign n4466 = ~n4453 & ~n4465;
  assign n4467 = ~n198 & ~n4466;
  assign n4468 = n198 & ~n4453;
  assign n4469 = ~n4465 & n4468;
  assign n4470 = ~n4093 & ~n32754;
  assign n4471 = ~n4093 & ~n4155;
  assign n4472 = ~n32754 & n4471;
  assign n4473 = ~n4155 & n4470;
  assign n4474 = n32756 & ~n32807;
  assign n4475 = n4108 & n4471;
  assign n4476 = ~n32756 & n32807;
  assign n4477 = ~n4093 & n32756;
  assign n4478 = ~n32754 & n4477;
  assign n4479 = ~n4155 & n4478;
  assign n4480 = ~n32756 & ~n32807;
  assign n4481 = ~n4479 & ~n4480;
  assign n4482 = ~n4474 & ~n32808;
  assign n4483 = ~n4469 & ~n32809;
  assign n4484 = ~n4467 & ~n4483;
  assign n4485 = ~n4110 & ~n4112;
  assign n4486 = ~n4155 & n4485;
  assign n4487 = ~n32758 & ~n4486;
  assign n4488 = ~n4112 & n32758;
  assign n4489 = ~n4110 & n4488;
  assign n4490 = n32758 & n4486;
  assign n4491 = ~n4155 & n4489;
  assign n4492 = ~n4487 & ~n32810;
  assign n4493 = ~n4126 & ~n32761;
  assign n4494 = ~n32761 & ~n4155;
  assign n4495 = ~n4126 & n4494;
  assign n4496 = ~n4155 & n4493;
  assign n4497 = ~n32763 & ~n32811;
  assign n4498 = ~n4492 & n4497;
  assign n4499 = ~n4484 & n4498;
  assign n4500 = n193 & ~n4499;
  assign n4501 = ~n4467 & n4492;
  assign n4502 = n4484 & n4492;
  assign n4503 = ~n4483 & n4501;
  assign n4504 = n4126 & ~n4494;
  assign n4505 = ~n193 & ~n4493;
  assign n4506 = ~n4504 & n4505;
  assign n4507 = ~n32812 & ~n4506;
  assign n4508 = ~n4500 & n4507;
  assign n4509 = pi80  & ~n4508;
  assign n4510 = ~pi78  & ~pi79 ;
  assign n4511 = ~pi80  & n4510;
  assign n4512 = ~n4509 & ~n4511;
  assign n4513 = ~n4155 & ~n4512;
  assign n4514 = ~pi80  & ~n4508;
  assign n4515 = pi81  & ~n4514;
  assign n4516 = ~pi81  & n4514;
  assign n4517 = n4157 & ~n4508;
  assign n4518 = ~n4515 & ~n32813;
  assign n4519 = ~n32709 & ~n32764;
  assign n4520 = ~n3767 & n4519;
  assign n4521 = ~n3786 & n4520;
  assign n4522 = ~n32711 & n4521;
  assign n4523 = n3772 & n3788;
  assign n4524 = ~n3780 & n4522;
  assign n4525 = ~n4511 & ~n32814;
  assign n4526 = ~n4153 & n4525;
  assign n4527 = ~n32763 & n4526;
  assign n4528 = ~n4147 & n4527;
  assign n4529 = n4155 & n4512;
  assign n4530 = ~n4509 & n4528;
  assign n4531 = n4518 & ~n32815;
  assign n4532 = ~n4513 & ~n4531;
  assign n4533 = ~n3788 & ~n4532;
  assign n4534 = n3788 & ~n4513;
  assign n4535 = ~n4531 & n4534;
  assign n4536 = ~n4155 & ~n4506;
  assign n4537 = ~n32812 & n4536;
  assign n4538 = ~n4500 & n4537;
  assign n4539 = ~n32813 & ~n4538;
  assign n4540 = pi82  & ~n4539;
  assign n4541 = ~pi82  & ~n4538;
  assign n4542 = ~pi82  & n4539;
  assign n4543 = ~n32813 & n4541;
  assign n4544 = ~n4540 & ~n32816;
  assign n4545 = ~n4535 & ~n4544;
  assign n4546 = ~n4533 & ~n4545;
  assign n4547 = ~n3473 & ~n4546;
  assign n4548 = n3473 & ~n4533;
  assign n4549 = ~n4545 & n4548;
  assign n4550 = n3473 & n4546;
  assign n4551 = ~n4160 & ~n32765;
  assign n4552 = ~n4508 & n4551;
  assign n4553 = n4177 & ~n4552;
  assign n4554 = ~n4177 & n4551;
  assign n4555 = ~n4177 & n4552;
  assign n4556 = ~n4508 & n4554;
  assign n4557 = ~n4553 & ~n32818;
  assign n4558 = ~n32817 & ~n4557;
  assign n4559 = ~n4547 & ~n4558;
  assign n4560 = ~n3140 & ~n4559;
  assign n4561 = n3140 & ~n4547;
  assign n4562 = ~n4558 & n4561;
  assign n4563 = ~n4180 & ~n32768;
  assign n4564 = ~n4180 & ~n4508;
  assign n4565 = ~n32768 & n4564;
  assign n4566 = ~n4508 & n4563;
  assign n4567 = n4189 & ~n32819;
  assign n4568 = n4193 & n4564;
  assign n4569 = n4189 & ~n32768;
  assign n4570 = ~n4180 & n4569;
  assign n4571 = ~n4508 & n4570;
  assign n4572 = ~n4189 & ~n32819;
  assign n4573 = ~n4571 & ~n4572;
  assign n4574 = ~n4567 & ~n4568;
  assign n4575 = ~n4562 & ~n32820;
  assign n4576 = ~n4560 & ~n4575;
  assign n4577 = ~n2855 & ~n4576;
  assign n4578 = n2855 & ~n4560;
  assign n4579 = ~n4575 & n4578;
  assign n4580 = n2855 & n4576;
  assign n4581 = ~n4195 & ~n4197;
  assign n4582 = ~n4508 & n4581;
  assign n4583 = n4204 & ~n4582;
  assign n4584 = ~n4204 & n4582;
  assign n4585 = ~n4195 & n4204;
  assign n4586 = ~n4197 & n4585;
  assign n4587 = n4204 & n4582;
  assign n4588 = ~n4508 & n4586;
  assign n4589 = ~n4204 & ~n4582;
  assign n4590 = ~n32822 & ~n4589;
  assign n4591 = ~n4583 & ~n4584;
  assign n4592 = ~n32821 & ~n32823;
  assign n4593 = ~n4577 & ~n4592;
  assign n4594 = ~n2556 & ~n4593;
  assign n4595 = n2556 & ~n4577;
  assign n4596 = ~n4592 & n4595;
  assign n4597 = ~n4207 & ~n32771;
  assign n4598 = ~n4207 & ~n4508;
  assign n4599 = ~n32771 & n4598;
  assign n4600 = ~n4508 & n4597;
  assign n4601 = n4215 & ~n32824;
  assign n4602 = n4219 & n4598;
  assign n4603 = n4215 & ~n32771;
  assign n4604 = ~n4207 & n4603;
  assign n4605 = ~n4508 & n4604;
  assign n4606 = ~n4215 & ~n32824;
  assign n4607 = ~n4605 & ~n4606;
  assign n4608 = ~n4601 & ~n4602;
  assign n4609 = ~n4596 & ~n32825;
  assign n4610 = ~n4594 & ~n4609;
  assign n4611 = ~n2301 & ~n4610;
  assign n4612 = n2301 & ~n4594;
  assign n4613 = ~n4609 & n4612;
  assign n4614 = n2301 & n4610;
  assign n4615 = ~n4221 & ~n4223;
  assign n4616 = ~n4508 & n4615;
  assign n4617 = ~n32773 & n4616;
  assign n4618 = n32773 & ~n4616;
  assign n4619 = ~n4221 & n32773;
  assign n4620 = ~n4223 & n4619;
  assign n4621 = ~n4508 & n4620;
  assign n4622 = ~n32773 & ~n4616;
  assign n4623 = ~n4621 & ~n4622;
  assign n4624 = ~n4617 & ~n4618;
  assign n4625 = ~n32826 & ~n32827;
  assign n4626 = ~n4611 & ~n4625;
  assign n4627 = ~n2038 & ~n4626;
  assign n4628 = n2038 & ~n4611;
  assign n4629 = ~n4625 & n4628;
  assign n4630 = ~n4237 & ~n32775;
  assign n4631 = ~n4237 & ~n4508;
  assign n4632 = ~n32775 & n4631;
  assign n4633 = ~n4508 & n4630;
  assign n4634 = n4245 & ~n32828;
  assign n4635 = n4249 & n4631;
  assign n4636 = n4245 & ~n32775;
  assign n4637 = ~n4237 & n4636;
  assign n4638 = ~n4508 & n4637;
  assign n4639 = ~n4245 & ~n32828;
  assign n4640 = ~n4638 & ~n4639;
  assign n4641 = ~n4634 & ~n4635;
  assign n4642 = ~n4629 & ~n32829;
  assign n4643 = ~n4627 & ~n4642;
  assign n4644 = ~n1812 & ~n4643;
  assign n4645 = n1812 & ~n4627;
  assign n4646 = ~n4642 & n4645;
  assign n4647 = n1812 & n4643;
  assign n4648 = ~n4251 & ~n4253;
  assign n4649 = ~n4508 & n4648;
  assign n4650 = ~n32776 & ~n4649;
  assign n4651 = ~n4251 & n32776;
  assign n4652 = ~n4253 & n4651;
  assign n4653 = n32776 & n4649;
  assign n4654 = ~n4508 & n4652;
  assign n4655 = n32776 & ~n4649;
  assign n4656 = ~n32776 & n4649;
  assign n4657 = ~n4655 & ~n4656;
  assign n4658 = ~n4650 & ~n32831;
  assign n4659 = ~n32830 & n32832;
  assign n4660 = ~n4644 & ~n4659;
  assign n4661 = ~n1582 & ~n4660;
  assign n4662 = n1582 & ~n4644;
  assign n4663 = ~n4659 & n4662;
  assign n4664 = ~n4266 & ~n32778;
  assign n4665 = ~n4266 & ~n4508;
  assign n4666 = ~n32778 & n4665;
  assign n4667 = ~n4508 & n4664;
  assign n4668 = n4274 & ~n32833;
  assign n4669 = n4278 & n4665;
  assign n4670 = n4274 & ~n32778;
  assign n4671 = ~n4266 & n4670;
  assign n4672 = ~n4508 & n4671;
  assign n4673 = ~n4274 & ~n32833;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = ~n4668 & ~n4669;
  assign n4676 = ~n4663 & ~n32834;
  assign n4677 = ~n4661 & ~n4676;
  assign n4678 = ~n1388 & ~n4677;
  assign n4679 = n1388 & ~n4661;
  assign n4680 = ~n4676 & n4679;
  assign n4681 = n1388 & n4677;
  assign n4682 = ~n4280 & ~n4282;
  assign n4683 = ~n4508 & n4682;
  assign n4684 = n32780 & ~n4683;
  assign n4685 = ~n4280 & ~n32780;
  assign n4686 = ~n4282 & n4685;
  assign n4687 = ~n32780 & n4683;
  assign n4688 = ~n4508 & n4686;
  assign n4689 = n32780 & n4683;
  assign n4690 = ~n32780 & ~n4683;
  assign n4691 = ~n4689 & ~n4690;
  assign n4692 = ~n4684 & ~n32836;
  assign n4693 = ~n32835 & n32837;
  assign n4694 = ~n4678 & ~n4693;
  assign n4695 = ~n1192 & ~n4694;
  assign n4696 = n1192 & ~n4678;
  assign n4697 = ~n4693 & n4696;
  assign n4698 = ~n4296 & ~n32782;
  assign n4699 = ~n4296 & ~n4508;
  assign n4700 = ~n32782 & n4699;
  assign n4701 = ~n4508 & n4698;
  assign n4702 = n4304 & ~n32838;
  assign n4703 = n4308 & n4699;
  assign n4704 = n4304 & ~n32782;
  assign n4705 = ~n4296 & n4704;
  assign n4706 = ~n4508 & n4705;
  assign n4707 = ~n4304 & ~n32838;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = ~n4702 & ~n4703;
  assign n4710 = ~n4697 & ~n32839;
  assign n4711 = ~n4695 & ~n4710;
  assign n4712 = ~n1028 & ~n4711;
  assign n4713 = n1028 & ~n4695;
  assign n4714 = ~n4710 & n4713;
  assign n4715 = n1028 & n4711;
  assign n4716 = ~n4310 & ~n4312;
  assign n4717 = ~n4310 & ~n4508;
  assign n4718 = ~n4312 & n4717;
  assign n4719 = ~n4508 & n4716;
  assign n4720 = ~n32784 & ~n32841;
  assign n4721 = n4324 & n4717;
  assign n4722 = n32784 & n32841;
  assign n4723 = ~n4310 & ~n32784;
  assign n4724 = ~n4312 & n4723;
  assign n4725 = ~n4508 & n4724;
  assign n4726 = n32784 & ~n32841;
  assign n4727 = ~n4725 & ~n4726;
  assign n4728 = ~n4720 & ~n32842;
  assign n4729 = ~n32840 & ~n32843;
  assign n4730 = ~n4712 & ~n4729;
  assign n4731 = ~n866 & ~n4730;
  assign n4732 = n866 & ~n4712;
  assign n4733 = ~n4729 & n4732;
  assign n4734 = ~n4326 & ~n32786;
  assign n4735 = ~n4326 & ~n4508;
  assign n4736 = ~n32786 & n4735;
  assign n4737 = ~n4508 & n4734;
  assign n4738 = n4334 & ~n32844;
  assign n4739 = n4338 & n4735;
  assign n4740 = n4334 & ~n32786;
  assign n4741 = ~n4326 & n4740;
  assign n4742 = ~n4508 & n4741;
  assign n4743 = ~n4334 & ~n32844;
  assign n4744 = ~n4742 & ~n4743;
  assign n4745 = ~n4738 & ~n4739;
  assign n4746 = ~n4733 & ~n32845;
  assign n4747 = ~n4731 & ~n4746;
  assign n4748 = ~n730 & ~n4747;
  assign n4749 = n730 & ~n4731;
  assign n4750 = ~n4746 & n4749;
  assign n4751 = n730 & n4747;
  assign n4752 = ~n4340 & ~n4342;
  assign n4753 = ~n4508 & n4752;
  assign n4754 = ~n32789 & ~n4753;
  assign n4755 = ~n4340 & n32789;
  assign n4756 = ~n4342 & n4755;
  assign n4757 = n32789 & n4753;
  assign n4758 = ~n4508 & n4756;
  assign n4759 = ~n4754 & ~n32847;
  assign n4760 = ~n32846 & ~n4759;
  assign n4761 = ~n4748 & ~n4760;
  assign n4762 = ~n602 & ~n4761;
  assign n4763 = n602 & ~n4748;
  assign n4764 = ~n4760 & n4763;
  assign n4765 = ~n4358 & ~n32791;
  assign n4766 = ~n4358 & ~n4508;
  assign n4767 = ~n32791 & n4766;
  assign n4768 = ~n4508 & n4765;
  assign n4769 = n4366 & ~n32848;
  assign n4770 = n4370 & n4766;
  assign n4771 = n4366 & ~n32791;
  assign n4772 = ~n4358 & n4771;
  assign n4773 = ~n4508 & n4772;
  assign n4774 = ~n4366 & ~n32848;
  assign n4775 = ~n4773 & ~n4774;
  assign n4776 = ~n4769 & ~n4770;
  assign n4777 = ~n4764 & ~n32849;
  assign n4778 = ~n4762 & ~n4777;
  assign n4779 = ~n497 & ~n4778;
  assign n4780 = ~n4372 & ~n4374;
  assign n4781 = ~n4508 & n4780;
  assign n4782 = ~n32795 & ~n4781;
  assign n4783 = ~n4372 & n32795;
  assign n4784 = ~n4374 & n4783;
  assign n4785 = n32795 & n4781;
  assign n4786 = ~n4508 & n4784;
  assign n4787 = ~n4782 & ~n32850;
  assign n4788 = n497 & ~n4762;
  assign n4789 = ~n4777 & n4788;
  assign n4790 = n497 & n4778;
  assign n4791 = ~n4787 & ~n32851;
  assign n4792 = ~n4779 & ~n4791;
  assign n4793 = ~n403 & ~n4792;
  assign n4794 = n403 & ~n4779;
  assign n4795 = ~n4791 & n4794;
  assign n4796 = ~n4391 & ~n32797;
  assign n4797 = ~n4391 & ~n4508;
  assign n4798 = ~n32797 & n4797;
  assign n4799 = ~n4508 & n4796;
  assign n4800 = n4399 & ~n32852;
  assign n4801 = n4403 & n4797;
  assign n4802 = n4399 & ~n32797;
  assign n4803 = ~n4391 & n4802;
  assign n4804 = ~n4508 & n4803;
  assign n4805 = ~n4399 & ~n32852;
  assign n4806 = ~n4804 & ~n4805;
  assign n4807 = ~n4800 & ~n4801;
  assign n4808 = ~n4795 & ~n32853;
  assign n4809 = ~n4793 & ~n4808;
  assign n4810 = ~n330 & ~n4809;
  assign n4811 = n330 & ~n4793;
  assign n4812 = ~n4808 & n4811;
  assign n4813 = n330 & n4809;
  assign n4814 = ~n4405 & ~n4407;
  assign n4815 = ~n4508 & n4814;
  assign n4816 = ~n32800 & n4815;
  assign n4817 = n32800 & ~n4815;
  assign n4818 = ~n4405 & n32800;
  assign n4819 = ~n4407 & n4818;
  assign n4820 = n32800 & n4815;
  assign n4821 = ~n4508 & n4819;
  assign n4822 = ~n32800 & ~n4815;
  assign n4823 = ~n32855 & ~n4822;
  assign n4824 = ~n4816 & ~n4817;
  assign n4825 = ~n32854 & ~n32856;
  assign n4826 = ~n4810 & ~n4825;
  assign n4827 = ~n271 & ~n4826;
  assign n4828 = n271 & ~n4810;
  assign n4829 = ~n4825 & n4828;
  assign n4830 = ~n4423 & ~n32802;
  assign n4831 = ~n4423 & ~n4508;
  assign n4832 = ~n32802 & n4831;
  assign n4833 = ~n4508 & n4830;
  assign n4834 = n4431 & ~n32857;
  assign n4835 = n4435 & n4831;
  assign n4836 = n4431 & ~n32802;
  assign n4837 = ~n4423 & n4836;
  assign n4838 = ~n4508 & n4837;
  assign n4839 = ~n4431 & ~n32857;
  assign n4840 = ~n4838 & ~n4839;
  assign n4841 = ~n4834 & ~n4835;
  assign n4842 = ~n4829 & ~n32858;
  assign n4843 = ~n4827 & ~n4842;
  assign n4844 = ~n217 & ~n4843;
  assign n4845 = n217 & ~n4827;
  assign n4846 = ~n4842 & n4845;
  assign n4847 = n217 & n4843;
  assign n4848 = ~n4437 & ~n4439;
  assign n4849 = ~n4437 & ~n4508;
  assign n4850 = ~n4439 & n4849;
  assign n4851 = ~n4508 & n4848;
  assign n4852 = n32804 & ~n32860;
  assign n4853 = n4451 & n4849;
  assign n4854 = ~n32804 & n32860;
  assign n4855 = ~n4437 & n32804;
  assign n4856 = ~n4439 & n4855;
  assign n4857 = ~n4508 & n4856;
  assign n4858 = ~n32804 & ~n32860;
  assign n4859 = ~n4857 & ~n4858;
  assign n4860 = ~n4852 & ~n32861;
  assign n4861 = ~n32859 & ~n32862;
  assign n4862 = ~n4844 & ~n4861;
  assign n4863 = ~n198 & ~n4862;
  assign n4864 = n198 & ~n4844;
  assign n4865 = ~n4861 & n4864;
  assign n4866 = ~n4453 & ~n32806;
  assign n4867 = ~n4453 & ~n4508;
  assign n4868 = ~n32806 & n4867;
  assign n4869 = ~n4508 & n4866;
  assign n4870 = n4461 & ~n32863;
  assign n4871 = n4465 & n4867;
  assign n4872 = n4461 & ~n32806;
  assign n4873 = ~n4453 & n4872;
  assign n4874 = ~n4508 & n4873;
  assign n4875 = ~n4461 & ~n32863;
  assign n4876 = ~n4874 & ~n4875;
  assign n4877 = ~n4870 & ~n4871;
  assign n4878 = ~n4865 & ~n32864;
  assign n4879 = ~n4863 & ~n4878;
  assign n4880 = ~n4467 & ~n4469;
  assign n4881 = ~n4508 & n4880;
  assign n4882 = ~n32809 & ~n4881;
  assign n4883 = ~n4467 & n32809;
  assign n4884 = ~n4469 & n4883;
  assign n4885 = n32809 & n4881;
  assign n4886 = ~n4508 & n4884;
  assign n4887 = ~n4882 & ~n32865;
  assign n4888 = ~n4484 & ~n4492;
  assign n4889 = ~n4492 & ~n4508;
  assign n4890 = ~n4484 & n4889;
  assign n4891 = ~n4508 & n4888;
  assign n4892 = ~n32812 & ~n32866;
  assign n4893 = ~n4887 & n4892;
  assign n4894 = ~n4879 & n4893;
  assign n4895 = n193 & ~n4894;
  assign n4896 = ~n4863 & n4887;
  assign n4897 = ~n4878 & n4896;
  assign n4898 = n4879 & n4887;
  assign n4899 = n4484 & ~n4889;
  assign n4900 = ~n193 & ~n4888;
  assign n4901 = ~n4899 & n4900;
  assign n4902 = ~n32867 & ~n4901;
  assign n4903 = ~n4895 & n4902;
  assign n4904 = pi78  & ~n4903;
  assign n4905 = ~pi76  & ~pi77 ;
  assign n4906 = ~pi78  & n4905;
  assign n4907 = ~n4904 & ~n4906;
  assign n4908 = ~n4508 & ~n4907;
  assign n4909 = ~n4136 & ~n32814;
  assign n4910 = ~n4137 & n4909;
  assign n4911 = ~n4153 & n4910;
  assign n4912 = ~n32763 & n4911;
  assign n4913 = n32761 & n4155;
  assign n4914 = ~n4147 & n4912;
  assign n4915 = ~n4906 & ~n32868;
  assign n4916 = ~n4506 & n4915;
  assign n4917 = ~n32812 & n4916;
  assign n4918 = ~n4500 & n4917;
  assign n4919 = n4508 & n4907;
  assign n4920 = ~n4904 & n4918;
  assign n4921 = ~pi78  & ~n4903;
  assign n4922 = pi79  & ~n4921;
  assign n4923 = ~pi79  & n4921;
  assign n4924 = n4510 & ~n4903;
  assign n4925 = ~n4922 & ~n32870;
  assign n4926 = ~n32869 & n4925;
  assign n4927 = ~n4908 & ~n4926;
  assign n4928 = ~n4155 & ~n4927;
  assign n4929 = ~n4508 & ~n4901;
  assign n4930 = ~n32867 & n4929;
  assign n4931 = ~n4895 & n4930;
  assign n4932 = ~n32870 & ~n4931;
  assign n4933 = pi80  & ~n4932;
  assign n4934 = ~pi80  & ~n4931;
  assign n4935 = ~pi80  & n4932;
  assign n4936 = ~n32870 & n4934;
  assign n4937 = ~n4933 & ~n32871;
  assign n4938 = n4155 & ~n4908;
  assign n4939 = n4155 & n4927;
  assign n4940 = ~n4926 & n4938;
  assign n4941 = ~n4937 & ~n32872;
  assign n4942 = ~n4928 & ~n4941;
  assign n4943 = ~n3788 & ~n4942;
  assign n4944 = n3788 & ~n4928;
  assign n4945 = ~n4941 & n4944;
  assign n4946 = ~n4513 & ~n32815;
  assign n4947 = ~n4903 & n4946;
  assign n4948 = n4518 & ~n4947;
  assign n4949 = ~n4518 & n4946;
  assign n4950 = ~n4518 & n4947;
  assign n4951 = ~n4903 & n4949;
  assign n4952 = ~n4948 & ~n32873;
  assign n4953 = ~n4945 & ~n4952;
  assign n4954 = ~n4943 & ~n4953;
  assign n4955 = ~n3473 & ~n4954;
  assign n4956 = ~n4533 & ~n4535;
  assign n4957 = ~n4903 & n4956;
  assign n4958 = ~n4544 & ~n4957;
  assign n4959 = ~n4535 & n4544;
  assign n4960 = ~n4533 & n4959;
  assign n4961 = n4544 & n4957;
  assign n4962 = ~n4903 & n4960;
  assign n4963 = ~n4958 & ~n32874;
  assign n4964 = n3473 & ~n4943;
  assign n4965 = n3473 & n4954;
  assign n4966 = ~n4953 & n4964;
  assign n4967 = ~n4963 & ~n32875;
  assign n4968 = ~n4955 & ~n4967;
  assign n4969 = ~n3140 & ~n4968;
  assign n4970 = n3140 & ~n4955;
  assign n4971 = ~n4967 & n4970;
  assign n4972 = ~n4547 & ~n32817;
  assign n4973 = ~n4903 & n4972;
  assign n4974 = n4557 & ~n4973;
  assign n4975 = ~n4557 & n4973;
  assign n4976 = ~n4547 & n4557;
  assign n4977 = ~n32817 & n4976;
  assign n4978 = n4557 & n4973;
  assign n4979 = ~n4903 & n4977;
  assign n4980 = ~n4557 & ~n4973;
  assign n4981 = ~n32876 & ~n4980;
  assign n4982 = ~n4974 & ~n4975;
  assign n4983 = ~n4971 & ~n32877;
  assign n4984 = ~n4969 & ~n4983;
  assign n4985 = ~n2855 & ~n4984;
  assign n4986 = ~n4560 & ~n4562;
  assign n4987 = ~n4903 & n4986;
  assign n4988 = ~n32820 & ~n4987;
  assign n4989 = ~n4562 & n32820;
  assign n4990 = ~n4560 & n4989;
  assign n4991 = n32820 & n4987;
  assign n4992 = ~n4903 & n4990;
  assign n4993 = ~n4988 & ~n32878;
  assign n4994 = n2855 & ~n4969;
  assign n4995 = n2855 & n4984;
  assign n4996 = ~n4983 & n4994;
  assign n4997 = ~n4993 & ~n32879;
  assign n4998 = ~n4985 & ~n4997;
  assign n4999 = ~n2556 & ~n4998;
  assign n5000 = n2556 & ~n4985;
  assign n5001 = ~n4997 & n5000;
  assign n5002 = ~n4577 & ~n32821;
  assign n5003 = ~n4903 & n5002;
  assign n5004 = ~n32823 & n5003;
  assign n5005 = n32823 & ~n5003;
  assign n5006 = ~n4577 & n32823;
  assign n5007 = ~n32821 & n5006;
  assign n5008 = ~n4903 & n5007;
  assign n5009 = ~n32823 & ~n5003;
  assign n5010 = ~n5008 & ~n5009;
  assign n5011 = ~n5004 & ~n5005;
  assign n5012 = ~n5001 & ~n32880;
  assign n5013 = ~n4999 & ~n5012;
  assign n5014 = ~n2301 & ~n5013;
  assign n5015 = ~n4594 & ~n4596;
  assign n5016 = ~n4903 & n5015;
  assign n5017 = ~n32825 & ~n5016;
  assign n5018 = ~n4596 & n32825;
  assign n5019 = ~n4594 & n5018;
  assign n5020 = n32825 & n5016;
  assign n5021 = ~n4903 & n5019;
  assign n5022 = ~n5017 & ~n32881;
  assign n5023 = n2301 & ~n4999;
  assign n5024 = n2301 & n5013;
  assign n5025 = ~n5012 & n5023;
  assign n5026 = ~n5022 & ~n32882;
  assign n5027 = ~n5014 & ~n5026;
  assign n5028 = ~n2038 & ~n5027;
  assign n5029 = n2038 & ~n5014;
  assign n5030 = ~n5026 & n5029;
  assign n5031 = ~n4611 & ~n32826;
  assign n5032 = ~n4903 & n5031;
  assign n5033 = ~n32827 & ~n5032;
  assign n5034 = ~n4611 & n32827;
  assign n5035 = ~n32826 & n5034;
  assign n5036 = n32827 & n5032;
  assign n5037 = ~n4903 & n5035;
  assign n5038 = n32827 & ~n5032;
  assign n5039 = ~n32827 & n5032;
  assign n5040 = ~n5038 & ~n5039;
  assign n5041 = ~n5033 & ~n32883;
  assign n5042 = ~n5030 & n32884;
  assign n5043 = ~n5028 & ~n5042;
  assign n5044 = ~n1812 & ~n5043;
  assign n5045 = ~n4627 & ~n4629;
  assign n5046 = ~n4903 & n5045;
  assign n5047 = ~n32829 & ~n5046;
  assign n5048 = ~n4629 & n32829;
  assign n5049 = ~n4627 & n5048;
  assign n5050 = n32829 & n5046;
  assign n5051 = ~n4903 & n5049;
  assign n5052 = ~n5047 & ~n32885;
  assign n5053 = n1812 & ~n5028;
  assign n5054 = n1812 & n5043;
  assign n5055 = ~n5042 & n5053;
  assign n5056 = ~n5052 & ~n32886;
  assign n5057 = ~n5044 & ~n5056;
  assign n5058 = ~n1582 & ~n5057;
  assign n5059 = n1582 & ~n5044;
  assign n5060 = ~n5056 & n5059;
  assign n5061 = ~n4644 & ~n32830;
  assign n5062 = ~n4903 & n5061;
  assign n5063 = n32832 & ~n5062;
  assign n5064 = ~n4644 & ~n32832;
  assign n5065 = ~n32830 & n5064;
  assign n5066 = ~n32832 & n5062;
  assign n5067 = ~n4903 & n5065;
  assign n5068 = n32832 & n5062;
  assign n5069 = ~n32832 & ~n5062;
  assign n5070 = ~n5068 & ~n5069;
  assign n5071 = ~n5063 & ~n32887;
  assign n5072 = ~n5060 & n32888;
  assign n5073 = ~n5058 & ~n5072;
  assign n5074 = ~n1388 & ~n5073;
  assign n5075 = ~n4661 & ~n4663;
  assign n5076 = ~n4903 & n5075;
  assign n5077 = ~n32834 & ~n5076;
  assign n5078 = ~n4663 & n32834;
  assign n5079 = ~n4661 & n5078;
  assign n5080 = n32834 & n5076;
  assign n5081 = ~n4903 & n5079;
  assign n5082 = ~n5077 & ~n32889;
  assign n5083 = n1388 & ~n5058;
  assign n5084 = n1388 & n5073;
  assign n5085 = ~n5072 & n5083;
  assign n5086 = ~n5082 & ~n32890;
  assign n5087 = ~n5074 & ~n5086;
  assign n5088 = ~n1192 & ~n5087;
  assign n5089 = n1192 & ~n5074;
  assign n5090 = ~n5086 & n5089;
  assign n5091 = ~n4678 & ~n32835;
  assign n5092 = ~n4678 & ~n4903;
  assign n5093 = ~n32835 & n5092;
  assign n5094 = ~n4903 & n5091;
  assign n5095 = ~n32837 & ~n32891;
  assign n5096 = n4693 & n5092;
  assign n5097 = n32837 & n32891;
  assign n5098 = ~n4678 & ~n32837;
  assign n5099 = ~n32835 & n5098;
  assign n5100 = ~n4903 & n5099;
  assign n5101 = n32837 & ~n32891;
  assign n5102 = ~n5100 & ~n5101;
  assign n5103 = ~n5095 & ~n32892;
  assign n5104 = ~n5090 & ~n32893;
  assign n5105 = ~n5088 & ~n5104;
  assign n5106 = ~n1028 & ~n5105;
  assign n5107 = ~n4695 & ~n4697;
  assign n5108 = ~n4903 & n5107;
  assign n5109 = ~n32839 & ~n5108;
  assign n5110 = ~n4697 & n32839;
  assign n5111 = ~n4695 & n5110;
  assign n5112 = n32839 & n5108;
  assign n5113 = ~n4903 & n5111;
  assign n5114 = ~n5109 & ~n32894;
  assign n5115 = n1028 & ~n5088;
  assign n5116 = n1028 & n5105;
  assign n5117 = ~n5104 & n5115;
  assign n5118 = ~n5114 & ~n32895;
  assign n5119 = ~n5106 & ~n5118;
  assign n5120 = ~n866 & ~n5119;
  assign n5121 = n866 & ~n5106;
  assign n5122 = ~n5118 & n5121;
  assign n5123 = ~n4712 & ~n32840;
  assign n5124 = ~n4903 & n5123;
  assign n5125 = ~n32843 & ~n5124;
  assign n5126 = ~n4712 & n32843;
  assign n5127 = ~n32840 & n5126;
  assign n5128 = n32843 & n5124;
  assign n5129 = ~n4903 & n5127;
  assign n5130 = ~n5125 & ~n32896;
  assign n5131 = ~n5122 & ~n5130;
  assign n5132 = ~n5120 & ~n5131;
  assign n5133 = ~n730 & ~n5132;
  assign n5134 = ~n4731 & ~n4733;
  assign n5135 = ~n4903 & n5134;
  assign n5136 = ~n32845 & ~n5135;
  assign n5137 = ~n4733 & n32845;
  assign n5138 = ~n4731 & n5137;
  assign n5139 = n32845 & n5135;
  assign n5140 = ~n4903 & n5138;
  assign n5141 = ~n5136 & ~n32897;
  assign n5142 = n730 & ~n5120;
  assign n5143 = n730 & n5132;
  assign n5144 = ~n5131 & n5142;
  assign n5145 = ~n5141 & ~n32898;
  assign n5146 = ~n5133 & ~n5145;
  assign n5147 = ~n602 & ~n5146;
  assign n5148 = n602 & ~n5133;
  assign n5149 = ~n5145 & n5148;
  assign n5150 = ~n4748 & ~n32846;
  assign n5151 = ~n4748 & ~n4903;
  assign n5152 = ~n32846 & n5151;
  assign n5153 = ~n4903 & n5150;
  assign n5154 = n4759 & ~n32899;
  assign n5155 = n4760 & n5151;
  assign n5156 = ~n4759 & n32899;
  assign n5157 = ~n4748 & n4759;
  assign n5158 = ~n32846 & n5157;
  assign n5159 = ~n4903 & n5158;
  assign n5160 = ~n4759 & ~n32899;
  assign n5161 = ~n5159 & ~n5160;
  assign n5162 = ~n5154 & ~n32900;
  assign n5163 = ~n5149 & ~n32901;
  assign n5164 = ~n5147 & ~n5163;
  assign n5165 = ~n497 & ~n5164;
  assign n5166 = ~n4762 & ~n4764;
  assign n5167 = ~n4903 & n5166;
  assign n5168 = ~n32849 & ~n5167;
  assign n5169 = ~n4764 & n32849;
  assign n5170 = ~n4762 & n5169;
  assign n5171 = n32849 & n5167;
  assign n5172 = ~n4903 & n5170;
  assign n5173 = ~n5168 & ~n32902;
  assign n5174 = n497 & ~n5147;
  assign n5175 = n497 & n5164;
  assign n5176 = ~n5163 & n5174;
  assign n5177 = ~n5173 & ~n32903;
  assign n5178 = ~n5165 & ~n5177;
  assign n5179 = ~n403 & ~n5178;
  assign n5180 = n403 & ~n5165;
  assign n5181 = ~n5177 & n5180;
  assign n5182 = ~n4779 & ~n32851;
  assign n5183 = ~n4779 & ~n4903;
  assign n5184 = ~n32851 & n5183;
  assign n5185 = ~n4903 & n5182;
  assign n5186 = n4787 & ~n32904;
  assign n5187 = n4791 & n5183;
  assign n5188 = ~n4779 & n4787;
  assign n5189 = ~n32851 & n5188;
  assign n5190 = ~n4903 & n5189;
  assign n5191 = ~n4787 & ~n32904;
  assign n5192 = ~n5190 & ~n5191;
  assign n5193 = ~n5186 & ~n5187;
  assign n5194 = ~n5181 & ~n32905;
  assign n5195 = ~n5179 & ~n5194;
  assign n5196 = ~n330 & ~n5195;
  assign n5197 = ~n4793 & ~n4795;
  assign n5198 = ~n4903 & n5197;
  assign n5199 = ~n32853 & ~n5198;
  assign n5200 = ~n4795 & n32853;
  assign n5201 = ~n4793 & n5200;
  assign n5202 = n32853 & n5198;
  assign n5203 = ~n4903 & n5201;
  assign n5204 = ~n5199 & ~n32906;
  assign n5205 = n330 & ~n5179;
  assign n5206 = n330 & n5195;
  assign n5207 = ~n5194 & n5205;
  assign n5208 = ~n5204 & ~n32907;
  assign n5209 = ~n5196 & ~n5208;
  assign n5210 = ~n271 & ~n5209;
  assign n5211 = n271 & ~n5196;
  assign n5212 = ~n5208 & n5211;
  assign n5213 = ~n4810 & ~n32854;
  assign n5214 = ~n4810 & ~n4903;
  assign n5215 = ~n32854 & n5214;
  assign n5216 = ~n4903 & n5213;
  assign n5217 = n32856 & ~n32908;
  assign n5218 = n4825 & n5214;
  assign n5219 = ~n32856 & n32908;
  assign n5220 = ~n4810 & n32856;
  assign n5221 = ~n32854 & n5220;
  assign n5222 = ~n4903 & n5221;
  assign n5223 = ~n32856 & ~n32908;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = ~n5217 & ~n32909;
  assign n5226 = ~n5212 & ~n32910;
  assign n5227 = ~n5210 & ~n5226;
  assign n5228 = ~n217 & ~n5227;
  assign n5229 = ~n4827 & ~n4829;
  assign n5230 = ~n4903 & n5229;
  assign n5231 = ~n32858 & ~n5230;
  assign n5232 = ~n4829 & n32858;
  assign n5233 = ~n4827 & n5232;
  assign n5234 = n32858 & n5230;
  assign n5235 = ~n4903 & n5233;
  assign n5236 = ~n5231 & ~n32911;
  assign n5237 = n217 & ~n5210;
  assign n5238 = n217 & n5227;
  assign n5239 = ~n5226 & n5237;
  assign n5240 = ~n5236 & ~n32912;
  assign n5241 = ~n5228 & ~n5240;
  assign n5242 = ~n198 & ~n5241;
  assign n5243 = ~n4844 & ~n32859;
  assign n5244 = ~n4903 & n5243;
  assign n5245 = ~n32862 & ~n5244;
  assign n5246 = ~n4844 & n32862;
  assign n5247 = ~n32859 & n5246;
  assign n5248 = n32862 & n5244;
  assign n5249 = ~n4903 & n5247;
  assign n5250 = ~n5245 & ~n32913;
  assign n5251 = n198 & ~n5228;
  assign n5252 = ~n5240 & n5251;
  assign n5253 = ~n5250 & ~n5252;
  assign n5254 = ~n5242 & ~n5253;
  assign n5255 = ~n4863 & ~n4865;
  assign n5256 = ~n4903 & n5255;
  assign n5257 = ~n32864 & ~n5256;
  assign n5258 = ~n4865 & n32864;
  assign n5259 = ~n4863 & n5258;
  assign n5260 = n32864 & n5256;
  assign n5261 = ~n4903 & n5259;
  assign n5262 = ~n5257 & ~n32914;
  assign n5263 = ~n4879 & ~n4887;
  assign n5264 = ~n4887 & ~n4903;
  assign n5265 = ~n4879 & n5264;
  assign n5266 = ~n4903 & n5263;
  assign n5267 = ~n32867 & ~n32915;
  assign n5268 = ~n5262 & n5267;
  assign n5269 = ~n5254 & n5268;
  assign n5270 = n193 & ~n5269;
  assign n5271 = ~n5242 & n5262;
  assign n5272 = n5254 & n5262;
  assign n5273 = ~n5253 & n5271;
  assign n5274 = n4879 & ~n5264;
  assign n5275 = ~n193 & ~n5263;
  assign n5276 = ~n5274 & n5275;
  assign n5277 = ~n32916 & ~n5276;
  assign n5278 = ~n5270 & n5277;
  assign n5279 = pi76  & ~n5278;
  assign n5280 = ~pi74  & ~pi75 ;
  assign n5281 = ~pi76  & n5280;
  assign n5282 = ~n5279 & ~n5281;
  assign n5283 = ~n4903 & ~n5282;
  assign n5284 = ~pi76  & ~n5278;
  assign n5285 = pi77  & ~n5284;
  assign n5286 = ~pi77  & n5284;
  assign n5287 = n4905 & ~n5278;
  assign n5288 = ~n5285 & ~n32917;
  assign n5289 = ~n32810 & ~n32868;
  assign n5290 = ~n4487 & n5289;
  assign n5291 = ~n4506 & n5290;
  assign n5292 = ~n32812 & n5291;
  assign n5293 = n4492 & n4508;
  assign n5294 = ~n4500 & n5292;
  assign n5295 = ~n5281 & ~n32918;
  assign n5296 = ~n4901 & n5295;
  assign n5297 = ~n32867 & n5296;
  assign n5298 = ~n4895 & n5297;
  assign n5299 = n4903 & n5282;
  assign n5300 = ~n5279 & n5298;
  assign n5301 = n5288 & ~n32919;
  assign n5302 = ~n5283 & ~n5301;
  assign n5303 = ~n4508 & ~n5302;
  assign n5304 = n4508 & ~n5283;
  assign n5305 = ~n5301 & n5304;
  assign n5306 = ~n4903 & ~n5276;
  assign n5307 = ~n32916 & n5306;
  assign n5308 = ~n5270 & n5307;
  assign n5309 = ~n32917 & ~n5308;
  assign n5310 = pi78  & ~n5309;
  assign n5311 = ~pi78  & ~n5308;
  assign n5312 = ~pi78  & n5309;
  assign n5313 = ~n32917 & n5311;
  assign n5314 = ~n5310 & ~n32920;
  assign n5315 = ~n5305 & ~n5314;
  assign n5316 = ~n5303 & ~n5315;
  assign n5317 = ~n4155 & ~n5316;
  assign n5318 = n4155 & ~n5303;
  assign n5319 = ~n5315 & n5318;
  assign n5320 = n4155 & n5316;
  assign n5321 = ~n4908 & ~n32869;
  assign n5322 = ~n5278 & n5321;
  assign n5323 = n4925 & ~n5322;
  assign n5324 = ~n4925 & n5321;
  assign n5325 = ~n4925 & n5322;
  assign n5326 = ~n5278 & n5324;
  assign n5327 = ~n5323 & ~n32922;
  assign n5328 = ~n32921 & ~n5327;
  assign n5329 = ~n5317 & ~n5328;
  assign n5330 = ~n3788 & ~n5329;
  assign n5331 = n3788 & ~n5317;
  assign n5332 = ~n5328 & n5331;
  assign n5333 = ~n4928 & ~n32872;
  assign n5334 = ~n4928 & ~n5278;
  assign n5335 = ~n32872 & n5334;
  assign n5336 = ~n5278 & n5333;
  assign n5337 = n4937 & ~n32923;
  assign n5338 = n4941 & n5334;
  assign n5339 = n4937 & ~n32872;
  assign n5340 = ~n4928 & n5339;
  assign n5341 = ~n5278 & n5340;
  assign n5342 = ~n4937 & ~n32923;
  assign n5343 = ~n5341 & ~n5342;
  assign n5344 = ~n5337 & ~n5338;
  assign n5345 = ~n5332 & ~n32924;
  assign n5346 = ~n5330 & ~n5345;
  assign n5347 = ~n3473 & ~n5346;
  assign n5348 = n3473 & ~n5330;
  assign n5349 = ~n5345 & n5348;
  assign n5350 = n3473 & n5346;
  assign n5351 = ~n4943 & ~n4945;
  assign n5352 = ~n5278 & n5351;
  assign n5353 = n4952 & ~n5352;
  assign n5354 = ~n4952 & n5352;
  assign n5355 = ~n4943 & n4952;
  assign n5356 = ~n4945 & n5355;
  assign n5357 = n4952 & n5352;
  assign n5358 = ~n5278 & n5356;
  assign n5359 = ~n4952 & ~n5352;
  assign n5360 = ~n32926 & ~n5359;
  assign n5361 = ~n5353 & ~n5354;
  assign n5362 = ~n32925 & ~n32927;
  assign n5363 = ~n5347 & ~n5362;
  assign n5364 = ~n3140 & ~n5363;
  assign n5365 = n3140 & ~n5347;
  assign n5366 = ~n5362 & n5365;
  assign n5367 = ~n4955 & ~n32875;
  assign n5368 = ~n4955 & ~n5278;
  assign n5369 = ~n32875 & n5368;
  assign n5370 = ~n5278 & n5367;
  assign n5371 = n4963 & ~n32928;
  assign n5372 = n4967 & n5368;
  assign n5373 = n4963 & ~n32875;
  assign n5374 = ~n4955 & n5373;
  assign n5375 = ~n5278 & n5374;
  assign n5376 = ~n4963 & ~n32928;
  assign n5377 = ~n5375 & ~n5376;
  assign n5378 = ~n5371 & ~n5372;
  assign n5379 = ~n5366 & ~n32929;
  assign n5380 = ~n5364 & ~n5379;
  assign n5381 = ~n2855 & ~n5380;
  assign n5382 = n2855 & ~n5364;
  assign n5383 = ~n5379 & n5382;
  assign n5384 = n2855 & n5380;
  assign n5385 = ~n4969 & ~n4971;
  assign n5386 = ~n5278 & n5385;
  assign n5387 = ~n32877 & n5386;
  assign n5388 = n32877 & ~n5386;
  assign n5389 = ~n4969 & n32877;
  assign n5390 = ~n4971 & n5389;
  assign n5391 = ~n5278 & n5390;
  assign n5392 = ~n32877 & ~n5386;
  assign n5393 = ~n5391 & ~n5392;
  assign n5394 = ~n5387 & ~n5388;
  assign n5395 = ~n32930 & ~n32931;
  assign n5396 = ~n5381 & ~n5395;
  assign n5397 = ~n2556 & ~n5396;
  assign n5398 = n2556 & ~n5381;
  assign n5399 = ~n5395 & n5398;
  assign n5400 = ~n4985 & ~n32879;
  assign n5401 = ~n4985 & ~n5278;
  assign n5402 = ~n32879 & n5401;
  assign n5403 = ~n5278 & n5400;
  assign n5404 = n4993 & ~n32932;
  assign n5405 = n4997 & n5401;
  assign n5406 = n4993 & ~n32879;
  assign n5407 = ~n4985 & n5406;
  assign n5408 = ~n5278 & n5407;
  assign n5409 = ~n4993 & ~n32932;
  assign n5410 = ~n5408 & ~n5409;
  assign n5411 = ~n5404 & ~n5405;
  assign n5412 = ~n5399 & ~n32933;
  assign n5413 = ~n5397 & ~n5412;
  assign n5414 = ~n2301 & ~n5413;
  assign n5415 = n2301 & ~n5397;
  assign n5416 = ~n5412 & n5415;
  assign n5417 = n2301 & n5413;
  assign n5418 = ~n4999 & ~n5001;
  assign n5419 = ~n5278 & n5418;
  assign n5420 = ~n32880 & ~n5419;
  assign n5421 = ~n4999 & n32880;
  assign n5422 = ~n5001 & n5421;
  assign n5423 = n32880 & n5419;
  assign n5424 = ~n5278 & n5422;
  assign n5425 = n32880 & ~n5419;
  assign n5426 = ~n32880 & n5419;
  assign n5427 = ~n5425 & ~n5426;
  assign n5428 = ~n5420 & ~n32935;
  assign n5429 = ~n32934 & n32936;
  assign n5430 = ~n5414 & ~n5429;
  assign n5431 = ~n2038 & ~n5430;
  assign n5432 = n2038 & ~n5414;
  assign n5433 = ~n5429 & n5432;
  assign n5434 = ~n5014 & ~n32882;
  assign n5435 = ~n5014 & ~n5278;
  assign n5436 = ~n32882 & n5435;
  assign n5437 = ~n5278 & n5434;
  assign n5438 = n5022 & ~n32937;
  assign n5439 = n5026 & n5435;
  assign n5440 = n5022 & ~n32882;
  assign n5441 = ~n5014 & n5440;
  assign n5442 = ~n5278 & n5441;
  assign n5443 = ~n5022 & ~n32937;
  assign n5444 = ~n5442 & ~n5443;
  assign n5445 = ~n5438 & ~n5439;
  assign n5446 = ~n5433 & ~n32938;
  assign n5447 = ~n5431 & ~n5446;
  assign n5448 = ~n1812 & ~n5447;
  assign n5449 = n1812 & ~n5431;
  assign n5450 = ~n5446 & n5449;
  assign n5451 = n1812 & n5447;
  assign n5452 = ~n5028 & ~n5030;
  assign n5453 = ~n5278 & n5452;
  assign n5454 = n32884 & ~n5453;
  assign n5455 = ~n5028 & ~n32884;
  assign n5456 = ~n5030 & n5455;
  assign n5457 = ~n32884 & n5453;
  assign n5458 = ~n5278 & n5456;
  assign n5459 = n32884 & n5453;
  assign n5460 = ~n32884 & ~n5453;
  assign n5461 = ~n5459 & ~n5460;
  assign n5462 = ~n5454 & ~n32940;
  assign n5463 = ~n32939 & n32941;
  assign n5464 = ~n5448 & ~n5463;
  assign n5465 = ~n1582 & ~n5464;
  assign n5466 = n1582 & ~n5448;
  assign n5467 = ~n5463 & n5466;
  assign n5468 = ~n5044 & ~n32886;
  assign n5469 = ~n5044 & ~n5278;
  assign n5470 = ~n32886 & n5469;
  assign n5471 = ~n5278 & n5468;
  assign n5472 = n5052 & ~n32942;
  assign n5473 = n5056 & n5469;
  assign n5474 = n5052 & ~n32886;
  assign n5475 = ~n5044 & n5474;
  assign n5476 = ~n5278 & n5475;
  assign n5477 = ~n5052 & ~n32942;
  assign n5478 = ~n5476 & ~n5477;
  assign n5479 = ~n5472 & ~n5473;
  assign n5480 = ~n5467 & ~n32943;
  assign n5481 = ~n5465 & ~n5480;
  assign n5482 = ~n1388 & ~n5481;
  assign n5483 = n1388 & ~n5465;
  assign n5484 = ~n5480 & n5483;
  assign n5485 = n1388 & n5481;
  assign n5486 = ~n5058 & ~n5060;
  assign n5487 = ~n5058 & ~n5278;
  assign n5488 = ~n5060 & n5487;
  assign n5489 = ~n5278 & n5486;
  assign n5490 = ~n32888 & ~n32945;
  assign n5491 = n5072 & n5487;
  assign n5492 = n32888 & n32945;
  assign n5493 = ~n5058 & ~n32888;
  assign n5494 = ~n5060 & n5493;
  assign n5495 = ~n5278 & n5494;
  assign n5496 = n32888 & ~n32945;
  assign n5497 = ~n5495 & ~n5496;
  assign n5498 = ~n5490 & ~n32946;
  assign n5499 = ~n32944 & ~n32947;
  assign n5500 = ~n5482 & ~n5499;
  assign n5501 = ~n1192 & ~n5500;
  assign n5502 = n1192 & ~n5482;
  assign n5503 = ~n5499 & n5502;
  assign n5504 = ~n5074 & ~n32890;
  assign n5505 = ~n5074 & ~n5278;
  assign n5506 = ~n32890 & n5505;
  assign n5507 = ~n5278 & n5504;
  assign n5508 = n5082 & ~n32948;
  assign n5509 = n5086 & n5505;
  assign n5510 = n5082 & ~n32890;
  assign n5511 = ~n5074 & n5510;
  assign n5512 = ~n5278 & n5511;
  assign n5513 = ~n5082 & ~n32948;
  assign n5514 = ~n5512 & ~n5513;
  assign n5515 = ~n5508 & ~n5509;
  assign n5516 = ~n5503 & ~n32949;
  assign n5517 = ~n5501 & ~n5516;
  assign n5518 = ~n1028 & ~n5517;
  assign n5519 = n1028 & ~n5501;
  assign n5520 = ~n5516 & n5519;
  assign n5521 = n1028 & n5517;
  assign n5522 = ~n5088 & ~n5090;
  assign n5523 = ~n5278 & n5522;
  assign n5524 = ~n32893 & ~n5523;
  assign n5525 = ~n5088 & n32893;
  assign n5526 = ~n5090 & n5525;
  assign n5527 = n32893 & n5523;
  assign n5528 = ~n5278 & n5526;
  assign n5529 = ~n5524 & ~n32951;
  assign n5530 = ~n32950 & ~n5529;
  assign n5531 = ~n5518 & ~n5530;
  assign n5532 = ~n866 & ~n5531;
  assign n5533 = n866 & ~n5518;
  assign n5534 = ~n5530 & n5533;
  assign n5535 = ~n5106 & ~n32895;
  assign n5536 = ~n5106 & ~n5278;
  assign n5537 = ~n32895 & n5536;
  assign n5538 = ~n5278 & n5535;
  assign n5539 = n5114 & ~n32952;
  assign n5540 = n5118 & n5536;
  assign n5541 = n5114 & ~n32895;
  assign n5542 = ~n5106 & n5541;
  assign n5543 = ~n5278 & n5542;
  assign n5544 = ~n5114 & ~n32952;
  assign n5545 = ~n5543 & ~n5544;
  assign n5546 = ~n5539 & ~n5540;
  assign n5547 = ~n5534 & ~n32953;
  assign n5548 = ~n5532 & ~n5547;
  assign n5549 = ~n730 & ~n5548;
  assign n5550 = n730 & ~n5532;
  assign n5551 = ~n5547 & n5550;
  assign n5552 = n730 & n5548;
  assign n5553 = ~n5120 & ~n5122;
  assign n5554 = ~n5120 & ~n5278;
  assign n5555 = ~n5122 & n5554;
  assign n5556 = ~n5278 & n5553;
  assign n5557 = n5130 & ~n32955;
  assign n5558 = n5131 & n5554;
  assign n5559 = ~n5130 & n32955;
  assign n5560 = ~n5120 & n5130;
  assign n5561 = ~n5122 & n5560;
  assign n5562 = ~n5278 & n5561;
  assign n5563 = ~n5130 & ~n32955;
  assign n5564 = ~n5562 & ~n5563;
  assign n5565 = ~n5557 & ~n32956;
  assign n5566 = ~n32954 & ~n32957;
  assign n5567 = ~n5549 & ~n5566;
  assign n5568 = ~n602 & ~n5567;
  assign n5569 = n602 & ~n5549;
  assign n5570 = ~n5566 & n5569;
  assign n5571 = ~n5133 & ~n32898;
  assign n5572 = ~n5133 & ~n5278;
  assign n5573 = ~n32898 & n5572;
  assign n5574 = ~n5278 & n5571;
  assign n5575 = n5141 & ~n32958;
  assign n5576 = n5145 & n5572;
  assign n5577 = n5141 & ~n32898;
  assign n5578 = ~n5133 & n5577;
  assign n5579 = ~n5278 & n5578;
  assign n5580 = ~n5141 & ~n32958;
  assign n5581 = ~n5579 & ~n5580;
  assign n5582 = ~n5575 & ~n5576;
  assign n5583 = ~n5570 & ~n32959;
  assign n5584 = ~n5568 & ~n5583;
  assign n5585 = ~n497 & ~n5584;
  assign n5586 = n497 & ~n5568;
  assign n5587 = ~n5583 & n5586;
  assign n5588 = n497 & n5584;
  assign n5589 = ~n5147 & ~n5149;
  assign n5590 = ~n5278 & n5589;
  assign n5591 = ~n32901 & n5590;
  assign n5592 = n32901 & ~n5590;
  assign n5593 = ~n5147 & n32901;
  assign n5594 = ~n5149 & n5593;
  assign n5595 = n32901 & n5590;
  assign n5596 = ~n5278 & n5594;
  assign n5597 = ~n32901 & ~n5590;
  assign n5598 = ~n32961 & ~n5597;
  assign n5599 = ~n5591 & ~n5592;
  assign n5600 = ~n32960 & ~n32962;
  assign n5601 = ~n5585 & ~n5600;
  assign n5602 = ~n403 & ~n5601;
  assign n5603 = n403 & ~n5585;
  assign n5604 = ~n5600 & n5603;
  assign n5605 = ~n5165 & ~n32903;
  assign n5606 = ~n5165 & ~n5278;
  assign n5607 = ~n32903 & n5606;
  assign n5608 = ~n5278 & n5605;
  assign n5609 = n5173 & ~n32963;
  assign n5610 = n5177 & n5606;
  assign n5611 = n5173 & ~n32903;
  assign n5612 = ~n5165 & n5611;
  assign n5613 = ~n5278 & n5612;
  assign n5614 = ~n5173 & ~n32963;
  assign n5615 = ~n5613 & ~n5614;
  assign n5616 = ~n5609 & ~n5610;
  assign n5617 = ~n5604 & ~n32964;
  assign n5618 = ~n5602 & ~n5617;
  assign n5619 = ~n330 & ~n5618;
  assign n5620 = ~n5179 & ~n5181;
  assign n5621 = ~n5278 & n5620;
  assign n5622 = ~n32905 & ~n5621;
  assign n5623 = ~n5179 & n32905;
  assign n5624 = ~n5181 & n5623;
  assign n5625 = n32905 & n5621;
  assign n5626 = ~n5278 & n5624;
  assign n5627 = ~n5622 & ~n32965;
  assign n5628 = n330 & ~n5602;
  assign n5629 = ~n5617 & n5628;
  assign n5630 = n330 & n5618;
  assign n5631 = ~n5627 & ~n32966;
  assign n5632 = ~n5619 & ~n5631;
  assign n5633 = ~n271 & ~n5632;
  assign n5634 = n271 & ~n5619;
  assign n5635 = ~n5631 & n5634;
  assign n5636 = ~n5196 & ~n32907;
  assign n5637 = ~n5196 & ~n5278;
  assign n5638 = ~n32907 & n5637;
  assign n5639 = ~n5278 & n5636;
  assign n5640 = n5204 & ~n32967;
  assign n5641 = n5208 & n5637;
  assign n5642 = n5204 & ~n32907;
  assign n5643 = ~n5196 & n5642;
  assign n5644 = ~n5278 & n5643;
  assign n5645 = ~n5204 & ~n32967;
  assign n5646 = ~n5644 & ~n5645;
  assign n5647 = ~n5640 & ~n5641;
  assign n5648 = ~n5635 & ~n32968;
  assign n5649 = ~n5633 & ~n5648;
  assign n5650 = ~n217 & ~n5649;
  assign n5651 = ~n5210 & ~n5212;
  assign n5652 = ~n5278 & n5651;
  assign n5653 = ~n32910 & ~n5652;
  assign n5654 = ~n5210 & n32910;
  assign n5655 = ~n5212 & n5654;
  assign n5656 = n32910 & n5652;
  assign n5657 = ~n5278 & n5655;
  assign n5658 = ~n5653 & ~n32969;
  assign n5659 = n217 & ~n5633;
  assign n5660 = ~n5648 & n5659;
  assign n5661 = n217 & n5649;
  assign n5662 = ~n5658 & ~n32970;
  assign n5663 = ~n5650 & ~n5662;
  assign n5664 = ~n198 & ~n5663;
  assign n5665 = n198 & ~n5650;
  assign n5666 = ~n5662 & n5665;
  assign n5667 = ~n5228 & ~n32912;
  assign n5668 = ~n5228 & ~n5278;
  assign n5669 = ~n32912 & n5668;
  assign n5670 = ~n5278 & n5667;
  assign n5671 = n5236 & ~n32971;
  assign n5672 = n5240 & n5668;
  assign n5673 = n5236 & ~n32912;
  assign n5674 = ~n5228 & n5673;
  assign n5675 = ~n5278 & n5674;
  assign n5676 = ~n5236 & ~n32971;
  assign n5677 = ~n5675 & ~n5676;
  assign n5678 = ~n5671 & ~n5672;
  assign n5679 = ~n5666 & ~n32972;
  assign n5680 = ~n5664 & ~n5679;
  assign n5681 = ~n5242 & ~n5252;
  assign n5682 = ~n5242 & ~n5278;
  assign n5683 = ~n5252 & n5682;
  assign n5684 = ~n5278 & n5681;
  assign n5685 = n5250 & ~n32973;
  assign n5686 = n5253 & n5682;
  assign n5687 = ~n5242 & n5250;
  assign n5688 = ~n5252 & n5687;
  assign n5689 = ~n5278 & n5688;
  assign n5690 = ~n5250 & ~n32973;
  assign n5691 = ~n5689 & ~n5690;
  assign n5692 = ~n5685 & ~n5686;
  assign n5693 = ~n5254 & ~n5262;
  assign n5694 = ~n5262 & ~n5278;
  assign n5695 = ~n5254 & n5694;
  assign n5696 = ~n5278 & n5693;
  assign n5697 = ~n32916 & ~n32975;
  assign n5698 = ~n32974 & n5697;
  assign n5699 = ~n5680 & n5698;
  assign n5700 = n193 & ~n5699;
  assign n5701 = ~n5664 & n32974;
  assign n5702 = ~n5679 & n5701;
  assign n5703 = n5680 & n32974;
  assign n5704 = n5254 & ~n5694;
  assign n5705 = ~n193 & ~n5693;
  assign n5706 = ~n5704 & n5705;
  assign n5707 = ~n32976 & ~n5706;
  assign n5708 = ~n5700 & n5707;
  assign n5709 = pi74  & ~n5708;
  assign n5710 = ~pi72  & ~pi73 ;
  assign n5711 = ~pi74  & n5710;
  assign n5712 = ~n5709 & ~n5711;
  assign n5713 = ~n5278 & ~n5712;
  assign n5714 = ~n32865 & ~n32918;
  assign n5715 = ~n4882 & n5714;
  assign n5716 = ~n4901 & n5715;
  assign n5717 = ~n32867 & n5716;
  assign n5718 = n4887 & n4903;
  assign n5719 = ~n4895 & n5717;
  assign n5720 = ~n5711 & ~n32977;
  assign n5721 = ~n5276 & n5720;
  assign n5722 = ~n32916 & n5721;
  assign n5723 = ~n5270 & n5722;
  assign n5724 = n5278 & n5712;
  assign n5725 = ~n5709 & n5723;
  assign n5726 = ~pi74  & ~n5708;
  assign n5727 = pi75  & ~n5726;
  assign n5728 = ~pi75  & n5726;
  assign n5729 = n5280 & ~n5708;
  assign n5730 = ~n5727 & ~n32979;
  assign n5731 = ~n32978 & n5730;
  assign n5732 = ~n5713 & ~n5731;
  assign n5733 = ~n4903 & ~n5732;
  assign n5734 = ~n5278 & ~n5706;
  assign n5735 = ~n32976 & n5734;
  assign n5736 = ~n5700 & n5735;
  assign n5737 = ~n32979 & ~n5736;
  assign n5738 = pi76  & ~n5737;
  assign n5739 = ~pi76  & ~n5736;
  assign n5740 = ~pi76  & n5737;
  assign n5741 = ~n32979 & n5739;
  assign n5742 = ~n5738 & ~n32980;
  assign n5743 = n4903 & ~n5713;
  assign n5744 = n4903 & n5732;
  assign n5745 = ~n5731 & n5743;
  assign n5746 = ~n5742 & ~n32981;
  assign n5747 = ~n5733 & ~n5746;
  assign n5748 = ~n4508 & ~n5747;
  assign n5749 = n4508 & ~n5733;
  assign n5750 = ~n5746 & n5749;
  assign n5751 = ~n5283 & ~n32919;
  assign n5752 = ~n5708 & n5751;
  assign n5753 = n5288 & ~n5752;
  assign n5754 = ~n5288 & n5751;
  assign n5755 = ~n5288 & n5752;
  assign n5756 = ~n5708 & n5754;
  assign n5757 = ~n5753 & ~n32982;
  assign n5758 = ~n5750 & ~n5757;
  assign n5759 = ~n5748 & ~n5758;
  assign n5760 = ~n4155 & ~n5759;
  assign n5761 = ~n5303 & ~n5305;
  assign n5762 = ~n5708 & n5761;
  assign n5763 = ~n5314 & ~n5762;
  assign n5764 = ~n5305 & n5314;
  assign n5765 = ~n5303 & n5764;
  assign n5766 = n5314 & n5762;
  assign n5767 = ~n5708 & n5765;
  assign n5768 = ~n5763 & ~n32983;
  assign n5769 = n4155 & ~n5748;
  assign n5770 = n4155 & n5759;
  assign n5771 = ~n5758 & n5769;
  assign n5772 = ~n5768 & ~n32984;
  assign n5773 = ~n5760 & ~n5772;
  assign n5774 = ~n3788 & ~n5773;
  assign n5775 = n3788 & ~n5760;
  assign n5776 = ~n5772 & n5775;
  assign n5777 = ~n5317 & ~n32921;
  assign n5778 = ~n5708 & n5777;
  assign n5779 = n5327 & ~n5778;
  assign n5780 = ~n5327 & n5778;
  assign n5781 = ~n5317 & n5327;
  assign n5782 = ~n32921 & n5781;
  assign n5783 = n5327 & n5778;
  assign n5784 = ~n5708 & n5782;
  assign n5785 = ~n5327 & ~n5778;
  assign n5786 = ~n32985 & ~n5785;
  assign n5787 = ~n5779 & ~n5780;
  assign n5788 = ~n5776 & ~n32986;
  assign n5789 = ~n5774 & ~n5788;
  assign n5790 = ~n3473 & ~n5789;
  assign n5791 = ~n5330 & ~n5332;
  assign n5792 = ~n5708 & n5791;
  assign n5793 = ~n32924 & ~n5792;
  assign n5794 = ~n5332 & n32924;
  assign n5795 = ~n5330 & n5794;
  assign n5796 = n32924 & n5792;
  assign n5797 = ~n5708 & n5795;
  assign n5798 = ~n5793 & ~n32987;
  assign n5799 = n3473 & ~n5774;
  assign n5800 = n3473 & n5789;
  assign n5801 = ~n5788 & n5799;
  assign n5802 = ~n5798 & ~n32988;
  assign n5803 = ~n5790 & ~n5802;
  assign n5804 = ~n3140 & ~n5803;
  assign n5805 = n3140 & ~n5790;
  assign n5806 = ~n5802 & n5805;
  assign n5807 = ~n5347 & ~n32925;
  assign n5808 = ~n5708 & n5807;
  assign n5809 = ~n32927 & n5808;
  assign n5810 = n32927 & ~n5808;
  assign n5811 = ~n5347 & n32927;
  assign n5812 = ~n32925 & n5811;
  assign n5813 = ~n5708 & n5812;
  assign n5814 = ~n32927 & ~n5808;
  assign n5815 = ~n5813 & ~n5814;
  assign n5816 = ~n5809 & ~n5810;
  assign n5817 = ~n5806 & ~n32989;
  assign n5818 = ~n5804 & ~n5817;
  assign n5819 = ~n2855 & ~n5818;
  assign n5820 = ~n5364 & ~n5366;
  assign n5821 = ~n5708 & n5820;
  assign n5822 = ~n32929 & ~n5821;
  assign n5823 = ~n5366 & n32929;
  assign n5824 = ~n5364 & n5823;
  assign n5825 = n32929 & n5821;
  assign n5826 = ~n5708 & n5824;
  assign n5827 = ~n5822 & ~n32990;
  assign n5828 = n2855 & ~n5804;
  assign n5829 = n2855 & n5818;
  assign n5830 = ~n5817 & n5828;
  assign n5831 = ~n5827 & ~n32991;
  assign n5832 = ~n5819 & ~n5831;
  assign n5833 = ~n2556 & ~n5832;
  assign n5834 = n2556 & ~n5819;
  assign n5835 = ~n5831 & n5834;
  assign n5836 = ~n5381 & ~n32930;
  assign n5837 = ~n5708 & n5836;
  assign n5838 = ~n32931 & ~n5837;
  assign n5839 = ~n5381 & n32931;
  assign n5840 = ~n32930 & n5839;
  assign n5841 = n32931 & n5837;
  assign n5842 = ~n5708 & n5840;
  assign n5843 = n32931 & ~n5837;
  assign n5844 = ~n32931 & n5837;
  assign n5845 = ~n5843 & ~n5844;
  assign n5846 = ~n5838 & ~n32992;
  assign n5847 = ~n5835 & n32993;
  assign n5848 = ~n5833 & ~n5847;
  assign n5849 = ~n2301 & ~n5848;
  assign n5850 = ~n5397 & ~n5399;
  assign n5851 = ~n5708 & n5850;
  assign n5852 = ~n32933 & ~n5851;
  assign n5853 = ~n5399 & n32933;
  assign n5854 = ~n5397 & n5853;
  assign n5855 = n32933 & n5851;
  assign n5856 = ~n5708 & n5854;
  assign n5857 = ~n5852 & ~n32994;
  assign n5858 = n2301 & ~n5833;
  assign n5859 = n2301 & n5848;
  assign n5860 = ~n5847 & n5858;
  assign n5861 = ~n5857 & ~n32995;
  assign n5862 = ~n5849 & ~n5861;
  assign n5863 = ~n2038 & ~n5862;
  assign n5864 = n2038 & ~n5849;
  assign n5865 = ~n5861 & n5864;
  assign n5866 = ~n5414 & ~n32934;
  assign n5867 = ~n5708 & n5866;
  assign n5868 = n32936 & ~n5867;
  assign n5869 = ~n5414 & ~n32936;
  assign n5870 = ~n32934 & n5869;
  assign n5871 = ~n32936 & n5867;
  assign n5872 = ~n5708 & n5870;
  assign n5873 = n32936 & n5867;
  assign n5874 = ~n32936 & ~n5867;
  assign n5875 = ~n5873 & ~n5874;
  assign n5876 = ~n5868 & ~n32996;
  assign n5877 = ~n5865 & n32997;
  assign n5878 = ~n5863 & ~n5877;
  assign n5879 = ~n1812 & ~n5878;
  assign n5880 = ~n5431 & ~n5433;
  assign n5881 = ~n5708 & n5880;
  assign n5882 = ~n32938 & ~n5881;
  assign n5883 = ~n5433 & n32938;
  assign n5884 = ~n5431 & n5883;
  assign n5885 = n32938 & n5881;
  assign n5886 = ~n5708 & n5884;
  assign n5887 = ~n5882 & ~n32998;
  assign n5888 = n1812 & ~n5863;
  assign n5889 = n1812 & n5878;
  assign n5890 = ~n5877 & n5888;
  assign n5891 = ~n5887 & ~n32999;
  assign n5892 = ~n5879 & ~n5891;
  assign n5893 = ~n1582 & ~n5892;
  assign n5894 = n1582 & ~n5879;
  assign n5895 = ~n5891 & n5894;
  assign n5896 = ~n5448 & ~n32939;
  assign n5897 = ~n5448 & ~n5708;
  assign n5898 = ~n32939 & n5897;
  assign n5899 = ~n5708 & n5896;
  assign n5900 = ~n32941 & ~n33000;
  assign n5901 = n5463 & n5897;
  assign n5902 = n32941 & n33000;
  assign n5903 = ~n5448 & ~n32941;
  assign n5904 = ~n32939 & n5903;
  assign n5905 = ~n5708 & n5904;
  assign n5906 = n32941 & ~n33000;
  assign n5907 = ~n5905 & ~n5906;
  assign n5908 = ~n5900 & ~n33001;
  assign n5909 = ~n5895 & ~n33002;
  assign n5910 = ~n5893 & ~n5909;
  assign n5911 = ~n1388 & ~n5910;
  assign n5912 = ~n5465 & ~n5467;
  assign n5913 = ~n5708 & n5912;
  assign n5914 = ~n32943 & ~n5913;
  assign n5915 = ~n5467 & n32943;
  assign n5916 = ~n5465 & n5915;
  assign n5917 = n32943 & n5913;
  assign n5918 = ~n5708 & n5916;
  assign n5919 = ~n5914 & ~n33003;
  assign n5920 = n1388 & ~n5893;
  assign n5921 = n1388 & n5910;
  assign n5922 = ~n5909 & n5920;
  assign n5923 = ~n5919 & ~n33004;
  assign n5924 = ~n5911 & ~n5923;
  assign n5925 = ~n1192 & ~n5924;
  assign n5926 = n1192 & ~n5911;
  assign n5927 = ~n5923 & n5926;
  assign n5928 = ~n5482 & ~n32944;
  assign n5929 = ~n5708 & n5928;
  assign n5930 = ~n32947 & ~n5929;
  assign n5931 = ~n5482 & n32947;
  assign n5932 = ~n32944 & n5931;
  assign n5933 = n32947 & n5929;
  assign n5934 = ~n5708 & n5932;
  assign n5935 = ~n5930 & ~n33005;
  assign n5936 = ~n5927 & ~n5935;
  assign n5937 = ~n5925 & ~n5936;
  assign n5938 = ~n1028 & ~n5937;
  assign n5939 = ~n5501 & ~n5503;
  assign n5940 = ~n5708 & n5939;
  assign n5941 = ~n32949 & ~n5940;
  assign n5942 = ~n5503 & n32949;
  assign n5943 = ~n5501 & n5942;
  assign n5944 = n32949 & n5940;
  assign n5945 = ~n5708 & n5943;
  assign n5946 = ~n5941 & ~n33006;
  assign n5947 = n1028 & ~n5925;
  assign n5948 = n1028 & n5937;
  assign n5949 = ~n5936 & n5947;
  assign n5950 = ~n5946 & ~n33007;
  assign n5951 = ~n5938 & ~n5950;
  assign n5952 = ~n866 & ~n5951;
  assign n5953 = n866 & ~n5938;
  assign n5954 = ~n5950 & n5953;
  assign n5955 = ~n5518 & ~n32950;
  assign n5956 = ~n5518 & ~n5708;
  assign n5957 = ~n32950 & n5956;
  assign n5958 = ~n5708 & n5955;
  assign n5959 = n5529 & ~n33008;
  assign n5960 = n5530 & n5956;
  assign n5961 = ~n5529 & n33008;
  assign n5962 = ~n5518 & n5529;
  assign n5963 = ~n32950 & n5962;
  assign n5964 = ~n5708 & n5963;
  assign n5965 = ~n5529 & ~n33008;
  assign n5966 = ~n5964 & ~n5965;
  assign n5967 = ~n5959 & ~n33009;
  assign n5968 = ~n5954 & ~n33010;
  assign n5969 = ~n5952 & ~n5968;
  assign n5970 = ~n730 & ~n5969;
  assign n5971 = ~n5532 & ~n5534;
  assign n5972 = ~n5708 & n5971;
  assign n5973 = ~n32953 & ~n5972;
  assign n5974 = ~n5534 & n32953;
  assign n5975 = ~n5532 & n5974;
  assign n5976 = n32953 & n5972;
  assign n5977 = ~n5708 & n5975;
  assign n5978 = ~n5973 & ~n33011;
  assign n5979 = n730 & ~n5952;
  assign n5980 = n730 & n5969;
  assign n5981 = ~n5968 & n5979;
  assign n5982 = ~n5978 & ~n33012;
  assign n5983 = ~n5970 & ~n5982;
  assign n5984 = ~n602 & ~n5983;
  assign n5985 = n602 & ~n5970;
  assign n5986 = ~n5982 & n5985;
  assign n5987 = ~n5549 & ~n32954;
  assign n5988 = ~n5708 & n5987;
  assign n5989 = ~n32957 & n5988;
  assign n5990 = n32957 & ~n5988;
  assign n5991 = ~n5549 & n32957;
  assign n5992 = ~n32954 & n5991;
  assign n5993 = n32957 & n5988;
  assign n5994 = ~n5708 & n5992;
  assign n5995 = ~n32957 & ~n5988;
  assign n5996 = ~n33013 & ~n5995;
  assign n5997 = ~n5989 & ~n5990;
  assign n5998 = ~n5986 & ~n33014;
  assign n5999 = ~n5984 & ~n5998;
  assign n6000 = ~n497 & ~n5999;
  assign n6001 = ~n5568 & ~n5570;
  assign n6002 = ~n5708 & n6001;
  assign n6003 = ~n32959 & ~n6002;
  assign n6004 = ~n5570 & n32959;
  assign n6005 = ~n5568 & n6004;
  assign n6006 = n32959 & n6002;
  assign n6007 = ~n5708 & n6005;
  assign n6008 = ~n6003 & ~n33015;
  assign n6009 = n497 & ~n5984;
  assign n6010 = n497 & n5999;
  assign n6011 = ~n5998 & n6009;
  assign n6012 = ~n6008 & ~n33016;
  assign n6013 = ~n6000 & ~n6012;
  assign n6014 = ~n403 & ~n6013;
  assign n6015 = n403 & ~n6000;
  assign n6016 = ~n6012 & n6015;
  assign n6017 = ~n5585 & ~n32960;
  assign n6018 = ~n5585 & ~n5708;
  assign n6019 = ~n32960 & n6018;
  assign n6020 = ~n5708 & n6017;
  assign n6021 = n32962 & ~n33017;
  assign n6022 = n5600 & n6018;
  assign n6023 = ~n32962 & n33017;
  assign n6024 = ~n5585 & n32962;
  assign n6025 = ~n32960 & n6024;
  assign n6026 = ~n5708 & n6025;
  assign n6027 = ~n32962 & ~n33017;
  assign n6028 = ~n6026 & ~n6027;
  assign n6029 = ~n6021 & ~n33018;
  assign n6030 = ~n6016 & ~n33019;
  assign n6031 = ~n6014 & ~n6030;
  assign n6032 = ~n330 & ~n6031;
  assign n6033 = ~n5602 & ~n5604;
  assign n6034 = ~n5708 & n6033;
  assign n6035 = ~n32964 & ~n6034;
  assign n6036 = ~n5604 & n32964;
  assign n6037 = ~n5602 & n6036;
  assign n6038 = n32964 & n6034;
  assign n6039 = ~n5708 & n6037;
  assign n6040 = ~n6035 & ~n33020;
  assign n6041 = n330 & ~n6014;
  assign n6042 = n330 & n6031;
  assign n6043 = ~n6030 & n6041;
  assign n6044 = ~n6040 & ~n33021;
  assign n6045 = ~n6032 & ~n6044;
  assign n6046 = ~n271 & ~n6045;
  assign n6047 = n271 & ~n6032;
  assign n6048 = ~n6044 & n6047;
  assign n6049 = ~n5619 & ~n32966;
  assign n6050 = ~n5619 & ~n5708;
  assign n6051 = ~n32966 & n6050;
  assign n6052 = ~n5708 & n6049;
  assign n6053 = n5627 & ~n33022;
  assign n6054 = n5631 & n6050;
  assign n6055 = ~n5619 & n5627;
  assign n6056 = ~n32966 & n6055;
  assign n6057 = ~n5708 & n6056;
  assign n6058 = ~n5627 & ~n33022;
  assign n6059 = ~n6057 & ~n6058;
  assign n6060 = ~n6053 & ~n6054;
  assign n6061 = ~n6048 & ~n33023;
  assign n6062 = ~n6046 & ~n6061;
  assign n6063 = ~n217 & ~n6062;
  assign n6064 = ~n5633 & ~n5635;
  assign n6065 = ~n5708 & n6064;
  assign n6066 = ~n32968 & ~n6065;
  assign n6067 = ~n5635 & n32968;
  assign n6068 = ~n5633 & n6067;
  assign n6069 = n32968 & n6065;
  assign n6070 = ~n5708 & n6068;
  assign n6071 = ~n6066 & ~n33024;
  assign n6072 = n217 & ~n6046;
  assign n6073 = n217 & n6062;
  assign n6074 = ~n6061 & n6072;
  assign n6075 = ~n6071 & ~n33025;
  assign n6076 = ~n6063 & ~n6075;
  assign n6077 = ~n198 & ~n6076;
  assign n6078 = n198 & ~n6063;
  assign n6079 = ~n6075 & n6078;
  assign n6080 = ~n5650 & ~n32970;
  assign n6081 = ~n5650 & ~n5708;
  assign n6082 = ~n32970 & n6081;
  assign n6083 = ~n5708 & n6080;
  assign n6084 = n5658 & ~n33026;
  assign n6085 = n5662 & n6081;
  assign n6086 = ~n5650 & n5658;
  assign n6087 = ~n32970 & n6086;
  assign n6088 = ~n5708 & n6087;
  assign n6089 = ~n5658 & ~n33026;
  assign n6090 = ~n6088 & ~n6089;
  assign n6091 = ~n6084 & ~n6085;
  assign n6092 = ~n6079 & ~n33027;
  assign n6093 = ~n6077 & ~n6092;
  assign n6094 = ~n5664 & ~n5666;
  assign n6095 = ~n5708 & n6094;
  assign n6096 = ~n32972 & ~n6095;
  assign n6097 = ~n5666 & n32972;
  assign n6098 = ~n5664 & n6097;
  assign n6099 = n32972 & n6095;
  assign n6100 = ~n5708 & n6098;
  assign n6101 = ~n6096 & ~n33028;
  assign n6102 = ~n5680 & ~n32974;
  assign n6103 = ~n32974 & ~n5708;
  assign n6104 = ~n5680 & n6103;
  assign n6105 = ~n5708 & n6102;
  assign n6106 = ~n32976 & ~n33029;
  assign n6107 = ~n6101 & n6106;
  assign n6108 = ~n6093 & n6107;
  assign n6109 = n193 & ~n6108;
  assign n6110 = ~n6077 & n6101;
  assign n6111 = n6093 & n6101;
  assign n6112 = ~n6092 & n6110;
  assign n6113 = n5680 & ~n6103;
  assign n6114 = ~n193 & ~n6102;
  assign n6115 = ~n6113 & n6114;
  assign n6116 = ~n33030 & ~n6115;
  assign n6117 = ~n6109 & n6116;
  assign n6118 = pi72  & ~n6117;
  assign n6119 = ~pi70  & ~pi71 ;
  assign n6120 = ~pi72  & n6119;
  assign n6121 = ~n6118 & ~n6120;
  assign n6122 = ~n5708 & ~n6121;
  assign n6123 = ~pi72  & ~n6117;
  assign n6124 = pi73  & ~n6123;
  assign n6125 = ~pi73  & n6123;
  assign n6126 = n5710 & ~n6117;
  assign n6127 = ~n6124 & ~n33031;
  assign n6128 = ~n32914 & ~n32977;
  assign n6129 = ~n5257 & n6128;
  assign n6130 = ~n5276 & n6129;
  assign n6131 = ~n32916 & n6130;
  assign n6132 = n5262 & n5278;
  assign n6133 = ~n5270 & n6131;
  assign n6134 = ~n6120 & ~n33032;
  assign n6135 = ~n5706 & n6134;
  assign n6136 = ~n32976 & n6135;
  assign n6137 = ~n5700 & n6136;
  assign n6138 = n5708 & n6121;
  assign n6139 = ~n6118 & n6137;
  assign n6140 = n6127 & ~n33033;
  assign n6141 = ~n6122 & ~n6140;
  assign n6142 = ~n5278 & ~n6141;
  assign n6143 = n5278 & ~n6122;
  assign n6144 = ~n6140 & n6143;
  assign n6145 = ~n5708 & ~n6115;
  assign n6146 = ~n33030 & n6145;
  assign n6147 = ~n6109 & n6146;
  assign n6148 = ~n33031 & ~n6147;
  assign n6149 = pi74  & ~n6148;
  assign n6150 = ~pi74  & ~n6147;
  assign n6151 = ~pi74  & n6148;
  assign n6152 = ~n33031 & n6150;
  assign n6153 = ~n6149 & ~n33034;
  assign n6154 = ~n6144 & ~n6153;
  assign n6155 = ~n6142 & ~n6154;
  assign n6156 = ~n4903 & ~n6155;
  assign n6157 = n4903 & ~n6142;
  assign n6158 = ~n6154 & n6157;
  assign n6159 = n4903 & n6155;
  assign n6160 = ~n5713 & ~n32978;
  assign n6161 = ~n6117 & n6160;
  assign n6162 = n5730 & ~n6161;
  assign n6163 = ~n5730 & n6160;
  assign n6164 = ~n5730 & n6161;
  assign n6165 = ~n6117 & n6163;
  assign n6166 = ~n6162 & ~n33036;
  assign n6167 = ~n33035 & ~n6166;
  assign n6168 = ~n6156 & ~n6167;
  assign n6169 = ~n4508 & ~n6168;
  assign n6170 = n4508 & ~n6156;
  assign n6171 = ~n6167 & n6170;
  assign n6172 = ~n5733 & ~n32981;
  assign n6173 = ~n5733 & ~n6117;
  assign n6174 = ~n32981 & n6173;
  assign n6175 = ~n6117 & n6172;
  assign n6176 = n5742 & ~n33037;
  assign n6177 = n5746 & n6173;
  assign n6178 = n5742 & ~n32981;
  assign n6179 = ~n5733 & n6178;
  assign n6180 = ~n6117 & n6179;
  assign n6181 = ~n5742 & ~n33037;
  assign n6182 = ~n6180 & ~n6181;
  assign n6183 = ~n6176 & ~n6177;
  assign n6184 = ~n6171 & ~n33038;
  assign n6185 = ~n6169 & ~n6184;
  assign n6186 = ~n4155 & ~n6185;
  assign n6187 = n4155 & ~n6169;
  assign n6188 = ~n6184 & n6187;
  assign n6189 = n4155 & n6185;
  assign n6190 = ~n5748 & ~n5750;
  assign n6191 = ~n6117 & n6190;
  assign n6192 = n5757 & ~n6191;
  assign n6193 = ~n5757 & n6191;
  assign n6194 = ~n5748 & n5757;
  assign n6195 = ~n5750 & n6194;
  assign n6196 = n5757 & n6191;
  assign n6197 = ~n6117 & n6195;
  assign n6198 = ~n5757 & ~n6191;
  assign n6199 = ~n33040 & ~n6198;
  assign n6200 = ~n6192 & ~n6193;
  assign n6201 = ~n33039 & ~n33041;
  assign n6202 = ~n6186 & ~n6201;
  assign n6203 = ~n3788 & ~n6202;
  assign n6204 = n3788 & ~n6186;
  assign n6205 = ~n6201 & n6204;
  assign n6206 = ~n5760 & ~n32984;
  assign n6207 = ~n5760 & ~n6117;
  assign n6208 = ~n32984 & n6207;
  assign n6209 = ~n6117 & n6206;
  assign n6210 = n5768 & ~n33042;
  assign n6211 = n5772 & n6207;
  assign n6212 = n5768 & ~n32984;
  assign n6213 = ~n5760 & n6212;
  assign n6214 = ~n6117 & n6213;
  assign n6215 = ~n5768 & ~n33042;
  assign n6216 = ~n6214 & ~n6215;
  assign n6217 = ~n6210 & ~n6211;
  assign n6218 = ~n6205 & ~n33043;
  assign n6219 = ~n6203 & ~n6218;
  assign n6220 = ~n3473 & ~n6219;
  assign n6221 = n3473 & ~n6203;
  assign n6222 = ~n6218 & n6221;
  assign n6223 = n3473 & n6219;
  assign n6224 = ~n5774 & ~n5776;
  assign n6225 = ~n6117 & n6224;
  assign n6226 = ~n32986 & n6225;
  assign n6227 = n32986 & ~n6225;
  assign n6228 = ~n5774 & n32986;
  assign n6229 = ~n5776 & n6228;
  assign n6230 = ~n6117 & n6229;
  assign n6231 = ~n32986 & ~n6225;
  assign n6232 = ~n6230 & ~n6231;
  assign n6233 = ~n6226 & ~n6227;
  assign n6234 = ~n33044 & ~n33045;
  assign n6235 = ~n6220 & ~n6234;
  assign n6236 = ~n3140 & ~n6235;
  assign n6237 = n3140 & ~n6220;
  assign n6238 = ~n6234 & n6237;
  assign n6239 = ~n5790 & ~n32988;
  assign n6240 = ~n5790 & ~n6117;
  assign n6241 = ~n32988 & n6240;
  assign n6242 = ~n6117 & n6239;
  assign n6243 = n5798 & ~n33046;
  assign n6244 = n5802 & n6240;
  assign n6245 = n5798 & ~n32988;
  assign n6246 = ~n5790 & n6245;
  assign n6247 = ~n6117 & n6246;
  assign n6248 = ~n5798 & ~n33046;
  assign n6249 = ~n6247 & ~n6248;
  assign n6250 = ~n6243 & ~n6244;
  assign n6251 = ~n6238 & ~n33047;
  assign n6252 = ~n6236 & ~n6251;
  assign n6253 = ~n2855 & ~n6252;
  assign n6254 = n2855 & ~n6236;
  assign n6255 = ~n6251 & n6254;
  assign n6256 = n2855 & n6252;
  assign n6257 = ~n5804 & ~n5806;
  assign n6258 = ~n6117 & n6257;
  assign n6259 = ~n32989 & ~n6258;
  assign n6260 = ~n5804 & n32989;
  assign n6261 = ~n5806 & n6260;
  assign n6262 = n32989 & n6258;
  assign n6263 = ~n6117 & n6261;
  assign n6264 = n32989 & ~n6258;
  assign n6265 = ~n32989 & n6258;
  assign n6266 = ~n6264 & ~n6265;
  assign n6267 = ~n6259 & ~n33049;
  assign n6268 = ~n33048 & n33050;
  assign n6269 = ~n6253 & ~n6268;
  assign n6270 = ~n2556 & ~n6269;
  assign n6271 = n2556 & ~n6253;
  assign n6272 = ~n6268 & n6271;
  assign n6273 = ~n5819 & ~n32991;
  assign n6274 = ~n5819 & ~n6117;
  assign n6275 = ~n32991 & n6274;
  assign n6276 = ~n6117 & n6273;
  assign n6277 = n5827 & ~n33051;
  assign n6278 = n5831 & n6274;
  assign n6279 = n5827 & ~n32991;
  assign n6280 = ~n5819 & n6279;
  assign n6281 = ~n6117 & n6280;
  assign n6282 = ~n5827 & ~n33051;
  assign n6283 = ~n6281 & ~n6282;
  assign n6284 = ~n6277 & ~n6278;
  assign n6285 = ~n6272 & ~n33052;
  assign n6286 = ~n6270 & ~n6285;
  assign n6287 = ~n2301 & ~n6286;
  assign n6288 = n2301 & ~n6270;
  assign n6289 = ~n6285 & n6288;
  assign n6290 = n2301 & n6286;
  assign n6291 = ~n5833 & ~n5835;
  assign n6292 = ~n6117 & n6291;
  assign n6293 = n32993 & ~n6292;
  assign n6294 = ~n5833 & ~n32993;
  assign n6295 = ~n5835 & n6294;
  assign n6296 = ~n32993 & n6292;
  assign n6297 = ~n6117 & n6295;
  assign n6298 = n32993 & n6292;
  assign n6299 = ~n32993 & ~n6292;
  assign n6300 = ~n6298 & ~n6299;
  assign n6301 = ~n6293 & ~n33054;
  assign n6302 = ~n33053 & n33055;
  assign n6303 = ~n6287 & ~n6302;
  assign n6304 = ~n2038 & ~n6303;
  assign n6305 = n2038 & ~n6287;
  assign n6306 = ~n6302 & n6305;
  assign n6307 = ~n5849 & ~n32995;
  assign n6308 = ~n5849 & ~n6117;
  assign n6309 = ~n32995 & n6308;
  assign n6310 = ~n6117 & n6307;
  assign n6311 = n5857 & ~n33056;
  assign n6312 = n5861 & n6308;
  assign n6313 = n5857 & ~n32995;
  assign n6314 = ~n5849 & n6313;
  assign n6315 = ~n6117 & n6314;
  assign n6316 = ~n5857 & ~n33056;
  assign n6317 = ~n6315 & ~n6316;
  assign n6318 = ~n6311 & ~n6312;
  assign n6319 = ~n6306 & ~n33057;
  assign n6320 = ~n6304 & ~n6319;
  assign n6321 = ~n1812 & ~n6320;
  assign n6322 = n1812 & ~n6304;
  assign n6323 = ~n6319 & n6322;
  assign n6324 = n1812 & n6320;
  assign n6325 = ~n5863 & ~n5865;
  assign n6326 = ~n5863 & ~n6117;
  assign n6327 = ~n5865 & n6326;
  assign n6328 = ~n6117 & n6325;
  assign n6329 = ~n32997 & ~n33059;
  assign n6330 = n5877 & n6326;
  assign n6331 = n32997 & n33059;
  assign n6332 = ~n5863 & ~n32997;
  assign n6333 = ~n5865 & n6332;
  assign n6334 = ~n6117 & n6333;
  assign n6335 = n32997 & ~n33059;
  assign n6336 = ~n6334 & ~n6335;
  assign n6337 = ~n6329 & ~n33060;
  assign n6338 = ~n33058 & ~n33061;
  assign n6339 = ~n6321 & ~n6338;
  assign n6340 = ~n1582 & ~n6339;
  assign n6341 = n1582 & ~n6321;
  assign n6342 = ~n6338 & n6341;
  assign n6343 = ~n5879 & ~n32999;
  assign n6344 = ~n5879 & ~n6117;
  assign n6345 = ~n32999 & n6344;
  assign n6346 = ~n6117 & n6343;
  assign n6347 = n5887 & ~n33062;
  assign n6348 = n5891 & n6344;
  assign n6349 = n5887 & ~n32999;
  assign n6350 = ~n5879 & n6349;
  assign n6351 = ~n6117 & n6350;
  assign n6352 = ~n5887 & ~n33062;
  assign n6353 = ~n6351 & ~n6352;
  assign n6354 = ~n6347 & ~n6348;
  assign n6355 = ~n6342 & ~n33063;
  assign n6356 = ~n6340 & ~n6355;
  assign n6357 = ~n1388 & ~n6356;
  assign n6358 = n1388 & ~n6340;
  assign n6359 = ~n6355 & n6358;
  assign n6360 = n1388 & n6356;
  assign n6361 = ~n5893 & ~n5895;
  assign n6362 = ~n6117 & n6361;
  assign n6363 = ~n33002 & ~n6362;
  assign n6364 = ~n5893 & n33002;
  assign n6365 = ~n5895 & n6364;
  assign n6366 = n33002 & n6362;
  assign n6367 = ~n6117 & n6365;
  assign n6368 = ~n6363 & ~n33065;
  assign n6369 = ~n33064 & ~n6368;
  assign n6370 = ~n6357 & ~n6369;
  assign n6371 = ~n1192 & ~n6370;
  assign n6372 = n1192 & ~n6357;
  assign n6373 = ~n6369 & n6372;
  assign n6374 = ~n5911 & ~n33004;
  assign n6375 = ~n5911 & ~n6117;
  assign n6376 = ~n33004 & n6375;
  assign n6377 = ~n6117 & n6374;
  assign n6378 = n5919 & ~n33066;
  assign n6379 = n5923 & n6375;
  assign n6380 = n5919 & ~n33004;
  assign n6381 = ~n5911 & n6380;
  assign n6382 = ~n6117 & n6381;
  assign n6383 = ~n5919 & ~n33066;
  assign n6384 = ~n6382 & ~n6383;
  assign n6385 = ~n6378 & ~n6379;
  assign n6386 = ~n6373 & ~n33067;
  assign n6387 = ~n6371 & ~n6386;
  assign n6388 = ~n1028 & ~n6387;
  assign n6389 = n1028 & ~n6371;
  assign n6390 = ~n6386 & n6389;
  assign n6391 = n1028 & n6387;
  assign n6392 = ~n5925 & ~n5927;
  assign n6393 = ~n5925 & ~n6117;
  assign n6394 = ~n5927 & n6393;
  assign n6395 = ~n6117 & n6392;
  assign n6396 = n5935 & ~n33069;
  assign n6397 = n5936 & n6393;
  assign n6398 = ~n5935 & n33069;
  assign n6399 = ~n5925 & n5935;
  assign n6400 = ~n5927 & n6399;
  assign n6401 = ~n6117 & n6400;
  assign n6402 = ~n5935 & ~n33069;
  assign n6403 = ~n6401 & ~n6402;
  assign n6404 = ~n6396 & ~n33070;
  assign n6405 = ~n33068 & ~n33071;
  assign n6406 = ~n6388 & ~n6405;
  assign n6407 = ~n866 & ~n6406;
  assign n6408 = n866 & ~n6388;
  assign n6409 = ~n6405 & n6408;
  assign n6410 = ~n5938 & ~n33007;
  assign n6411 = ~n5938 & ~n6117;
  assign n6412 = ~n33007 & n6411;
  assign n6413 = ~n6117 & n6410;
  assign n6414 = n5946 & ~n33072;
  assign n6415 = n5950 & n6411;
  assign n6416 = n5946 & ~n33007;
  assign n6417 = ~n5938 & n6416;
  assign n6418 = ~n6117 & n6417;
  assign n6419 = ~n5946 & ~n33072;
  assign n6420 = ~n6418 & ~n6419;
  assign n6421 = ~n6414 & ~n6415;
  assign n6422 = ~n6409 & ~n33073;
  assign n6423 = ~n6407 & ~n6422;
  assign n6424 = ~n730 & ~n6423;
  assign n6425 = n730 & ~n6407;
  assign n6426 = ~n6422 & n6425;
  assign n6427 = n730 & n6423;
  assign n6428 = ~n5952 & ~n5954;
  assign n6429 = ~n6117 & n6428;
  assign n6430 = ~n33010 & n6429;
  assign n6431 = n33010 & ~n6429;
  assign n6432 = ~n5952 & n33010;
  assign n6433 = ~n5954 & n6432;
  assign n6434 = n33010 & n6429;
  assign n6435 = ~n6117 & n6433;
  assign n6436 = ~n33010 & ~n6429;
  assign n6437 = ~n33075 & ~n6436;
  assign n6438 = ~n6430 & ~n6431;
  assign n6439 = ~n33074 & ~n33076;
  assign n6440 = ~n6424 & ~n6439;
  assign n6441 = ~n602 & ~n6440;
  assign n6442 = n602 & ~n6424;
  assign n6443 = ~n6439 & n6442;
  assign n6444 = ~n5970 & ~n33012;
  assign n6445 = ~n5970 & ~n6117;
  assign n6446 = ~n33012 & n6445;
  assign n6447 = ~n6117 & n6444;
  assign n6448 = n5978 & ~n33077;
  assign n6449 = n5982 & n6445;
  assign n6450 = n5978 & ~n33012;
  assign n6451 = ~n5970 & n6450;
  assign n6452 = ~n6117 & n6451;
  assign n6453 = ~n5978 & ~n33077;
  assign n6454 = ~n6452 & ~n6453;
  assign n6455 = ~n6448 & ~n6449;
  assign n6456 = ~n6443 & ~n33078;
  assign n6457 = ~n6441 & ~n6456;
  assign n6458 = ~n497 & ~n6457;
  assign n6459 = n497 & ~n6441;
  assign n6460 = ~n6456 & n6459;
  assign n6461 = n497 & n6457;
  assign n6462 = ~n5984 & ~n5986;
  assign n6463 = ~n5984 & ~n6117;
  assign n6464 = ~n5986 & n6463;
  assign n6465 = ~n6117 & n6462;
  assign n6466 = n33014 & ~n33080;
  assign n6467 = n5998 & n6463;
  assign n6468 = ~n33014 & n33080;
  assign n6469 = ~n5984 & n33014;
  assign n6470 = ~n5986 & n6469;
  assign n6471 = ~n6117 & n6470;
  assign n6472 = ~n33014 & ~n33080;
  assign n6473 = ~n6471 & ~n6472;
  assign n6474 = ~n6466 & ~n33081;
  assign n6475 = ~n33079 & ~n33082;
  assign n6476 = ~n6458 & ~n6475;
  assign n6477 = ~n403 & ~n6476;
  assign n6478 = n403 & ~n6458;
  assign n6479 = ~n6475 & n6478;
  assign n6480 = ~n6000 & ~n33016;
  assign n6481 = ~n6000 & ~n6117;
  assign n6482 = ~n33016 & n6481;
  assign n6483 = ~n6117 & n6480;
  assign n6484 = n6008 & ~n33083;
  assign n6485 = n6012 & n6481;
  assign n6486 = n6008 & ~n33016;
  assign n6487 = ~n6000 & n6486;
  assign n6488 = ~n6117 & n6487;
  assign n6489 = ~n6008 & ~n33083;
  assign n6490 = ~n6488 & ~n6489;
  assign n6491 = ~n6484 & ~n6485;
  assign n6492 = ~n6479 & ~n33084;
  assign n6493 = ~n6477 & ~n6492;
  assign n6494 = ~n330 & ~n6493;
  assign n6495 = ~n6014 & ~n6016;
  assign n6496 = ~n6117 & n6495;
  assign n6497 = ~n33019 & ~n6496;
  assign n6498 = ~n6014 & n33019;
  assign n6499 = ~n6016 & n6498;
  assign n6500 = n33019 & n6496;
  assign n6501 = ~n6117 & n6499;
  assign n6502 = ~n6497 & ~n33085;
  assign n6503 = n330 & ~n6477;
  assign n6504 = ~n6492 & n6503;
  assign n6505 = n330 & n6493;
  assign n6506 = ~n6502 & ~n33086;
  assign n6507 = ~n6494 & ~n6506;
  assign n6508 = ~n271 & ~n6507;
  assign n6509 = n271 & ~n6494;
  assign n6510 = ~n6506 & n6509;
  assign n6511 = ~n6032 & ~n33021;
  assign n6512 = ~n6032 & ~n6117;
  assign n6513 = ~n33021 & n6512;
  assign n6514 = ~n6117 & n6511;
  assign n6515 = n6040 & ~n33087;
  assign n6516 = n6044 & n6512;
  assign n6517 = n6040 & ~n33021;
  assign n6518 = ~n6032 & n6517;
  assign n6519 = ~n6117 & n6518;
  assign n6520 = ~n6040 & ~n33087;
  assign n6521 = ~n6519 & ~n6520;
  assign n6522 = ~n6515 & ~n6516;
  assign n6523 = ~n6510 & ~n33088;
  assign n6524 = ~n6508 & ~n6523;
  assign n6525 = ~n217 & ~n6524;
  assign n6526 = ~n6046 & ~n6048;
  assign n6527 = ~n6117 & n6526;
  assign n6528 = ~n33023 & ~n6527;
  assign n6529 = ~n6046 & n33023;
  assign n6530 = ~n6048 & n6529;
  assign n6531 = n33023 & n6527;
  assign n6532 = ~n6117 & n6530;
  assign n6533 = ~n6528 & ~n33089;
  assign n6534 = n217 & ~n6508;
  assign n6535 = ~n6523 & n6534;
  assign n6536 = n217 & n6524;
  assign n6537 = ~n6533 & ~n33090;
  assign n6538 = ~n6525 & ~n6537;
  assign n6539 = ~n198 & ~n6538;
  assign n6540 = n198 & ~n6525;
  assign n6541 = ~n6537 & n6540;
  assign n6542 = ~n6063 & ~n33025;
  assign n6543 = ~n6063 & ~n6117;
  assign n6544 = ~n33025 & n6543;
  assign n6545 = ~n6117 & n6542;
  assign n6546 = n6071 & ~n33091;
  assign n6547 = n6075 & n6543;
  assign n6548 = n6071 & ~n33025;
  assign n6549 = ~n6063 & n6548;
  assign n6550 = ~n6117 & n6549;
  assign n6551 = ~n6071 & ~n33091;
  assign n6552 = ~n6550 & ~n6551;
  assign n6553 = ~n6546 & ~n6547;
  assign n6554 = ~n6541 & ~n33092;
  assign n6555 = ~n6539 & ~n6554;
  assign n6556 = ~n6077 & ~n6079;
  assign n6557 = ~n6117 & n6556;
  assign n6558 = ~n33027 & ~n6557;
  assign n6559 = ~n6077 & n33027;
  assign n6560 = ~n6079 & n6559;
  assign n6561 = n33027 & n6557;
  assign n6562 = ~n6117 & n6560;
  assign n6563 = ~n6558 & ~n33093;
  assign n6564 = ~n6093 & ~n6101;
  assign n6565 = ~n6101 & ~n6117;
  assign n6566 = ~n6093 & n6565;
  assign n6567 = ~n6117 & n6564;
  assign n6568 = ~n33030 & ~n33094;
  assign n6569 = ~n6563 & n6568;
  assign n6570 = ~n6555 & n6569;
  assign n6571 = n193 & ~n6570;
  assign n6572 = ~n6539 & n6563;
  assign n6573 = ~n6554 & n6572;
  assign n6574 = n6555 & n6563;
  assign n6575 = n6093 & ~n6565;
  assign n6576 = ~n193 & ~n6564;
  assign n6577 = ~n6575 & n6576;
  assign n6578 = ~n33095 & ~n6577;
  assign n6579 = ~n6571 & n6578;
  assign n6580 = pi70  & ~n6579;
  assign n6581 = ~pi68  & ~pi69 ;
  assign n6582 = ~pi70  & n6581;
  assign n6583 = ~n6580 & ~n6582;
  assign n6584 = ~n6117 & ~n6583;
  assign n6585 = ~n5689 & ~n33032;
  assign n6586 = ~n5690 & n6585;
  assign n6587 = ~n5706 & n6586;
  assign n6588 = ~n32976 & n6587;
  assign n6589 = n32974 & n5708;
  assign n6590 = ~n5700 & n6588;
  assign n6591 = ~n6582 & ~n33096;
  assign n6592 = ~n6115 & n6591;
  assign n6593 = ~n33030 & n6592;
  assign n6594 = ~n6109 & n6593;
  assign n6595 = n6117 & n6583;
  assign n6596 = ~n6580 & n6594;
  assign n6597 = ~pi70  & ~n6579;
  assign n6598 = pi71  & ~n6597;
  assign n6599 = ~pi71  & n6597;
  assign n6600 = n6119 & ~n6579;
  assign n6601 = ~n6598 & ~n33098;
  assign n6602 = ~n33097 & n6601;
  assign n6603 = ~n6584 & ~n6602;
  assign n6604 = ~n5708 & ~n6603;
  assign n6605 = ~n6117 & ~n6577;
  assign n6606 = ~n33095 & n6605;
  assign n6607 = ~n6571 & n6606;
  assign n6608 = ~n33098 & ~n6607;
  assign n6609 = pi72  & ~n6608;
  assign n6610 = ~pi72  & ~n6607;
  assign n6611 = ~pi72  & n6608;
  assign n6612 = ~n33098 & n6610;
  assign n6613 = ~n6609 & ~n33099;
  assign n6614 = n5708 & ~n6584;
  assign n6615 = n5708 & n6603;
  assign n6616 = ~n6602 & n6614;
  assign n6617 = ~n6613 & ~n33100;
  assign n6618 = ~n6604 & ~n6617;
  assign n6619 = ~n5278 & ~n6618;
  assign n6620 = n5278 & ~n6604;
  assign n6621 = ~n6617 & n6620;
  assign n6622 = ~n6122 & ~n33033;
  assign n6623 = ~n6579 & n6622;
  assign n6624 = n6127 & ~n6623;
  assign n6625 = ~n6127 & n6622;
  assign n6626 = ~n6127 & n6623;
  assign n6627 = ~n6579 & n6625;
  assign n6628 = ~n6624 & ~n33101;
  assign n6629 = ~n6621 & ~n6628;
  assign n6630 = ~n6619 & ~n6629;
  assign n6631 = ~n4903 & ~n6630;
  assign n6632 = ~n6142 & ~n6144;
  assign n6633 = ~n6579 & n6632;
  assign n6634 = ~n6153 & ~n6633;
  assign n6635 = ~n6144 & n6153;
  assign n6636 = ~n6142 & n6635;
  assign n6637 = n6153 & n6633;
  assign n6638 = ~n6579 & n6636;
  assign n6639 = ~n6634 & ~n33102;
  assign n6640 = n4903 & ~n6619;
  assign n6641 = n4903 & n6630;
  assign n6642 = ~n6629 & n6640;
  assign n6643 = ~n6639 & ~n33103;
  assign n6644 = ~n6631 & ~n6643;
  assign n6645 = ~n4508 & ~n6644;
  assign n6646 = n4508 & ~n6631;
  assign n6647 = ~n6643 & n6646;
  assign n6648 = ~n6156 & ~n33035;
  assign n6649 = ~n6579 & n6648;
  assign n6650 = n6166 & ~n6649;
  assign n6651 = ~n6166 & n6649;
  assign n6652 = ~n6156 & n6166;
  assign n6653 = ~n33035 & n6652;
  assign n6654 = n6166 & n6649;
  assign n6655 = ~n6579 & n6653;
  assign n6656 = ~n6166 & ~n6649;
  assign n6657 = ~n33104 & ~n6656;
  assign n6658 = ~n6650 & ~n6651;
  assign n6659 = ~n6647 & ~n33105;
  assign n6660 = ~n6645 & ~n6659;
  assign n6661 = ~n4155 & ~n6660;
  assign n6662 = ~n6169 & ~n6171;
  assign n6663 = ~n6579 & n6662;
  assign n6664 = ~n33038 & ~n6663;
  assign n6665 = ~n6171 & n33038;
  assign n6666 = ~n6169 & n6665;
  assign n6667 = n33038 & n6663;
  assign n6668 = ~n6579 & n6666;
  assign n6669 = ~n6664 & ~n33106;
  assign n6670 = n4155 & ~n6645;
  assign n6671 = n4155 & n6660;
  assign n6672 = ~n6659 & n6670;
  assign n6673 = ~n6669 & ~n33107;
  assign n6674 = ~n6661 & ~n6673;
  assign n6675 = ~n3788 & ~n6674;
  assign n6676 = n3788 & ~n6661;
  assign n6677 = ~n6673 & n6676;
  assign n6678 = ~n6186 & ~n33039;
  assign n6679 = ~n6579 & n6678;
  assign n6680 = ~n33041 & n6679;
  assign n6681 = n33041 & ~n6679;
  assign n6682 = ~n6186 & n33041;
  assign n6683 = ~n33039 & n6682;
  assign n6684 = ~n6579 & n6683;
  assign n6685 = ~n33041 & ~n6679;
  assign n6686 = ~n6684 & ~n6685;
  assign n6687 = ~n6680 & ~n6681;
  assign n6688 = ~n6677 & ~n33108;
  assign n6689 = ~n6675 & ~n6688;
  assign n6690 = ~n3473 & ~n6689;
  assign n6691 = ~n6203 & ~n6205;
  assign n6692 = ~n6579 & n6691;
  assign n6693 = ~n33043 & ~n6692;
  assign n6694 = ~n6205 & n33043;
  assign n6695 = ~n6203 & n6694;
  assign n6696 = n33043 & n6692;
  assign n6697 = ~n6579 & n6695;
  assign n6698 = ~n6693 & ~n33109;
  assign n6699 = n3473 & ~n6675;
  assign n6700 = n3473 & n6689;
  assign n6701 = ~n6688 & n6699;
  assign n6702 = ~n6698 & ~n33110;
  assign n6703 = ~n6690 & ~n6702;
  assign n6704 = ~n3140 & ~n6703;
  assign n6705 = n3140 & ~n6690;
  assign n6706 = ~n6702 & n6705;
  assign n6707 = ~n6220 & ~n33044;
  assign n6708 = ~n6579 & n6707;
  assign n6709 = ~n33045 & ~n6708;
  assign n6710 = ~n6220 & n33045;
  assign n6711 = ~n33044 & n6710;
  assign n6712 = n33045 & n6708;
  assign n6713 = ~n6579 & n6711;
  assign n6714 = n33045 & ~n6708;
  assign n6715 = ~n33045 & n6708;
  assign n6716 = ~n6714 & ~n6715;
  assign n6717 = ~n6709 & ~n33111;
  assign n6718 = ~n6706 & n33112;
  assign n6719 = ~n6704 & ~n6718;
  assign n6720 = ~n2855 & ~n6719;
  assign n6721 = ~n6236 & ~n6238;
  assign n6722 = ~n6579 & n6721;
  assign n6723 = ~n33047 & ~n6722;
  assign n6724 = ~n6238 & n33047;
  assign n6725 = ~n6236 & n6724;
  assign n6726 = n33047 & n6722;
  assign n6727 = ~n6579 & n6725;
  assign n6728 = ~n6723 & ~n33113;
  assign n6729 = n2855 & ~n6704;
  assign n6730 = n2855 & n6719;
  assign n6731 = ~n6718 & n6729;
  assign n6732 = ~n6728 & ~n33114;
  assign n6733 = ~n6720 & ~n6732;
  assign n6734 = ~n2556 & ~n6733;
  assign n6735 = n2556 & ~n6720;
  assign n6736 = ~n6732 & n6735;
  assign n6737 = ~n6253 & ~n33048;
  assign n6738 = ~n6579 & n6737;
  assign n6739 = n33050 & ~n6738;
  assign n6740 = ~n6253 & ~n33050;
  assign n6741 = ~n33048 & n6740;
  assign n6742 = ~n33050 & n6738;
  assign n6743 = ~n6579 & n6741;
  assign n6744 = n33050 & n6738;
  assign n6745 = ~n33050 & ~n6738;
  assign n6746 = ~n6744 & ~n6745;
  assign n6747 = ~n6739 & ~n33115;
  assign n6748 = ~n6736 & n33116;
  assign n6749 = ~n6734 & ~n6748;
  assign n6750 = ~n2301 & ~n6749;
  assign n6751 = ~n6270 & ~n6272;
  assign n6752 = ~n6579 & n6751;
  assign n6753 = ~n33052 & ~n6752;
  assign n6754 = ~n6272 & n33052;
  assign n6755 = ~n6270 & n6754;
  assign n6756 = n33052 & n6752;
  assign n6757 = ~n6579 & n6755;
  assign n6758 = ~n6753 & ~n33117;
  assign n6759 = n2301 & ~n6734;
  assign n6760 = n2301 & n6749;
  assign n6761 = ~n6748 & n6759;
  assign n6762 = ~n6758 & ~n33118;
  assign n6763 = ~n6750 & ~n6762;
  assign n6764 = ~n2038 & ~n6763;
  assign n6765 = n2038 & ~n6750;
  assign n6766 = ~n6762 & n6765;
  assign n6767 = ~n6287 & ~n33053;
  assign n6768 = ~n6287 & ~n6579;
  assign n6769 = ~n33053 & n6768;
  assign n6770 = ~n6579 & n6767;
  assign n6771 = ~n33055 & ~n33119;
  assign n6772 = n6302 & n6768;
  assign n6773 = n33055 & n33119;
  assign n6774 = ~n6287 & ~n33055;
  assign n6775 = ~n33053 & n6774;
  assign n6776 = ~n6579 & n6775;
  assign n6777 = n33055 & ~n33119;
  assign n6778 = ~n6776 & ~n6777;
  assign n6779 = ~n6771 & ~n33120;
  assign n6780 = ~n6766 & ~n33121;
  assign n6781 = ~n6764 & ~n6780;
  assign n6782 = ~n1812 & ~n6781;
  assign n6783 = ~n6304 & ~n6306;
  assign n6784 = ~n6579 & n6783;
  assign n6785 = ~n33057 & ~n6784;
  assign n6786 = ~n6306 & n33057;
  assign n6787 = ~n6304 & n6786;
  assign n6788 = n33057 & n6784;
  assign n6789 = ~n6579 & n6787;
  assign n6790 = ~n6785 & ~n33122;
  assign n6791 = n1812 & ~n6764;
  assign n6792 = n1812 & n6781;
  assign n6793 = ~n6780 & n6791;
  assign n6794 = ~n6790 & ~n33123;
  assign n6795 = ~n6782 & ~n6794;
  assign n6796 = ~n1582 & ~n6795;
  assign n6797 = n1582 & ~n6782;
  assign n6798 = ~n6794 & n6797;
  assign n6799 = ~n6321 & ~n33058;
  assign n6800 = ~n6579 & n6799;
  assign n6801 = ~n33061 & ~n6800;
  assign n6802 = ~n6321 & n33061;
  assign n6803 = ~n33058 & n6802;
  assign n6804 = n33061 & n6800;
  assign n6805 = ~n6579 & n6803;
  assign n6806 = ~n6801 & ~n33124;
  assign n6807 = ~n6798 & ~n6806;
  assign n6808 = ~n6796 & ~n6807;
  assign n6809 = ~n1388 & ~n6808;
  assign n6810 = ~n6340 & ~n6342;
  assign n6811 = ~n6579 & n6810;
  assign n6812 = ~n33063 & ~n6811;
  assign n6813 = ~n6342 & n33063;
  assign n6814 = ~n6340 & n6813;
  assign n6815 = n33063 & n6811;
  assign n6816 = ~n6579 & n6814;
  assign n6817 = ~n6812 & ~n33125;
  assign n6818 = n1388 & ~n6796;
  assign n6819 = n1388 & n6808;
  assign n6820 = ~n6807 & n6818;
  assign n6821 = ~n6817 & ~n33126;
  assign n6822 = ~n6809 & ~n6821;
  assign n6823 = ~n1192 & ~n6822;
  assign n6824 = n1192 & ~n6809;
  assign n6825 = ~n6821 & n6824;
  assign n6826 = ~n6357 & ~n33064;
  assign n6827 = ~n6357 & ~n6579;
  assign n6828 = ~n33064 & n6827;
  assign n6829 = ~n6579 & n6826;
  assign n6830 = n6368 & ~n33127;
  assign n6831 = n6369 & n6827;
  assign n6832 = ~n6368 & n33127;
  assign n6833 = ~n6357 & n6368;
  assign n6834 = ~n33064 & n6833;
  assign n6835 = ~n6579 & n6834;
  assign n6836 = ~n6368 & ~n33127;
  assign n6837 = ~n6835 & ~n6836;
  assign n6838 = ~n6830 & ~n33128;
  assign n6839 = ~n6825 & ~n33129;
  assign n6840 = ~n6823 & ~n6839;
  assign n6841 = ~n1028 & ~n6840;
  assign n6842 = ~n6371 & ~n6373;
  assign n6843 = ~n6579 & n6842;
  assign n6844 = ~n33067 & ~n6843;
  assign n6845 = ~n6373 & n33067;
  assign n6846 = ~n6371 & n6845;
  assign n6847 = n33067 & n6843;
  assign n6848 = ~n6579 & n6846;
  assign n6849 = ~n6844 & ~n33130;
  assign n6850 = n1028 & ~n6823;
  assign n6851 = n1028 & n6840;
  assign n6852 = ~n6839 & n6850;
  assign n6853 = ~n6849 & ~n33131;
  assign n6854 = ~n6841 & ~n6853;
  assign n6855 = ~n866 & ~n6854;
  assign n6856 = n866 & ~n6841;
  assign n6857 = ~n6853 & n6856;
  assign n6858 = ~n6388 & ~n33068;
  assign n6859 = ~n6579 & n6858;
  assign n6860 = ~n33071 & n6859;
  assign n6861 = n33071 & ~n6859;
  assign n6862 = ~n6388 & n33071;
  assign n6863 = ~n33068 & n6862;
  assign n6864 = n33071 & n6859;
  assign n6865 = ~n6579 & n6863;
  assign n6866 = ~n33071 & ~n6859;
  assign n6867 = ~n33132 & ~n6866;
  assign n6868 = ~n6860 & ~n6861;
  assign n6869 = ~n6857 & ~n33133;
  assign n6870 = ~n6855 & ~n6869;
  assign n6871 = ~n730 & ~n6870;
  assign n6872 = ~n6407 & ~n6409;
  assign n6873 = ~n6579 & n6872;
  assign n6874 = ~n33073 & ~n6873;
  assign n6875 = ~n6409 & n33073;
  assign n6876 = ~n6407 & n6875;
  assign n6877 = n33073 & n6873;
  assign n6878 = ~n6579 & n6876;
  assign n6879 = ~n6874 & ~n33134;
  assign n6880 = n730 & ~n6855;
  assign n6881 = n730 & n6870;
  assign n6882 = ~n6869 & n6880;
  assign n6883 = ~n6879 & ~n33135;
  assign n6884 = ~n6871 & ~n6883;
  assign n6885 = ~n602 & ~n6884;
  assign n6886 = n602 & ~n6871;
  assign n6887 = ~n6883 & n6886;
  assign n6888 = ~n6424 & ~n33074;
  assign n6889 = ~n6424 & ~n6579;
  assign n6890 = ~n33074 & n6889;
  assign n6891 = ~n6579 & n6888;
  assign n6892 = n33076 & ~n33136;
  assign n6893 = n6439 & n6889;
  assign n6894 = ~n33076 & n33136;
  assign n6895 = ~n6424 & n33076;
  assign n6896 = ~n33074 & n6895;
  assign n6897 = ~n6579 & n6896;
  assign n6898 = ~n33076 & ~n33136;
  assign n6899 = ~n6897 & ~n6898;
  assign n6900 = ~n6892 & ~n33137;
  assign n6901 = ~n6887 & ~n33138;
  assign n6902 = ~n6885 & ~n6901;
  assign n6903 = ~n497 & ~n6902;
  assign n6904 = ~n6441 & ~n6443;
  assign n6905 = ~n6579 & n6904;
  assign n6906 = ~n33078 & ~n6905;
  assign n6907 = ~n6443 & n33078;
  assign n6908 = ~n6441 & n6907;
  assign n6909 = n33078 & n6905;
  assign n6910 = ~n6579 & n6908;
  assign n6911 = ~n6906 & ~n33139;
  assign n6912 = n497 & ~n6885;
  assign n6913 = n497 & n6902;
  assign n6914 = ~n6901 & n6912;
  assign n6915 = ~n6911 & ~n33140;
  assign n6916 = ~n6903 & ~n6915;
  assign n6917 = ~n403 & ~n6916;
  assign n6918 = ~n6458 & ~n33079;
  assign n6919 = ~n6579 & n6918;
  assign n6920 = ~n33082 & ~n6919;
  assign n6921 = ~n6458 & n33082;
  assign n6922 = ~n33079 & n6921;
  assign n6923 = n33082 & n6919;
  assign n6924 = ~n6579 & n6922;
  assign n6925 = ~n6920 & ~n33141;
  assign n6926 = n403 & ~n6903;
  assign n6927 = ~n6915 & n6926;
  assign n6928 = ~n6925 & ~n6927;
  assign n6929 = ~n6917 & ~n6928;
  assign n6930 = ~n330 & ~n6929;
  assign n6931 = ~n6477 & ~n6479;
  assign n6932 = ~n6579 & n6931;
  assign n6933 = ~n33084 & ~n6932;
  assign n6934 = ~n6479 & n33084;
  assign n6935 = ~n6477 & n6934;
  assign n6936 = n33084 & n6932;
  assign n6937 = ~n6579 & n6935;
  assign n6938 = ~n6933 & ~n33142;
  assign n6939 = n330 & ~n6917;
  assign n6940 = n330 & n6929;
  assign n6941 = ~n6928 & n6939;
  assign n6942 = ~n6938 & ~n33143;
  assign n6943 = ~n6930 & ~n6942;
  assign n6944 = ~n271 & ~n6943;
  assign n6945 = n271 & ~n6930;
  assign n6946 = ~n6942 & n6945;
  assign n6947 = ~n6494 & ~n33086;
  assign n6948 = ~n6494 & ~n6579;
  assign n6949 = ~n33086 & n6948;
  assign n6950 = ~n6579 & n6947;
  assign n6951 = n6502 & ~n33144;
  assign n6952 = n6506 & n6948;
  assign n6953 = ~n6494 & n6502;
  assign n6954 = ~n33086 & n6953;
  assign n6955 = ~n6579 & n6954;
  assign n6956 = ~n6502 & ~n33144;
  assign n6957 = ~n6955 & ~n6956;
  assign n6958 = ~n6951 & ~n6952;
  assign n6959 = ~n6946 & ~n33145;
  assign n6960 = ~n6944 & ~n6959;
  assign n6961 = ~n217 & ~n6960;
  assign n6962 = ~n6508 & ~n6510;
  assign n6963 = ~n6579 & n6962;
  assign n6964 = ~n33088 & ~n6963;
  assign n6965 = ~n6510 & n33088;
  assign n6966 = ~n6508 & n6965;
  assign n6967 = n33088 & n6963;
  assign n6968 = ~n6579 & n6966;
  assign n6969 = ~n6964 & ~n33146;
  assign n6970 = n217 & ~n6944;
  assign n6971 = n217 & n6960;
  assign n6972 = ~n6959 & n6970;
  assign n6973 = ~n6969 & ~n33147;
  assign n6974 = ~n6961 & ~n6973;
  assign n6975 = ~n198 & ~n6974;
  assign n6976 = n198 & ~n6961;
  assign n6977 = ~n6973 & n6976;
  assign n6978 = ~n6525 & ~n33090;
  assign n6979 = ~n6525 & ~n6579;
  assign n6980 = ~n33090 & n6979;
  assign n6981 = ~n6579 & n6978;
  assign n6982 = n6533 & ~n33148;
  assign n6983 = n6537 & n6979;
  assign n6984 = ~n6525 & n6533;
  assign n6985 = ~n33090 & n6984;
  assign n6986 = ~n6579 & n6985;
  assign n6987 = ~n6533 & ~n33148;
  assign n6988 = ~n6986 & ~n6987;
  assign n6989 = ~n6982 & ~n6983;
  assign n6990 = ~n6977 & ~n33149;
  assign n6991 = ~n6975 & ~n6990;
  assign n6992 = ~n6539 & ~n6541;
  assign n6993 = ~n6579 & n6992;
  assign n6994 = ~n33092 & ~n6993;
  assign n6995 = ~n6541 & n33092;
  assign n6996 = ~n6539 & n6995;
  assign n6997 = n33092 & n6993;
  assign n6998 = ~n6579 & n6996;
  assign n6999 = ~n6994 & ~n33150;
  assign n7000 = ~n6555 & ~n6563;
  assign n7001 = ~n6563 & ~n6579;
  assign n7002 = ~n6555 & n7001;
  assign n7003 = ~n6579 & n7000;
  assign n7004 = ~n33095 & ~n33151;
  assign n7005 = ~n6999 & n7004;
  assign n7006 = ~n6991 & n7005;
  assign n7007 = n193 & ~n7006;
  assign n7008 = ~n6975 & n6999;
  assign n7009 = n6991 & n6999;
  assign n7010 = ~n6990 & n7008;
  assign n7011 = n6555 & ~n7001;
  assign n7012 = ~n193 & ~n7000;
  assign n7013 = ~n7011 & n7012;
  assign n7014 = ~n33152 & ~n7013;
  assign n7015 = ~n7007 & n7014;
  assign n7016 = pi68  & ~n7015;
  assign n7017 = ~pi66  & ~pi67 ;
  assign n7018 = ~pi68  & n7017;
  assign n7019 = ~n7016 & ~n7018;
  assign n7020 = ~n6579 & ~n7019;
  assign n7021 = ~pi68  & ~n7015;
  assign n7022 = pi69  & ~n7021;
  assign n7023 = ~pi69  & n7021;
  assign n7024 = n6581 & ~n7015;
  assign n7025 = ~n7022 & ~n33153;
  assign n7026 = ~n33028 & ~n33096;
  assign n7027 = ~n6096 & n7026;
  assign n7028 = ~n6115 & n7027;
  assign n7029 = ~n33030 & n7028;
  assign n7030 = n6101 & n6117;
  assign n7031 = ~n6109 & n7029;
  assign n7032 = ~n7018 & ~n33154;
  assign n7033 = ~n6577 & n7032;
  assign n7034 = ~n33095 & n7033;
  assign n7035 = ~n6571 & n7034;
  assign n7036 = n6579 & n7019;
  assign n7037 = ~n7016 & n7035;
  assign n7038 = n7025 & ~n33155;
  assign n7039 = ~n7020 & ~n7038;
  assign n7040 = ~n6117 & ~n7039;
  assign n7041 = n6117 & ~n7020;
  assign n7042 = ~n7038 & n7041;
  assign n7043 = ~n6579 & ~n7013;
  assign n7044 = ~n33152 & n7043;
  assign n7045 = ~n7007 & n7044;
  assign n7046 = ~n33153 & ~n7045;
  assign n7047 = pi70  & ~n7046;
  assign n7048 = ~pi70  & ~n7045;
  assign n7049 = ~pi70  & n7046;
  assign n7050 = ~n33153 & n7048;
  assign n7051 = ~n7047 & ~n33156;
  assign n7052 = ~n7042 & ~n7051;
  assign n7053 = ~n7040 & ~n7052;
  assign n7054 = ~n5708 & ~n7053;
  assign n7055 = n5708 & ~n7040;
  assign n7056 = ~n7052 & n7055;
  assign n7057 = n5708 & n7053;
  assign n7058 = ~n6584 & ~n33097;
  assign n7059 = ~n7015 & n7058;
  assign n7060 = n6601 & ~n7059;
  assign n7061 = ~n6601 & n7058;
  assign n7062 = ~n6601 & n7059;
  assign n7063 = ~n7015 & n7061;
  assign n7064 = ~n7060 & ~n33158;
  assign n7065 = ~n33157 & ~n7064;
  assign n7066 = ~n7054 & ~n7065;
  assign n7067 = ~n5278 & ~n7066;
  assign n7068 = n5278 & ~n7054;
  assign n7069 = ~n7065 & n7068;
  assign n7070 = ~n6604 & ~n33100;
  assign n7071 = ~n6604 & ~n7015;
  assign n7072 = ~n33100 & n7071;
  assign n7073 = ~n7015 & n7070;
  assign n7074 = n6613 & ~n33159;
  assign n7075 = n6617 & n7071;
  assign n7076 = n6613 & ~n33100;
  assign n7077 = ~n6604 & n7076;
  assign n7078 = ~n7015 & n7077;
  assign n7079 = ~n6613 & ~n33159;
  assign n7080 = ~n7078 & ~n7079;
  assign n7081 = ~n7074 & ~n7075;
  assign n7082 = ~n7069 & ~n33160;
  assign n7083 = ~n7067 & ~n7082;
  assign n7084 = ~n4903 & ~n7083;
  assign n7085 = n4903 & ~n7067;
  assign n7086 = ~n7082 & n7085;
  assign n7087 = n4903 & n7083;
  assign n7088 = ~n6619 & ~n6621;
  assign n7089 = ~n7015 & n7088;
  assign n7090 = n6628 & ~n7089;
  assign n7091 = ~n6628 & n7089;
  assign n7092 = ~n6619 & n6628;
  assign n7093 = ~n6621 & n7092;
  assign n7094 = n6628 & n7089;
  assign n7095 = ~n7015 & n7093;
  assign n7096 = ~n6628 & ~n7089;
  assign n7097 = ~n33162 & ~n7096;
  assign n7098 = ~n7090 & ~n7091;
  assign n7099 = ~n33161 & ~n33163;
  assign n7100 = ~n7084 & ~n7099;
  assign n7101 = ~n4508 & ~n7100;
  assign n7102 = n4508 & ~n7084;
  assign n7103 = ~n7099 & n7102;
  assign n7104 = ~n6631 & ~n33103;
  assign n7105 = ~n6631 & ~n7015;
  assign n7106 = ~n33103 & n7105;
  assign n7107 = ~n7015 & n7104;
  assign n7108 = n6639 & ~n33164;
  assign n7109 = n6643 & n7105;
  assign n7110 = n6639 & ~n33103;
  assign n7111 = ~n6631 & n7110;
  assign n7112 = ~n7015 & n7111;
  assign n7113 = ~n6639 & ~n33164;
  assign n7114 = ~n7112 & ~n7113;
  assign n7115 = ~n7108 & ~n7109;
  assign n7116 = ~n7103 & ~n33165;
  assign n7117 = ~n7101 & ~n7116;
  assign n7118 = ~n4155 & ~n7117;
  assign n7119 = n4155 & ~n7101;
  assign n7120 = ~n7116 & n7119;
  assign n7121 = n4155 & n7117;
  assign n7122 = ~n6645 & ~n6647;
  assign n7123 = ~n7015 & n7122;
  assign n7124 = ~n33105 & n7123;
  assign n7125 = n33105 & ~n7123;
  assign n7126 = ~n6645 & n33105;
  assign n7127 = ~n6647 & n7126;
  assign n7128 = ~n7015 & n7127;
  assign n7129 = ~n33105 & ~n7123;
  assign n7130 = ~n7128 & ~n7129;
  assign n7131 = ~n7124 & ~n7125;
  assign n7132 = ~n33166 & ~n33167;
  assign n7133 = ~n7118 & ~n7132;
  assign n7134 = ~n3788 & ~n7133;
  assign n7135 = n3788 & ~n7118;
  assign n7136 = ~n7132 & n7135;
  assign n7137 = ~n6661 & ~n33107;
  assign n7138 = ~n6661 & ~n7015;
  assign n7139 = ~n33107 & n7138;
  assign n7140 = ~n7015 & n7137;
  assign n7141 = n6669 & ~n33168;
  assign n7142 = n6673 & n7138;
  assign n7143 = n6669 & ~n33107;
  assign n7144 = ~n6661 & n7143;
  assign n7145 = ~n7015 & n7144;
  assign n7146 = ~n6669 & ~n33168;
  assign n7147 = ~n7145 & ~n7146;
  assign n7148 = ~n7141 & ~n7142;
  assign n7149 = ~n7136 & ~n33169;
  assign n7150 = ~n7134 & ~n7149;
  assign n7151 = ~n3473 & ~n7150;
  assign n7152 = n3473 & ~n7134;
  assign n7153 = ~n7149 & n7152;
  assign n7154 = n3473 & n7150;
  assign n7155 = ~n6675 & ~n6677;
  assign n7156 = ~n7015 & n7155;
  assign n7157 = ~n33108 & ~n7156;
  assign n7158 = ~n6675 & n33108;
  assign n7159 = ~n6677 & n7158;
  assign n7160 = n33108 & n7156;
  assign n7161 = ~n7015 & n7159;
  assign n7162 = n33108 & ~n7156;
  assign n7163 = ~n33108 & n7156;
  assign n7164 = ~n7162 & ~n7163;
  assign n7165 = ~n7157 & ~n33171;
  assign n7166 = ~n33170 & n33172;
  assign n7167 = ~n7151 & ~n7166;
  assign n7168 = ~n3140 & ~n7167;
  assign n7169 = n3140 & ~n7151;
  assign n7170 = ~n7166 & n7169;
  assign n7171 = ~n6690 & ~n33110;
  assign n7172 = ~n6690 & ~n7015;
  assign n7173 = ~n33110 & n7172;
  assign n7174 = ~n7015 & n7171;
  assign n7175 = n6698 & ~n33173;
  assign n7176 = n6702 & n7172;
  assign n7177 = n6698 & ~n33110;
  assign n7178 = ~n6690 & n7177;
  assign n7179 = ~n7015 & n7178;
  assign n7180 = ~n6698 & ~n33173;
  assign n7181 = ~n7179 & ~n7180;
  assign n7182 = ~n7175 & ~n7176;
  assign n7183 = ~n7170 & ~n33174;
  assign n7184 = ~n7168 & ~n7183;
  assign n7185 = ~n2855 & ~n7184;
  assign n7186 = n2855 & ~n7168;
  assign n7187 = ~n7183 & n7186;
  assign n7188 = n2855 & n7184;
  assign n7189 = ~n6704 & ~n6706;
  assign n7190 = ~n7015 & n7189;
  assign n7191 = n33112 & ~n7190;
  assign n7192 = ~n6704 & ~n33112;
  assign n7193 = ~n6706 & n7192;
  assign n7194 = ~n33112 & n7190;
  assign n7195 = ~n7015 & n7193;
  assign n7196 = n33112 & n7190;
  assign n7197 = ~n33112 & ~n7190;
  assign n7198 = ~n7196 & ~n7197;
  assign n7199 = ~n7191 & ~n33176;
  assign n7200 = ~n33175 & n33177;
  assign n7201 = ~n7185 & ~n7200;
  assign n7202 = ~n2556 & ~n7201;
  assign n7203 = n2556 & ~n7185;
  assign n7204 = ~n7200 & n7203;
  assign n7205 = ~n6720 & ~n33114;
  assign n7206 = ~n6720 & ~n7015;
  assign n7207 = ~n33114 & n7206;
  assign n7208 = ~n7015 & n7205;
  assign n7209 = n6728 & ~n33178;
  assign n7210 = n6732 & n7206;
  assign n7211 = n6728 & ~n33114;
  assign n7212 = ~n6720 & n7211;
  assign n7213 = ~n7015 & n7212;
  assign n7214 = ~n6728 & ~n33178;
  assign n7215 = ~n7213 & ~n7214;
  assign n7216 = ~n7209 & ~n7210;
  assign n7217 = ~n7204 & ~n33179;
  assign n7218 = ~n7202 & ~n7217;
  assign n7219 = ~n2301 & ~n7218;
  assign n7220 = n2301 & ~n7202;
  assign n7221 = ~n7217 & n7220;
  assign n7222 = n2301 & n7218;
  assign n7223 = ~n6734 & ~n6736;
  assign n7224 = ~n6734 & ~n7015;
  assign n7225 = ~n6736 & n7224;
  assign n7226 = ~n7015 & n7223;
  assign n7227 = ~n33116 & ~n33181;
  assign n7228 = n6748 & n7224;
  assign n7229 = n33116 & n33181;
  assign n7230 = ~n6734 & ~n33116;
  assign n7231 = ~n6736 & n7230;
  assign n7232 = ~n7015 & n7231;
  assign n7233 = n33116 & ~n33181;
  assign n7234 = ~n7232 & ~n7233;
  assign n7235 = ~n7227 & ~n33182;
  assign n7236 = ~n33180 & ~n33183;
  assign n7237 = ~n7219 & ~n7236;
  assign n7238 = ~n2038 & ~n7237;
  assign n7239 = n2038 & ~n7219;
  assign n7240 = ~n7236 & n7239;
  assign n7241 = ~n6750 & ~n33118;
  assign n7242 = ~n6750 & ~n7015;
  assign n7243 = ~n33118 & n7242;
  assign n7244 = ~n7015 & n7241;
  assign n7245 = n6758 & ~n33184;
  assign n7246 = n6762 & n7242;
  assign n7247 = n6758 & ~n33118;
  assign n7248 = ~n6750 & n7247;
  assign n7249 = ~n7015 & n7248;
  assign n7250 = ~n6758 & ~n33184;
  assign n7251 = ~n7249 & ~n7250;
  assign n7252 = ~n7245 & ~n7246;
  assign n7253 = ~n7240 & ~n33185;
  assign n7254 = ~n7238 & ~n7253;
  assign n7255 = ~n1812 & ~n7254;
  assign n7256 = n1812 & ~n7238;
  assign n7257 = ~n7253 & n7256;
  assign n7258 = n1812 & n7254;
  assign n7259 = ~n6764 & ~n6766;
  assign n7260 = ~n7015 & n7259;
  assign n7261 = ~n33121 & ~n7260;
  assign n7262 = ~n6764 & n33121;
  assign n7263 = ~n6766 & n7262;
  assign n7264 = n33121 & n7260;
  assign n7265 = ~n7015 & n7263;
  assign n7266 = ~n7261 & ~n33187;
  assign n7267 = ~n33186 & ~n7266;
  assign n7268 = ~n7255 & ~n7267;
  assign n7269 = ~n1582 & ~n7268;
  assign n7270 = n1582 & ~n7255;
  assign n7271 = ~n7267 & n7270;
  assign n7272 = ~n6782 & ~n33123;
  assign n7273 = ~n6782 & ~n7015;
  assign n7274 = ~n33123 & n7273;
  assign n7275 = ~n7015 & n7272;
  assign n7276 = n6790 & ~n33188;
  assign n7277 = n6794 & n7273;
  assign n7278 = n6790 & ~n33123;
  assign n7279 = ~n6782 & n7278;
  assign n7280 = ~n7015 & n7279;
  assign n7281 = ~n6790 & ~n33188;
  assign n7282 = ~n7280 & ~n7281;
  assign n7283 = ~n7276 & ~n7277;
  assign n7284 = ~n7271 & ~n33189;
  assign n7285 = ~n7269 & ~n7284;
  assign n7286 = ~n1388 & ~n7285;
  assign n7287 = n1388 & ~n7269;
  assign n7288 = ~n7284 & n7287;
  assign n7289 = n1388 & n7285;
  assign n7290 = ~n6796 & ~n6798;
  assign n7291 = ~n6796 & ~n7015;
  assign n7292 = ~n6798 & n7291;
  assign n7293 = ~n7015 & n7290;
  assign n7294 = n6806 & ~n33191;
  assign n7295 = n6807 & n7291;
  assign n7296 = ~n6806 & n33191;
  assign n7297 = ~n6796 & n6806;
  assign n7298 = ~n6798 & n7297;
  assign n7299 = ~n7015 & n7298;
  assign n7300 = ~n6806 & ~n33191;
  assign n7301 = ~n7299 & ~n7300;
  assign n7302 = ~n7294 & ~n33192;
  assign n7303 = ~n33190 & ~n33193;
  assign n7304 = ~n7286 & ~n7303;
  assign n7305 = ~n1192 & ~n7304;
  assign n7306 = n1192 & ~n7286;
  assign n7307 = ~n7303 & n7306;
  assign n7308 = ~n6809 & ~n33126;
  assign n7309 = ~n6809 & ~n7015;
  assign n7310 = ~n33126 & n7309;
  assign n7311 = ~n7015 & n7308;
  assign n7312 = n6817 & ~n33194;
  assign n7313 = n6821 & n7309;
  assign n7314 = n6817 & ~n33126;
  assign n7315 = ~n6809 & n7314;
  assign n7316 = ~n7015 & n7315;
  assign n7317 = ~n6817 & ~n33194;
  assign n7318 = ~n7316 & ~n7317;
  assign n7319 = ~n7312 & ~n7313;
  assign n7320 = ~n7307 & ~n33195;
  assign n7321 = ~n7305 & ~n7320;
  assign n7322 = ~n1028 & ~n7321;
  assign n7323 = n1028 & ~n7305;
  assign n7324 = ~n7320 & n7323;
  assign n7325 = n1028 & n7321;
  assign n7326 = ~n6823 & ~n6825;
  assign n7327 = ~n7015 & n7326;
  assign n7328 = ~n33129 & n7327;
  assign n7329 = n33129 & ~n7327;
  assign n7330 = ~n6823 & n33129;
  assign n7331 = ~n6825 & n7330;
  assign n7332 = n33129 & n7327;
  assign n7333 = ~n7015 & n7331;
  assign n7334 = ~n33129 & ~n7327;
  assign n7335 = ~n33197 & ~n7334;
  assign n7336 = ~n7328 & ~n7329;
  assign n7337 = ~n33196 & ~n33198;
  assign n7338 = ~n7322 & ~n7337;
  assign n7339 = ~n866 & ~n7338;
  assign n7340 = n866 & ~n7322;
  assign n7341 = ~n7337 & n7340;
  assign n7342 = ~n6841 & ~n33131;
  assign n7343 = ~n6841 & ~n7015;
  assign n7344 = ~n33131 & n7343;
  assign n7345 = ~n7015 & n7342;
  assign n7346 = n6849 & ~n33199;
  assign n7347 = n6853 & n7343;
  assign n7348 = n6849 & ~n33131;
  assign n7349 = ~n6841 & n7348;
  assign n7350 = ~n7015 & n7349;
  assign n7351 = ~n6849 & ~n33199;
  assign n7352 = ~n7350 & ~n7351;
  assign n7353 = ~n7346 & ~n7347;
  assign n7354 = ~n7341 & ~n33200;
  assign n7355 = ~n7339 & ~n7354;
  assign n7356 = ~n730 & ~n7355;
  assign n7357 = n730 & ~n7339;
  assign n7358 = ~n7354 & n7357;
  assign n7359 = n730 & n7355;
  assign n7360 = ~n6855 & ~n6857;
  assign n7361 = ~n6855 & ~n7015;
  assign n7362 = ~n6857 & n7361;
  assign n7363 = ~n7015 & n7360;
  assign n7364 = n33133 & ~n33202;
  assign n7365 = n6869 & n7361;
  assign n7366 = ~n33133 & n33202;
  assign n7367 = ~n6855 & n33133;
  assign n7368 = ~n6857 & n7367;
  assign n7369 = ~n7015 & n7368;
  assign n7370 = ~n33133 & ~n33202;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = ~n7364 & ~n33203;
  assign n7373 = ~n33201 & ~n33204;
  assign n7374 = ~n7356 & ~n7373;
  assign n7375 = ~n602 & ~n7374;
  assign n7376 = n602 & ~n7356;
  assign n7377 = ~n7373 & n7376;
  assign n7378 = ~n6871 & ~n33135;
  assign n7379 = ~n6871 & ~n7015;
  assign n7380 = ~n33135 & n7379;
  assign n7381 = ~n7015 & n7378;
  assign n7382 = n6879 & ~n33205;
  assign n7383 = n6883 & n7379;
  assign n7384 = n6879 & ~n33135;
  assign n7385 = ~n6871 & n7384;
  assign n7386 = ~n7015 & n7385;
  assign n7387 = ~n6879 & ~n33205;
  assign n7388 = ~n7386 & ~n7387;
  assign n7389 = ~n7382 & ~n7383;
  assign n7390 = ~n7377 & ~n33206;
  assign n7391 = ~n7375 & ~n7390;
  assign n7392 = ~n497 & ~n7391;
  assign n7393 = ~n6885 & ~n6887;
  assign n7394 = ~n7015 & n7393;
  assign n7395 = ~n33138 & ~n7394;
  assign n7396 = ~n6885 & n33138;
  assign n7397 = ~n6887 & n7396;
  assign n7398 = n33138 & n7394;
  assign n7399 = ~n7015 & n7397;
  assign n7400 = ~n7395 & ~n33207;
  assign n7401 = n497 & ~n7375;
  assign n7402 = ~n7390 & n7401;
  assign n7403 = n497 & n7391;
  assign n7404 = ~n7400 & ~n33208;
  assign n7405 = ~n7392 & ~n7404;
  assign n7406 = ~n403 & ~n7405;
  assign n7407 = n403 & ~n7392;
  assign n7408 = ~n7404 & n7407;
  assign n7409 = ~n6903 & ~n33140;
  assign n7410 = ~n6903 & ~n7015;
  assign n7411 = ~n33140 & n7410;
  assign n7412 = ~n7015 & n7409;
  assign n7413 = n6911 & ~n33209;
  assign n7414 = n6915 & n7410;
  assign n7415 = n6911 & ~n33140;
  assign n7416 = ~n6903 & n7415;
  assign n7417 = ~n7015 & n7416;
  assign n7418 = ~n6911 & ~n33209;
  assign n7419 = ~n7417 & ~n7418;
  assign n7420 = ~n7413 & ~n7414;
  assign n7421 = ~n7408 & ~n33210;
  assign n7422 = ~n7406 & ~n7421;
  assign n7423 = ~n330 & ~n7422;
  assign n7424 = n330 & ~n7406;
  assign n7425 = ~n7421 & n7424;
  assign n7426 = n330 & n7422;
  assign n7427 = ~n6917 & ~n6927;
  assign n7428 = ~n6917 & ~n7015;
  assign n7429 = ~n6927 & n7428;
  assign n7430 = ~n7015 & n7427;
  assign n7431 = n6925 & ~n33212;
  assign n7432 = n6928 & n7428;
  assign n7433 = ~n6917 & n6925;
  assign n7434 = ~n6927 & n7433;
  assign n7435 = ~n7015 & n7434;
  assign n7436 = ~n6925 & ~n33212;
  assign n7437 = ~n7435 & ~n7436;
  assign n7438 = ~n7431 & ~n7432;
  assign n7439 = ~n33211 & ~n33213;
  assign n7440 = ~n7423 & ~n7439;
  assign n7441 = ~n271 & ~n7440;
  assign n7442 = n271 & ~n7423;
  assign n7443 = ~n7439 & n7442;
  assign n7444 = ~n6930 & ~n33143;
  assign n7445 = ~n6930 & ~n7015;
  assign n7446 = ~n33143 & n7445;
  assign n7447 = ~n7015 & n7444;
  assign n7448 = n6938 & ~n33214;
  assign n7449 = n6942 & n7445;
  assign n7450 = n6938 & ~n33143;
  assign n7451 = ~n6930 & n7450;
  assign n7452 = ~n7015 & n7451;
  assign n7453 = ~n6938 & ~n33214;
  assign n7454 = ~n7452 & ~n7453;
  assign n7455 = ~n7448 & ~n7449;
  assign n7456 = ~n7443 & ~n33215;
  assign n7457 = ~n7441 & ~n7456;
  assign n7458 = ~n217 & ~n7457;
  assign n7459 = ~n6944 & ~n6946;
  assign n7460 = ~n7015 & n7459;
  assign n7461 = ~n33145 & ~n7460;
  assign n7462 = ~n6944 & n33145;
  assign n7463 = ~n6946 & n7462;
  assign n7464 = n33145 & n7460;
  assign n7465 = ~n7015 & n7463;
  assign n7466 = ~n7461 & ~n33216;
  assign n7467 = n217 & ~n7441;
  assign n7468 = ~n7456 & n7467;
  assign n7469 = n217 & n7457;
  assign n7470 = ~n7466 & ~n33217;
  assign n7471 = ~n7458 & ~n7470;
  assign n7472 = ~n198 & ~n7471;
  assign n7473 = n198 & ~n7458;
  assign n7474 = ~n7470 & n7473;
  assign n7475 = ~n6961 & ~n33147;
  assign n7476 = ~n6961 & ~n7015;
  assign n7477 = ~n33147 & n7476;
  assign n7478 = ~n7015 & n7475;
  assign n7479 = n6969 & ~n33218;
  assign n7480 = n6973 & n7476;
  assign n7481 = n6969 & ~n33147;
  assign n7482 = ~n6961 & n7481;
  assign n7483 = ~n7015 & n7482;
  assign n7484 = ~n6969 & ~n33218;
  assign n7485 = ~n7483 & ~n7484;
  assign n7486 = ~n7479 & ~n7480;
  assign n7487 = ~n7474 & ~n33219;
  assign n7488 = ~n7472 & ~n7487;
  assign n7489 = ~n6975 & ~n6977;
  assign n7490 = ~n7015 & n7489;
  assign n7491 = ~n33149 & ~n7490;
  assign n7492 = ~n6975 & n33149;
  assign n7493 = ~n6977 & n7492;
  assign n7494 = n33149 & n7490;
  assign n7495 = ~n7015 & n7493;
  assign n7496 = ~n7491 & ~n33220;
  assign n7497 = ~n6991 & ~n6999;
  assign n7498 = ~n6999 & ~n7015;
  assign n7499 = ~n6991 & n7498;
  assign n7500 = ~n7015 & n7497;
  assign n7501 = ~n33152 & ~n33221;
  assign n7502 = ~n7496 & n7501;
  assign n7503 = ~n7488 & n7502;
  assign n7504 = n193 & ~n7503;
  assign n7505 = ~n7472 & n7496;
  assign n7506 = ~n7487 & n7505;
  assign n7507 = n7488 & n7496;
  assign n7508 = n6991 & ~n7498;
  assign n7509 = ~n193 & ~n7497;
  assign n7510 = ~n7508 & n7509;
  assign n7511 = ~n33222 & ~n7510;
  assign n7512 = ~n7504 & n7511;
  assign n7513 = pi66  & ~n7512;
  assign n7514 = ~pi64  & ~pi65 ;
  assign n7515 = ~pi66  & n7514;
  assign n7516 = ~n7513 & ~n7515;
  assign n7517 = ~n7015 & ~n7516;
  assign n7518 = ~n33093 & ~n33154;
  assign n7519 = ~n6558 & n7518;
  assign n7520 = ~n6577 & n7519;
  assign n7521 = ~n33095 & n7520;
  assign n7522 = n6563 & n6579;
  assign n7523 = ~n6571 & n7521;
  assign n7524 = ~n7515 & ~n33223;
  assign n7525 = ~n7013 & n7524;
  assign n7526 = ~n33152 & n7525;
  assign n7527 = ~n7007 & n7526;
  assign n7528 = n7015 & n7516;
  assign n7529 = ~n7513 & n7527;
  assign n7530 = ~pi66  & ~n7512;
  assign n7531 = pi67  & ~n7530;
  assign n7532 = ~pi67  & n7530;
  assign n7533 = n7017 & ~n7512;
  assign n7534 = ~n7531 & ~n33225;
  assign n7535 = ~n33224 & n7534;
  assign n7536 = ~n7517 & ~n7535;
  assign n7537 = ~n6579 & ~n7536;
  assign n7538 = ~n7015 & ~n7510;
  assign n7539 = ~n33222 & n7538;
  assign n7540 = ~n7504 & n7539;
  assign n7541 = ~n33225 & ~n7540;
  assign n7542 = pi68  & ~n7541;
  assign n7543 = ~pi68  & ~n7540;
  assign n7544 = ~pi68  & n7541;
  assign n7545 = ~n33225 & n7543;
  assign n7546 = ~n7542 & ~n33226;
  assign n7547 = n6579 & ~n7517;
  assign n7548 = n6579 & n7536;
  assign n7549 = ~n7535 & n7547;
  assign n7550 = ~n7546 & ~n33227;
  assign n7551 = ~n7537 & ~n7550;
  assign n7552 = ~n6117 & ~n7551;
  assign n7553 = n6117 & ~n7537;
  assign n7554 = ~n7550 & n7553;
  assign n7555 = ~n7020 & ~n33155;
  assign n7556 = ~n7512 & n7555;
  assign n7557 = n7025 & ~n7556;
  assign n7558 = ~n7025 & n7555;
  assign n7559 = ~n7025 & n7556;
  assign n7560 = ~n7512 & n7558;
  assign n7561 = ~n7557 & ~n33228;
  assign n7562 = ~n7554 & ~n7561;
  assign n7563 = ~n7552 & ~n7562;
  assign n7564 = ~n5708 & ~n7563;
  assign n7565 = ~n7040 & ~n7042;
  assign n7566 = ~n7512 & n7565;
  assign n7567 = ~n7051 & ~n7566;
  assign n7568 = ~n7042 & n7051;
  assign n7569 = ~n7040 & n7568;
  assign n7570 = n7051 & n7566;
  assign n7571 = ~n7512 & n7569;
  assign n7572 = ~n7567 & ~n33229;
  assign n7573 = n5708 & ~n7552;
  assign n7574 = n5708 & n7563;
  assign n7575 = ~n7562 & n7573;
  assign n7576 = ~n7572 & ~n33230;
  assign n7577 = ~n7564 & ~n7576;
  assign n7578 = ~n5278 & ~n7577;
  assign n7579 = n5278 & ~n7564;
  assign n7580 = ~n7576 & n7579;
  assign n7581 = ~n7054 & ~n33157;
  assign n7582 = ~n7512 & n7581;
  assign n7583 = n7064 & ~n7582;
  assign n7584 = ~n7064 & n7582;
  assign n7585 = ~n7054 & n7064;
  assign n7586 = ~n33157 & n7585;
  assign n7587 = n7064 & n7582;
  assign n7588 = ~n7512 & n7586;
  assign n7589 = ~n7064 & ~n7582;
  assign n7590 = ~n33231 & ~n7589;
  assign n7591 = ~n7583 & ~n7584;
  assign n7592 = ~n7580 & ~n33232;
  assign n7593 = ~n7578 & ~n7592;
  assign n7594 = ~n4903 & ~n7593;
  assign n7595 = ~n7067 & ~n7069;
  assign n7596 = ~n7512 & n7595;
  assign n7597 = ~n33160 & ~n7596;
  assign n7598 = ~n7069 & n33160;
  assign n7599 = ~n7067 & n7598;
  assign n7600 = n33160 & n7596;
  assign n7601 = ~n7512 & n7599;
  assign n7602 = ~n7597 & ~n33233;
  assign n7603 = n4903 & ~n7578;
  assign n7604 = n4903 & n7593;
  assign n7605 = ~n7592 & n7603;
  assign n7606 = ~n7602 & ~n33234;
  assign n7607 = ~n7594 & ~n7606;
  assign n7608 = ~n4508 & ~n7607;
  assign n7609 = n4508 & ~n7594;
  assign n7610 = ~n7606 & n7609;
  assign n7611 = ~n7084 & ~n33161;
  assign n7612 = ~n7512 & n7611;
  assign n7613 = ~n33163 & n7612;
  assign n7614 = n33163 & ~n7612;
  assign n7615 = ~n7084 & n33163;
  assign n7616 = ~n33161 & n7615;
  assign n7617 = ~n7512 & n7616;
  assign n7618 = ~n33163 & ~n7612;
  assign n7619 = ~n7617 & ~n7618;
  assign n7620 = ~n7613 & ~n7614;
  assign n7621 = ~n7610 & ~n33235;
  assign n7622 = ~n7608 & ~n7621;
  assign n7623 = ~n4155 & ~n7622;
  assign n7624 = ~n7101 & ~n7103;
  assign n7625 = ~n7512 & n7624;
  assign n7626 = ~n33165 & ~n7625;
  assign n7627 = ~n7103 & n33165;
  assign n7628 = ~n7101 & n7627;
  assign n7629 = n33165 & n7625;
  assign n7630 = ~n7512 & n7628;
  assign n7631 = ~n7626 & ~n33236;
  assign n7632 = n4155 & ~n7608;
  assign n7633 = n4155 & n7622;
  assign n7634 = ~n7621 & n7632;
  assign n7635 = ~n7631 & ~n33237;
  assign n7636 = ~n7623 & ~n7635;
  assign n7637 = ~n3788 & ~n7636;
  assign n7638 = n3788 & ~n7623;
  assign n7639 = ~n7635 & n7638;
  assign n7640 = ~n7118 & ~n33166;
  assign n7641 = ~n7512 & n7640;
  assign n7642 = ~n33167 & ~n7641;
  assign n7643 = ~n7118 & n33167;
  assign n7644 = ~n33166 & n7643;
  assign n7645 = n33167 & n7641;
  assign n7646 = ~n7512 & n7644;
  assign n7647 = n33167 & ~n7641;
  assign n7648 = ~n33167 & n7641;
  assign n7649 = ~n7647 & ~n7648;
  assign n7650 = ~n7642 & ~n33238;
  assign n7651 = ~n7639 & n33239;
  assign n7652 = ~n7637 & ~n7651;
  assign n7653 = ~n3473 & ~n7652;
  assign n7654 = ~n7134 & ~n7136;
  assign n7655 = ~n7512 & n7654;
  assign n7656 = ~n33169 & ~n7655;
  assign n7657 = ~n7136 & n33169;
  assign n7658 = ~n7134 & n7657;
  assign n7659 = n33169 & n7655;
  assign n7660 = ~n7512 & n7658;
  assign n7661 = ~n7656 & ~n33240;
  assign n7662 = n3473 & ~n7637;
  assign n7663 = n3473 & n7652;
  assign n7664 = ~n7651 & n7662;
  assign n7665 = ~n7661 & ~n33241;
  assign n7666 = ~n7653 & ~n7665;
  assign n7667 = ~n3140 & ~n7666;
  assign n7668 = n3140 & ~n7653;
  assign n7669 = ~n7665 & n7668;
  assign n7670 = ~n7151 & ~n33170;
  assign n7671 = ~n7512 & n7670;
  assign n7672 = n33172 & ~n7671;
  assign n7673 = ~n7151 & ~n33172;
  assign n7674 = ~n33170 & n7673;
  assign n7675 = ~n33172 & n7671;
  assign n7676 = ~n7512 & n7674;
  assign n7677 = n33172 & n7671;
  assign n7678 = ~n33172 & ~n7671;
  assign n7679 = ~n7677 & ~n7678;
  assign n7680 = ~n7672 & ~n33242;
  assign n7681 = ~n7669 & n33243;
  assign n7682 = ~n7667 & ~n7681;
  assign n7683 = ~n2855 & ~n7682;
  assign n7684 = ~n7168 & ~n7170;
  assign n7685 = ~n7512 & n7684;
  assign n7686 = ~n33174 & ~n7685;
  assign n7687 = ~n7170 & n33174;
  assign n7688 = ~n7168 & n7687;
  assign n7689 = n33174 & n7685;
  assign n7690 = ~n7512 & n7688;
  assign n7691 = ~n7686 & ~n33244;
  assign n7692 = n2855 & ~n7667;
  assign n7693 = n2855 & n7682;
  assign n7694 = ~n7681 & n7692;
  assign n7695 = ~n7691 & ~n33245;
  assign n7696 = ~n7683 & ~n7695;
  assign n7697 = ~n2556 & ~n7696;
  assign n7698 = n2556 & ~n7683;
  assign n7699 = ~n7695 & n7698;
  assign n7700 = ~n7185 & ~n33175;
  assign n7701 = ~n7185 & ~n7512;
  assign n7702 = ~n33175 & n7701;
  assign n7703 = ~n7512 & n7700;
  assign n7704 = ~n33177 & ~n33246;
  assign n7705 = n7200 & n7701;
  assign n7706 = n33177 & n33246;
  assign n7707 = ~n7185 & ~n33177;
  assign n7708 = ~n33175 & n7707;
  assign n7709 = ~n7512 & n7708;
  assign n7710 = n33177 & ~n33246;
  assign n7711 = ~n7709 & ~n7710;
  assign n7712 = ~n7704 & ~n33247;
  assign n7713 = ~n7699 & ~n33248;
  assign n7714 = ~n7697 & ~n7713;
  assign n7715 = ~n2301 & ~n7714;
  assign n7716 = ~n7202 & ~n7204;
  assign n7717 = ~n7512 & n7716;
  assign n7718 = ~n33179 & ~n7717;
  assign n7719 = ~n7204 & n33179;
  assign n7720 = ~n7202 & n7719;
  assign n7721 = n33179 & n7717;
  assign n7722 = ~n7512 & n7720;
  assign n7723 = ~n7718 & ~n33249;
  assign n7724 = n2301 & ~n7697;
  assign n7725 = n2301 & n7714;
  assign n7726 = ~n7713 & n7724;
  assign n7727 = ~n7723 & ~n33250;
  assign n7728 = ~n7715 & ~n7727;
  assign n7729 = ~n2038 & ~n7728;
  assign n7730 = n2038 & ~n7715;
  assign n7731 = ~n7727 & n7730;
  assign n7732 = ~n7219 & ~n33180;
  assign n7733 = ~n7512 & n7732;
  assign n7734 = ~n33183 & ~n7733;
  assign n7735 = ~n7219 & n33183;
  assign n7736 = ~n33180 & n7735;
  assign n7737 = n33183 & n7733;
  assign n7738 = ~n7512 & n7736;
  assign n7739 = ~n7734 & ~n33251;
  assign n7740 = ~n7731 & ~n7739;
  assign n7741 = ~n7729 & ~n7740;
  assign n7742 = ~n1812 & ~n7741;
  assign n7743 = ~n7238 & ~n7240;
  assign n7744 = ~n7512 & n7743;
  assign n7745 = ~n33185 & ~n7744;
  assign n7746 = ~n7240 & n33185;
  assign n7747 = ~n7238 & n7746;
  assign n7748 = n33185 & n7744;
  assign n7749 = ~n7512 & n7747;
  assign n7750 = ~n7745 & ~n33252;
  assign n7751 = n1812 & ~n7729;
  assign n7752 = n1812 & n7741;
  assign n7753 = ~n7740 & n7751;
  assign n7754 = ~n7750 & ~n33253;
  assign n7755 = ~n7742 & ~n7754;
  assign n7756 = ~n1582 & ~n7755;
  assign n7757 = n1582 & ~n7742;
  assign n7758 = ~n7754 & n7757;
  assign n7759 = ~n7255 & ~n33186;
  assign n7760 = ~n7255 & ~n7512;
  assign n7761 = ~n33186 & n7760;
  assign n7762 = ~n7512 & n7759;
  assign n7763 = n7266 & ~n33254;
  assign n7764 = n7267 & n7760;
  assign n7765 = ~n7266 & n33254;
  assign n7766 = ~n7255 & n7266;
  assign n7767 = ~n33186 & n7766;
  assign n7768 = ~n7512 & n7767;
  assign n7769 = ~n7266 & ~n33254;
  assign n7770 = ~n7768 & ~n7769;
  assign n7771 = ~n7763 & ~n33255;
  assign n7772 = ~n7758 & ~n33256;
  assign n7773 = ~n7756 & ~n7772;
  assign n7774 = ~n1388 & ~n7773;
  assign n7775 = ~n7269 & ~n7271;
  assign n7776 = ~n7512 & n7775;
  assign n7777 = ~n33189 & ~n7776;
  assign n7778 = ~n7271 & n33189;
  assign n7779 = ~n7269 & n7778;
  assign n7780 = n33189 & n7776;
  assign n7781 = ~n7512 & n7779;
  assign n7782 = ~n7777 & ~n33257;
  assign n7783 = n1388 & ~n7756;
  assign n7784 = n1388 & n7773;
  assign n7785 = ~n7772 & n7783;
  assign n7786 = ~n7782 & ~n33258;
  assign n7787 = ~n7774 & ~n7786;
  assign n7788 = ~n1192 & ~n7787;
  assign n7789 = n1192 & ~n7774;
  assign n7790 = ~n7786 & n7789;
  assign n7791 = ~n7286 & ~n33190;
  assign n7792 = ~n7512 & n7791;
  assign n7793 = ~n33193 & n7792;
  assign n7794 = n33193 & ~n7792;
  assign n7795 = ~n7286 & n33193;
  assign n7796 = ~n33190 & n7795;
  assign n7797 = n33193 & n7792;
  assign n7798 = ~n7512 & n7796;
  assign n7799 = ~n33193 & ~n7792;
  assign n7800 = ~n33259 & ~n7799;
  assign n7801 = ~n7793 & ~n7794;
  assign n7802 = ~n7790 & ~n33260;
  assign n7803 = ~n7788 & ~n7802;
  assign n7804 = ~n1028 & ~n7803;
  assign n7805 = ~n7305 & ~n7307;
  assign n7806 = ~n7512 & n7805;
  assign n7807 = ~n33195 & ~n7806;
  assign n7808 = ~n7307 & n33195;
  assign n7809 = ~n7305 & n7808;
  assign n7810 = n33195 & n7806;
  assign n7811 = ~n7512 & n7809;
  assign n7812 = ~n7807 & ~n33261;
  assign n7813 = n1028 & ~n7788;
  assign n7814 = n1028 & n7803;
  assign n7815 = ~n7802 & n7813;
  assign n7816 = ~n7812 & ~n33262;
  assign n7817 = ~n7804 & ~n7816;
  assign n7818 = ~n866 & ~n7817;
  assign n7819 = n866 & ~n7804;
  assign n7820 = ~n7816 & n7819;
  assign n7821 = ~n7322 & ~n33196;
  assign n7822 = ~n7322 & ~n7512;
  assign n7823 = ~n33196 & n7822;
  assign n7824 = ~n7512 & n7821;
  assign n7825 = n33198 & ~n33263;
  assign n7826 = n7337 & n7822;
  assign n7827 = ~n33198 & n33263;
  assign n7828 = ~n7322 & n33198;
  assign n7829 = ~n33196 & n7828;
  assign n7830 = ~n7512 & n7829;
  assign n7831 = ~n33198 & ~n33263;
  assign n7832 = ~n7830 & ~n7831;
  assign n7833 = ~n7825 & ~n33264;
  assign n7834 = ~n7820 & ~n33265;
  assign n7835 = ~n7818 & ~n7834;
  assign n7836 = ~n730 & ~n7835;
  assign n7837 = ~n7339 & ~n7341;
  assign n7838 = ~n7512 & n7837;
  assign n7839 = ~n33200 & ~n7838;
  assign n7840 = ~n7341 & n33200;
  assign n7841 = ~n7339 & n7840;
  assign n7842 = n33200 & n7838;
  assign n7843 = ~n7512 & n7841;
  assign n7844 = ~n7839 & ~n33266;
  assign n7845 = n730 & ~n7818;
  assign n7846 = n730 & n7835;
  assign n7847 = ~n7834 & n7845;
  assign n7848 = ~n7844 & ~n33267;
  assign n7849 = ~n7836 & ~n7848;
  assign n7850 = ~n602 & ~n7849;
  assign n7851 = ~n7356 & ~n33201;
  assign n7852 = ~n7512 & n7851;
  assign n7853 = ~n33204 & ~n7852;
  assign n7854 = ~n7356 & n33204;
  assign n7855 = ~n33201 & n7854;
  assign n7856 = n33204 & n7852;
  assign n7857 = ~n7512 & n7855;
  assign n7858 = ~n7853 & ~n33268;
  assign n7859 = n602 & ~n7836;
  assign n7860 = ~n7848 & n7859;
  assign n7861 = ~n7858 & ~n7860;
  assign n7862 = ~n7850 & ~n7861;
  assign n7863 = ~n497 & ~n7862;
  assign n7864 = ~n7375 & ~n7377;
  assign n7865 = ~n7512 & n7864;
  assign n7866 = ~n33206 & ~n7865;
  assign n7867 = ~n7377 & n33206;
  assign n7868 = ~n7375 & n7867;
  assign n7869 = n33206 & n7865;
  assign n7870 = ~n7512 & n7868;
  assign n7871 = ~n7866 & ~n33269;
  assign n7872 = n497 & ~n7850;
  assign n7873 = n497 & n7862;
  assign n7874 = ~n7861 & n7872;
  assign n7875 = ~n7871 & ~n33270;
  assign n7876 = ~n7863 & ~n7875;
  assign n7877 = ~n403 & ~n7876;
  assign n7878 = n403 & ~n7863;
  assign n7879 = ~n7875 & n7878;
  assign n7880 = ~n7392 & ~n33208;
  assign n7881 = ~n7392 & ~n7512;
  assign n7882 = ~n33208 & n7881;
  assign n7883 = ~n7512 & n7880;
  assign n7884 = n7400 & ~n33271;
  assign n7885 = n7404 & n7881;
  assign n7886 = ~n7392 & n7400;
  assign n7887 = ~n33208 & n7886;
  assign n7888 = ~n7512 & n7887;
  assign n7889 = ~n7400 & ~n33271;
  assign n7890 = ~n7888 & ~n7889;
  assign n7891 = ~n7884 & ~n7885;
  assign n7892 = ~n7879 & ~n33272;
  assign n7893 = ~n7877 & ~n7892;
  assign n7894 = ~n330 & ~n7893;
  assign n7895 = ~n7406 & ~n7408;
  assign n7896 = ~n7512 & n7895;
  assign n7897 = ~n33210 & ~n7896;
  assign n7898 = ~n7408 & n33210;
  assign n7899 = ~n7406 & n7898;
  assign n7900 = n33210 & n7896;
  assign n7901 = ~n7512 & n7899;
  assign n7902 = ~n7897 & ~n33273;
  assign n7903 = n330 & ~n7877;
  assign n7904 = n330 & n7893;
  assign n7905 = ~n7892 & n7903;
  assign n7906 = ~n7902 & ~n33274;
  assign n7907 = ~n7894 & ~n7906;
  assign n7908 = ~n271 & ~n7907;
  assign n7909 = ~n7423 & ~n33211;
  assign n7910 = ~n7512 & n7909;
  assign n7911 = ~n33213 & ~n7910;
  assign n7912 = ~n7423 & n33213;
  assign n7913 = ~n33211 & n7912;
  assign n7914 = n33213 & n7910;
  assign n7915 = ~n7512 & n7913;
  assign n7916 = ~n7911 & ~n33275;
  assign n7917 = n271 & ~n7894;
  assign n7918 = ~n7906 & n7917;
  assign n7919 = ~n7916 & ~n7918;
  assign n7920 = ~n7908 & ~n7919;
  assign n7921 = ~n217 & ~n7920;
  assign n7922 = ~n7441 & ~n7443;
  assign n7923 = ~n7512 & n7922;
  assign n7924 = ~n33215 & ~n7923;
  assign n7925 = ~n7443 & n33215;
  assign n7926 = ~n7441 & n7925;
  assign n7927 = n33215 & n7923;
  assign n7928 = ~n7512 & n7926;
  assign n7929 = ~n7924 & ~n33276;
  assign n7930 = n217 & ~n7908;
  assign n7931 = n217 & n7920;
  assign n7932 = ~n7919 & n7930;
  assign n7933 = ~n7929 & ~n33277;
  assign n7934 = ~n7921 & ~n7933;
  assign n7935 = ~n198 & ~n7934;
  assign n7936 = n198 & ~n7921;
  assign n7937 = ~n7933 & n7936;
  assign n7938 = ~n7458 & ~n33217;
  assign n7939 = ~n7458 & ~n7512;
  assign n7940 = ~n33217 & n7939;
  assign n7941 = ~n7512 & n7938;
  assign n7942 = n7466 & ~n33278;
  assign n7943 = n7470 & n7939;
  assign n7944 = ~n7458 & n7466;
  assign n7945 = ~n33217 & n7944;
  assign n7946 = ~n7512 & n7945;
  assign n7947 = ~n7466 & ~n33278;
  assign n7948 = ~n7946 & ~n7947;
  assign n7949 = ~n7942 & ~n7943;
  assign n7950 = ~n7937 & ~n33279;
  assign n7951 = ~n7935 & ~n7950;
  assign n7952 = ~n7472 & ~n7474;
  assign n7953 = ~n7512 & n7952;
  assign n7954 = ~n33219 & ~n7953;
  assign n7955 = ~n7474 & n33219;
  assign n7956 = ~n7472 & n7955;
  assign n7957 = n33219 & n7953;
  assign n7958 = ~n7512 & n7956;
  assign n7959 = ~n7954 & ~n33280;
  assign n7960 = ~n7488 & ~n7496;
  assign n7961 = ~n7496 & ~n7512;
  assign n7962 = ~n7488 & n7961;
  assign n7963 = ~n7512 & n7960;
  assign n7964 = ~n33222 & ~n33281;
  assign n7965 = ~n7959 & n7964;
  assign n7966 = ~n7951 & n7965;
  assign n7967 = n193 & ~n7966;
  assign n7968 = ~n7935 & n7959;
  assign n7969 = n7951 & n7959;
  assign n7970 = ~n7950 & n7968;
  assign n7971 = n7488 & ~n7961;
  assign n7972 = ~n193 & ~n7960;
  assign n7973 = ~n7971 & n7972;
  assign n7974 = ~n33282 & ~n7973;
  assign n7975 = ~n7967 & n7974;
  assign n7976 = pi64  & ~n7975;
  assign n7977 = ~pi64  & n194;
  assign n7978 = ~n7976 & ~n7977;
  assign n7979 = ~n7512 & ~n7978;
  assign n7980 = ~pi64  & ~n7975;
  assign n7981 = pi65  & ~n7980;
  assign n7982 = ~pi65  & n7980;
  assign n7983 = n7514 & ~n7975;
  assign n7984 = ~n7981 & ~n33283;
  assign n7985 = ~n33150 & ~n33223;
  assign n7986 = ~n6994 & n7985;
  assign n7987 = ~n7013 & n7986;
  assign n7988 = ~n33152 & n7987;
  assign n7989 = n6999 & n7015;
  assign n7990 = ~n7007 & n7988;
  assign n7991 = ~n7977 & ~n33284;
  assign n7992 = ~n7510 & n7991;
  assign n7993 = ~n33222 & n7992;
  assign n7994 = ~n7504 & n7993;
  assign n7995 = n7512 & n7978;
  assign n7996 = ~n7976 & n7994;
  assign n7997 = n7984 & ~n33285;
  assign n7998 = ~n7979 & ~n7997;
  assign n7999 = ~n7015 & ~n7998;
  assign n8000 = n7015 & ~n7979;
  assign n8001 = ~n7997 & n8000;
  assign n8002 = ~n7512 & ~n7973;
  assign n8003 = ~n33282 & n8002;
  assign n8004 = ~n7967 & n8003;
  assign n8005 = ~n33283 & ~n8004;
  assign n8006 = pi66  & ~n8005;
  assign n8007 = ~pi66  & ~n8004;
  assign n8008 = ~pi66  & n8005;
  assign n8009 = ~n33283 & n8007;
  assign n8010 = ~n8006 & ~n33286;
  assign n8011 = ~n8001 & ~n8010;
  assign n8012 = ~n7999 & ~n8011;
  assign n8013 = ~n6579 & ~n8012;
  assign n8014 = n6579 & ~n7999;
  assign n8015 = ~n8011 & n8014;
  assign n8016 = n6579 & n8012;
  assign n8017 = ~n7517 & ~n33224;
  assign n8018 = ~n7975 & n8017;
  assign n8019 = n7534 & ~n8018;
  assign n8020 = ~n7534 & n8017;
  assign n8021 = ~n7534 & n8018;
  assign n8022 = ~n7975 & n8020;
  assign n8023 = ~n8019 & ~n33288;
  assign n8024 = ~n33287 & ~n8023;
  assign n8025 = ~n8013 & ~n8024;
  assign n8026 = ~n6117 & ~n8025;
  assign n8027 = n6117 & ~n8013;
  assign n8028 = ~n8024 & n8027;
  assign n8029 = ~n7537 & ~n33227;
  assign n8030 = ~n7537 & ~n7975;
  assign n8031 = ~n33227 & n8030;
  assign n8032 = ~n7975 & n8029;
  assign n8033 = n7546 & ~n33289;
  assign n8034 = n7550 & n8030;
  assign n8035 = n7546 & ~n33227;
  assign n8036 = ~n7537 & n8035;
  assign n8037 = ~n7975 & n8036;
  assign n8038 = ~n7546 & ~n33289;
  assign n8039 = ~n8037 & ~n8038;
  assign n8040 = ~n8033 & ~n8034;
  assign n8041 = ~n8028 & ~n33290;
  assign n8042 = ~n8026 & ~n8041;
  assign n8043 = ~n5708 & ~n8042;
  assign n8044 = n5708 & ~n8026;
  assign n8045 = ~n8041 & n8044;
  assign n8046 = n5708 & n8042;
  assign n8047 = ~n7552 & ~n7554;
  assign n8048 = ~n7975 & n8047;
  assign n8049 = n7561 & ~n8048;
  assign n8050 = ~n7561 & n8048;
  assign n8051 = ~n7552 & n7561;
  assign n8052 = ~n7554 & n8051;
  assign n8053 = n7561 & n8048;
  assign n8054 = ~n7975 & n8052;
  assign n8055 = ~n7561 & ~n8048;
  assign n8056 = ~n33292 & ~n8055;
  assign n8057 = ~n8049 & ~n8050;
  assign n8058 = ~n33291 & ~n33293;
  assign n8059 = ~n8043 & ~n8058;
  assign n8060 = ~n5278 & ~n8059;
  assign n8061 = n5278 & ~n8043;
  assign n8062 = ~n8058 & n8061;
  assign n8063 = ~n7564 & ~n33230;
  assign n8064 = ~n7564 & ~n7975;
  assign n8065 = ~n33230 & n8064;
  assign n8066 = ~n7975 & n8063;
  assign n8067 = n7572 & ~n33294;
  assign n8068 = n7576 & n8064;
  assign n8069 = n7572 & ~n33230;
  assign n8070 = ~n7564 & n8069;
  assign n8071 = ~n7975 & n8070;
  assign n8072 = ~n7572 & ~n33294;
  assign n8073 = ~n8071 & ~n8072;
  assign n8074 = ~n8067 & ~n8068;
  assign n8075 = ~n8062 & ~n33295;
  assign n8076 = ~n8060 & ~n8075;
  assign n8077 = ~n4903 & ~n8076;
  assign n8078 = n4903 & ~n8060;
  assign n8079 = ~n8075 & n8078;
  assign n8080 = n4903 & n8076;
  assign n8081 = ~n7578 & ~n7580;
  assign n8082 = ~n7975 & n8081;
  assign n8083 = ~n33232 & n8082;
  assign n8084 = n33232 & ~n8082;
  assign n8085 = ~n7578 & n33232;
  assign n8086 = ~n7580 & n8085;
  assign n8087 = ~n7975 & n8086;
  assign n8088 = ~n33232 & ~n8082;
  assign n8089 = ~n8087 & ~n8088;
  assign n8090 = ~n8083 & ~n8084;
  assign n8091 = ~n33296 & ~n33297;
  assign n8092 = ~n8077 & ~n8091;
  assign n8093 = ~n4508 & ~n8092;
  assign n8094 = n4508 & ~n8077;
  assign n8095 = ~n8091 & n8094;
  assign n8096 = ~n7594 & ~n33234;
  assign n8097 = ~n7594 & ~n7975;
  assign n8098 = ~n33234 & n8097;
  assign n8099 = ~n7975 & n8096;
  assign n8100 = n7602 & ~n33298;
  assign n8101 = n7606 & n8097;
  assign n8102 = n7602 & ~n33234;
  assign n8103 = ~n7594 & n8102;
  assign n8104 = ~n7975 & n8103;
  assign n8105 = ~n7602 & ~n33298;
  assign n8106 = ~n8104 & ~n8105;
  assign n8107 = ~n8100 & ~n8101;
  assign n8108 = ~n8095 & ~n33299;
  assign n8109 = ~n8093 & ~n8108;
  assign n8110 = ~n4155 & ~n8109;
  assign n8111 = n4155 & ~n8093;
  assign n8112 = ~n8108 & n8111;
  assign n8113 = n4155 & n8109;
  assign n8114 = ~n7608 & ~n7610;
  assign n8115 = ~n7975 & n8114;
  assign n8116 = ~n33235 & ~n8115;
  assign n8117 = ~n7608 & n33235;
  assign n8118 = ~n7610 & n8117;
  assign n8119 = n33235 & n8115;
  assign n8120 = ~n7975 & n8118;
  assign n8121 = n33235 & ~n8115;
  assign n8122 = ~n33235 & n8115;
  assign n8123 = ~n8121 & ~n8122;
  assign n8124 = ~n8116 & ~n33301;
  assign n8125 = ~n33300 & n33302;
  assign n8126 = ~n8110 & ~n8125;
  assign n8127 = ~n3788 & ~n8126;
  assign n8128 = n3788 & ~n8110;
  assign n8129 = ~n8125 & n8128;
  assign n8130 = ~n7623 & ~n33237;
  assign n8131 = ~n7623 & ~n7975;
  assign n8132 = ~n33237 & n8131;
  assign n8133 = ~n7975 & n8130;
  assign n8134 = n7631 & ~n33303;
  assign n8135 = n7635 & n8131;
  assign n8136 = n7631 & ~n33237;
  assign n8137 = ~n7623 & n8136;
  assign n8138 = ~n7975 & n8137;
  assign n8139 = ~n7631 & ~n33303;
  assign n8140 = ~n8138 & ~n8139;
  assign n8141 = ~n8134 & ~n8135;
  assign n8142 = ~n8129 & ~n33304;
  assign n8143 = ~n8127 & ~n8142;
  assign n8144 = ~n3473 & ~n8143;
  assign n8145 = n3473 & ~n8127;
  assign n8146 = ~n8142 & n8145;
  assign n8147 = n3473 & n8143;
  assign n8148 = ~n7637 & ~n7639;
  assign n8149 = ~n7975 & n8148;
  assign n8150 = n33239 & ~n8149;
  assign n8151 = ~n7637 & ~n33239;
  assign n8152 = ~n7639 & n8151;
  assign n8153 = ~n33239 & n8149;
  assign n8154 = ~n7975 & n8152;
  assign n8155 = n33239 & n8149;
  assign n8156 = ~n33239 & ~n8149;
  assign n8157 = ~n8155 & ~n8156;
  assign n8158 = ~n8150 & ~n33306;
  assign n8159 = ~n33305 & n33307;
  assign n8160 = ~n8144 & ~n8159;
  assign n8161 = ~n3140 & ~n8160;
  assign n8162 = n3140 & ~n8144;
  assign n8163 = ~n8159 & n8162;
  assign n8164 = ~n7653 & ~n33241;
  assign n8165 = ~n7653 & ~n7975;
  assign n8166 = ~n33241 & n8165;
  assign n8167 = ~n7975 & n8164;
  assign n8168 = n7661 & ~n33308;
  assign n8169 = n7665 & n8165;
  assign n8170 = n7661 & ~n33241;
  assign n8171 = ~n7653 & n8170;
  assign n8172 = ~n7975 & n8171;
  assign n8173 = ~n7661 & ~n33308;
  assign n8174 = ~n8172 & ~n8173;
  assign n8175 = ~n8168 & ~n8169;
  assign n8176 = ~n8163 & ~n33309;
  assign n8177 = ~n8161 & ~n8176;
  assign n8178 = ~n2855 & ~n8177;
  assign n8179 = n2855 & ~n8161;
  assign n8180 = ~n8176 & n8179;
  assign n8181 = n2855 & n8177;
  assign n8182 = ~n7667 & ~n7669;
  assign n8183 = ~n7667 & ~n7975;
  assign n8184 = ~n7669 & n8183;
  assign n8185 = ~n7975 & n8182;
  assign n8186 = ~n33243 & ~n33311;
  assign n8187 = n7681 & n8183;
  assign n8188 = n33243 & n33311;
  assign n8189 = ~n7667 & ~n33243;
  assign n8190 = ~n7669 & n8189;
  assign n8191 = ~n7975 & n8190;
  assign n8192 = n33243 & ~n33311;
  assign n8193 = ~n8191 & ~n8192;
  assign n8194 = ~n8186 & ~n33312;
  assign n8195 = ~n33310 & ~n33313;
  assign n8196 = ~n8178 & ~n8195;
  assign n8197 = ~n2556 & ~n8196;
  assign n8198 = n2556 & ~n8178;
  assign n8199 = ~n8195 & n8198;
  assign n8200 = ~n7683 & ~n33245;
  assign n8201 = ~n7683 & ~n7975;
  assign n8202 = ~n33245 & n8201;
  assign n8203 = ~n7975 & n8200;
  assign n8204 = n7691 & ~n33314;
  assign n8205 = n7695 & n8201;
  assign n8206 = n7691 & ~n33245;
  assign n8207 = ~n7683 & n8206;
  assign n8208 = ~n7975 & n8207;
  assign n8209 = ~n7691 & ~n33314;
  assign n8210 = ~n8208 & ~n8209;
  assign n8211 = ~n8204 & ~n8205;
  assign n8212 = ~n8199 & ~n33315;
  assign n8213 = ~n8197 & ~n8212;
  assign n8214 = ~n2301 & ~n8213;
  assign n8215 = n2301 & ~n8197;
  assign n8216 = ~n8212 & n8215;
  assign n8217 = n2301 & n8213;
  assign n8218 = ~n7697 & ~n7699;
  assign n8219 = ~n7975 & n8218;
  assign n8220 = ~n33248 & ~n8219;
  assign n8221 = ~n7697 & n33248;
  assign n8222 = ~n7699 & n8221;
  assign n8223 = n33248 & n8219;
  assign n8224 = ~n7975 & n8222;
  assign n8225 = ~n8220 & ~n33317;
  assign n8226 = ~n33316 & ~n8225;
  assign n8227 = ~n8214 & ~n8226;
  assign n8228 = ~n2038 & ~n8227;
  assign n8229 = n2038 & ~n8214;
  assign n8230 = ~n8226 & n8229;
  assign n8231 = ~n7715 & ~n33250;
  assign n8232 = ~n7715 & ~n7975;
  assign n8233 = ~n33250 & n8232;
  assign n8234 = ~n7975 & n8231;
  assign n8235 = n7723 & ~n33318;
  assign n8236 = n7727 & n8232;
  assign n8237 = n7723 & ~n33250;
  assign n8238 = ~n7715 & n8237;
  assign n8239 = ~n7975 & n8238;
  assign n8240 = ~n7723 & ~n33318;
  assign n8241 = ~n8239 & ~n8240;
  assign n8242 = ~n8235 & ~n8236;
  assign n8243 = ~n8230 & ~n33319;
  assign n8244 = ~n8228 & ~n8243;
  assign n8245 = ~n1812 & ~n8244;
  assign n8246 = n1812 & ~n8228;
  assign n8247 = ~n8243 & n8246;
  assign n8248 = n1812 & n8244;
  assign n8249 = ~n7729 & ~n7731;
  assign n8250 = ~n7729 & ~n7975;
  assign n8251 = ~n7731 & n8250;
  assign n8252 = ~n7975 & n8249;
  assign n8253 = n7739 & ~n33321;
  assign n8254 = n7740 & n8250;
  assign n8255 = ~n7739 & n33321;
  assign n8256 = ~n7729 & n7739;
  assign n8257 = ~n7731 & n8256;
  assign n8258 = ~n7975 & n8257;
  assign n8259 = ~n7739 & ~n33321;
  assign n8260 = ~n8258 & ~n8259;
  assign n8261 = ~n8253 & ~n33322;
  assign n8262 = ~n33320 & ~n33323;
  assign n8263 = ~n8245 & ~n8262;
  assign n8264 = ~n1582 & ~n8263;
  assign n8265 = n1582 & ~n8245;
  assign n8266 = ~n8262 & n8265;
  assign n8267 = ~n7742 & ~n33253;
  assign n8268 = ~n7742 & ~n7975;
  assign n8269 = ~n33253 & n8268;
  assign n8270 = ~n7975 & n8267;
  assign n8271 = n7750 & ~n33324;
  assign n8272 = n7754 & n8268;
  assign n8273 = n7750 & ~n33253;
  assign n8274 = ~n7742 & n8273;
  assign n8275 = ~n7975 & n8274;
  assign n8276 = ~n7750 & ~n33324;
  assign n8277 = ~n8275 & ~n8276;
  assign n8278 = ~n8271 & ~n8272;
  assign n8279 = ~n8266 & ~n33325;
  assign n8280 = ~n8264 & ~n8279;
  assign n8281 = ~n1388 & ~n8280;
  assign n8282 = n1388 & ~n8264;
  assign n8283 = ~n8279 & n8282;
  assign n8284 = n1388 & n8280;
  assign n8285 = ~n7756 & ~n7758;
  assign n8286 = ~n7975 & n8285;
  assign n8287 = ~n33256 & n8286;
  assign n8288 = n33256 & ~n8286;
  assign n8289 = ~n7756 & n33256;
  assign n8290 = ~n7758 & n8289;
  assign n8291 = n33256 & n8286;
  assign n8292 = ~n7975 & n8290;
  assign n8293 = ~n33256 & ~n8286;
  assign n8294 = ~n33327 & ~n8293;
  assign n8295 = ~n8287 & ~n8288;
  assign n8296 = ~n33326 & ~n33328;
  assign n8297 = ~n8281 & ~n8296;
  assign n8298 = ~n1192 & ~n8297;
  assign n8299 = n1192 & ~n8281;
  assign n8300 = ~n8296 & n8299;
  assign n8301 = ~n7774 & ~n33258;
  assign n8302 = ~n7774 & ~n7975;
  assign n8303 = ~n33258 & n8302;
  assign n8304 = ~n7975 & n8301;
  assign n8305 = n7782 & ~n33329;
  assign n8306 = n7786 & n8302;
  assign n8307 = n7782 & ~n33258;
  assign n8308 = ~n7774 & n8307;
  assign n8309 = ~n7975 & n8308;
  assign n8310 = ~n7782 & ~n33329;
  assign n8311 = ~n8309 & ~n8310;
  assign n8312 = ~n8305 & ~n8306;
  assign n8313 = ~n8300 & ~n33330;
  assign n8314 = ~n8298 & ~n8313;
  assign n8315 = ~n1028 & ~n8314;
  assign n8316 = n1028 & ~n8298;
  assign n8317 = ~n8313 & n8316;
  assign n8318 = n1028 & n8314;
  assign n8319 = ~n7788 & ~n7790;
  assign n8320 = ~n7788 & ~n7975;
  assign n8321 = ~n7790 & n8320;
  assign n8322 = ~n7975 & n8319;
  assign n8323 = n33260 & ~n33332;
  assign n8324 = n7802 & n8320;
  assign n8325 = ~n33260 & n33332;
  assign n8326 = ~n7788 & n33260;
  assign n8327 = ~n7790 & n8326;
  assign n8328 = ~n7975 & n8327;
  assign n8329 = ~n33260 & ~n33332;
  assign n8330 = ~n8328 & ~n8329;
  assign n8331 = ~n8323 & ~n33333;
  assign n8332 = ~n33331 & ~n33334;
  assign n8333 = ~n8315 & ~n8332;
  assign n8334 = ~n866 & ~n8333;
  assign n8335 = n866 & ~n8315;
  assign n8336 = ~n8332 & n8335;
  assign n8337 = ~n7804 & ~n33262;
  assign n8338 = ~n7804 & ~n7975;
  assign n8339 = ~n33262 & n8338;
  assign n8340 = ~n7975 & n8337;
  assign n8341 = n7812 & ~n33335;
  assign n8342 = n7816 & n8338;
  assign n8343 = n7812 & ~n33262;
  assign n8344 = ~n7804 & n8343;
  assign n8345 = ~n7975 & n8344;
  assign n8346 = ~n7812 & ~n33335;
  assign n8347 = ~n8345 & ~n8346;
  assign n8348 = ~n8341 & ~n8342;
  assign n8349 = ~n8336 & ~n33336;
  assign n8350 = ~n8334 & ~n8349;
  assign n8351 = ~n730 & ~n8350;
  assign n8352 = ~n7818 & ~n7820;
  assign n8353 = ~n7975 & n8352;
  assign n8354 = ~n33265 & ~n8353;
  assign n8355 = ~n7818 & n33265;
  assign n8356 = ~n7820 & n8355;
  assign n8357 = n33265 & n8353;
  assign n8358 = ~n7975 & n8356;
  assign n8359 = ~n8354 & ~n33337;
  assign n8360 = n730 & ~n8334;
  assign n8361 = ~n8349 & n8360;
  assign n8362 = n730 & n8350;
  assign n8363 = ~n8359 & ~n33338;
  assign n8364 = ~n8351 & ~n8363;
  assign n8365 = ~n602 & ~n8364;
  assign n8366 = n602 & ~n8351;
  assign n8367 = ~n8363 & n8366;
  assign n8368 = ~n7836 & ~n33267;
  assign n8369 = ~n7836 & ~n7975;
  assign n8370 = ~n33267 & n8369;
  assign n8371 = ~n7975 & n8368;
  assign n8372 = n7844 & ~n33339;
  assign n8373 = n7848 & n8369;
  assign n8374 = n7844 & ~n33267;
  assign n8375 = ~n7836 & n8374;
  assign n8376 = ~n7975 & n8375;
  assign n8377 = ~n7844 & ~n33339;
  assign n8378 = ~n8376 & ~n8377;
  assign n8379 = ~n8372 & ~n8373;
  assign n8380 = ~n8367 & ~n33340;
  assign n8381 = ~n8365 & ~n8380;
  assign n8382 = ~n497 & ~n8381;
  assign n8383 = n497 & ~n8365;
  assign n8384 = ~n8380 & n8383;
  assign n8385 = n497 & n8381;
  assign n8386 = ~n7850 & ~n7860;
  assign n8387 = ~n7850 & ~n7975;
  assign n8388 = ~n7860 & n8387;
  assign n8389 = ~n7975 & n8386;
  assign n8390 = n7858 & ~n33342;
  assign n8391 = n7861 & n8387;
  assign n8392 = ~n7850 & n7858;
  assign n8393 = ~n7860 & n8392;
  assign n8394 = ~n7975 & n8393;
  assign n8395 = ~n7858 & ~n33342;
  assign n8396 = ~n8394 & ~n8395;
  assign n8397 = ~n8390 & ~n8391;
  assign n8398 = ~n33341 & ~n33343;
  assign n8399 = ~n8382 & ~n8398;
  assign n8400 = ~n403 & ~n8399;
  assign n8401 = n403 & ~n8382;
  assign n8402 = ~n8398 & n8401;
  assign n8403 = ~n7863 & ~n33270;
  assign n8404 = ~n7863 & ~n7975;
  assign n8405 = ~n33270 & n8404;
  assign n8406 = ~n7975 & n8403;
  assign n8407 = n7871 & ~n33344;
  assign n8408 = n7875 & n8404;
  assign n8409 = n7871 & ~n33270;
  assign n8410 = ~n7863 & n8409;
  assign n8411 = ~n7975 & n8410;
  assign n8412 = ~n7871 & ~n33344;
  assign n8413 = ~n8411 & ~n8412;
  assign n8414 = ~n8407 & ~n8408;
  assign n8415 = ~n8402 & ~n33345;
  assign n8416 = ~n8400 & ~n8415;
  assign n8417 = ~n330 & ~n8416;
  assign n8418 = ~n7877 & ~n7879;
  assign n8419 = ~n7975 & n8418;
  assign n8420 = ~n33272 & ~n8419;
  assign n8421 = ~n7877 & n33272;
  assign n8422 = ~n7879 & n8421;
  assign n8423 = n33272 & n8419;
  assign n8424 = ~n7975 & n8422;
  assign n8425 = ~n8420 & ~n33346;
  assign n8426 = n330 & ~n8400;
  assign n8427 = ~n8415 & n8426;
  assign n8428 = n330 & n8416;
  assign n8429 = ~n8425 & ~n33347;
  assign n8430 = ~n8417 & ~n8429;
  assign n8431 = ~n271 & ~n8430;
  assign n8432 = n271 & ~n8417;
  assign n8433 = ~n8429 & n8432;
  assign n8434 = ~n7894 & ~n33274;
  assign n8435 = ~n7894 & ~n7975;
  assign n8436 = ~n33274 & n8435;
  assign n8437 = ~n7975 & n8434;
  assign n8438 = n7902 & ~n33348;
  assign n8439 = n7906 & n8435;
  assign n8440 = n7902 & ~n33274;
  assign n8441 = ~n7894 & n8440;
  assign n8442 = ~n7975 & n8441;
  assign n8443 = ~n7902 & ~n33348;
  assign n8444 = ~n8442 & ~n8443;
  assign n8445 = ~n8438 & ~n8439;
  assign n8446 = ~n8433 & ~n33349;
  assign n8447 = ~n8431 & ~n8446;
  assign n8448 = ~n217 & ~n8447;
  assign n8449 = n217 & ~n8431;
  assign n8450 = ~n8446 & n8449;
  assign n8451 = n217 & n8447;
  assign n8452 = ~n7908 & ~n7918;
  assign n8453 = ~n7908 & ~n7975;
  assign n8454 = ~n7918 & n8453;
  assign n8455 = ~n7975 & n8452;
  assign n8456 = n7916 & ~n33351;
  assign n8457 = n7919 & n8453;
  assign n8458 = ~n7908 & n7916;
  assign n8459 = ~n7918 & n8458;
  assign n8460 = ~n7975 & n8459;
  assign n8461 = ~n7916 & ~n33351;
  assign n8462 = ~n8460 & ~n8461;
  assign n8463 = ~n8456 & ~n8457;
  assign n8464 = ~n33350 & ~n33352;
  assign n8465 = ~n8448 & ~n8464;
  assign n8466 = ~n198 & ~n8465;
  assign n8467 = n198 & ~n8448;
  assign n8468 = ~n8464 & n8467;
  assign n8469 = ~n7921 & ~n33277;
  assign n8470 = ~n7921 & ~n7975;
  assign n8471 = ~n33277 & n8470;
  assign n8472 = ~n7975 & n8469;
  assign n8473 = n7929 & ~n33353;
  assign n8474 = n7933 & n8470;
  assign n8475 = n7929 & ~n33277;
  assign n8476 = ~n7921 & n8475;
  assign n8477 = ~n7975 & n8476;
  assign n8478 = ~n7929 & ~n33353;
  assign n8479 = ~n8477 & ~n8478;
  assign n8480 = ~n8473 & ~n8474;
  assign n8481 = ~n8468 & ~n33354;
  assign n8482 = ~n8466 & ~n8481;
  assign n8483 = ~n7935 & ~n7937;
  assign n8484 = ~n7975 & n8483;
  assign n8485 = ~n33279 & ~n8484;
  assign n8486 = ~n7935 & n33279;
  assign n8487 = ~n7937 & n8486;
  assign n8488 = n33279 & n8484;
  assign n8489 = ~n7975 & n8487;
  assign n8490 = ~n8485 & ~n33355;
  assign n8491 = ~n7951 & ~n7959;
  assign n8492 = ~n7959 & ~n7975;
  assign n8493 = ~n7951 & n8492;
  assign n8494 = ~n7975 & n8491;
  assign n8495 = ~n33282 & ~n33356;
  assign n8496 = ~n8490 & n8495;
  assign n8497 = ~n8482 & n8496;
  assign n8498 = n193 & ~n8497;
  assign n8499 = ~n8466 & n8490;
  assign n8500 = ~n8481 & n8499;
  assign n8501 = n8482 & n8490;
  assign n8502 = n7951 & ~n8492;
  assign n8503 = ~n193 & ~n8491;
  assign n8504 = ~n8502 & n8503;
  assign n8505 = ~n33357 & ~n8504;
  assign n8506 = ~n8498 & n8505;
  assign n8507 = ~pi62  & ~n8506;
  assign n8508 = ~pi63  & n8507;
  assign n8509 = n194 & ~n8506;
  assign n8510 = ~n7975 & ~n8504;
  assign n8511 = ~n33357 & n8510;
  assign n8512 = ~n8498 & n8511;
  assign n8513 = ~n33358 & ~n8512;
  assign n8514 = pi64  & ~n8513;
  assign n8515 = ~pi64  & ~n8512;
  assign n8516 = ~pi64  & n8513;
  assign n8517 = ~n33358 & n8515;
  assign n8518 = ~n8514 & ~n33359;
  assign n8519 = pi62  & ~n8506;
  assign n8520 = ~pi60  & ~pi61 ;
  assign n8521 = ~pi62  & n8520;
  assign n8522 = ~n8519 & ~n8521;
  assign n8523 = ~n7975 & ~n8522;
  assign n8524 = ~n33220 & ~n33284;
  assign n8525 = ~n7491 & n8524;
  assign n8526 = ~n7510 & n8525;
  assign n8527 = ~n33222 & n8526;
  assign n8528 = n7496 & n7512;
  assign n8529 = ~n7504 & n8527;
  assign n8530 = ~n8521 & ~n33360;
  assign n8531 = ~n7973 & n8530;
  assign n8532 = ~n33282 & n8531;
  assign n8533 = ~n7967 & n8532;
  assign n8534 = n7975 & n8522;
  assign n8535 = ~n8519 & n8533;
  assign n8536 = pi63  & ~n8507;
  assign n8537 = ~n33358 & ~n8536;
  assign n8538 = ~n33361 & n8537;
  assign n8539 = ~n8523 & ~n8538;
  assign n8540 = ~n7512 & ~n8539;
  assign n8541 = n7512 & ~n8523;
  assign n8542 = n7512 & n8539;
  assign n8543 = ~n8538 & n8541;
  assign n8544 = ~n8518 & ~n33362;
  assign n8545 = ~n8540 & ~n8544;
  assign n8546 = ~n7015 & ~n8545;
  assign n8547 = n7015 & ~n8540;
  assign n8548 = ~n8544 & n8547;
  assign n8549 = ~n7979 & ~n33285;
  assign n8550 = ~n8506 & n8549;
  assign n8551 = n7984 & ~n8550;
  assign n8552 = ~n7984 & ~n33285;
  assign n8553 = ~n7979 & n8552;
  assign n8554 = ~n7984 & n8549;
  assign n8555 = ~n7984 & n8550;
  assign n8556 = ~n8506 & n33363;
  assign n8557 = ~n8551 & ~n33364;
  assign n8558 = ~n8548 & ~n8557;
  assign n8559 = ~n8546 & ~n8558;
  assign n8560 = ~n6579 & ~n8559;
  assign n8561 = ~n7999 & ~n8001;
  assign n8562 = ~n8506 & n8561;
  assign n8563 = ~n8010 & ~n8562;
  assign n8564 = ~n8001 & n8010;
  assign n8565 = ~n7999 & n8564;
  assign n8566 = n8010 & n8562;
  assign n8567 = ~n8506 & n8565;
  assign n8568 = ~n8563 & ~n33365;
  assign n8569 = n6579 & ~n8546;
  assign n8570 = n6579 & n8559;
  assign n8571 = ~n8558 & n8569;
  assign n8572 = ~n8568 & ~n33366;
  assign n8573 = ~n8560 & ~n8572;
  assign n8574 = ~n6117 & ~n8573;
  assign n8575 = n6117 & ~n8560;
  assign n8576 = ~n8572 & n8575;
  assign n8577 = ~n8013 & ~n33287;
  assign n8578 = ~n8506 & n8577;
  assign n8579 = n8023 & ~n8578;
  assign n8580 = ~n8023 & n8578;
  assign n8581 = ~n8013 & n8023;
  assign n8582 = ~n33287 & n8581;
  assign n8583 = n8023 & n8578;
  assign n8584 = ~n8506 & n8582;
  assign n8585 = ~n8023 & ~n8578;
  assign n8586 = ~n33367 & ~n8585;
  assign n8587 = ~n8579 & ~n8580;
  assign n8588 = ~n8576 & ~n33368;
  assign n8589 = ~n8574 & ~n8588;
  assign n8590 = ~n5708 & ~n8589;
  assign n8591 = ~n8026 & ~n8028;
  assign n8592 = ~n8506 & n8591;
  assign n8593 = ~n33290 & ~n8592;
  assign n8594 = ~n8028 & n33290;
  assign n8595 = ~n8026 & n8594;
  assign n8596 = n33290 & n8592;
  assign n8597 = ~n8506 & n8595;
  assign n8598 = ~n8593 & ~n33369;
  assign n8599 = n5708 & ~n8574;
  assign n8600 = n5708 & n8589;
  assign n8601 = ~n8588 & n8599;
  assign n8602 = ~n8598 & ~n33370;
  assign n8603 = ~n8590 & ~n8602;
  assign n8604 = ~n5278 & ~n8603;
  assign n8605 = n5278 & ~n8590;
  assign n8606 = ~n8602 & n8605;
  assign n8607 = ~n8043 & ~n33291;
  assign n8608 = ~n8506 & n8607;
  assign n8609 = ~n33293 & n8608;
  assign n8610 = n33293 & ~n8608;
  assign n8611 = ~n8043 & n33293;
  assign n8612 = ~n33291 & n8611;
  assign n8613 = ~n8506 & n8612;
  assign n8614 = ~n33293 & ~n8608;
  assign n8615 = ~n8613 & ~n8614;
  assign n8616 = ~n8609 & ~n8610;
  assign n8617 = ~n8606 & ~n33371;
  assign n8618 = ~n8604 & ~n8617;
  assign n8619 = ~n4903 & ~n8618;
  assign n8620 = ~n8060 & ~n8062;
  assign n8621 = ~n8506 & n8620;
  assign n8622 = ~n33295 & ~n8621;
  assign n8623 = ~n8062 & n33295;
  assign n8624 = ~n8060 & n8623;
  assign n8625 = n33295 & n8621;
  assign n8626 = ~n8506 & n8624;
  assign n8627 = ~n8622 & ~n33372;
  assign n8628 = n4903 & ~n8604;
  assign n8629 = n4903 & n8618;
  assign n8630 = ~n8617 & n8628;
  assign n8631 = ~n8627 & ~n33373;
  assign n8632 = ~n8619 & ~n8631;
  assign n8633 = ~n4508 & ~n8632;
  assign n8634 = n4508 & ~n8619;
  assign n8635 = ~n8631 & n8634;
  assign n8636 = ~n8077 & ~n33296;
  assign n8637 = ~n8506 & n8636;
  assign n8638 = ~n33297 & ~n8637;
  assign n8639 = ~n8077 & n33297;
  assign n8640 = ~n33296 & n8639;
  assign n8641 = n33297 & n8637;
  assign n8642 = ~n8506 & n8640;
  assign n8643 = n33297 & ~n8637;
  assign n8644 = ~n33297 & n8637;
  assign n8645 = ~n8643 & ~n8644;
  assign n8646 = ~n8638 & ~n33374;
  assign n8647 = ~n8635 & n33375;
  assign n8648 = ~n8633 & ~n8647;
  assign n8649 = ~n4155 & ~n8648;
  assign n8650 = ~n8093 & ~n8095;
  assign n8651 = ~n8506 & n8650;
  assign n8652 = ~n33299 & ~n8651;
  assign n8653 = ~n8095 & n33299;
  assign n8654 = ~n8093 & n8653;
  assign n8655 = n33299 & n8651;
  assign n8656 = ~n8506 & n8654;
  assign n8657 = ~n8652 & ~n33376;
  assign n8658 = n4155 & ~n8633;
  assign n8659 = n4155 & n8648;
  assign n8660 = ~n8647 & n8658;
  assign n8661 = ~n8657 & ~n33377;
  assign n8662 = ~n8649 & ~n8661;
  assign n8663 = ~n3788 & ~n8662;
  assign n8664 = n3788 & ~n8649;
  assign n8665 = ~n8661 & n8664;
  assign n8666 = ~n8110 & ~n33300;
  assign n8667 = ~n8506 & n8666;
  assign n8668 = n33302 & ~n8667;
  assign n8669 = ~n8110 & ~n33302;
  assign n8670 = ~n33300 & n8669;
  assign n8671 = ~n33302 & n8667;
  assign n8672 = ~n8506 & n8670;
  assign n8673 = n33302 & n8667;
  assign n8674 = ~n33302 & ~n8667;
  assign n8675 = ~n8673 & ~n8674;
  assign n8676 = ~n8668 & ~n33378;
  assign n8677 = ~n8665 & n33379;
  assign n8678 = ~n8663 & ~n8677;
  assign n8679 = ~n3473 & ~n8678;
  assign n8680 = ~n8127 & ~n8129;
  assign n8681 = ~n8506 & n8680;
  assign n8682 = ~n33304 & ~n8681;
  assign n8683 = ~n8129 & n33304;
  assign n8684 = ~n8127 & n8683;
  assign n8685 = n33304 & n8681;
  assign n8686 = ~n8506 & n8684;
  assign n8687 = ~n8682 & ~n33380;
  assign n8688 = n3473 & ~n8663;
  assign n8689 = n3473 & n8678;
  assign n8690 = ~n8677 & n8688;
  assign n8691 = ~n8687 & ~n33381;
  assign n8692 = ~n8679 & ~n8691;
  assign n8693 = ~n3140 & ~n8692;
  assign n8694 = n3140 & ~n8679;
  assign n8695 = ~n8691 & n8694;
  assign n8696 = ~n8144 & ~n33305;
  assign n8697 = ~n8144 & ~n8506;
  assign n8698 = ~n33305 & n8697;
  assign n8699 = ~n8506 & n8696;
  assign n8700 = ~n33307 & ~n33382;
  assign n8701 = n8159 & n8697;
  assign n8702 = n33307 & n33382;
  assign n8703 = ~n8144 & ~n33307;
  assign n8704 = ~n33305 & n8703;
  assign n8705 = ~n8506 & n8704;
  assign n8706 = n33307 & ~n33382;
  assign n8707 = ~n8705 & ~n8706;
  assign n8708 = ~n8700 & ~n33383;
  assign n8709 = ~n8695 & ~n33384;
  assign n8710 = ~n8693 & ~n8709;
  assign n8711 = ~n2855 & ~n8710;
  assign n8712 = ~n8161 & ~n8163;
  assign n8713 = ~n8506 & n8712;
  assign n8714 = ~n33309 & ~n8713;
  assign n8715 = ~n8163 & n33309;
  assign n8716 = ~n8161 & n8715;
  assign n8717 = n33309 & n8713;
  assign n8718 = ~n8506 & n8716;
  assign n8719 = ~n8714 & ~n33385;
  assign n8720 = n2855 & ~n8693;
  assign n8721 = n2855 & n8710;
  assign n8722 = ~n8709 & n8720;
  assign n8723 = ~n8719 & ~n33386;
  assign n8724 = ~n8711 & ~n8723;
  assign n8725 = ~n2556 & ~n8724;
  assign n8726 = n2556 & ~n8711;
  assign n8727 = ~n8723 & n8726;
  assign n8728 = ~n8178 & ~n33310;
  assign n8729 = ~n8506 & n8728;
  assign n8730 = ~n33313 & ~n8729;
  assign n8731 = ~n8178 & n33313;
  assign n8732 = ~n33310 & n8731;
  assign n8733 = n33313 & n8729;
  assign n8734 = ~n8506 & n8732;
  assign n8735 = ~n8730 & ~n33387;
  assign n8736 = ~n8727 & ~n8735;
  assign n8737 = ~n8725 & ~n8736;
  assign n8738 = ~n2301 & ~n8737;
  assign n8739 = ~n8197 & ~n8199;
  assign n8740 = ~n8506 & n8739;
  assign n8741 = ~n33315 & ~n8740;
  assign n8742 = ~n8199 & n33315;
  assign n8743 = ~n8197 & n8742;
  assign n8744 = n33315 & n8740;
  assign n8745 = ~n8506 & n8743;
  assign n8746 = ~n8741 & ~n33388;
  assign n8747 = n2301 & ~n8725;
  assign n8748 = n2301 & n8737;
  assign n8749 = ~n8736 & n8747;
  assign n8750 = ~n8746 & ~n33389;
  assign n8751 = ~n8738 & ~n8750;
  assign n8752 = ~n2038 & ~n8751;
  assign n8753 = n2038 & ~n8738;
  assign n8754 = ~n8750 & n8753;
  assign n8755 = ~n8214 & ~n33316;
  assign n8756 = ~n8214 & ~n8506;
  assign n8757 = ~n33316 & n8756;
  assign n8758 = ~n8506 & n8755;
  assign n8759 = n8225 & ~n33390;
  assign n8760 = n8226 & n8756;
  assign n8761 = ~n8225 & n33390;
  assign n8762 = ~n8214 & n8225;
  assign n8763 = ~n33316 & n8762;
  assign n8764 = ~n8506 & n8763;
  assign n8765 = ~n8225 & ~n33390;
  assign n8766 = ~n8764 & ~n8765;
  assign n8767 = ~n8759 & ~n33391;
  assign n8768 = ~n8754 & ~n33392;
  assign n8769 = ~n8752 & ~n8768;
  assign n8770 = ~n1812 & ~n8769;
  assign n8771 = ~n8228 & ~n8230;
  assign n8772 = ~n8506 & n8771;
  assign n8773 = ~n33319 & ~n8772;
  assign n8774 = ~n8230 & n33319;
  assign n8775 = ~n8228 & n8774;
  assign n8776 = n33319 & n8772;
  assign n8777 = ~n8506 & n8775;
  assign n8778 = ~n8773 & ~n33393;
  assign n8779 = n1812 & ~n8752;
  assign n8780 = n1812 & n8769;
  assign n8781 = ~n8768 & n8779;
  assign n8782 = ~n8778 & ~n33394;
  assign n8783 = ~n8770 & ~n8782;
  assign n8784 = ~n1582 & ~n8783;
  assign n8785 = n1582 & ~n8770;
  assign n8786 = ~n8782 & n8785;
  assign n8787 = ~n8245 & ~n33320;
  assign n8788 = ~n8506 & n8787;
  assign n8789 = ~n33323 & n8788;
  assign n8790 = n33323 & ~n8788;
  assign n8791 = ~n8245 & n33323;
  assign n8792 = ~n33320 & n8791;
  assign n8793 = n33323 & n8788;
  assign n8794 = ~n8506 & n8792;
  assign n8795 = ~n33323 & ~n8788;
  assign n8796 = ~n33395 & ~n8795;
  assign n8797 = ~n8789 & ~n8790;
  assign n8798 = ~n8786 & ~n33396;
  assign n8799 = ~n8784 & ~n8798;
  assign n8800 = ~n1388 & ~n8799;
  assign n8801 = ~n8264 & ~n8266;
  assign n8802 = ~n8506 & n8801;
  assign n8803 = ~n33325 & ~n8802;
  assign n8804 = ~n8266 & n33325;
  assign n8805 = ~n8264 & n8804;
  assign n8806 = n33325 & n8802;
  assign n8807 = ~n8506 & n8805;
  assign n8808 = ~n8803 & ~n33397;
  assign n8809 = n1388 & ~n8784;
  assign n8810 = n1388 & n8799;
  assign n8811 = ~n8798 & n8809;
  assign n8812 = ~n8808 & ~n33398;
  assign n8813 = ~n8800 & ~n8812;
  assign n8814 = ~n1192 & ~n8813;
  assign n8815 = n1192 & ~n8800;
  assign n8816 = ~n8812 & n8815;
  assign n8817 = ~n8281 & ~n33326;
  assign n8818 = ~n8281 & ~n8506;
  assign n8819 = ~n33326 & n8818;
  assign n8820 = ~n8506 & n8817;
  assign n8821 = n33328 & ~n33399;
  assign n8822 = n8296 & n8818;
  assign n8823 = ~n33328 & n33399;
  assign n8824 = ~n8281 & n33328;
  assign n8825 = ~n33326 & n8824;
  assign n8826 = ~n8506 & n8825;
  assign n8827 = ~n33328 & ~n33399;
  assign n8828 = ~n8826 & ~n8827;
  assign n8829 = ~n8821 & ~n33400;
  assign n8830 = ~n8816 & ~n33401;
  assign n8831 = ~n8814 & ~n8830;
  assign n8832 = ~n1028 & ~n8831;
  assign n8833 = ~n8298 & ~n8300;
  assign n8834 = ~n8506 & n8833;
  assign n8835 = ~n33330 & ~n8834;
  assign n8836 = ~n8300 & n33330;
  assign n8837 = ~n8298 & n8836;
  assign n8838 = n33330 & n8834;
  assign n8839 = ~n8506 & n8837;
  assign n8840 = ~n8835 & ~n33402;
  assign n8841 = n1028 & ~n8814;
  assign n8842 = n1028 & n8831;
  assign n8843 = ~n8830 & n8841;
  assign n8844 = ~n8840 & ~n33403;
  assign n8845 = ~n8832 & ~n8844;
  assign n8846 = ~n866 & ~n8845;
  assign n8847 = ~n8315 & ~n33331;
  assign n8848 = ~n8506 & n8847;
  assign n8849 = ~n33334 & ~n8848;
  assign n8850 = ~n8315 & n33334;
  assign n8851 = ~n33331 & n8850;
  assign n8852 = n33334 & n8848;
  assign n8853 = ~n8506 & n8851;
  assign n8854 = ~n8849 & ~n33404;
  assign n8855 = n866 & ~n8832;
  assign n8856 = ~n8844 & n8855;
  assign n8857 = ~n8854 & ~n8856;
  assign n8858 = ~n8846 & ~n8857;
  assign n8859 = ~n730 & ~n8858;
  assign n8860 = ~n8334 & ~n8336;
  assign n8861 = ~n8506 & n8860;
  assign n8862 = ~n33336 & ~n8861;
  assign n8863 = ~n8336 & n33336;
  assign n8864 = ~n8334 & n8863;
  assign n8865 = n33336 & n8861;
  assign n8866 = ~n8506 & n8864;
  assign n8867 = ~n8862 & ~n33405;
  assign n8868 = n730 & ~n8846;
  assign n8869 = n730 & n8858;
  assign n8870 = ~n8857 & n8868;
  assign n8871 = ~n8867 & ~n33406;
  assign n8872 = ~n8859 & ~n8871;
  assign n8873 = ~n602 & ~n8872;
  assign n8874 = n602 & ~n8859;
  assign n8875 = ~n8871 & n8874;
  assign n8876 = ~n8351 & ~n33338;
  assign n8877 = ~n8351 & ~n8506;
  assign n8878 = ~n33338 & n8877;
  assign n8879 = ~n8506 & n8876;
  assign n8880 = n8359 & ~n33407;
  assign n8881 = n8363 & n8877;
  assign n8882 = ~n8351 & n8359;
  assign n8883 = ~n33338 & n8882;
  assign n8884 = ~n8506 & n8883;
  assign n8885 = ~n8359 & ~n33407;
  assign n8886 = ~n8884 & ~n8885;
  assign n8887 = ~n8880 & ~n8881;
  assign n8888 = ~n8875 & ~n33408;
  assign n8889 = ~n8873 & ~n8888;
  assign n8890 = ~n497 & ~n8889;
  assign n8891 = ~n8365 & ~n8367;
  assign n8892 = ~n8506 & n8891;
  assign n8893 = ~n33340 & ~n8892;
  assign n8894 = ~n8367 & n33340;
  assign n8895 = ~n8365 & n8894;
  assign n8896 = n33340 & n8892;
  assign n8897 = ~n8506 & n8895;
  assign n8898 = ~n8893 & ~n33409;
  assign n8899 = n497 & ~n8873;
  assign n8900 = n497 & n8889;
  assign n8901 = ~n8888 & n8899;
  assign n8902 = ~n8898 & ~n33410;
  assign n8903 = ~n8890 & ~n8902;
  assign n8904 = ~n403 & ~n8903;
  assign n8905 = ~n8382 & ~n33341;
  assign n8906 = ~n8506 & n8905;
  assign n8907 = ~n33343 & ~n8906;
  assign n8908 = ~n8382 & n33343;
  assign n8909 = ~n33341 & n8908;
  assign n8910 = n33343 & n8906;
  assign n8911 = ~n8506 & n8909;
  assign n8912 = ~n8907 & ~n33411;
  assign n8913 = n403 & ~n8890;
  assign n8914 = ~n8902 & n8913;
  assign n8915 = ~n8912 & ~n8914;
  assign n8916 = ~n8904 & ~n8915;
  assign n8917 = ~n330 & ~n8916;
  assign n8918 = ~n8400 & ~n8402;
  assign n8919 = ~n8506 & n8918;
  assign n8920 = ~n33345 & ~n8919;
  assign n8921 = ~n8402 & n33345;
  assign n8922 = ~n8400 & n8921;
  assign n8923 = n33345 & n8919;
  assign n8924 = ~n8506 & n8922;
  assign n8925 = ~n8920 & ~n33412;
  assign n8926 = n330 & ~n8904;
  assign n8927 = n330 & n8916;
  assign n8928 = ~n8915 & n8926;
  assign n8929 = ~n8925 & ~n33413;
  assign n8930 = ~n8917 & ~n8929;
  assign n8931 = ~n271 & ~n8930;
  assign n8932 = n271 & ~n8917;
  assign n8933 = ~n8929 & n8932;
  assign n8934 = ~n8417 & ~n33347;
  assign n8935 = ~n8417 & ~n8506;
  assign n8936 = ~n33347 & n8935;
  assign n8937 = ~n8506 & n8934;
  assign n8938 = n8425 & ~n33414;
  assign n8939 = n8429 & n8935;
  assign n8940 = ~n8417 & n8425;
  assign n8941 = ~n33347 & n8940;
  assign n8942 = ~n8506 & n8941;
  assign n8943 = ~n8425 & ~n33414;
  assign n8944 = ~n8942 & ~n8943;
  assign n8945 = ~n8938 & ~n8939;
  assign n8946 = ~n8933 & ~n33415;
  assign n8947 = ~n8931 & ~n8946;
  assign n8948 = ~n217 & ~n8947;
  assign n8949 = ~n8431 & ~n8433;
  assign n8950 = ~n8506 & n8949;
  assign n8951 = ~n33349 & ~n8950;
  assign n8952 = ~n8433 & n33349;
  assign n8953 = ~n8431 & n8952;
  assign n8954 = n33349 & n8950;
  assign n8955 = ~n8506 & n8953;
  assign n8956 = ~n8951 & ~n33416;
  assign n8957 = n217 & ~n8931;
  assign n8958 = n217 & n8947;
  assign n8959 = ~n8946 & n8957;
  assign n8960 = ~n8956 & ~n33417;
  assign n8961 = ~n8948 & ~n8960;
  assign n8962 = ~n198 & ~n8961;
  assign n8963 = ~n8448 & ~n33350;
  assign n8964 = ~n8506 & n8963;
  assign n8965 = ~n33352 & ~n8964;
  assign n8966 = ~n8448 & n33352;
  assign n8967 = ~n33350 & n8966;
  assign n8968 = n33352 & n8964;
  assign n8969 = ~n8506 & n8967;
  assign n8970 = ~n8965 & ~n33418;
  assign n8971 = n198 & ~n8948;
  assign n8972 = ~n8960 & n8971;
  assign n8973 = ~n8970 & ~n8972;
  assign n8974 = ~n8962 & ~n8973;
  assign n8975 = ~n8466 & ~n8468;
  assign n8976 = ~n8506 & n8975;
  assign n8977 = ~n33354 & ~n8976;
  assign n8978 = ~n8468 & n33354;
  assign n8979 = ~n8466 & n8978;
  assign n8980 = n33354 & n8976;
  assign n8981 = ~n8506 & n8979;
  assign n8982 = ~n8977 & ~n33419;
  assign n8983 = ~n8482 & ~n8490;
  assign n8984 = ~n8490 & ~n8506;
  assign n8985 = ~n8482 & n8984;
  assign n8986 = ~n8506 & n8983;
  assign n8987 = ~n33357 & ~n33420;
  assign n8988 = ~n8982 & n8987;
  assign n8989 = ~n8974 & n8988;
  assign n8990 = n193 & ~n8989;
  assign n8991 = ~n8962 & n8982;
  assign n8992 = n8974 & n8982;
  assign n8993 = ~n8973 & n8991;
  assign n8994 = n8482 & ~n8984;
  assign n8995 = ~n193 & ~n8983;
  assign n8996 = ~n8994 & n8995;
  assign n8997 = ~n33421 & ~n8996;
  assign n8998 = ~n8990 & n8997;
  assign n8999 = ~n8540 & ~n33362;
  assign n9000 = ~n8540 & ~n8998;
  assign n9001 = ~n33362 & n9000;
  assign n9002 = ~n8998 & n8999;
  assign n9003 = n8518 & ~n33422;
  assign n9004 = n8544 & n9000;
  assign n9005 = n8518 & ~n33362;
  assign n9006 = ~n8540 & n9005;
  assign n9007 = ~n8998 & n9006;
  assign n9008 = ~n8518 & ~n33422;
  assign n9009 = ~n9007 & ~n9008;
  assign n9010 = ~n9003 & ~n9004;
  assign n9011 = pi60  & ~n8998;
  assign n9012 = ~pi58  & ~pi59 ;
  assign n9013 = ~pi60  & n9012;
  assign n9014 = ~n9011 & ~n9013;
  assign n9015 = ~n8506 & ~n9014;
  assign n9016 = ~pi60  & ~n8998;
  assign n9017 = pi61  & ~n9016;
  assign n9018 = ~pi61  & n9016;
  assign n9019 = n8520 & ~n8998;
  assign n9020 = ~n9017 & ~n33424;
  assign n9021 = ~n33280 & ~n33360;
  assign n9022 = ~n7954 & n9021;
  assign n9023 = ~n7973 & n9022;
  assign n9024 = ~n33282 & n9023;
  assign n9025 = n7959 & n7975;
  assign n9026 = ~n7967 & n9024;
  assign n9027 = ~n9013 & ~n33425;
  assign n9028 = ~n8504 & n9027;
  assign n9029 = ~n33357 & n9028;
  assign n9030 = ~n8498 & n9029;
  assign n9031 = n8506 & n9014;
  assign n9032 = ~n9011 & n9030;
  assign n9033 = n9020 & ~n33426;
  assign n9034 = ~n9015 & ~n9033;
  assign n9035 = ~n7975 & ~n9034;
  assign n9036 = n7975 & ~n9015;
  assign n9037 = ~n9033 & n9036;
  assign n9038 = ~n8506 & ~n8996;
  assign n9039 = ~n33421 & n9038;
  assign n9040 = ~n8990 & n9039;
  assign n9041 = ~n33424 & ~n9040;
  assign n9042 = pi62  & ~n9041;
  assign n9043 = ~pi62  & ~n9040;
  assign n9044 = ~pi62  & n9041;
  assign n9045 = ~n33424 & n9043;
  assign n9046 = ~n9042 & ~n33427;
  assign n9047 = ~n9037 & ~n9046;
  assign n9048 = ~n9035 & ~n9047;
  assign n9049 = ~n7512 & ~n9048;
  assign n9050 = n7512 & ~n9035;
  assign n9051 = ~n9047 & n9050;
  assign n9052 = n7512 & n9048;
  assign n9053 = ~n8523 & ~n33361;
  assign n9054 = ~n8998 & n9053;
  assign n9055 = n8537 & ~n9054;
  assign n9056 = ~n8537 & n9053;
  assign n9057 = ~n8537 & n9054;
  assign n9058 = ~n8998 & n9056;
  assign n9059 = ~n9055 & ~n33429;
  assign n9060 = ~n33428 & ~n9059;
  assign n9061 = ~n9049 & ~n9060;
  assign n9062 = ~n7015 & ~n9061;
  assign n9063 = n7015 & ~n9049;
  assign n9064 = ~n9060 & n9063;
  assign n9065 = ~n33423 & ~n9064;
  assign n9066 = ~n9062 & ~n9065;
  assign n9067 = ~n6579 & ~n9066;
  assign n9068 = n6579 & ~n9062;
  assign n9069 = ~n9065 & n9068;
  assign n9070 = n6579 & n9066;
  assign n9071 = ~n8546 & ~n8548;
  assign n9072 = ~n8998 & n9071;
  assign n9073 = n8557 & ~n9072;
  assign n9074 = ~n8557 & n9072;
  assign n9075 = ~n8546 & n8557;
  assign n9076 = ~n8548 & n9075;
  assign n9077 = n8557 & n9072;
  assign n9078 = ~n8998 & n9076;
  assign n9079 = ~n8557 & ~n9072;
  assign n9080 = ~n33431 & ~n9079;
  assign n9081 = ~n9073 & ~n9074;
  assign n9082 = ~n33430 & ~n33432;
  assign n9083 = ~n9067 & ~n9082;
  assign n9084 = ~n6117 & ~n9083;
  assign n9085 = n6117 & ~n9067;
  assign n9086 = ~n9082 & n9085;
  assign n9087 = ~n8560 & ~n33366;
  assign n9088 = ~n8560 & ~n8998;
  assign n9089 = ~n33366 & n9088;
  assign n9090 = ~n8998 & n9087;
  assign n9091 = n8568 & ~n33433;
  assign n9092 = n8572 & n9088;
  assign n9093 = n8568 & ~n33366;
  assign n9094 = ~n8560 & n9093;
  assign n9095 = ~n8998 & n9094;
  assign n9096 = ~n8568 & ~n33433;
  assign n9097 = ~n9095 & ~n9096;
  assign n9098 = ~n9091 & ~n9092;
  assign n9099 = ~n9086 & ~n33434;
  assign n9100 = ~n9084 & ~n9099;
  assign n9101 = ~n5708 & ~n9100;
  assign n9102 = n5708 & ~n9084;
  assign n9103 = ~n9099 & n9102;
  assign n9104 = n5708 & n9100;
  assign n9105 = ~n8574 & ~n8576;
  assign n9106 = ~n8998 & n9105;
  assign n9107 = ~n33368 & n9106;
  assign n9108 = n33368 & ~n9106;
  assign n9109 = ~n8574 & n33368;
  assign n9110 = ~n8576 & n9109;
  assign n9111 = ~n8998 & n9110;
  assign n9112 = ~n33368 & ~n9106;
  assign n9113 = ~n9111 & ~n9112;
  assign n9114 = ~n9107 & ~n9108;
  assign n9115 = ~n33435 & ~n33436;
  assign n9116 = ~n9101 & ~n9115;
  assign n9117 = ~n5278 & ~n9116;
  assign n9118 = n5278 & ~n9101;
  assign n9119 = ~n9115 & n9118;
  assign n9120 = ~n8590 & ~n33370;
  assign n9121 = ~n8590 & ~n8998;
  assign n9122 = ~n33370 & n9121;
  assign n9123 = ~n8998 & n9120;
  assign n9124 = n8598 & ~n33437;
  assign n9125 = n8602 & n9121;
  assign n9126 = n8598 & ~n33370;
  assign n9127 = ~n8590 & n9126;
  assign n9128 = ~n8998 & n9127;
  assign n9129 = ~n8598 & ~n33437;
  assign n9130 = ~n9128 & ~n9129;
  assign n9131 = ~n9124 & ~n9125;
  assign n9132 = ~n9119 & ~n33438;
  assign n9133 = ~n9117 & ~n9132;
  assign n9134 = ~n4903 & ~n9133;
  assign n9135 = n4903 & ~n9117;
  assign n9136 = ~n9132 & n9135;
  assign n9137 = n4903 & n9133;
  assign n9138 = ~n8604 & ~n8606;
  assign n9139 = ~n8998 & n9138;
  assign n9140 = ~n33371 & ~n9139;
  assign n9141 = ~n8604 & n33371;
  assign n9142 = ~n8606 & n9141;
  assign n9143 = n33371 & n9139;
  assign n9144 = ~n8998 & n9142;
  assign n9145 = n33371 & ~n9139;
  assign n9146 = ~n33371 & n9139;
  assign n9147 = ~n9145 & ~n9146;
  assign n9148 = ~n9140 & ~n33440;
  assign n9149 = ~n33439 & n33441;
  assign n9150 = ~n9134 & ~n9149;
  assign n9151 = ~n4508 & ~n9150;
  assign n9152 = n4508 & ~n9134;
  assign n9153 = ~n9149 & n9152;
  assign n9154 = ~n8619 & ~n33373;
  assign n9155 = ~n8619 & ~n8998;
  assign n9156 = ~n33373 & n9155;
  assign n9157 = ~n8998 & n9154;
  assign n9158 = n8627 & ~n33442;
  assign n9159 = n8631 & n9155;
  assign n9160 = n8627 & ~n33373;
  assign n9161 = ~n8619 & n9160;
  assign n9162 = ~n8998 & n9161;
  assign n9163 = ~n8627 & ~n33442;
  assign n9164 = ~n9162 & ~n9163;
  assign n9165 = ~n9158 & ~n9159;
  assign n9166 = ~n9153 & ~n33443;
  assign n9167 = ~n9151 & ~n9166;
  assign n9168 = ~n4155 & ~n9167;
  assign n9169 = n4155 & ~n9151;
  assign n9170 = ~n9166 & n9169;
  assign n9171 = n4155 & n9167;
  assign n9172 = ~n8633 & ~n8635;
  assign n9173 = ~n8998 & n9172;
  assign n9174 = n33375 & ~n9173;
  assign n9175 = ~n8633 & ~n33375;
  assign n9176 = ~n8635 & n9175;
  assign n9177 = ~n33375 & n9173;
  assign n9178 = ~n8998 & n9176;
  assign n9179 = n33375 & n9173;
  assign n9180 = ~n33375 & ~n9173;
  assign n9181 = ~n9179 & ~n9180;
  assign n9182 = ~n9174 & ~n33445;
  assign n9183 = ~n33444 & n33446;
  assign n9184 = ~n9168 & ~n9183;
  assign n9185 = ~n3788 & ~n9184;
  assign n9186 = n3788 & ~n9168;
  assign n9187 = ~n9183 & n9186;
  assign n9188 = ~n8649 & ~n33377;
  assign n9189 = ~n8649 & ~n8998;
  assign n9190 = ~n33377 & n9189;
  assign n9191 = ~n8998 & n9188;
  assign n9192 = n8657 & ~n33447;
  assign n9193 = n8661 & n9189;
  assign n9194 = n8657 & ~n33377;
  assign n9195 = ~n8649 & n9194;
  assign n9196 = ~n8998 & n9195;
  assign n9197 = ~n8657 & ~n33447;
  assign n9198 = ~n9196 & ~n9197;
  assign n9199 = ~n9192 & ~n9193;
  assign n9200 = ~n9187 & ~n33448;
  assign n9201 = ~n9185 & ~n9200;
  assign n9202 = ~n3473 & ~n9201;
  assign n9203 = n3473 & ~n9185;
  assign n9204 = ~n9200 & n9203;
  assign n9205 = n3473 & n9201;
  assign n9206 = ~n8663 & ~n8665;
  assign n9207 = ~n8663 & ~n8998;
  assign n9208 = ~n8665 & n9207;
  assign n9209 = ~n8998 & n9206;
  assign n9210 = ~n33379 & ~n33450;
  assign n9211 = n8677 & n9207;
  assign n9212 = n33379 & n33450;
  assign n9213 = ~n8663 & ~n33379;
  assign n9214 = ~n8665 & n9213;
  assign n9215 = ~n8998 & n9214;
  assign n9216 = n33379 & ~n33450;
  assign n9217 = ~n9215 & ~n9216;
  assign n9218 = ~n9210 & ~n33451;
  assign n9219 = ~n33449 & ~n33452;
  assign n9220 = ~n9202 & ~n9219;
  assign n9221 = ~n3140 & ~n9220;
  assign n9222 = n3140 & ~n9202;
  assign n9223 = ~n9219 & n9222;
  assign n9224 = ~n8679 & ~n33381;
  assign n9225 = ~n8679 & ~n8998;
  assign n9226 = ~n33381 & n9225;
  assign n9227 = ~n8998 & n9224;
  assign n9228 = n8687 & ~n33453;
  assign n9229 = n8691 & n9225;
  assign n9230 = n8687 & ~n33381;
  assign n9231 = ~n8679 & n9230;
  assign n9232 = ~n8998 & n9231;
  assign n9233 = ~n8687 & ~n33453;
  assign n9234 = ~n9232 & ~n9233;
  assign n9235 = ~n9228 & ~n9229;
  assign n9236 = ~n9223 & ~n33454;
  assign n9237 = ~n9221 & ~n9236;
  assign n9238 = ~n2855 & ~n9237;
  assign n9239 = n2855 & ~n9221;
  assign n9240 = ~n9236 & n9239;
  assign n9241 = n2855 & n9237;
  assign n9242 = ~n8693 & ~n8695;
  assign n9243 = ~n8998 & n9242;
  assign n9244 = ~n33384 & ~n9243;
  assign n9245 = ~n8693 & n33384;
  assign n9246 = ~n8695 & n9245;
  assign n9247 = n33384 & n9243;
  assign n9248 = ~n8998 & n9246;
  assign n9249 = ~n9244 & ~n33456;
  assign n9250 = ~n33455 & ~n9249;
  assign n9251 = ~n9238 & ~n9250;
  assign n9252 = ~n2556 & ~n9251;
  assign n9253 = n2556 & ~n9238;
  assign n9254 = ~n9250 & n9253;
  assign n9255 = ~n8711 & ~n33386;
  assign n9256 = ~n8711 & ~n8998;
  assign n9257 = ~n33386 & n9256;
  assign n9258 = ~n8998 & n9255;
  assign n9259 = n8719 & ~n33457;
  assign n9260 = n8723 & n9256;
  assign n9261 = n8719 & ~n33386;
  assign n9262 = ~n8711 & n9261;
  assign n9263 = ~n8998 & n9262;
  assign n9264 = ~n8719 & ~n33457;
  assign n9265 = ~n9263 & ~n9264;
  assign n9266 = ~n9259 & ~n9260;
  assign n9267 = ~n9254 & ~n33458;
  assign n9268 = ~n9252 & ~n9267;
  assign n9269 = ~n2301 & ~n9268;
  assign n9270 = n2301 & ~n9252;
  assign n9271 = ~n9267 & n9270;
  assign n9272 = n2301 & n9268;
  assign n9273 = ~n8725 & ~n8727;
  assign n9274 = ~n8725 & ~n8998;
  assign n9275 = ~n8727 & n9274;
  assign n9276 = ~n8998 & n9273;
  assign n9277 = n8735 & ~n33460;
  assign n9278 = n8736 & n9274;
  assign n9279 = ~n8735 & n33460;
  assign n9280 = ~n8725 & n8735;
  assign n9281 = ~n8727 & n9280;
  assign n9282 = ~n8998 & n9281;
  assign n9283 = ~n8735 & ~n33460;
  assign n9284 = ~n9282 & ~n9283;
  assign n9285 = ~n9277 & ~n33461;
  assign n9286 = ~n33459 & ~n33462;
  assign n9287 = ~n9269 & ~n9286;
  assign n9288 = ~n2038 & ~n9287;
  assign n9289 = n2038 & ~n9269;
  assign n9290 = ~n9286 & n9289;
  assign n9291 = ~n8738 & ~n33389;
  assign n9292 = ~n8738 & ~n8998;
  assign n9293 = ~n33389 & n9292;
  assign n9294 = ~n8998 & n9291;
  assign n9295 = n8746 & ~n33463;
  assign n9296 = n8750 & n9292;
  assign n9297 = n8746 & ~n33389;
  assign n9298 = ~n8738 & n9297;
  assign n9299 = ~n8998 & n9298;
  assign n9300 = ~n8746 & ~n33463;
  assign n9301 = ~n9299 & ~n9300;
  assign n9302 = ~n9295 & ~n9296;
  assign n9303 = ~n9290 & ~n33464;
  assign n9304 = ~n9288 & ~n9303;
  assign n9305 = ~n1812 & ~n9304;
  assign n9306 = n1812 & ~n9288;
  assign n9307 = ~n9303 & n9306;
  assign n9308 = n1812 & n9304;
  assign n9309 = ~n8752 & ~n8754;
  assign n9310 = ~n8998 & n9309;
  assign n9311 = ~n33392 & n9310;
  assign n9312 = n33392 & ~n9310;
  assign n9313 = ~n8752 & n33392;
  assign n9314 = ~n8754 & n9313;
  assign n9315 = n33392 & n9310;
  assign n9316 = ~n8998 & n9314;
  assign n9317 = ~n33392 & ~n9310;
  assign n9318 = ~n33466 & ~n9317;
  assign n9319 = ~n9311 & ~n9312;
  assign n9320 = ~n33465 & ~n33467;
  assign n9321 = ~n9305 & ~n9320;
  assign n9322 = ~n1582 & ~n9321;
  assign n9323 = n1582 & ~n9305;
  assign n9324 = ~n9320 & n9323;
  assign n9325 = ~n8770 & ~n33394;
  assign n9326 = ~n8770 & ~n8998;
  assign n9327 = ~n33394 & n9326;
  assign n9328 = ~n8998 & n9325;
  assign n9329 = n8778 & ~n33468;
  assign n9330 = n8782 & n9326;
  assign n9331 = n8778 & ~n33394;
  assign n9332 = ~n8770 & n9331;
  assign n9333 = ~n8998 & n9332;
  assign n9334 = ~n8778 & ~n33468;
  assign n9335 = ~n9333 & ~n9334;
  assign n9336 = ~n9329 & ~n9330;
  assign n9337 = ~n9324 & ~n33469;
  assign n9338 = ~n9322 & ~n9337;
  assign n9339 = ~n1388 & ~n9338;
  assign n9340 = n1388 & ~n9322;
  assign n9341 = ~n9337 & n9340;
  assign n9342 = n1388 & n9338;
  assign n9343 = ~n8784 & ~n8786;
  assign n9344 = ~n8784 & ~n8998;
  assign n9345 = ~n8786 & n9344;
  assign n9346 = ~n8998 & n9343;
  assign n9347 = n33396 & ~n33471;
  assign n9348 = n8798 & n9344;
  assign n9349 = ~n33396 & n33471;
  assign n9350 = ~n8784 & n33396;
  assign n9351 = ~n8786 & n9350;
  assign n9352 = ~n8998 & n9351;
  assign n9353 = ~n33396 & ~n33471;
  assign n9354 = ~n9352 & ~n9353;
  assign n9355 = ~n9347 & ~n33472;
  assign n9356 = ~n33470 & ~n33473;
  assign n9357 = ~n9339 & ~n9356;
  assign n9358 = ~n1192 & ~n9357;
  assign n9359 = n1192 & ~n9339;
  assign n9360 = ~n9356 & n9359;
  assign n9361 = ~n8800 & ~n33398;
  assign n9362 = ~n8800 & ~n8998;
  assign n9363 = ~n33398 & n9362;
  assign n9364 = ~n8998 & n9361;
  assign n9365 = n8808 & ~n33474;
  assign n9366 = n8812 & n9362;
  assign n9367 = n8808 & ~n33398;
  assign n9368 = ~n8800 & n9367;
  assign n9369 = ~n8998 & n9368;
  assign n9370 = ~n8808 & ~n33474;
  assign n9371 = ~n9369 & ~n9370;
  assign n9372 = ~n9365 & ~n9366;
  assign n9373 = ~n9360 & ~n33475;
  assign n9374 = ~n9358 & ~n9373;
  assign n9375 = ~n1028 & ~n9374;
  assign n9376 = ~n8814 & ~n8816;
  assign n9377 = ~n8998 & n9376;
  assign n9378 = ~n33401 & ~n9377;
  assign n9379 = ~n8814 & n33401;
  assign n9380 = ~n8816 & n9379;
  assign n9381 = n33401 & n9377;
  assign n9382 = ~n8998 & n9380;
  assign n9383 = ~n9378 & ~n33476;
  assign n9384 = n1028 & ~n9358;
  assign n9385 = ~n9373 & n9384;
  assign n9386 = n1028 & n9374;
  assign n9387 = ~n9383 & ~n33477;
  assign n9388 = ~n9375 & ~n9387;
  assign n9389 = ~n866 & ~n9388;
  assign n9390 = n866 & ~n9375;
  assign n9391 = ~n9387 & n9390;
  assign n9392 = ~n8832 & ~n33403;
  assign n9393 = ~n8832 & ~n8998;
  assign n9394 = ~n33403 & n9393;
  assign n9395 = ~n8998 & n9392;
  assign n9396 = n8840 & ~n33478;
  assign n9397 = n8844 & n9393;
  assign n9398 = n8840 & ~n33403;
  assign n9399 = ~n8832 & n9398;
  assign n9400 = ~n8998 & n9399;
  assign n9401 = ~n8840 & ~n33478;
  assign n9402 = ~n9400 & ~n9401;
  assign n9403 = ~n9396 & ~n9397;
  assign n9404 = ~n9391 & ~n33479;
  assign n9405 = ~n9389 & ~n9404;
  assign n9406 = ~n730 & ~n9405;
  assign n9407 = n730 & ~n9389;
  assign n9408 = ~n9404 & n9407;
  assign n9409 = n730 & n9405;
  assign n9410 = ~n8846 & ~n8856;
  assign n9411 = ~n8846 & ~n8998;
  assign n9412 = ~n8856 & n9411;
  assign n9413 = ~n8998 & n9410;
  assign n9414 = n8854 & ~n33481;
  assign n9415 = n8857 & n9411;
  assign n9416 = ~n8846 & n8854;
  assign n9417 = ~n8856 & n9416;
  assign n9418 = ~n8998 & n9417;
  assign n9419 = ~n8854 & ~n33481;
  assign n9420 = ~n9418 & ~n9419;
  assign n9421 = ~n9414 & ~n9415;
  assign n9422 = ~n33480 & ~n33482;
  assign n9423 = ~n9406 & ~n9422;
  assign n9424 = ~n602 & ~n9423;
  assign n9425 = n602 & ~n9406;
  assign n9426 = ~n9422 & n9425;
  assign n9427 = ~n8859 & ~n33406;
  assign n9428 = ~n8859 & ~n8998;
  assign n9429 = ~n33406 & n9428;
  assign n9430 = ~n8998 & n9427;
  assign n9431 = n8867 & ~n33483;
  assign n9432 = n8871 & n9428;
  assign n9433 = n8867 & ~n33406;
  assign n9434 = ~n8859 & n9433;
  assign n9435 = ~n8998 & n9434;
  assign n9436 = ~n8867 & ~n33483;
  assign n9437 = ~n9435 & ~n9436;
  assign n9438 = ~n9431 & ~n9432;
  assign n9439 = ~n9426 & ~n33484;
  assign n9440 = ~n9424 & ~n9439;
  assign n9441 = ~n497 & ~n9440;
  assign n9442 = ~n8873 & ~n8875;
  assign n9443 = ~n8998 & n9442;
  assign n9444 = ~n33408 & ~n9443;
  assign n9445 = ~n8873 & n33408;
  assign n9446 = ~n8875 & n9445;
  assign n9447 = n33408 & n9443;
  assign n9448 = ~n8998 & n9446;
  assign n9449 = ~n9444 & ~n33485;
  assign n9450 = n497 & ~n9424;
  assign n9451 = ~n9439 & n9450;
  assign n9452 = n497 & n9440;
  assign n9453 = ~n9449 & ~n33486;
  assign n9454 = ~n9441 & ~n9453;
  assign n9455 = ~n403 & ~n9454;
  assign n9456 = n403 & ~n9441;
  assign n9457 = ~n9453 & n9456;
  assign n9458 = ~n8890 & ~n33410;
  assign n9459 = ~n8890 & ~n8998;
  assign n9460 = ~n33410 & n9459;
  assign n9461 = ~n8998 & n9458;
  assign n9462 = n8898 & ~n33487;
  assign n9463 = n8902 & n9459;
  assign n9464 = n8898 & ~n33410;
  assign n9465 = ~n8890 & n9464;
  assign n9466 = ~n8998 & n9465;
  assign n9467 = ~n8898 & ~n33487;
  assign n9468 = ~n9466 & ~n9467;
  assign n9469 = ~n9462 & ~n9463;
  assign n9470 = ~n9457 & ~n33488;
  assign n9471 = ~n9455 & ~n9470;
  assign n9472 = ~n330 & ~n9471;
  assign n9473 = n330 & ~n9455;
  assign n9474 = ~n9470 & n9473;
  assign n9475 = n330 & n9471;
  assign n9476 = ~n8904 & ~n8914;
  assign n9477 = ~n8904 & ~n8998;
  assign n9478 = ~n8914 & n9477;
  assign n9479 = ~n8998 & n9476;
  assign n9480 = n8912 & ~n33490;
  assign n9481 = n8915 & n9477;
  assign n9482 = ~n8904 & n8912;
  assign n9483 = ~n8914 & n9482;
  assign n9484 = ~n8998 & n9483;
  assign n9485 = ~n8912 & ~n33490;
  assign n9486 = ~n9484 & ~n9485;
  assign n9487 = ~n9480 & ~n9481;
  assign n9488 = ~n33489 & ~n33491;
  assign n9489 = ~n9472 & ~n9488;
  assign n9490 = ~n271 & ~n9489;
  assign n9491 = n271 & ~n9472;
  assign n9492 = ~n9488 & n9491;
  assign n9493 = ~n8917 & ~n33413;
  assign n9494 = ~n8917 & ~n8998;
  assign n9495 = ~n33413 & n9494;
  assign n9496 = ~n8998 & n9493;
  assign n9497 = n8925 & ~n33492;
  assign n9498 = n8929 & n9494;
  assign n9499 = n8925 & ~n33413;
  assign n9500 = ~n8917 & n9499;
  assign n9501 = ~n8998 & n9500;
  assign n9502 = ~n8925 & ~n33492;
  assign n9503 = ~n9501 & ~n9502;
  assign n9504 = ~n9497 & ~n9498;
  assign n9505 = ~n9492 & ~n33493;
  assign n9506 = ~n9490 & ~n9505;
  assign n9507 = ~n217 & ~n9506;
  assign n9508 = ~n8931 & ~n8933;
  assign n9509 = ~n8998 & n9508;
  assign n9510 = ~n33415 & ~n9509;
  assign n9511 = ~n8931 & n33415;
  assign n9512 = ~n8933 & n9511;
  assign n9513 = n33415 & n9509;
  assign n9514 = ~n8998 & n9512;
  assign n9515 = ~n9510 & ~n33494;
  assign n9516 = n217 & ~n9490;
  assign n9517 = ~n9505 & n9516;
  assign n9518 = n217 & n9506;
  assign n9519 = ~n9515 & ~n33495;
  assign n9520 = ~n9507 & ~n9519;
  assign n9521 = ~n198 & ~n9520;
  assign n9522 = n198 & ~n9507;
  assign n9523 = ~n9519 & n9522;
  assign n9524 = ~n8948 & ~n33417;
  assign n9525 = ~n8948 & ~n8998;
  assign n9526 = ~n33417 & n9525;
  assign n9527 = ~n8998 & n9524;
  assign n9528 = n8956 & ~n33496;
  assign n9529 = n8960 & n9525;
  assign n9530 = n8956 & ~n33417;
  assign n9531 = ~n8948 & n9530;
  assign n9532 = ~n8998 & n9531;
  assign n9533 = ~n8956 & ~n33496;
  assign n9534 = ~n9532 & ~n9533;
  assign n9535 = ~n9528 & ~n9529;
  assign n9536 = ~n9523 & ~n33497;
  assign n9537 = ~n9521 & ~n9536;
  assign n9538 = ~n8962 & ~n8972;
  assign n9539 = ~n8962 & ~n8998;
  assign n9540 = ~n8972 & n9539;
  assign n9541 = ~n8998 & n9538;
  assign n9542 = n8970 & ~n33498;
  assign n9543 = n8973 & n9539;
  assign n9544 = ~n8962 & n8970;
  assign n9545 = ~n8972 & n9544;
  assign n9546 = ~n8998 & n9545;
  assign n9547 = ~n8970 & ~n33498;
  assign n9548 = ~n9546 & ~n9547;
  assign n9549 = ~n9542 & ~n9543;
  assign n9550 = ~n8974 & ~n8982;
  assign n9551 = ~n8982 & ~n8998;
  assign n9552 = ~n8974 & n9551;
  assign n9553 = ~n8998 & n9550;
  assign n9554 = ~n33421 & ~n33500;
  assign n9555 = ~n33499 & n9554;
  assign n9556 = ~n9537 & n9555;
  assign n9557 = n193 & ~n9556;
  assign n9558 = ~n9521 & n33499;
  assign n9559 = ~n9536 & n9558;
  assign n9560 = n9537 & n33499;
  assign n9561 = n8974 & ~n9551;
  assign n9562 = ~n193 & ~n9550;
  assign n9563 = ~n9561 & n9562;
  assign n9564 = ~n33501 & ~n9563;
  assign n9565 = ~n9557 & n9564;
  assign n9566 = ~n9062 & ~n9064;
  assign n9567 = ~n9565 & n9566;
  assign n9568 = ~n33423 & ~n9567;
  assign n9569 = n33423 & ~n9064;
  assign n9570 = ~n9062 & n9569;
  assign n9571 = n33423 & n9567;
  assign n9572 = ~n9565 & n9570;
  assign n9573 = ~n9568 & ~n33502;
  assign n9574 = ~n9035 & ~n9037;
  assign n9575 = ~n9565 & n9574;
  assign n9576 = ~n9046 & ~n9575;
  assign n9577 = ~n9037 & n9046;
  assign n9578 = ~n9035 & n9577;
  assign n9579 = n9046 & n9575;
  assign n9580 = ~n9565 & n9578;
  assign n9581 = ~n9576 & ~n33503;
  assign n9582 = ~pi58  & ~n9565;
  assign n9583 = ~pi59  & n9582;
  assign n9584 = n9012 & ~n9565;
  assign n9585 = ~n8998 & ~n9563;
  assign n9586 = ~n33501 & n9585;
  assign n9587 = ~n9557 & n9586;
  assign n9588 = ~n33504 & ~n9587;
  assign n9589 = pi60  & ~n9588;
  assign n9590 = ~pi60  & ~n9587;
  assign n9591 = ~pi60  & n9588;
  assign n9592 = ~n33504 & n9590;
  assign n9593 = ~n9589 & ~n33505;
  assign n9594 = pi58  & ~n9565;
  assign n9595 = ~pi56  & ~pi57 ;
  assign n9596 = ~pi58  & n9595;
  assign n9597 = ~n33355 & ~n33425;
  assign n9598 = ~n8485 & n9597;
  assign n9599 = ~n8504 & n9598;
  assign n9600 = ~n33357 & n9599;
  assign n9601 = n8490 & n8506;
  assign n9602 = ~n8498 & n9600;
  assign n9603 = ~n9596 & ~n33506;
  assign n9604 = ~n8996 & n9603;
  assign n9605 = ~n33421 & n9604;
  assign n9606 = ~n8990 & n9605;
  assign n9607 = ~n9594 & ~n9596;
  assign n9608 = n8998 & n9607;
  assign n9609 = ~n9594 & n9606;
  assign n9610 = pi59  & ~n9582;
  assign n9611 = ~n33504 & ~n9610;
  assign n9612 = ~n33507 & n9611;
  assign n9613 = ~n8998 & ~n9607;
  assign n9614 = n8506 & ~n9613;
  assign n9615 = ~n9612 & ~n9613;
  assign n9616 = n8506 & n9615;
  assign n9617 = ~n9612 & n9614;
  assign n9618 = ~n9593 & ~n33508;
  assign n9619 = ~n8506 & ~n9615;
  assign n9620 = n7975 & ~n9619;
  assign n9621 = ~n9618 & n9620;
  assign n9622 = ~n9015 & ~n33426;
  assign n9623 = ~n9565 & n9622;
  assign n9624 = n9020 & ~n9623;
  assign n9625 = ~n9020 & n9622;
  assign n9626 = ~n9020 & n9623;
  assign n9627 = ~n9565 & n9625;
  assign n9628 = ~n9624 & ~n33509;
  assign n9629 = ~n9621 & ~n9628;
  assign n9630 = ~n9618 & ~n9619;
  assign n9631 = ~n7975 & ~n9630;
  assign n9632 = n7512 & ~n9631;
  assign n9633 = ~n9629 & ~n9631;
  assign n9634 = n7512 & n9633;
  assign n9635 = ~n9629 & n9632;
  assign n9636 = ~n9581 & ~n33510;
  assign n9637 = ~n7512 & ~n9633;
  assign n9638 = ~n9636 & ~n9637;
  assign n9639 = ~n7015 & ~n9638;
  assign n9640 = n7015 & ~n9637;
  assign n9641 = ~n9636 & n9640;
  assign n9642 = ~n9049 & ~n33428;
  assign n9643 = ~n9565 & n9642;
  assign n9644 = n9059 & ~n9643;
  assign n9645 = ~n9059 & n9643;
  assign n9646 = ~n9049 & n9059;
  assign n9647 = ~n33428 & n9646;
  assign n9648 = n9059 & n9643;
  assign n9649 = ~n9565 & n9647;
  assign n9650 = ~n9059 & ~n9643;
  assign n9651 = ~n33511 & ~n9650;
  assign n9652 = ~n9644 & ~n9645;
  assign n9653 = ~n9641 & ~n33512;
  assign n9654 = ~n9639 & ~n9653;
  assign n9655 = ~n6579 & ~n9654;
  assign n9656 = n6579 & ~n9639;
  assign n9657 = n6579 & n9654;
  assign n9658 = ~n9653 & n9656;
  assign n9659 = ~n9573 & ~n33513;
  assign n9660 = ~n9655 & ~n9659;
  assign n9661 = ~n6117 & ~n9660;
  assign n9662 = n6117 & ~n9655;
  assign n9663 = ~n9659 & n9662;
  assign n9664 = ~n9067 & ~n33430;
  assign n9665 = ~n9565 & n9664;
  assign n9666 = ~n33432 & n9665;
  assign n9667 = n33432 & ~n9665;
  assign n9668 = ~n9067 & n33432;
  assign n9669 = ~n33430 & n9668;
  assign n9670 = ~n9565 & n9669;
  assign n9671 = ~n33432 & ~n9665;
  assign n9672 = ~n9670 & ~n9671;
  assign n9673 = ~n9666 & ~n9667;
  assign n9674 = ~n9663 & ~n33514;
  assign n9675 = ~n9661 & ~n9674;
  assign n9676 = ~n5708 & ~n9675;
  assign n9677 = ~n9084 & ~n9086;
  assign n9678 = ~n9565 & n9677;
  assign n9679 = ~n33434 & ~n9678;
  assign n9680 = ~n9086 & n33434;
  assign n9681 = ~n9084 & n9680;
  assign n9682 = n33434 & n9678;
  assign n9683 = ~n9565 & n9681;
  assign n9684 = ~n9679 & ~n33515;
  assign n9685 = n5708 & ~n9661;
  assign n9686 = n5708 & n9675;
  assign n9687 = ~n9674 & n9685;
  assign n9688 = ~n9684 & ~n33516;
  assign n9689 = ~n9676 & ~n9688;
  assign n9690 = ~n5278 & ~n9689;
  assign n9691 = n5278 & ~n9676;
  assign n9692 = ~n9688 & n9691;
  assign n9693 = ~n9101 & ~n33435;
  assign n9694 = ~n9565 & n9693;
  assign n9695 = ~n33436 & ~n9694;
  assign n9696 = ~n9101 & n33436;
  assign n9697 = ~n33435 & n9696;
  assign n9698 = n33436 & n9694;
  assign n9699 = ~n9565 & n9697;
  assign n9700 = n33436 & ~n9694;
  assign n9701 = ~n33436 & n9694;
  assign n9702 = ~n9700 & ~n9701;
  assign n9703 = ~n9695 & ~n33517;
  assign n9704 = ~n9692 & n33518;
  assign n9705 = ~n9690 & ~n9704;
  assign n9706 = ~n4903 & ~n9705;
  assign n9707 = ~n9117 & ~n9119;
  assign n9708 = ~n9565 & n9707;
  assign n9709 = ~n33438 & ~n9708;
  assign n9710 = ~n9119 & n33438;
  assign n9711 = ~n9117 & n9710;
  assign n9712 = n33438 & n9708;
  assign n9713 = ~n9565 & n9711;
  assign n9714 = ~n9709 & ~n33519;
  assign n9715 = n4903 & ~n9690;
  assign n9716 = n4903 & n9705;
  assign n9717 = ~n9704 & n9715;
  assign n9718 = ~n9714 & ~n33520;
  assign n9719 = ~n9706 & ~n9718;
  assign n9720 = ~n4508 & ~n9719;
  assign n9721 = n4508 & ~n9706;
  assign n9722 = ~n9718 & n9721;
  assign n9723 = ~n9134 & ~n33439;
  assign n9724 = ~n9565 & n9723;
  assign n9725 = n33441 & ~n9724;
  assign n9726 = ~n9134 & ~n33441;
  assign n9727 = ~n33439 & n9726;
  assign n9728 = ~n33441 & n9724;
  assign n9729 = ~n9565 & n9727;
  assign n9730 = n33441 & n9724;
  assign n9731 = ~n33441 & ~n9724;
  assign n9732 = ~n9730 & ~n9731;
  assign n9733 = ~n9725 & ~n33521;
  assign n9734 = ~n9722 & n33522;
  assign n9735 = ~n9720 & ~n9734;
  assign n9736 = ~n4155 & ~n9735;
  assign n9737 = ~n9151 & ~n9153;
  assign n9738 = ~n9565 & n9737;
  assign n9739 = ~n33443 & ~n9738;
  assign n9740 = ~n9153 & n33443;
  assign n9741 = ~n9151 & n9740;
  assign n9742 = n33443 & n9738;
  assign n9743 = ~n9565 & n9741;
  assign n9744 = ~n9739 & ~n33523;
  assign n9745 = n4155 & ~n9720;
  assign n9746 = n4155 & n9735;
  assign n9747 = ~n9734 & n9745;
  assign n9748 = ~n9744 & ~n33524;
  assign n9749 = ~n9736 & ~n9748;
  assign n9750 = ~n3788 & ~n9749;
  assign n9751 = n3788 & ~n9736;
  assign n9752 = ~n9748 & n9751;
  assign n9753 = ~n9168 & ~n33444;
  assign n9754 = ~n9168 & ~n9565;
  assign n9755 = ~n33444 & n9754;
  assign n9756 = ~n9565 & n9753;
  assign n9757 = ~n33446 & ~n33525;
  assign n9758 = n9183 & n9754;
  assign n9759 = n33446 & n33525;
  assign n9760 = ~n9168 & ~n33446;
  assign n9761 = ~n33444 & n9760;
  assign n9762 = ~n9565 & n9761;
  assign n9763 = n33446 & ~n33525;
  assign n9764 = ~n9762 & ~n9763;
  assign n9765 = ~n9757 & ~n33526;
  assign n9766 = ~n9752 & ~n33527;
  assign n9767 = ~n9750 & ~n9766;
  assign n9768 = ~n3473 & ~n9767;
  assign n9769 = ~n9185 & ~n9187;
  assign n9770 = ~n9565 & n9769;
  assign n9771 = ~n33448 & ~n9770;
  assign n9772 = ~n9187 & n33448;
  assign n9773 = ~n9185 & n9772;
  assign n9774 = n33448 & n9770;
  assign n9775 = ~n9565 & n9773;
  assign n9776 = ~n9771 & ~n33528;
  assign n9777 = n3473 & ~n9750;
  assign n9778 = n3473 & n9767;
  assign n9779 = ~n9766 & n9777;
  assign n9780 = ~n9776 & ~n33529;
  assign n9781 = ~n9768 & ~n9780;
  assign n9782 = ~n3140 & ~n9781;
  assign n9783 = n3140 & ~n9768;
  assign n9784 = ~n9780 & n9783;
  assign n9785 = ~n9202 & ~n33449;
  assign n9786 = ~n9565 & n9785;
  assign n9787 = ~n33452 & ~n9786;
  assign n9788 = ~n9202 & n33452;
  assign n9789 = ~n33449 & n9788;
  assign n9790 = n33452 & n9786;
  assign n9791 = ~n9565 & n9789;
  assign n9792 = ~n9787 & ~n33530;
  assign n9793 = ~n9784 & ~n9792;
  assign n9794 = ~n9782 & ~n9793;
  assign n9795 = ~n2855 & ~n9794;
  assign n9796 = ~n9221 & ~n9223;
  assign n9797 = ~n9565 & n9796;
  assign n9798 = ~n33454 & ~n9797;
  assign n9799 = ~n9223 & n33454;
  assign n9800 = ~n9221 & n9799;
  assign n9801 = n33454 & n9797;
  assign n9802 = ~n9565 & n9800;
  assign n9803 = ~n9798 & ~n33531;
  assign n9804 = n2855 & ~n9782;
  assign n9805 = n2855 & n9794;
  assign n9806 = ~n9793 & n9804;
  assign n9807 = ~n9803 & ~n33532;
  assign n9808 = ~n9795 & ~n9807;
  assign n9809 = ~n2556 & ~n9808;
  assign n9810 = n2556 & ~n9795;
  assign n9811 = ~n9807 & n9810;
  assign n9812 = ~n9238 & ~n33455;
  assign n9813 = ~n9238 & ~n9565;
  assign n9814 = ~n33455 & n9813;
  assign n9815 = ~n9565 & n9812;
  assign n9816 = n9249 & ~n33533;
  assign n9817 = n9250 & n9813;
  assign n9818 = ~n9249 & n33533;
  assign n9819 = ~n9238 & n9249;
  assign n9820 = ~n33455 & n9819;
  assign n9821 = ~n9565 & n9820;
  assign n9822 = ~n9249 & ~n33533;
  assign n9823 = ~n9821 & ~n9822;
  assign n9824 = ~n9816 & ~n33534;
  assign n9825 = ~n9811 & ~n33535;
  assign n9826 = ~n9809 & ~n9825;
  assign n9827 = ~n2301 & ~n9826;
  assign n9828 = ~n9252 & ~n9254;
  assign n9829 = ~n9565 & n9828;
  assign n9830 = ~n33458 & ~n9829;
  assign n9831 = ~n9254 & n33458;
  assign n9832 = ~n9252 & n9831;
  assign n9833 = n33458 & n9829;
  assign n9834 = ~n9565 & n9832;
  assign n9835 = ~n9830 & ~n33536;
  assign n9836 = n2301 & ~n9809;
  assign n9837 = n2301 & n9826;
  assign n9838 = ~n9825 & n9836;
  assign n9839 = ~n9835 & ~n33537;
  assign n9840 = ~n9827 & ~n9839;
  assign n9841 = ~n2038 & ~n9840;
  assign n9842 = n2038 & ~n9827;
  assign n9843 = ~n9839 & n9842;
  assign n9844 = ~n9269 & ~n33459;
  assign n9845 = ~n9565 & n9844;
  assign n9846 = ~n33462 & n9845;
  assign n9847 = n33462 & ~n9845;
  assign n9848 = ~n9269 & n33462;
  assign n9849 = ~n33459 & n9848;
  assign n9850 = n33462 & n9845;
  assign n9851 = ~n9565 & n9849;
  assign n9852 = ~n33462 & ~n9845;
  assign n9853 = ~n33538 & ~n9852;
  assign n9854 = ~n9846 & ~n9847;
  assign n9855 = ~n9843 & ~n33539;
  assign n9856 = ~n9841 & ~n9855;
  assign n9857 = ~n1812 & ~n9856;
  assign n9858 = ~n9288 & ~n9290;
  assign n9859 = ~n9565 & n9858;
  assign n9860 = ~n33464 & ~n9859;
  assign n9861 = ~n9290 & n33464;
  assign n9862 = ~n9288 & n9861;
  assign n9863 = n33464 & n9859;
  assign n9864 = ~n9565 & n9862;
  assign n9865 = ~n9860 & ~n33540;
  assign n9866 = n1812 & ~n9841;
  assign n9867 = n1812 & n9856;
  assign n9868 = ~n9855 & n9866;
  assign n9869 = ~n9865 & ~n33541;
  assign n9870 = ~n9857 & ~n9869;
  assign n9871 = ~n1582 & ~n9870;
  assign n9872 = n1582 & ~n9857;
  assign n9873 = ~n9869 & n9872;
  assign n9874 = ~n9305 & ~n33465;
  assign n9875 = ~n9305 & ~n9565;
  assign n9876 = ~n33465 & n9875;
  assign n9877 = ~n9565 & n9874;
  assign n9878 = n33467 & ~n33542;
  assign n9879 = n9320 & n9875;
  assign n9880 = ~n33467 & n33542;
  assign n9881 = ~n9305 & n33467;
  assign n9882 = ~n33465 & n9881;
  assign n9883 = ~n9565 & n9882;
  assign n9884 = ~n33467 & ~n33542;
  assign n9885 = ~n9883 & ~n9884;
  assign n9886 = ~n9878 & ~n33543;
  assign n9887 = ~n9873 & ~n33544;
  assign n9888 = ~n9871 & ~n9887;
  assign n9889 = ~n1388 & ~n9888;
  assign n9890 = ~n9322 & ~n9324;
  assign n9891 = ~n9565 & n9890;
  assign n9892 = ~n33469 & ~n9891;
  assign n9893 = ~n9324 & n33469;
  assign n9894 = ~n9322 & n9893;
  assign n9895 = n33469 & n9891;
  assign n9896 = ~n9565 & n9894;
  assign n9897 = ~n9892 & ~n33545;
  assign n9898 = n1388 & ~n9871;
  assign n9899 = n1388 & n9888;
  assign n9900 = ~n9887 & n9898;
  assign n9901 = ~n9897 & ~n33546;
  assign n9902 = ~n9889 & ~n9901;
  assign n9903 = ~n1192 & ~n9902;
  assign n9904 = ~n9339 & ~n33470;
  assign n9905 = ~n9565 & n9904;
  assign n9906 = ~n33473 & ~n9905;
  assign n9907 = ~n9339 & n33473;
  assign n9908 = ~n33470 & n9907;
  assign n9909 = n33473 & n9905;
  assign n9910 = ~n9565 & n9908;
  assign n9911 = ~n9906 & ~n33547;
  assign n9912 = n1192 & ~n9889;
  assign n9913 = ~n9901 & n9912;
  assign n9914 = ~n9911 & ~n9913;
  assign n9915 = ~n9903 & ~n9914;
  assign n9916 = ~n1028 & ~n9915;
  assign n9917 = ~n9358 & ~n9360;
  assign n9918 = ~n9565 & n9917;
  assign n9919 = ~n33475 & ~n9918;
  assign n9920 = ~n9360 & n33475;
  assign n9921 = ~n9358 & n9920;
  assign n9922 = n33475 & n9918;
  assign n9923 = ~n9565 & n9921;
  assign n9924 = ~n9919 & ~n33548;
  assign n9925 = n1028 & ~n9903;
  assign n9926 = n1028 & n9915;
  assign n9927 = ~n9914 & n9925;
  assign n9928 = ~n9924 & ~n33549;
  assign n9929 = ~n9916 & ~n9928;
  assign n9930 = ~n866 & ~n9929;
  assign n9931 = n866 & ~n9916;
  assign n9932 = ~n9928 & n9931;
  assign n9933 = ~n9375 & ~n33477;
  assign n9934 = ~n9375 & ~n9565;
  assign n9935 = ~n33477 & n9934;
  assign n9936 = ~n9565 & n9933;
  assign n9937 = n9383 & ~n33550;
  assign n9938 = n9387 & n9934;
  assign n9939 = ~n9375 & n9383;
  assign n9940 = ~n33477 & n9939;
  assign n9941 = ~n9565 & n9940;
  assign n9942 = ~n9383 & ~n33550;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = ~n9937 & ~n9938;
  assign n9945 = ~n9932 & ~n33551;
  assign n9946 = ~n9930 & ~n9945;
  assign n9947 = ~n730 & ~n9946;
  assign n9948 = ~n9389 & ~n9391;
  assign n9949 = ~n9565 & n9948;
  assign n9950 = ~n33479 & ~n9949;
  assign n9951 = ~n9391 & n33479;
  assign n9952 = ~n9389 & n9951;
  assign n9953 = n33479 & n9949;
  assign n9954 = ~n9565 & n9952;
  assign n9955 = ~n9950 & ~n33552;
  assign n9956 = n730 & ~n9930;
  assign n9957 = n730 & n9946;
  assign n9958 = ~n9945 & n9956;
  assign n9959 = ~n9955 & ~n33553;
  assign n9960 = ~n9947 & ~n9959;
  assign n9961 = ~n602 & ~n9960;
  assign n9962 = ~n9406 & ~n33480;
  assign n9963 = ~n9565 & n9962;
  assign n9964 = ~n33482 & ~n9963;
  assign n9965 = ~n9406 & n33482;
  assign n9966 = ~n33480 & n9965;
  assign n9967 = n33482 & n9963;
  assign n9968 = ~n9565 & n9966;
  assign n9969 = ~n9964 & ~n33554;
  assign n9970 = n602 & ~n9947;
  assign n9971 = ~n9959 & n9970;
  assign n9972 = ~n9969 & ~n9971;
  assign n9973 = ~n9961 & ~n9972;
  assign n9974 = ~n497 & ~n9973;
  assign n9975 = ~n9424 & ~n9426;
  assign n9976 = ~n9565 & n9975;
  assign n9977 = ~n33484 & ~n9976;
  assign n9978 = ~n9426 & n33484;
  assign n9979 = ~n9424 & n9978;
  assign n9980 = n33484 & n9976;
  assign n9981 = ~n9565 & n9979;
  assign n9982 = ~n9977 & ~n33555;
  assign n9983 = n497 & ~n9961;
  assign n9984 = n497 & n9973;
  assign n9985 = ~n9972 & n9983;
  assign n9986 = ~n9982 & ~n33556;
  assign n9987 = ~n9974 & ~n9986;
  assign n9988 = ~n403 & ~n9987;
  assign n9989 = n403 & ~n9974;
  assign n9990 = ~n9986 & n9989;
  assign n9991 = ~n9441 & ~n33486;
  assign n9992 = ~n9441 & ~n9565;
  assign n9993 = ~n33486 & n9992;
  assign n9994 = ~n9565 & n9991;
  assign n9995 = n9449 & ~n33557;
  assign n9996 = n9453 & n9992;
  assign n9997 = ~n9441 & n9449;
  assign n9998 = ~n33486 & n9997;
  assign n9999 = ~n9565 & n9998;
  assign n10000 = ~n9449 & ~n33557;
  assign n10001 = ~n9999 & ~n10000;
  assign n10002 = ~n9995 & ~n9996;
  assign n10003 = ~n9990 & ~n33558;
  assign n10004 = ~n9988 & ~n10003;
  assign n10005 = ~n330 & ~n10004;
  assign n10006 = ~n9455 & ~n9457;
  assign n10007 = ~n9565 & n10006;
  assign n10008 = ~n33488 & ~n10007;
  assign n10009 = ~n9457 & n33488;
  assign n10010 = ~n9455 & n10009;
  assign n10011 = n33488 & n10007;
  assign n10012 = ~n9565 & n10010;
  assign n10013 = ~n10008 & ~n33559;
  assign n10014 = n330 & ~n9988;
  assign n10015 = n330 & n10004;
  assign n10016 = ~n10003 & n10014;
  assign n10017 = ~n10013 & ~n33560;
  assign n10018 = ~n10005 & ~n10017;
  assign n10019 = ~n271 & ~n10018;
  assign n10020 = ~n9472 & ~n33489;
  assign n10021 = ~n9565 & n10020;
  assign n10022 = ~n33491 & ~n10021;
  assign n10023 = ~n9472 & n33491;
  assign n10024 = ~n33489 & n10023;
  assign n10025 = n33491 & n10021;
  assign n10026 = ~n9565 & n10024;
  assign n10027 = ~n10022 & ~n33561;
  assign n10028 = n271 & ~n10005;
  assign n10029 = ~n10017 & n10028;
  assign n10030 = ~n10027 & ~n10029;
  assign n10031 = ~n10019 & ~n10030;
  assign n10032 = ~n217 & ~n10031;
  assign n10033 = ~n9490 & ~n9492;
  assign n10034 = ~n9565 & n10033;
  assign n10035 = ~n33493 & ~n10034;
  assign n10036 = ~n9492 & n33493;
  assign n10037 = ~n9490 & n10036;
  assign n10038 = n33493 & n10034;
  assign n10039 = ~n9565 & n10037;
  assign n10040 = ~n10035 & ~n33562;
  assign n10041 = n217 & ~n10019;
  assign n10042 = n217 & n10031;
  assign n10043 = ~n10030 & n10041;
  assign n10044 = ~n10040 & ~n33563;
  assign n10045 = ~n10032 & ~n10044;
  assign n10046 = ~n198 & ~n10045;
  assign n10047 = n198 & ~n10032;
  assign n10048 = ~n10044 & n10047;
  assign n10049 = ~n9507 & ~n33495;
  assign n10050 = ~n9507 & ~n9565;
  assign n10051 = ~n33495 & n10050;
  assign n10052 = ~n9565 & n10049;
  assign n10053 = n9515 & ~n33564;
  assign n10054 = n9519 & n10050;
  assign n10055 = ~n9507 & n9515;
  assign n10056 = ~n33495 & n10055;
  assign n10057 = ~n9565 & n10056;
  assign n10058 = ~n9515 & ~n33564;
  assign n10059 = ~n10057 & ~n10058;
  assign n10060 = ~n10053 & ~n10054;
  assign n10061 = ~n10048 & ~n33565;
  assign n10062 = ~n10046 & ~n10061;
  assign n10063 = ~n9521 & ~n9523;
  assign n10064 = ~n9565 & n10063;
  assign n10065 = ~n33497 & ~n10064;
  assign n10066 = ~n9523 & n33497;
  assign n10067 = ~n9521 & n10066;
  assign n10068 = n33497 & n10064;
  assign n10069 = ~n9565 & n10067;
  assign n10070 = ~n10065 & ~n33566;
  assign n10071 = ~n9537 & ~n33499;
  assign n10072 = ~n33499 & ~n9565;
  assign n10073 = ~n9537 & n10072;
  assign n10074 = ~n9565 & n10071;
  assign n10075 = ~n33501 & ~n33567;
  assign n10076 = ~n10070 & n10075;
  assign n10077 = ~n10062 & n10076;
  assign n10078 = n193 & ~n10077;
  assign n10079 = ~n10046 & n10070;
  assign n10080 = n10062 & n10070;
  assign n10081 = ~n10061 & n10079;
  assign n10082 = n9537 & ~n10072;
  assign n10083 = ~n193 & ~n10071;
  assign n10084 = ~n10082 & n10083;
  assign n10085 = ~n33568 & ~n10084;
  assign n10086 = ~n10078 & n10085;
  assign n10087 = ~n9655 & ~n33513;
  assign n10088 = ~n9655 & ~n10086;
  assign n10089 = ~n33513 & n10088;
  assign n10090 = ~n10086 & n10087;
  assign n10091 = n9573 & ~n33569;
  assign n10092 = n9659 & n10088;
  assign n10093 = n9573 & ~n33513;
  assign n10094 = ~n9655 & n10093;
  assign n10095 = ~n10086 & n10094;
  assign n10096 = ~n9573 & ~n33569;
  assign n10097 = ~n10095 & ~n10096;
  assign n10098 = ~n10091 & ~n10092;
  assign n10099 = pi56  & ~n10086;
  assign n10100 = ~pi54  & ~pi55 ;
  assign n10101 = ~pi56  & n10100;
  assign n10102 = ~n10099 & ~n10101;
  assign n10103 = ~n9565 & ~n10102;
  assign n10104 = ~pi56  & ~n10086;
  assign n10105 = pi57  & ~n10104;
  assign n10106 = ~pi57  & n10104;
  assign n10107 = n9595 & ~n10086;
  assign n10108 = ~n10105 & ~n33571;
  assign n10109 = ~n33419 & ~n33506;
  assign n10110 = ~n8977 & n10109;
  assign n10111 = ~n8996 & n10110;
  assign n10112 = ~n33421 & n10111;
  assign n10113 = n8982 & n8998;
  assign n10114 = ~n8990 & n10112;
  assign n10115 = ~n10101 & ~n33572;
  assign n10116 = ~n9563 & n10115;
  assign n10117 = ~n33501 & n10116;
  assign n10118 = ~n9557 & n10117;
  assign n10119 = n9565 & n10102;
  assign n10120 = ~n10099 & n10118;
  assign n10121 = n10108 & ~n33573;
  assign n10122 = ~n10103 & ~n10121;
  assign n10123 = ~n8998 & ~n10122;
  assign n10124 = n8998 & ~n10103;
  assign n10125 = ~n10121 & n10124;
  assign n10126 = ~n9565 & ~n10084;
  assign n10127 = ~n33568 & n10126;
  assign n10128 = ~n10078 & n10127;
  assign n10129 = ~n33571 & ~n10128;
  assign n10130 = pi58  & ~n10129;
  assign n10131 = ~pi58  & ~n10128;
  assign n10132 = ~pi58  & n10129;
  assign n10133 = ~n33571 & n10131;
  assign n10134 = ~n10130 & ~n33574;
  assign n10135 = ~n10125 & ~n10134;
  assign n10136 = ~n10123 & ~n10135;
  assign n10137 = ~n8506 & ~n10136;
  assign n10138 = n8506 & ~n10123;
  assign n10139 = ~n10135 & n10138;
  assign n10140 = n8506 & n10136;
  assign n10141 = ~n33507 & ~n9613;
  assign n10142 = ~n10086 & n10141;
  assign n10143 = n9611 & ~n10142;
  assign n10144 = ~n9611 & n10141;
  assign n10145 = ~n9611 & n10142;
  assign n10146 = ~n10086 & n10144;
  assign n10147 = ~n10143 & ~n33576;
  assign n10148 = ~n33575 & ~n10147;
  assign n10149 = ~n10137 & ~n10148;
  assign n10150 = ~n7975 & ~n10149;
  assign n10151 = n7975 & ~n10137;
  assign n10152 = ~n10148 & n10151;
  assign n10153 = ~n33508 & ~n9619;
  assign n10154 = ~n9619 & ~n10086;
  assign n10155 = ~n33508 & n10154;
  assign n10156 = ~n10086 & n10153;
  assign n10157 = n9593 & ~n33577;
  assign n10158 = n9618 & n10154;
  assign n10159 = n9593 & ~n33508;
  assign n10160 = ~n9619 & n10159;
  assign n10161 = ~n10086 & n10160;
  assign n10162 = ~n9593 & ~n33577;
  assign n10163 = ~n10161 & ~n10162;
  assign n10164 = ~n10157 & ~n10158;
  assign n10165 = ~n10152 & ~n33578;
  assign n10166 = ~n10150 & ~n10165;
  assign n10167 = ~n7512 & ~n10166;
  assign n10168 = n7512 & ~n10150;
  assign n10169 = ~n10165 & n10168;
  assign n10170 = n7512 & n10166;
  assign n10171 = ~n9621 & ~n9631;
  assign n10172 = ~n10086 & n10171;
  assign n10173 = n9628 & ~n10172;
  assign n10174 = ~n9628 & n10172;
  assign n10175 = n9628 & ~n9631;
  assign n10176 = ~n9621 & n10175;
  assign n10177 = n9628 & n10172;
  assign n10178 = ~n10086 & n10176;
  assign n10179 = ~n9628 & ~n10172;
  assign n10180 = ~n33580 & ~n10179;
  assign n10181 = ~n10173 & ~n10174;
  assign n10182 = ~n33579 & ~n33581;
  assign n10183 = ~n10167 & ~n10182;
  assign n10184 = ~n7015 & ~n10183;
  assign n10185 = n7015 & ~n10167;
  assign n10186 = ~n10182 & n10185;
  assign n10187 = n9581 & ~n33510;
  assign n10188 = ~n9637 & n10187;
  assign n10189 = ~n33510 & ~n9637;
  assign n10190 = ~n10086 & n10189;
  assign n10191 = n9581 & n10190;
  assign n10192 = ~n10086 & n10188;
  assign n10193 = ~n9581 & ~n10190;
  assign n10194 = ~n33582 & ~n10193;
  assign n10195 = ~n10186 & ~n10194;
  assign n10196 = ~n10184 & ~n10195;
  assign n10197 = ~n6579 & ~n10196;
  assign n10198 = n6579 & ~n10184;
  assign n10199 = ~n10195 & n10198;
  assign n10200 = n6579 & n10196;
  assign n10201 = ~n9639 & ~n9641;
  assign n10202 = ~n10086 & n10201;
  assign n10203 = ~n33512 & n10202;
  assign n10204 = n33512 & ~n10202;
  assign n10205 = ~n9639 & n33512;
  assign n10206 = ~n9641 & n10205;
  assign n10207 = n33512 & n10202;
  assign n10208 = ~n10086 & n10206;
  assign n10209 = ~n33512 & ~n10202;
  assign n10210 = ~n33584 & ~n10209;
  assign n10211 = ~n10203 & ~n10204;
  assign n10212 = ~n33583 & ~n33585;
  assign n10213 = ~n10197 & ~n10212;
  assign n10214 = ~n6117 & ~n10213;
  assign n10215 = n6117 & ~n10197;
  assign n10216 = ~n10212 & n10215;
  assign n10217 = ~n33570 & ~n10216;
  assign n10218 = ~n10214 & ~n10217;
  assign n10219 = ~n5708 & ~n10218;
  assign n10220 = n5708 & ~n10214;
  assign n10221 = ~n10217 & n10220;
  assign n10222 = n5708 & n10218;
  assign n10223 = ~n9661 & ~n9663;
  assign n10224 = ~n10086 & n10223;
  assign n10225 = ~n33514 & ~n10224;
  assign n10226 = ~n9661 & n33514;
  assign n10227 = ~n9663 & n10226;
  assign n10228 = n33514 & n10224;
  assign n10229 = ~n10086 & n10227;
  assign n10230 = ~n33514 & n10224;
  assign n10231 = n33514 & ~n10224;
  assign n10232 = ~n10230 & ~n10231;
  assign n10233 = ~n10225 & ~n33587;
  assign n10234 = ~n33586 & n33588;
  assign n10235 = ~n10219 & ~n10234;
  assign n10236 = ~n5278 & ~n10235;
  assign n10237 = n5278 & ~n10219;
  assign n10238 = ~n10234 & n10237;
  assign n10239 = ~n9676 & ~n33516;
  assign n10240 = ~n9676 & ~n10086;
  assign n10241 = ~n33516 & n10240;
  assign n10242 = ~n10086 & n10239;
  assign n10243 = n9684 & ~n33589;
  assign n10244 = n9688 & n10240;
  assign n10245 = n9684 & ~n33516;
  assign n10246 = ~n9676 & n10245;
  assign n10247 = ~n10086 & n10246;
  assign n10248 = ~n9684 & ~n33589;
  assign n10249 = ~n10247 & ~n10248;
  assign n10250 = ~n10243 & ~n10244;
  assign n10251 = ~n10238 & ~n33590;
  assign n10252 = ~n10236 & ~n10251;
  assign n10253 = ~n4903 & ~n10252;
  assign n10254 = n4903 & ~n10236;
  assign n10255 = ~n10251 & n10254;
  assign n10256 = n4903 & n10252;
  assign n10257 = ~n9690 & ~n9692;
  assign n10258 = ~n10086 & n10257;
  assign n10259 = n33518 & ~n10258;
  assign n10260 = ~n9690 & ~n33518;
  assign n10261 = ~n9692 & n10260;
  assign n10262 = ~n33518 & n10258;
  assign n10263 = ~n10086 & n10261;
  assign n10264 = n33518 & n10258;
  assign n10265 = ~n33518 & ~n10258;
  assign n10266 = ~n10264 & ~n10265;
  assign n10267 = ~n10259 & ~n33592;
  assign n10268 = ~n33591 & n33593;
  assign n10269 = ~n10253 & ~n10268;
  assign n10270 = ~n4508 & ~n10269;
  assign n10271 = n4508 & ~n10253;
  assign n10272 = ~n10268 & n10271;
  assign n10273 = ~n9706 & ~n33520;
  assign n10274 = ~n9706 & ~n10086;
  assign n10275 = ~n33520 & n10274;
  assign n10276 = ~n10086 & n10273;
  assign n10277 = n9714 & ~n33594;
  assign n10278 = n9718 & n10274;
  assign n10279 = n9714 & ~n33520;
  assign n10280 = ~n9706 & n10279;
  assign n10281 = ~n10086 & n10280;
  assign n10282 = ~n9714 & ~n33594;
  assign n10283 = ~n10281 & ~n10282;
  assign n10284 = ~n10277 & ~n10278;
  assign n10285 = ~n10272 & ~n33595;
  assign n10286 = ~n10270 & ~n10285;
  assign n10287 = ~n4155 & ~n10286;
  assign n10288 = n4155 & ~n10270;
  assign n10289 = ~n10285 & n10288;
  assign n10290 = n4155 & n10286;
  assign n10291 = ~n9720 & ~n9722;
  assign n10292 = ~n9720 & ~n10086;
  assign n10293 = ~n9722 & n10292;
  assign n10294 = ~n10086 & n10291;
  assign n10295 = ~n33522 & ~n33597;
  assign n10296 = n9734 & n10292;
  assign n10297 = n33522 & n33597;
  assign n10298 = ~n9720 & ~n33522;
  assign n10299 = ~n9722 & n10298;
  assign n10300 = ~n10086 & n10299;
  assign n10301 = n33522 & ~n33597;
  assign n10302 = ~n10300 & ~n10301;
  assign n10303 = ~n10295 & ~n33598;
  assign n10304 = ~n33596 & ~n33599;
  assign n10305 = ~n10287 & ~n10304;
  assign n10306 = ~n3788 & ~n10305;
  assign n10307 = n3788 & ~n10287;
  assign n10308 = ~n10304 & n10307;
  assign n10309 = ~n9736 & ~n33524;
  assign n10310 = ~n9736 & ~n10086;
  assign n10311 = ~n33524 & n10310;
  assign n10312 = ~n10086 & n10309;
  assign n10313 = n9744 & ~n33600;
  assign n10314 = n9748 & n10310;
  assign n10315 = n9744 & ~n33524;
  assign n10316 = ~n9736 & n10315;
  assign n10317 = ~n10086 & n10316;
  assign n10318 = ~n9744 & ~n33600;
  assign n10319 = ~n10317 & ~n10318;
  assign n10320 = ~n10313 & ~n10314;
  assign n10321 = ~n10308 & ~n33601;
  assign n10322 = ~n10306 & ~n10321;
  assign n10323 = ~n3473 & ~n10322;
  assign n10324 = n3473 & ~n10306;
  assign n10325 = ~n10321 & n10324;
  assign n10326 = n3473 & n10322;
  assign n10327 = ~n9750 & ~n9752;
  assign n10328 = ~n10086 & n10327;
  assign n10329 = ~n33527 & ~n10328;
  assign n10330 = ~n9750 & n33527;
  assign n10331 = ~n9752 & n10330;
  assign n10332 = n33527 & n10328;
  assign n10333 = ~n10086 & n10331;
  assign n10334 = ~n10329 & ~n33603;
  assign n10335 = ~n33602 & ~n10334;
  assign n10336 = ~n10323 & ~n10335;
  assign n10337 = ~n3140 & ~n10336;
  assign n10338 = n3140 & ~n10323;
  assign n10339 = ~n10335 & n10338;
  assign n10340 = ~n9768 & ~n33529;
  assign n10341 = ~n9768 & ~n10086;
  assign n10342 = ~n33529 & n10341;
  assign n10343 = ~n10086 & n10340;
  assign n10344 = n9776 & ~n33604;
  assign n10345 = n9780 & n10341;
  assign n10346 = n9776 & ~n33529;
  assign n10347 = ~n9768 & n10346;
  assign n10348 = ~n10086 & n10347;
  assign n10349 = ~n9776 & ~n33604;
  assign n10350 = ~n10348 & ~n10349;
  assign n10351 = ~n10344 & ~n10345;
  assign n10352 = ~n10339 & ~n33605;
  assign n10353 = ~n10337 & ~n10352;
  assign n10354 = ~n2855 & ~n10353;
  assign n10355 = n2855 & ~n10337;
  assign n10356 = ~n10352 & n10355;
  assign n10357 = n2855 & n10353;
  assign n10358 = ~n9782 & ~n9784;
  assign n10359 = ~n9782 & ~n10086;
  assign n10360 = ~n9784 & n10359;
  assign n10361 = ~n10086 & n10358;
  assign n10362 = n9792 & ~n33607;
  assign n10363 = n9793 & n10359;
  assign n10364 = ~n9792 & n33607;
  assign n10365 = ~n9782 & n9792;
  assign n10366 = ~n9784 & n10365;
  assign n10367 = ~n10086 & n10366;
  assign n10368 = ~n9792 & ~n33607;
  assign n10369 = ~n10367 & ~n10368;
  assign n10370 = ~n10362 & ~n33608;
  assign n10371 = ~n33606 & ~n33609;
  assign n10372 = ~n10354 & ~n10371;
  assign n10373 = ~n2556 & ~n10372;
  assign n10374 = n2556 & ~n10354;
  assign n10375 = ~n10371 & n10374;
  assign n10376 = ~n9795 & ~n33532;
  assign n10377 = ~n9795 & ~n10086;
  assign n10378 = ~n33532 & n10377;
  assign n10379 = ~n10086 & n10376;
  assign n10380 = n9803 & ~n33610;
  assign n10381 = n9807 & n10377;
  assign n10382 = n9803 & ~n33532;
  assign n10383 = ~n9795 & n10382;
  assign n10384 = ~n10086 & n10383;
  assign n10385 = ~n9803 & ~n33610;
  assign n10386 = ~n10384 & ~n10385;
  assign n10387 = ~n10380 & ~n10381;
  assign n10388 = ~n10375 & ~n33611;
  assign n10389 = ~n10373 & ~n10388;
  assign n10390 = ~n2301 & ~n10389;
  assign n10391 = n2301 & ~n10373;
  assign n10392 = ~n10388 & n10391;
  assign n10393 = n2301 & n10389;
  assign n10394 = ~n9809 & ~n9811;
  assign n10395 = ~n10086 & n10394;
  assign n10396 = ~n33535 & n10395;
  assign n10397 = n33535 & ~n10395;
  assign n10398 = ~n9809 & n33535;
  assign n10399 = ~n9811 & n10398;
  assign n10400 = n33535 & n10395;
  assign n10401 = ~n10086 & n10399;
  assign n10402 = ~n33535 & ~n10395;
  assign n10403 = ~n33613 & ~n10402;
  assign n10404 = ~n10396 & ~n10397;
  assign n10405 = ~n33612 & ~n33614;
  assign n10406 = ~n10390 & ~n10405;
  assign n10407 = ~n2038 & ~n10406;
  assign n10408 = n2038 & ~n10390;
  assign n10409 = ~n10405 & n10408;
  assign n10410 = ~n9827 & ~n33537;
  assign n10411 = ~n9827 & ~n10086;
  assign n10412 = ~n33537 & n10411;
  assign n10413 = ~n10086 & n10410;
  assign n10414 = n9835 & ~n33615;
  assign n10415 = n9839 & n10411;
  assign n10416 = n9835 & ~n33537;
  assign n10417 = ~n9827 & n10416;
  assign n10418 = ~n10086 & n10417;
  assign n10419 = ~n9835 & ~n33615;
  assign n10420 = ~n10418 & ~n10419;
  assign n10421 = ~n10414 & ~n10415;
  assign n10422 = ~n10409 & ~n33616;
  assign n10423 = ~n10407 & ~n10422;
  assign n10424 = ~n1812 & ~n10423;
  assign n10425 = n1812 & ~n10407;
  assign n10426 = ~n10422 & n10425;
  assign n10427 = n1812 & n10423;
  assign n10428 = ~n9841 & ~n9843;
  assign n10429 = ~n9841 & ~n10086;
  assign n10430 = ~n9843 & n10429;
  assign n10431 = ~n10086 & n10428;
  assign n10432 = n33539 & ~n33618;
  assign n10433 = n9855 & n10429;
  assign n10434 = ~n33539 & n33618;
  assign n10435 = ~n9841 & n33539;
  assign n10436 = ~n9843 & n10435;
  assign n10437 = ~n10086 & n10436;
  assign n10438 = ~n33539 & ~n33618;
  assign n10439 = ~n10437 & ~n10438;
  assign n10440 = ~n10432 & ~n33619;
  assign n10441 = ~n33617 & ~n33620;
  assign n10442 = ~n10424 & ~n10441;
  assign n10443 = ~n1582 & ~n10442;
  assign n10444 = n1582 & ~n10424;
  assign n10445 = ~n10441 & n10444;
  assign n10446 = ~n9857 & ~n33541;
  assign n10447 = ~n9857 & ~n10086;
  assign n10448 = ~n33541 & n10447;
  assign n10449 = ~n10086 & n10446;
  assign n10450 = n9865 & ~n33621;
  assign n10451 = n9869 & n10447;
  assign n10452 = n9865 & ~n33541;
  assign n10453 = ~n9857 & n10452;
  assign n10454 = ~n10086 & n10453;
  assign n10455 = ~n9865 & ~n33621;
  assign n10456 = ~n10454 & ~n10455;
  assign n10457 = ~n10450 & ~n10451;
  assign n10458 = ~n10445 & ~n33622;
  assign n10459 = ~n10443 & ~n10458;
  assign n10460 = ~n1388 & ~n10459;
  assign n10461 = ~n9871 & ~n9873;
  assign n10462 = ~n10086 & n10461;
  assign n10463 = ~n33544 & ~n10462;
  assign n10464 = ~n9871 & n33544;
  assign n10465 = ~n9873 & n10464;
  assign n10466 = n33544 & n10462;
  assign n10467 = ~n10086 & n10465;
  assign n10468 = ~n10463 & ~n33623;
  assign n10469 = n1388 & ~n10443;
  assign n10470 = ~n10458 & n10469;
  assign n10471 = n1388 & n10459;
  assign n10472 = ~n10468 & ~n33624;
  assign n10473 = ~n10460 & ~n10472;
  assign n10474 = ~n1192 & ~n10473;
  assign n10475 = n1192 & ~n10460;
  assign n10476 = ~n10472 & n10475;
  assign n10477 = ~n9889 & ~n33546;
  assign n10478 = ~n9889 & ~n10086;
  assign n10479 = ~n33546 & n10478;
  assign n10480 = ~n10086 & n10477;
  assign n10481 = n9897 & ~n33625;
  assign n10482 = n9901 & n10478;
  assign n10483 = n9897 & ~n33546;
  assign n10484 = ~n9889 & n10483;
  assign n10485 = ~n10086 & n10484;
  assign n10486 = ~n9897 & ~n33625;
  assign n10487 = ~n10485 & ~n10486;
  assign n10488 = ~n10481 & ~n10482;
  assign n10489 = ~n10476 & ~n33626;
  assign n10490 = ~n10474 & ~n10489;
  assign n10491 = ~n1028 & ~n10490;
  assign n10492 = n1028 & ~n10474;
  assign n10493 = ~n10489 & n10492;
  assign n10494 = n1028 & n10490;
  assign n10495 = ~n9903 & ~n9913;
  assign n10496 = ~n9903 & ~n10086;
  assign n10497 = ~n9913 & n10496;
  assign n10498 = ~n10086 & n10495;
  assign n10499 = n9911 & ~n33628;
  assign n10500 = n9914 & n10496;
  assign n10501 = ~n9903 & n9911;
  assign n10502 = ~n9913 & n10501;
  assign n10503 = ~n10086 & n10502;
  assign n10504 = ~n9911 & ~n33628;
  assign n10505 = ~n10503 & ~n10504;
  assign n10506 = ~n10499 & ~n10500;
  assign n10507 = ~n33627 & ~n33629;
  assign n10508 = ~n10491 & ~n10507;
  assign n10509 = ~n866 & ~n10508;
  assign n10510 = n866 & ~n10491;
  assign n10511 = ~n10507 & n10510;
  assign n10512 = ~n9916 & ~n33549;
  assign n10513 = ~n9916 & ~n10086;
  assign n10514 = ~n33549 & n10513;
  assign n10515 = ~n10086 & n10512;
  assign n10516 = n9924 & ~n33630;
  assign n10517 = n9928 & n10513;
  assign n10518 = n9924 & ~n33549;
  assign n10519 = ~n9916 & n10518;
  assign n10520 = ~n10086 & n10519;
  assign n10521 = ~n9924 & ~n33630;
  assign n10522 = ~n10520 & ~n10521;
  assign n10523 = ~n10516 & ~n10517;
  assign n10524 = ~n10511 & ~n33631;
  assign n10525 = ~n10509 & ~n10524;
  assign n10526 = ~n730 & ~n10525;
  assign n10527 = ~n9930 & ~n9932;
  assign n10528 = ~n10086 & n10527;
  assign n10529 = ~n33551 & ~n10528;
  assign n10530 = ~n9930 & n33551;
  assign n10531 = ~n9932 & n10530;
  assign n10532 = n33551 & n10528;
  assign n10533 = ~n10086 & n10531;
  assign n10534 = ~n10529 & ~n33632;
  assign n10535 = n730 & ~n10509;
  assign n10536 = ~n10524 & n10535;
  assign n10537 = n730 & n10525;
  assign n10538 = ~n10534 & ~n33633;
  assign n10539 = ~n10526 & ~n10538;
  assign n10540 = ~n602 & ~n10539;
  assign n10541 = n602 & ~n10526;
  assign n10542 = ~n10538 & n10541;
  assign n10543 = ~n9947 & ~n33553;
  assign n10544 = ~n9947 & ~n10086;
  assign n10545 = ~n33553 & n10544;
  assign n10546 = ~n10086 & n10543;
  assign n10547 = n9955 & ~n33634;
  assign n10548 = n9959 & n10544;
  assign n10549 = n9955 & ~n33553;
  assign n10550 = ~n9947 & n10549;
  assign n10551 = ~n10086 & n10550;
  assign n10552 = ~n9955 & ~n33634;
  assign n10553 = ~n10551 & ~n10552;
  assign n10554 = ~n10547 & ~n10548;
  assign n10555 = ~n10542 & ~n33635;
  assign n10556 = ~n10540 & ~n10555;
  assign n10557 = ~n497 & ~n10556;
  assign n10558 = n497 & ~n10540;
  assign n10559 = ~n10555 & n10558;
  assign n10560 = n497 & n10556;
  assign n10561 = ~n9961 & ~n9971;
  assign n10562 = ~n9961 & ~n10086;
  assign n10563 = ~n9971 & n10562;
  assign n10564 = ~n10086 & n10561;
  assign n10565 = n9969 & ~n33637;
  assign n10566 = n9972 & n10562;
  assign n10567 = ~n9961 & n9969;
  assign n10568 = ~n9971 & n10567;
  assign n10569 = ~n10086 & n10568;
  assign n10570 = ~n9969 & ~n33637;
  assign n10571 = ~n10569 & ~n10570;
  assign n10572 = ~n10565 & ~n10566;
  assign n10573 = ~n33636 & ~n33638;
  assign n10574 = ~n10557 & ~n10573;
  assign n10575 = ~n403 & ~n10574;
  assign n10576 = n403 & ~n10557;
  assign n10577 = ~n10573 & n10576;
  assign n10578 = ~n9974 & ~n33556;
  assign n10579 = ~n9974 & ~n10086;
  assign n10580 = ~n33556 & n10579;
  assign n10581 = ~n10086 & n10578;
  assign n10582 = n9982 & ~n33639;
  assign n10583 = n9986 & n10579;
  assign n10584 = n9982 & ~n33556;
  assign n10585 = ~n9974 & n10584;
  assign n10586 = ~n10086 & n10585;
  assign n10587 = ~n9982 & ~n33639;
  assign n10588 = ~n10586 & ~n10587;
  assign n10589 = ~n10582 & ~n10583;
  assign n10590 = ~n10577 & ~n33640;
  assign n10591 = ~n10575 & ~n10590;
  assign n10592 = ~n330 & ~n10591;
  assign n10593 = ~n9988 & ~n9990;
  assign n10594 = ~n10086 & n10593;
  assign n10595 = ~n33558 & ~n10594;
  assign n10596 = ~n9988 & n33558;
  assign n10597 = ~n9990 & n10596;
  assign n10598 = n33558 & n10594;
  assign n10599 = ~n10086 & n10597;
  assign n10600 = ~n10595 & ~n33641;
  assign n10601 = n330 & ~n10575;
  assign n10602 = ~n10590 & n10601;
  assign n10603 = n330 & n10591;
  assign n10604 = ~n10600 & ~n33642;
  assign n10605 = ~n10592 & ~n10604;
  assign n10606 = ~n271 & ~n10605;
  assign n10607 = n271 & ~n10592;
  assign n10608 = ~n10604 & n10607;
  assign n10609 = ~n10005 & ~n33560;
  assign n10610 = ~n10005 & ~n10086;
  assign n10611 = ~n33560 & n10610;
  assign n10612 = ~n10086 & n10609;
  assign n10613 = n10013 & ~n33643;
  assign n10614 = n10017 & n10610;
  assign n10615 = n10013 & ~n33560;
  assign n10616 = ~n10005 & n10615;
  assign n10617 = ~n10086 & n10616;
  assign n10618 = ~n10013 & ~n33643;
  assign n10619 = ~n10617 & ~n10618;
  assign n10620 = ~n10613 & ~n10614;
  assign n10621 = ~n10608 & ~n33644;
  assign n10622 = ~n10606 & ~n10621;
  assign n10623 = ~n217 & ~n10622;
  assign n10624 = n217 & ~n10606;
  assign n10625 = ~n10621 & n10624;
  assign n10626 = n217 & n10622;
  assign n10627 = ~n10019 & ~n10029;
  assign n10628 = ~n10019 & ~n10086;
  assign n10629 = ~n10029 & n10628;
  assign n10630 = ~n10086 & n10627;
  assign n10631 = n10027 & ~n33646;
  assign n10632 = n10030 & n10628;
  assign n10633 = ~n10019 & n10027;
  assign n10634 = ~n10029 & n10633;
  assign n10635 = ~n10086 & n10634;
  assign n10636 = ~n10027 & ~n33646;
  assign n10637 = ~n10635 & ~n10636;
  assign n10638 = ~n10631 & ~n10632;
  assign n10639 = ~n33645 & ~n33647;
  assign n10640 = ~n10623 & ~n10639;
  assign n10641 = ~n198 & ~n10640;
  assign n10642 = n198 & ~n10623;
  assign n10643 = ~n10639 & n10642;
  assign n10644 = ~n10032 & ~n33563;
  assign n10645 = ~n10032 & ~n10086;
  assign n10646 = ~n33563 & n10645;
  assign n10647 = ~n10086 & n10644;
  assign n10648 = n10040 & ~n33648;
  assign n10649 = n10044 & n10645;
  assign n10650 = n10040 & ~n33563;
  assign n10651 = ~n10032 & n10650;
  assign n10652 = ~n10086 & n10651;
  assign n10653 = ~n10040 & ~n33648;
  assign n10654 = ~n10652 & ~n10653;
  assign n10655 = ~n10648 & ~n10649;
  assign n10656 = ~n10643 & ~n33649;
  assign n10657 = ~n10641 & ~n10656;
  assign n10658 = ~n10046 & ~n10048;
  assign n10659 = ~n10086 & n10658;
  assign n10660 = ~n33565 & ~n10659;
  assign n10661 = ~n10046 & n33565;
  assign n10662 = ~n10048 & n10661;
  assign n10663 = n33565 & n10659;
  assign n10664 = ~n10086 & n10662;
  assign n10665 = ~n10660 & ~n33650;
  assign n10666 = ~n10062 & ~n10070;
  assign n10667 = ~n10070 & ~n10086;
  assign n10668 = ~n10062 & n10667;
  assign n10669 = ~n10086 & n10666;
  assign n10670 = ~n33568 & ~n33651;
  assign n10671 = ~n10665 & n10670;
  assign n10672 = ~n10657 & n10671;
  assign n10673 = n193 & ~n10672;
  assign n10674 = ~n10641 & n10665;
  assign n10675 = ~n10656 & n10674;
  assign n10676 = n10657 & n10665;
  assign n10677 = n10062 & ~n10667;
  assign n10678 = ~n193 & ~n10666;
  assign n10679 = ~n10677 & n10678;
  assign n10680 = ~n33652 & ~n10679;
  assign n10681 = ~n10673 & n10680;
  assign n10682 = ~n10214 & ~n10216;
  assign n10683 = ~n10681 & n10682;
  assign n10684 = ~n33570 & ~n10683;
  assign n10685 = n33570 & ~n10216;
  assign n10686 = ~n10214 & n10685;
  assign n10687 = n33570 & n10683;
  assign n10688 = ~n10681 & n10686;
  assign n10689 = ~n10684 & ~n33653;
  assign n10690 = ~n10184 & ~n10186;
  assign n10691 = ~n10681 & n10690;
  assign n10692 = ~n10194 & ~n10691;
  assign n10693 = ~n10186 & n10194;
  assign n10694 = ~n10184 & n10693;
  assign n10695 = n10194 & n10691;
  assign n10696 = ~n10681 & n10694;
  assign n10697 = ~n10692 & ~n33654;
  assign n10698 = ~n10150 & ~n10152;
  assign n10699 = ~n10681 & n10698;
  assign n10700 = ~n33578 & ~n10699;
  assign n10701 = ~n10152 & n33578;
  assign n10702 = ~n10150 & n10701;
  assign n10703 = n33578 & n10699;
  assign n10704 = ~n10681 & n10702;
  assign n10705 = ~n10700 & ~n33655;
  assign n10706 = ~n10123 & ~n10125;
  assign n10707 = ~n10681 & n10706;
  assign n10708 = ~n10134 & ~n10707;
  assign n10709 = ~n10125 & n10134;
  assign n10710 = ~n10123 & n10709;
  assign n10711 = n10134 & n10707;
  assign n10712 = ~n10681 & n10710;
  assign n10713 = ~n10708 & ~n33656;
  assign n10714 = ~pi54  & ~n10681;
  assign n10715 = ~pi55  & n10714;
  assign n10716 = n10100 & ~n10681;
  assign n10717 = ~n10086 & ~n10679;
  assign n10718 = ~n33652 & n10717;
  assign n10719 = ~n10673 & n10718;
  assign n10720 = ~n33657 & ~n10719;
  assign n10721 = pi56  & ~n10720;
  assign n10722 = ~pi56  & ~n10719;
  assign n10723 = ~pi56  & n10720;
  assign n10724 = ~n33657 & n10722;
  assign n10725 = ~n10721 & ~n33658;
  assign n10726 = pi54  & ~n10681;
  assign n10727 = ~pi52  & ~pi53 ;
  assign n10728 = ~pi54  & n10727;
  assign n10729 = ~n9546 & ~n33572;
  assign n10730 = ~n9547 & n10729;
  assign n10731 = ~n9563 & n10730;
  assign n10732 = ~n33501 & n10731;
  assign n10733 = n33499 & n9565;
  assign n10734 = ~n9557 & n10732;
  assign n10735 = ~n10728 & ~n33659;
  assign n10736 = ~n10084 & n10735;
  assign n10737 = ~n33568 & n10736;
  assign n10738 = ~n10078 & n10737;
  assign n10739 = ~n10726 & ~n10728;
  assign n10740 = n10086 & n10739;
  assign n10741 = ~n10726 & n10738;
  assign n10742 = pi55  & ~n10714;
  assign n10743 = ~n33657 & ~n10742;
  assign n10744 = ~n33660 & n10743;
  assign n10745 = ~n10086 & ~n10739;
  assign n10746 = n9565 & ~n10745;
  assign n10747 = ~n10744 & ~n10745;
  assign n10748 = n9565 & n10747;
  assign n10749 = ~n10744 & n10746;
  assign n10750 = ~n10725 & ~n33661;
  assign n10751 = ~n9565 & ~n10747;
  assign n10752 = n8998 & ~n10751;
  assign n10753 = ~n10750 & n10752;
  assign n10754 = ~n10103 & ~n33573;
  assign n10755 = ~n10681 & n10754;
  assign n10756 = n10108 & ~n10755;
  assign n10757 = ~n10108 & n10754;
  assign n10758 = ~n10108 & n10755;
  assign n10759 = ~n10681 & n10757;
  assign n10760 = ~n10756 & ~n33662;
  assign n10761 = ~n10753 & ~n10760;
  assign n10762 = ~n10750 & ~n10751;
  assign n10763 = ~n8998 & ~n10762;
  assign n10764 = n8506 & ~n10763;
  assign n10765 = ~n10761 & ~n10763;
  assign n10766 = n8506 & n10765;
  assign n10767 = ~n10761 & n10764;
  assign n10768 = ~n10713 & ~n33663;
  assign n10769 = ~n8506 & ~n10765;
  assign n10770 = n7975 & ~n10769;
  assign n10771 = ~n10768 & n10770;
  assign n10772 = ~n10137 & ~n33575;
  assign n10773 = ~n10681 & n10772;
  assign n10774 = n10147 & ~n10773;
  assign n10775 = ~n10147 & n10773;
  assign n10776 = ~n10137 & n10147;
  assign n10777 = ~n33575 & n10776;
  assign n10778 = n10147 & n10773;
  assign n10779 = ~n10681 & n10777;
  assign n10780 = ~n10147 & ~n10773;
  assign n10781 = ~n33664 & ~n10780;
  assign n10782 = ~n10774 & ~n10775;
  assign n10783 = ~n10771 & ~n33665;
  assign n10784 = ~n10768 & ~n10769;
  assign n10785 = ~n7975 & ~n10784;
  assign n10786 = n7512 & ~n10785;
  assign n10787 = ~n10783 & ~n10785;
  assign n10788 = n7512 & n10787;
  assign n10789 = ~n10783 & n10786;
  assign n10790 = ~n10705 & ~n33666;
  assign n10791 = ~n7512 & ~n10787;
  assign n10792 = n7015 & ~n10791;
  assign n10793 = ~n10790 & n10792;
  assign n10794 = ~n10167 & ~n33579;
  assign n10795 = ~n10681 & n10794;
  assign n10796 = ~n33581 & n10795;
  assign n10797 = n33581 & ~n10795;
  assign n10798 = ~n10167 & n33581;
  assign n10799 = ~n33579 & n10798;
  assign n10800 = ~n10681 & n10799;
  assign n10801 = ~n33581 & ~n10795;
  assign n10802 = ~n10800 & ~n10801;
  assign n10803 = ~n10796 & ~n10797;
  assign n10804 = ~n10793 & ~n33667;
  assign n10805 = ~n10790 & ~n10791;
  assign n10806 = ~n7015 & ~n10805;
  assign n10807 = n6579 & ~n10806;
  assign n10808 = ~n10804 & ~n10806;
  assign n10809 = n6579 & n10808;
  assign n10810 = ~n10804 & n10807;
  assign n10811 = ~n10697 & ~n33668;
  assign n10812 = ~n6579 & ~n10808;
  assign n10813 = ~n10811 & ~n10812;
  assign n10814 = ~n6117 & ~n10813;
  assign n10815 = n6117 & ~n10812;
  assign n10816 = ~n10811 & n10815;
  assign n10817 = ~n10197 & ~n33583;
  assign n10818 = ~n10681 & n10817;
  assign n10819 = ~n33585 & ~n10818;
  assign n10820 = ~n10197 & n33585;
  assign n10821 = ~n33583 & n10820;
  assign n10822 = n33585 & n10818;
  assign n10823 = ~n10681 & n10821;
  assign n10824 = n33585 & ~n10818;
  assign n10825 = ~n33585 & n10818;
  assign n10826 = ~n10824 & ~n10825;
  assign n10827 = ~n10819 & ~n33669;
  assign n10828 = ~n10816 & n33670;
  assign n10829 = ~n10814 & ~n10828;
  assign n10830 = ~n5708 & ~n10829;
  assign n10831 = n5708 & ~n10814;
  assign n10832 = n5708 & n10829;
  assign n10833 = ~n10828 & n10831;
  assign n10834 = ~n10689 & ~n33671;
  assign n10835 = ~n10830 & ~n10834;
  assign n10836 = ~n5278 & ~n10835;
  assign n10837 = n5278 & ~n10830;
  assign n10838 = ~n10834 & n10837;
  assign n10839 = ~n10219 & ~n33586;
  assign n10840 = ~n10681 & n10839;
  assign n10841 = ~n33588 & ~n10840;
  assign n10842 = n33588 & n10840;
  assign n10843 = ~n10219 & ~n33588;
  assign n10844 = ~n33586 & n10843;
  assign n10845 = ~n33588 & n10840;
  assign n10846 = ~n10681 & n10844;
  assign n10847 = n33588 & ~n10840;
  assign n10848 = ~n33672 & ~n10847;
  assign n10849 = ~n10841 & ~n10842;
  assign n10850 = ~n10838 & ~n33673;
  assign n10851 = ~n10836 & ~n10850;
  assign n10852 = ~n4903 & ~n10851;
  assign n10853 = ~n10236 & ~n10238;
  assign n10854 = ~n10681 & n10853;
  assign n10855 = ~n33590 & ~n10854;
  assign n10856 = ~n10238 & n33590;
  assign n10857 = ~n10236 & n10856;
  assign n10858 = n33590 & n10854;
  assign n10859 = ~n10681 & n10857;
  assign n10860 = ~n10855 & ~n33674;
  assign n10861 = n4903 & ~n10836;
  assign n10862 = n4903 & n10851;
  assign n10863 = ~n10850 & n10861;
  assign n10864 = ~n10860 & ~n33675;
  assign n10865 = ~n10852 & ~n10864;
  assign n10866 = ~n4508 & ~n10865;
  assign n10867 = n4508 & ~n10852;
  assign n10868 = ~n10864 & n10867;
  assign n10869 = ~n10253 & ~n33591;
  assign n10870 = ~n10253 & ~n10681;
  assign n10871 = ~n33591 & n10870;
  assign n10872 = ~n10681 & n10869;
  assign n10873 = ~n33593 & ~n33676;
  assign n10874 = n10268 & n10870;
  assign n10875 = n33593 & n33676;
  assign n10876 = ~n10253 & ~n33593;
  assign n10877 = ~n33591 & n10876;
  assign n10878 = ~n10681 & n10877;
  assign n10879 = n33593 & ~n33676;
  assign n10880 = ~n10878 & ~n10879;
  assign n10881 = ~n10873 & ~n33677;
  assign n10882 = ~n10868 & ~n33678;
  assign n10883 = ~n10866 & ~n10882;
  assign n10884 = ~n4155 & ~n10883;
  assign n10885 = ~n10270 & ~n10272;
  assign n10886 = ~n10681 & n10885;
  assign n10887 = ~n33595 & ~n10886;
  assign n10888 = ~n10272 & n33595;
  assign n10889 = ~n10270 & n10888;
  assign n10890 = n33595 & n10886;
  assign n10891 = ~n10681 & n10889;
  assign n10892 = ~n10887 & ~n33679;
  assign n10893 = n4155 & ~n10866;
  assign n10894 = n4155 & n10883;
  assign n10895 = ~n10882 & n10893;
  assign n10896 = ~n10892 & ~n33680;
  assign n10897 = ~n10884 & ~n10896;
  assign n10898 = ~n3788 & ~n10897;
  assign n10899 = n3788 & ~n10884;
  assign n10900 = ~n10896 & n10899;
  assign n10901 = ~n10287 & ~n33596;
  assign n10902 = ~n10681 & n10901;
  assign n10903 = ~n33599 & ~n10902;
  assign n10904 = ~n10287 & n33599;
  assign n10905 = ~n33596 & n10904;
  assign n10906 = n33599 & n10902;
  assign n10907 = ~n10681 & n10905;
  assign n10908 = ~n10903 & ~n33681;
  assign n10909 = ~n10900 & ~n10908;
  assign n10910 = ~n10898 & ~n10909;
  assign n10911 = ~n3473 & ~n10910;
  assign n10912 = ~n10306 & ~n10308;
  assign n10913 = ~n10681 & n10912;
  assign n10914 = ~n33601 & ~n10913;
  assign n10915 = ~n10308 & n33601;
  assign n10916 = ~n10306 & n10915;
  assign n10917 = n33601 & n10913;
  assign n10918 = ~n10681 & n10916;
  assign n10919 = ~n10914 & ~n33682;
  assign n10920 = n3473 & ~n10898;
  assign n10921 = n3473 & n10910;
  assign n10922 = ~n10909 & n10920;
  assign n10923 = ~n10919 & ~n33683;
  assign n10924 = ~n10911 & ~n10923;
  assign n10925 = ~n3140 & ~n10924;
  assign n10926 = n3140 & ~n10911;
  assign n10927 = ~n10923 & n10926;
  assign n10928 = ~n10323 & ~n33602;
  assign n10929 = ~n10323 & ~n10681;
  assign n10930 = ~n33602 & n10929;
  assign n10931 = ~n10681 & n10928;
  assign n10932 = n10334 & ~n33684;
  assign n10933 = n10335 & n10929;
  assign n10934 = ~n10334 & n33684;
  assign n10935 = ~n10323 & n10334;
  assign n10936 = ~n33602 & n10935;
  assign n10937 = ~n10681 & n10936;
  assign n10938 = ~n10334 & ~n33684;
  assign n10939 = ~n10937 & ~n10938;
  assign n10940 = ~n10932 & ~n33685;
  assign n10941 = ~n10927 & ~n33686;
  assign n10942 = ~n10925 & ~n10941;
  assign n10943 = ~n2855 & ~n10942;
  assign n10944 = ~n10337 & ~n10339;
  assign n10945 = ~n10681 & n10944;
  assign n10946 = ~n33605 & ~n10945;
  assign n10947 = ~n10339 & n33605;
  assign n10948 = ~n10337 & n10947;
  assign n10949 = n33605 & n10945;
  assign n10950 = ~n10681 & n10948;
  assign n10951 = ~n10946 & ~n33687;
  assign n10952 = n2855 & ~n10925;
  assign n10953 = n2855 & n10942;
  assign n10954 = ~n10941 & n10952;
  assign n10955 = ~n10951 & ~n33688;
  assign n10956 = ~n10943 & ~n10955;
  assign n10957 = ~n2556 & ~n10956;
  assign n10958 = n2556 & ~n10943;
  assign n10959 = ~n10955 & n10958;
  assign n10960 = ~n10354 & ~n33606;
  assign n10961 = ~n10681 & n10960;
  assign n10962 = ~n33609 & n10961;
  assign n10963 = n33609 & ~n10961;
  assign n10964 = ~n10354 & n33609;
  assign n10965 = ~n33606 & n10964;
  assign n10966 = n33609 & n10961;
  assign n10967 = ~n10681 & n10965;
  assign n10968 = ~n33609 & ~n10961;
  assign n10969 = ~n33689 & ~n10968;
  assign n10970 = ~n10962 & ~n10963;
  assign n10971 = ~n10959 & ~n33690;
  assign n10972 = ~n10957 & ~n10971;
  assign n10973 = ~n2301 & ~n10972;
  assign n10974 = ~n10373 & ~n10375;
  assign n10975 = ~n10681 & n10974;
  assign n10976 = ~n33611 & ~n10975;
  assign n10977 = ~n10375 & n33611;
  assign n10978 = ~n10373 & n10977;
  assign n10979 = n33611 & n10975;
  assign n10980 = ~n10681 & n10978;
  assign n10981 = ~n10976 & ~n33691;
  assign n10982 = n2301 & ~n10957;
  assign n10983 = n2301 & n10972;
  assign n10984 = ~n10971 & n10982;
  assign n10985 = ~n10981 & ~n33692;
  assign n10986 = ~n10973 & ~n10985;
  assign n10987 = ~n2038 & ~n10986;
  assign n10988 = n2038 & ~n10973;
  assign n10989 = ~n10985 & n10988;
  assign n10990 = ~n10390 & ~n33612;
  assign n10991 = ~n10390 & ~n10681;
  assign n10992 = ~n33612 & n10991;
  assign n10993 = ~n10681 & n10990;
  assign n10994 = n33614 & ~n33693;
  assign n10995 = n10405 & n10991;
  assign n10996 = ~n33614 & n33693;
  assign n10997 = ~n10390 & n33614;
  assign n10998 = ~n33612 & n10997;
  assign n10999 = ~n10681 & n10998;
  assign n11000 = ~n33614 & ~n33693;
  assign n11001 = ~n10999 & ~n11000;
  assign n11002 = ~n10994 & ~n33694;
  assign n11003 = ~n10989 & ~n33695;
  assign n11004 = ~n10987 & ~n11003;
  assign n11005 = ~n1812 & ~n11004;
  assign n11006 = ~n10407 & ~n10409;
  assign n11007 = ~n10681 & n11006;
  assign n11008 = ~n33616 & ~n11007;
  assign n11009 = ~n10409 & n33616;
  assign n11010 = ~n10407 & n11009;
  assign n11011 = n33616 & n11007;
  assign n11012 = ~n10681 & n11010;
  assign n11013 = ~n11008 & ~n33696;
  assign n11014 = n1812 & ~n10987;
  assign n11015 = n1812 & n11004;
  assign n11016 = ~n11003 & n11014;
  assign n11017 = ~n11013 & ~n33697;
  assign n11018 = ~n11005 & ~n11017;
  assign n11019 = ~n1582 & ~n11018;
  assign n11020 = ~n10424 & ~n33617;
  assign n11021 = ~n10681 & n11020;
  assign n11022 = ~n33620 & ~n11021;
  assign n11023 = ~n10424 & n33620;
  assign n11024 = ~n33617 & n11023;
  assign n11025 = n33620 & n11021;
  assign n11026 = ~n10681 & n11024;
  assign n11027 = ~n11022 & ~n33698;
  assign n11028 = n1582 & ~n11005;
  assign n11029 = ~n11017 & n11028;
  assign n11030 = ~n11027 & ~n11029;
  assign n11031 = ~n11019 & ~n11030;
  assign n11032 = ~n1388 & ~n11031;
  assign n11033 = ~n10443 & ~n10445;
  assign n11034 = ~n10681 & n11033;
  assign n11035 = ~n33622 & ~n11034;
  assign n11036 = ~n10445 & n33622;
  assign n11037 = ~n10443 & n11036;
  assign n11038 = n33622 & n11034;
  assign n11039 = ~n10681 & n11037;
  assign n11040 = ~n11035 & ~n33699;
  assign n11041 = n1388 & ~n11019;
  assign n11042 = n1388 & n11031;
  assign n11043 = ~n11030 & n11041;
  assign n11044 = ~n11040 & ~n33700;
  assign n11045 = ~n11032 & ~n11044;
  assign n11046 = ~n1192 & ~n11045;
  assign n11047 = n1192 & ~n11032;
  assign n11048 = ~n11044 & n11047;
  assign n11049 = ~n10460 & ~n33624;
  assign n11050 = ~n10460 & ~n10681;
  assign n11051 = ~n33624 & n11050;
  assign n11052 = ~n10681 & n11049;
  assign n11053 = n10468 & ~n33701;
  assign n11054 = n10472 & n11050;
  assign n11055 = ~n10460 & n10468;
  assign n11056 = ~n33624 & n11055;
  assign n11057 = ~n10681 & n11056;
  assign n11058 = ~n10468 & ~n33701;
  assign n11059 = ~n11057 & ~n11058;
  assign n11060 = ~n11053 & ~n11054;
  assign n11061 = ~n11048 & ~n33702;
  assign n11062 = ~n11046 & ~n11061;
  assign n11063 = ~n1028 & ~n11062;
  assign n11064 = ~n10474 & ~n10476;
  assign n11065 = ~n10681 & n11064;
  assign n11066 = ~n33626 & ~n11065;
  assign n11067 = ~n10476 & n33626;
  assign n11068 = ~n10474 & n11067;
  assign n11069 = n33626 & n11065;
  assign n11070 = ~n10681 & n11068;
  assign n11071 = ~n11066 & ~n33703;
  assign n11072 = n1028 & ~n11046;
  assign n11073 = n1028 & n11062;
  assign n11074 = ~n11061 & n11072;
  assign n11075 = ~n11071 & ~n33704;
  assign n11076 = ~n11063 & ~n11075;
  assign n11077 = ~n866 & ~n11076;
  assign n11078 = ~n10491 & ~n33627;
  assign n11079 = ~n10681 & n11078;
  assign n11080 = ~n33629 & ~n11079;
  assign n11081 = ~n10491 & n33629;
  assign n11082 = ~n33627 & n11081;
  assign n11083 = n33629 & n11079;
  assign n11084 = ~n10681 & n11082;
  assign n11085 = ~n11080 & ~n33705;
  assign n11086 = n866 & ~n11063;
  assign n11087 = ~n11075 & n11086;
  assign n11088 = ~n11085 & ~n11087;
  assign n11089 = ~n11077 & ~n11088;
  assign n11090 = ~n730 & ~n11089;
  assign n11091 = ~n10509 & ~n10511;
  assign n11092 = ~n10681 & n11091;
  assign n11093 = ~n33631 & ~n11092;
  assign n11094 = ~n10511 & n33631;
  assign n11095 = ~n10509 & n11094;
  assign n11096 = n33631 & n11092;
  assign n11097 = ~n10681 & n11095;
  assign n11098 = ~n11093 & ~n33706;
  assign n11099 = n730 & ~n11077;
  assign n11100 = n730 & n11089;
  assign n11101 = ~n11088 & n11099;
  assign n11102 = ~n11098 & ~n33707;
  assign n11103 = ~n11090 & ~n11102;
  assign n11104 = ~n602 & ~n11103;
  assign n11105 = n602 & ~n11090;
  assign n11106 = ~n11102 & n11105;
  assign n11107 = ~n10526 & ~n33633;
  assign n11108 = ~n10526 & ~n10681;
  assign n11109 = ~n33633 & n11108;
  assign n11110 = ~n10681 & n11107;
  assign n11111 = n10534 & ~n33708;
  assign n11112 = n10538 & n11108;
  assign n11113 = ~n10526 & n10534;
  assign n11114 = ~n33633 & n11113;
  assign n11115 = ~n10681 & n11114;
  assign n11116 = ~n10534 & ~n33708;
  assign n11117 = ~n11115 & ~n11116;
  assign n11118 = ~n11111 & ~n11112;
  assign n11119 = ~n11106 & ~n33709;
  assign n11120 = ~n11104 & ~n11119;
  assign n11121 = ~n497 & ~n11120;
  assign n11122 = ~n10540 & ~n10542;
  assign n11123 = ~n10681 & n11122;
  assign n11124 = ~n33635 & ~n11123;
  assign n11125 = ~n10542 & n33635;
  assign n11126 = ~n10540 & n11125;
  assign n11127 = n33635 & n11123;
  assign n11128 = ~n10681 & n11126;
  assign n11129 = ~n11124 & ~n33710;
  assign n11130 = n497 & ~n11104;
  assign n11131 = n497 & n11120;
  assign n11132 = ~n11119 & n11130;
  assign n11133 = ~n11129 & ~n33711;
  assign n11134 = ~n11121 & ~n11133;
  assign n11135 = ~n403 & ~n11134;
  assign n11136 = ~n10557 & ~n33636;
  assign n11137 = ~n10681 & n11136;
  assign n11138 = ~n33638 & ~n11137;
  assign n11139 = ~n10557 & n33638;
  assign n11140 = ~n33636 & n11139;
  assign n11141 = n33638 & n11137;
  assign n11142 = ~n10681 & n11140;
  assign n11143 = ~n11138 & ~n33712;
  assign n11144 = n403 & ~n11121;
  assign n11145 = ~n11133 & n11144;
  assign n11146 = ~n11143 & ~n11145;
  assign n11147 = ~n11135 & ~n11146;
  assign n11148 = ~n330 & ~n11147;
  assign n11149 = ~n10575 & ~n10577;
  assign n11150 = ~n10681 & n11149;
  assign n11151 = ~n33640 & ~n11150;
  assign n11152 = ~n10577 & n33640;
  assign n11153 = ~n10575 & n11152;
  assign n11154 = n33640 & n11150;
  assign n11155 = ~n10681 & n11153;
  assign n11156 = ~n11151 & ~n33713;
  assign n11157 = n330 & ~n11135;
  assign n11158 = n330 & n11147;
  assign n11159 = ~n11146 & n11157;
  assign n11160 = ~n11156 & ~n33714;
  assign n11161 = ~n11148 & ~n11160;
  assign n11162 = ~n271 & ~n11161;
  assign n11163 = n271 & ~n11148;
  assign n11164 = ~n11160 & n11163;
  assign n11165 = ~n10592 & ~n33642;
  assign n11166 = ~n10592 & ~n10681;
  assign n11167 = ~n33642 & n11166;
  assign n11168 = ~n10681 & n11165;
  assign n11169 = n10600 & ~n33715;
  assign n11170 = n10604 & n11166;
  assign n11171 = ~n10592 & n10600;
  assign n11172 = ~n33642 & n11171;
  assign n11173 = ~n10681 & n11172;
  assign n11174 = ~n10600 & ~n33715;
  assign n11175 = ~n11173 & ~n11174;
  assign n11176 = ~n11169 & ~n11170;
  assign n11177 = ~n11164 & ~n33716;
  assign n11178 = ~n11162 & ~n11177;
  assign n11179 = ~n217 & ~n11178;
  assign n11180 = ~n10606 & ~n10608;
  assign n11181 = ~n10681 & n11180;
  assign n11182 = ~n33644 & ~n11181;
  assign n11183 = ~n10608 & n33644;
  assign n11184 = ~n10606 & n11183;
  assign n11185 = n33644 & n11181;
  assign n11186 = ~n10681 & n11184;
  assign n11187 = ~n11182 & ~n33717;
  assign n11188 = n217 & ~n11162;
  assign n11189 = n217 & n11178;
  assign n11190 = ~n11177 & n11188;
  assign n11191 = ~n11187 & ~n33718;
  assign n11192 = ~n11179 & ~n11191;
  assign n11193 = ~n198 & ~n11192;
  assign n11194 = ~n10623 & ~n33645;
  assign n11195 = ~n10681 & n11194;
  assign n11196 = ~n33647 & ~n11195;
  assign n11197 = ~n10623 & n33647;
  assign n11198 = ~n33645 & n11197;
  assign n11199 = n33647 & n11195;
  assign n11200 = ~n10681 & n11198;
  assign n11201 = ~n11196 & ~n33719;
  assign n11202 = n198 & ~n11179;
  assign n11203 = ~n11191 & n11202;
  assign n11204 = ~n11201 & ~n11203;
  assign n11205 = ~n11193 & ~n11204;
  assign n11206 = ~n10641 & ~n10643;
  assign n11207 = ~n10681 & n11206;
  assign n11208 = ~n33649 & ~n11207;
  assign n11209 = ~n10643 & n33649;
  assign n11210 = ~n10641 & n11209;
  assign n11211 = n33649 & n11207;
  assign n11212 = ~n10681 & n11210;
  assign n11213 = ~n11208 & ~n33720;
  assign n11214 = ~n10657 & ~n10665;
  assign n11215 = ~n10665 & ~n10681;
  assign n11216 = ~n10657 & n11215;
  assign n11217 = ~n10681 & n11214;
  assign n11218 = ~n33652 & ~n33721;
  assign n11219 = ~n11213 & n11218;
  assign n11220 = ~n11205 & n11219;
  assign n11221 = n193 & ~n11220;
  assign n11222 = ~n11193 & n11213;
  assign n11223 = n11205 & n11213;
  assign n11224 = ~n11204 & n11222;
  assign n11225 = n10657 & ~n11215;
  assign n11226 = ~n193 & ~n11214;
  assign n11227 = ~n11225 & n11226;
  assign n11228 = ~n33722 & ~n11227;
  assign n11229 = ~n11221 & n11228;
  assign n11230 = ~n10830 & ~n33671;
  assign n11231 = ~n10830 & ~n11229;
  assign n11232 = ~n33671 & n11231;
  assign n11233 = ~n11229 & n11230;
  assign n11234 = n10689 & ~n33723;
  assign n11235 = n10834 & n11231;
  assign n11236 = n10689 & ~n33671;
  assign n11237 = ~n10830 & n11236;
  assign n11238 = ~n11229 & n11237;
  assign n11239 = ~n10689 & ~n33723;
  assign n11240 = ~n11238 & ~n11239;
  assign n11241 = ~n11234 & ~n11235;
  assign n11242 = pi52  & ~n11229;
  assign n11243 = ~pi50  & ~pi51 ;
  assign n11244 = ~pi52  & n11243;
  assign n11245 = ~n11242 & ~n11244;
  assign n11246 = ~n10681 & ~n11245;
  assign n11247 = ~pi52  & ~n11229;
  assign n11248 = pi53  & ~n11247;
  assign n11249 = ~pi53  & n11247;
  assign n11250 = n10727 & ~n11229;
  assign n11251 = ~n11248 & ~n33725;
  assign n11252 = ~n33566 & ~n33659;
  assign n11253 = ~n10065 & n11252;
  assign n11254 = ~n10084 & n11253;
  assign n11255 = ~n33568 & n11254;
  assign n11256 = n10070 & n10086;
  assign n11257 = ~n10078 & n11255;
  assign n11258 = ~n11244 & ~n33726;
  assign n11259 = ~n10679 & n11258;
  assign n11260 = ~n33652 & n11259;
  assign n11261 = ~n10673 & n11260;
  assign n11262 = n10681 & n11245;
  assign n11263 = ~n11242 & n11261;
  assign n11264 = n11251 & ~n33727;
  assign n11265 = ~n11246 & ~n11264;
  assign n11266 = ~n10086 & ~n11265;
  assign n11267 = n10086 & ~n11246;
  assign n11268 = ~n11264 & n11267;
  assign n11269 = ~n10681 & ~n11227;
  assign n11270 = ~n33722 & n11269;
  assign n11271 = ~n11221 & n11270;
  assign n11272 = ~n33725 & ~n11271;
  assign n11273 = pi54  & ~n11272;
  assign n11274 = ~pi54  & ~n11271;
  assign n11275 = ~pi54  & n11272;
  assign n11276 = ~n33725 & n11274;
  assign n11277 = ~n11273 & ~n33728;
  assign n11278 = ~n11268 & ~n11277;
  assign n11279 = ~n11266 & ~n11278;
  assign n11280 = ~n9565 & ~n11279;
  assign n11281 = n9565 & ~n11266;
  assign n11282 = ~n11278 & n11281;
  assign n11283 = n9565 & n11279;
  assign n11284 = ~n33660 & ~n10745;
  assign n11285 = ~n11229 & n11284;
  assign n11286 = n10743 & ~n11285;
  assign n11287 = ~n10743 & n11284;
  assign n11288 = ~n10743 & n11285;
  assign n11289 = ~n11229 & n11287;
  assign n11290 = ~n11286 & ~n33730;
  assign n11291 = ~n33729 & ~n11290;
  assign n11292 = ~n11280 & ~n11291;
  assign n11293 = ~n8998 & ~n11292;
  assign n11294 = n8998 & ~n11280;
  assign n11295 = ~n11291 & n11294;
  assign n11296 = ~n33661 & ~n10751;
  assign n11297 = ~n10751 & ~n11229;
  assign n11298 = ~n33661 & n11297;
  assign n11299 = ~n11229 & n11296;
  assign n11300 = n10725 & ~n33731;
  assign n11301 = n10750 & n11297;
  assign n11302 = n10725 & ~n33661;
  assign n11303 = ~n10751 & n11302;
  assign n11304 = ~n11229 & n11303;
  assign n11305 = ~n10725 & ~n33731;
  assign n11306 = ~n11304 & ~n11305;
  assign n11307 = ~n11300 & ~n11301;
  assign n11308 = ~n11295 & ~n33732;
  assign n11309 = ~n11293 & ~n11308;
  assign n11310 = ~n8506 & ~n11309;
  assign n11311 = n8506 & ~n11293;
  assign n11312 = ~n11308 & n11311;
  assign n11313 = n8506 & n11309;
  assign n11314 = ~n10753 & ~n10763;
  assign n11315 = ~n11229 & n11314;
  assign n11316 = n10760 & ~n11315;
  assign n11317 = ~n10760 & n11315;
  assign n11318 = n10760 & ~n10763;
  assign n11319 = ~n10753 & n11318;
  assign n11320 = n10760 & n11315;
  assign n11321 = ~n11229 & n11319;
  assign n11322 = ~n10760 & ~n11315;
  assign n11323 = ~n33734 & ~n11322;
  assign n11324 = ~n11316 & ~n11317;
  assign n11325 = ~n33733 & ~n33735;
  assign n11326 = ~n11310 & ~n11325;
  assign n11327 = ~n7975 & ~n11326;
  assign n11328 = n7975 & ~n11310;
  assign n11329 = ~n11325 & n11328;
  assign n11330 = ~n33663 & ~n10769;
  assign n11331 = ~n10769 & ~n11229;
  assign n11332 = ~n33663 & n11331;
  assign n11333 = ~n11229 & n11330;
  assign n11334 = n10713 & ~n33736;
  assign n11335 = n10768 & n11331;
  assign n11336 = n10713 & ~n33663;
  assign n11337 = ~n10769 & n11336;
  assign n11338 = ~n11229 & n11337;
  assign n11339 = ~n10713 & ~n33736;
  assign n11340 = ~n11338 & ~n11339;
  assign n11341 = ~n11334 & ~n11335;
  assign n11342 = ~n11329 & ~n33737;
  assign n11343 = ~n11327 & ~n11342;
  assign n11344 = ~n7512 & ~n11343;
  assign n11345 = n7512 & ~n11327;
  assign n11346 = ~n11342 & n11345;
  assign n11347 = n7512 & n11343;
  assign n11348 = ~n10771 & ~n10785;
  assign n11349 = ~n11229 & n11348;
  assign n11350 = ~n33665 & n11349;
  assign n11351 = n33665 & ~n11349;
  assign n11352 = n33665 & ~n10785;
  assign n11353 = ~n10771 & n11352;
  assign n11354 = ~n11229 & n11353;
  assign n11355 = ~n33665 & ~n11349;
  assign n11356 = ~n11354 & ~n11355;
  assign n11357 = ~n11350 & ~n11351;
  assign n11358 = ~n33738 & ~n33739;
  assign n11359 = ~n11344 & ~n11358;
  assign n11360 = ~n7015 & ~n11359;
  assign n11361 = n7015 & ~n11344;
  assign n11362 = ~n11358 & n11361;
  assign n11363 = ~n33666 & ~n10791;
  assign n11364 = ~n10791 & ~n11229;
  assign n11365 = ~n33666 & n11364;
  assign n11366 = ~n11229 & n11363;
  assign n11367 = n10705 & ~n33740;
  assign n11368 = n10790 & n11364;
  assign n11369 = n10705 & ~n33666;
  assign n11370 = ~n10791 & n11369;
  assign n11371 = ~n11229 & n11370;
  assign n11372 = ~n10705 & ~n33740;
  assign n11373 = ~n11371 & ~n11372;
  assign n11374 = ~n11367 & ~n11368;
  assign n11375 = ~n11362 & ~n33741;
  assign n11376 = ~n11360 & ~n11375;
  assign n11377 = ~n6579 & ~n11376;
  assign n11378 = n6579 & ~n11360;
  assign n11379 = ~n11375 & n11378;
  assign n11380 = n6579 & n11376;
  assign n11381 = ~n10793 & ~n10806;
  assign n11382 = ~n11229 & n11381;
  assign n11383 = ~n33667 & ~n11382;
  assign n11384 = n33667 & ~n10806;
  assign n11385 = ~n10793 & n11384;
  assign n11386 = n33667 & n11382;
  assign n11387 = ~n11229 & n11385;
  assign n11388 = n33667 & ~n11382;
  assign n11389 = ~n33667 & n11382;
  assign n11390 = ~n11388 & ~n11389;
  assign n11391 = ~n11383 & ~n33743;
  assign n11392 = ~n33742 & n33744;
  assign n11393 = ~n11377 & ~n11392;
  assign n11394 = ~n6117 & ~n11393;
  assign n11395 = n6117 & ~n11377;
  assign n11396 = ~n11392 & n11395;
  assign n11397 = ~n33668 & ~n10812;
  assign n11398 = ~n11229 & n11397;
  assign n11399 = n10697 & ~n11398;
  assign n11400 = ~n10697 & n11398;
  assign n11401 = n10697 & ~n33668;
  assign n11402 = ~n10812 & n11401;
  assign n11403 = ~n11229 & n11402;
  assign n11404 = ~n10697 & ~n11398;
  assign n11405 = ~n11403 & ~n11404;
  assign n11406 = ~n11399 & ~n11400;
  assign n11407 = ~n11396 & ~n33745;
  assign n11408 = ~n11394 & ~n11407;
  assign n11409 = ~n5708 & ~n11408;
  assign n11410 = ~n10814 & ~n10816;
  assign n11411 = ~n11229 & n11410;
  assign n11412 = n33670 & ~n11411;
  assign n11413 = ~n10814 & ~n33670;
  assign n11414 = ~n10816 & n11413;
  assign n11415 = ~n33670 & n11411;
  assign n11416 = ~n11229 & n11414;
  assign n11417 = n33670 & n11411;
  assign n11418 = ~n33670 & ~n11411;
  assign n11419 = ~n11417 & ~n11418;
  assign n11420 = ~n11412 & ~n33746;
  assign n11421 = n5708 & ~n11394;
  assign n11422 = ~n11407 & n11421;
  assign n11423 = n5708 & n11408;
  assign n11424 = n33747 & ~n33748;
  assign n11425 = ~n11409 & ~n11424;
  assign n11426 = ~n5278 & ~n11425;
  assign n11427 = n5278 & ~n11409;
  assign n11428 = ~n11424 & n11427;
  assign n11429 = ~n33724 & ~n11428;
  assign n11430 = ~n11426 & ~n11429;
  assign n11431 = ~n4903 & ~n11430;
  assign n11432 = n4903 & ~n11426;
  assign n11433 = ~n11429 & n11432;
  assign n11434 = n4903 & n11430;
  assign n11435 = ~n10836 & ~n10838;
  assign n11436 = ~n11229 & n11435;
  assign n11437 = ~n33673 & n11436;
  assign n11438 = n33673 & ~n11436;
  assign n11439 = ~n10836 & n33673;
  assign n11440 = ~n10838 & n11439;
  assign n11441 = n33673 & n11436;
  assign n11442 = ~n11229 & n11440;
  assign n11443 = ~n33673 & ~n11436;
  assign n11444 = ~n33750 & ~n11443;
  assign n11445 = ~n11437 & ~n11438;
  assign n11446 = ~n33749 & ~n33751;
  assign n11447 = ~n11431 & ~n11446;
  assign n11448 = ~n4508 & ~n11447;
  assign n11449 = n4508 & ~n11431;
  assign n11450 = ~n11446 & n11449;
  assign n11451 = ~n10852 & ~n33675;
  assign n11452 = ~n10852 & ~n11229;
  assign n11453 = ~n33675 & n11452;
  assign n11454 = ~n11229 & n11451;
  assign n11455 = n10860 & ~n33752;
  assign n11456 = n10864 & n11452;
  assign n11457 = n10860 & ~n33675;
  assign n11458 = ~n10852 & n11457;
  assign n11459 = ~n11229 & n11458;
  assign n11460 = ~n10860 & ~n33752;
  assign n11461 = ~n11459 & ~n11460;
  assign n11462 = ~n11455 & ~n11456;
  assign n11463 = ~n11450 & ~n33753;
  assign n11464 = ~n11448 & ~n11463;
  assign n11465 = ~n4155 & ~n11464;
  assign n11466 = n4155 & ~n11448;
  assign n11467 = ~n11463 & n11466;
  assign n11468 = n4155 & n11464;
  assign n11469 = ~n10866 & ~n10868;
  assign n11470 = ~n11229 & n11469;
  assign n11471 = ~n33678 & ~n11470;
  assign n11472 = ~n10866 & n33678;
  assign n11473 = ~n10868 & n11472;
  assign n11474 = n33678 & n11470;
  assign n11475 = ~n11229 & n11473;
  assign n11476 = ~n11471 & ~n33755;
  assign n11477 = ~n33754 & ~n11476;
  assign n11478 = ~n11465 & ~n11477;
  assign n11479 = ~n3788 & ~n11478;
  assign n11480 = n3788 & ~n11465;
  assign n11481 = ~n11477 & n11480;
  assign n11482 = ~n10884 & ~n33680;
  assign n11483 = ~n10884 & ~n11229;
  assign n11484 = ~n33680 & n11483;
  assign n11485 = ~n11229 & n11482;
  assign n11486 = n10892 & ~n33756;
  assign n11487 = n10896 & n11483;
  assign n11488 = n10892 & ~n33680;
  assign n11489 = ~n10884 & n11488;
  assign n11490 = ~n11229 & n11489;
  assign n11491 = ~n10892 & ~n33756;
  assign n11492 = ~n11490 & ~n11491;
  assign n11493 = ~n11486 & ~n11487;
  assign n11494 = ~n11481 & ~n33757;
  assign n11495 = ~n11479 & ~n11494;
  assign n11496 = ~n3473 & ~n11495;
  assign n11497 = n3473 & ~n11479;
  assign n11498 = ~n11494 & n11497;
  assign n11499 = n3473 & n11495;
  assign n11500 = ~n10898 & ~n10900;
  assign n11501 = ~n10898 & ~n11229;
  assign n11502 = ~n10900 & n11501;
  assign n11503 = ~n11229 & n11500;
  assign n11504 = n10908 & ~n33759;
  assign n11505 = n10909 & n11501;
  assign n11506 = ~n10908 & n33759;
  assign n11507 = ~n10898 & n10908;
  assign n11508 = ~n10900 & n11507;
  assign n11509 = ~n11229 & n11508;
  assign n11510 = ~n10908 & ~n33759;
  assign n11511 = ~n11509 & ~n11510;
  assign n11512 = ~n11504 & ~n33760;
  assign n11513 = ~n33758 & ~n33761;
  assign n11514 = ~n11496 & ~n11513;
  assign n11515 = ~n3140 & ~n11514;
  assign n11516 = n3140 & ~n11496;
  assign n11517 = ~n11513 & n11516;
  assign n11518 = ~n10911 & ~n33683;
  assign n11519 = ~n10911 & ~n11229;
  assign n11520 = ~n33683 & n11519;
  assign n11521 = ~n11229 & n11518;
  assign n11522 = n10919 & ~n33762;
  assign n11523 = n10923 & n11519;
  assign n11524 = n10919 & ~n33683;
  assign n11525 = ~n10911 & n11524;
  assign n11526 = ~n11229 & n11525;
  assign n11527 = ~n10919 & ~n33762;
  assign n11528 = ~n11526 & ~n11527;
  assign n11529 = ~n11522 & ~n11523;
  assign n11530 = ~n11517 & ~n33763;
  assign n11531 = ~n11515 & ~n11530;
  assign n11532 = ~n2855 & ~n11531;
  assign n11533 = n2855 & ~n11515;
  assign n11534 = ~n11530 & n11533;
  assign n11535 = n2855 & n11531;
  assign n11536 = ~n10925 & ~n10927;
  assign n11537 = ~n11229 & n11536;
  assign n11538 = ~n33686 & n11537;
  assign n11539 = n33686 & ~n11537;
  assign n11540 = ~n10925 & n33686;
  assign n11541 = ~n10927 & n11540;
  assign n11542 = n33686 & n11537;
  assign n11543 = ~n11229 & n11541;
  assign n11544 = ~n33686 & ~n11537;
  assign n11545 = ~n33765 & ~n11544;
  assign n11546 = ~n11538 & ~n11539;
  assign n11547 = ~n33764 & ~n33766;
  assign n11548 = ~n11532 & ~n11547;
  assign n11549 = ~n2556 & ~n11548;
  assign n11550 = n2556 & ~n11532;
  assign n11551 = ~n11547 & n11550;
  assign n11552 = ~n10943 & ~n33688;
  assign n11553 = ~n10943 & ~n11229;
  assign n11554 = ~n33688 & n11553;
  assign n11555 = ~n11229 & n11552;
  assign n11556 = n10951 & ~n33767;
  assign n11557 = n10955 & n11553;
  assign n11558 = n10951 & ~n33688;
  assign n11559 = ~n10943 & n11558;
  assign n11560 = ~n11229 & n11559;
  assign n11561 = ~n10951 & ~n33767;
  assign n11562 = ~n11560 & ~n11561;
  assign n11563 = ~n11556 & ~n11557;
  assign n11564 = ~n11551 & ~n33768;
  assign n11565 = ~n11549 & ~n11564;
  assign n11566 = ~n2301 & ~n11565;
  assign n11567 = n2301 & ~n11549;
  assign n11568 = ~n11564 & n11567;
  assign n11569 = n2301 & n11565;
  assign n11570 = ~n10957 & ~n10959;
  assign n11571 = ~n10957 & ~n11229;
  assign n11572 = ~n10959 & n11571;
  assign n11573 = ~n11229 & n11570;
  assign n11574 = n33690 & ~n33770;
  assign n11575 = n10971 & n11571;
  assign n11576 = ~n33690 & n33770;
  assign n11577 = ~n10957 & n33690;
  assign n11578 = ~n10959 & n11577;
  assign n11579 = ~n11229 & n11578;
  assign n11580 = ~n33690 & ~n33770;
  assign n11581 = ~n11579 & ~n11580;
  assign n11582 = ~n11574 & ~n33771;
  assign n11583 = ~n33769 & ~n33772;
  assign n11584 = ~n11566 & ~n11583;
  assign n11585 = ~n2038 & ~n11584;
  assign n11586 = n2038 & ~n11566;
  assign n11587 = ~n11583 & n11586;
  assign n11588 = ~n10973 & ~n33692;
  assign n11589 = ~n10973 & ~n11229;
  assign n11590 = ~n33692 & n11589;
  assign n11591 = ~n11229 & n11588;
  assign n11592 = n10981 & ~n33773;
  assign n11593 = n10985 & n11589;
  assign n11594 = n10981 & ~n33692;
  assign n11595 = ~n10973 & n11594;
  assign n11596 = ~n11229 & n11595;
  assign n11597 = ~n10981 & ~n33773;
  assign n11598 = ~n11596 & ~n11597;
  assign n11599 = ~n11592 & ~n11593;
  assign n11600 = ~n11587 & ~n33774;
  assign n11601 = ~n11585 & ~n11600;
  assign n11602 = ~n1812 & ~n11601;
  assign n11603 = ~n10987 & ~n10989;
  assign n11604 = ~n11229 & n11603;
  assign n11605 = ~n33695 & ~n11604;
  assign n11606 = ~n10987 & n33695;
  assign n11607 = ~n10989 & n11606;
  assign n11608 = n33695 & n11604;
  assign n11609 = ~n11229 & n11607;
  assign n11610 = ~n11605 & ~n33775;
  assign n11611 = n1812 & ~n11585;
  assign n11612 = ~n11600 & n11611;
  assign n11613 = n1812 & n11601;
  assign n11614 = ~n11610 & ~n33776;
  assign n11615 = ~n11602 & ~n11614;
  assign n11616 = ~n1582 & ~n11615;
  assign n11617 = n1582 & ~n11602;
  assign n11618 = ~n11614 & n11617;
  assign n11619 = ~n11005 & ~n33697;
  assign n11620 = ~n11005 & ~n11229;
  assign n11621 = ~n33697 & n11620;
  assign n11622 = ~n11229 & n11619;
  assign n11623 = n11013 & ~n33777;
  assign n11624 = n11017 & n11620;
  assign n11625 = n11013 & ~n33697;
  assign n11626 = ~n11005 & n11625;
  assign n11627 = ~n11229 & n11626;
  assign n11628 = ~n11013 & ~n33777;
  assign n11629 = ~n11627 & ~n11628;
  assign n11630 = ~n11623 & ~n11624;
  assign n11631 = ~n11618 & ~n33778;
  assign n11632 = ~n11616 & ~n11631;
  assign n11633 = ~n1388 & ~n11632;
  assign n11634 = n1388 & ~n11616;
  assign n11635 = ~n11631 & n11634;
  assign n11636 = n1388 & n11632;
  assign n11637 = ~n11019 & ~n11029;
  assign n11638 = ~n11019 & ~n11229;
  assign n11639 = ~n11029 & n11638;
  assign n11640 = ~n11229 & n11637;
  assign n11641 = n11027 & ~n33780;
  assign n11642 = n11030 & n11638;
  assign n11643 = ~n11019 & n11027;
  assign n11644 = ~n11029 & n11643;
  assign n11645 = ~n11229 & n11644;
  assign n11646 = ~n11027 & ~n33780;
  assign n11647 = ~n11645 & ~n11646;
  assign n11648 = ~n11641 & ~n11642;
  assign n11649 = ~n33779 & ~n33781;
  assign n11650 = ~n11633 & ~n11649;
  assign n11651 = ~n1192 & ~n11650;
  assign n11652 = n1192 & ~n11633;
  assign n11653 = ~n11649 & n11652;
  assign n11654 = ~n11032 & ~n33700;
  assign n11655 = ~n11032 & ~n11229;
  assign n11656 = ~n33700 & n11655;
  assign n11657 = ~n11229 & n11654;
  assign n11658 = n11040 & ~n33782;
  assign n11659 = n11044 & n11655;
  assign n11660 = n11040 & ~n33700;
  assign n11661 = ~n11032 & n11660;
  assign n11662 = ~n11229 & n11661;
  assign n11663 = ~n11040 & ~n33782;
  assign n11664 = ~n11662 & ~n11663;
  assign n11665 = ~n11658 & ~n11659;
  assign n11666 = ~n11653 & ~n33783;
  assign n11667 = ~n11651 & ~n11666;
  assign n11668 = ~n1028 & ~n11667;
  assign n11669 = ~n11046 & ~n11048;
  assign n11670 = ~n11229 & n11669;
  assign n11671 = ~n33702 & ~n11670;
  assign n11672 = ~n11046 & n33702;
  assign n11673 = ~n11048 & n11672;
  assign n11674 = n33702 & n11670;
  assign n11675 = ~n11229 & n11673;
  assign n11676 = ~n11671 & ~n33784;
  assign n11677 = n1028 & ~n11651;
  assign n11678 = ~n11666 & n11677;
  assign n11679 = n1028 & n11667;
  assign n11680 = ~n11676 & ~n33785;
  assign n11681 = ~n11668 & ~n11680;
  assign n11682 = ~n866 & ~n11681;
  assign n11683 = n866 & ~n11668;
  assign n11684 = ~n11680 & n11683;
  assign n11685 = ~n11063 & ~n33704;
  assign n11686 = ~n11063 & ~n11229;
  assign n11687 = ~n33704 & n11686;
  assign n11688 = ~n11229 & n11685;
  assign n11689 = n11071 & ~n33786;
  assign n11690 = n11075 & n11686;
  assign n11691 = n11071 & ~n33704;
  assign n11692 = ~n11063 & n11691;
  assign n11693 = ~n11229 & n11692;
  assign n11694 = ~n11071 & ~n33786;
  assign n11695 = ~n11693 & ~n11694;
  assign n11696 = ~n11689 & ~n11690;
  assign n11697 = ~n11684 & ~n33787;
  assign n11698 = ~n11682 & ~n11697;
  assign n11699 = ~n730 & ~n11698;
  assign n11700 = n730 & ~n11682;
  assign n11701 = ~n11697 & n11700;
  assign n11702 = n730 & n11698;
  assign n11703 = ~n11077 & ~n11087;
  assign n11704 = ~n11077 & ~n11229;
  assign n11705 = ~n11087 & n11704;
  assign n11706 = ~n11229 & n11703;
  assign n11707 = n11085 & ~n33789;
  assign n11708 = n11088 & n11704;
  assign n11709 = ~n11077 & n11085;
  assign n11710 = ~n11087 & n11709;
  assign n11711 = ~n11229 & n11710;
  assign n11712 = ~n11085 & ~n33789;
  assign n11713 = ~n11711 & ~n11712;
  assign n11714 = ~n11707 & ~n11708;
  assign n11715 = ~n33788 & ~n33790;
  assign n11716 = ~n11699 & ~n11715;
  assign n11717 = ~n602 & ~n11716;
  assign n11718 = n602 & ~n11699;
  assign n11719 = ~n11715 & n11718;
  assign n11720 = ~n11090 & ~n33707;
  assign n11721 = ~n11090 & ~n11229;
  assign n11722 = ~n33707 & n11721;
  assign n11723 = ~n11229 & n11720;
  assign n11724 = n11098 & ~n33791;
  assign n11725 = n11102 & n11721;
  assign n11726 = n11098 & ~n33707;
  assign n11727 = ~n11090 & n11726;
  assign n11728 = ~n11229 & n11727;
  assign n11729 = ~n11098 & ~n33791;
  assign n11730 = ~n11728 & ~n11729;
  assign n11731 = ~n11724 & ~n11725;
  assign n11732 = ~n11719 & ~n33792;
  assign n11733 = ~n11717 & ~n11732;
  assign n11734 = ~n497 & ~n11733;
  assign n11735 = ~n11104 & ~n11106;
  assign n11736 = ~n11229 & n11735;
  assign n11737 = ~n33709 & ~n11736;
  assign n11738 = ~n11104 & n33709;
  assign n11739 = ~n11106 & n11738;
  assign n11740 = n33709 & n11736;
  assign n11741 = ~n11229 & n11739;
  assign n11742 = ~n11737 & ~n33793;
  assign n11743 = n497 & ~n11717;
  assign n11744 = ~n11732 & n11743;
  assign n11745 = n497 & n11733;
  assign n11746 = ~n11742 & ~n33794;
  assign n11747 = ~n11734 & ~n11746;
  assign n11748 = ~n403 & ~n11747;
  assign n11749 = n403 & ~n11734;
  assign n11750 = ~n11746 & n11749;
  assign n11751 = ~n11121 & ~n33711;
  assign n11752 = ~n11121 & ~n11229;
  assign n11753 = ~n33711 & n11752;
  assign n11754 = ~n11229 & n11751;
  assign n11755 = n11129 & ~n33795;
  assign n11756 = n11133 & n11752;
  assign n11757 = n11129 & ~n33711;
  assign n11758 = ~n11121 & n11757;
  assign n11759 = ~n11229 & n11758;
  assign n11760 = ~n11129 & ~n33795;
  assign n11761 = ~n11759 & ~n11760;
  assign n11762 = ~n11755 & ~n11756;
  assign n11763 = ~n11750 & ~n33796;
  assign n11764 = ~n11748 & ~n11763;
  assign n11765 = ~n330 & ~n11764;
  assign n11766 = n330 & ~n11748;
  assign n11767 = ~n11763 & n11766;
  assign n11768 = n330 & n11764;
  assign n11769 = ~n11135 & ~n11145;
  assign n11770 = ~n11135 & ~n11229;
  assign n11771 = ~n11145 & n11770;
  assign n11772 = ~n11229 & n11769;
  assign n11773 = n11143 & ~n33798;
  assign n11774 = n11146 & n11770;
  assign n11775 = ~n11135 & n11143;
  assign n11776 = ~n11145 & n11775;
  assign n11777 = ~n11229 & n11776;
  assign n11778 = ~n11143 & ~n33798;
  assign n11779 = ~n11777 & ~n11778;
  assign n11780 = ~n11773 & ~n11774;
  assign n11781 = ~n33797 & ~n33799;
  assign n11782 = ~n11765 & ~n11781;
  assign n11783 = ~n271 & ~n11782;
  assign n11784 = n271 & ~n11765;
  assign n11785 = ~n11781 & n11784;
  assign n11786 = ~n11148 & ~n33714;
  assign n11787 = ~n11148 & ~n11229;
  assign n11788 = ~n33714 & n11787;
  assign n11789 = ~n11229 & n11786;
  assign n11790 = n11156 & ~n33800;
  assign n11791 = n11160 & n11787;
  assign n11792 = n11156 & ~n33714;
  assign n11793 = ~n11148 & n11792;
  assign n11794 = ~n11229 & n11793;
  assign n11795 = ~n11156 & ~n33800;
  assign n11796 = ~n11794 & ~n11795;
  assign n11797 = ~n11790 & ~n11791;
  assign n11798 = ~n11785 & ~n33801;
  assign n11799 = ~n11783 & ~n11798;
  assign n11800 = ~n217 & ~n11799;
  assign n11801 = ~n11162 & ~n11164;
  assign n11802 = ~n11229 & n11801;
  assign n11803 = ~n33716 & ~n11802;
  assign n11804 = ~n11162 & n33716;
  assign n11805 = ~n11164 & n11804;
  assign n11806 = n33716 & n11802;
  assign n11807 = ~n11229 & n11805;
  assign n11808 = ~n11803 & ~n33802;
  assign n11809 = n217 & ~n11783;
  assign n11810 = ~n11798 & n11809;
  assign n11811 = n217 & n11799;
  assign n11812 = ~n11808 & ~n33803;
  assign n11813 = ~n11800 & ~n11812;
  assign n11814 = ~n198 & ~n11813;
  assign n11815 = n198 & ~n11800;
  assign n11816 = ~n11812 & n11815;
  assign n11817 = ~n11179 & ~n33718;
  assign n11818 = ~n11179 & ~n11229;
  assign n11819 = ~n33718 & n11818;
  assign n11820 = ~n11229 & n11817;
  assign n11821 = n11187 & ~n33804;
  assign n11822 = n11191 & n11818;
  assign n11823 = n11187 & ~n33718;
  assign n11824 = ~n11179 & n11823;
  assign n11825 = ~n11229 & n11824;
  assign n11826 = ~n11187 & ~n33804;
  assign n11827 = ~n11825 & ~n11826;
  assign n11828 = ~n11821 & ~n11822;
  assign n11829 = ~n11816 & ~n33805;
  assign n11830 = ~n11814 & ~n11829;
  assign n11831 = ~n11193 & ~n11203;
  assign n11832 = ~n11193 & ~n11229;
  assign n11833 = ~n11203 & n11832;
  assign n11834 = ~n11229 & n11831;
  assign n11835 = n11201 & ~n33806;
  assign n11836 = n11204 & n11832;
  assign n11837 = ~n11193 & n11201;
  assign n11838 = ~n11203 & n11837;
  assign n11839 = ~n11229 & n11838;
  assign n11840 = ~n11201 & ~n33806;
  assign n11841 = ~n11839 & ~n11840;
  assign n11842 = ~n11835 & ~n11836;
  assign n11843 = ~n11205 & ~n11213;
  assign n11844 = ~n11213 & ~n11229;
  assign n11845 = ~n11205 & n11844;
  assign n11846 = ~n11229 & n11843;
  assign n11847 = ~n33722 & ~n33808;
  assign n11848 = ~n33807 & n11847;
  assign n11849 = ~n11830 & n11848;
  assign n11850 = n193 & ~n11849;
  assign n11851 = ~n11814 & n33807;
  assign n11852 = ~n11829 & n11851;
  assign n11853 = n11830 & n33807;
  assign n11854 = n11205 & ~n11844;
  assign n11855 = ~n193 & ~n11843;
  assign n11856 = ~n11854 & n11855;
  assign n11857 = ~n33809 & ~n11856;
  assign n11858 = ~n11850 & n11857;
  assign n11859 = ~n11426 & ~n11428;
  assign n11860 = ~n11858 & n11859;
  assign n11861 = ~n33724 & ~n11860;
  assign n11862 = n33724 & ~n11428;
  assign n11863 = ~n11426 & n11862;
  assign n11864 = n33724 & n11860;
  assign n11865 = ~n11858 & n11863;
  assign n11866 = ~n11861 & ~n33810;
  assign n11867 = ~n11360 & ~n11362;
  assign n11868 = ~n11858 & n11867;
  assign n11869 = ~n33741 & ~n11868;
  assign n11870 = ~n11362 & n33741;
  assign n11871 = ~n11360 & n11870;
  assign n11872 = n33741 & n11868;
  assign n11873 = ~n11858 & n11871;
  assign n11874 = ~n11869 & ~n33811;
  assign n11875 = ~n11327 & ~n11329;
  assign n11876 = ~n11858 & n11875;
  assign n11877 = ~n33737 & ~n11876;
  assign n11878 = ~n11329 & n33737;
  assign n11879 = ~n11327 & n11878;
  assign n11880 = n33737 & n11876;
  assign n11881 = ~n11858 & n11879;
  assign n11882 = ~n11877 & ~n33812;
  assign n11883 = ~n11293 & ~n11295;
  assign n11884 = ~n11858 & n11883;
  assign n11885 = ~n33732 & ~n11884;
  assign n11886 = ~n11295 & n33732;
  assign n11887 = ~n11293 & n11886;
  assign n11888 = n33732 & n11884;
  assign n11889 = ~n11858 & n11887;
  assign n11890 = ~n11885 & ~n33813;
  assign n11891 = ~n11266 & ~n11268;
  assign n11892 = ~n11858 & n11891;
  assign n11893 = ~n11277 & ~n11892;
  assign n11894 = ~n11268 & n11277;
  assign n11895 = ~n11266 & n11894;
  assign n11896 = n11277 & n11892;
  assign n11897 = ~n11858 & n11895;
  assign n11898 = ~n11893 & ~n33814;
  assign n11899 = ~pi50  & ~n11858;
  assign n11900 = ~pi51  & n11899;
  assign n11901 = n11243 & ~n11858;
  assign n11902 = ~n11229 & ~n11856;
  assign n11903 = ~n33809 & n11902;
  assign n11904 = ~n11850 & n11903;
  assign n11905 = ~n33815 & ~n11904;
  assign n11906 = pi52  & ~n11905;
  assign n11907 = ~pi52  & ~n11904;
  assign n11908 = ~pi52  & n11905;
  assign n11909 = ~n33815 & n11907;
  assign n11910 = ~n11906 & ~n33816;
  assign n11911 = pi50  & ~n11858;
  assign n11912 = ~pi48  & ~pi49 ;
  assign n11913 = ~pi50  & n11912;
  assign n11914 = ~n33650 & ~n33726;
  assign n11915 = ~n10660 & n11914;
  assign n11916 = ~n10679 & n11915;
  assign n11917 = ~n33652 & n11916;
  assign n11918 = n10665 & n10681;
  assign n11919 = ~n10673 & n11917;
  assign n11920 = ~n11913 & ~n33817;
  assign n11921 = ~n11227 & n11920;
  assign n11922 = ~n33722 & n11921;
  assign n11923 = ~n11221 & n11922;
  assign n11924 = ~n11911 & ~n11913;
  assign n11925 = n11229 & n11924;
  assign n11926 = ~n11911 & n11923;
  assign n11927 = pi51  & ~n11899;
  assign n11928 = ~n33815 & ~n11927;
  assign n11929 = ~n33818 & n11928;
  assign n11930 = ~n11229 & ~n11924;
  assign n11931 = n10681 & ~n11930;
  assign n11932 = ~n11929 & ~n11930;
  assign n11933 = n10681 & n11932;
  assign n11934 = ~n11929 & n11931;
  assign n11935 = ~n11910 & ~n33819;
  assign n11936 = ~n10681 & ~n11932;
  assign n11937 = n10086 & ~n11936;
  assign n11938 = ~n11935 & n11937;
  assign n11939 = ~n11246 & ~n33727;
  assign n11940 = ~n11858 & n11939;
  assign n11941 = n11251 & ~n11940;
  assign n11942 = ~n11251 & n11939;
  assign n11943 = ~n11251 & n11940;
  assign n11944 = ~n11858 & n11942;
  assign n11945 = ~n11941 & ~n33820;
  assign n11946 = ~n11938 & ~n11945;
  assign n11947 = ~n11935 & ~n11936;
  assign n11948 = ~n10086 & ~n11947;
  assign n11949 = n9565 & ~n11948;
  assign n11950 = ~n11946 & ~n11948;
  assign n11951 = n9565 & n11950;
  assign n11952 = ~n11946 & n11949;
  assign n11953 = ~n11898 & ~n33821;
  assign n11954 = ~n9565 & ~n11950;
  assign n11955 = n8998 & ~n11954;
  assign n11956 = ~n11953 & n11955;
  assign n11957 = ~n11280 & ~n33729;
  assign n11958 = ~n11858 & n11957;
  assign n11959 = n11290 & ~n11958;
  assign n11960 = ~n11290 & n11958;
  assign n11961 = ~n11280 & n11290;
  assign n11962 = ~n33729 & n11961;
  assign n11963 = n11290 & n11958;
  assign n11964 = ~n11858 & n11962;
  assign n11965 = ~n11290 & ~n11958;
  assign n11966 = ~n33822 & ~n11965;
  assign n11967 = ~n11959 & ~n11960;
  assign n11968 = ~n11956 & ~n33823;
  assign n11969 = ~n11953 & ~n11954;
  assign n11970 = ~n8998 & ~n11969;
  assign n11971 = n8506 & ~n11970;
  assign n11972 = ~n11968 & ~n11970;
  assign n11973 = n8506 & n11972;
  assign n11974 = ~n11968 & n11971;
  assign n11975 = ~n11890 & ~n33824;
  assign n11976 = ~n8506 & ~n11972;
  assign n11977 = n7975 & ~n11976;
  assign n11978 = ~n11975 & n11977;
  assign n11979 = ~n11310 & ~n33733;
  assign n11980 = ~n11858 & n11979;
  assign n11981 = ~n33735 & n11980;
  assign n11982 = n33735 & ~n11980;
  assign n11983 = ~n11310 & n33735;
  assign n11984 = ~n33733 & n11983;
  assign n11985 = ~n11858 & n11984;
  assign n11986 = ~n33735 & ~n11980;
  assign n11987 = ~n11985 & ~n11986;
  assign n11988 = ~n11981 & ~n11982;
  assign n11989 = ~n11978 & ~n33825;
  assign n11990 = ~n11975 & ~n11976;
  assign n11991 = ~n7975 & ~n11990;
  assign n11992 = n7512 & ~n11991;
  assign n11993 = ~n11989 & ~n11991;
  assign n11994 = n7512 & n11993;
  assign n11995 = ~n11989 & n11992;
  assign n11996 = ~n11882 & ~n33826;
  assign n11997 = ~n7512 & ~n11993;
  assign n11998 = n7015 & ~n11997;
  assign n11999 = ~n11996 & n11998;
  assign n12000 = ~n11344 & ~n33738;
  assign n12001 = ~n11858 & n12000;
  assign n12002 = ~n33739 & ~n12001;
  assign n12003 = ~n11344 & n33739;
  assign n12004 = ~n33738 & n12003;
  assign n12005 = n33739 & n12001;
  assign n12006 = ~n11858 & n12004;
  assign n12007 = n33739 & ~n12001;
  assign n12008 = ~n33739 & n12001;
  assign n12009 = ~n12007 & ~n12008;
  assign n12010 = ~n12002 & ~n33827;
  assign n12011 = ~n11999 & n33828;
  assign n12012 = ~n11996 & ~n11997;
  assign n12013 = ~n7015 & ~n12012;
  assign n12014 = n6579 & ~n12013;
  assign n12015 = ~n12011 & ~n12013;
  assign n12016 = n6579 & n12015;
  assign n12017 = ~n12011 & n12014;
  assign n12018 = ~n11874 & ~n33829;
  assign n12019 = ~n6579 & ~n12015;
  assign n12020 = n6117 & ~n12019;
  assign n12021 = ~n12018 & n12020;
  assign n12022 = ~n11377 & ~n33742;
  assign n12023 = ~n11858 & n12022;
  assign n12024 = n33744 & ~n12023;
  assign n12025 = ~n11377 & ~n33744;
  assign n12026 = ~n33742 & n12025;
  assign n12027 = ~n33744 & n12023;
  assign n12028 = ~n11858 & n12026;
  assign n12029 = n33744 & n12023;
  assign n12030 = ~n33744 & ~n12023;
  assign n12031 = ~n12029 & ~n12030;
  assign n12032 = ~n12024 & ~n33830;
  assign n12033 = ~n12021 & n33831;
  assign n12034 = ~n12018 & ~n12019;
  assign n12035 = ~n6117 & ~n12034;
  assign n12036 = n5708 & ~n12035;
  assign n12037 = ~n12033 & ~n12035;
  assign n12038 = n5708 & n12037;
  assign n12039 = ~n12033 & n12036;
  assign n12040 = ~n11394 & ~n11396;
  assign n12041 = ~n11858 & n12040;
  assign n12042 = ~n33745 & n12041;
  assign n12043 = n33745 & ~n12041;
  assign n12044 = ~n11396 & n33745;
  assign n12045 = ~n11394 & n12044;
  assign n12046 = ~n11858 & n12045;
  assign n12047 = ~n33745 & ~n12041;
  assign n12048 = ~n12046 & ~n12047;
  assign n12049 = ~n12042 & ~n12043;
  assign n12050 = ~n33832 & ~n33833;
  assign n12051 = ~n5708 & ~n12037;
  assign n12052 = ~n12050 & ~n12051;
  assign n12053 = ~n5278 & ~n12052;
  assign n12054 = n5278 & ~n12051;
  assign n12055 = ~n12050 & n12054;
  assign n12056 = ~n11409 & ~n33748;
  assign n12057 = ~n11858 & n12056;
  assign n12058 = ~n33747 & ~n12057;
  assign n12059 = n33747 & n12057;
  assign n12060 = ~n11409 & ~n33747;
  assign n12061 = ~n33748 & n12060;
  assign n12062 = ~n11858 & n12061;
  assign n12063 = n33747 & ~n12057;
  assign n12064 = ~n12062 & ~n12063;
  assign n12065 = ~n12058 & ~n12059;
  assign n12066 = ~n12055 & ~n33834;
  assign n12067 = ~n12053 & ~n12066;
  assign n12068 = ~n4903 & ~n12067;
  assign n12069 = n4903 & ~n12053;
  assign n12070 = n4903 & n12067;
  assign n12071 = ~n12066 & n12069;
  assign n12072 = ~n11866 & ~n33835;
  assign n12073 = ~n12068 & ~n12072;
  assign n12074 = ~n4508 & ~n12073;
  assign n12075 = n4508 & ~n12068;
  assign n12076 = ~n12072 & n12075;
  assign n12077 = ~n11431 & ~n33749;
  assign n12078 = ~n11431 & ~n11858;
  assign n12079 = ~n33749 & n12078;
  assign n12080 = ~n11858 & n12077;
  assign n12081 = n11446 & n12078;
  assign n12082 = ~n33751 & n33836;
  assign n12083 = n33751 & ~n33836;
  assign n12084 = ~n11431 & n33751;
  assign n12085 = ~n33749 & n12084;
  assign n12086 = n33751 & n33836;
  assign n12087 = ~n11858 & n12085;
  assign n12088 = ~n33751 & ~n33836;
  assign n12089 = ~n33838 & ~n12088;
  assign n12090 = ~n33837 & ~n12083;
  assign n12091 = ~n12076 & ~n33839;
  assign n12092 = ~n12074 & ~n12091;
  assign n12093 = ~n4155 & ~n12092;
  assign n12094 = ~n11448 & ~n11450;
  assign n12095 = ~n11858 & n12094;
  assign n12096 = ~n33753 & ~n12095;
  assign n12097 = ~n11450 & n33753;
  assign n12098 = ~n11448 & n12097;
  assign n12099 = n33753 & n12095;
  assign n12100 = ~n11858 & n12098;
  assign n12101 = ~n12096 & ~n33840;
  assign n12102 = n4155 & ~n12074;
  assign n12103 = n4155 & n12092;
  assign n12104 = ~n12091 & n12102;
  assign n12105 = ~n12101 & ~n33841;
  assign n12106 = ~n12093 & ~n12105;
  assign n12107 = ~n3788 & ~n12106;
  assign n12108 = n3788 & ~n12093;
  assign n12109 = ~n12105 & n12108;
  assign n12110 = ~n11465 & ~n33754;
  assign n12111 = ~n11465 & ~n11858;
  assign n12112 = ~n33754 & n12111;
  assign n12113 = ~n11858 & n12110;
  assign n12114 = n11476 & ~n33842;
  assign n12115 = n11477 & n12111;
  assign n12116 = ~n11476 & n33842;
  assign n12117 = ~n11465 & n11476;
  assign n12118 = ~n33754 & n12117;
  assign n12119 = ~n11858 & n12118;
  assign n12120 = ~n11476 & ~n33842;
  assign n12121 = ~n12119 & ~n12120;
  assign n12122 = ~n12114 & ~n33843;
  assign n12123 = ~n12109 & ~n33844;
  assign n12124 = ~n12107 & ~n12123;
  assign n12125 = ~n3473 & ~n12124;
  assign n12126 = ~n11479 & ~n11481;
  assign n12127 = ~n11858 & n12126;
  assign n12128 = ~n33757 & ~n12127;
  assign n12129 = ~n11481 & n33757;
  assign n12130 = ~n11479 & n12129;
  assign n12131 = n33757 & n12127;
  assign n12132 = ~n11858 & n12130;
  assign n12133 = ~n12128 & ~n33845;
  assign n12134 = n3473 & ~n12107;
  assign n12135 = n3473 & n12124;
  assign n12136 = ~n12123 & n12134;
  assign n12137 = ~n12133 & ~n33846;
  assign n12138 = ~n12125 & ~n12137;
  assign n12139 = ~n3140 & ~n12138;
  assign n12140 = n3140 & ~n12125;
  assign n12141 = ~n12137 & n12140;
  assign n12142 = ~n11496 & ~n33758;
  assign n12143 = ~n11858 & n12142;
  assign n12144 = ~n33761 & n12143;
  assign n12145 = n33761 & ~n12143;
  assign n12146 = ~n11496 & n33761;
  assign n12147 = ~n33758 & n12146;
  assign n12148 = n33761 & n12143;
  assign n12149 = ~n11858 & n12147;
  assign n12150 = ~n33761 & ~n12143;
  assign n12151 = ~n33847 & ~n12150;
  assign n12152 = ~n12144 & ~n12145;
  assign n12153 = ~n12141 & ~n33848;
  assign n12154 = ~n12139 & ~n12153;
  assign n12155 = ~n2855 & ~n12154;
  assign n12156 = ~n11515 & ~n11517;
  assign n12157 = ~n11858 & n12156;
  assign n12158 = ~n33763 & ~n12157;
  assign n12159 = ~n11517 & n33763;
  assign n12160 = ~n11515 & n12159;
  assign n12161 = n33763 & n12157;
  assign n12162 = ~n11858 & n12160;
  assign n12163 = ~n12158 & ~n33849;
  assign n12164 = n2855 & ~n12139;
  assign n12165 = n2855 & n12154;
  assign n12166 = ~n12153 & n12164;
  assign n12167 = ~n12163 & ~n33850;
  assign n12168 = ~n12155 & ~n12167;
  assign n12169 = ~n2556 & ~n12168;
  assign n12170 = n2556 & ~n12155;
  assign n12171 = ~n12167 & n12170;
  assign n12172 = ~n11532 & ~n33764;
  assign n12173 = ~n11532 & ~n11858;
  assign n12174 = ~n33764 & n12173;
  assign n12175 = ~n11858 & n12172;
  assign n12176 = n33766 & ~n33851;
  assign n12177 = n11547 & n12173;
  assign n12178 = ~n33766 & n33851;
  assign n12179 = ~n11532 & n33766;
  assign n12180 = ~n33764 & n12179;
  assign n12181 = ~n11858 & n12180;
  assign n12182 = ~n33766 & ~n33851;
  assign n12183 = ~n12181 & ~n12182;
  assign n12184 = ~n12176 & ~n33852;
  assign n12185 = ~n12171 & ~n33853;
  assign n12186 = ~n12169 & ~n12185;
  assign n12187 = ~n2301 & ~n12186;
  assign n12188 = ~n11549 & ~n11551;
  assign n12189 = ~n11858 & n12188;
  assign n12190 = ~n33768 & ~n12189;
  assign n12191 = ~n11551 & n33768;
  assign n12192 = ~n11549 & n12191;
  assign n12193 = n33768 & n12189;
  assign n12194 = ~n11858 & n12192;
  assign n12195 = ~n12190 & ~n33854;
  assign n12196 = n2301 & ~n12169;
  assign n12197 = n2301 & n12186;
  assign n12198 = ~n12185 & n12196;
  assign n12199 = ~n12195 & ~n33855;
  assign n12200 = ~n12187 & ~n12199;
  assign n12201 = ~n2038 & ~n12200;
  assign n12202 = ~n11566 & ~n33769;
  assign n12203 = ~n11858 & n12202;
  assign n12204 = ~n33772 & ~n12203;
  assign n12205 = ~n11566 & n33772;
  assign n12206 = ~n33769 & n12205;
  assign n12207 = n33772 & n12203;
  assign n12208 = ~n11858 & n12206;
  assign n12209 = ~n12204 & ~n33856;
  assign n12210 = n2038 & ~n12187;
  assign n12211 = ~n12199 & n12210;
  assign n12212 = ~n12209 & ~n12211;
  assign n12213 = ~n12201 & ~n12212;
  assign n12214 = ~n1812 & ~n12213;
  assign n12215 = ~n11585 & ~n11587;
  assign n12216 = ~n11858 & n12215;
  assign n12217 = ~n33774 & ~n12216;
  assign n12218 = ~n11587 & n33774;
  assign n12219 = ~n11585 & n12218;
  assign n12220 = n33774 & n12216;
  assign n12221 = ~n11858 & n12219;
  assign n12222 = ~n12217 & ~n33857;
  assign n12223 = n1812 & ~n12201;
  assign n12224 = n1812 & n12213;
  assign n12225 = ~n12212 & n12223;
  assign n12226 = ~n12222 & ~n33858;
  assign n12227 = ~n12214 & ~n12226;
  assign n12228 = ~n1582 & ~n12227;
  assign n12229 = n1582 & ~n12214;
  assign n12230 = ~n12226 & n12229;
  assign n12231 = ~n11602 & ~n33776;
  assign n12232 = ~n11602 & ~n11858;
  assign n12233 = ~n33776 & n12232;
  assign n12234 = ~n11858 & n12231;
  assign n12235 = n11610 & ~n33859;
  assign n12236 = n11614 & n12232;
  assign n12237 = ~n11602 & n11610;
  assign n12238 = ~n33776 & n12237;
  assign n12239 = ~n11858 & n12238;
  assign n12240 = ~n11610 & ~n33859;
  assign n12241 = ~n12239 & ~n12240;
  assign n12242 = ~n12235 & ~n12236;
  assign n12243 = ~n12230 & ~n33860;
  assign n12244 = ~n12228 & ~n12243;
  assign n12245 = ~n1388 & ~n12244;
  assign n12246 = ~n11616 & ~n11618;
  assign n12247 = ~n11858 & n12246;
  assign n12248 = ~n33778 & ~n12247;
  assign n12249 = ~n11618 & n33778;
  assign n12250 = ~n11616 & n12249;
  assign n12251 = n33778 & n12247;
  assign n12252 = ~n11858 & n12250;
  assign n12253 = ~n12248 & ~n33861;
  assign n12254 = n1388 & ~n12228;
  assign n12255 = n1388 & n12244;
  assign n12256 = ~n12243 & n12254;
  assign n12257 = ~n12253 & ~n33862;
  assign n12258 = ~n12245 & ~n12257;
  assign n12259 = ~n1192 & ~n12258;
  assign n12260 = ~n11633 & ~n33779;
  assign n12261 = ~n11858 & n12260;
  assign n12262 = ~n33781 & ~n12261;
  assign n12263 = ~n11633 & n33781;
  assign n12264 = ~n33779 & n12263;
  assign n12265 = n33781 & n12261;
  assign n12266 = ~n11858 & n12264;
  assign n12267 = ~n12262 & ~n33863;
  assign n12268 = n1192 & ~n12245;
  assign n12269 = ~n12257 & n12268;
  assign n12270 = ~n12267 & ~n12269;
  assign n12271 = ~n12259 & ~n12270;
  assign n12272 = ~n1028 & ~n12271;
  assign n12273 = ~n11651 & ~n11653;
  assign n12274 = ~n11858 & n12273;
  assign n12275 = ~n33783 & ~n12274;
  assign n12276 = ~n11653 & n33783;
  assign n12277 = ~n11651 & n12276;
  assign n12278 = n33783 & n12274;
  assign n12279 = ~n11858 & n12277;
  assign n12280 = ~n12275 & ~n33864;
  assign n12281 = n1028 & ~n12259;
  assign n12282 = n1028 & n12271;
  assign n12283 = ~n12270 & n12281;
  assign n12284 = ~n12280 & ~n33865;
  assign n12285 = ~n12272 & ~n12284;
  assign n12286 = ~n866 & ~n12285;
  assign n12287 = n866 & ~n12272;
  assign n12288 = ~n12284 & n12287;
  assign n12289 = ~n11668 & ~n33785;
  assign n12290 = ~n11668 & ~n11858;
  assign n12291 = ~n33785 & n12290;
  assign n12292 = ~n11858 & n12289;
  assign n12293 = n11676 & ~n33866;
  assign n12294 = n11680 & n12290;
  assign n12295 = ~n11668 & n11676;
  assign n12296 = ~n33785 & n12295;
  assign n12297 = ~n11858 & n12296;
  assign n12298 = ~n11676 & ~n33866;
  assign n12299 = ~n12297 & ~n12298;
  assign n12300 = ~n12293 & ~n12294;
  assign n12301 = ~n12288 & ~n33867;
  assign n12302 = ~n12286 & ~n12301;
  assign n12303 = ~n730 & ~n12302;
  assign n12304 = ~n11682 & ~n11684;
  assign n12305 = ~n11858 & n12304;
  assign n12306 = ~n33787 & ~n12305;
  assign n12307 = ~n11684 & n33787;
  assign n12308 = ~n11682 & n12307;
  assign n12309 = n33787 & n12305;
  assign n12310 = ~n11858 & n12308;
  assign n12311 = ~n12306 & ~n33868;
  assign n12312 = n730 & ~n12286;
  assign n12313 = n730 & n12302;
  assign n12314 = ~n12301 & n12312;
  assign n12315 = ~n12311 & ~n33869;
  assign n12316 = ~n12303 & ~n12315;
  assign n12317 = ~n602 & ~n12316;
  assign n12318 = ~n11699 & ~n33788;
  assign n12319 = ~n11858 & n12318;
  assign n12320 = ~n33790 & ~n12319;
  assign n12321 = ~n11699 & n33790;
  assign n12322 = ~n33788 & n12321;
  assign n12323 = n33790 & n12319;
  assign n12324 = ~n11858 & n12322;
  assign n12325 = ~n12320 & ~n33870;
  assign n12326 = n602 & ~n12303;
  assign n12327 = ~n12315 & n12326;
  assign n12328 = ~n12325 & ~n12327;
  assign n12329 = ~n12317 & ~n12328;
  assign n12330 = ~n497 & ~n12329;
  assign n12331 = ~n11717 & ~n11719;
  assign n12332 = ~n11858 & n12331;
  assign n12333 = ~n33792 & ~n12332;
  assign n12334 = ~n11719 & n33792;
  assign n12335 = ~n11717 & n12334;
  assign n12336 = n33792 & n12332;
  assign n12337 = ~n11858 & n12335;
  assign n12338 = ~n12333 & ~n33871;
  assign n12339 = n497 & ~n12317;
  assign n12340 = n497 & n12329;
  assign n12341 = ~n12328 & n12339;
  assign n12342 = ~n12338 & ~n33872;
  assign n12343 = ~n12330 & ~n12342;
  assign n12344 = ~n403 & ~n12343;
  assign n12345 = n403 & ~n12330;
  assign n12346 = ~n12342 & n12345;
  assign n12347 = ~n11734 & ~n33794;
  assign n12348 = ~n11734 & ~n11858;
  assign n12349 = ~n33794 & n12348;
  assign n12350 = ~n11858 & n12347;
  assign n12351 = n11742 & ~n33873;
  assign n12352 = n11746 & n12348;
  assign n12353 = ~n11734 & n11742;
  assign n12354 = ~n33794 & n12353;
  assign n12355 = ~n11858 & n12354;
  assign n12356 = ~n11742 & ~n33873;
  assign n12357 = ~n12355 & ~n12356;
  assign n12358 = ~n12351 & ~n12352;
  assign n12359 = ~n12346 & ~n33874;
  assign n12360 = ~n12344 & ~n12359;
  assign n12361 = ~n330 & ~n12360;
  assign n12362 = ~n11748 & ~n11750;
  assign n12363 = ~n11858 & n12362;
  assign n12364 = ~n33796 & ~n12363;
  assign n12365 = ~n11750 & n33796;
  assign n12366 = ~n11748 & n12365;
  assign n12367 = n33796 & n12363;
  assign n12368 = ~n11858 & n12366;
  assign n12369 = ~n12364 & ~n33875;
  assign n12370 = n330 & ~n12344;
  assign n12371 = n330 & n12360;
  assign n12372 = ~n12359 & n12370;
  assign n12373 = ~n12369 & ~n33876;
  assign n12374 = ~n12361 & ~n12373;
  assign n12375 = ~n271 & ~n12374;
  assign n12376 = ~n11765 & ~n33797;
  assign n12377 = ~n11858 & n12376;
  assign n12378 = ~n33799 & ~n12377;
  assign n12379 = ~n11765 & n33799;
  assign n12380 = ~n33797 & n12379;
  assign n12381 = n33799 & n12377;
  assign n12382 = ~n11858 & n12380;
  assign n12383 = ~n12378 & ~n33877;
  assign n12384 = n271 & ~n12361;
  assign n12385 = ~n12373 & n12384;
  assign n12386 = ~n12383 & ~n12385;
  assign n12387 = ~n12375 & ~n12386;
  assign n12388 = ~n217 & ~n12387;
  assign n12389 = ~n11783 & ~n11785;
  assign n12390 = ~n11858 & n12389;
  assign n12391 = ~n33801 & ~n12390;
  assign n12392 = ~n11785 & n33801;
  assign n12393 = ~n11783 & n12392;
  assign n12394 = n33801 & n12390;
  assign n12395 = ~n11858 & n12393;
  assign n12396 = ~n12391 & ~n33878;
  assign n12397 = n217 & ~n12375;
  assign n12398 = n217 & n12387;
  assign n12399 = ~n12386 & n12397;
  assign n12400 = ~n12396 & ~n33879;
  assign n12401 = ~n12388 & ~n12400;
  assign n12402 = ~n198 & ~n12401;
  assign n12403 = n198 & ~n12388;
  assign n12404 = ~n12400 & n12403;
  assign n12405 = ~n11800 & ~n33803;
  assign n12406 = ~n11800 & ~n11858;
  assign n12407 = ~n33803 & n12406;
  assign n12408 = ~n11858 & n12405;
  assign n12409 = n11808 & ~n33880;
  assign n12410 = n11812 & n12406;
  assign n12411 = ~n11800 & n11808;
  assign n12412 = ~n33803 & n12411;
  assign n12413 = ~n11858 & n12412;
  assign n12414 = ~n11808 & ~n33880;
  assign n12415 = ~n12413 & ~n12414;
  assign n12416 = ~n12409 & ~n12410;
  assign n12417 = ~n12404 & ~n33881;
  assign n12418 = ~n12402 & ~n12417;
  assign n12419 = ~n11814 & ~n11816;
  assign n12420 = ~n11858 & n12419;
  assign n12421 = ~n33805 & ~n12420;
  assign n12422 = ~n11816 & n33805;
  assign n12423 = ~n11814 & n12422;
  assign n12424 = n33805 & n12420;
  assign n12425 = ~n11858 & n12423;
  assign n12426 = ~n12421 & ~n33882;
  assign n12427 = ~n11830 & ~n33807;
  assign n12428 = ~n33807 & ~n11858;
  assign n12429 = ~n11830 & n12428;
  assign n12430 = ~n11858 & n12427;
  assign n12431 = ~n33809 & ~n33883;
  assign n12432 = ~n12426 & n12431;
  assign n12433 = ~n12418 & n12432;
  assign n12434 = n193 & ~n12433;
  assign n12435 = ~n12402 & n12426;
  assign n12436 = n12418 & n12426;
  assign n12437 = ~n12417 & n12435;
  assign n12438 = n11830 & ~n12428;
  assign n12439 = ~n193 & ~n12427;
  assign n12440 = ~n12438 & n12439;
  assign n12441 = ~n33884 & ~n12440;
  assign n12442 = ~n12434 & n12441;
  assign n12443 = ~n12068 & ~n33835;
  assign n12444 = ~n12068 & ~n12442;
  assign n12445 = ~n33835 & n12444;
  assign n12446 = ~n12442 & n12443;
  assign n12447 = n11866 & ~n33885;
  assign n12448 = n12072 & n12444;
  assign n12449 = n11866 & ~n33835;
  assign n12450 = ~n12068 & n12449;
  assign n12451 = ~n12442 & n12450;
  assign n12452 = ~n11866 & ~n33885;
  assign n12453 = ~n12451 & ~n12452;
  assign n12454 = ~n12447 & ~n12448;
  assign n12455 = pi48  & ~n12442;
  assign n12456 = ~pi46  & ~pi47 ;
  assign n12457 = ~pi48  & n12456;
  assign n12458 = ~n12455 & ~n12457;
  assign n12459 = ~n11858 & ~n12458;
  assign n12460 = ~pi48  & ~n12442;
  assign n12461 = pi49  & ~n12460;
  assign n12462 = ~pi49  & n12460;
  assign n12463 = n11912 & ~n12442;
  assign n12464 = ~n12461 & ~n33887;
  assign n12465 = ~n33720 & ~n33817;
  assign n12466 = ~n11208 & n12465;
  assign n12467 = ~n11227 & n12466;
  assign n12468 = ~n33722 & n12467;
  assign n12469 = n11213 & n11229;
  assign n12470 = ~n11221 & n12468;
  assign n12471 = ~n12457 & ~n33888;
  assign n12472 = ~n11856 & n12471;
  assign n12473 = ~n33809 & n12472;
  assign n12474 = ~n11850 & n12473;
  assign n12475 = n11858 & n12458;
  assign n12476 = ~n12455 & n12474;
  assign n12477 = n12464 & ~n33889;
  assign n12478 = ~n12459 & ~n12477;
  assign n12479 = ~n11229 & ~n12478;
  assign n12480 = n11229 & ~n12459;
  assign n12481 = ~n12477 & n12480;
  assign n12482 = ~n11858 & ~n12440;
  assign n12483 = ~n33884 & n12482;
  assign n12484 = ~n12434 & n12483;
  assign n12485 = ~n33887 & ~n12484;
  assign n12486 = pi50  & ~n12485;
  assign n12487 = ~pi50  & ~n12484;
  assign n12488 = ~pi50  & n12485;
  assign n12489 = ~n33887 & n12487;
  assign n12490 = ~n12486 & ~n33890;
  assign n12491 = ~n12481 & ~n12490;
  assign n12492 = ~n12479 & ~n12491;
  assign n12493 = ~n10681 & ~n12492;
  assign n12494 = n10681 & ~n12479;
  assign n12495 = ~n12491 & n12494;
  assign n12496 = n10681 & n12492;
  assign n12497 = ~n33818 & ~n11930;
  assign n12498 = ~n12442 & n12497;
  assign n12499 = n11928 & ~n12498;
  assign n12500 = ~n11928 & n12497;
  assign n12501 = ~n11928 & n12498;
  assign n12502 = ~n12442 & n12500;
  assign n12503 = ~n12499 & ~n33892;
  assign n12504 = ~n33891 & ~n12503;
  assign n12505 = ~n12493 & ~n12504;
  assign n12506 = ~n10086 & ~n12505;
  assign n12507 = n10086 & ~n12493;
  assign n12508 = ~n12504 & n12507;
  assign n12509 = ~n33819 & ~n11936;
  assign n12510 = ~n11936 & ~n12442;
  assign n12511 = ~n33819 & n12510;
  assign n12512 = ~n12442 & n12509;
  assign n12513 = n11910 & ~n33893;
  assign n12514 = n11935 & n12510;
  assign n12515 = n11910 & ~n33819;
  assign n12516 = ~n11936 & n12515;
  assign n12517 = ~n12442 & n12516;
  assign n12518 = ~n11910 & ~n33893;
  assign n12519 = ~n12517 & ~n12518;
  assign n12520 = ~n12513 & ~n12514;
  assign n12521 = ~n12508 & ~n33894;
  assign n12522 = ~n12506 & ~n12521;
  assign n12523 = ~n9565 & ~n12522;
  assign n12524 = n9565 & ~n12506;
  assign n12525 = ~n12521 & n12524;
  assign n12526 = n9565 & n12522;
  assign n12527 = ~n11938 & ~n11948;
  assign n12528 = ~n12442 & n12527;
  assign n12529 = n11945 & ~n12528;
  assign n12530 = ~n11945 & n12528;
  assign n12531 = n11945 & ~n11948;
  assign n12532 = ~n11938 & n12531;
  assign n12533 = n11945 & n12528;
  assign n12534 = ~n12442 & n12532;
  assign n12535 = ~n11945 & ~n12528;
  assign n12536 = ~n33896 & ~n12535;
  assign n12537 = ~n12529 & ~n12530;
  assign n12538 = ~n33895 & ~n33897;
  assign n12539 = ~n12523 & ~n12538;
  assign n12540 = ~n8998 & ~n12539;
  assign n12541 = n8998 & ~n12523;
  assign n12542 = ~n12538 & n12541;
  assign n12543 = ~n33821 & ~n11954;
  assign n12544 = ~n11954 & ~n12442;
  assign n12545 = ~n33821 & n12544;
  assign n12546 = ~n12442 & n12543;
  assign n12547 = n11898 & ~n33898;
  assign n12548 = n11953 & n12544;
  assign n12549 = n11898 & ~n33821;
  assign n12550 = ~n11954 & n12549;
  assign n12551 = ~n12442 & n12550;
  assign n12552 = ~n11898 & ~n33898;
  assign n12553 = ~n12551 & ~n12552;
  assign n12554 = ~n12547 & ~n12548;
  assign n12555 = ~n12542 & ~n33899;
  assign n12556 = ~n12540 & ~n12555;
  assign n12557 = ~n8506 & ~n12556;
  assign n12558 = n8506 & ~n12540;
  assign n12559 = ~n12555 & n12558;
  assign n12560 = n8506 & n12556;
  assign n12561 = ~n11956 & ~n11970;
  assign n12562 = ~n12442 & n12561;
  assign n12563 = ~n33823 & n12562;
  assign n12564 = n33823 & ~n12562;
  assign n12565 = n33823 & ~n11970;
  assign n12566 = ~n11956 & n12565;
  assign n12567 = ~n12442 & n12566;
  assign n12568 = ~n33823 & ~n12562;
  assign n12569 = ~n12567 & ~n12568;
  assign n12570 = ~n12563 & ~n12564;
  assign n12571 = ~n33900 & ~n33901;
  assign n12572 = ~n12557 & ~n12571;
  assign n12573 = ~n7975 & ~n12572;
  assign n12574 = n7975 & ~n12557;
  assign n12575 = ~n12571 & n12574;
  assign n12576 = ~n33824 & ~n11976;
  assign n12577 = ~n11976 & ~n12442;
  assign n12578 = ~n33824 & n12577;
  assign n12579 = ~n12442 & n12576;
  assign n12580 = n11890 & ~n33902;
  assign n12581 = n11975 & n12577;
  assign n12582 = n11890 & ~n33824;
  assign n12583 = ~n11976 & n12582;
  assign n12584 = ~n12442 & n12583;
  assign n12585 = ~n11890 & ~n33902;
  assign n12586 = ~n12584 & ~n12585;
  assign n12587 = ~n12580 & ~n12581;
  assign n12588 = ~n12575 & ~n33903;
  assign n12589 = ~n12573 & ~n12588;
  assign n12590 = ~n7512 & ~n12589;
  assign n12591 = n7512 & ~n12573;
  assign n12592 = ~n12588 & n12591;
  assign n12593 = n7512 & n12589;
  assign n12594 = ~n11978 & ~n11991;
  assign n12595 = ~n12442 & n12594;
  assign n12596 = ~n33825 & ~n12595;
  assign n12597 = n33825 & ~n11991;
  assign n12598 = ~n11978 & n12597;
  assign n12599 = n33825 & n12595;
  assign n12600 = ~n12442 & n12598;
  assign n12601 = n33825 & ~n12595;
  assign n12602 = ~n33825 & n12595;
  assign n12603 = ~n12601 & ~n12602;
  assign n12604 = ~n12596 & ~n33905;
  assign n12605 = ~n33904 & n33906;
  assign n12606 = ~n12590 & ~n12605;
  assign n12607 = ~n7015 & ~n12606;
  assign n12608 = n7015 & ~n12590;
  assign n12609 = ~n12605 & n12608;
  assign n12610 = ~n33826 & ~n11997;
  assign n12611 = ~n11997 & ~n12442;
  assign n12612 = ~n33826 & n12611;
  assign n12613 = ~n12442 & n12610;
  assign n12614 = n11882 & ~n33907;
  assign n12615 = n11996 & n12611;
  assign n12616 = n11882 & ~n33826;
  assign n12617 = ~n11997 & n12616;
  assign n12618 = ~n12442 & n12617;
  assign n12619 = ~n11882 & ~n33907;
  assign n12620 = ~n12618 & ~n12619;
  assign n12621 = ~n12614 & ~n12615;
  assign n12622 = ~n12609 & ~n33908;
  assign n12623 = ~n12607 & ~n12622;
  assign n12624 = ~n6579 & ~n12623;
  assign n12625 = n6579 & ~n12607;
  assign n12626 = ~n12622 & n12625;
  assign n12627 = n6579 & n12623;
  assign n12628 = ~n11999 & ~n12013;
  assign n12629 = ~n12442 & n12628;
  assign n12630 = n33828 & ~n12629;
  assign n12631 = ~n33828 & ~n12013;
  assign n12632 = ~n11999 & n12631;
  assign n12633 = ~n33828 & n12629;
  assign n12634 = ~n12442 & n12632;
  assign n12635 = n33828 & n12629;
  assign n12636 = ~n33828 & ~n12629;
  assign n12637 = ~n12635 & ~n12636;
  assign n12638 = ~n12630 & ~n33910;
  assign n12639 = ~n33909 & n33911;
  assign n12640 = ~n12624 & ~n12639;
  assign n12641 = ~n6117 & ~n12640;
  assign n12642 = n6117 & ~n12624;
  assign n12643 = ~n12639 & n12642;
  assign n12644 = ~n33829 & ~n12019;
  assign n12645 = ~n12019 & ~n12442;
  assign n12646 = ~n33829 & n12645;
  assign n12647 = ~n12442 & n12644;
  assign n12648 = n11874 & ~n33912;
  assign n12649 = n12018 & n12645;
  assign n12650 = n11874 & ~n33829;
  assign n12651 = ~n12019 & n12650;
  assign n12652 = ~n12442 & n12651;
  assign n12653 = ~n11874 & ~n33912;
  assign n12654 = ~n12652 & ~n12653;
  assign n12655 = ~n12648 & ~n12649;
  assign n12656 = ~n12643 & ~n33913;
  assign n12657 = ~n12641 & ~n12656;
  assign n12658 = ~n5708 & ~n12657;
  assign n12659 = n5708 & ~n12641;
  assign n12660 = ~n12656 & n12659;
  assign n12661 = n5708 & n12657;
  assign n12662 = ~n12021 & ~n12035;
  assign n12663 = ~n12035 & ~n12442;
  assign n12664 = ~n12021 & n12663;
  assign n12665 = ~n12442 & n12662;
  assign n12666 = ~n33831 & ~n33915;
  assign n12667 = n12033 & n12663;
  assign n12668 = n33831 & n33915;
  assign n12669 = ~n33831 & ~n12035;
  assign n12670 = ~n12021 & n12669;
  assign n12671 = ~n12442 & n12670;
  assign n12672 = n33831 & ~n33915;
  assign n12673 = ~n12671 & ~n12672;
  assign n12674 = ~n12666 & ~n33916;
  assign n12675 = ~n33914 & ~n33917;
  assign n12676 = ~n12658 & ~n12675;
  assign n12677 = ~n5278 & ~n12676;
  assign n12678 = n5278 & ~n12658;
  assign n12679 = ~n12675 & n12678;
  assign n12680 = ~n33832 & ~n12051;
  assign n12681 = ~n12442 & n12680;
  assign n12682 = ~n33833 & n12681;
  assign n12683 = n33833 & ~n12681;
  assign n12684 = ~n33832 & n33833;
  assign n12685 = ~n12051 & n12684;
  assign n12686 = ~n12442 & n12685;
  assign n12687 = ~n33833 & ~n12681;
  assign n12688 = ~n12686 & ~n12687;
  assign n12689 = ~n12682 & ~n12683;
  assign n12690 = ~n12679 & ~n33918;
  assign n12691 = ~n12677 & ~n12690;
  assign n12692 = ~n4903 & ~n12691;
  assign n12693 = n4903 & ~n12677;
  assign n12694 = ~n12690 & n12693;
  assign n12695 = n4903 & n12691;
  assign n12696 = ~n12053 & ~n12055;
  assign n12697 = ~n12442 & n12696;
  assign n12698 = ~n33834 & ~n12697;
  assign n12699 = ~n12053 & n33834;
  assign n12700 = ~n12055 & n12699;
  assign n12701 = n33834 & n12697;
  assign n12702 = ~n12442 & n12700;
  assign n12703 = ~n12698 & ~n33920;
  assign n12704 = ~n33919 & ~n12703;
  assign n12705 = ~n12692 & ~n12704;
  assign n12706 = ~n4508 & ~n12705;
  assign n12707 = n4508 & ~n12692;
  assign n12708 = ~n12704 & n12707;
  assign n12709 = ~n33886 & ~n12708;
  assign n12710 = ~n12706 & ~n12709;
  assign n12711 = ~n4155 & ~n12710;
  assign n12712 = ~n12074 & ~n12076;
  assign n12713 = ~n12442 & n12712;
  assign n12714 = ~n33839 & ~n12713;
  assign n12715 = ~n12074 & n33839;
  assign n12716 = ~n12076 & n12715;
  assign n12717 = n33839 & n12713;
  assign n12718 = ~n12442 & n12716;
  assign n12719 = ~n12714 & ~n33921;
  assign n12720 = n4155 & ~n12706;
  assign n12721 = ~n12709 & n12720;
  assign n12722 = n4155 & n12710;
  assign n12723 = ~n12719 & ~n33922;
  assign n12724 = ~n12711 & ~n12723;
  assign n12725 = ~n3788 & ~n12724;
  assign n12726 = n3788 & ~n12711;
  assign n12727 = ~n12723 & n12726;
  assign n12728 = ~n12093 & ~n33841;
  assign n12729 = ~n12093 & ~n12442;
  assign n12730 = ~n33841 & n12729;
  assign n12731 = ~n12442 & n12728;
  assign n12732 = n12101 & ~n33923;
  assign n12733 = n12105 & n12729;
  assign n12734 = n12101 & ~n33841;
  assign n12735 = ~n12093 & n12734;
  assign n12736 = ~n12442 & n12735;
  assign n12737 = ~n12101 & ~n33923;
  assign n12738 = ~n12736 & ~n12737;
  assign n12739 = ~n12732 & ~n12733;
  assign n12740 = ~n12727 & ~n33924;
  assign n12741 = ~n12725 & ~n12740;
  assign n12742 = ~n3473 & ~n12741;
  assign n12743 = n3473 & ~n12725;
  assign n12744 = ~n12740 & n12743;
  assign n12745 = n3473 & n12741;
  assign n12746 = ~n12107 & ~n12109;
  assign n12747 = ~n12442 & n12746;
  assign n12748 = ~n33844 & n12747;
  assign n12749 = n33844 & ~n12747;
  assign n12750 = ~n12107 & n33844;
  assign n12751 = ~n12109 & n12750;
  assign n12752 = n33844 & n12747;
  assign n12753 = ~n12442 & n12751;
  assign n12754 = ~n33844 & ~n12747;
  assign n12755 = ~n33926 & ~n12754;
  assign n12756 = ~n12748 & ~n12749;
  assign n12757 = ~n33925 & ~n33927;
  assign n12758 = ~n12742 & ~n12757;
  assign n12759 = ~n3140 & ~n12758;
  assign n12760 = n3140 & ~n12742;
  assign n12761 = ~n12757 & n12760;
  assign n12762 = ~n12125 & ~n33846;
  assign n12763 = ~n12125 & ~n12442;
  assign n12764 = ~n33846 & n12763;
  assign n12765 = ~n12442 & n12762;
  assign n12766 = n12133 & ~n33928;
  assign n12767 = n12137 & n12763;
  assign n12768 = n12133 & ~n33846;
  assign n12769 = ~n12125 & n12768;
  assign n12770 = ~n12442 & n12769;
  assign n12771 = ~n12133 & ~n33928;
  assign n12772 = ~n12770 & ~n12771;
  assign n12773 = ~n12766 & ~n12767;
  assign n12774 = ~n12761 & ~n33929;
  assign n12775 = ~n12759 & ~n12774;
  assign n12776 = ~n2855 & ~n12775;
  assign n12777 = n2855 & ~n12759;
  assign n12778 = ~n12774 & n12777;
  assign n12779 = n2855 & n12775;
  assign n12780 = ~n12139 & ~n12141;
  assign n12781 = ~n12139 & ~n12442;
  assign n12782 = ~n12141 & n12781;
  assign n12783 = ~n12442 & n12780;
  assign n12784 = n33848 & ~n33931;
  assign n12785 = n12153 & n12781;
  assign n12786 = ~n33848 & n33931;
  assign n12787 = ~n12139 & n33848;
  assign n12788 = ~n12141 & n12787;
  assign n12789 = ~n12442 & n12788;
  assign n12790 = ~n33848 & ~n33931;
  assign n12791 = ~n12789 & ~n12790;
  assign n12792 = ~n12784 & ~n33932;
  assign n12793 = ~n33930 & ~n33933;
  assign n12794 = ~n12776 & ~n12793;
  assign n12795 = ~n2556 & ~n12794;
  assign n12796 = n2556 & ~n12776;
  assign n12797 = ~n12793 & n12796;
  assign n12798 = ~n12155 & ~n33850;
  assign n12799 = ~n12155 & ~n12442;
  assign n12800 = ~n33850 & n12799;
  assign n12801 = ~n12442 & n12798;
  assign n12802 = n12163 & ~n33934;
  assign n12803 = n12167 & n12799;
  assign n12804 = n12163 & ~n33850;
  assign n12805 = ~n12155 & n12804;
  assign n12806 = ~n12442 & n12805;
  assign n12807 = ~n12163 & ~n33934;
  assign n12808 = ~n12806 & ~n12807;
  assign n12809 = ~n12802 & ~n12803;
  assign n12810 = ~n12797 & ~n33935;
  assign n12811 = ~n12795 & ~n12810;
  assign n12812 = ~n2301 & ~n12811;
  assign n12813 = ~n12169 & ~n12171;
  assign n12814 = ~n12442 & n12813;
  assign n12815 = ~n33853 & ~n12814;
  assign n12816 = ~n12169 & n33853;
  assign n12817 = ~n12171 & n12816;
  assign n12818 = n33853 & n12814;
  assign n12819 = ~n12442 & n12817;
  assign n12820 = ~n12815 & ~n33936;
  assign n12821 = n2301 & ~n12795;
  assign n12822 = ~n12810 & n12821;
  assign n12823 = n2301 & n12811;
  assign n12824 = ~n12820 & ~n33937;
  assign n12825 = ~n12812 & ~n12824;
  assign n12826 = ~n2038 & ~n12825;
  assign n12827 = n2038 & ~n12812;
  assign n12828 = ~n12824 & n12827;
  assign n12829 = ~n12187 & ~n33855;
  assign n12830 = ~n12187 & ~n12442;
  assign n12831 = ~n33855 & n12830;
  assign n12832 = ~n12442 & n12829;
  assign n12833 = n12195 & ~n33938;
  assign n12834 = n12199 & n12830;
  assign n12835 = n12195 & ~n33855;
  assign n12836 = ~n12187 & n12835;
  assign n12837 = ~n12442 & n12836;
  assign n12838 = ~n12195 & ~n33938;
  assign n12839 = ~n12837 & ~n12838;
  assign n12840 = ~n12833 & ~n12834;
  assign n12841 = ~n12828 & ~n33939;
  assign n12842 = ~n12826 & ~n12841;
  assign n12843 = ~n1812 & ~n12842;
  assign n12844 = n1812 & ~n12826;
  assign n12845 = ~n12841 & n12844;
  assign n12846 = n1812 & n12842;
  assign n12847 = ~n12201 & ~n12211;
  assign n12848 = ~n12201 & ~n12442;
  assign n12849 = ~n12211 & n12848;
  assign n12850 = ~n12442 & n12847;
  assign n12851 = n12209 & ~n33941;
  assign n12852 = n12212 & n12848;
  assign n12853 = ~n12201 & n12209;
  assign n12854 = ~n12211 & n12853;
  assign n12855 = ~n12442 & n12854;
  assign n12856 = ~n12209 & ~n33941;
  assign n12857 = ~n12855 & ~n12856;
  assign n12858 = ~n12851 & ~n12852;
  assign n12859 = ~n33940 & ~n33942;
  assign n12860 = ~n12843 & ~n12859;
  assign n12861 = ~n1582 & ~n12860;
  assign n12862 = n1582 & ~n12843;
  assign n12863 = ~n12859 & n12862;
  assign n12864 = ~n12214 & ~n33858;
  assign n12865 = ~n12214 & ~n12442;
  assign n12866 = ~n33858 & n12865;
  assign n12867 = ~n12442 & n12864;
  assign n12868 = n12222 & ~n33943;
  assign n12869 = n12226 & n12865;
  assign n12870 = n12222 & ~n33858;
  assign n12871 = ~n12214 & n12870;
  assign n12872 = ~n12442 & n12871;
  assign n12873 = ~n12222 & ~n33943;
  assign n12874 = ~n12872 & ~n12873;
  assign n12875 = ~n12868 & ~n12869;
  assign n12876 = ~n12863 & ~n33944;
  assign n12877 = ~n12861 & ~n12876;
  assign n12878 = ~n1388 & ~n12877;
  assign n12879 = ~n12228 & ~n12230;
  assign n12880 = ~n12442 & n12879;
  assign n12881 = ~n33860 & ~n12880;
  assign n12882 = ~n12228 & n33860;
  assign n12883 = ~n12230 & n12882;
  assign n12884 = n33860 & n12880;
  assign n12885 = ~n12442 & n12883;
  assign n12886 = ~n12881 & ~n33945;
  assign n12887 = n1388 & ~n12861;
  assign n12888 = ~n12876 & n12887;
  assign n12889 = n1388 & n12877;
  assign n12890 = ~n12886 & ~n33946;
  assign n12891 = ~n12878 & ~n12890;
  assign n12892 = ~n1192 & ~n12891;
  assign n12893 = n1192 & ~n12878;
  assign n12894 = ~n12890 & n12893;
  assign n12895 = ~n12245 & ~n33862;
  assign n12896 = ~n12245 & ~n12442;
  assign n12897 = ~n33862 & n12896;
  assign n12898 = ~n12442 & n12895;
  assign n12899 = n12253 & ~n33947;
  assign n12900 = n12257 & n12896;
  assign n12901 = n12253 & ~n33862;
  assign n12902 = ~n12245 & n12901;
  assign n12903 = ~n12442 & n12902;
  assign n12904 = ~n12253 & ~n33947;
  assign n12905 = ~n12903 & ~n12904;
  assign n12906 = ~n12899 & ~n12900;
  assign n12907 = ~n12894 & ~n33948;
  assign n12908 = ~n12892 & ~n12907;
  assign n12909 = ~n1028 & ~n12908;
  assign n12910 = n1028 & ~n12892;
  assign n12911 = ~n12907 & n12910;
  assign n12912 = n1028 & n12908;
  assign n12913 = ~n12259 & ~n12269;
  assign n12914 = ~n12259 & ~n12442;
  assign n12915 = ~n12269 & n12914;
  assign n12916 = ~n12442 & n12913;
  assign n12917 = n12267 & ~n33950;
  assign n12918 = n12270 & n12914;
  assign n12919 = ~n12259 & n12267;
  assign n12920 = ~n12269 & n12919;
  assign n12921 = ~n12442 & n12920;
  assign n12922 = ~n12267 & ~n33950;
  assign n12923 = ~n12921 & ~n12922;
  assign n12924 = ~n12917 & ~n12918;
  assign n12925 = ~n33949 & ~n33951;
  assign n12926 = ~n12909 & ~n12925;
  assign n12927 = ~n866 & ~n12926;
  assign n12928 = n866 & ~n12909;
  assign n12929 = ~n12925 & n12928;
  assign n12930 = ~n12272 & ~n33865;
  assign n12931 = ~n12272 & ~n12442;
  assign n12932 = ~n33865 & n12931;
  assign n12933 = ~n12442 & n12930;
  assign n12934 = n12280 & ~n33952;
  assign n12935 = n12284 & n12931;
  assign n12936 = n12280 & ~n33865;
  assign n12937 = ~n12272 & n12936;
  assign n12938 = ~n12442 & n12937;
  assign n12939 = ~n12280 & ~n33952;
  assign n12940 = ~n12938 & ~n12939;
  assign n12941 = ~n12934 & ~n12935;
  assign n12942 = ~n12929 & ~n33953;
  assign n12943 = ~n12927 & ~n12942;
  assign n12944 = ~n730 & ~n12943;
  assign n12945 = ~n12286 & ~n12288;
  assign n12946 = ~n12442 & n12945;
  assign n12947 = ~n33867 & ~n12946;
  assign n12948 = ~n12286 & n33867;
  assign n12949 = ~n12288 & n12948;
  assign n12950 = n33867 & n12946;
  assign n12951 = ~n12442 & n12949;
  assign n12952 = ~n12947 & ~n33954;
  assign n12953 = n730 & ~n12927;
  assign n12954 = ~n12942 & n12953;
  assign n12955 = n730 & n12943;
  assign n12956 = ~n12952 & ~n33955;
  assign n12957 = ~n12944 & ~n12956;
  assign n12958 = ~n602 & ~n12957;
  assign n12959 = n602 & ~n12944;
  assign n12960 = ~n12956 & n12959;
  assign n12961 = ~n12303 & ~n33869;
  assign n12962 = ~n12303 & ~n12442;
  assign n12963 = ~n33869 & n12962;
  assign n12964 = ~n12442 & n12961;
  assign n12965 = n12311 & ~n33956;
  assign n12966 = n12315 & n12962;
  assign n12967 = n12311 & ~n33869;
  assign n12968 = ~n12303 & n12967;
  assign n12969 = ~n12442 & n12968;
  assign n12970 = ~n12311 & ~n33956;
  assign n12971 = ~n12969 & ~n12970;
  assign n12972 = ~n12965 & ~n12966;
  assign n12973 = ~n12960 & ~n33957;
  assign n12974 = ~n12958 & ~n12973;
  assign n12975 = ~n497 & ~n12974;
  assign n12976 = n497 & ~n12958;
  assign n12977 = ~n12973 & n12976;
  assign n12978 = n497 & n12974;
  assign n12979 = ~n12317 & ~n12327;
  assign n12980 = ~n12317 & ~n12442;
  assign n12981 = ~n12327 & n12980;
  assign n12982 = ~n12442 & n12979;
  assign n12983 = n12325 & ~n33959;
  assign n12984 = n12328 & n12980;
  assign n12985 = ~n12317 & n12325;
  assign n12986 = ~n12327 & n12985;
  assign n12987 = ~n12442 & n12986;
  assign n12988 = ~n12325 & ~n33959;
  assign n12989 = ~n12987 & ~n12988;
  assign n12990 = ~n12983 & ~n12984;
  assign n12991 = ~n33958 & ~n33960;
  assign n12992 = ~n12975 & ~n12991;
  assign n12993 = ~n403 & ~n12992;
  assign n12994 = n403 & ~n12975;
  assign n12995 = ~n12991 & n12994;
  assign n12996 = ~n12330 & ~n33872;
  assign n12997 = ~n12330 & ~n12442;
  assign n12998 = ~n33872 & n12997;
  assign n12999 = ~n12442 & n12996;
  assign n13000 = n12338 & ~n33961;
  assign n13001 = n12342 & n12997;
  assign n13002 = n12338 & ~n33872;
  assign n13003 = ~n12330 & n13002;
  assign n13004 = ~n12442 & n13003;
  assign n13005 = ~n12338 & ~n33961;
  assign n13006 = ~n13004 & ~n13005;
  assign n13007 = ~n13000 & ~n13001;
  assign n13008 = ~n12995 & ~n33962;
  assign n13009 = ~n12993 & ~n13008;
  assign n13010 = ~n330 & ~n13009;
  assign n13011 = ~n12344 & ~n12346;
  assign n13012 = ~n12442 & n13011;
  assign n13013 = ~n33874 & ~n13012;
  assign n13014 = ~n12344 & n33874;
  assign n13015 = ~n12346 & n13014;
  assign n13016 = n33874 & n13012;
  assign n13017 = ~n12442 & n13015;
  assign n13018 = ~n13013 & ~n33963;
  assign n13019 = n330 & ~n12993;
  assign n13020 = ~n13008 & n13019;
  assign n13021 = n330 & n13009;
  assign n13022 = ~n13018 & ~n33964;
  assign n13023 = ~n13010 & ~n13022;
  assign n13024 = ~n271 & ~n13023;
  assign n13025 = n271 & ~n13010;
  assign n13026 = ~n13022 & n13025;
  assign n13027 = ~n12361 & ~n33876;
  assign n13028 = ~n12361 & ~n12442;
  assign n13029 = ~n33876 & n13028;
  assign n13030 = ~n12442 & n13027;
  assign n13031 = n12369 & ~n33965;
  assign n13032 = n12373 & n13028;
  assign n13033 = n12369 & ~n33876;
  assign n13034 = ~n12361 & n13033;
  assign n13035 = ~n12442 & n13034;
  assign n13036 = ~n12369 & ~n33965;
  assign n13037 = ~n13035 & ~n13036;
  assign n13038 = ~n13031 & ~n13032;
  assign n13039 = ~n13026 & ~n33966;
  assign n13040 = ~n13024 & ~n13039;
  assign n13041 = ~n217 & ~n13040;
  assign n13042 = n217 & ~n13024;
  assign n13043 = ~n13039 & n13042;
  assign n13044 = n217 & n13040;
  assign n13045 = ~n12375 & ~n12385;
  assign n13046 = ~n12375 & ~n12442;
  assign n13047 = ~n12385 & n13046;
  assign n13048 = ~n12442 & n13045;
  assign n13049 = n12383 & ~n33968;
  assign n13050 = n12386 & n13046;
  assign n13051 = ~n12375 & n12383;
  assign n13052 = ~n12385 & n13051;
  assign n13053 = ~n12442 & n13052;
  assign n13054 = ~n12383 & ~n33968;
  assign n13055 = ~n13053 & ~n13054;
  assign n13056 = ~n13049 & ~n13050;
  assign n13057 = ~n33967 & ~n33969;
  assign n13058 = ~n13041 & ~n13057;
  assign n13059 = ~n198 & ~n13058;
  assign n13060 = n198 & ~n13041;
  assign n13061 = ~n13057 & n13060;
  assign n13062 = ~n12388 & ~n33879;
  assign n13063 = ~n12388 & ~n12442;
  assign n13064 = ~n33879 & n13063;
  assign n13065 = ~n12442 & n13062;
  assign n13066 = n12396 & ~n33970;
  assign n13067 = n12400 & n13063;
  assign n13068 = n12396 & ~n33879;
  assign n13069 = ~n12388 & n13068;
  assign n13070 = ~n12442 & n13069;
  assign n13071 = ~n12396 & ~n33970;
  assign n13072 = ~n13070 & ~n13071;
  assign n13073 = ~n13066 & ~n13067;
  assign n13074 = ~n13061 & ~n33971;
  assign n13075 = ~n13059 & ~n13074;
  assign n13076 = ~n12402 & ~n12404;
  assign n13077 = ~n12442 & n13076;
  assign n13078 = ~n33881 & ~n13077;
  assign n13079 = ~n12402 & n33881;
  assign n13080 = ~n12404 & n13079;
  assign n13081 = n33881 & n13077;
  assign n13082 = ~n12442 & n13080;
  assign n13083 = ~n13078 & ~n33972;
  assign n13084 = ~n12418 & ~n12426;
  assign n13085 = ~n12426 & ~n12442;
  assign n13086 = ~n12418 & n13085;
  assign n13087 = ~n12442 & n13084;
  assign n13088 = ~n33884 & ~n33973;
  assign n13089 = ~n13083 & n13088;
  assign n13090 = ~n13075 & n13089;
  assign n13091 = n193 & ~n13090;
  assign n13092 = ~n13059 & n13083;
  assign n13093 = ~n13074 & n13092;
  assign n13094 = n13075 & n13083;
  assign n13095 = n12418 & ~n13085;
  assign n13096 = ~n193 & ~n13084;
  assign n13097 = ~n13095 & n13096;
  assign n13098 = ~n33974 & ~n13097;
  assign n13099 = ~n13091 & n13098;
  assign n13100 = ~n12706 & ~n12708;
  assign n13101 = ~n13099 & n13100;
  assign n13102 = ~n33886 & ~n13101;
  assign n13103 = n33886 & ~n12708;
  assign n13104 = ~n12706 & n13103;
  assign n13105 = n33886 & n13101;
  assign n13106 = ~n13099 & n13104;
  assign n13107 = ~n13102 & ~n33975;
  assign n13108 = ~n12677 & ~n12679;
  assign n13109 = ~n13099 & n13108;
  assign n13110 = ~n33918 & ~n13109;
  assign n13111 = ~n12679 & n33918;
  assign n13112 = ~n12677 & n13111;
  assign n13113 = n33918 & n13109;
  assign n13114 = ~n13099 & n13112;
  assign n13115 = ~n13110 & ~n33976;
  assign n13116 = ~n12641 & ~n12643;
  assign n13117 = ~n13099 & n13116;
  assign n13118 = ~n33913 & ~n13117;
  assign n13119 = ~n12643 & n33913;
  assign n13120 = ~n12641 & n13119;
  assign n13121 = n33913 & n13117;
  assign n13122 = ~n13099 & n13120;
  assign n13123 = ~n13118 & ~n33977;
  assign n13124 = ~n12607 & ~n12609;
  assign n13125 = ~n13099 & n13124;
  assign n13126 = ~n33908 & ~n13125;
  assign n13127 = ~n12609 & n33908;
  assign n13128 = ~n12607 & n13127;
  assign n13129 = n33908 & n13125;
  assign n13130 = ~n13099 & n13128;
  assign n13131 = ~n13126 & ~n33978;
  assign n13132 = ~n12573 & ~n12575;
  assign n13133 = ~n13099 & n13132;
  assign n13134 = ~n33903 & ~n13133;
  assign n13135 = ~n12575 & n33903;
  assign n13136 = ~n12573 & n13135;
  assign n13137 = n33903 & n13133;
  assign n13138 = ~n13099 & n13136;
  assign n13139 = ~n13134 & ~n33979;
  assign n13140 = ~n12540 & ~n12542;
  assign n13141 = ~n13099 & n13140;
  assign n13142 = ~n33899 & ~n13141;
  assign n13143 = ~n12542 & n33899;
  assign n13144 = ~n12540 & n13143;
  assign n13145 = n33899 & n13141;
  assign n13146 = ~n13099 & n13144;
  assign n13147 = ~n13142 & ~n33980;
  assign n13148 = ~n12506 & ~n12508;
  assign n13149 = ~n13099 & n13148;
  assign n13150 = ~n33894 & ~n13149;
  assign n13151 = ~n12508 & n33894;
  assign n13152 = ~n12506 & n13151;
  assign n13153 = n33894 & n13149;
  assign n13154 = ~n13099 & n13152;
  assign n13155 = ~n13150 & ~n33981;
  assign n13156 = ~n12479 & ~n12481;
  assign n13157 = ~n13099 & n13156;
  assign n13158 = ~n12490 & ~n13157;
  assign n13159 = ~n12481 & n12490;
  assign n13160 = ~n12479 & n13159;
  assign n13161 = n12490 & n13157;
  assign n13162 = ~n13099 & n13160;
  assign n13163 = ~n13158 & ~n33982;
  assign n13164 = ~pi46  & ~n13099;
  assign n13165 = ~pi47  & n13164;
  assign n13166 = n12456 & ~n13099;
  assign n13167 = ~n12442 & ~n13097;
  assign n13168 = ~n33974 & n13167;
  assign n13169 = ~n13091 & n13168;
  assign n13170 = ~n33983 & ~n13169;
  assign n13171 = pi48  & ~n13170;
  assign n13172 = ~pi48  & ~n13169;
  assign n13173 = ~pi48  & n13170;
  assign n13174 = ~n33983 & n13172;
  assign n13175 = ~n13171 & ~n33984;
  assign n13176 = pi46  & ~n13099;
  assign n13177 = ~pi44  & ~pi45 ;
  assign n13178 = ~pi46  & n13177;
  assign n13179 = ~n11839 & ~n33888;
  assign n13180 = ~n11840 & n13179;
  assign n13181 = ~n11856 & n13180;
  assign n13182 = ~n33809 & n13181;
  assign n13183 = n33807 & n11858;
  assign n13184 = ~n11850 & n13182;
  assign n13185 = ~n13178 & ~n33985;
  assign n13186 = ~n12440 & n13185;
  assign n13187 = ~n33884 & n13186;
  assign n13188 = ~n12434 & n13187;
  assign n13189 = ~n13176 & ~n13178;
  assign n13190 = n12442 & n13189;
  assign n13191 = ~n13176 & n13188;
  assign n13192 = pi47  & ~n13164;
  assign n13193 = ~n33983 & ~n13192;
  assign n13194 = ~n33986 & n13193;
  assign n13195 = ~n12442 & ~n13189;
  assign n13196 = n11858 & ~n13195;
  assign n13197 = ~n13194 & ~n13195;
  assign n13198 = n11858 & n13197;
  assign n13199 = ~n13194 & n13196;
  assign n13200 = ~n13175 & ~n33987;
  assign n13201 = ~n11858 & ~n13197;
  assign n13202 = n11229 & ~n13201;
  assign n13203 = ~n13200 & n13202;
  assign n13204 = ~n12459 & ~n33889;
  assign n13205 = ~n13099 & n13204;
  assign n13206 = n12464 & ~n13205;
  assign n13207 = ~n12464 & n13204;
  assign n13208 = ~n12464 & n13205;
  assign n13209 = ~n13099 & n13207;
  assign n13210 = ~n13206 & ~n33988;
  assign n13211 = ~n13203 & ~n13210;
  assign n13212 = ~n13200 & ~n13201;
  assign n13213 = ~n11229 & ~n13212;
  assign n13214 = n10681 & ~n13213;
  assign n13215 = ~n13211 & ~n13213;
  assign n13216 = n10681 & n13215;
  assign n13217 = ~n13211 & n13214;
  assign n13218 = ~n13163 & ~n33989;
  assign n13219 = ~n10681 & ~n13215;
  assign n13220 = n10086 & ~n13219;
  assign n13221 = ~n13218 & n13220;
  assign n13222 = ~n12493 & ~n33891;
  assign n13223 = ~n13099 & n13222;
  assign n13224 = n12503 & ~n13223;
  assign n13225 = ~n12503 & n13223;
  assign n13226 = ~n12493 & n12503;
  assign n13227 = ~n33891 & n13226;
  assign n13228 = n12503 & n13223;
  assign n13229 = ~n13099 & n13227;
  assign n13230 = ~n12503 & ~n13223;
  assign n13231 = ~n33990 & ~n13230;
  assign n13232 = ~n13224 & ~n13225;
  assign n13233 = ~n13221 & ~n33991;
  assign n13234 = ~n13218 & ~n13219;
  assign n13235 = ~n10086 & ~n13234;
  assign n13236 = n9565 & ~n13235;
  assign n13237 = ~n13233 & ~n13235;
  assign n13238 = n9565 & n13237;
  assign n13239 = ~n13233 & n13236;
  assign n13240 = ~n13155 & ~n33992;
  assign n13241 = ~n9565 & ~n13237;
  assign n13242 = n8998 & ~n13241;
  assign n13243 = ~n13240 & n13242;
  assign n13244 = ~n12523 & ~n33895;
  assign n13245 = ~n13099 & n13244;
  assign n13246 = ~n33897 & n13245;
  assign n13247 = n33897 & ~n13245;
  assign n13248 = ~n12523 & n33897;
  assign n13249 = ~n33895 & n13248;
  assign n13250 = ~n13099 & n13249;
  assign n13251 = ~n33897 & ~n13245;
  assign n13252 = ~n13250 & ~n13251;
  assign n13253 = ~n13246 & ~n13247;
  assign n13254 = ~n13243 & ~n33993;
  assign n13255 = ~n13240 & ~n13241;
  assign n13256 = ~n8998 & ~n13255;
  assign n13257 = n8506 & ~n13256;
  assign n13258 = ~n13254 & ~n13256;
  assign n13259 = n8506 & n13258;
  assign n13260 = ~n13254 & n13257;
  assign n13261 = ~n13147 & ~n33994;
  assign n13262 = ~n8506 & ~n13258;
  assign n13263 = n7975 & ~n13262;
  assign n13264 = ~n13261 & n13263;
  assign n13265 = ~n12557 & ~n33900;
  assign n13266 = ~n13099 & n13265;
  assign n13267 = ~n33901 & ~n13266;
  assign n13268 = ~n12557 & n33901;
  assign n13269 = ~n33900 & n13268;
  assign n13270 = n33901 & n13266;
  assign n13271 = ~n13099 & n13269;
  assign n13272 = n33901 & ~n13266;
  assign n13273 = ~n33901 & n13266;
  assign n13274 = ~n13272 & ~n13273;
  assign n13275 = ~n13267 & ~n33995;
  assign n13276 = ~n13264 & n33996;
  assign n13277 = ~n13261 & ~n13262;
  assign n13278 = ~n7975 & ~n13277;
  assign n13279 = n7512 & ~n13278;
  assign n13280 = ~n13276 & ~n13278;
  assign n13281 = n7512 & n13280;
  assign n13282 = ~n13276 & n13279;
  assign n13283 = ~n13139 & ~n33997;
  assign n13284 = ~n7512 & ~n13280;
  assign n13285 = n7015 & ~n13284;
  assign n13286 = ~n13283 & n13285;
  assign n13287 = ~n12590 & ~n33904;
  assign n13288 = ~n13099 & n13287;
  assign n13289 = n33906 & ~n13288;
  assign n13290 = ~n12590 & ~n33906;
  assign n13291 = ~n33904 & n13290;
  assign n13292 = ~n33906 & n13288;
  assign n13293 = ~n13099 & n13291;
  assign n13294 = n33906 & n13288;
  assign n13295 = ~n33906 & ~n13288;
  assign n13296 = ~n13294 & ~n13295;
  assign n13297 = ~n13289 & ~n33998;
  assign n13298 = ~n13286 & n33999;
  assign n13299 = ~n13283 & ~n13284;
  assign n13300 = ~n7015 & ~n13299;
  assign n13301 = n6579 & ~n13300;
  assign n13302 = ~n13298 & ~n13300;
  assign n13303 = n6579 & n13302;
  assign n13304 = ~n13298 & n13301;
  assign n13305 = ~n13131 & ~n34000;
  assign n13306 = ~n6579 & ~n13302;
  assign n13307 = n6117 & ~n13306;
  assign n13308 = ~n13305 & n13307;
  assign n13309 = ~n12624 & ~n33909;
  assign n13310 = ~n12624 & ~n13099;
  assign n13311 = ~n33909 & n13310;
  assign n13312 = ~n13099 & n13309;
  assign n13313 = ~n33911 & ~n34001;
  assign n13314 = n12639 & n13310;
  assign n13315 = n33911 & n34001;
  assign n13316 = ~n12624 & ~n33911;
  assign n13317 = ~n33909 & n13316;
  assign n13318 = ~n13099 & n13317;
  assign n13319 = n33911 & ~n34001;
  assign n13320 = ~n13318 & ~n13319;
  assign n13321 = ~n13313 & ~n34002;
  assign n13322 = ~n13308 & ~n34003;
  assign n13323 = ~n13305 & ~n13306;
  assign n13324 = ~n6117 & ~n13323;
  assign n13325 = n5708 & ~n13324;
  assign n13326 = ~n13322 & ~n13324;
  assign n13327 = n5708 & n13326;
  assign n13328 = ~n13322 & n13325;
  assign n13329 = ~n13123 & ~n34004;
  assign n13330 = ~n5708 & ~n13326;
  assign n13331 = n5278 & ~n13330;
  assign n13332 = ~n13329 & n13331;
  assign n13333 = ~n12658 & ~n33914;
  assign n13334 = ~n13099 & n13333;
  assign n13335 = ~n33917 & ~n13334;
  assign n13336 = ~n12658 & n33917;
  assign n13337 = ~n33914 & n13336;
  assign n13338 = n33917 & n13334;
  assign n13339 = ~n13099 & n13337;
  assign n13340 = ~n13335 & ~n34005;
  assign n13341 = ~n13332 & ~n13340;
  assign n13342 = ~n13329 & ~n13330;
  assign n13343 = ~n5278 & ~n13342;
  assign n13344 = n4903 & ~n13343;
  assign n13345 = ~n13341 & ~n13343;
  assign n13346 = n4903 & n13345;
  assign n13347 = ~n13341 & n13344;
  assign n13348 = ~n13115 & ~n34006;
  assign n13349 = ~n4903 & ~n13345;
  assign n13350 = ~n13348 & ~n13349;
  assign n13351 = ~n4508 & ~n13350;
  assign n13352 = n4508 & ~n13349;
  assign n13353 = ~n13348 & n13352;
  assign n13354 = ~n12692 & ~n33919;
  assign n13355 = ~n13099 & n13354;
  assign n13356 = n12703 & ~n13355;
  assign n13357 = ~n12703 & n13355;
  assign n13358 = ~n12692 & n12703;
  assign n13359 = ~n33919 & n13358;
  assign n13360 = n12703 & n13355;
  assign n13361 = ~n13099 & n13359;
  assign n13362 = ~n12703 & ~n13355;
  assign n13363 = ~n34007 & ~n13362;
  assign n13364 = ~n13356 & ~n13357;
  assign n13365 = ~n13353 & ~n34008;
  assign n13366 = ~n13351 & ~n13365;
  assign n13367 = ~n4155 & ~n13366;
  assign n13368 = n4155 & ~n13351;
  assign n13369 = n4155 & n13366;
  assign n13370 = ~n13365 & n13368;
  assign n13371 = ~n13107 & ~n34009;
  assign n13372 = ~n13367 & ~n13371;
  assign n13373 = ~n3788 & ~n13372;
  assign n13374 = n3788 & ~n13367;
  assign n13375 = ~n13371 & n13374;
  assign n13376 = ~n12711 & ~n33922;
  assign n13377 = ~n12711 & ~n13099;
  assign n13378 = ~n33922 & n13377;
  assign n13379 = ~n13099 & n13376;
  assign n13380 = n12719 & ~n34010;
  assign n13381 = n12723 & n13377;
  assign n13382 = ~n12711 & n12719;
  assign n13383 = ~n33922 & n13382;
  assign n13384 = ~n13099 & n13383;
  assign n13385 = ~n12719 & ~n34010;
  assign n13386 = ~n13384 & ~n13385;
  assign n13387 = ~n13380 & ~n13381;
  assign n13388 = ~n13375 & ~n34011;
  assign n13389 = ~n13373 & ~n13388;
  assign n13390 = ~n3473 & ~n13389;
  assign n13391 = ~n12725 & ~n12727;
  assign n13392 = ~n13099 & n13391;
  assign n13393 = ~n33924 & ~n13392;
  assign n13394 = ~n12727 & n33924;
  assign n13395 = ~n12725 & n13394;
  assign n13396 = n33924 & n13392;
  assign n13397 = ~n13099 & n13395;
  assign n13398 = ~n13393 & ~n34012;
  assign n13399 = n3473 & ~n13373;
  assign n13400 = n3473 & n13389;
  assign n13401 = ~n13388 & n13399;
  assign n13402 = ~n13398 & ~n34013;
  assign n13403 = ~n13390 & ~n13402;
  assign n13404 = ~n3140 & ~n13403;
  assign n13405 = n3140 & ~n13390;
  assign n13406 = ~n13402 & n13405;
  assign n13407 = ~n12742 & ~n33925;
  assign n13408 = ~n12742 & ~n13099;
  assign n13409 = ~n33925 & n13408;
  assign n13410 = ~n13099 & n13407;
  assign n13411 = n33927 & ~n34014;
  assign n13412 = n12757 & n13408;
  assign n13413 = ~n33927 & n34014;
  assign n13414 = ~n12742 & n33927;
  assign n13415 = ~n33925 & n13414;
  assign n13416 = ~n13099 & n13415;
  assign n13417 = ~n33927 & ~n34014;
  assign n13418 = ~n13416 & ~n13417;
  assign n13419 = ~n13411 & ~n34015;
  assign n13420 = ~n13406 & ~n34016;
  assign n13421 = ~n13404 & ~n13420;
  assign n13422 = ~n2855 & ~n13421;
  assign n13423 = ~n12759 & ~n12761;
  assign n13424 = ~n13099 & n13423;
  assign n13425 = ~n33929 & ~n13424;
  assign n13426 = ~n12761 & n33929;
  assign n13427 = ~n12759 & n13426;
  assign n13428 = n33929 & n13424;
  assign n13429 = ~n13099 & n13427;
  assign n13430 = ~n13425 & ~n34017;
  assign n13431 = n2855 & ~n13404;
  assign n13432 = n2855 & n13421;
  assign n13433 = ~n13420 & n13431;
  assign n13434 = ~n13430 & ~n34018;
  assign n13435 = ~n13422 & ~n13434;
  assign n13436 = ~n2556 & ~n13435;
  assign n13437 = ~n12776 & ~n33930;
  assign n13438 = ~n13099 & n13437;
  assign n13439 = ~n33933 & ~n13438;
  assign n13440 = ~n12776 & n33933;
  assign n13441 = ~n33930 & n13440;
  assign n13442 = n33933 & n13438;
  assign n13443 = ~n13099 & n13441;
  assign n13444 = ~n13439 & ~n34019;
  assign n13445 = n2556 & ~n13422;
  assign n13446 = ~n13434 & n13445;
  assign n13447 = ~n13444 & ~n13446;
  assign n13448 = ~n13436 & ~n13447;
  assign n13449 = ~n2301 & ~n13448;
  assign n13450 = ~n12795 & ~n12797;
  assign n13451 = ~n13099 & n13450;
  assign n13452 = ~n33935 & ~n13451;
  assign n13453 = ~n12797 & n33935;
  assign n13454 = ~n12795 & n13453;
  assign n13455 = n33935 & n13451;
  assign n13456 = ~n13099 & n13454;
  assign n13457 = ~n13452 & ~n34020;
  assign n13458 = n2301 & ~n13436;
  assign n13459 = n2301 & n13448;
  assign n13460 = ~n13447 & n13458;
  assign n13461 = ~n13457 & ~n34021;
  assign n13462 = ~n13449 & ~n13461;
  assign n13463 = ~n2038 & ~n13462;
  assign n13464 = n2038 & ~n13449;
  assign n13465 = ~n13461 & n13464;
  assign n13466 = ~n12812 & ~n33937;
  assign n13467 = ~n12812 & ~n13099;
  assign n13468 = ~n33937 & n13467;
  assign n13469 = ~n13099 & n13466;
  assign n13470 = n12820 & ~n34022;
  assign n13471 = n12824 & n13467;
  assign n13472 = ~n12812 & n12820;
  assign n13473 = ~n33937 & n13472;
  assign n13474 = ~n13099 & n13473;
  assign n13475 = ~n12820 & ~n34022;
  assign n13476 = ~n13474 & ~n13475;
  assign n13477 = ~n13470 & ~n13471;
  assign n13478 = ~n13465 & ~n34023;
  assign n13479 = ~n13463 & ~n13478;
  assign n13480 = ~n1812 & ~n13479;
  assign n13481 = ~n12826 & ~n12828;
  assign n13482 = ~n13099 & n13481;
  assign n13483 = ~n33939 & ~n13482;
  assign n13484 = ~n12828 & n33939;
  assign n13485 = ~n12826 & n13484;
  assign n13486 = n33939 & n13482;
  assign n13487 = ~n13099 & n13485;
  assign n13488 = ~n13483 & ~n34024;
  assign n13489 = n1812 & ~n13463;
  assign n13490 = n1812 & n13479;
  assign n13491 = ~n13478 & n13489;
  assign n13492 = ~n13488 & ~n34025;
  assign n13493 = ~n13480 & ~n13492;
  assign n13494 = ~n1582 & ~n13493;
  assign n13495 = ~n12843 & ~n33940;
  assign n13496 = ~n13099 & n13495;
  assign n13497 = ~n33942 & ~n13496;
  assign n13498 = ~n12843 & n33942;
  assign n13499 = ~n33940 & n13498;
  assign n13500 = n33942 & n13496;
  assign n13501 = ~n13099 & n13499;
  assign n13502 = ~n13497 & ~n34026;
  assign n13503 = n1582 & ~n13480;
  assign n13504 = ~n13492 & n13503;
  assign n13505 = ~n13502 & ~n13504;
  assign n13506 = ~n13494 & ~n13505;
  assign n13507 = ~n1388 & ~n13506;
  assign n13508 = ~n12861 & ~n12863;
  assign n13509 = ~n13099 & n13508;
  assign n13510 = ~n33944 & ~n13509;
  assign n13511 = ~n12863 & n33944;
  assign n13512 = ~n12861 & n13511;
  assign n13513 = n33944 & n13509;
  assign n13514 = ~n13099 & n13512;
  assign n13515 = ~n13510 & ~n34027;
  assign n13516 = n1388 & ~n13494;
  assign n13517 = n1388 & n13506;
  assign n13518 = ~n13505 & n13516;
  assign n13519 = ~n13515 & ~n34028;
  assign n13520 = ~n13507 & ~n13519;
  assign n13521 = ~n1192 & ~n13520;
  assign n13522 = n1192 & ~n13507;
  assign n13523 = ~n13519 & n13522;
  assign n13524 = ~n12878 & ~n33946;
  assign n13525 = ~n12878 & ~n13099;
  assign n13526 = ~n33946 & n13525;
  assign n13527 = ~n13099 & n13524;
  assign n13528 = n12886 & ~n34029;
  assign n13529 = n12890 & n13525;
  assign n13530 = ~n12878 & n12886;
  assign n13531 = ~n33946 & n13530;
  assign n13532 = ~n13099 & n13531;
  assign n13533 = ~n12886 & ~n34029;
  assign n13534 = ~n13532 & ~n13533;
  assign n13535 = ~n13528 & ~n13529;
  assign n13536 = ~n13523 & ~n34030;
  assign n13537 = ~n13521 & ~n13536;
  assign n13538 = ~n1028 & ~n13537;
  assign n13539 = ~n12892 & ~n12894;
  assign n13540 = ~n13099 & n13539;
  assign n13541 = ~n33948 & ~n13540;
  assign n13542 = ~n12894 & n33948;
  assign n13543 = ~n12892 & n13542;
  assign n13544 = n33948 & n13540;
  assign n13545 = ~n13099 & n13543;
  assign n13546 = ~n13541 & ~n34031;
  assign n13547 = n1028 & ~n13521;
  assign n13548 = n1028 & n13537;
  assign n13549 = ~n13536 & n13547;
  assign n13550 = ~n13546 & ~n34032;
  assign n13551 = ~n13538 & ~n13550;
  assign n13552 = ~n866 & ~n13551;
  assign n13553 = ~n12909 & ~n33949;
  assign n13554 = ~n13099 & n13553;
  assign n13555 = ~n33951 & ~n13554;
  assign n13556 = ~n12909 & n33951;
  assign n13557 = ~n33949 & n13556;
  assign n13558 = n33951 & n13554;
  assign n13559 = ~n13099 & n13557;
  assign n13560 = ~n13555 & ~n34033;
  assign n13561 = n866 & ~n13538;
  assign n13562 = ~n13550 & n13561;
  assign n13563 = ~n13560 & ~n13562;
  assign n13564 = ~n13552 & ~n13563;
  assign n13565 = ~n730 & ~n13564;
  assign n13566 = ~n12927 & ~n12929;
  assign n13567 = ~n13099 & n13566;
  assign n13568 = ~n33953 & ~n13567;
  assign n13569 = ~n12929 & n33953;
  assign n13570 = ~n12927 & n13569;
  assign n13571 = n33953 & n13567;
  assign n13572 = ~n13099 & n13570;
  assign n13573 = ~n13568 & ~n34034;
  assign n13574 = n730 & ~n13552;
  assign n13575 = n730 & n13564;
  assign n13576 = ~n13563 & n13574;
  assign n13577 = ~n13573 & ~n34035;
  assign n13578 = ~n13565 & ~n13577;
  assign n13579 = ~n602 & ~n13578;
  assign n13580 = n602 & ~n13565;
  assign n13581 = ~n13577 & n13580;
  assign n13582 = ~n12944 & ~n33955;
  assign n13583 = ~n12944 & ~n13099;
  assign n13584 = ~n33955 & n13583;
  assign n13585 = ~n13099 & n13582;
  assign n13586 = n12952 & ~n34036;
  assign n13587 = n12956 & n13583;
  assign n13588 = ~n12944 & n12952;
  assign n13589 = ~n33955 & n13588;
  assign n13590 = ~n13099 & n13589;
  assign n13591 = ~n12952 & ~n34036;
  assign n13592 = ~n13590 & ~n13591;
  assign n13593 = ~n13586 & ~n13587;
  assign n13594 = ~n13581 & ~n34037;
  assign n13595 = ~n13579 & ~n13594;
  assign n13596 = ~n497 & ~n13595;
  assign n13597 = ~n12958 & ~n12960;
  assign n13598 = ~n13099 & n13597;
  assign n13599 = ~n33957 & ~n13598;
  assign n13600 = ~n12960 & n33957;
  assign n13601 = ~n12958 & n13600;
  assign n13602 = n33957 & n13598;
  assign n13603 = ~n13099 & n13601;
  assign n13604 = ~n13599 & ~n34038;
  assign n13605 = n497 & ~n13579;
  assign n13606 = n497 & n13595;
  assign n13607 = ~n13594 & n13605;
  assign n13608 = ~n13604 & ~n34039;
  assign n13609 = ~n13596 & ~n13608;
  assign n13610 = ~n403 & ~n13609;
  assign n13611 = ~n12975 & ~n33958;
  assign n13612 = ~n13099 & n13611;
  assign n13613 = ~n33960 & ~n13612;
  assign n13614 = ~n12975 & n33960;
  assign n13615 = ~n33958 & n13614;
  assign n13616 = n33960 & n13612;
  assign n13617 = ~n13099 & n13615;
  assign n13618 = ~n13613 & ~n34040;
  assign n13619 = n403 & ~n13596;
  assign n13620 = ~n13608 & n13619;
  assign n13621 = ~n13618 & ~n13620;
  assign n13622 = ~n13610 & ~n13621;
  assign n13623 = ~n330 & ~n13622;
  assign n13624 = ~n12993 & ~n12995;
  assign n13625 = ~n13099 & n13624;
  assign n13626 = ~n33962 & ~n13625;
  assign n13627 = ~n12995 & n33962;
  assign n13628 = ~n12993 & n13627;
  assign n13629 = n33962 & n13625;
  assign n13630 = ~n13099 & n13628;
  assign n13631 = ~n13626 & ~n34041;
  assign n13632 = n330 & ~n13610;
  assign n13633 = n330 & n13622;
  assign n13634 = ~n13621 & n13632;
  assign n13635 = ~n13631 & ~n34042;
  assign n13636 = ~n13623 & ~n13635;
  assign n13637 = ~n271 & ~n13636;
  assign n13638 = n271 & ~n13623;
  assign n13639 = ~n13635 & n13638;
  assign n13640 = ~n13010 & ~n33964;
  assign n13641 = ~n13010 & ~n13099;
  assign n13642 = ~n33964 & n13641;
  assign n13643 = ~n13099 & n13640;
  assign n13644 = n13018 & ~n34043;
  assign n13645 = n13022 & n13641;
  assign n13646 = ~n13010 & n13018;
  assign n13647 = ~n33964 & n13646;
  assign n13648 = ~n13099 & n13647;
  assign n13649 = ~n13018 & ~n34043;
  assign n13650 = ~n13648 & ~n13649;
  assign n13651 = ~n13644 & ~n13645;
  assign n13652 = ~n13639 & ~n34044;
  assign n13653 = ~n13637 & ~n13652;
  assign n13654 = ~n217 & ~n13653;
  assign n13655 = ~n13024 & ~n13026;
  assign n13656 = ~n13099 & n13655;
  assign n13657 = ~n33966 & ~n13656;
  assign n13658 = ~n13026 & n33966;
  assign n13659 = ~n13024 & n13658;
  assign n13660 = n33966 & n13656;
  assign n13661 = ~n13099 & n13659;
  assign n13662 = ~n13657 & ~n34045;
  assign n13663 = n217 & ~n13637;
  assign n13664 = n217 & n13653;
  assign n13665 = ~n13652 & n13663;
  assign n13666 = ~n13662 & ~n34046;
  assign n13667 = ~n13654 & ~n13666;
  assign n13668 = ~n198 & ~n13667;
  assign n13669 = ~n13041 & ~n33967;
  assign n13670 = ~n13099 & n13669;
  assign n13671 = ~n33969 & ~n13670;
  assign n13672 = ~n13041 & n33969;
  assign n13673 = ~n33967 & n13672;
  assign n13674 = n33969 & n13670;
  assign n13675 = ~n13099 & n13673;
  assign n13676 = ~n13671 & ~n34047;
  assign n13677 = n198 & ~n13654;
  assign n13678 = ~n13666 & n13677;
  assign n13679 = ~n13676 & ~n13678;
  assign n13680 = ~n13668 & ~n13679;
  assign n13681 = ~n13059 & ~n13061;
  assign n13682 = ~n13099 & n13681;
  assign n13683 = ~n33971 & ~n13682;
  assign n13684 = ~n13061 & n33971;
  assign n13685 = ~n13059 & n13684;
  assign n13686 = n33971 & n13682;
  assign n13687 = ~n13099 & n13685;
  assign n13688 = ~n13683 & ~n34048;
  assign n13689 = ~n13075 & ~n13083;
  assign n13690 = ~n13083 & ~n13099;
  assign n13691 = ~n13075 & n13690;
  assign n13692 = ~n13099 & n13689;
  assign n13693 = ~n33974 & ~n34049;
  assign n13694 = ~n13688 & n13693;
  assign n13695 = ~n13680 & n13694;
  assign n13696 = n193 & ~n13695;
  assign n13697 = ~n13668 & n13688;
  assign n13698 = n13680 & n13688;
  assign n13699 = ~n13679 & n13697;
  assign n13700 = n13075 & ~n13690;
  assign n13701 = ~n193 & ~n13689;
  assign n13702 = ~n13700 & n13701;
  assign n13703 = ~n34050 & ~n13702;
  assign n13704 = ~n13696 & n13703;
  assign n13705 = ~n13367 & ~n34009;
  assign n13706 = ~n13367 & ~n13704;
  assign n13707 = ~n34009 & n13706;
  assign n13708 = ~n13704 & n13705;
  assign n13709 = n13107 & ~n34051;
  assign n13710 = n13371 & n13706;
  assign n13711 = n13107 & ~n34009;
  assign n13712 = ~n13367 & n13711;
  assign n13713 = ~n13704 & n13712;
  assign n13714 = ~n13107 & ~n34051;
  assign n13715 = ~n13713 & ~n13714;
  assign n13716 = ~n13709 & ~n13710;
  assign n13717 = pi44  & ~n13704;
  assign n13718 = ~pi42  & ~pi43 ;
  assign n13719 = ~pi44  & n13718;
  assign n13720 = ~n13717 & ~n13719;
  assign n13721 = ~n13099 & ~n13720;
  assign n13722 = ~pi44  & ~n13704;
  assign n13723 = pi45  & ~n13722;
  assign n13724 = ~pi45  & n13722;
  assign n13725 = n13177 & ~n13704;
  assign n13726 = ~n13723 & ~n34053;
  assign n13727 = ~n33882 & ~n33985;
  assign n13728 = ~n12421 & n13727;
  assign n13729 = ~n12440 & n13728;
  assign n13730 = ~n33884 & n13729;
  assign n13731 = n12426 & n12442;
  assign n13732 = ~n12434 & n13730;
  assign n13733 = ~n13719 & ~n34054;
  assign n13734 = ~n13097 & n13733;
  assign n13735 = ~n33974 & n13734;
  assign n13736 = ~n13091 & n13735;
  assign n13737 = n13099 & n13720;
  assign n13738 = ~n13717 & n13736;
  assign n13739 = n13726 & ~n34055;
  assign n13740 = ~n13721 & ~n13739;
  assign n13741 = ~n12442 & ~n13740;
  assign n13742 = n12442 & ~n13721;
  assign n13743 = ~n13739 & n13742;
  assign n13744 = ~n13099 & ~n13702;
  assign n13745 = ~n34050 & n13744;
  assign n13746 = ~n13696 & n13745;
  assign n13747 = ~n34053 & ~n13746;
  assign n13748 = pi46  & ~n13747;
  assign n13749 = ~pi46  & ~n13746;
  assign n13750 = ~pi46  & n13747;
  assign n13751 = ~n34053 & n13749;
  assign n13752 = ~n13748 & ~n34056;
  assign n13753 = ~n13743 & ~n13752;
  assign n13754 = ~n13741 & ~n13753;
  assign n13755 = ~n11858 & ~n13754;
  assign n13756 = n11858 & ~n13741;
  assign n13757 = ~n13753 & n13756;
  assign n13758 = n11858 & n13754;
  assign n13759 = ~n33986 & ~n13195;
  assign n13760 = ~n13704 & n13759;
  assign n13761 = n13193 & ~n13760;
  assign n13762 = ~n13193 & n13759;
  assign n13763 = ~n13193 & n13760;
  assign n13764 = ~n13704 & n13762;
  assign n13765 = ~n13761 & ~n34058;
  assign n13766 = ~n34057 & ~n13765;
  assign n13767 = ~n13755 & ~n13766;
  assign n13768 = ~n11229 & ~n13767;
  assign n13769 = n11229 & ~n13755;
  assign n13770 = ~n13766 & n13769;
  assign n13771 = ~n33987 & ~n13201;
  assign n13772 = ~n13201 & ~n13704;
  assign n13773 = ~n33987 & n13772;
  assign n13774 = ~n13704 & n13771;
  assign n13775 = n13175 & ~n34059;
  assign n13776 = n13200 & n13772;
  assign n13777 = n13175 & ~n33987;
  assign n13778 = ~n13201 & n13777;
  assign n13779 = ~n13704 & n13778;
  assign n13780 = ~n13175 & ~n34059;
  assign n13781 = ~n13779 & ~n13780;
  assign n13782 = ~n13775 & ~n13776;
  assign n13783 = ~n13770 & ~n34060;
  assign n13784 = ~n13768 & ~n13783;
  assign n13785 = ~n10681 & ~n13784;
  assign n13786 = n10681 & ~n13768;
  assign n13787 = ~n13783 & n13786;
  assign n13788 = n10681 & n13784;
  assign n13789 = ~n13203 & ~n13213;
  assign n13790 = ~n13704 & n13789;
  assign n13791 = n13210 & ~n13790;
  assign n13792 = ~n13210 & n13790;
  assign n13793 = n13210 & ~n13213;
  assign n13794 = ~n13203 & n13793;
  assign n13795 = n13210 & n13790;
  assign n13796 = ~n13704 & n13794;
  assign n13797 = ~n13210 & ~n13790;
  assign n13798 = ~n34062 & ~n13797;
  assign n13799 = ~n13791 & ~n13792;
  assign n13800 = ~n34061 & ~n34063;
  assign n13801 = ~n13785 & ~n13800;
  assign n13802 = ~n10086 & ~n13801;
  assign n13803 = n10086 & ~n13785;
  assign n13804 = ~n13800 & n13803;
  assign n13805 = ~n33989 & ~n13219;
  assign n13806 = ~n13219 & ~n13704;
  assign n13807 = ~n33989 & n13806;
  assign n13808 = ~n13704 & n13805;
  assign n13809 = n13163 & ~n34064;
  assign n13810 = n13218 & n13806;
  assign n13811 = n13163 & ~n33989;
  assign n13812 = ~n13219 & n13811;
  assign n13813 = ~n13704 & n13812;
  assign n13814 = ~n13163 & ~n34064;
  assign n13815 = ~n13813 & ~n13814;
  assign n13816 = ~n13809 & ~n13810;
  assign n13817 = ~n13804 & ~n34065;
  assign n13818 = ~n13802 & ~n13817;
  assign n13819 = ~n9565 & ~n13818;
  assign n13820 = n9565 & ~n13802;
  assign n13821 = ~n13817 & n13820;
  assign n13822 = n9565 & n13818;
  assign n13823 = ~n13221 & ~n13235;
  assign n13824 = ~n13704 & n13823;
  assign n13825 = ~n33991 & n13824;
  assign n13826 = n33991 & ~n13824;
  assign n13827 = n33991 & ~n13235;
  assign n13828 = ~n13221 & n13827;
  assign n13829 = ~n13704 & n13828;
  assign n13830 = ~n33991 & ~n13824;
  assign n13831 = ~n13829 & ~n13830;
  assign n13832 = ~n13825 & ~n13826;
  assign n13833 = ~n34066 & ~n34067;
  assign n13834 = ~n13819 & ~n13833;
  assign n13835 = ~n8998 & ~n13834;
  assign n13836 = n8998 & ~n13819;
  assign n13837 = ~n13833 & n13836;
  assign n13838 = ~n33992 & ~n13241;
  assign n13839 = ~n13241 & ~n13704;
  assign n13840 = ~n33992 & n13839;
  assign n13841 = ~n13704 & n13838;
  assign n13842 = n13155 & ~n34068;
  assign n13843 = n13240 & n13839;
  assign n13844 = n13155 & ~n33992;
  assign n13845 = ~n13241 & n13844;
  assign n13846 = ~n13704 & n13845;
  assign n13847 = ~n13155 & ~n34068;
  assign n13848 = ~n13846 & ~n13847;
  assign n13849 = ~n13842 & ~n13843;
  assign n13850 = ~n13837 & ~n34069;
  assign n13851 = ~n13835 & ~n13850;
  assign n13852 = ~n8506 & ~n13851;
  assign n13853 = n8506 & ~n13835;
  assign n13854 = ~n13850 & n13853;
  assign n13855 = n8506 & n13851;
  assign n13856 = ~n13243 & ~n13256;
  assign n13857 = ~n13704 & n13856;
  assign n13858 = ~n33993 & ~n13857;
  assign n13859 = n33993 & ~n13256;
  assign n13860 = ~n13243 & n13859;
  assign n13861 = n33993 & n13857;
  assign n13862 = ~n13704 & n13860;
  assign n13863 = n33993 & ~n13857;
  assign n13864 = ~n33993 & n13857;
  assign n13865 = ~n13863 & ~n13864;
  assign n13866 = ~n13858 & ~n34071;
  assign n13867 = ~n34070 & n34072;
  assign n13868 = ~n13852 & ~n13867;
  assign n13869 = ~n7975 & ~n13868;
  assign n13870 = n7975 & ~n13852;
  assign n13871 = ~n13867 & n13870;
  assign n13872 = ~n33994 & ~n13262;
  assign n13873 = ~n13262 & ~n13704;
  assign n13874 = ~n33994 & n13873;
  assign n13875 = ~n13704 & n13872;
  assign n13876 = n13147 & ~n34073;
  assign n13877 = n13261 & n13873;
  assign n13878 = n13147 & ~n33994;
  assign n13879 = ~n13262 & n13878;
  assign n13880 = ~n13704 & n13879;
  assign n13881 = ~n13147 & ~n34073;
  assign n13882 = ~n13880 & ~n13881;
  assign n13883 = ~n13876 & ~n13877;
  assign n13884 = ~n13871 & ~n34074;
  assign n13885 = ~n13869 & ~n13884;
  assign n13886 = ~n7512 & ~n13885;
  assign n13887 = n7512 & ~n13869;
  assign n13888 = ~n13884 & n13887;
  assign n13889 = n7512 & n13885;
  assign n13890 = ~n13264 & ~n13278;
  assign n13891 = ~n13704 & n13890;
  assign n13892 = n33996 & ~n13891;
  assign n13893 = ~n33996 & ~n13278;
  assign n13894 = ~n13264 & n13893;
  assign n13895 = ~n33996 & n13891;
  assign n13896 = ~n13704 & n13894;
  assign n13897 = n33996 & n13891;
  assign n13898 = ~n33996 & ~n13891;
  assign n13899 = ~n13897 & ~n13898;
  assign n13900 = ~n13892 & ~n34076;
  assign n13901 = ~n34075 & n34077;
  assign n13902 = ~n13886 & ~n13901;
  assign n13903 = ~n7015 & ~n13902;
  assign n13904 = n7015 & ~n13886;
  assign n13905 = ~n13901 & n13904;
  assign n13906 = ~n33997 & ~n13284;
  assign n13907 = ~n13284 & ~n13704;
  assign n13908 = ~n33997 & n13907;
  assign n13909 = ~n13704 & n13906;
  assign n13910 = n13139 & ~n34078;
  assign n13911 = n13283 & n13907;
  assign n13912 = n13139 & ~n33997;
  assign n13913 = ~n13284 & n13912;
  assign n13914 = ~n13704 & n13913;
  assign n13915 = ~n13139 & ~n34078;
  assign n13916 = ~n13914 & ~n13915;
  assign n13917 = ~n13910 & ~n13911;
  assign n13918 = ~n13905 & ~n34079;
  assign n13919 = ~n13903 & ~n13918;
  assign n13920 = ~n6579 & ~n13919;
  assign n13921 = n6579 & ~n13903;
  assign n13922 = ~n13918 & n13921;
  assign n13923 = n6579 & n13919;
  assign n13924 = ~n13286 & ~n13300;
  assign n13925 = ~n13300 & ~n13704;
  assign n13926 = ~n13286 & n13925;
  assign n13927 = ~n13704 & n13924;
  assign n13928 = ~n33999 & ~n34081;
  assign n13929 = n13298 & n13925;
  assign n13930 = n33999 & n34081;
  assign n13931 = ~n33999 & ~n13300;
  assign n13932 = ~n13286 & n13931;
  assign n13933 = ~n13704 & n13932;
  assign n13934 = n33999 & ~n34081;
  assign n13935 = ~n13933 & ~n13934;
  assign n13936 = ~n13928 & ~n34082;
  assign n13937 = ~n34080 & ~n34083;
  assign n13938 = ~n13920 & ~n13937;
  assign n13939 = ~n6117 & ~n13938;
  assign n13940 = n6117 & ~n13920;
  assign n13941 = ~n13937 & n13940;
  assign n13942 = ~n34000 & ~n13306;
  assign n13943 = ~n13306 & ~n13704;
  assign n13944 = ~n34000 & n13943;
  assign n13945 = ~n13704 & n13942;
  assign n13946 = n13131 & ~n34084;
  assign n13947 = n13305 & n13943;
  assign n13948 = n13131 & ~n34000;
  assign n13949 = ~n13306 & n13948;
  assign n13950 = ~n13704 & n13949;
  assign n13951 = ~n13131 & ~n34084;
  assign n13952 = ~n13950 & ~n13951;
  assign n13953 = ~n13946 & ~n13947;
  assign n13954 = ~n13941 & ~n34085;
  assign n13955 = ~n13939 & ~n13954;
  assign n13956 = ~n5708 & ~n13955;
  assign n13957 = n5708 & ~n13939;
  assign n13958 = ~n13954 & n13957;
  assign n13959 = n5708 & n13955;
  assign n13960 = ~n13308 & ~n13324;
  assign n13961 = ~n13704 & n13960;
  assign n13962 = ~n34003 & ~n13961;
  assign n13963 = n34003 & ~n13324;
  assign n13964 = ~n13308 & n13963;
  assign n13965 = n34003 & n13961;
  assign n13966 = ~n13704 & n13964;
  assign n13967 = ~n13962 & ~n34087;
  assign n13968 = ~n34086 & ~n13967;
  assign n13969 = ~n13956 & ~n13968;
  assign n13970 = ~n5278 & ~n13969;
  assign n13971 = n5278 & ~n13956;
  assign n13972 = ~n13968 & n13971;
  assign n13973 = ~n34004 & ~n13330;
  assign n13974 = ~n13330 & ~n13704;
  assign n13975 = ~n34004 & n13974;
  assign n13976 = ~n13704 & n13973;
  assign n13977 = n13123 & ~n34088;
  assign n13978 = n13329 & n13974;
  assign n13979 = n13123 & ~n34004;
  assign n13980 = ~n13330 & n13979;
  assign n13981 = ~n13704 & n13980;
  assign n13982 = ~n13123 & ~n34088;
  assign n13983 = ~n13981 & ~n13982;
  assign n13984 = ~n13977 & ~n13978;
  assign n13985 = ~n13972 & ~n34089;
  assign n13986 = ~n13970 & ~n13985;
  assign n13987 = ~n4903 & ~n13986;
  assign n13988 = n4903 & ~n13970;
  assign n13989 = ~n13985 & n13988;
  assign n13990 = n4903 & n13986;
  assign n13991 = ~n13332 & ~n13343;
  assign n13992 = ~n13343 & ~n13704;
  assign n13993 = ~n13332 & n13992;
  assign n13994 = ~n13704 & n13991;
  assign n13995 = n13340 & ~n34091;
  assign n13996 = n13341 & n13992;
  assign n13997 = ~n13340 & n34091;
  assign n13998 = n13340 & ~n13343;
  assign n13999 = ~n13332 & n13998;
  assign n14000 = ~n13704 & n13999;
  assign n14001 = ~n13340 & ~n34091;
  assign n14002 = ~n14000 & ~n14001;
  assign n14003 = ~n13995 & ~n34092;
  assign n14004 = ~n34090 & ~n34093;
  assign n14005 = ~n13987 & ~n14004;
  assign n14006 = ~n4508 & ~n14005;
  assign n14007 = n4508 & ~n13987;
  assign n14008 = ~n14004 & n14007;
  assign n14009 = n13115 & ~n34006;
  assign n14010 = ~n13349 & n14009;
  assign n14011 = ~n34006 & ~n13349;
  assign n14012 = ~n13704 & n14011;
  assign n14013 = n13115 & n14012;
  assign n14014 = ~n13704 & n14010;
  assign n14015 = ~n13115 & ~n14012;
  assign n14016 = ~n34094 & ~n14015;
  assign n14017 = ~n14008 & ~n14016;
  assign n14018 = ~n14006 & ~n14017;
  assign n14019 = ~n4155 & ~n14018;
  assign n14020 = n4155 & ~n14006;
  assign n14021 = ~n14017 & n14020;
  assign n14022 = n4155 & n14018;
  assign n14023 = ~n13351 & ~n13353;
  assign n14024 = ~n13704 & n14023;
  assign n14025 = ~n34008 & n14024;
  assign n14026 = n34008 & ~n14024;
  assign n14027 = ~n13351 & n34008;
  assign n14028 = ~n13353 & n14027;
  assign n14029 = n34008 & n14024;
  assign n14030 = ~n13704 & n14028;
  assign n14031 = ~n34008 & ~n14024;
  assign n14032 = ~n34096 & ~n14031;
  assign n14033 = ~n14025 & ~n14026;
  assign n14034 = ~n34095 & ~n34097;
  assign n14035 = ~n14019 & ~n14034;
  assign n14036 = ~n3788 & ~n14035;
  assign n14037 = n3788 & ~n14019;
  assign n14038 = ~n14034 & n14037;
  assign n14039 = ~n34052 & ~n14038;
  assign n14040 = ~n14036 & ~n14039;
  assign n14041 = ~n3473 & ~n14040;
  assign n14042 = ~n13373 & ~n13375;
  assign n14043 = ~n13704 & n14042;
  assign n14044 = ~n34011 & ~n14043;
  assign n14045 = ~n13373 & n34011;
  assign n14046 = ~n13375 & n14045;
  assign n14047 = n34011 & n14043;
  assign n14048 = ~n13704 & n14046;
  assign n14049 = ~n14044 & ~n34098;
  assign n14050 = n3473 & ~n14036;
  assign n14051 = ~n14039 & n14050;
  assign n14052 = n3473 & n14040;
  assign n14053 = ~n14049 & ~n34099;
  assign n14054 = ~n14041 & ~n14053;
  assign n14055 = ~n3140 & ~n14054;
  assign n14056 = n3140 & ~n14041;
  assign n14057 = ~n14053 & n14056;
  assign n14058 = ~n13390 & ~n34013;
  assign n14059 = ~n13390 & ~n13704;
  assign n14060 = ~n34013 & n14059;
  assign n14061 = ~n13704 & n14058;
  assign n14062 = n13398 & ~n34100;
  assign n14063 = n13402 & n14059;
  assign n14064 = n13398 & ~n34013;
  assign n14065 = ~n13390 & n14064;
  assign n14066 = ~n13704 & n14065;
  assign n14067 = ~n13398 & ~n34100;
  assign n14068 = ~n14066 & ~n14067;
  assign n14069 = ~n14062 & ~n14063;
  assign n14070 = ~n14057 & ~n34101;
  assign n14071 = ~n14055 & ~n14070;
  assign n14072 = ~n2855 & ~n14071;
  assign n14073 = ~n13404 & ~n13406;
  assign n14074 = ~n13704 & n14073;
  assign n14075 = ~n34016 & ~n14074;
  assign n14076 = ~n13404 & n34016;
  assign n14077 = ~n13406 & n14076;
  assign n14078 = n34016 & n14074;
  assign n14079 = ~n13704 & n14077;
  assign n14080 = ~n14075 & ~n34102;
  assign n14081 = n2855 & ~n14055;
  assign n14082 = ~n14070 & n14081;
  assign n14083 = n2855 & n14071;
  assign n14084 = ~n14080 & ~n34103;
  assign n14085 = ~n14072 & ~n14084;
  assign n14086 = ~n2556 & ~n14085;
  assign n14087 = n2556 & ~n14072;
  assign n14088 = ~n14084 & n14087;
  assign n14089 = ~n13422 & ~n34018;
  assign n14090 = ~n13422 & ~n13704;
  assign n14091 = ~n34018 & n14090;
  assign n14092 = ~n13704 & n14089;
  assign n14093 = n13430 & ~n34104;
  assign n14094 = n13434 & n14090;
  assign n14095 = n13430 & ~n34018;
  assign n14096 = ~n13422 & n14095;
  assign n14097 = ~n13704 & n14096;
  assign n14098 = ~n13430 & ~n34104;
  assign n14099 = ~n14097 & ~n14098;
  assign n14100 = ~n14093 & ~n14094;
  assign n14101 = ~n14088 & ~n34105;
  assign n14102 = ~n14086 & ~n14101;
  assign n14103 = ~n2301 & ~n14102;
  assign n14104 = n2301 & ~n14086;
  assign n14105 = ~n14101 & n14104;
  assign n14106 = n2301 & n14102;
  assign n14107 = ~n13436 & ~n13446;
  assign n14108 = ~n13436 & ~n13704;
  assign n14109 = ~n13446 & n14108;
  assign n14110 = ~n13704 & n14107;
  assign n14111 = n13444 & ~n34107;
  assign n14112 = n13447 & n14108;
  assign n14113 = ~n13436 & n13444;
  assign n14114 = ~n13446 & n14113;
  assign n14115 = ~n13704 & n14114;
  assign n14116 = ~n13444 & ~n34107;
  assign n14117 = ~n14115 & ~n14116;
  assign n14118 = ~n14111 & ~n14112;
  assign n14119 = ~n34106 & ~n34108;
  assign n14120 = ~n14103 & ~n14119;
  assign n14121 = ~n2038 & ~n14120;
  assign n14122 = n2038 & ~n14103;
  assign n14123 = ~n14119 & n14122;
  assign n14124 = ~n13449 & ~n34021;
  assign n14125 = ~n13449 & ~n13704;
  assign n14126 = ~n34021 & n14125;
  assign n14127 = ~n13704 & n14124;
  assign n14128 = n13457 & ~n34109;
  assign n14129 = n13461 & n14125;
  assign n14130 = n13457 & ~n34021;
  assign n14131 = ~n13449 & n14130;
  assign n14132 = ~n13704 & n14131;
  assign n14133 = ~n13457 & ~n34109;
  assign n14134 = ~n14132 & ~n14133;
  assign n14135 = ~n14128 & ~n14129;
  assign n14136 = ~n14123 & ~n34110;
  assign n14137 = ~n14121 & ~n14136;
  assign n14138 = ~n1812 & ~n14137;
  assign n14139 = ~n13463 & ~n13465;
  assign n14140 = ~n13704 & n14139;
  assign n14141 = ~n34023 & ~n14140;
  assign n14142 = ~n13463 & n34023;
  assign n14143 = ~n13465 & n14142;
  assign n14144 = n34023 & n14140;
  assign n14145 = ~n13704 & n14143;
  assign n14146 = ~n14141 & ~n34111;
  assign n14147 = n1812 & ~n14121;
  assign n14148 = ~n14136 & n14147;
  assign n14149 = n1812 & n14137;
  assign n14150 = ~n14146 & ~n34112;
  assign n14151 = ~n14138 & ~n14150;
  assign n14152 = ~n1582 & ~n14151;
  assign n14153 = n1582 & ~n14138;
  assign n14154 = ~n14150 & n14153;
  assign n14155 = ~n13480 & ~n34025;
  assign n14156 = ~n13480 & ~n13704;
  assign n14157 = ~n34025 & n14156;
  assign n14158 = ~n13704 & n14155;
  assign n14159 = n13488 & ~n34113;
  assign n14160 = n13492 & n14156;
  assign n14161 = n13488 & ~n34025;
  assign n14162 = ~n13480 & n14161;
  assign n14163 = ~n13704 & n14162;
  assign n14164 = ~n13488 & ~n34113;
  assign n14165 = ~n14163 & ~n14164;
  assign n14166 = ~n14159 & ~n14160;
  assign n14167 = ~n14154 & ~n34114;
  assign n14168 = ~n14152 & ~n14167;
  assign n14169 = ~n1388 & ~n14168;
  assign n14170 = n1388 & ~n14152;
  assign n14171 = ~n14167 & n14170;
  assign n14172 = n1388 & n14168;
  assign n14173 = ~n13494 & ~n13504;
  assign n14174 = ~n13494 & ~n13704;
  assign n14175 = ~n13504 & n14174;
  assign n14176 = ~n13704 & n14173;
  assign n14177 = n13502 & ~n34116;
  assign n14178 = n13505 & n14174;
  assign n14179 = ~n13494 & n13502;
  assign n14180 = ~n13504 & n14179;
  assign n14181 = ~n13704 & n14180;
  assign n14182 = ~n13502 & ~n34116;
  assign n14183 = ~n14181 & ~n14182;
  assign n14184 = ~n14177 & ~n14178;
  assign n14185 = ~n34115 & ~n34117;
  assign n14186 = ~n14169 & ~n14185;
  assign n14187 = ~n1192 & ~n14186;
  assign n14188 = n1192 & ~n14169;
  assign n14189 = ~n14185 & n14188;
  assign n14190 = ~n13507 & ~n34028;
  assign n14191 = ~n13507 & ~n13704;
  assign n14192 = ~n34028 & n14191;
  assign n14193 = ~n13704 & n14190;
  assign n14194 = n13515 & ~n34118;
  assign n14195 = n13519 & n14191;
  assign n14196 = n13515 & ~n34028;
  assign n14197 = ~n13507 & n14196;
  assign n14198 = ~n13704 & n14197;
  assign n14199 = ~n13515 & ~n34118;
  assign n14200 = ~n14198 & ~n14199;
  assign n14201 = ~n14194 & ~n14195;
  assign n14202 = ~n14189 & ~n34119;
  assign n14203 = ~n14187 & ~n14202;
  assign n14204 = ~n1028 & ~n14203;
  assign n14205 = ~n13521 & ~n13523;
  assign n14206 = ~n13704 & n14205;
  assign n14207 = ~n34030 & ~n14206;
  assign n14208 = ~n13521 & n34030;
  assign n14209 = ~n13523 & n14208;
  assign n14210 = n34030 & n14206;
  assign n14211 = ~n13704 & n14209;
  assign n14212 = ~n14207 & ~n34120;
  assign n14213 = n1028 & ~n14187;
  assign n14214 = ~n14202 & n14213;
  assign n14215 = n1028 & n14203;
  assign n14216 = ~n14212 & ~n34121;
  assign n14217 = ~n14204 & ~n14216;
  assign n14218 = ~n866 & ~n14217;
  assign n14219 = n866 & ~n14204;
  assign n14220 = ~n14216 & n14219;
  assign n14221 = ~n13538 & ~n34032;
  assign n14222 = ~n13538 & ~n13704;
  assign n14223 = ~n34032 & n14222;
  assign n14224 = ~n13704 & n14221;
  assign n14225 = n13546 & ~n34122;
  assign n14226 = n13550 & n14222;
  assign n14227 = n13546 & ~n34032;
  assign n14228 = ~n13538 & n14227;
  assign n14229 = ~n13704 & n14228;
  assign n14230 = ~n13546 & ~n34122;
  assign n14231 = ~n14229 & ~n14230;
  assign n14232 = ~n14225 & ~n14226;
  assign n14233 = ~n14220 & ~n34123;
  assign n14234 = ~n14218 & ~n14233;
  assign n14235 = ~n730 & ~n14234;
  assign n14236 = n730 & ~n14218;
  assign n14237 = ~n14233 & n14236;
  assign n14238 = n730 & n14234;
  assign n14239 = ~n13552 & ~n13562;
  assign n14240 = ~n13552 & ~n13704;
  assign n14241 = ~n13562 & n14240;
  assign n14242 = ~n13704 & n14239;
  assign n14243 = n13560 & ~n34125;
  assign n14244 = n13563 & n14240;
  assign n14245 = ~n13552 & n13560;
  assign n14246 = ~n13562 & n14245;
  assign n14247 = ~n13704 & n14246;
  assign n14248 = ~n13560 & ~n34125;
  assign n14249 = ~n14247 & ~n14248;
  assign n14250 = ~n14243 & ~n14244;
  assign n14251 = ~n34124 & ~n34126;
  assign n14252 = ~n14235 & ~n14251;
  assign n14253 = ~n602 & ~n14252;
  assign n14254 = n602 & ~n14235;
  assign n14255 = ~n14251 & n14254;
  assign n14256 = ~n13565 & ~n34035;
  assign n14257 = ~n13565 & ~n13704;
  assign n14258 = ~n34035 & n14257;
  assign n14259 = ~n13704 & n14256;
  assign n14260 = n13573 & ~n34127;
  assign n14261 = n13577 & n14257;
  assign n14262 = n13573 & ~n34035;
  assign n14263 = ~n13565 & n14262;
  assign n14264 = ~n13704 & n14263;
  assign n14265 = ~n13573 & ~n34127;
  assign n14266 = ~n14264 & ~n14265;
  assign n14267 = ~n14260 & ~n14261;
  assign n14268 = ~n14255 & ~n34128;
  assign n14269 = ~n14253 & ~n14268;
  assign n14270 = ~n497 & ~n14269;
  assign n14271 = ~n13579 & ~n13581;
  assign n14272 = ~n13704 & n14271;
  assign n14273 = ~n34037 & ~n14272;
  assign n14274 = ~n13579 & n34037;
  assign n14275 = ~n13581 & n14274;
  assign n14276 = n34037 & n14272;
  assign n14277 = ~n13704 & n14275;
  assign n14278 = ~n14273 & ~n34129;
  assign n14279 = n497 & ~n14253;
  assign n14280 = ~n14268 & n14279;
  assign n14281 = n497 & n14269;
  assign n14282 = ~n14278 & ~n34130;
  assign n14283 = ~n14270 & ~n14282;
  assign n14284 = ~n403 & ~n14283;
  assign n14285 = n403 & ~n14270;
  assign n14286 = ~n14282 & n14285;
  assign n14287 = ~n13596 & ~n34039;
  assign n14288 = ~n13596 & ~n13704;
  assign n14289 = ~n34039 & n14288;
  assign n14290 = ~n13704 & n14287;
  assign n14291 = n13604 & ~n34131;
  assign n14292 = n13608 & n14288;
  assign n14293 = n13604 & ~n34039;
  assign n14294 = ~n13596 & n14293;
  assign n14295 = ~n13704 & n14294;
  assign n14296 = ~n13604 & ~n34131;
  assign n14297 = ~n14295 & ~n14296;
  assign n14298 = ~n14291 & ~n14292;
  assign n14299 = ~n14286 & ~n34132;
  assign n14300 = ~n14284 & ~n14299;
  assign n14301 = ~n330 & ~n14300;
  assign n14302 = n330 & ~n14284;
  assign n14303 = ~n14299 & n14302;
  assign n14304 = n330 & n14300;
  assign n14305 = ~n13610 & ~n13620;
  assign n14306 = ~n13610 & ~n13704;
  assign n14307 = ~n13620 & n14306;
  assign n14308 = ~n13704 & n14305;
  assign n14309 = n13618 & ~n34134;
  assign n14310 = n13621 & n14306;
  assign n14311 = ~n13610 & n13618;
  assign n14312 = ~n13620 & n14311;
  assign n14313 = ~n13704 & n14312;
  assign n14314 = ~n13618 & ~n34134;
  assign n14315 = ~n14313 & ~n14314;
  assign n14316 = ~n14309 & ~n14310;
  assign n14317 = ~n34133 & ~n34135;
  assign n14318 = ~n14301 & ~n14317;
  assign n14319 = ~n271 & ~n14318;
  assign n14320 = n271 & ~n14301;
  assign n14321 = ~n14317 & n14320;
  assign n14322 = ~n13623 & ~n34042;
  assign n14323 = ~n13623 & ~n13704;
  assign n14324 = ~n34042 & n14323;
  assign n14325 = ~n13704 & n14322;
  assign n14326 = n13631 & ~n34136;
  assign n14327 = n13635 & n14323;
  assign n14328 = n13631 & ~n34042;
  assign n14329 = ~n13623 & n14328;
  assign n14330 = ~n13704 & n14329;
  assign n14331 = ~n13631 & ~n34136;
  assign n14332 = ~n14330 & ~n14331;
  assign n14333 = ~n14326 & ~n14327;
  assign n14334 = ~n14321 & ~n34137;
  assign n14335 = ~n14319 & ~n14334;
  assign n14336 = ~n217 & ~n14335;
  assign n14337 = ~n13637 & ~n13639;
  assign n14338 = ~n13704 & n14337;
  assign n14339 = ~n34044 & ~n14338;
  assign n14340 = ~n13637 & n34044;
  assign n14341 = ~n13639 & n14340;
  assign n14342 = n34044 & n14338;
  assign n14343 = ~n13704 & n14341;
  assign n14344 = ~n14339 & ~n34138;
  assign n14345 = n217 & ~n14319;
  assign n14346 = ~n14334 & n14345;
  assign n14347 = n217 & n14335;
  assign n14348 = ~n14344 & ~n34139;
  assign n14349 = ~n14336 & ~n14348;
  assign n14350 = ~n198 & ~n14349;
  assign n14351 = n198 & ~n14336;
  assign n14352 = ~n14348 & n14351;
  assign n14353 = ~n13654 & ~n34046;
  assign n14354 = ~n13654 & ~n13704;
  assign n14355 = ~n34046 & n14354;
  assign n14356 = ~n13704 & n14353;
  assign n14357 = n13662 & ~n34140;
  assign n14358 = n13666 & n14354;
  assign n14359 = n13662 & ~n34046;
  assign n14360 = ~n13654 & n14359;
  assign n14361 = ~n13704 & n14360;
  assign n14362 = ~n13662 & ~n34140;
  assign n14363 = ~n14361 & ~n14362;
  assign n14364 = ~n14357 & ~n14358;
  assign n14365 = ~n14352 & ~n34141;
  assign n14366 = ~n14350 & ~n14365;
  assign n14367 = ~n13668 & ~n13678;
  assign n14368 = ~n13668 & ~n13704;
  assign n14369 = ~n13678 & n14368;
  assign n14370 = ~n13704 & n14367;
  assign n14371 = n13676 & ~n34142;
  assign n14372 = n13679 & n14368;
  assign n14373 = ~n13668 & n13676;
  assign n14374 = ~n13678 & n14373;
  assign n14375 = ~n13704 & n14374;
  assign n14376 = ~n13676 & ~n34142;
  assign n14377 = ~n14375 & ~n14376;
  assign n14378 = ~n14371 & ~n14372;
  assign n14379 = ~n13680 & ~n13688;
  assign n14380 = ~n13688 & ~n13704;
  assign n14381 = ~n13680 & n14380;
  assign n14382 = ~n13704 & n14379;
  assign n14383 = ~n34050 & ~n34144;
  assign n14384 = ~n34143 & n14383;
  assign n14385 = ~n14366 & n14384;
  assign n14386 = n193 & ~n14385;
  assign n14387 = ~n14350 & n34143;
  assign n14388 = ~n14365 & n14387;
  assign n14389 = n14366 & n34143;
  assign n14390 = n13680 & ~n14380;
  assign n14391 = ~n193 & ~n14379;
  assign n14392 = ~n14390 & n14391;
  assign n14393 = ~n34145 & ~n14392;
  assign n14394 = ~n14386 & n14393;
  assign n14395 = ~n14036 & ~n14038;
  assign n14396 = ~n14394 & n14395;
  assign n14397 = ~n34052 & ~n14396;
  assign n14398 = n34052 & ~n14038;
  assign n14399 = ~n14036 & n14398;
  assign n14400 = n34052 & n14396;
  assign n14401 = ~n14394 & n14399;
  assign n14402 = ~n14397 & ~n34146;
  assign n14403 = ~n14006 & ~n14008;
  assign n14404 = ~n14394 & n14403;
  assign n14405 = ~n14016 & ~n14404;
  assign n14406 = ~n14008 & n14016;
  assign n14407 = ~n14006 & n14406;
  assign n14408 = n14016 & n14404;
  assign n14409 = ~n14394 & n14407;
  assign n14410 = ~n14405 & ~n34147;
  assign n14411 = ~n13970 & ~n13972;
  assign n14412 = ~n14394 & n14411;
  assign n14413 = ~n34089 & ~n14412;
  assign n14414 = ~n13972 & n34089;
  assign n14415 = ~n13970 & n14414;
  assign n14416 = n34089 & n14412;
  assign n14417 = ~n14394 & n14415;
  assign n14418 = ~n14413 & ~n34148;
  assign n14419 = ~n13939 & ~n13941;
  assign n14420 = ~n14394 & n14419;
  assign n14421 = ~n34085 & ~n14420;
  assign n14422 = ~n13941 & n34085;
  assign n14423 = ~n13939 & n14422;
  assign n14424 = n34085 & n14420;
  assign n14425 = ~n14394 & n14423;
  assign n14426 = ~n14421 & ~n34149;
  assign n14427 = ~n13903 & ~n13905;
  assign n14428 = ~n14394 & n14427;
  assign n14429 = ~n34079 & ~n14428;
  assign n14430 = ~n13905 & n34079;
  assign n14431 = ~n13903 & n14430;
  assign n14432 = n34079 & n14428;
  assign n14433 = ~n14394 & n14431;
  assign n14434 = ~n14429 & ~n34150;
  assign n14435 = ~n13869 & ~n13871;
  assign n14436 = ~n14394 & n14435;
  assign n14437 = ~n34074 & ~n14436;
  assign n14438 = ~n13871 & n34074;
  assign n14439 = ~n13869 & n14438;
  assign n14440 = n34074 & n14436;
  assign n14441 = ~n14394 & n14439;
  assign n14442 = ~n14437 & ~n34151;
  assign n14443 = ~n13835 & ~n13837;
  assign n14444 = ~n14394 & n14443;
  assign n14445 = ~n34069 & ~n14444;
  assign n14446 = ~n13837 & n34069;
  assign n14447 = ~n13835 & n14446;
  assign n14448 = n34069 & n14444;
  assign n14449 = ~n14394 & n14447;
  assign n14450 = ~n14445 & ~n34152;
  assign n14451 = ~n13802 & ~n13804;
  assign n14452 = ~n14394 & n14451;
  assign n14453 = ~n34065 & ~n14452;
  assign n14454 = ~n13804 & n34065;
  assign n14455 = ~n13802 & n14454;
  assign n14456 = n34065 & n14452;
  assign n14457 = ~n14394 & n14455;
  assign n14458 = ~n14453 & ~n34153;
  assign n14459 = ~n13768 & ~n13770;
  assign n14460 = ~n14394 & n14459;
  assign n14461 = ~n34060 & ~n14460;
  assign n14462 = ~n13770 & n34060;
  assign n14463 = ~n13768 & n14462;
  assign n14464 = n34060 & n14460;
  assign n14465 = ~n14394 & n14463;
  assign n14466 = ~n14461 & ~n34154;
  assign n14467 = ~n13741 & ~n13743;
  assign n14468 = ~n14394 & n14467;
  assign n14469 = ~n13752 & ~n14468;
  assign n14470 = ~n13743 & n13752;
  assign n14471 = ~n13741 & n14470;
  assign n14472 = n13752 & n14468;
  assign n14473 = ~n14394 & n14471;
  assign n14474 = ~n14469 & ~n34155;
  assign n14475 = ~pi42  & ~n14394;
  assign n14476 = ~pi43  & n14475;
  assign n14477 = n13718 & ~n14394;
  assign n14478 = ~n13704 & ~n14392;
  assign n14479 = ~n34145 & n14478;
  assign n14480 = ~n14386 & n14479;
  assign n14481 = ~n34156 & ~n14480;
  assign n14482 = pi44  & ~n14481;
  assign n14483 = ~pi44  & ~n14480;
  assign n14484 = ~pi44  & n14481;
  assign n14485 = ~n34156 & n14483;
  assign n14486 = ~n14482 & ~n34157;
  assign n14487 = pi42  & ~n14394;
  assign n14488 = ~pi40  & ~pi41 ;
  assign n14489 = ~pi42  & n14488;
  assign n14490 = ~n33972 & ~n34054;
  assign n14491 = ~n13078 & n14490;
  assign n14492 = ~n13097 & n14491;
  assign n14493 = ~n33974 & n14492;
  assign n14494 = n13083 & n13099;
  assign n14495 = ~n13091 & n14493;
  assign n14496 = ~n14489 & ~n34158;
  assign n14497 = ~n13702 & n14496;
  assign n14498 = ~n34050 & n14497;
  assign n14499 = ~n13696 & n14498;
  assign n14500 = ~n14487 & ~n14489;
  assign n14501 = n13704 & n14500;
  assign n14502 = ~n14487 & n14499;
  assign n14503 = pi43  & ~n14475;
  assign n14504 = ~n34156 & ~n14503;
  assign n14505 = ~n34159 & n14504;
  assign n14506 = ~n13704 & ~n14500;
  assign n14507 = n13099 & ~n14506;
  assign n14508 = ~n14505 & ~n14506;
  assign n14509 = n13099 & n14508;
  assign n14510 = ~n14505 & n14507;
  assign n14511 = ~n14486 & ~n34160;
  assign n14512 = ~n13099 & ~n14508;
  assign n14513 = n12442 & ~n14512;
  assign n14514 = ~n14511 & n14513;
  assign n14515 = ~n13721 & ~n34055;
  assign n14516 = ~n14394 & n14515;
  assign n14517 = n13726 & ~n14516;
  assign n14518 = ~n13726 & n14515;
  assign n14519 = ~n13726 & n14516;
  assign n14520 = ~n14394 & n14518;
  assign n14521 = ~n14517 & ~n34161;
  assign n14522 = ~n14514 & ~n14521;
  assign n14523 = ~n14511 & ~n14512;
  assign n14524 = ~n12442 & ~n14523;
  assign n14525 = n11858 & ~n14524;
  assign n14526 = ~n14522 & ~n14524;
  assign n14527 = n11858 & n14526;
  assign n14528 = ~n14522 & n14525;
  assign n14529 = ~n14474 & ~n34162;
  assign n14530 = ~n11858 & ~n14526;
  assign n14531 = n11229 & ~n14530;
  assign n14532 = ~n14529 & n14531;
  assign n14533 = ~n13755 & ~n34057;
  assign n14534 = ~n14394 & n14533;
  assign n14535 = n13765 & ~n14534;
  assign n14536 = ~n13765 & n14534;
  assign n14537 = ~n13755 & n13765;
  assign n14538 = ~n34057 & n14537;
  assign n14539 = n13765 & n14534;
  assign n14540 = ~n14394 & n14538;
  assign n14541 = ~n13765 & ~n14534;
  assign n14542 = ~n34163 & ~n14541;
  assign n14543 = ~n14535 & ~n14536;
  assign n14544 = ~n14532 & ~n34164;
  assign n14545 = ~n14529 & ~n14530;
  assign n14546 = ~n11229 & ~n14545;
  assign n14547 = n10681 & ~n14546;
  assign n14548 = ~n14544 & ~n14546;
  assign n14549 = n10681 & n14548;
  assign n14550 = ~n14544 & n14547;
  assign n14551 = ~n14466 & ~n34165;
  assign n14552 = ~n10681 & ~n14548;
  assign n14553 = n10086 & ~n14552;
  assign n14554 = ~n14551 & n14553;
  assign n14555 = ~n13785 & ~n34061;
  assign n14556 = ~n14394 & n14555;
  assign n14557 = ~n34063 & n14556;
  assign n14558 = n34063 & ~n14556;
  assign n14559 = ~n13785 & n34063;
  assign n14560 = ~n34061 & n14559;
  assign n14561 = ~n14394 & n14560;
  assign n14562 = ~n34063 & ~n14556;
  assign n14563 = ~n14561 & ~n14562;
  assign n14564 = ~n14557 & ~n14558;
  assign n14565 = ~n14554 & ~n34166;
  assign n14566 = ~n14551 & ~n14552;
  assign n14567 = ~n10086 & ~n14566;
  assign n14568 = n9565 & ~n14567;
  assign n14569 = ~n14565 & ~n14567;
  assign n14570 = n9565 & n14569;
  assign n14571 = ~n14565 & n14568;
  assign n14572 = ~n14458 & ~n34167;
  assign n14573 = ~n9565 & ~n14569;
  assign n14574 = n8998 & ~n14573;
  assign n14575 = ~n14572 & n14574;
  assign n14576 = ~n13819 & ~n34066;
  assign n14577 = ~n14394 & n14576;
  assign n14578 = ~n34067 & ~n14577;
  assign n14579 = ~n13819 & n34067;
  assign n14580 = ~n34066 & n14579;
  assign n14581 = n34067 & n14577;
  assign n14582 = ~n14394 & n14580;
  assign n14583 = n34067 & ~n14577;
  assign n14584 = ~n34067 & n14577;
  assign n14585 = ~n14583 & ~n14584;
  assign n14586 = ~n14578 & ~n34168;
  assign n14587 = ~n14575 & n34169;
  assign n14588 = ~n14572 & ~n14573;
  assign n14589 = ~n8998 & ~n14588;
  assign n14590 = n8506 & ~n14589;
  assign n14591 = ~n14587 & ~n14589;
  assign n14592 = n8506 & n14591;
  assign n14593 = ~n14587 & n14590;
  assign n14594 = ~n14450 & ~n34170;
  assign n14595 = ~n8506 & ~n14591;
  assign n14596 = n7975 & ~n14595;
  assign n14597 = ~n14594 & n14596;
  assign n14598 = ~n13852 & ~n34070;
  assign n14599 = ~n14394 & n14598;
  assign n14600 = n34072 & ~n14599;
  assign n14601 = ~n13852 & ~n34072;
  assign n14602 = ~n34070 & n14601;
  assign n14603 = ~n34072 & n14599;
  assign n14604 = ~n14394 & n14602;
  assign n14605 = n34072 & n14599;
  assign n14606 = ~n34072 & ~n14599;
  assign n14607 = ~n14605 & ~n14606;
  assign n14608 = ~n14600 & ~n34171;
  assign n14609 = ~n14597 & n34172;
  assign n14610 = ~n14594 & ~n14595;
  assign n14611 = ~n7975 & ~n14610;
  assign n14612 = n7512 & ~n14611;
  assign n14613 = ~n14609 & ~n14611;
  assign n14614 = n7512 & n14613;
  assign n14615 = ~n14609 & n14612;
  assign n14616 = ~n14442 & ~n34173;
  assign n14617 = ~n7512 & ~n14613;
  assign n14618 = n7015 & ~n14617;
  assign n14619 = ~n14616 & n14618;
  assign n14620 = ~n13886 & ~n34075;
  assign n14621 = ~n13886 & ~n14394;
  assign n14622 = ~n34075 & n14621;
  assign n14623 = ~n14394 & n14620;
  assign n14624 = ~n34077 & ~n34174;
  assign n14625 = n13901 & n14621;
  assign n14626 = n34077 & n34174;
  assign n14627 = ~n13886 & ~n34077;
  assign n14628 = ~n34075 & n14627;
  assign n14629 = ~n14394 & n14628;
  assign n14630 = n34077 & ~n34174;
  assign n14631 = ~n14629 & ~n14630;
  assign n14632 = ~n14624 & ~n34175;
  assign n14633 = ~n14619 & ~n34176;
  assign n14634 = ~n14616 & ~n14617;
  assign n14635 = ~n7015 & ~n14634;
  assign n14636 = n6579 & ~n14635;
  assign n14637 = ~n14633 & ~n14635;
  assign n14638 = n6579 & n14637;
  assign n14639 = ~n14633 & n14636;
  assign n14640 = ~n14434 & ~n34177;
  assign n14641 = ~n6579 & ~n14637;
  assign n14642 = n6117 & ~n14641;
  assign n14643 = ~n14640 & n14642;
  assign n14644 = ~n13920 & ~n34080;
  assign n14645 = ~n14394 & n14644;
  assign n14646 = ~n34083 & ~n14645;
  assign n14647 = ~n13920 & n34083;
  assign n14648 = ~n34080 & n14647;
  assign n14649 = n34083 & n14645;
  assign n14650 = ~n14394 & n14648;
  assign n14651 = ~n14646 & ~n34178;
  assign n14652 = ~n14643 & ~n14651;
  assign n14653 = ~n14640 & ~n14641;
  assign n14654 = ~n6117 & ~n14653;
  assign n14655 = n5708 & ~n14654;
  assign n14656 = ~n14652 & ~n14654;
  assign n14657 = n5708 & n14656;
  assign n14658 = ~n14652 & n14655;
  assign n14659 = ~n14426 & ~n34179;
  assign n14660 = ~n5708 & ~n14656;
  assign n14661 = n5278 & ~n14660;
  assign n14662 = ~n14659 & n14661;
  assign n14663 = ~n13956 & ~n34086;
  assign n14664 = ~n13956 & ~n14394;
  assign n14665 = ~n34086 & n14664;
  assign n14666 = ~n14394 & n14663;
  assign n14667 = n13967 & ~n34180;
  assign n14668 = n13968 & n14664;
  assign n14669 = ~n13967 & n34180;
  assign n14670 = ~n13956 & n13967;
  assign n14671 = ~n34086 & n14670;
  assign n14672 = ~n14394 & n14671;
  assign n14673 = ~n13967 & ~n34180;
  assign n14674 = ~n14672 & ~n14673;
  assign n14675 = ~n14667 & ~n34181;
  assign n14676 = ~n14662 & ~n34182;
  assign n14677 = ~n14659 & ~n14660;
  assign n14678 = ~n5278 & ~n14677;
  assign n14679 = n4903 & ~n14678;
  assign n14680 = ~n14676 & ~n14678;
  assign n14681 = n4903 & n14680;
  assign n14682 = ~n14676 & n14679;
  assign n14683 = ~n14418 & ~n34183;
  assign n14684 = ~n4903 & ~n14680;
  assign n14685 = n4508 & ~n14684;
  assign n14686 = ~n14683 & n14685;
  assign n14687 = ~n13987 & ~n34090;
  assign n14688 = ~n14394 & n14687;
  assign n14689 = ~n34093 & n14688;
  assign n14690 = n34093 & ~n14688;
  assign n14691 = ~n13987 & n34093;
  assign n14692 = ~n34090 & n14691;
  assign n14693 = n34093 & n14688;
  assign n14694 = ~n14394 & n14692;
  assign n14695 = ~n34093 & ~n14688;
  assign n14696 = ~n34184 & ~n14695;
  assign n14697 = ~n14689 & ~n14690;
  assign n14698 = ~n14686 & ~n34185;
  assign n14699 = ~n14683 & ~n14684;
  assign n14700 = ~n4508 & ~n14699;
  assign n14701 = n4155 & ~n14700;
  assign n14702 = ~n14698 & ~n14700;
  assign n14703 = n4155 & n14702;
  assign n14704 = ~n14698 & n14701;
  assign n14705 = ~n14410 & ~n34186;
  assign n14706 = ~n4155 & ~n14702;
  assign n14707 = ~n14705 & ~n14706;
  assign n14708 = ~n3788 & ~n14707;
  assign n14709 = n3788 & ~n14706;
  assign n14710 = ~n14705 & n14709;
  assign n14711 = ~n14019 & ~n34095;
  assign n14712 = ~n14394 & n14711;
  assign n14713 = ~n34097 & ~n14712;
  assign n14714 = ~n14019 & n34097;
  assign n14715 = ~n34095 & n14714;
  assign n14716 = n34097 & n14712;
  assign n14717 = ~n14394 & n14715;
  assign n14718 = n34097 & ~n14712;
  assign n14719 = ~n34097 & n14712;
  assign n14720 = ~n14718 & ~n14719;
  assign n14721 = ~n14713 & ~n34187;
  assign n14722 = ~n14710 & n34188;
  assign n14723 = ~n14708 & ~n14722;
  assign n14724 = ~n3473 & ~n14723;
  assign n14725 = n3473 & ~n14708;
  assign n14726 = n3473 & n14723;
  assign n14727 = ~n14722 & n14725;
  assign n14728 = ~n14402 & ~n34189;
  assign n14729 = ~n14724 & ~n14728;
  assign n14730 = ~n3140 & ~n14729;
  assign n14731 = n3140 & ~n14724;
  assign n14732 = ~n14728 & n14731;
  assign n14733 = ~n14041 & ~n34099;
  assign n14734 = ~n14041 & ~n14394;
  assign n14735 = ~n34099 & n14734;
  assign n14736 = ~n14394 & n14733;
  assign n14737 = n14049 & ~n34190;
  assign n14738 = n14053 & n14734;
  assign n14739 = ~n14041 & n14049;
  assign n14740 = ~n34099 & n14739;
  assign n14741 = ~n14394 & n14740;
  assign n14742 = ~n14049 & ~n34190;
  assign n14743 = ~n14741 & ~n14742;
  assign n14744 = ~n14737 & ~n14738;
  assign n14745 = ~n14732 & ~n34191;
  assign n14746 = ~n14730 & ~n14745;
  assign n14747 = ~n2855 & ~n14746;
  assign n14748 = ~n14055 & ~n14057;
  assign n14749 = ~n14394 & n14748;
  assign n14750 = ~n34101 & ~n14749;
  assign n14751 = ~n14057 & n34101;
  assign n14752 = ~n14055 & n14751;
  assign n14753 = n34101 & n14749;
  assign n14754 = ~n14394 & n14752;
  assign n14755 = ~n14750 & ~n34192;
  assign n14756 = n2855 & ~n14730;
  assign n14757 = n2855 & n14746;
  assign n14758 = ~n14745 & n14756;
  assign n14759 = ~n14755 & ~n34193;
  assign n14760 = ~n14747 & ~n14759;
  assign n14761 = ~n2556 & ~n14760;
  assign n14762 = n2556 & ~n14747;
  assign n14763 = ~n14759 & n14762;
  assign n14764 = ~n14072 & ~n34103;
  assign n14765 = ~n14072 & ~n14394;
  assign n14766 = ~n34103 & n14765;
  assign n14767 = ~n14394 & n14764;
  assign n14768 = n14080 & ~n34194;
  assign n14769 = n14084 & n14765;
  assign n14770 = ~n14072 & n14080;
  assign n14771 = ~n34103 & n14770;
  assign n14772 = ~n14394 & n14771;
  assign n14773 = ~n14080 & ~n34194;
  assign n14774 = ~n14772 & ~n14773;
  assign n14775 = ~n14768 & ~n14769;
  assign n14776 = ~n14763 & ~n34195;
  assign n14777 = ~n14761 & ~n14776;
  assign n14778 = ~n2301 & ~n14777;
  assign n14779 = ~n14086 & ~n14088;
  assign n14780 = ~n14394 & n14779;
  assign n14781 = ~n34105 & ~n14780;
  assign n14782 = ~n14088 & n34105;
  assign n14783 = ~n14086 & n14782;
  assign n14784 = n34105 & n14780;
  assign n14785 = ~n14394 & n14783;
  assign n14786 = ~n14781 & ~n34196;
  assign n14787 = n2301 & ~n14761;
  assign n14788 = n2301 & n14777;
  assign n14789 = ~n14776 & n14787;
  assign n14790 = ~n14786 & ~n34197;
  assign n14791 = ~n14778 & ~n14790;
  assign n14792 = ~n2038 & ~n14791;
  assign n14793 = ~n14103 & ~n34106;
  assign n14794 = ~n14394 & n14793;
  assign n14795 = ~n34108 & ~n14794;
  assign n14796 = ~n14103 & n34108;
  assign n14797 = ~n34106 & n14796;
  assign n14798 = n34108 & n14794;
  assign n14799 = ~n14394 & n14797;
  assign n14800 = ~n14795 & ~n34198;
  assign n14801 = n2038 & ~n14778;
  assign n14802 = ~n14790 & n14801;
  assign n14803 = ~n14800 & ~n14802;
  assign n14804 = ~n14792 & ~n14803;
  assign n14805 = ~n1812 & ~n14804;
  assign n14806 = ~n14121 & ~n14123;
  assign n14807 = ~n14394 & n14806;
  assign n14808 = ~n34110 & ~n14807;
  assign n14809 = ~n14123 & n34110;
  assign n14810 = ~n14121 & n14809;
  assign n14811 = n34110 & n14807;
  assign n14812 = ~n14394 & n14810;
  assign n14813 = ~n14808 & ~n34199;
  assign n14814 = n1812 & ~n14792;
  assign n14815 = n1812 & n14804;
  assign n14816 = ~n14803 & n14814;
  assign n14817 = ~n14813 & ~n34200;
  assign n14818 = ~n14805 & ~n14817;
  assign n14819 = ~n1582 & ~n14818;
  assign n14820 = n1582 & ~n14805;
  assign n14821 = ~n14817 & n14820;
  assign n14822 = ~n14138 & ~n34112;
  assign n14823 = ~n14138 & ~n14394;
  assign n14824 = ~n34112 & n14823;
  assign n14825 = ~n14394 & n14822;
  assign n14826 = n14146 & ~n34201;
  assign n14827 = n14150 & n14823;
  assign n14828 = ~n14138 & n14146;
  assign n14829 = ~n34112 & n14828;
  assign n14830 = ~n14394 & n14829;
  assign n14831 = ~n14146 & ~n34201;
  assign n14832 = ~n14830 & ~n14831;
  assign n14833 = ~n14826 & ~n14827;
  assign n14834 = ~n14821 & ~n34202;
  assign n14835 = ~n14819 & ~n14834;
  assign n14836 = ~n1388 & ~n14835;
  assign n14837 = ~n14152 & ~n14154;
  assign n14838 = ~n14394 & n14837;
  assign n14839 = ~n34114 & ~n14838;
  assign n14840 = ~n14154 & n34114;
  assign n14841 = ~n14152 & n14840;
  assign n14842 = n34114 & n14838;
  assign n14843 = ~n14394 & n14841;
  assign n14844 = ~n14839 & ~n34203;
  assign n14845 = n1388 & ~n14819;
  assign n14846 = n1388 & n14835;
  assign n14847 = ~n14834 & n14845;
  assign n14848 = ~n14844 & ~n34204;
  assign n14849 = ~n14836 & ~n14848;
  assign n14850 = ~n1192 & ~n14849;
  assign n14851 = ~n14169 & ~n34115;
  assign n14852 = ~n14394 & n14851;
  assign n14853 = ~n34117 & ~n14852;
  assign n14854 = ~n14169 & n34117;
  assign n14855 = ~n34115 & n14854;
  assign n14856 = n34117 & n14852;
  assign n14857 = ~n14394 & n14855;
  assign n14858 = ~n14853 & ~n34205;
  assign n14859 = n1192 & ~n14836;
  assign n14860 = ~n14848 & n14859;
  assign n14861 = ~n14858 & ~n14860;
  assign n14862 = ~n14850 & ~n14861;
  assign n14863 = ~n1028 & ~n14862;
  assign n14864 = ~n14187 & ~n14189;
  assign n14865 = ~n14394 & n14864;
  assign n14866 = ~n34119 & ~n14865;
  assign n14867 = ~n14189 & n34119;
  assign n14868 = ~n14187 & n14867;
  assign n14869 = n34119 & n14865;
  assign n14870 = ~n14394 & n14868;
  assign n14871 = ~n14866 & ~n34206;
  assign n14872 = n1028 & ~n14850;
  assign n14873 = n1028 & n14862;
  assign n14874 = ~n14861 & n14872;
  assign n14875 = ~n14871 & ~n34207;
  assign n14876 = ~n14863 & ~n14875;
  assign n14877 = ~n866 & ~n14876;
  assign n14878 = n866 & ~n14863;
  assign n14879 = ~n14875 & n14878;
  assign n14880 = ~n14204 & ~n34121;
  assign n14881 = ~n14204 & ~n14394;
  assign n14882 = ~n34121 & n14881;
  assign n14883 = ~n14394 & n14880;
  assign n14884 = n14212 & ~n34208;
  assign n14885 = n14216 & n14881;
  assign n14886 = ~n14204 & n14212;
  assign n14887 = ~n34121 & n14886;
  assign n14888 = ~n14394 & n14887;
  assign n14889 = ~n14212 & ~n34208;
  assign n14890 = ~n14888 & ~n14889;
  assign n14891 = ~n14884 & ~n14885;
  assign n14892 = ~n14879 & ~n34209;
  assign n14893 = ~n14877 & ~n14892;
  assign n14894 = ~n730 & ~n14893;
  assign n14895 = ~n14218 & ~n14220;
  assign n14896 = ~n14394 & n14895;
  assign n14897 = ~n34123 & ~n14896;
  assign n14898 = ~n14220 & n34123;
  assign n14899 = ~n14218 & n14898;
  assign n14900 = n34123 & n14896;
  assign n14901 = ~n14394 & n14899;
  assign n14902 = ~n14897 & ~n34210;
  assign n14903 = n730 & ~n14877;
  assign n14904 = n730 & n14893;
  assign n14905 = ~n14892 & n14903;
  assign n14906 = ~n14902 & ~n34211;
  assign n14907 = ~n14894 & ~n14906;
  assign n14908 = ~n602 & ~n14907;
  assign n14909 = ~n14235 & ~n34124;
  assign n14910 = ~n14394 & n14909;
  assign n14911 = ~n34126 & ~n14910;
  assign n14912 = ~n14235 & n34126;
  assign n14913 = ~n34124 & n14912;
  assign n14914 = n34126 & n14910;
  assign n14915 = ~n14394 & n14913;
  assign n14916 = ~n14911 & ~n34212;
  assign n14917 = n602 & ~n14894;
  assign n14918 = ~n14906 & n14917;
  assign n14919 = ~n14916 & ~n14918;
  assign n14920 = ~n14908 & ~n14919;
  assign n14921 = ~n497 & ~n14920;
  assign n14922 = ~n14253 & ~n14255;
  assign n14923 = ~n14394 & n14922;
  assign n14924 = ~n34128 & ~n14923;
  assign n14925 = ~n14255 & n34128;
  assign n14926 = ~n14253 & n14925;
  assign n14927 = n34128 & n14923;
  assign n14928 = ~n14394 & n14926;
  assign n14929 = ~n14924 & ~n34213;
  assign n14930 = n497 & ~n14908;
  assign n14931 = n497 & n14920;
  assign n14932 = ~n14919 & n14930;
  assign n14933 = ~n14929 & ~n34214;
  assign n14934 = ~n14921 & ~n14933;
  assign n14935 = ~n403 & ~n14934;
  assign n14936 = n403 & ~n14921;
  assign n14937 = ~n14933 & n14936;
  assign n14938 = ~n14270 & ~n34130;
  assign n14939 = ~n14270 & ~n14394;
  assign n14940 = ~n34130 & n14939;
  assign n14941 = ~n14394 & n14938;
  assign n14942 = n14278 & ~n34215;
  assign n14943 = n14282 & n14939;
  assign n14944 = ~n14270 & n14278;
  assign n14945 = ~n34130 & n14944;
  assign n14946 = ~n14394 & n14945;
  assign n14947 = ~n14278 & ~n34215;
  assign n14948 = ~n14946 & ~n14947;
  assign n14949 = ~n14942 & ~n14943;
  assign n14950 = ~n14937 & ~n34216;
  assign n14951 = ~n14935 & ~n14950;
  assign n14952 = ~n330 & ~n14951;
  assign n14953 = ~n14284 & ~n14286;
  assign n14954 = ~n14394 & n14953;
  assign n14955 = ~n34132 & ~n14954;
  assign n14956 = ~n14286 & n34132;
  assign n14957 = ~n14284 & n14956;
  assign n14958 = n34132 & n14954;
  assign n14959 = ~n14394 & n14957;
  assign n14960 = ~n14955 & ~n34217;
  assign n14961 = n330 & ~n14935;
  assign n14962 = n330 & n14951;
  assign n14963 = ~n14950 & n14961;
  assign n14964 = ~n14960 & ~n34218;
  assign n14965 = ~n14952 & ~n14964;
  assign n14966 = ~n271 & ~n14965;
  assign n14967 = ~n14301 & ~n34133;
  assign n14968 = ~n14394 & n14967;
  assign n14969 = ~n34135 & ~n14968;
  assign n14970 = ~n14301 & n34135;
  assign n14971 = ~n34133 & n14970;
  assign n14972 = n34135 & n14968;
  assign n14973 = ~n14394 & n14971;
  assign n14974 = ~n14969 & ~n34219;
  assign n14975 = n271 & ~n14952;
  assign n14976 = ~n14964 & n14975;
  assign n14977 = ~n14974 & ~n14976;
  assign n14978 = ~n14966 & ~n14977;
  assign n14979 = ~n217 & ~n14978;
  assign n14980 = ~n14319 & ~n14321;
  assign n14981 = ~n14394 & n14980;
  assign n14982 = ~n34137 & ~n14981;
  assign n14983 = ~n14321 & n34137;
  assign n14984 = ~n14319 & n14983;
  assign n14985 = n34137 & n14981;
  assign n14986 = ~n14394 & n14984;
  assign n14987 = ~n14982 & ~n34220;
  assign n14988 = n217 & ~n14966;
  assign n14989 = n217 & n14978;
  assign n14990 = ~n14977 & n14988;
  assign n14991 = ~n14987 & ~n34221;
  assign n14992 = ~n14979 & ~n14991;
  assign n14993 = ~n198 & ~n14992;
  assign n14994 = n198 & ~n14979;
  assign n14995 = ~n14991 & n14994;
  assign n14996 = ~n14336 & ~n34139;
  assign n14997 = ~n14336 & ~n14394;
  assign n14998 = ~n34139 & n14997;
  assign n14999 = ~n14394 & n14996;
  assign n15000 = n14344 & ~n34222;
  assign n15001 = n14348 & n14997;
  assign n15002 = ~n14336 & n14344;
  assign n15003 = ~n34139 & n15002;
  assign n15004 = ~n14394 & n15003;
  assign n15005 = ~n14344 & ~n34222;
  assign n15006 = ~n15004 & ~n15005;
  assign n15007 = ~n15000 & ~n15001;
  assign n15008 = ~n14995 & ~n34223;
  assign n15009 = ~n14993 & ~n15008;
  assign n15010 = ~n14350 & ~n14352;
  assign n15011 = ~n14394 & n15010;
  assign n15012 = ~n34141 & ~n15011;
  assign n15013 = ~n14352 & n34141;
  assign n15014 = ~n14350 & n15013;
  assign n15015 = n34141 & n15011;
  assign n15016 = ~n14394 & n15014;
  assign n15017 = ~n15012 & ~n34224;
  assign n15018 = ~n14366 & ~n34143;
  assign n15019 = ~n34143 & ~n14394;
  assign n15020 = ~n14366 & n15019;
  assign n15021 = ~n14394 & n15018;
  assign n15022 = ~n34145 & ~n34225;
  assign n15023 = ~n15017 & n15022;
  assign n15024 = ~n15009 & n15023;
  assign n15025 = n193 & ~n15024;
  assign n15026 = ~n14993 & n15017;
  assign n15027 = n15009 & n15017;
  assign n15028 = ~n15008 & n15026;
  assign n15029 = n14366 & ~n15019;
  assign n15030 = ~n193 & ~n15018;
  assign n15031 = ~n15029 & n15030;
  assign n15032 = ~n34226 & ~n15031;
  assign n15033 = ~n15025 & n15032;
  assign n15034 = ~n14724 & ~n34189;
  assign n15035 = ~n14724 & ~n15033;
  assign n15036 = ~n34189 & n15035;
  assign n15037 = ~n15033 & n15034;
  assign n15038 = n14402 & ~n34227;
  assign n15039 = n14728 & n15035;
  assign n15040 = n14402 & ~n34189;
  assign n15041 = ~n14724 & n15040;
  assign n15042 = ~n15033 & n15041;
  assign n15043 = ~n14402 & ~n34227;
  assign n15044 = ~n15042 & ~n15043;
  assign n15045 = ~n15038 & ~n15039;
  assign n15046 = pi40  & ~n15033;
  assign n15047 = ~pi38  & ~pi39 ;
  assign n15048 = ~pi40  & n15047;
  assign n15049 = ~n15046 & ~n15048;
  assign n15050 = ~n14394 & ~n15049;
  assign n15051 = ~pi40  & ~n15033;
  assign n15052 = pi41  & ~n15051;
  assign n15053 = ~pi41  & n15051;
  assign n15054 = n14488 & ~n15033;
  assign n15055 = ~n15052 & ~n34229;
  assign n15056 = ~n34048 & ~n34158;
  assign n15057 = ~n13683 & n15056;
  assign n15058 = ~n13702 & n15057;
  assign n15059 = ~n34050 & n15058;
  assign n15060 = n13688 & n13704;
  assign n15061 = ~n13696 & n15059;
  assign n15062 = ~n15048 & ~n34230;
  assign n15063 = ~n14392 & n15062;
  assign n15064 = ~n34145 & n15063;
  assign n15065 = ~n14386 & n15064;
  assign n15066 = n14394 & n15049;
  assign n15067 = ~n15046 & n15065;
  assign n15068 = n15055 & ~n34231;
  assign n15069 = ~n15050 & ~n15068;
  assign n15070 = ~n13704 & ~n15069;
  assign n15071 = n13704 & ~n15050;
  assign n15072 = ~n15068 & n15071;
  assign n15073 = ~n14394 & ~n15031;
  assign n15074 = ~n34226 & n15073;
  assign n15075 = ~n15025 & n15074;
  assign n15076 = ~n34229 & ~n15075;
  assign n15077 = pi42  & ~n15076;
  assign n15078 = ~pi42  & ~n15075;
  assign n15079 = ~pi42  & n15076;
  assign n15080 = ~n34229 & n15078;
  assign n15081 = ~n15077 & ~n34232;
  assign n15082 = ~n15072 & ~n15081;
  assign n15083 = ~n15070 & ~n15082;
  assign n15084 = ~n13099 & ~n15083;
  assign n15085 = n13099 & ~n15070;
  assign n15086 = ~n15082 & n15085;
  assign n15087 = n13099 & n15083;
  assign n15088 = ~n34159 & ~n14506;
  assign n15089 = ~n15033 & n15088;
  assign n15090 = n14504 & ~n15089;
  assign n15091 = ~n14504 & n15088;
  assign n15092 = ~n14504 & n15089;
  assign n15093 = ~n15033 & n15091;
  assign n15094 = ~n15090 & ~n34234;
  assign n15095 = ~n34233 & ~n15094;
  assign n15096 = ~n15084 & ~n15095;
  assign n15097 = ~n12442 & ~n15096;
  assign n15098 = n12442 & ~n15084;
  assign n15099 = ~n15095 & n15098;
  assign n15100 = ~n34160 & ~n14512;
  assign n15101 = ~n14512 & ~n15033;
  assign n15102 = ~n34160 & n15101;
  assign n15103 = ~n15033 & n15100;
  assign n15104 = n14486 & ~n34235;
  assign n15105 = n14511 & n15101;
  assign n15106 = n14486 & ~n34160;
  assign n15107 = ~n14512 & n15106;
  assign n15108 = ~n15033 & n15107;
  assign n15109 = ~n14486 & ~n34235;
  assign n15110 = ~n15108 & ~n15109;
  assign n15111 = ~n15104 & ~n15105;
  assign n15112 = ~n15099 & ~n34236;
  assign n15113 = ~n15097 & ~n15112;
  assign n15114 = ~n11858 & ~n15113;
  assign n15115 = n11858 & ~n15097;
  assign n15116 = ~n15112 & n15115;
  assign n15117 = n11858 & n15113;
  assign n15118 = ~n14514 & ~n14524;
  assign n15119 = ~n15033 & n15118;
  assign n15120 = n14521 & ~n15119;
  assign n15121 = ~n14521 & n15119;
  assign n15122 = n14521 & ~n14524;
  assign n15123 = ~n14514 & n15122;
  assign n15124 = n14521 & n15119;
  assign n15125 = ~n15033 & n15123;
  assign n15126 = ~n14521 & ~n15119;
  assign n15127 = ~n34238 & ~n15126;
  assign n15128 = ~n15120 & ~n15121;
  assign n15129 = ~n34237 & ~n34239;
  assign n15130 = ~n15114 & ~n15129;
  assign n15131 = ~n11229 & ~n15130;
  assign n15132 = n11229 & ~n15114;
  assign n15133 = ~n15129 & n15132;
  assign n15134 = ~n34162 & ~n14530;
  assign n15135 = ~n14530 & ~n15033;
  assign n15136 = ~n34162 & n15135;
  assign n15137 = ~n15033 & n15134;
  assign n15138 = n14474 & ~n34240;
  assign n15139 = n14529 & n15135;
  assign n15140 = n14474 & ~n34162;
  assign n15141 = ~n14530 & n15140;
  assign n15142 = ~n15033 & n15141;
  assign n15143 = ~n14474 & ~n34240;
  assign n15144 = ~n15142 & ~n15143;
  assign n15145 = ~n15138 & ~n15139;
  assign n15146 = ~n15133 & ~n34241;
  assign n15147 = ~n15131 & ~n15146;
  assign n15148 = ~n10681 & ~n15147;
  assign n15149 = n10681 & ~n15131;
  assign n15150 = ~n15146 & n15149;
  assign n15151 = n10681 & n15147;
  assign n15152 = ~n14532 & ~n14546;
  assign n15153 = ~n15033 & n15152;
  assign n15154 = ~n34164 & n15153;
  assign n15155 = n34164 & ~n15153;
  assign n15156 = n34164 & ~n14546;
  assign n15157 = ~n14532 & n15156;
  assign n15158 = ~n15033 & n15157;
  assign n15159 = ~n34164 & ~n15153;
  assign n15160 = ~n15158 & ~n15159;
  assign n15161 = ~n15154 & ~n15155;
  assign n15162 = ~n34242 & ~n34243;
  assign n15163 = ~n15148 & ~n15162;
  assign n15164 = ~n10086 & ~n15163;
  assign n15165 = n10086 & ~n15148;
  assign n15166 = ~n15162 & n15165;
  assign n15167 = ~n34165 & ~n14552;
  assign n15168 = ~n14552 & ~n15033;
  assign n15169 = ~n34165 & n15168;
  assign n15170 = ~n15033 & n15167;
  assign n15171 = n14466 & ~n34244;
  assign n15172 = n14551 & n15168;
  assign n15173 = n14466 & ~n34165;
  assign n15174 = ~n14552 & n15173;
  assign n15175 = ~n15033 & n15174;
  assign n15176 = ~n14466 & ~n34244;
  assign n15177 = ~n15175 & ~n15176;
  assign n15178 = ~n15171 & ~n15172;
  assign n15179 = ~n15166 & ~n34245;
  assign n15180 = ~n15164 & ~n15179;
  assign n15181 = ~n9565 & ~n15180;
  assign n15182 = n9565 & ~n15164;
  assign n15183 = ~n15179 & n15182;
  assign n15184 = n9565 & n15180;
  assign n15185 = ~n14554 & ~n14567;
  assign n15186 = ~n15033 & n15185;
  assign n15187 = ~n34166 & ~n15186;
  assign n15188 = n34166 & ~n14567;
  assign n15189 = ~n14554 & n15188;
  assign n15190 = n34166 & n15186;
  assign n15191 = ~n15033 & n15189;
  assign n15192 = n34166 & ~n15186;
  assign n15193 = ~n34166 & n15186;
  assign n15194 = ~n15192 & ~n15193;
  assign n15195 = ~n15187 & ~n34247;
  assign n15196 = ~n34246 & n34248;
  assign n15197 = ~n15181 & ~n15196;
  assign n15198 = ~n8998 & ~n15197;
  assign n15199 = n8998 & ~n15181;
  assign n15200 = ~n15196 & n15199;
  assign n15201 = ~n34167 & ~n14573;
  assign n15202 = ~n14573 & ~n15033;
  assign n15203 = ~n34167 & n15202;
  assign n15204 = ~n15033 & n15201;
  assign n15205 = n14458 & ~n34249;
  assign n15206 = n14572 & n15202;
  assign n15207 = n14458 & ~n34167;
  assign n15208 = ~n14573 & n15207;
  assign n15209 = ~n15033 & n15208;
  assign n15210 = ~n14458 & ~n34249;
  assign n15211 = ~n15209 & ~n15210;
  assign n15212 = ~n15205 & ~n15206;
  assign n15213 = ~n15200 & ~n34250;
  assign n15214 = ~n15198 & ~n15213;
  assign n15215 = ~n8506 & ~n15214;
  assign n15216 = n8506 & ~n15198;
  assign n15217 = ~n15213 & n15216;
  assign n15218 = n8506 & n15214;
  assign n15219 = ~n14575 & ~n14589;
  assign n15220 = ~n15033 & n15219;
  assign n15221 = n34169 & ~n15220;
  assign n15222 = ~n34169 & ~n14589;
  assign n15223 = ~n14575 & n15222;
  assign n15224 = ~n34169 & n15220;
  assign n15225 = ~n15033 & n15223;
  assign n15226 = n34169 & n15220;
  assign n15227 = ~n34169 & ~n15220;
  assign n15228 = ~n15226 & ~n15227;
  assign n15229 = ~n15221 & ~n34252;
  assign n15230 = ~n34251 & n34253;
  assign n15231 = ~n15215 & ~n15230;
  assign n15232 = ~n7975 & ~n15231;
  assign n15233 = n7975 & ~n15215;
  assign n15234 = ~n15230 & n15233;
  assign n15235 = ~n34170 & ~n14595;
  assign n15236 = ~n14595 & ~n15033;
  assign n15237 = ~n34170 & n15236;
  assign n15238 = ~n15033 & n15235;
  assign n15239 = n14450 & ~n34254;
  assign n15240 = n14594 & n15236;
  assign n15241 = n14450 & ~n34170;
  assign n15242 = ~n14595 & n15241;
  assign n15243 = ~n15033 & n15242;
  assign n15244 = ~n14450 & ~n34254;
  assign n15245 = ~n15243 & ~n15244;
  assign n15246 = ~n15239 & ~n15240;
  assign n15247 = ~n15234 & ~n34255;
  assign n15248 = ~n15232 & ~n15247;
  assign n15249 = ~n7512 & ~n15248;
  assign n15250 = n7512 & ~n15232;
  assign n15251 = ~n15247 & n15250;
  assign n15252 = n7512 & n15248;
  assign n15253 = ~n14597 & ~n14611;
  assign n15254 = ~n14611 & ~n15033;
  assign n15255 = ~n14597 & n15254;
  assign n15256 = ~n15033 & n15253;
  assign n15257 = ~n34172 & ~n34257;
  assign n15258 = n14609 & n15254;
  assign n15259 = n34172 & n34257;
  assign n15260 = ~n34172 & ~n14611;
  assign n15261 = ~n14597 & n15260;
  assign n15262 = ~n15033 & n15261;
  assign n15263 = n34172 & ~n34257;
  assign n15264 = ~n15262 & ~n15263;
  assign n15265 = ~n15257 & ~n34258;
  assign n15266 = ~n34256 & ~n34259;
  assign n15267 = ~n15249 & ~n15266;
  assign n15268 = ~n7015 & ~n15267;
  assign n15269 = n7015 & ~n15249;
  assign n15270 = ~n15266 & n15269;
  assign n15271 = ~n34173 & ~n14617;
  assign n15272 = ~n14617 & ~n15033;
  assign n15273 = ~n34173 & n15272;
  assign n15274 = ~n15033 & n15271;
  assign n15275 = n14442 & ~n34260;
  assign n15276 = n14616 & n15272;
  assign n15277 = n14442 & ~n34173;
  assign n15278 = ~n14617 & n15277;
  assign n15279 = ~n15033 & n15278;
  assign n15280 = ~n14442 & ~n34260;
  assign n15281 = ~n15279 & ~n15280;
  assign n15282 = ~n15275 & ~n15276;
  assign n15283 = ~n15270 & ~n34261;
  assign n15284 = ~n15268 & ~n15283;
  assign n15285 = ~n6579 & ~n15284;
  assign n15286 = n6579 & ~n15268;
  assign n15287 = ~n15283 & n15286;
  assign n15288 = n6579 & n15284;
  assign n15289 = ~n14619 & ~n14635;
  assign n15290 = ~n15033 & n15289;
  assign n15291 = ~n34176 & ~n15290;
  assign n15292 = n34176 & ~n14635;
  assign n15293 = ~n14619 & n15292;
  assign n15294 = n34176 & n15290;
  assign n15295 = ~n15033 & n15293;
  assign n15296 = ~n15291 & ~n34263;
  assign n15297 = ~n34262 & ~n15296;
  assign n15298 = ~n15285 & ~n15297;
  assign n15299 = ~n6117 & ~n15298;
  assign n15300 = n6117 & ~n15285;
  assign n15301 = ~n15297 & n15300;
  assign n15302 = ~n34177 & ~n14641;
  assign n15303 = ~n14641 & ~n15033;
  assign n15304 = ~n34177 & n15303;
  assign n15305 = ~n15033 & n15302;
  assign n15306 = n14434 & ~n34264;
  assign n15307 = n14640 & n15303;
  assign n15308 = n14434 & ~n34177;
  assign n15309 = ~n14641 & n15308;
  assign n15310 = ~n15033 & n15309;
  assign n15311 = ~n14434 & ~n34264;
  assign n15312 = ~n15310 & ~n15311;
  assign n15313 = ~n15306 & ~n15307;
  assign n15314 = ~n15301 & ~n34265;
  assign n15315 = ~n15299 & ~n15314;
  assign n15316 = ~n5708 & ~n15315;
  assign n15317 = n5708 & ~n15299;
  assign n15318 = ~n15314 & n15317;
  assign n15319 = n5708 & n15315;
  assign n15320 = ~n14643 & ~n14654;
  assign n15321 = ~n14654 & ~n15033;
  assign n15322 = ~n14643 & n15321;
  assign n15323 = ~n15033 & n15320;
  assign n15324 = n14651 & ~n34267;
  assign n15325 = n14652 & n15321;
  assign n15326 = ~n14651 & n34267;
  assign n15327 = n14651 & ~n14654;
  assign n15328 = ~n14643 & n15327;
  assign n15329 = ~n15033 & n15328;
  assign n15330 = ~n14651 & ~n34267;
  assign n15331 = ~n15329 & ~n15330;
  assign n15332 = ~n15324 & ~n34268;
  assign n15333 = ~n34266 & ~n34269;
  assign n15334 = ~n15316 & ~n15333;
  assign n15335 = ~n5278 & ~n15334;
  assign n15336 = n5278 & ~n15316;
  assign n15337 = ~n15333 & n15336;
  assign n15338 = ~n34179 & ~n14660;
  assign n15339 = ~n14660 & ~n15033;
  assign n15340 = ~n34179 & n15339;
  assign n15341 = ~n15033 & n15338;
  assign n15342 = n14426 & ~n34270;
  assign n15343 = n14659 & n15339;
  assign n15344 = n14426 & ~n34179;
  assign n15345 = ~n14660 & n15344;
  assign n15346 = ~n15033 & n15345;
  assign n15347 = ~n14426 & ~n34270;
  assign n15348 = ~n15346 & ~n15347;
  assign n15349 = ~n15342 & ~n15343;
  assign n15350 = ~n15337 & ~n34271;
  assign n15351 = ~n15335 & ~n15350;
  assign n15352 = ~n4903 & ~n15351;
  assign n15353 = n4903 & ~n15335;
  assign n15354 = ~n15350 & n15353;
  assign n15355 = n4903 & n15351;
  assign n15356 = ~n14662 & ~n14678;
  assign n15357 = ~n15033 & n15356;
  assign n15358 = ~n34182 & n15357;
  assign n15359 = n34182 & ~n15357;
  assign n15360 = n34182 & ~n14678;
  assign n15361 = ~n14662 & n15360;
  assign n15362 = n34182 & n15357;
  assign n15363 = ~n15033 & n15361;
  assign n15364 = ~n34182 & ~n15357;
  assign n15365 = ~n34273 & ~n15364;
  assign n15366 = ~n15358 & ~n15359;
  assign n15367 = ~n34272 & ~n34274;
  assign n15368 = ~n15352 & ~n15367;
  assign n15369 = ~n4508 & ~n15368;
  assign n15370 = n4508 & ~n15352;
  assign n15371 = ~n15367 & n15370;
  assign n15372 = ~n34183 & ~n14684;
  assign n15373 = ~n14684 & ~n15033;
  assign n15374 = ~n34183 & n15373;
  assign n15375 = ~n15033 & n15372;
  assign n15376 = n14418 & ~n34275;
  assign n15377 = n14683 & n15373;
  assign n15378 = n14418 & ~n34183;
  assign n15379 = ~n14684 & n15378;
  assign n15380 = ~n15033 & n15379;
  assign n15381 = ~n14418 & ~n34275;
  assign n15382 = ~n15380 & ~n15381;
  assign n15383 = ~n15376 & ~n15377;
  assign n15384 = ~n15371 & ~n34276;
  assign n15385 = ~n15369 & ~n15384;
  assign n15386 = ~n4155 & ~n15385;
  assign n15387 = n4155 & ~n15369;
  assign n15388 = ~n15384 & n15387;
  assign n15389 = n4155 & n15385;
  assign n15390 = ~n14686 & ~n14700;
  assign n15391 = ~n14700 & ~n15033;
  assign n15392 = ~n14686 & n15391;
  assign n15393 = ~n15033 & n15390;
  assign n15394 = n34185 & ~n34278;
  assign n15395 = n14698 & n15391;
  assign n15396 = ~n34185 & n34278;
  assign n15397 = n34185 & ~n14700;
  assign n15398 = ~n14686 & n15397;
  assign n15399 = ~n15033 & n15398;
  assign n15400 = ~n34185 & ~n34278;
  assign n15401 = ~n15399 & ~n15400;
  assign n15402 = ~n15394 & ~n34279;
  assign n15403 = ~n34277 & ~n34280;
  assign n15404 = ~n15386 & ~n15403;
  assign n15405 = ~n3788 & ~n15404;
  assign n15406 = n3788 & ~n15386;
  assign n15407 = ~n15403 & n15406;
  assign n15408 = ~n34186 & ~n14706;
  assign n15409 = ~n15033 & n15408;
  assign n15410 = n14410 & ~n15409;
  assign n15411 = ~n14410 & n15409;
  assign n15412 = n14410 & ~n34186;
  assign n15413 = ~n14706 & n15412;
  assign n15414 = ~n15033 & n15413;
  assign n15415 = ~n14410 & ~n15409;
  assign n15416 = ~n15414 & ~n15415;
  assign n15417 = ~n15410 & ~n15411;
  assign n15418 = ~n15407 & ~n34281;
  assign n15419 = ~n15405 & ~n15418;
  assign n15420 = ~n3473 & ~n15419;
  assign n15421 = ~n14708 & ~n14710;
  assign n15422 = ~n15033 & n15421;
  assign n15423 = n34188 & ~n15422;
  assign n15424 = ~n14708 & ~n34188;
  assign n15425 = ~n14710 & n15424;
  assign n15426 = ~n34188 & n15422;
  assign n15427 = ~n15033 & n15425;
  assign n15428 = n34188 & n15422;
  assign n15429 = ~n34188 & ~n15422;
  assign n15430 = ~n15428 & ~n15429;
  assign n15431 = ~n15423 & ~n34282;
  assign n15432 = n3473 & ~n15405;
  assign n15433 = ~n15418 & n15432;
  assign n15434 = n3473 & n15419;
  assign n15435 = n34283 & ~n34284;
  assign n15436 = ~n15420 & ~n15435;
  assign n15437 = ~n3140 & ~n15436;
  assign n15438 = n3140 & ~n15420;
  assign n15439 = ~n15435 & n15438;
  assign n15440 = ~n34228 & ~n15439;
  assign n15441 = ~n15437 & ~n15440;
  assign n15442 = ~n2855 & ~n15441;
  assign n15443 = ~n14730 & ~n14732;
  assign n15444 = ~n15033 & n15443;
  assign n15445 = ~n34191 & ~n15444;
  assign n15446 = ~n14730 & n34191;
  assign n15447 = ~n14732 & n15446;
  assign n15448 = n34191 & n15444;
  assign n15449 = ~n15033 & n15447;
  assign n15450 = ~n15445 & ~n34285;
  assign n15451 = n2855 & ~n15437;
  assign n15452 = ~n15440 & n15451;
  assign n15453 = n2855 & n15441;
  assign n15454 = ~n15450 & ~n34286;
  assign n15455 = ~n15442 & ~n15454;
  assign n15456 = ~n2556 & ~n15455;
  assign n15457 = n2556 & ~n15442;
  assign n15458 = ~n15454 & n15457;
  assign n15459 = ~n14747 & ~n34193;
  assign n15460 = ~n14747 & ~n15033;
  assign n15461 = ~n34193 & n15460;
  assign n15462 = ~n15033 & n15459;
  assign n15463 = n14755 & ~n34287;
  assign n15464 = n14759 & n15460;
  assign n15465 = n14755 & ~n34193;
  assign n15466 = ~n14747 & n15465;
  assign n15467 = ~n15033 & n15466;
  assign n15468 = ~n14755 & ~n34287;
  assign n15469 = ~n15467 & ~n15468;
  assign n15470 = ~n15463 & ~n15464;
  assign n15471 = ~n15458 & ~n34288;
  assign n15472 = ~n15456 & ~n15471;
  assign n15473 = ~n2301 & ~n15472;
  assign n15474 = ~n14761 & ~n14763;
  assign n15475 = ~n15033 & n15474;
  assign n15476 = ~n34195 & ~n15475;
  assign n15477 = ~n14761 & n34195;
  assign n15478 = ~n14763 & n15477;
  assign n15479 = n34195 & n15475;
  assign n15480 = ~n15033 & n15478;
  assign n15481 = ~n15476 & ~n34289;
  assign n15482 = n2301 & ~n15456;
  assign n15483 = ~n15471 & n15482;
  assign n15484 = n2301 & n15472;
  assign n15485 = ~n15481 & ~n34290;
  assign n15486 = ~n15473 & ~n15485;
  assign n15487 = ~n2038 & ~n15486;
  assign n15488 = n2038 & ~n15473;
  assign n15489 = ~n15485 & n15488;
  assign n15490 = ~n14778 & ~n34197;
  assign n15491 = ~n14778 & ~n15033;
  assign n15492 = ~n34197 & n15491;
  assign n15493 = ~n15033 & n15490;
  assign n15494 = n14786 & ~n34291;
  assign n15495 = n14790 & n15491;
  assign n15496 = n14786 & ~n34197;
  assign n15497 = ~n14778 & n15496;
  assign n15498 = ~n15033 & n15497;
  assign n15499 = ~n14786 & ~n34291;
  assign n15500 = ~n15498 & ~n15499;
  assign n15501 = ~n15494 & ~n15495;
  assign n15502 = ~n15489 & ~n34292;
  assign n15503 = ~n15487 & ~n15502;
  assign n15504 = ~n1812 & ~n15503;
  assign n15505 = n1812 & ~n15487;
  assign n15506 = ~n15502 & n15505;
  assign n15507 = n1812 & n15503;
  assign n15508 = ~n14792 & ~n14802;
  assign n15509 = ~n14792 & ~n15033;
  assign n15510 = ~n14802 & n15509;
  assign n15511 = ~n15033 & n15508;
  assign n15512 = n14800 & ~n34294;
  assign n15513 = n14803 & n15509;
  assign n15514 = ~n14792 & n14800;
  assign n15515 = ~n14802 & n15514;
  assign n15516 = ~n15033 & n15515;
  assign n15517 = ~n14800 & ~n34294;
  assign n15518 = ~n15516 & ~n15517;
  assign n15519 = ~n15512 & ~n15513;
  assign n15520 = ~n34293 & ~n34295;
  assign n15521 = ~n15504 & ~n15520;
  assign n15522 = ~n1582 & ~n15521;
  assign n15523 = n1582 & ~n15504;
  assign n15524 = ~n15520 & n15523;
  assign n15525 = ~n14805 & ~n34200;
  assign n15526 = ~n14805 & ~n15033;
  assign n15527 = ~n34200 & n15526;
  assign n15528 = ~n15033 & n15525;
  assign n15529 = n14813 & ~n34296;
  assign n15530 = n14817 & n15526;
  assign n15531 = n14813 & ~n34200;
  assign n15532 = ~n14805 & n15531;
  assign n15533 = ~n15033 & n15532;
  assign n15534 = ~n14813 & ~n34296;
  assign n15535 = ~n15533 & ~n15534;
  assign n15536 = ~n15529 & ~n15530;
  assign n15537 = ~n15524 & ~n34297;
  assign n15538 = ~n15522 & ~n15537;
  assign n15539 = ~n1388 & ~n15538;
  assign n15540 = ~n14819 & ~n14821;
  assign n15541 = ~n15033 & n15540;
  assign n15542 = ~n34202 & ~n15541;
  assign n15543 = ~n14819 & n34202;
  assign n15544 = ~n14821 & n15543;
  assign n15545 = n34202 & n15541;
  assign n15546 = ~n15033 & n15544;
  assign n15547 = ~n15542 & ~n34298;
  assign n15548 = n1388 & ~n15522;
  assign n15549 = ~n15537 & n15548;
  assign n15550 = n1388 & n15538;
  assign n15551 = ~n15547 & ~n34299;
  assign n15552 = ~n15539 & ~n15551;
  assign n15553 = ~n1192 & ~n15552;
  assign n15554 = n1192 & ~n15539;
  assign n15555 = ~n15551 & n15554;
  assign n15556 = ~n14836 & ~n34204;
  assign n15557 = ~n14836 & ~n15033;
  assign n15558 = ~n34204 & n15557;
  assign n15559 = ~n15033 & n15556;
  assign n15560 = n14844 & ~n34300;
  assign n15561 = n14848 & n15557;
  assign n15562 = n14844 & ~n34204;
  assign n15563 = ~n14836 & n15562;
  assign n15564 = ~n15033 & n15563;
  assign n15565 = ~n14844 & ~n34300;
  assign n15566 = ~n15564 & ~n15565;
  assign n15567 = ~n15560 & ~n15561;
  assign n15568 = ~n15555 & ~n34301;
  assign n15569 = ~n15553 & ~n15568;
  assign n15570 = ~n1028 & ~n15569;
  assign n15571 = n1028 & ~n15553;
  assign n15572 = ~n15568 & n15571;
  assign n15573 = n1028 & n15569;
  assign n15574 = ~n14850 & ~n14860;
  assign n15575 = ~n14850 & ~n15033;
  assign n15576 = ~n14860 & n15575;
  assign n15577 = ~n15033 & n15574;
  assign n15578 = n14858 & ~n34303;
  assign n15579 = n14861 & n15575;
  assign n15580 = ~n14850 & n14858;
  assign n15581 = ~n14860 & n15580;
  assign n15582 = ~n15033 & n15581;
  assign n15583 = ~n14858 & ~n34303;
  assign n15584 = ~n15582 & ~n15583;
  assign n15585 = ~n15578 & ~n15579;
  assign n15586 = ~n34302 & ~n34304;
  assign n15587 = ~n15570 & ~n15586;
  assign n15588 = ~n866 & ~n15587;
  assign n15589 = n866 & ~n15570;
  assign n15590 = ~n15586 & n15589;
  assign n15591 = ~n14863 & ~n34207;
  assign n15592 = ~n14863 & ~n15033;
  assign n15593 = ~n34207 & n15592;
  assign n15594 = ~n15033 & n15591;
  assign n15595 = n14871 & ~n34305;
  assign n15596 = n14875 & n15592;
  assign n15597 = n14871 & ~n34207;
  assign n15598 = ~n14863 & n15597;
  assign n15599 = ~n15033 & n15598;
  assign n15600 = ~n14871 & ~n34305;
  assign n15601 = ~n15599 & ~n15600;
  assign n15602 = ~n15595 & ~n15596;
  assign n15603 = ~n15590 & ~n34306;
  assign n15604 = ~n15588 & ~n15603;
  assign n15605 = ~n730 & ~n15604;
  assign n15606 = ~n14877 & ~n14879;
  assign n15607 = ~n15033 & n15606;
  assign n15608 = ~n34209 & ~n15607;
  assign n15609 = ~n14877 & n34209;
  assign n15610 = ~n14879 & n15609;
  assign n15611 = n34209 & n15607;
  assign n15612 = ~n15033 & n15610;
  assign n15613 = ~n15608 & ~n34307;
  assign n15614 = n730 & ~n15588;
  assign n15615 = ~n15603 & n15614;
  assign n15616 = n730 & n15604;
  assign n15617 = ~n15613 & ~n34308;
  assign n15618 = ~n15605 & ~n15617;
  assign n15619 = ~n602 & ~n15618;
  assign n15620 = n602 & ~n15605;
  assign n15621 = ~n15617 & n15620;
  assign n15622 = ~n14894 & ~n34211;
  assign n15623 = ~n14894 & ~n15033;
  assign n15624 = ~n34211 & n15623;
  assign n15625 = ~n15033 & n15622;
  assign n15626 = n14902 & ~n34309;
  assign n15627 = n14906 & n15623;
  assign n15628 = n14902 & ~n34211;
  assign n15629 = ~n14894 & n15628;
  assign n15630 = ~n15033 & n15629;
  assign n15631 = ~n14902 & ~n34309;
  assign n15632 = ~n15630 & ~n15631;
  assign n15633 = ~n15626 & ~n15627;
  assign n15634 = ~n15621 & ~n34310;
  assign n15635 = ~n15619 & ~n15634;
  assign n15636 = ~n497 & ~n15635;
  assign n15637 = n497 & ~n15619;
  assign n15638 = ~n15634 & n15637;
  assign n15639 = n497 & n15635;
  assign n15640 = ~n14908 & ~n14918;
  assign n15641 = ~n14908 & ~n15033;
  assign n15642 = ~n14918 & n15641;
  assign n15643 = ~n15033 & n15640;
  assign n15644 = n14916 & ~n34312;
  assign n15645 = n14919 & n15641;
  assign n15646 = ~n14908 & n14916;
  assign n15647 = ~n14918 & n15646;
  assign n15648 = ~n15033 & n15647;
  assign n15649 = ~n14916 & ~n34312;
  assign n15650 = ~n15648 & ~n15649;
  assign n15651 = ~n15644 & ~n15645;
  assign n15652 = ~n34311 & ~n34313;
  assign n15653 = ~n15636 & ~n15652;
  assign n15654 = ~n403 & ~n15653;
  assign n15655 = n403 & ~n15636;
  assign n15656 = ~n15652 & n15655;
  assign n15657 = ~n14921 & ~n34214;
  assign n15658 = ~n14921 & ~n15033;
  assign n15659 = ~n34214 & n15658;
  assign n15660 = ~n15033 & n15657;
  assign n15661 = n14929 & ~n34314;
  assign n15662 = n14933 & n15658;
  assign n15663 = n14929 & ~n34214;
  assign n15664 = ~n14921 & n15663;
  assign n15665 = ~n15033 & n15664;
  assign n15666 = ~n14929 & ~n34314;
  assign n15667 = ~n15665 & ~n15666;
  assign n15668 = ~n15661 & ~n15662;
  assign n15669 = ~n15656 & ~n34315;
  assign n15670 = ~n15654 & ~n15669;
  assign n15671 = ~n330 & ~n15670;
  assign n15672 = ~n14935 & ~n14937;
  assign n15673 = ~n15033 & n15672;
  assign n15674 = ~n34216 & ~n15673;
  assign n15675 = ~n14935 & n34216;
  assign n15676 = ~n14937 & n15675;
  assign n15677 = n34216 & n15673;
  assign n15678 = ~n15033 & n15676;
  assign n15679 = ~n15674 & ~n34316;
  assign n15680 = n330 & ~n15654;
  assign n15681 = ~n15669 & n15680;
  assign n15682 = n330 & n15670;
  assign n15683 = ~n15679 & ~n34317;
  assign n15684 = ~n15671 & ~n15683;
  assign n15685 = ~n271 & ~n15684;
  assign n15686 = n271 & ~n15671;
  assign n15687 = ~n15683 & n15686;
  assign n15688 = ~n14952 & ~n34218;
  assign n15689 = ~n14952 & ~n15033;
  assign n15690 = ~n34218 & n15689;
  assign n15691 = ~n15033 & n15688;
  assign n15692 = n14960 & ~n34318;
  assign n15693 = n14964 & n15689;
  assign n15694 = n14960 & ~n34218;
  assign n15695 = ~n14952 & n15694;
  assign n15696 = ~n15033 & n15695;
  assign n15697 = ~n14960 & ~n34318;
  assign n15698 = ~n15696 & ~n15697;
  assign n15699 = ~n15692 & ~n15693;
  assign n15700 = ~n15687 & ~n34319;
  assign n15701 = ~n15685 & ~n15700;
  assign n15702 = ~n217 & ~n15701;
  assign n15703 = n217 & ~n15685;
  assign n15704 = ~n15700 & n15703;
  assign n15705 = n217 & n15701;
  assign n15706 = ~n14966 & ~n14976;
  assign n15707 = ~n14966 & ~n15033;
  assign n15708 = ~n14976 & n15707;
  assign n15709 = ~n15033 & n15706;
  assign n15710 = n14974 & ~n34321;
  assign n15711 = n14977 & n15707;
  assign n15712 = ~n14966 & n14974;
  assign n15713 = ~n14976 & n15712;
  assign n15714 = ~n15033 & n15713;
  assign n15715 = ~n14974 & ~n34321;
  assign n15716 = ~n15714 & ~n15715;
  assign n15717 = ~n15710 & ~n15711;
  assign n15718 = ~n34320 & ~n34322;
  assign n15719 = ~n15702 & ~n15718;
  assign n15720 = ~n198 & ~n15719;
  assign n15721 = n198 & ~n15702;
  assign n15722 = ~n15718 & n15721;
  assign n15723 = ~n14979 & ~n34221;
  assign n15724 = ~n14979 & ~n15033;
  assign n15725 = ~n34221 & n15724;
  assign n15726 = ~n15033 & n15723;
  assign n15727 = n14987 & ~n34323;
  assign n15728 = n14991 & n15724;
  assign n15729 = n14987 & ~n34221;
  assign n15730 = ~n14979 & n15729;
  assign n15731 = ~n15033 & n15730;
  assign n15732 = ~n14987 & ~n34323;
  assign n15733 = ~n15731 & ~n15732;
  assign n15734 = ~n15727 & ~n15728;
  assign n15735 = ~n15722 & ~n34324;
  assign n15736 = ~n15720 & ~n15735;
  assign n15737 = ~n14993 & ~n14995;
  assign n15738 = ~n15033 & n15737;
  assign n15739 = ~n34223 & ~n15738;
  assign n15740 = ~n14993 & n34223;
  assign n15741 = ~n14995 & n15740;
  assign n15742 = n34223 & n15738;
  assign n15743 = ~n15033 & n15741;
  assign n15744 = ~n15739 & ~n34325;
  assign n15745 = ~n15009 & ~n15017;
  assign n15746 = ~n15017 & ~n15033;
  assign n15747 = ~n15009 & n15746;
  assign n15748 = ~n15033 & n15745;
  assign n15749 = ~n34226 & ~n34326;
  assign n15750 = ~n15744 & n15749;
  assign n15751 = ~n15736 & n15750;
  assign n15752 = n193 & ~n15751;
  assign n15753 = ~n15720 & n15744;
  assign n15754 = ~n15735 & n15753;
  assign n15755 = n15736 & n15744;
  assign n15756 = n15009 & ~n15746;
  assign n15757 = ~n193 & ~n15745;
  assign n15758 = ~n15756 & n15757;
  assign n15759 = ~n34327 & ~n15758;
  assign n15760 = ~n15752 & n15759;
  assign n15761 = ~n15437 & ~n15439;
  assign n15762 = ~n15760 & n15761;
  assign n15763 = ~n34228 & ~n15762;
  assign n15764 = n34228 & ~n15439;
  assign n15765 = ~n15437 & n15764;
  assign n15766 = n34228 & n15762;
  assign n15767 = ~n15760 & n15765;
  assign n15768 = ~n15763 & ~n34328;
  assign n15769 = ~n15386 & ~n34277;
  assign n15770 = ~n15760 & n15769;
  assign n15771 = ~n34280 & ~n15770;
  assign n15772 = ~n15386 & n34280;
  assign n15773 = ~n34277 & n15772;
  assign n15774 = n34280 & n15770;
  assign n15775 = ~n15760 & n15773;
  assign n15776 = ~n15771 & ~n34329;
  assign n15777 = ~n15369 & ~n15371;
  assign n15778 = ~n15760 & n15777;
  assign n15779 = ~n34276 & ~n15778;
  assign n15780 = ~n15371 & n34276;
  assign n15781 = ~n15369 & n15780;
  assign n15782 = n34276 & n15778;
  assign n15783 = ~n15760 & n15781;
  assign n15784 = ~n15779 & ~n34330;
  assign n15785 = ~n15335 & ~n15337;
  assign n15786 = ~n15760 & n15785;
  assign n15787 = ~n34271 & ~n15786;
  assign n15788 = ~n15337 & n34271;
  assign n15789 = ~n15335 & n15788;
  assign n15790 = n34271 & n15786;
  assign n15791 = ~n15760 & n15789;
  assign n15792 = ~n15787 & ~n34331;
  assign n15793 = ~n15299 & ~n15301;
  assign n15794 = ~n15760 & n15793;
  assign n15795 = ~n34265 & ~n15794;
  assign n15796 = ~n15301 & n34265;
  assign n15797 = ~n15299 & n15796;
  assign n15798 = n34265 & n15794;
  assign n15799 = ~n15760 & n15797;
  assign n15800 = ~n15795 & ~n34332;
  assign n15801 = ~n15268 & ~n15270;
  assign n15802 = ~n15760 & n15801;
  assign n15803 = ~n34261 & ~n15802;
  assign n15804 = ~n15270 & n34261;
  assign n15805 = ~n15268 & n15804;
  assign n15806 = n34261 & n15802;
  assign n15807 = ~n15760 & n15805;
  assign n15808 = ~n15803 & ~n34333;
  assign n15809 = ~n15232 & ~n15234;
  assign n15810 = ~n15760 & n15809;
  assign n15811 = ~n34255 & ~n15810;
  assign n15812 = ~n15234 & n34255;
  assign n15813 = ~n15232 & n15812;
  assign n15814 = n34255 & n15810;
  assign n15815 = ~n15760 & n15813;
  assign n15816 = ~n15811 & ~n34334;
  assign n15817 = ~n15198 & ~n15200;
  assign n15818 = ~n15760 & n15817;
  assign n15819 = ~n34250 & ~n15818;
  assign n15820 = ~n15200 & n34250;
  assign n15821 = ~n15198 & n15820;
  assign n15822 = n34250 & n15818;
  assign n15823 = ~n15760 & n15821;
  assign n15824 = ~n15819 & ~n34335;
  assign n15825 = ~n15164 & ~n15166;
  assign n15826 = ~n15760 & n15825;
  assign n15827 = ~n34245 & ~n15826;
  assign n15828 = ~n15166 & n34245;
  assign n15829 = ~n15164 & n15828;
  assign n15830 = n34245 & n15826;
  assign n15831 = ~n15760 & n15829;
  assign n15832 = ~n15827 & ~n34336;
  assign n15833 = ~n15131 & ~n15133;
  assign n15834 = ~n15760 & n15833;
  assign n15835 = ~n34241 & ~n15834;
  assign n15836 = ~n15133 & n34241;
  assign n15837 = ~n15131 & n15836;
  assign n15838 = n34241 & n15834;
  assign n15839 = ~n15760 & n15837;
  assign n15840 = ~n15835 & ~n34337;
  assign n15841 = ~n15097 & ~n15099;
  assign n15842 = ~n15760 & n15841;
  assign n15843 = ~n34236 & ~n15842;
  assign n15844 = ~n15099 & n34236;
  assign n15845 = ~n15097 & n15844;
  assign n15846 = n34236 & n15842;
  assign n15847 = ~n15760 & n15845;
  assign n15848 = ~n15843 & ~n34338;
  assign n15849 = ~n15070 & ~n15072;
  assign n15850 = ~n15760 & n15849;
  assign n15851 = ~n15081 & ~n15850;
  assign n15852 = ~n15072 & n15081;
  assign n15853 = ~n15070 & n15852;
  assign n15854 = n15081 & n15850;
  assign n15855 = ~n15760 & n15853;
  assign n15856 = ~n15851 & ~n34339;
  assign n15857 = ~pi38  & ~n15760;
  assign n15858 = ~pi39  & n15857;
  assign n15859 = n15047 & ~n15760;
  assign n15860 = ~n15033 & ~n15758;
  assign n15861 = ~n34327 & n15860;
  assign n15862 = ~n15752 & n15861;
  assign n15863 = ~n34340 & ~n15862;
  assign n15864 = pi40  & ~n15863;
  assign n15865 = ~pi40  & ~n15862;
  assign n15866 = ~pi40  & n15863;
  assign n15867 = ~n34340 & n15865;
  assign n15868 = ~n15864 & ~n34341;
  assign n15869 = pi38  & ~n15760;
  assign n15870 = ~pi36  & ~pi37 ;
  assign n15871 = ~pi38  & n15870;
  assign n15872 = ~n14375 & ~n34230;
  assign n15873 = ~n14376 & n15872;
  assign n15874 = ~n14392 & n15873;
  assign n15875 = ~n34145 & n15874;
  assign n15876 = n34143 & n14394;
  assign n15877 = ~n14386 & n15875;
  assign n15878 = ~n15871 & ~n34342;
  assign n15879 = ~n15031 & n15878;
  assign n15880 = ~n34226 & n15879;
  assign n15881 = ~n15025 & n15880;
  assign n15882 = ~n15869 & ~n15871;
  assign n15883 = n15033 & n15882;
  assign n15884 = ~n15869 & n15881;
  assign n15885 = pi39  & ~n15857;
  assign n15886 = ~n34340 & ~n15885;
  assign n15887 = ~n34343 & n15886;
  assign n15888 = ~n15033 & ~n15882;
  assign n15889 = n14394 & ~n15888;
  assign n15890 = ~n15887 & ~n15888;
  assign n15891 = n14394 & n15890;
  assign n15892 = ~n15887 & n15889;
  assign n15893 = ~n15868 & ~n34344;
  assign n15894 = ~n14394 & ~n15890;
  assign n15895 = n13704 & ~n15894;
  assign n15896 = ~n15893 & n15895;
  assign n15897 = ~n15050 & ~n34231;
  assign n15898 = ~n15760 & n15897;
  assign n15899 = n15055 & ~n15898;
  assign n15900 = ~n15055 & n15897;
  assign n15901 = ~n15055 & n15898;
  assign n15902 = ~n15760 & n15900;
  assign n15903 = ~n15899 & ~n34345;
  assign n15904 = ~n15896 & ~n15903;
  assign n15905 = ~n15893 & ~n15894;
  assign n15906 = ~n13704 & ~n15905;
  assign n15907 = n13099 & ~n15906;
  assign n15908 = ~n15904 & ~n15906;
  assign n15909 = n13099 & n15908;
  assign n15910 = ~n15904 & n15907;
  assign n15911 = ~n15856 & ~n34346;
  assign n15912 = ~n13099 & ~n15908;
  assign n15913 = n12442 & ~n15912;
  assign n15914 = ~n15911 & n15913;
  assign n15915 = ~n15084 & ~n34233;
  assign n15916 = ~n15760 & n15915;
  assign n15917 = n15094 & ~n15916;
  assign n15918 = ~n15094 & n15916;
  assign n15919 = ~n15084 & n15094;
  assign n15920 = ~n34233 & n15919;
  assign n15921 = n15094 & n15916;
  assign n15922 = ~n15760 & n15920;
  assign n15923 = ~n15094 & ~n15916;
  assign n15924 = ~n34347 & ~n15923;
  assign n15925 = ~n15917 & ~n15918;
  assign n15926 = ~n15914 & ~n34348;
  assign n15927 = ~n15911 & ~n15912;
  assign n15928 = ~n12442 & ~n15927;
  assign n15929 = n11858 & ~n15928;
  assign n15930 = ~n15926 & ~n15928;
  assign n15931 = n11858 & n15930;
  assign n15932 = ~n15926 & n15929;
  assign n15933 = ~n15848 & ~n34349;
  assign n15934 = ~n11858 & ~n15930;
  assign n15935 = n11229 & ~n15934;
  assign n15936 = ~n15933 & n15935;
  assign n15937 = ~n15114 & ~n34237;
  assign n15938 = ~n15760 & n15937;
  assign n15939 = ~n34239 & n15938;
  assign n15940 = n34239 & ~n15938;
  assign n15941 = ~n15114 & n34239;
  assign n15942 = ~n34237 & n15941;
  assign n15943 = ~n15760 & n15942;
  assign n15944 = ~n34239 & ~n15938;
  assign n15945 = ~n15943 & ~n15944;
  assign n15946 = ~n15939 & ~n15940;
  assign n15947 = ~n15936 & ~n34350;
  assign n15948 = ~n15933 & ~n15934;
  assign n15949 = ~n11229 & ~n15948;
  assign n15950 = n10681 & ~n15949;
  assign n15951 = ~n15947 & ~n15949;
  assign n15952 = n10681 & n15951;
  assign n15953 = ~n15947 & n15950;
  assign n15954 = ~n15840 & ~n34351;
  assign n15955 = ~n10681 & ~n15951;
  assign n15956 = n10086 & ~n15955;
  assign n15957 = ~n15954 & n15956;
  assign n15958 = ~n15148 & ~n34242;
  assign n15959 = ~n15760 & n15958;
  assign n15960 = ~n34243 & ~n15959;
  assign n15961 = ~n15148 & n34243;
  assign n15962 = ~n34242 & n15961;
  assign n15963 = n34243 & n15959;
  assign n15964 = ~n15760 & n15962;
  assign n15965 = n34243 & ~n15959;
  assign n15966 = ~n34243 & n15959;
  assign n15967 = ~n15965 & ~n15966;
  assign n15968 = ~n15960 & ~n34352;
  assign n15969 = ~n15957 & n34353;
  assign n15970 = ~n15954 & ~n15955;
  assign n15971 = ~n10086 & ~n15970;
  assign n15972 = n9565 & ~n15971;
  assign n15973 = ~n15969 & ~n15971;
  assign n15974 = n9565 & n15973;
  assign n15975 = ~n15969 & n15972;
  assign n15976 = ~n15832 & ~n34354;
  assign n15977 = ~n9565 & ~n15973;
  assign n15978 = n8998 & ~n15977;
  assign n15979 = ~n15976 & n15978;
  assign n15980 = ~n15181 & ~n34246;
  assign n15981 = ~n15760 & n15980;
  assign n15982 = n34248 & ~n15981;
  assign n15983 = ~n15181 & ~n34248;
  assign n15984 = ~n34246 & n15983;
  assign n15985 = ~n34248 & n15981;
  assign n15986 = ~n15760 & n15984;
  assign n15987 = n34248 & n15981;
  assign n15988 = ~n34248 & ~n15981;
  assign n15989 = ~n15987 & ~n15988;
  assign n15990 = ~n15982 & ~n34355;
  assign n15991 = ~n15979 & n34356;
  assign n15992 = ~n15976 & ~n15977;
  assign n15993 = ~n8998 & ~n15992;
  assign n15994 = n8506 & ~n15993;
  assign n15995 = ~n15991 & ~n15993;
  assign n15996 = n8506 & n15995;
  assign n15997 = ~n15991 & n15994;
  assign n15998 = ~n15824 & ~n34357;
  assign n15999 = ~n8506 & ~n15995;
  assign n16000 = n7975 & ~n15999;
  assign n16001 = ~n15998 & n16000;
  assign n16002 = ~n15215 & ~n34251;
  assign n16003 = ~n15215 & ~n15760;
  assign n16004 = ~n34251 & n16003;
  assign n16005 = ~n15760 & n16002;
  assign n16006 = ~n34253 & ~n34358;
  assign n16007 = n15230 & n16003;
  assign n16008 = n34253 & n34358;
  assign n16009 = ~n15215 & ~n34253;
  assign n16010 = ~n34251 & n16009;
  assign n16011 = ~n15760 & n16010;
  assign n16012 = n34253 & ~n34358;
  assign n16013 = ~n16011 & ~n16012;
  assign n16014 = ~n16006 & ~n34359;
  assign n16015 = ~n16001 & ~n34360;
  assign n16016 = ~n15998 & ~n15999;
  assign n16017 = ~n7975 & ~n16016;
  assign n16018 = n7512 & ~n16017;
  assign n16019 = ~n16015 & ~n16017;
  assign n16020 = n7512 & n16019;
  assign n16021 = ~n16015 & n16018;
  assign n16022 = ~n15816 & ~n34361;
  assign n16023 = ~n7512 & ~n16019;
  assign n16024 = n7015 & ~n16023;
  assign n16025 = ~n16022 & n16024;
  assign n16026 = ~n15249 & ~n34256;
  assign n16027 = ~n15760 & n16026;
  assign n16028 = ~n34259 & ~n16027;
  assign n16029 = ~n15249 & n34259;
  assign n16030 = ~n34256 & n16029;
  assign n16031 = n34259 & n16027;
  assign n16032 = ~n15760 & n16030;
  assign n16033 = ~n16028 & ~n34362;
  assign n16034 = ~n16025 & ~n16033;
  assign n16035 = ~n16022 & ~n16023;
  assign n16036 = ~n7015 & ~n16035;
  assign n16037 = n6579 & ~n16036;
  assign n16038 = ~n16034 & ~n16036;
  assign n16039 = n6579 & n16038;
  assign n16040 = ~n16034 & n16037;
  assign n16041 = ~n15808 & ~n34363;
  assign n16042 = ~n6579 & ~n16038;
  assign n16043 = n6117 & ~n16042;
  assign n16044 = ~n16041 & n16043;
  assign n16045 = ~n15285 & ~n34262;
  assign n16046 = ~n15285 & ~n15760;
  assign n16047 = ~n34262 & n16046;
  assign n16048 = ~n15760 & n16045;
  assign n16049 = n15296 & ~n34364;
  assign n16050 = n15297 & n16046;
  assign n16051 = ~n15296 & n34364;
  assign n16052 = ~n15285 & n15296;
  assign n16053 = ~n34262 & n16052;
  assign n16054 = ~n15760 & n16053;
  assign n16055 = ~n15296 & ~n34364;
  assign n16056 = ~n16054 & ~n16055;
  assign n16057 = ~n16049 & ~n34365;
  assign n16058 = ~n16044 & ~n34366;
  assign n16059 = ~n16041 & ~n16042;
  assign n16060 = ~n6117 & ~n16059;
  assign n16061 = n5708 & ~n16060;
  assign n16062 = ~n16058 & ~n16060;
  assign n16063 = n5708 & n16062;
  assign n16064 = ~n16058 & n16061;
  assign n16065 = ~n15800 & ~n34367;
  assign n16066 = ~n5708 & ~n16062;
  assign n16067 = n5278 & ~n16066;
  assign n16068 = ~n16065 & n16067;
  assign n16069 = ~n15316 & ~n34266;
  assign n16070 = ~n15760 & n16069;
  assign n16071 = ~n34269 & n16070;
  assign n16072 = n34269 & ~n16070;
  assign n16073 = ~n15316 & n34269;
  assign n16074 = ~n34266 & n16073;
  assign n16075 = n34269 & n16070;
  assign n16076 = ~n15760 & n16074;
  assign n16077 = ~n34269 & ~n16070;
  assign n16078 = ~n34368 & ~n16077;
  assign n16079 = ~n16071 & ~n16072;
  assign n16080 = ~n16068 & ~n34369;
  assign n16081 = ~n16065 & ~n16066;
  assign n16082 = ~n5278 & ~n16081;
  assign n16083 = n4903 & ~n16082;
  assign n16084 = ~n16080 & ~n16082;
  assign n16085 = n4903 & n16084;
  assign n16086 = ~n16080 & n16083;
  assign n16087 = ~n15792 & ~n34370;
  assign n16088 = ~n4903 & ~n16084;
  assign n16089 = n4508 & ~n16088;
  assign n16090 = ~n16087 & n16089;
  assign n16091 = ~n15352 & ~n34272;
  assign n16092 = ~n15352 & ~n15760;
  assign n16093 = ~n34272 & n16092;
  assign n16094 = ~n15760 & n16091;
  assign n16095 = n34274 & ~n34371;
  assign n16096 = n15367 & n16092;
  assign n16097 = ~n34274 & n34371;
  assign n16098 = ~n15352 & n34274;
  assign n16099 = ~n34272 & n16098;
  assign n16100 = ~n15760 & n16099;
  assign n16101 = ~n34274 & ~n34371;
  assign n16102 = ~n16100 & ~n16101;
  assign n16103 = ~n16095 & ~n34372;
  assign n16104 = ~n16090 & ~n34373;
  assign n16105 = ~n16087 & ~n16088;
  assign n16106 = ~n4508 & ~n16105;
  assign n16107 = n4155 & ~n16106;
  assign n16108 = ~n16104 & ~n16106;
  assign n16109 = n4155 & n16108;
  assign n16110 = ~n16104 & n16107;
  assign n16111 = ~n15784 & ~n34374;
  assign n16112 = ~n4155 & ~n16108;
  assign n16113 = n3788 & ~n16112;
  assign n16114 = ~n16111 & n16113;
  assign n16115 = ~n15776 & ~n16114;
  assign n16116 = ~n16111 & ~n16112;
  assign n16117 = ~n3788 & ~n16116;
  assign n16118 = n3473 & ~n16117;
  assign n16119 = ~n16115 & ~n16117;
  assign n16120 = n3473 & n16119;
  assign n16121 = ~n16115 & n16118;
  assign n16122 = ~n15405 & ~n15407;
  assign n16123 = ~n15760 & n16122;
  assign n16124 = ~n34281 & n16123;
  assign n16125 = n34281 & ~n16123;
  assign n16126 = ~n15407 & n34281;
  assign n16127 = ~n15405 & n16126;
  assign n16128 = ~n15760 & n16127;
  assign n16129 = ~n34281 & ~n16123;
  assign n16130 = ~n16128 & ~n16129;
  assign n16131 = ~n16124 & ~n16125;
  assign n16132 = ~n34375 & ~n34376;
  assign n16133 = ~n3473 & ~n16119;
  assign n16134 = ~n16132 & ~n16133;
  assign n16135 = ~n3140 & ~n16134;
  assign n16136 = n3140 & ~n16133;
  assign n16137 = ~n16132 & n16136;
  assign n16138 = ~n15420 & ~n34284;
  assign n16139 = ~n15760 & n16138;
  assign n16140 = ~n34283 & ~n16139;
  assign n16141 = n34283 & n16139;
  assign n16142 = ~n15420 & ~n34283;
  assign n16143 = ~n34284 & n16142;
  assign n16144 = ~n15760 & n16143;
  assign n16145 = n34283 & ~n16139;
  assign n16146 = ~n16144 & ~n16145;
  assign n16147 = ~n16140 & ~n16141;
  assign n16148 = ~n16137 & ~n34377;
  assign n16149 = ~n16135 & ~n16148;
  assign n16150 = ~n2855 & ~n16149;
  assign n16151 = n2855 & ~n16135;
  assign n16152 = n2855 & n16149;
  assign n16153 = ~n16148 & n16151;
  assign n16154 = ~n15768 & ~n34378;
  assign n16155 = ~n16150 & ~n16154;
  assign n16156 = ~n2556 & ~n16155;
  assign n16157 = n2556 & ~n16150;
  assign n16158 = ~n16154 & n16157;
  assign n16159 = ~n15442 & ~n34286;
  assign n16160 = ~n15442 & ~n15760;
  assign n16161 = ~n34286 & n16160;
  assign n16162 = ~n15760 & n16159;
  assign n16163 = n15450 & ~n34379;
  assign n16164 = n15454 & n16160;
  assign n16165 = ~n15442 & n15450;
  assign n16166 = ~n34286 & n16165;
  assign n16167 = ~n15760 & n16166;
  assign n16168 = ~n15450 & ~n34379;
  assign n16169 = ~n16167 & ~n16168;
  assign n16170 = ~n16163 & ~n16164;
  assign n16171 = ~n16158 & ~n34380;
  assign n16172 = ~n16156 & ~n16171;
  assign n16173 = ~n2301 & ~n16172;
  assign n16174 = ~n15456 & ~n15458;
  assign n16175 = ~n15760 & n16174;
  assign n16176 = ~n34288 & ~n16175;
  assign n16177 = ~n15458 & n34288;
  assign n16178 = ~n15456 & n16177;
  assign n16179 = n34288 & n16175;
  assign n16180 = ~n15760 & n16178;
  assign n16181 = ~n16176 & ~n34381;
  assign n16182 = n2301 & ~n16156;
  assign n16183 = n2301 & n16172;
  assign n16184 = ~n16171 & n16182;
  assign n16185 = ~n16181 & ~n34382;
  assign n16186 = ~n16173 & ~n16185;
  assign n16187 = ~n2038 & ~n16186;
  assign n16188 = n2038 & ~n16173;
  assign n16189 = ~n16185 & n16188;
  assign n16190 = ~n15473 & ~n34290;
  assign n16191 = ~n15473 & ~n15760;
  assign n16192 = ~n34290 & n16191;
  assign n16193 = ~n15760 & n16190;
  assign n16194 = n15481 & ~n34383;
  assign n16195 = n15485 & n16191;
  assign n16196 = ~n15473 & n15481;
  assign n16197 = ~n34290 & n16196;
  assign n16198 = ~n15760 & n16197;
  assign n16199 = ~n15481 & ~n34383;
  assign n16200 = ~n16198 & ~n16199;
  assign n16201 = ~n16194 & ~n16195;
  assign n16202 = ~n16189 & ~n34384;
  assign n16203 = ~n16187 & ~n16202;
  assign n16204 = ~n1812 & ~n16203;
  assign n16205 = ~n15487 & ~n15489;
  assign n16206 = ~n15760 & n16205;
  assign n16207 = ~n34292 & ~n16206;
  assign n16208 = ~n15489 & n34292;
  assign n16209 = ~n15487 & n16208;
  assign n16210 = n34292 & n16206;
  assign n16211 = ~n15760 & n16209;
  assign n16212 = ~n16207 & ~n34385;
  assign n16213 = n1812 & ~n16187;
  assign n16214 = n1812 & n16203;
  assign n16215 = ~n16202 & n16213;
  assign n16216 = ~n16212 & ~n34386;
  assign n16217 = ~n16204 & ~n16216;
  assign n16218 = ~n1582 & ~n16217;
  assign n16219 = ~n15504 & ~n34293;
  assign n16220 = ~n15760 & n16219;
  assign n16221 = ~n34295 & ~n16220;
  assign n16222 = ~n15504 & n34295;
  assign n16223 = ~n34293 & n16222;
  assign n16224 = n34295 & n16220;
  assign n16225 = ~n15760 & n16223;
  assign n16226 = ~n16221 & ~n34387;
  assign n16227 = n1582 & ~n16204;
  assign n16228 = ~n16216 & n16227;
  assign n16229 = ~n16226 & ~n16228;
  assign n16230 = ~n16218 & ~n16229;
  assign n16231 = ~n1388 & ~n16230;
  assign n16232 = ~n15522 & ~n15524;
  assign n16233 = ~n15760 & n16232;
  assign n16234 = ~n34297 & ~n16233;
  assign n16235 = ~n15524 & n34297;
  assign n16236 = ~n15522 & n16235;
  assign n16237 = n34297 & n16233;
  assign n16238 = ~n15760 & n16236;
  assign n16239 = ~n16234 & ~n34388;
  assign n16240 = n1388 & ~n16218;
  assign n16241 = n1388 & n16230;
  assign n16242 = ~n16229 & n16240;
  assign n16243 = ~n16239 & ~n34389;
  assign n16244 = ~n16231 & ~n16243;
  assign n16245 = ~n1192 & ~n16244;
  assign n16246 = n1192 & ~n16231;
  assign n16247 = ~n16243 & n16246;
  assign n16248 = ~n15539 & ~n34299;
  assign n16249 = ~n15539 & ~n15760;
  assign n16250 = ~n34299 & n16249;
  assign n16251 = ~n15760 & n16248;
  assign n16252 = n15547 & ~n34390;
  assign n16253 = n15551 & n16249;
  assign n16254 = ~n15539 & n15547;
  assign n16255 = ~n34299 & n16254;
  assign n16256 = ~n15760 & n16255;
  assign n16257 = ~n15547 & ~n34390;
  assign n16258 = ~n16256 & ~n16257;
  assign n16259 = ~n16252 & ~n16253;
  assign n16260 = ~n16247 & ~n34391;
  assign n16261 = ~n16245 & ~n16260;
  assign n16262 = ~n1028 & ~n16261;
  assign n16263 = ~n15553 & ~n15555;
  assign n16264 = ~n15760 & n16263;
  assign n16265 = ~n34301 & ~n16264;
  assign n16266 = ~n15555 & n34301;
  assign n16267 = ~n15553 & n16266;
  assign n16268 = n34301 & n16264;
  assign n16269 = ~n15760 & n16267;
  assign n16270 = ~n16265 & ~n34392;
  assign n16271 = n1028 & ~n16245;
  assign n16272 = n1028 & n16261;
  assign n16273 = ~n16260 & n16271;
  assign n16274 = ~n16270 & ~n34393;
  assign n16275 = ~n16262 & ~n16274;
  assign n16276 = ~n866 & ~n16275;
  assign n16277 = ~n15570 & ~n34302;
  assign n16278 = ~n15760 & n16277;
  assign n16279 = ~n34304 & ~n16278;
  assign n16280 = ~n15570 & n34304;
  assign n16281 = ~n34302 & n16280;
  assign n16282 = n34304 & n16278;
  assign n16283 = ~n15760 & n16281;
  assign n16284 = ~n16279 & ~n34394;
  assign n16285 = n866 & ~n16262;
  assign n16286 = ~n16274 & n16285;
  assign n16287 = ~n16284 & ~n16286;
  assign n16288 = ~n16276 & ~n16287;
  assign n16289 = ~n730 & ~n16288;
  assign n16290 = ~n15588 & ~n15590;
  assign n16291 = ~n15760 & n16290;
  assign n16292 = ~n34306 & ~n16291;
  assign n16293 = ~n15590 & n34306;
  assign n16294 = ~n15588 & n16293;
  assign n16295 = n34306 & n16291;
  assign n16296 = ~n15760 & n16294;
  assign n16297 = ~n16292 & ~n34395;
  assign n16298 = n730 & ~n16276;
  assign n16299 = n730 & n16288;
  assign n16300 = ~n16287 & n16298;
  assign n16301 = ~n16297 & ~n34396;
  assign n16302 = ~n16289 & ~n16301;
  assign n16303 = ~n602 & ~n16302;
  assign n16304 = n602 & ~n16289;
  assign n16305 = ~n16301 & n16304;
  assign n16306 = ~n15605 & ~n34308;
  assign n16307 = ~n15605 & ~n15760;
  assign n16308 = ~n34308 & n16307;
  assign n16309 = ~n15760 & n16306;
  assign n16310 = n15613 & ~n34397;
  assign n16311 = n15617 & n16307;
  assign n16312 = ~n15605 & n15613;
  assign n16313 = ~n34308 & n16312;
  assign n16314 = ~n15760 & n16313;
  assign n16315 = ~n15613 & ~n34397;
  assign n16316 = ~n16314 & ~n16315;
  assign n16317 = ~n16310 & ~n16311;
  assign n16318 = ~n16305 & ~n34398;
  assign n16319 = ~n16303 & ~n16318;
  assign n16320 = ~n497 & ~n16319;
  assign n16321 = ~n15619 & ~n15621;
  assign n16322 = ~n15760 & n16321;
  assign n16323 = ~n34310 & ~n16322;
  assign n16324 = ~n15621 & n34310;
  assign n16325 = ~n15619 & n16324;
  assign n16326 = n34310 & n16322;
  assign n16327 = ~n15760 & n16325;
  assign n16328 = ~n16323 & ~n34399;
  assign n16329 = n497 & ~n16303;
  assign n16330 = n497 & n16319;
  assign n16331 = ~n16318 & n16329;
  assign n16332 = ~n16328 & ~n34400;
  assign n16333 = ~n16320 & ~n16332;
  assign n16334 = ~n403 & ~n16333;
  assign n16335 = ~n15636 & ~n34311;
  assign n16336 = ~n15760 & n16335;
  assign n16337 = ~n34313 & ~n16336;
  assign n16338 = ~n15636 & n34313;
  assign n16339 = ~n34311 & n16338;
  assign n16340 = n34313 & n16336;
  assign n16341 = ~n15760 & n16339;
  assign n16342 = ~n16337 & ~n34401;
  assign n16343 = n403 & ~n16320;
  assign n16344 = ~n16332 & n16343;
  assign n16345 = ~n16342 & ~n16344;
  assign n16346 = ~n16334 & ~n16345;
  assign n16347 = ~n330 & ~n16346;
  assign n16348 = ~n15654 & ~n15656;
  assign n16349 = ~n15760 & n16348;
  assign n16350 = ~n34315 & ~n16349;
  assign n16351 = ~n15656 & n34315;
  assign n16352 = ~n15654 & n16351;
  assign n16353 = n34315 & n16349;
  assign n16354 = ~n15760 & n16352;
  assign n16355 = ~n16350 & ~n34402;
  assign n16356 = n330 & ~n16334;
  assign n16357 = n330 & n16346;
  assign n16358 = ~n16345 & n16356;
  assign n16359 = ~n16355 & ~n34403;
  assign n16360 = ~n16347 & ~n16359;
  assign n16361 = ~n271 & ~n16360;
  assign n16362 = n271 & ~n16347;
  assign n16363 = ~n16359 & n16362;
  assign n16364 = ~n15671 & ~n34317;
  assign n16365 = ~n15671 & ~n15760;
  assign n16366 = ~n34317 & n16365;
  assign n16367 = ~n15760 & n16364;
  assign n16368 = n15679 & ~n34404;
  assign n16369 = n15683 & n16365;
  assign n16370 = ~n15671 & n15679;
  assign n16371 = ~n34317 & n16370;
  assign n16372 = ~n15760 & n16371;
  assign n16373 = ~n15679 & ~n34404;
  assign n16374 = ~n16372 & ~n16373;
  assign n16375 = ~n16368 & ~n16369;
  assign n16376 = ~n16363 & ~n34405;
  assign n16377 = ~n16361 & ~n16376;
  assign n16378 = ~n217 & ~n16377;
  assign n16379 = ~n15685 & ~n15687;
  assign n16380 = ~n15760 & n16379;
  assign n16381 = ~n34319 & ~n16380;
  assign n16382 = ~n15687 & n34319;
  assign n16383 = ~n15685 & n16382;
  assign n16384 = n34319 & n16380;
  assign n16385 = ~n15760 & n16383;
  assign n16386 = ~n16381 & ~n34406;
  assign n16387 = n217 & ~n16361;
  assign n16388 = n217 & n16377;
  assign n16389 = ~n16376 & n16387;
  assign n16390 = ~n16386 & ~n34407;
  assign n16391 = ~n16378 & ~n16390;
  assign n16392 = ~n198 & ~n16391;
  assign n16393 = ~n15702 & ~n34320;
  assign n16394 = ~n15760 & n16393;
  assign n16395 = ~n34322 & ~n16394;
  assign n16396 = ~n15702 & n34322;
  assign n16397 = ~n34320 & n16396;
  assign n16398 = n34322 & n16394;
  assign n16399 = ~n15760 & n16397;
  assign n16400 = ~n16395 & ~n34408;
  assign n16401 = n198 & ~n16378;
  assign n16402 = ~n16390 & n16401;
  assign n16403 = ~n16400 & ~n16402;
  assign n16404 = ~n16392 & ~n16403;
  assign n16405 = ~n15720 & ~n15722;
  assign n16406 = ~n15760 & n16405;
  assign n16407 = ~n34324 & ~n16406;
  assign n16408 = ~n15722 & n34324;
  assign n16409 = ~n15720 & n16408;
  assign n16410 = n34324 & n16406;
  assign n16411 = ~n15760 & n16409;
  assign n16412 = ~n16407 & ~n34409;
  assign n16413 = ~n15736 & ~n15744;
  assign n16414 = ~n15744 & ~n15760;
  assign n16415 = ~n15736 & n16414;
  assign n16416 = ~n15760 & n16413;
  assign n16417 = ~n34327 & ~n34410;
  assign n16418 = ~n16412 & n16417;
  assign n16419 = ~n16404 & n16418;
  assign n16420 = n193 & ~n16419;
  assign n16421 = ~n16392 & n16412;
  assign n16422 = n16404 & n16412;
  assign n16423 = ~n16403 & n16421;
  assign n16424 = n15736 & ~n16414;
  assign n16425 = ~n193 & ~n16413;
  assign n16426 = ~n16424 & n16425;
  assign n16427 = ~n34411 & ~n16426;
  assign n16428 = ~n16420 & n16427;
  assign n16429 = ~n16150 & ~n34378;
  assign n16430 = ~n16150 & ~n16428;
  assign n16431 = ~n34378 & n16430;
  assign n16432 = ~n16428 & n16429;
  assign n16433 = n15768 & ~n34412;
  assign n16434 = n16154 & n16430;
  assign n16435 = n15768 & ~n34378;
  assign n16436 = ~n16150 & n16435;
  assign n16437 = ~n16428 & n16436;
  assign n16438 = ~n15768 & ~n34412;
  assign n16439 = ~n16437 & ~n16438;
  assign n16440 = ~n16433 & ~n16434;
  assign n16441 = pi36  & ~n16428;
  assign n16442 = ~pi34  & ~pi35 ;
  assign n16443 = ~pi36  & n16442;
  assign n16444 = ~n16441 & ~n16443;
  assign n16445 = ~n15760 & ~n16444;
  assign n16446 = ~pi36  & ~n16428;
  assign n16447 = pi37  & ~n16446;
  assign n16448 = ~pi37  & n16446;
  assign n16449 = n15870 & ~n16428;
  assign n16450 = ~n16447 & ~n34414;
  assign n16451 = ~n34224 & ~n34342;
  assign n16452 = ~n15012 & n16451;
  assign n16453 = ~n15031 & n16452;
  assign n16454 = ~n34226 & n16453;
  assign n16455 = n15017 & n15033;
  assign n16456 = ~n15025 & n16454;
  assign n16457 = ~n16443 & ~n34415;
  assign n16458 = ~n15758 & n16457;
  assign n16459 = ~n34327 & n16458;
  assign n16460 = ~n15752 & n16459;
  assign n16461 = n15760 & n16444;
  assign n16462 = ~n16441 & n16460;
  assign n16463 = n16450 & ~n34416;
  assign n16464 = ~n16445 & ~n16463;
  assign n16465 = ~n15033 & ~n16464;
  assign n16466 = n15033 & ~n16445;
  assign n16467 = ~n16463 & n16466;
  assign n16468 = ~n15760 & ~n16426;
  assign n16469 = ~n34411 & n16468;
  assign n16470 = ~n16420 & n16469;
  assign n16471 = ~n34414 & ~n16470;
  assign n16472 = pi38  & ~n16471;
  assign n16473 = ~pi38  & ~n16470;
  assign n16474 = ~pi38  & n16471;
  assign n16475 = ~n34414 & n16473;
  assign n16476 = ~n16472 & ~n34417;
  assign n16477 = ~n16467 & ~n16476;
  assign n16478 = ~n16465 & ~n16477;
  assign n16479 = ~n14394 & ~n16478;
  assign n16480 = n14394 & ~n16465;
  assign n16481 = ~n16477 & n16480;
  assign n16482 = n14394 & n16478;
  assign n16483 = ~n34343 & ~n15888;
  assign n16484 = ~n16428 & n16483;
  assign n16485 = n15886 & ~n16484;
  assign n16486 = ~n15886 & n16483;
  assign n16487 = ~n15886 & n16484;
  assign n16488 = ~n16428 & n16486;
  assign n16489 = ~n16485 & ~n34419;
  assign n16490 = ~n34418 & ~n16489;
  assign n16491 = ~n16479 & ~n16490;
  assign n16492 = ~n13704 & ~n16491;
  assign n16493 = n13704 & ~n16479;
  assign n16494 = ~n16490 & n16493;
  assign n16495 = ~n34344 & ~n15894;
  assign n16496 = ~n15894 & ~n16428;
  assign n16497 = ~n34344 & n16496;
  assign n16498 = ~n16428 & n16495;
  assign n16499 = n15868 & ~n34420;
  assign n16500 = n15893 & n16496;
  assign n16501 = n15868 & ~n34344;
  assign n16502 = ~n15894 & n16501;
  assign n16503 = ~n16428 & n16502;
  assign n16504 = ~n15868 & ~n34420;
  assign n16505 = ~n16503 & ~n16504;
  assign n16506 = ~n16499 & ~n16500;
  assign n16507 = ~n16494 & ~n34421;
  assign n16508 = ~n16492 & ~n16507;
  assign n16509 = ~n13099 & ~n16508;
  assign n16510 = n13099 & ~n16492;
  assign n16511 = ~n16507 & n16510;
  assign n16512 = n13099 & n16508;
  assign n16513 = ~n15896 & ~n15906;
  assign n16514 = ~n16428 & n16513;
  assign n16515 = n15903 & ~n16514;
  assign n16516 = ~n15903 & n16514;
  assign n16517 = n15903 & ~n15906;
  assign n16518 = ~n15896 & n16517;
  assign n16519 = n15903 & n16514;
  assign n16520 = ~n16428 & n16518;
  assign n16521 = ~n15903 & ~n16514;
  assign n16522 = ~n34423 & ~n16521;
  assign n16523 = ~n16515 & ~n16516;
  assign n16524 = ~n34422 & ~n34424;
  assign n16525 = ~n16509 & ~n16524;
  assign n16526 = ~n12442 & ~n16525;
  assign n16527 = n12442 & ~n16509;
  assign n16528 = ~n16524 & n16527;
  assign n16529 = ~n34346 & ~n15912;
  assign n16530 = ~n15912 & ~n16428;
  assign n16531 = ~n34346 & n16530;
  assign n16532 = ~n16428 & n16529;
  assign n16533 = n15856 & ~n34425;
  assign n16534 = n15911 & n16530;
  assign n16535 = n15856 & ~n34346;
  assign n16536 = ~n15912 & n16535;
  assign n16537 = ~n16428 & n16536;
  assign n16538 = ~n15856 & ~n34425;
  assign n16539 = ~n16537 & ~n16538;
  assign n16540 = ~n16533 & ~n16534;
  assign n16541 = ~n16528 & ~n34426;
  assign n16542 = ~n16526 & ~n16541;
  assign n16543 = ~n11858 & ~n16542;
  assign n16544 = n11858 & ~n16526;
  assign n16545 = ~n16541 & n16544;
  assign n16546 = n11858 & n16542;
  assign n16547 = ~n15914 & ~n15928;
  assign n16548 = ~n16428 & n16547;
  assign n16549 = ~n34348 & n16548;
  assign n16550 = n34348 & ~n16548;
  assign n16551 = n34348 & ~n15928;
  assign n16552 = ~n15914 & n16551;
  assign n16553 = ~n16428 & n16552;
  assign n16554 = ~n34348 & ~n16548;
  assign n16555 = ~n16553 & ~n16554;
  assign n16556 = ~n16549 & ~n16550;
  assign n16557 = ~n34427 & ~n34428;
  assign n16558 = ~n16543 & ~n16557;
  assign n16559 = ~n11229 & ~n16558;
  assign n16560 = n11229 & ~n16543;
  assign n16561 = ~n16557 & n16560;
  assign n16562 = ~n34349 & ~n15934;
  assign n16563 = ~n15934 & ~n16428;
  assign n16564 = ~n34349 & n16563;
  assign n16565 = ~n16428 & n16562;
  assign n16566 = n15848 & ~n34429;
  assign n16567 = n15933 & n16563;
  assign n16568 = n15848 & ~n34349;
  assign n16569 = ~n15934 & n16568;
  assign n16570 = ~n16428 & n16569;
  assign n16571 = ~n15848 & ~n34429;
  assign n16572 = ~n16570 & ~n16571;
  assign n16573 = ~n16566 & ~n16567;
  assign n16574 = ~n16561 & ~n34430;
  assign n16575 = ~n16559 & ~n16574;
  assign n16576 = ~n10681 & ~n16575;
  assign n16577 = n10681 & ~n16559;
  assign n16578 = ~n16574 & n16577;
  assign n16579 = n10681 & n16575;
  assign n16580 = ~n15936 & ~n15949;
  assign n16581 = ~n16428 & n16580;
  assign n16582 = ~n34350 & ~n16581;
  assign n16583 = n34350 & ~n15949;
  assign n16584 = ~n15936 & n16583;
  assign n16585 = n34350 & n16581;
  assign n16586 = ~n16428 & n16584;
  assign n16587 = n34350 & ~n16581;
  assign n16588 = ~n34350 & n16581;
  assign n16589 = ~n16587 & ~n16588;
  assign n16590 = ~n16582 & ~n34432;
  assign n16591 = ~n34431 & n34433;
  assign n16592 = ~n16576 & ~n16591;
  assign n16593 = ~n10086 & ~n16592;
  assign n16594 = n10086 & ~n16576;
  assign n16595 = ~n16591 & n16594;
  assign n16596 = ~n34351 & ~n15955;
  assign n16597 = ~n15955 & ~n16428;
  assign n16598 = ~n34351 & n16597;
  assign n16599 = ~n16428 & n16596;
  assign n16600 = n15840 & ~n34434;
  assign n16601 = n15954 & n16597;
  assign n16602 = n15840 & ~n34351;
  assign n16603 = ~n15955 & n16602;
  assign n16604 = ~n16428 & n16603;
  assign n16605 = ~n15840 & ~n34434;
  assign n16606 = ~n16604 & ~n16605;
  assign n16607 = ~n16600 & ~n16601;
  assign n16608 = ~n16595 & ~n34435;
  assign n16609 = ~n16593 & ~n16608;
  assign n16610 = ~n9565 & ~n16609;
  assign n16611 = n9565 & ~n16593;
  assign n16612 = ~n16608 & n16611;
  assign n16613 = n9565 & n16609;
  assign n16614 = ~n15957 & ~n15971;
  assign n16615 = ~n16428 & n16614;
  assign n16616 = n34353 & ~n16615;
  assign n16617 = ~n34353 & ~n15971;
  assign n16618 = ~n15957 & n16617;
  assign n16619 = ~n34353 & n16615;
  assign n16620 = ~n16428 & n16618;
  assign n16621 = n34353 & n16615;
  assign n16622 = ~n34353 & ~n16615;
  assign n16623 = ~n16621 & ~n16622;
  assign n16624 = ~n16616 & ~n34437;
  assign n16625 = ~n34436 & n34438;
  assign n16626 = ~n16610 & ~n16625;
  assign n16627 = ~n8998 & ~n16626;
  assign n16628 = n8998 & ~n16610;
  assign n16629 = ~n16625 & n16628;
  assign n16630 = ~n34354 & ~n15977;
  assign n16631 = ~n15977 & ~n16428;
  assign n16632 = ~n34354 & n16631;
  assign n16633 = ~n16428 & n16630;
  assign n16634 = n15832 & ~n34439;
  assign n16635 = n15976 & n16631;
  assign n16636 = n15832 & ~n34354;
  assign n16637 = ~n15977 & n16636;
  assign n16638 = ~n16428 & n16637;
  assign n16639 = ~n15832 & ~n34439;
  assign n16640 = ~n16638 & ~n16639;
  assign n16641 = ~n16634 & ~n16635;
  assign n16642 = ~n16629 & ~n34440;
  assign n16643 = ~n16627 & ~n16642;
  assign n16644 = ~n8506 & ~n16643;
  assign n16645 = n8506 & ~n16627;
  assign n16646 = ~n16642 & n16645;
  assign n16647 = n8506 & n16643;
  assign n16648 = ~n15979 & ~n15993;
  assign n16649 = ~n15993 & ~n16428;
  assign n16650 = ~n15979 & n16649;
  assign n16651 = ~n16428 & n16648;
  assign n16652 = ~n34356 & ~n34442;
  assign n16653 = n15991 & n16649;
  assign n16654 = n34356 & n34442;
  assign n16655 = ~n34356 & ~n15993;
  assign n16656 = ~n15979 & n16655;
  assign n16657 = ~n16428 & n16656;
  assign n16658 = n34356 & ~n34442;
  assign n16659 = ~n16657 & ~n16658;
  assign n16660 = ~n16652 & ~n34443;
  assign n16661 = ~n34441 & ~n34444;
  assign n16662 = ~n16644 & ~n16661;
  assign n16663 = ~n7975 & ~n16662;
  assign n16664 = n7975 & ~n16644;
  assign n16665 = ~n16661 & n16664;
  assign n16666 = ~n34357 & ~n15999;
  assign n16667 = ~n15999 & ~n16428;
  assign n16668 = ~n34357 & n16667;
  assign n16669 = ~n16428 & n16666;
  assign n16670 = n15824 & ~n34445;
  assign n16671 = n15998 & n16667;
  assign n16672 = n15824 & ~n34357;
  assign n16673 = ~n15999 & n16672;
  assign n16674 = ~n16428 & n16673;
  assign n16675 = ~n15824 & ~n34445;
  assign n16676 = ~n16674 & ~n16675;
  assign n16677 = ~n16670 & ~n16671;
  assign n16678 = ~n16665 & ~n34446;
  assign n16679 = ~n16663 & ~n16678;
  assign n16680 = ~n7512 & ~n16679;
  assign n16681 = n7512 & ~n16663;
  assign n16682 = ~n16678 & n16681;
  assign n16683 = n7512 & n16679;
  assign n16684 = ~n16001 & ~n16017;
  assign n16685 = ~n16428 & n16684;
  assign n16686 = ~n34360 & ~n16685;
  assign n16687 = n34360 & ~n16017;
  assign n16688 = ~n16001 & n16687;
  assign n16689 = n34360 & n16685;
  assign n16690 = ~n16428 & n16688;
  assign n16691 = ~n16686 & ~n34448;
  assign n16692 = ~n34447 & ~n16691;
  assign n16693 = ~n16680 & ~n16692;
  assign n16694 = ~n7015 & ~n16693;
  assign n16695 = n7015 & ~n16680;
  assign n16696 = ~n16692 & n16695;
  assign n16697 = ~n34361 & ~n16023;
  assign n16698 = ~n16023 & ~n16428;
  assign n16699 = ~n34361 & n16698;
  assign n16700 = ~n16428 & n16697;
  assign n16701 = n15816 & ~n34449;
  assign n16702 = n16022 & n16698;
  assign n16703 = n15816 & ~n34361;
  assign n16704 = ~n16023 & n16703;
  assign n16705 = ~n16428 & n16704;
  assign n16706 = ~n15816 & ~n34449;
  assign n16707 = ~n16705 & ~n16706;
  assign n16708 = ~n16701 & ~n16702;
  assign n16709 = ~n16696 & ~n34450;
  assign n16710 = ~n16694 & ~n16709;
  assign n16711 = ~n6579 & ~n16710;
  assign n16712 = n6579 & ~n16694;
  assign n16713 = ~n16709 & n16712;
  assign n16714 = n6579 & n16710;
  assign n16715 = ~n16025 & ~n16036;
  assign n16716 = ~n16036 & ~n16428;
  assign n16717 = ~n16025 & n16716;
  assign n16718 = ~n16428 & n16715;
  assign n16719 = n16033 & ~n34452;
  assign n16720 = n16034 & n16716;
  assign n16721 = ~n16033 & n34452;
  assign n16722 = n16033 & ~n16036;
  assign n16723 = ~n16025 & n16722;
  assign n16724 = ~n16428 & n16723;
  assign n16725 = ~n16033 & ~n34452;
  assign n16726 = ~n16724 & ~n16725;
  assign n16727 = ~n16719 & ~n34453;
  assign n16728 = ~n34451 & ~n34454;
  assign n16729 = ~n16711 & ~n16728;
  assign n16730 = ~n6117 & ~n16729;
  assign n16731 = n6117 & ~n16711;
  assign n16732 = ~n16728 & n16731;
  assign n16733 = ~n34363 & ~n16042;
  assign n16734 = ~n16042 & ~n16428;
  assign n16735 = ~n34363 & n16734;
  assign n16736 = ~n16428 & n16733;
  assign n16737 = n15808 & ~n34455;
  assign n16738 = n16041 & n16734;
  assign n16739 = n15808 & ~n34363;
  assign n16740 = ~n16042 & n16739;
  assign n16741 = ~n16428 & n16740;
  assign n16742 = ~n15808 & ~n34455;
  assign n16743 = ~n16741 & ~n16742;
  assign n16744 = ~n16737 & ~n16738;
  assign n16745 = ~n16732 & ~n34456;
  assign n16746 = ~n16730 & ~n16745;
  assign n16747 = ~n5708 & ~n16746;
  assign n16748 = n5708 & ~n16730;
  assign n16749 = ~n16745 & n16748;
  assign n16750 = n5708 & n16746;
  assign n16751 = ~n16044 & ~n16060;
  assign n16752 = ~n16428 & n16751;
  assign n16753 = ~n34366 & n16752;
  assign n16754 = n34366 & ~n16752;
  assign n16755 = n34366 & ~n16060;
  assign n16756 = ~n16044 & n16755;
  assign n16757 = n34366 & n16752;
  assign n16758 = ~n16428 & n16756;
  assign n16759 = ~n34366 & ~n16752;
  assign n16760 = ~n34458 & ~n16759;
  assign n16761 = ~n16753 & ~n16754;
  assign n16762 = ~n34457 & ~n34459;
  assign n16763 = ~n16747 & ~n16762;
  assign n16764 = ~n5278 & ~n16763;
  assign n16765 = n5278 & ~n16747;
  assign n16766 = ~n16762 & n16765;
  assign n16767 = ~n34367 & ~n16066;
  assign n16768 = ~n16066 & ~n16428;
  assign n16769 = ~n34367 & n16768;
  assign n16770 = ~n16428 & n16767;
  assign n16771 = n15800 & ~n34460;
  assign n16772 = n16065 & n16768;
  assign n16773 = n15800 & ~n34367;
  assign n16774 = ~n16066 & n16773;
  assign n16775 = ~n16428 & n16774;
  assign n16776 = ~n15800 & ~n34460;
  assign n16777 = ~n16775 & ~n16776;
  assign n16778 = ~n16771 & ~n16772;
  assign n16779 = ~n16766 & ~n34461;
  assign n16780 = ~n16764 & ~n16779;
  assign n16781 = ~n4903 & ~n16780;
  assign n16782 = n4903 & ~n16764;
  assign n16783 = ~n16779 & n16782;
  assign n16784 = n4903 & n16780;
  assign n16785 = ~n16068 & ~n16082;
  assign n16786 = ~n16082 & ~n16428;
  assign n16787 = ~n16068 & n16786;
  assign n16788 = ~n16428 & n16785;
  assign n16789 = n34369 & ~n34463;
  assign n16790 = n16080 & n16786;
  assign n16791 = ~n34369 & n34463;
  assign n16792 = n34369 & ~n16082;
  assign n16793 = ~n16068 & n16792;
  assign n16794 = ~n16428 & n16793;
  assign n16795 = ~n34369 & ~n34463;
  assign n16796 = ~n16794 & ~n16795;
  assign n16797 = ~n16789 & ~n34464;
  assign n16798 = ~n34462 & ~n34465;
  assign n16799 = ~n16781 & ~n16798;
  assign n16800 = ~n4508 & ~n16799;
  assign n16801 = n4508 & ~n16781;
  assign n16802 = ~n16798 & n16801;
  assign n16803 = ~n34370 & ~n16088;
  assign n16804 = ~n16088 & ~n16428;
  assign n16805 = ~n34370 & n16804;
  assign n16806 = ~n16428 & n16803;
  assign n16807 = n15792 & ~n34466;
  assign n16808 = n16087 & n16804;
  assign n16809 = n15792 & ~n34370;
  assign n16810 = ~n16088 & n16809;
  assign n16811 = ~n16428 & n16810;
  assign n16812 = ~n15792 & ~n34466;
  assign n16813 = ~n16811 & ~n16812;
  assign n16814 = ~n16807 & ~n16808;
  assign n16815 = ~n16802 & ~n34467;
  assign n16816 = ~n16800 & ~n16815;
  assign n16817 = ~n4155 & ~n16816;
  assign n16818 = ~n16090 & ~n16106;
  assign n16819 = ~n16428 & n16818;
  assign n16820 = ~n34373 & ~n16819;
  assign n16821 = n34373 & ~n16106;
  assign n16822 = ~n16090 & n16821;
  assign n16823 = n34373 & n16819;
  assign n16824 = ~n16428 & n16822;
  assign n16825 = ~n16820 & ~n34468;
  assign n16826 = n4155 & ~n16800;
  assign n16827 = ~n16815 & n16826;
  assign n16828 = n4155 & n16816;
  assign n16829 = ~n16825 & ~n34469;
  assign n16830 = ~n16817 & ~n16829;
  assign n16831 = ~n3788 & ~n16830;
  assign n16832 = n3788 & ~n16817;
  assign n16833 = ~n16829 & n16832;
  assign n16834 = ~n34374 & ~n16112;
  assign n16835 = ~n16112 & ~n16428;
  assign n16836 = ~n34374 & n16835;
  assign n16837 = ~n16428 & n16834;
  assign n16838 = n15784 & ~n34470;
  assign n16839 = n16111 & n16835;
  assign n16840 = n15784 & ~n34374;
  assign n16841 = ~n16112 & n16840;
  assign n16842 = ~n16428 & n16841;
  assign n16843 = ~n15784 & ~n34470;
  assign n16844 = ~n16842 & ~n16843;
  assign n16845 = ~n16838 & ~n16839;
  assign n16846 = ~n16833 & ~n34471;
  assign n16847 = ~n16831 & ~n16846;
  assign n16848 = ~n3473 & ~n16847;
  assign n16849 = n3473 & ~n16831;
  assign n16850 = ~n16846 & n16849;
  assign n16851 = n3473 & n16847;
  assign n16852 = ~n16114 & ~n16117;
  assign n16853 = ~n16117 & ~n16428;
  assign n16854 = ~n16114 & n16853;
  assign n16855 = ~n16428 & n16852;
  assign n16856 = n15776 & ~n34473;
  assign n16857 = n16115 & n16853;
  assign n16858 = n15776 & ~n16117;
  assign n16859 = ~n16114 & n16858;
  assign n16860 = ~n16428 & n16859;
  assign n16861 = ~n15776 & ~n34473;
  assign n16862 = ~n16860 & ~n16861;
  assign n16863 = ~n16856 & ~n16857;
  assign n16864 = ~n34472 & ~n34474;
  assign n16865 = ~n16848 & ~n16864;
  assign n16866 = ~n3140 & ~n16865;
  assign n16867 = n3140 & ~n16848;
  assign n16868 = ~n16864 & n16867;
  assign n16869 = ~n34375 & ~n16133;
  assign n16870 = ~n16428 & n16869;
  assign n16871 = ~n34376 & n16870;
  assign n16872 = n34376 & ~n16870;
  assign n16873 = ~n34375 & n34376;
  assign n16874 = ~n16133 & n16873;
  assign n16875 = ~n16428 & n16874;
  assign n16876 = ~n34376 & ~n16870;
  assign n16877 = ~n16875 & ~n16876;
  assign n16878 = ~n16871 & ~n16872;
  assign n16879 = ~n16868 & ~n34475;
  assign n16880 = ~n16866 & ~n16879;
  assign n16881 = ~n2855 & ~n16880;
  assign n16882 = n2855 & ~n16866;
  assign n16883 = ~n16879 & n16882;
  assign n16884 = n2855 & n16880;
  assign n16885 = ~n16135 & ~n16137;
  assign n16886 = ~n16428 & n16885;
  assign n16887 = ~n34377 & ~n16886;
  assign n16888 = ~n16135 & n34377;
  assign n16889 = ~n16137 & n16888;
  assign n16890 = n34377 & n16886;
  assign n16891 = ~n16428 & n16889;
  assign n16892 = ~n16887 & ~n34477;
  assign n16893 = ~n34476 & ~n16892;
  assign n16894 = ~n16881 & ~n16893;
  assign n16895 = ~n2556 & ~n16894;
  assign n16896 = n2556 & ~n16881;
  assign n16897 = ~n16893 & n16896;
  assign n16898 = ~n34413 & ~n16897;
  assign n16899 = ~n16895 & ~n16898;
  assign n16900 = ~n2301 & ~n16899;
  assign n16901 = ~n16156 & ~n16158;
  assign n16902 = ~n16428 & n16901;
  assign n16903 = ~n34380 & ~n16902;
  assign n16904 = ~n16156 & n34380;
  assign n16905 = ~n16158 & n16904;
  assign n16906 = n34380 & n16902;
  assign n16907 = ~n16428 & n16905;
  assign n16908 = ~n16903 & ~n34478;
  assign n16909 = n2301 & ~n16895;
  assign n16910 = ~n16898 & n16909;
  assign n16911 = n2301 & n16899;
  assign n16912 = ~n16908 & ~n34479;
  assign n16913 = ~n16900 & ~n16912;
  assign n16914 = ~n2038 & ~n16913;
  assign n16915 = n2038 & ~n16900;
  assign n16916 = ~n16912 & n16915;
  assign n16917 = ~n16173 & ~n34382;
  assign n16918 = ~n16173 & ~n16428;
  assign n16919 = ~n34382 & n16918;
  assign n16920 = ~n16428 & n16917;
  assign n16921 = n16181 & ~n34480;
  assign n16922 = n16185 & n16918;
  assign n16923 = n16181 & ~n34382;
  assign n16924 = ~n16173 & n16923;
  assign n16925 = ~n16428 & n16924;
  assign n16926 = ~n16181 & ~n34480;
  assign n16927 = ~n16925 & ~n16926;
  assign n16928 = ~n16921 & ~n16922;
  assign n16929 = ~n16916 & ~n34481;
  assign n16930 = ~n16914 & ~n16929;
  assign n16931 = ~n1812 & ~n16930;
  assign n16932 = ~n16187 & ~n16189;
  assign n16933 = ~n16428 & n16932;
  assign n16934 = ~n34384 & ~n16933;
  assign n16935 = ~n16187 & n34384;
  assign n16936 = ~n16189 & n16935;
  assign n16937 = n34384 & n16933;
  assign n16938 = ~n16428 & n16936;
  assign n16939 = ~n16934 & ~n34482;
  assign n16940 = n1812 & ~n16914;
  assign n16941 = ~n16929 & n16940;
  assign n16942 = n1812 & n16930;
  assign n16943 = ~n16939 & ~n34483;
  assign n16944 = ~n16931 & ~n16943;
  assign n16945 = ~n1582 & ~n16944;
  assign n16946 = n1582 & ~n16931;
  assign n16947 = ~n16943 & n16946;
  assign n16948 = ~n16204 & ~n34386;
  assign n16949 = ~n16204 & ~n16428;
  assign n16950 = ~n34386 & n16949;
  assign n16951 = ~n16428 & n16948;
  assign n16952 = n16212 & ~n34484;
  assign n16953 = n16216 & n16949;
  assign n16954 = n16212 & ~n34386;
  assign n16955 = ~n16204 & n16954;
  assign n16956 = ~n16428 & n16955;
  assign n16957 = ~n16212 & ~n34484;
  assign n16958 = ~n16956 & ~n16957;
  assign n16959 = ~n16952 & ~n16953;
  assign n16960 = ~n16947 & ~n34485;
  assign n16961 = ~n16945 & ~n16960;
  assign n16962 = ~n1388 & ~n16961;
  assign n16963 = n1388 & ~n16945;
  assign n16964 = ~n16960 & n16963;
  assign n16965 = n1388 & n16961;
  assign n16966 = ~n16218 & ~n16228;
  assign n16967 = ~n16218 & ~n16428;
  assign n16968 = ~n16228 & n16967;
  assign n16969 = ~n16428 & n16966;
  assign n16970 = n16226 & ~n34487;
  assign n16971 = n16229 & n16967;
  assign n16972 = ~n16218 & n16226;
  assign n16973 = ~n16228 & n16972;
  assign n16974 = ~n16428 & n16973;
  assign n16975 = ~n16226 & ~n34487;
  assign n16976 = ~n16974 & ~n16975;
  assign n16977 = ~n16970 & ~n16971;
  assign n16978 = ~n34486 & ~n34488;
  assign n16979 = ~n16962 & ~n16978;
  assign n16980 = ~n1192 & ~n16979;
  assign n16981 = n1192 & ~n16962;
  assign n16982 = ~n16978 & n16981;
  assign n16983 = ~n16231 & ~n34389;
  assign n16984 = ~n16231 & ~n16428;
  assign n16985 = ~n34389 & n16984;
  assign n16986 = ~n16428 & n16983;
  assign n16987 = n16239 & ~n34489;
  assign n16988 = n16243 & n16984;
  assign n16989 = n16239 & ~n34389;
  assign n16990 = ~n16231 & n16989;
  assign n16991 = ~n16428 & n16990;
  assign n16992 = ~n16239 & ~n34489;
  assign n16993 = ~n16991 & ~n16992;
  assign n16994 = ~n16987 & ~n16988;
  assign n16995 = ~n16982 & ~n34490;
  assign n16996 = ~n16980 & ~n16995;
  assign n16997 = ~n1028 & ~n16996;
  assign n16998 = ~n16245 & ~n16247;
  assign n16999 = ~n16428 & n16998;
  assign n17000 = ~n34391 & ~n16999;
  assign n17001 = ~n16245 & n34391;
  assign n17002 = ~n16247 & n17001;
  assign n17003 = n34391 & n16999;
  assign n17004 = ~n16428 & n17002;
  assign n17005 = ~n17000 & ~n34491;
  assign n17006 = n1028 & ~n16980;
  assign n17007 = ~n16995 & n17006;
  assign n17008 = n1028 & n16996;
  assign n17009 = ~n17005 & ~n34492;
  assign n17010 = ~n16997 & ~n17009;
  assign n17011 = ~n866 & ~n17010;
  assign n17012 = n866 & ~n16997;
  assign n17013 = ~n17009 & n17012;
  assign n17014 = ~n16262 & ~n34393;
  assign n17015 = ~n16262 & ~n16428;
  assign n17016 = ~n34393 & n17015;
  assign n17017 = ~n16428 & n17014;
  assign n17018 = n16270 & ~n34493;
  assign n17019 = n16274 & n17015;
  assign n17020 = n16270 & ~n34393;
  assign n17021 = ~n16262 & n17020;
  assign n17022 = ~n16428 & n17021;
  assign n17023 = ~n16270 & ~n34493;
  assign n17024 = ~n17022 & ~n17023;
  assign n17025 = ~n17018 & ~n17019;
  assign n17026 = ~n17013 & ~n34494;
  assign n17027 = ~n17011 & ~n17026;
  assign n17028 = ~n730 & ~n17027;
  assign n17029 = n730 & ~n17011;
  assign n17030 = ~n17026 & n17029;
  assign n17031 = n730 & n17027;
  assign n17032 = ~n16276 & ~n16286;
  assign n17033 = ~n16276 & ~n16428;
  assign n17034 = ~n16286 & n17033;
  assign n17035 = ~n16428 & n17032;
  assign n17036 = n16284 & ~n34496;
  assign n17037 = n16287 & n17033;
  assign n17038 = ~n16276 & n16284;
  assign n17039 = ~n16286 & n17038;
  assign n17040 = ~n16428 & n17039;
  assign n17041 = ~n16284 & ~n34496;
  assign n17042 = ~n17040 & ~n17041;
  assign n17043 = ~n17036 & ~n17037;
  assign n17044 = ~n34495 & ~n34497;
  assign n17045 = ~n17028 & ~n17044;
  assign n17046 = ~n602 & ~n17045;
  assign n17047 = n602 & ~n17028;
  assign n17048 = ~n17044 & n17047;
  assign n17049 = ~n16289 & ~n34396;
  assign n17050 = ~n16289 & ~n16428;
  assign n17051 = ~n34396 & n17050;
  assign n17052 = ~n16428 & n17049;
  assign n17053 = n16297 & ~n34498;
  assign n17054 = n16301 & n17050;
  assign n17055 = n16297 & ~n34396;
  assign n17056 = ~n16289 & n17055;
  assign n17057 = ~n16428 & n17056;
  assign n17058 = ~n16297 & ~n34498;
  assign n17059 = ~n17057 & ~n17058;
  assign n17060 = ~n17053 & ~n17054;
  assign n17061 = ~n17048 & ~n34499;
  assign n17062 = ~n17046 & ~n17061;
  assign n17063 = ~n497 & ~n17062;
  assign n17064 = ~n16303 & ~n16305;
  assign n17065 = ~n16428 & n17064;
  assign n17066 = ~n34398 & ~n17065;
  assign n17067 = ~n16303 & n34398;
  assign n17068 = ~n16305 & n17067;
  assign n17069 = n34398 & n17065;
  assign n17070 = ~n16428 & n17068;
  assign n17071 = ~n17066 & ~n34500;
  assign n17072 = n497 & ~n17046;
  assign n17073 = ~n17061 & n17072;
  assign n17074 = n497 & n17062;
  assign n17075 = ~n17071 & ~n34501;
  assign n17076 = ~n17063 & ~n17075;
  assign n17077 = ~n403 & ~n17076;
  assign n17078 = n403 & ~n17063;
  assign n17079 = ~n17075 & n17078;
  assign n17080 = ~n16320 & ~n34400;
  assign n17081 = ~n16320 & ~n16428;
  assign n17082 = ~n34400 & n17081;
  assign n17083 = ~n16428 & n17080;
  assign n17084 = n16328 & ~n34502;
  assign n17085 = n16332 & n17081;
  assign n17086 = n16328 & ~n34400;
  assign n17087 = ~n16320 & n17086;
  assign n17088 = ~n16428 & n17087;
  assign n17089 = ~n16328 & ~n34502;
  assign n17090 = ~n17088 & ~n17089;
  assign n17091 = ~n17084 & ~n17085;
  assign n17092 = ~n17079 & ~n34503;
  assign n17093 = ~n17077 & ~n17092;
  assign n17094 = ~n330 & ~n17093;
  assign n17095 = n330 & ~n17077;
  assign n17096 = ~n17092 & n17095;
  assign n17097 = n330 & n17093;
  assign n17098 = ~n16334 & ~n16344;
  assign n17099 = ~n16334 & ~n16428;
  assign n17100 = ~n16344 & n17099;
  assign n17101 = ~n16428 & n17098;
  assign n17102 = n16342 & ~n34505;
  assign n17103 = n16345 & n17099;
  assign n17104 = ~n16334 & n16342;
  assign n17105 = ~n16344 & n17104;
  assign n17106 = ~n16428 & n17105;
  assign n17107 = ~n16342 & ~n34505;
  assign n17108 = ~n17106 & ~n17107;
  assign n17109 = ~n17102 & ~n17103;
  assign n17110 = ~n34504 & ~n34506;
  assign n17111 = ~n17094 & ~n17110;
  assign n17112 = ~n271 & ~n17111;
  assign n17113 = n271 & ~n17094;
  assign n17114 = ~n17110 & n17113;
  assign n17115 = ~n16347 & ~n34403;
  assign n17116 = ~n16347 & ~n16428;
  assign n17117 = ~n34403 & n17116;
  assign n17118 = ~n16428 & n17115;
  assign n17119 = n16355 & ~n34507;
  assign n17120 = n16359 & n17116;
  assign n17121 = n16355 & ~n34403;
  assign n17122 = ~n16347 & n17121;
  assign n17123 = ~n16428 & n17122;
  assign n17124 = ~n16355 & ~n34507;
  assign n17125 = ~n17123 & ~n17124;
  assign n17126 = ~n17119 & ~n17120;
  assign n17127 = ~n17114 & ~n34508;
  assign n17128 = ~n17112 & ~n17127;
  assign n17129 = ~n217 & ~n17128;
  assign n17130 = ~n16361 & ~n16363;
  assign n17131 = ~n16428 & n17130;
  assign n17132 = ~n34405 & ~n17131;
  assign n17133 = ~n16361 & n34405;
  assign n17134 = ~n16363 & n17133;
  assign n17135 = n34405 & n17131;
  assign n17136 = ~n16428 & n17134;
  assign n17137 = ~n17132 & ~n34509;
  assign n17138 = n217 & ~n17112;
  assign n17139 = ~n17127 & n17138;
  assign n17140 = n217 & n17128;
  assign n17141 = ~n17137 & ~n34510;
  assign n17142 = ~n17129 & ~n17141;
  assign n17143 = ~n198 & ~n17142;
  assign n17144 = n198 & ~n17129;
  assign n17145 = ~n17141 & n17144;
  assign n17146 = ~n16378 & ~n34407;
  assign n17147 = ~n16378 & ~n16428;
  assign n17148 = ~n34407 & n17147;
  assign n17149 = ~n16428 & n17146;
  assign n17150 = n16386 & ~n34511;
  assign n17151 = n16390 & n17147;
  assign n17152 = n16386 & ~n34407;
  assign n17153 = ~n16378 & n17152;
  assign n17154 = ~n16428 & n17153;
  assign n17155 = ~n16386 & ~n34511;
  assign n17156 = ~n17154 & ~n17155;
  assign n17157 = ~n17150 & ~n17151;
  assign n17158 = ~n17145 & ~n34512;
  assign n17159 = ~n17143 & ~n17158;
  assign n17160 = ~n16392 & ~n16402;
  assign n17161 = ~n16392 & ~n16428;
  assign n17162 = ~n16402 & n17161;
  assign n17163 = ~n16428 & n17160;
  assign n17164 = n16400 & ~n34513;
  assign n17165 = n16403 & n17161;
  assign n17166 = ~n16392 & n16400;
  assign n17167 = ~n16402 & n17166;
  assign n17168 = ~n16428 & n17167;
  assign n17169 = ~n16400 & ~n34513;
  assign n17170 = ~n17168 & ~n17169;
  assign n17171 = ~n17164 & ~n17165;
  assign n17172 = ~n16404 & ~n16412;
  assign n17173 = ~n16412 & ~n16428;
  assign n17174 = ~n16404 & n17173;
  assign n17175 = ~n16428 & n17172;
  assign n17176 = ~n34411 & ~n34515;
  assign n17177 = ~n34514 & n17176;
  assign n17178 = ~n17159 & n17177;
  assign n17179 = n193 & ~n17178;
  assign n17180 = ~n17143 & n34514;
  assign n17181 = ~n17158 & n17180;
  assign n17182 = n17159 & n34514;
  assign n17183 = n16404 & ~n17173;
  assign n17184 = ~n193 & ~n17172;
  assign n17185 = ~n17183 & n17184;
  assign n17186 = ~n34516 & ~n17185;
  assign n17187 = ~n17179 & n17186;
  assign n17188 = ~n16895 & ~n16897;
  assign n17189 = ~n17187 & n17188;
  assign n17190 = ~n34413 & ~n17189;
  assign n17191 = n34413 & ~n16897;
  assign n17192 = ~n16895 & n17191;
  assign n17193 = n34413 & n17189;
  assign n17194 = ~n17187 & n17192;
  assign n17195 = ~n17190 & ~n34517;
  assign n17196 = ~n16866 & ~n16868;
  assign n17197 = ~n17187 & n17196;
  assign n17198 = ~n34475 & ~n17197;
  assign n17199 = ~n16868 & n34475;
  assign n17200 = ~n16866 & n17199;
  assign n17201 = n34475 & n17197;
  assign n17202 = ~n17187 & n17200;
  assign n17203 = ~n17198 & ~n34518;
  assign n17204 = ~n16848 & ~n34472;
  assign n17205 = ~n17187 & n17204;
  assign n17206 = ~n34474 & ~n17205;
  assign n17207 = ~n16848 & n34474;
  assign n17208 = ~n34472 & n17207;
  assign n17209 = n34474 & n17205;
  assign n17210 = ~n17187 & n17208;
  assign n17211 = ~n17206 & ~n34519;
  assign n17212 = ~n16831 & ~n16833;
  assign n17213 = ~n17187 & n17212;
  assign n17214 = ~n34471 & ~n17213;
  assign n17215 = ~n16833 & n34471;
  assign n17216 = ~n16831 & n17215;
  assign n17217 = n34471 & n17213;
  assign n17218 = ~n17187 & n17216;
  assign n17219 = ~n17214 & ~n34520;
  assign n17220 = ~n16800 & ~n16802;
  assign n17221 = ~n17187 & n17220;
  assign n17222 = ~n34467 & ~n17221;
  assign n17223 = ~n16802 & n34467;
  assign n17224 = ~n16800 & n17223;
  assign n17225 = n34467 & n17221;
  assign n17226 = ~n17187 & n17224;
  assign n17227 = ~n17222 & ~n34521;
  assign n17228 = ~n16781 & ~n34462;
  assign n17229 = ~n17187 & n17228;
  assign n17230 = ~n34465 & ~n17229;
  assign n17231 = ~n16781 & n34465;
  assign n17232 = ~n34462 & n17231;
  assign n17233 = n34465 & n17229;
  assign n17234 = ~n17187 & n17232;
  assign n17235 = ~n17230 & ~n34522;
  assign n17236 = ~n16764 & ~n16766;
  assign n17237 = ~n17187 & n17236;
  assign n17238 = ~n34461 & ~n17237;
  assign n17239 = ~n16766 & n34461;
  assign n17240 = ~n16764 & n17239;
  assign n17241 = n34461 & n17237;
  assign n17242 = ~n17187 & n17240;
  assign n17243 = ~n17238 & ~n34523;
  assign n17244 = ~n16730 & ~n16732;
  assign n17245 = ~n17187 & n17244;
  assign n17246 = ~n34456 & ~n17245;
  assign n17247 = ~n16732 & n34456;
  assign n17248 = ~n16730 & n17247;
  assign n17249 = n34456 & n17245;
  assign n17250 = ~n17187 & n17248;
  assign n17251 = ~n17246 & ~n34524;
  assign n17252 = ~n16694 & ~n16696;
  assign n17253 = ~n17187 & n17252;
  assign n17254 = ~n34450 & ~n17253;
  assign n17255 = ~n16696 & n34450;
  assign n17256 = ~n16694 & n17255;
  assign n17257 = n34450 & n17253;
  assign n17258 = ~n17187 & n17256;
  assign n17259 = ~n17254 & ~n34525;
  assign n17260 = ~n16663 & ~n16665;
  assign n17261 = ~n17187 & n17260;
  assign n17262 = ~n34446 & ~n17261;
  assign n17263 = ~n16665 & n34446;
  assign n17264 = ~n16663 & n17263;
  assign n17265 = n34446 & n17261;
  assign n17266 = ~n17187 & n17264;
  assign n17267 = ~n17262 & ~n34526;
  assign n17268 = ~n16627 & ~n16629;
  assign n17269 = ~n17187 & n17268;
  assign n17270 = ~n34440 & ~n17269;
  assign n17271 = ~n16629 & n34440;
  assign n17272 = ~n16627 & n17271;
  assign n17273 = n34440 & n17269;
  assign n17274 = ~n17187 & n17272;
  assign n17275 = ~n17270 & ~n34527;
  assign n17276 = ~n16593 & ~n16595;
  assign n17277 = ~n17187 & n17276;
  assign n17278 = ~n34435 & ~n17277;
  assign n17279 = ~n16595 & n34435;
  assign n17280 = ~n16593 & n17279;
  assign n17281 = n34435 & n17277;
  assign n17282 = ~n17187 & n17280;
  assign n17283 = ~n17278 & ~n34528;
  assign n17284 = ~n16559 & ~n16561;
  assign n17285 = ~n17187 & n17284;
  assign n17286 = ~n34430 & ~n17285;
  assign n17287 = ~n16561 & n34430;
  assign n17288 = ~n16559 & n17287;
  assign n17289 = n34430 & n17285;
  assign n17290 = ~n17187 & n17288;
  assign n17291 = ~n17286 & ~n34529;
  assign n17292 = ~n16526 & ~n16528;
  assign n17293 = ~n17187 & n17292;
  assign n17294 = ~n34426 & ~n17293;
  assign n17295 = ~n16528 & n34426;
  assign n17296 = ~n16526 & n17295;
  assign n17297 = n34426 & n17293;
  assign n17298 = ~n17187 & n17296;
  assign n17299 = ~n17294 & ~n34530;
  assign n17300 = ~n16492 & ~n16494;
  assign n17301 = ~n17187 & n17300;
  assign n17302 = ~n34421 & ~n17301;
  assign n17303 = ~n16494 & n34421;
  assign n17304 = ~n16492 & n17303;
  assign n17305 = n34421 & n17301;
  assign n17306 = ~n17187 & n17304;
  assign n17307 = ~n17302 & ~n34531;
  assign n17308 = ~n16465 & ~n16467;
  assign n17309 = ~n17187 & n17308;
  assign n17310 = ~n16476 & ~n17309;
  assign n17311 = ~n16467 & n16476;
  assign n17312 = ~n16465 & n17311;
  assign n17313 = n16476 & n17309;
  assign n17314 = ~n17187 & n17312;
  assign n17315 = ~n17310 & ~n34532;
  assign n17316 = ~pi34  & ~n17187;
  assign n17317 = ~pi35  & n17316;
  assign n17318 = n16442 & ~n17187;
  assign n17319 = ~n16428 & ~n17185;
  assign n17320 = ~n34516 & n17319;
  assign n17321 = ~n17179 & n17320;
  assign n17322 = ~n34533 & ~n17321;
  assign n17323 = pi36  & ~n17322;
  assign n17324 = ~pi36  & ~n17321;
  assign n17325 = ~pi36  & n17322;
  assign n17326 = ~n34533 & n17324;
  assign n17327 = ~n17323 & ~n34534;
  assign n17328 = pi34  & ~n17187;
  assign n17329 = ~pi32  & ~pi33 ;
  assign n17330 = ~pi34  & n17329;
  assign n17331 = ~n34325 & ~n34415;
  assign n17332 = ~n15739 & n17331;
  assign n17333 = ~n15758 & n17332;
  assign n17334 = ~n34327 & n17333;
  assign n17335 = n15744 & n15760;
  assign n17336 = ~n15752 & n17334;
  assign n17337 = ~n17330 & ~n34535;
  assign n17338 = ~n16426 & n17337;
  assign n17339 = ~n34411 & n17338;
  assign n17340 = ~n16420 & n17339;
  assign n17341 = ~n17328 & ~n17330;
  assign n17342 = n16428 & n17341;
  assign n17343 = ~n17328 & n17340;
  assign n17344 = pi35  & ~n17316;
  assign n17345 = ~n34533 & ~n17344;
  assign n17346 = ~n34536 & n17345;
  assign n17347 = ~n16428 & ~n17341;
  assign n17348 = n15760 & ~n17347;
  assign n17349 = ~n17346 & ~n17347;
  assign n17350 = n15760 & n17349;
  assign n17351 = ~n17346 & n17348;
  assign n17352 = ~n17327 & ~n34537;
  assign n17353 = ~n15760 & ~n17349;
  assign n17354 = n15033 & ~n17353;
  assign n17355 = ~n17352 & n17354;
  assign n17356 = ~n16445 & ~n34416;
  assign n17357 = ~n17187 & n17356;
  assign n17358 = n16450 & ~n17357;
  assign n17359 = ~n16450 & n17356;
  assign n17360 = ~n16450 & n17357;
  assign n17361 = ~n17187 & n17359;
  assign n17362 = ~n17358 & ~n34538;
  assign n17363 = ~n17355 & ~n17362;
  assign n17364 = ~n17352 & ~n17353;
  assign n17365 = ~n15033 & ~n17364;
  assign n17366 = n14394 & ~n17365;
  assign n17367 = ~n17363 & ~n17365;
  assign n17368 = n14394 & n17367;
  assign n17369 = ~n17363 & n17366;
  assign n17370 = ~n17315 & ~n34539;
  assign n17371 = ~n14394 & ~n17367;
  assign n17372 = n13704 & ~n17371;
  assign n17373 = ~n17370 & n17372;
  assign n17374 = ~n16479 & ~n34418;
  assign n17375 = ~n17187 & n17374;
  assign n17376 = n16489 & ~n17375;
  assign n17377 = ~n16489 & n17375;
  assign n17378 = ~n16479 & n16489;
  assign n17379 = ~n34418 & n17378;
  assign n17380 = n16489 & n17375;
  assign n17381 = ~n17187 & n17379;
  assign n17382 = ~n16489 & ~n17375;
  assign n17383 = ~n34540 & ~n17382;
  assign n17384 = ~n17376 & ~n17377;
  assign n17385 = ~n17373 & ~n34541;
  assign n17386 = ~n17370 & ~n17371;
  assign n17387 = ~n13704 & ~n17386;
  assign n17388 = n13099 & ~n17387;
  assign n17389 = ~n17385 & ~n17387;
  assign n17390 = n13099 & n17389;
  assign n17391 = ~n17385 & n17388;
  assign n17392 = ~n17307 & ~n34542;
  assign n17393 = ~n13099 & ~n17389;
  assign n17394 = n12442 & ~n17393;
  assign n17395 = ~n17392 & n17394;
  assign n17396 = ~n16509 & ~n34422;
  assign n17397 = ~n17187 & n17396;
  assign n17398 = ~n34424 & n17397;
  assign n17399 = n34424 & ~n17397;
  assign n17400 = ~n16509 & n34424;
  assign n17401 = ~n34422 & n17400;
  assign n17402 = ~n17187 & n17401;
  assign n17403 = ~n34424 & ~n17397;
  assign n17404 = ~n17402 & ~n17403;
  assign n17405 = ~n17398 & ~n17399;
  assign n17406 = ~n17395 & ~n34543;
  assign n17407 = ~n17392 & ~n17393;
  assign n17408 = ~n12442 & ~n17407;
  assign n17409 = n11858 & ~n17408;
  assign n17410 = ~n17406 & ~n17408;
  assign n17411 = n11858 & n17410;
  assign n17412 = ~n17406 & n17409;
  assign n17413 = ~n17299 & ~n34544;
  assign n17414 = ~n11858 & ~n17410;
  assign n17415 = n11229 & ~n17414;
  assign n17416 = ~n17413 & n17415;
  assign n17417 = ~n16543 & ~n34427;
  assign n17418 = ~n17187 & n17417;
  assign n17419 = ~n34428 & ~n17418;
  assign n17420 = ~n16543 & n34428;
  assign n17421 = ~n34427 & n17420;
  assign n17422 = n34428 & n17418;
  assign n17423 = ~n17187 & n17421;
  assign n17424 = n34428 & ~n17418;
  assign n17425 = ~n34428 & n17418;
  assign n17426 = ~n17424 & ~n17425;
  assign n17427 = ~n17419 & ~n34545;
  assign n17428 = ~n17416 & n34546;
  assign n17429 = ~n17413 & ~n17414;
  assign n17430 = ~n11229 & ~n17429;
  assign n17431 = n10681 & ~n17430;
  assign n17432 = ~n17428 & ~n17430;
  assign n17433 = n10681 & n17432;
  assign n17434 = ~n17428 & n17431;
  assign n17435 = ~n17291 & ~n34547;
  assign n17436 = ~n10681 & ~n17432;
  assign n17437 = n10086 & ~n17436;
  assign n17438 = ~n17435 & n17437;
  assign n17439 = ~n16576 & ~n34431;
  assign n17440 = ~n17187 & n17439;
  assign n17441 = n34433 & ~n17440;
  assign n17442 = ~n16576 & ~n34433;
  assign n17443 = ~n34431 & n17442;
  assign n17444 = ~n34433 & n17440;
  assign n17445 = ~n17187 & n17443;
  assign n17446 = n34433 & n17440;
  assign n17447 = ~n34433 & ~n17440;
  assign n17448 = ~n17446 & ~n17447;
  assign n17449 = ~n17441 & ~n34548;
  assign n17450 = ~n17438 & n34549;
  assign n17451 = ~n17435 & ~n17436;
  assign n17452 = ~n10086 & ~n17451;
  assign n17453 = n9565 & ~n17452;
  assign n17454 = ~n17450 & ~n17452;
  assign n17455 = n9565 & n17454;
  assign n17456 = ~n17450 & n17453;
  assign n17457 = ~n17283 & ~n34550;
  assign n17458 = ~n9565 & ~n17454;
  assign n17459 = n8998 & ~n17458;
  assign n17460 = ~n17457 & n17459;
  assign n17461 = ~n16610 & ~n34436;
  assign n17462 = ~n16610 & ~n17187;
  assign n17463 = ~n34436 & n17462;
  assign n17464 = ~n17187 & n17461;
  assign n17465 = ~n34438 & ~n34551;
  assign n17466 = n16625 & n17462;
  assign n17467 = n34438 & n34551;
  assign n17468 = ~n16610 & ~n34438;
  assign n17469 = ~n34436 & n17468;
  assign n17470 = ~n17187 & n17469;
  assign n17471 = n34438 & ~n34551;
  assign n17472 = ~n17470 & ~n17471;
  assign n17473 = ~n17465 & ~n34552;
  assign n17474 = ~n17460 & ~n34553;
  assign n17475 = ~n17457 & ~n17458;
  assign n17476 = ~n8998 & ~n17475;
  assign n17477 = n8506 & ~n17476;
  assign n17478 = ~n17474 & ~n17476;
  assign n17479 = n8506 & n17478;
  assign n17480 = ~n17474 & n17477;
  assign n17481 = ~n17275 & ~n34554;
  assign n17482 = ~n8506 & ~n17478;
  assign n17483 = n7975 & ~n17482;
  assign n17484 = ~n17481 & n17483;
  assign n17485 = ~n16644 & ~n34441;
  assign n17486 = ~n17187 & n17485;
  assign n17487 = ~n34444 & ~n17486;
  assign n17488 = ~n16644 & n34444;
  assign n17489 = ~n34441 & n17488;
  assign n17490 = n34444 & n17486;
  assign n17491 = ~n17187 & n17489;
  assign n17492 = ~n17487 & ~n34555;
  assign n17493 = ~n17484 & ~n17492;
  assign n17494 = ~n17481 & ~n17482;
  assign n17495 = ~n7975 & ~n17494;
  assign n17496 = n7512 & ~n17495;
  assign n17497 = ~n17493 & ~n17495;
  assign n17498 = n7512 & n17497;
  assign n17499 = ~n17493 & n17496;
  assign n17500 = ~n17267 & ~n34556;
  assign n17501 = ~n7512 & ~n17497;
  assign n17502 = n7015 & ~n17501;
  assign n17503 = ~n17500 & n17502;
  assign n17504 = ~n16680 & ~n34447;
  assign n17505 = ~n16680 & ~n17187;
  assign n17506 = ~n34447 & n17505;
  assign n17507 = ~n17187 & n17504;
  assign n17508 = n16691 & ~n34557;
  assign n17509 = n16692 & n17505;
  assign n17510 = ~n16691 & n34557;
  assign n17511 = ~n16680 & n16691;
  assign n17512 = ~n34447 & n17511;
  assign n17513 = ~n17187 & n17512;
  assign n17514 = ~n16691 & ~n34557;
  assign n17515 = ~n17513 & ~n17514;
  assign n17516 = ~n17508 & ~n34558;
  assign n17517 = ~n17503 & ~n34559;
  assign n17518 = ~n17500 & ~n17501;
  assign n17519 = ~n7015 & ~n17518;
  assign n17520 = n6579 & ~n17519;
  assign n17521 = ~n17517 & ~n17519;
  assign n17522 = n6579 & n17521;
  assign n17523 = ~n17517 & n17520;
  assign n17524 = ~n17259 & ~n34560;
  assign n17525 = ~n6579 & ~n17521;
  assign n17526 = n6117 & ~n17525;
  assign n17527 = ~n17524 & n17526;
  assign n17528 = ~n16711 & ~n34451;
  assign n17529 = ~n17187 & n17528;
  assign n17530 = ~n34454 & n17529;
  assign n17531 = n34454 & ~n17529;
  assign n17532 = ~n16711 & n34454;
  assign n17533 = ~n34451 & n17532;
  assign n17534 = n34454 & n17529;
  assign n17535 = ~n17187 & n17533;
  assign n17536 = ~n34454 & ~n17529;
  assign n17537 = ~n34561 & ~n17536;
  assign n17538 = ~n17530 & ~n17531;
  assign n17539 = ~n17527 & ~n34562;
  assign n17540 = ~n17524 & ~n17525;
  assign n17541 = ~n6117 & ~n17540;
  assign n17542 = n5708 & ~n17541;
  assign n17543 = ~n17539 & ~n17541;
  assign n17544 = n5708 & n17543;
  assign n17545 = ~n17539 & n17542;
  assign n17546 = ~n17251 & ~n34563;
  assign n17547 = ~n5708 & ~n17543;
  assign n17548 = n5278 & ~n17547;
  assign n17549 = ~n17546 & n17548;
  assign n17550 = ~n16747 & ~n34457;
  assign n17551 = ~n16747 & ~n17187;
  assign n17552 = ~n34457 & n17551;
  assign n17553 = ~n17187 & n17550;
  assign n17554 = n34459 & ~n34564;
  assign n17555 = n16762 & n17551;
  assign n17556 = ~n34459 & n34564;
  assign n17557 = ~n16747 & n34459;
  assign n17558 = ~n34457 & n17557;
  assign n17559 = ~n17187 & n17558;
  assign n17560 = ~n34459 & ~n34564;
  assign n17561 = ~n17559 & ~n17560;
  assign n17562 = ~n17554 & ~n34565;
  assign n17563 = ~n17549 & ~n34566;
  assign n17564 = ~n17546 & ~n17547;
  assign n17565 = ~n5278 & ~n17564;
  assign n17566 = n4903 & ~n17565;
  assign n17567 = ~n17563 & ~n17565;
  assign n17568 = n4903 & n17567;
  assign n17569 = ~n17563 & n17566;
  assign n17570 = ~n17243 & ~n34567;
  assign n17571 = ~n4903 & ~n17567;
  assign n17572 = n4508 & ~n17571;
  assign n17573 = ~n17570 & n17572;
  assign n17574 = ~n17235 & ~n17573;
  assign n17575 = ~n17570 & ~n17571;
  assign n17576 = ~n4508 & ~n17575;
  assign n17577 = n4155 & ~n17576;
  assign n17578 = ~n17574 & ~n17576;
  assign n17579 = n4155 & n17578;
  assign n17580 = ~n17574 & n17577;
  assign n17581 = ~n17227 & ~n34568;
  assign n17582 = ~n4155 & ~n17578;
  assign n17583 = n3788 & ~n17582;
  assign n17584 = ~n17581 & n17583;
  assign n17585 = ~n16817 & ~n34469;
  assign n17586 = ~n16817 & ~n17187;
  assign n17587 = ~n34469 & n17586;
  assign n17588 = ~n17187 & n17585;
  assign n17589 = n16825 & ~n34569;
  assign n17590 = n16829 & n17586;
  assign n17591 = ~n16817 & n16825;
  assign n17592 = ~n34469 & n17591;
  assign n17593 = ~n17187 & n17592;
  assign n17594 = ~n16825 & ~n34569;
  assign n17595 = ~n17593 & ~n17594;
  assign n17596 = ~n17589 & ~n17590;
  assign n17597 = ~n17584 & ~n34570;
  assign n17598 = ~n17581 & ~n17582;
  assign n17599 = ~n3788 & ~n17598;
  assign n17600 = n3473 & ~n17599;
  assign n17601 = ~n17597 & ~n17599;
  assign n17602 = n3473 & n17601;
  assign n17603 = ~n17597 & n17600;
  assign n17604 = ~n17219 & ~n34571;
  assign n17605 = ~n3473 & ~n17601;
  assign n17606 = n3140 & ~n17605;
  assign n17607 = ~n17604 & n17606;
  assign n17608 = ~n17211 & ~n17607;
  assign n17609 = ~n17604 & ~n17605;
  assign n17610 = ~n3140 & ~n17609;
  assign n17611 = n2855 & ~n17610;
  assign n17612 = ~n17608 & ~n17610;
  assign n17613 = n2855 & n17612;
  assign n17614 = ~n17608 & n17611;
  assign n17615 = ~n17203 & ~n34572;
  assign n17616 = ~n2855 & ~n17612;
  assign n17617 = ~n17615 & ~n17616;
  assign n17618 = ~n2556 & ~n17617;
  assign n17619 = n2556 & ~n17616;
  assign n17620 = ~n17615 & n17619;
  assign n17621 = ~n16881 & ~n34476;
  assign n17622 = ~n17187 & n17621;
  assign n17623 = n16892 & ~n17622;
  assign n17624 = ~n16892 & n17622;
  assign n17625 = ~n16881 & n16892;
  assign n17626 = ~n34476 & n17625;
  assign n17627 = n16892 & n17622;
  assign n17628 = ~n17187 & n17626;
  assign n17629 = ~n16892 & ~n17622;
  assign n17630 = ~n34573 & ~n17629;
  assign n17631 = ~n17623 & ~n17624;
  assign n17632 = ~n17620 & ~n34574;
  assign n17633 = ~n17618 & ~n17632;
  assign n17634 = ~n2301 & ~n17633;
  assign n17635 = n2301 & ~n17618;
  assign n17636 = n2301 & n17633;
  assign n17637 = ~n17632 & n17635;
  assign n17638 = ~n17195 & ~n34575;
  assign n17639 = ~n17634 & ~n17638;
  assign n17640 = ~n2038 & ~n17639;
  assign n17641 = n2038 & ~n17634;
  assign n17642 = ~n17638 & n17641;
  assign n17643 = ~n16900 & ~n34479;
  assign n17644 = ~n16900 & ~n17187;
  assign n17645 = ~n34479 & n17644;
  assign n17646 = ~n17187 & n17643;
  assign n17647 = n16908 & ~n34576;
  assign n17648 = n16912 & n17644;
  assign n17649 = ~n16900 & n16908;
  assign n17650 = ~n34479 & n17649;
  assign n17651 = ~n17187 & n17650;
  assign n17652 = ~n16908 & ~n34576;
  assign n17653 = ~n17651 & ~n17652;
  assign n17654 = ~n17647 & ~n17648;
  assign n17655 = ~n17642 & ~n34577;
  assign n17656 = ~n17640 & ~n17655;
  assign n17657 = ~n1812 & ~n17656;
  assign n17658 = ~n16914 & ~n16916;
  assign n17659 = ~n17187 & n17658;
  assign n17660 = ~n34481 & ~n17659;
  assign n17661 = ~n16916 & n34481;
  assign n17662 = ~n16914 & n17661;
  assign n17663 = n34481 & n17659;
  assign n17664 = ~n17187 & n17662;
  assign n17665 = ~n17660 & ~n34578;
  assign n17666 = n1812 & ~n17640;
  assign n17667 = n1812 & n17656;
  assign n17668 = ~n17655 & n17666;
  assign n17669 = ~n17665 & ~n34579;
  assign n17670 = ~n17657 & ~n17669;
  assign n17671 = ~n1582 & ~n17670;
  assign n17672 = n1582 & ~n17657;
  assign n17673 = ~n17669 & n17672;
  assign n17674 = ~n16931 & ~n34483;
  assign n17675 = ~n16931 & ~n17187;
  assign n17676 = ~n34483 & n17675;
  assign n17677 = ~n17187 & n17674;
  assign n17678 = n16939 & ~n34580;
  assign n17679 = n16943 & n17675;
  assign n17680 = ~n16931 & n16939;
  assign n17681 = ~n34483 & n17680;
  assign n17682 = ~n17187 & n17681;
  assign n17683 = ~n16939 & ~n34580;
  assign n17684 = ~n17682 & ~n17683;
  assign n17685 = ~n17678 & ~n17679;
  assign n17686 = ~n17673 & ~n34581;
  assign n17687 = ~n17671 & ~n17686;
  assign n17688 = ~n1388 & ~n17687;
  assign n17689 = ~n16945 & ~n16947;
  assign n17690 = ~n17187 & n17689;
  assign n17691 = ~n34485 & ~n17690;
  assign n17692 = ~n16947 & n34485;
  assign n17693 = ~n16945 & n17692;
  assign n17694 = n34485 & n17690;
  assign n17695 = ~n17187 & n17693;
  assign n17696 = ~n17691 & ~n34582;
  assign n17697 = n1388 & ~n17671;
  assign n17698 = n1388 & n17687;
  assign n17699 = ~n17686 & n17697;
  assign n17700 = ~n17696 & ~n34583;
  assign n17701 = ~n17688 & ~n17700;
  assign n17702 = ~n1192 & ~n17701;
  assign n17703 = ~n16962 & ~n34486;
  assign n17704 = ~n17187 & n17703;
  assign n17705 = ~n34488 & ~n17704;
  assign n17706 = ~n16962 & n34488;
  assign n17707 = ~n34486 & n17706;
  assign n17708 = n34488 & n17704;
  assign n17709 = ~n17187 & n17707;
  assign n17710 = ~n17705 & ~n34584;
  assign n17711 = n1192 & ~n17688;
  assign n17712 = ~n17700 & n17711;
  assign n17713 = ~n17710 & ~n17712;
  assign n17714 = ~n17702 & ~n17713;
  assign n17715 = ~n1028 & ~n17714;
  assign n17716 = ~n16980 & ~n16982;
  assign n17717 = ~n17187 & n17716;
  assign n17718 = ~n34490 & ~n17717;
  assign n17719 = ~n16982 & n34490;
  assign n17720 = ~n16980 & n17719;
  assign n17721 = n34490 & n17717;
  assign n17722 = ~n17187 & n17720;
  assign n17723 = ~n17718 & ~n34585;
  assign n17724 = n1028 & ~n17702;
  assign n17725 = n1028 & n17714;
  assign n17726 = ~n17713 & n17724;
  assign n17727 = ~n17723 & ~n34586;
  assign n17728 = ~n17715 & ~n17727;
  assign n17729 = ~n866 & ~n17728;
  assign n17730 = n866 & ~n17715;
  assign n17731 = ~n17727 & n17730;
  assign n17732 = ~n16997 & ~n34492;
  assign n17733 = ~n16997 & ~n17187;
  assign n17734 = ~n34492 & n17733;
  assign n17735 = ~n17187 & n17732;
  assign n17736 = n17005 & ~n34587;
  assign n17737 = n17009 & n17733;
  assign n17738 = ~n16997 & n17005;
  assign n17739 = ~n34492 & n17738;
  assign n17740 = ~n17187 & n17739;
  assign n17741 = ~n17005 & ~n34587;
  assign n17742 = ~n17740 & ~n17741;
  assign n17743 = ~n17736 & ~n17737;
  assign n17744 = ~n17731 & ~n34588;
  assign n17745 = ~n17729 & ~n17744;
  assign n17746 = ~n730 & ~n17745;
  assign n17747 = ~n17011 & ~n17013;
  assign n17748 = ~n17187 & n17747;
  assign n17749 = ~n34494 & ~n17748;
  assign n17750 = ~n17013 & n34494;
  assign n17751 = ~n17011 & n17750;
  assign n17752 = n34494 & n17748;
  assign n17753 = ~n17187 & n17751;
  assign n17754 = ~n17749 & ~n34589;
  assign n17755 = n730 & ~n17729;
  assign n17756 = n730 & n17745;
  assign n17757 = ~n17744 & n17755;
  assign n17758 = ~n17754 & ~n34590;
  assign n17759 = ~n17746 & ~n17758;
  assign n17760 = ~n602 & ~n17759;
  assign n17761 = ~n17028 & ~n34495;
  assign n17762 = ~n17187 & n17761;
  assign n17763 = ~n34497 & ~n17762;
  assign n17764 = ~n17028 & n34497;
  assign n17765 = ~n34495 & n17764;
  assign n17766 = n34497 & n17762;
  assign n17767 = ~n17187 & n17765;
  assign n17768 = ~n17763 & ~n34591;
  assign n17769 = n602 & ~n17746;
  assign n17770 = ~n17758 & n17769;
  assign n17771 = ~n17768 & ~n17770;
  assign n17772 = ~n17760 & ~n17771;
  assign n17773 = ~n497 & ~n17772;
  assign n17774 = ~n17046 & ~n17048;
  assign n17775 = ~n17187 & n17774;
  assign n17776 = ~n34499 & ~n17775;
  assign n17777 = ~n17048 & n34499;
  assign n17778 = ~n17046 & n17777;
  assign n17779 = n34499 & n17775;
  assign n17780 = ~n17187 & n17778;
  assign n17781 = ~n17776 & ~n34592;
  assign n17782 = n497 & ~n17760;
  assign n17783 = n497 & n17772;
  assign n17784 = ~n17771 & n17782;
  assign n17785 = ~n17781 & ~n34593;
  assign n17786 = ~n17773 & ~n17785;
  assign n17787 = ~n403 & ~n17786;
  assign n17788 = n403 & ~n17773;
  assign n17789 = ~n17785 & n17788;
  assign n17790 = ~n17063 & ~n34501;
  assign n17791 = ~n17063 & ~n17187;
  assign n17792 = ~n34501 & n17791;
  assign n17793 = ~n17187 & n17790;
  assign n17794 = n17071 & ~n34594;
  assign n17795 = n17075 & n17791;
  assign n17796 = ~n17063 & n17071;
  assign n17797 = ~n34501 & n17796;
  assign n17798 = ~n17187 & n17797;
  assign n17799 = ~n17071 & ~n34594;
  assign n17800 = ~n17798 & ~n17799;
  assign n17801 = ~n17794 & ~n17795;
  assign n17802 = ~n17789 & ~n34595;
  assign n17803 = ~n17787 & ~n17802;
  assign n17804 = ~n330 & ~n17803;
  assign n17805 = ~n17077 & ~n17079;
  assign n17806 = ~n17187 & n17805;
  assign n17807 = ~n34503 & ~n17806;
  assign n17808 = ~n17079 & n34503;
  assign n17809 = ~n17077 & n17808;
  assign n17810 = n34503 & n17806;
  assign n17811 = ~n17187 & n17809;
  assign n17812 = ~n17807 & ~n34596;
  assign n17813 = n330 & ~n17787;
  assign n17814 = n330 & n17803;
  assign n17815 = ~n17802 & n17813;
  assign n17816 = ~n17812 & ~n34597;
  assign n17817 = ~n17804 & ~n17816;
  assign n17818 = ~n271 & ~n17817;
  assign n17819 = ~n17094 & ~n34504;
  assign n17820 = ~n17187 & n17819;
  assign n17821 = ~n34506 & ~n17820;
  assign n17822 = ~n17094 & n34506;
  assign n17823 = ~n34504 & n17822;
  assign n17824 = n34506 & n17820;
  assign n17825 = ~n17187 & n17823;
  assign n17826 = ~n17821 & ~n34598;
  assign n17827 = n271 & ~n17804;
  assign n17828 = ~n17816 & n17827;
  assign n17829 = ~n17826 & ~n17828;
  assign n17830 = ~n17818 & ~n17829;
  assign n17831 = ~n217 & ~n17830;
  assign n17832 = ~n17112 & ~n17114;
  assign n17833 = ~n17187 & n17832;
  assign n17834 = ~n34508 & ~n17833;
  assign n17835 = ~n17114 & n34508;
  assign n17836 = ~n17112 & n17835;
  assign n17837 = n34508 & n17833;
  assign n17838 = ~n17187 & n17836;
  assign n17839 = ~n17834 & ~n34599;
  assign n17840 = n217 & ~n17818;
  assign n17841 = n217 & n17830;
  assign n17842 = ~n17829 & n17840;
  assign n17843 = ~n17839 & ~n34600;
  assign n17844 = ~n17831 & ~n17843;
  assign n17845 = ~n198 & ~n17844;
  assign n17846 = n198 & ~n17831;
  assign n17847 = ~n17843 & n17846;
  assign n17848 = ~n17129 & ~n34510;
  assign n17849 = ~n17129 & ~n17187;
  assign n17850 = ~n34510 & n17849;
  assign n17851 = ~n17187 & n17848;
  assign n17852 = n17137 & ~n34601;
  assign n17853 = n17141 & n17849;
  assign n17854 = ~n17129 & n17137;
  assign n17855 = ~n34510 & n17854;
  assign n17856 = ~n17187 & n17855;
  assign n17857 = ~n17137 & ~n34601;
  assign n17858 = ~n17856 & ~n17857;
  assign n17859 = ~n17852 & ~n17853;
  assign n17860 = ~n17847 & ~n34602;
  assign n17861 = ~n17845 & ~n17860;
  assign n17862 = ~n17143 & ~n17145;
  assign n17863 = ~n17187 & n17862;
  assign n17864 = ~n34512 & ~n17863;
  assign n17865 = ~n17145 & n34512;
  assign n17866 = ~n17143 & n17865;
  assign n17867 = n34512 & n17863;
  assign n17868 = ~n17187 & n17866;
  assign n17869 = ~n17864 & ~n34603;
  assign n17870 = ~n17159 & ~n34514;
  assign n17871 = ~n34514 & ~n17187;
  assign n17872 = ~n17159 & n17871;
  assign n17873 = ~n17187 & n17870;
  assign n17874 = ~n34516 & ~n34604;
  assign n17875 = ~n17869 & n17874;
  assign n17876 = ~n17861 & n17875;
  assign n17877 = n193 & ~n17876;
  assign n17878 = ~n17845 & n17869;
  assign n17879 = n17861 & n17869;
  assign n17880 = ~n17860 & n17878;
  assign n17881 = n17159 & ~n17871;
  assign n17882 = ~n193 & ~n17870;
  assign n17883 = ~n17881 & n17882;
  assign n17884 = ~n34605 & ~n17883;
  assign n17885 = ~n17877 & n17884;
  assign n17886 = ~n17634 & ~n34575;
  assign n17887 = ~n17634 & ~n17885;
  assign n17888 = ~n34575 & n17887;
  assign n17889 = ~n17885 & n17886;
  assign n17890 = n17195 & ~n34606;
  assign n17891 = n17638 & n17887;
  assign n17892 = n17195 & ~n34575;
  assign n17893 = ~n17634 & n17892;
  assign n17894 = ~n17885 & n17893;
  assign n17895 = ~n17195 & ~n34606;
  assign n17896 = ~n17894 & ~n17895;
  assign n17897 = ~n17890 & ~n17891;
  assign n17898 = pi32  & ~n17885;
  assign n17899 = ~pi30  & ~pi31 ;
  assign n17900 = ~pi32  & n17899;
  assign n17901 = ~n17898 & ~n17900;
  assign n17902 = ~n17187 & ~n17901;
  assign n17903 = ~pi32  & ~n17885;
  assign n17904 = pi33  & ~n17903;
  assign n17905 = ~pi33  & n17903;
  assign n17906 = n17329 & ~n17885;
  assign n17907 = ~n17904 & ~n34608;
  assign n17908 = ~n34409 & ~n34535;
  assign n17909 = ~n16407 & n17908;
  assign n17910 = ~n16426 & n17909;
  assign n17911 = ~n34411 & n17910;
  assign n17912 = n16412 & n16428;
  assign n17913 = ~n16420 & n17911;
  assign n17914 = ~n17900 & ~n34609;
  assign n17915 = ~n17185 & n17914;
  assign n17916 = ~n34516 & n17915;
  assign n17917 = ~n17179 & n17916;
  assign n17918 = n17187 & n17901;
  assign n17919 = ~n17898 & n17917;
  assign n17920 = n17907 & ~n34610;
  assign n17921 = ~n17902 & ~n17920;
  assign n17922 = ~n16428 & ~n17921;
  assign n17923 = n16428 & ~n17902;
  assign n17924 = ~n17920 & n17923;
  assign n17925 = ~n17187 & ~n17883;
  assign n17926 = ~n34605 & n17925;
  assign n17927 = ~n17877 & n17926;
  assign n17928 = ~n34608 & ~n17927;
  assign n17929 = pi34  & ~n17928;
  assign n17930 = ~pi34  & ~n17927;
  assign n17931 = ~pi34  & n17928;
  assign n17932 = ~n34608 & n17930;
  assign n17933 = ~n17929 & ~n34611;
  assign n17934 = ~n17924 & ~n17933;
  assign n17935 = ~n17922 & ~n17934;
  assign n17936 = ~n15760 & ~n17935;
  assign n17937 = n15760 & ~n17922;
  assign n17938 = ~n17934 & n17937;
  assign n17939 = n15760 & n17935;
  assign n17940 = ~n34536 & ~n17347;
  assign n17941 = ~n17885 & n17940;
  assign n17942 = n17345 & ~n17941;
  assign n17943 = ~n17345 & n17940;
  assign n17944 = ~n17345 & n17941;
  assign n17945 = ~n17885 & n17943;
  assign n17946 = ~n17942 & ~n34613;
  assign n17947 = ~n34612 & ~n17946;
  assign n17948 = ~n17936 & ~n17947;
  assign n17949 = ~n15033 & ~n17948;
  assign n17950 = n15033 & ~n17936;
  assign n17951 = ~n17947 & n17950;
  assign n17952 = ~n34537 & ~n17353;
  assign n17953 = ~n17353 & ~n17885;
  assign n17954 = ~n34537 & n17953;
  assign n17955 = ~n17885 & n17952;
  assign n17956 = n17327 & ~n34614;
  assign n17957 = n17352 & n17953;
  assign n17958 = n17327 & ~n34537;
  assign n17959 = ~n17353 & n17958;
  assign n17960 = ~n17885 & n17959;
  assign n17961 = ~n17327 & ~n34614;
  assign n17962 = ~n17960 & ~n17961;
  assign n17963 = ~n17956 & ~n17957;
  assign n17964 = ~n17951 & ~n34615;
  assign n17965 = ~n17949 & ~n17964;
  assign n17966 = ~n14394 & ~n17965;
  assign n17967 = n14394 & ~n17949;
  assign n17968 = ~n17964 & n17967;
  assign n17969 = n14394 & n17965;
  assign n17970 = ~n17355 & ~n17365;
  assign n17971 = ~n17885 & n17970;
  assign n17972 = n17362 & ~n17971;
  assign n17973 = ~n17362 & n17971;
  assign n17974 = n17362 & ~n17365;
  assign n17975 = ~n17355 & n17974;
  assign n17976 = n17362 & n17971;
  assign n17977 = ~n17885 & n17975;
  assign n17978 = ~n17362 & ~n17971;
  assign n17979 = ~n34617 & ~n17978;
  assign n17980 = ~n17972 & ~n17973;
  assign n17981 = ~n34616 & ~n34618;
  assign n17982 = ~n17966 & ~n17981;
  assign n17983 = ~n13704 & ~n17982;
  assign n17984 = n13704 & ~n17966;
  assign n17985 = ~n17981 & n17984;
  assign n17986 = ~n34539 & ~n17371;
  assign n17987 = ~n17371 & ~n17885;
  assign n17988 = ~n34539 & n17987;
  assign n17989 = ~n17885 & n17986;
  assign n17990 = n17315 & ~n34619;
  assign n17991 = n17370 & n17987;
  assign n17992 = n17315 & ~n34539;
  assign n17993 = ~n17371 & n17992;
  assign n17994 = ~n17885 & n17993;
  assign n17995 = ~n17315 & ~n34619;
  assign n17996 = ~n17994 & ~n17995;
  assign n17997 = ~n17990 & ~n17991;
  assign n17998 = ~n17985 & ~n34620;
  assign n17999 = ~n17983 & ~n17998;
  assign n18000 = ~n13099 & ~n17999;
  assign n18001 = n13099 & ~n17983;
  assign n18002 = ~n17998 & n18001;
  assign n18003 = n13099 & n17999;
  assign n18004 = ~n17373 & ~n17387;
  assign n18005 = ~n17885 & n18004;
  assign n18006 = ~n34541 & n18005;
  assign n18007 = n34541 & ~n18005;
  assign n18008 = n34541 & ~n17387;
  assign n18009 = ~n17373 & n18008;
  assign n18010 = ~n17885 & n18009;
  assign n18011 = ~n34541 & ~n18005;
  assign n18012 = ~n18010 & ~n18011;
  assign n18013 = ~n18006 & ~n18007;
  assign n18014 = ~n34621 & ~n34622;
  assign n18015 = ~n18000 & ~n18014;
  assign n18016 = ~n12442 & ~n18015;
  assign n18017 = n12442 & ~n18000;
  assign n18018 = ~n18014 & n18017;
  assign n18019 = ~n34542 & ~n17393;
  assign n18020 = ~n17393 & ~n17885;
  assign n18021 = ~n34542 & n18020;
  assign n18022 = ~n17885 & n18019;
  assign n18023 = n17307 & ~n34623;
  assign n18024 = n17392 & n18020;
  assign n18025 = n17307 & ~n34542;
  assign n18026 = ~n17393 & n18025;
  assign n18027 = ~n17885 & n18026;
  assign n18028 = ~n17307 & ~n34623;
  assign n18029 = ~n18027 & ~n18028;
  assign n18030 = ~n18023 & ~n18024;
  assign n18031 = ~n18018 & ~n34624;
  assign n18032 = ~n18016 & ~n18031;
  assign n18033 = ~n11858 & ~n18032;
  assign n18034 = n11858 & ~n18016;
  assign n18035 = ~n18031 & n18034;
  assign n18036 = n11858 & n18032;
  assign n18037 = ~n17395 & ~n17408;
  assign n18038 = ~n17885 & n18037;
  assign n18039 = ~n34543 & ~n18038;
  assign n18040 = n34543 & ~n17408;
  assign n18041 = ~n17395 & n18040;
  assign n18042 = n34543 & n18038;
  assign n18043 = ~n17885 & n18041;
  assign n18044 = n34543 & ~n18038;
  assign n18045 = ~n34543 & n18038;
  assign n18046 = ~n18044 & ~n18045;
  assign n18047 = ~n18039 & ~n34626;
  assign n18048 = ~n34625 & n34627;
  assign n18049 = ~n18033 & ~n18048;
  assign n18050 = ~n11229 & ~n18049;
  assign n18051 = n11229 & ~n18033;
  assign n18052 = ~n18048 & n18051;
  assign n18053 = ~n34544 & ~n17414;
  assign n18054 = ~n17414 & ~n17885;
  assign n18055 = ~n34544 & n18054;
  assign n18056 = ~n17885 & n18053;
  assign n18057 = n17299 & ~n34628;
  assign n18058 = n17413 & n18054;
  assign n18059 = n17299 & ~n34544;
  assign n18060 = ~n17414 & n18059;
  assign n18061 = ~n17885 & n18060;
  assign n18062 = ~n17299 & ~n34628;
  assign n18063 = ~n18061 & ~n18062;
  assign n18064 = ~n18057 & ~n18058;
  assign n18065 = ~n18052 & ~n34629;
  assign n18066 = ~n18050 & ~n18065;
  assign n18067 = ~n10681 & ~n18066;
  assign n18068 = n10681 & ~n18050;
  assign n18069 = ~n18065 & n18068;
  assign n18070 = n10681 & n18066;
  assign n18071 = ~n17416 & ~n17430;
  assign n18072 = ~n17885 & n18071;
  assign n18073 = n34546 & ~n18072;
  assign n18074 = ~n34546 & ~n17430;
  assign n18075 = ~n17416 & n18074;
  assign n18076 = ~n34546 & n18072;
  assign n18077 = ~n17885 & n18075;
  assign n18078 = n34546 & n18072;
  assign n18079 = ~n34546 & ~n18072;
  assign n18080 = ~n18078 & ~n18079;
  assign n18081 = ~n18073 & ~n34631;
  assign n18082 = ~n34630 & n34632;
  assign n18083 = ~n18067 & ~n18082;
  assign n18084 = ~n10086 & ~n18083;
  assign n18085 = n10086 & ~n18067;
  assign n18086 = ~n18082 & n18085;
  assign n18087 = ~n34547 & ~n17436;
  assign n18088 = ~n17436 & ~n17885;
  assign n18089 = ~n34547 & n18088;
  assign n18090 = ~n17885 & n18087;
  assign n18091 = n17291 & ~n34633;
  assign n18092 = n17435 & n18088;
  assign n18093 = n17291 & ~n34547;
  assign n18094 = ~n17436 & n18093;
  assign n18095 = ~n17885 & n18094;
  assign n18096 = ~n17291 & ~n34633;
  assign n18097 = ~n18095 & ~n18096;
  assign n18098 = ~n18091 & ~n18092;
  assign n18099 = ~n18086 & ~n34634;
  assign n18100 = ~n18084 & ~n18099;
  assign n18101 = ~n9565 & ~n18100;
  assign n18102 = n9565 & ~n18084;
  assign n18103 = ~n18099 & n18102;
  assign n18104 = n9565 & n18100;
  assign n18105 = ~n17438 & ~n17452;
  assign n18106 = ~n17452 & ~n17885;
  assign n18107 = ~n17438 & n18106;
  assign n18108 = ~n17885 & n18105;
  assign n18109 = ~n34549 & ~n34636;
  assign n18110 = n17450 & n18106;
  assign n18111 = n34549 & n34636;
  assign n18112 = ~n34549 & ~n17452;
  assign n18113 = ~n17438 & n18112;
  assign n18114 = ~n17885 & n18113;
  assign n18115 = n34549 & ~n34636;
  assign n18116 = ~n18114 & ~n18115;
  assign n18117 = ~n18109 & ~n34637;
  assign n18118 = ~n34635 & ~n34638;
  assign n18119 = ~n18101 & ~n18118;
  assign n18120 = ~n8998 & ~n18119;
  assign n18121 = n8998 & ~n18101;
  assign n18122 = ~n18118 & n18121;
  assign n18123 = ~n34550 & ~n17458;
  assign n18124 = ~n17458 & ~n17885;
  assign n18125 = ~n34550 & n18124;
  assign n18126 = ~n17885 & n18123;
  assign n18127 = n17283 & ~n34639;
  assign n18128 = n17457 & n18124;
  assign n18129 = n17283 & ~n34550;
  assign n18130 = ~n17458 & n18129;
  assign n18131 = ~n17885 & n18130;
  assign n18132 = ~n17283 & ~n34639;
  assign n18133 = ~n18131 & ~n18132;
  assign n18134 = ~n18127 & ~n18128;
  assign n18135 = ~n18122 & ~n34640;
  assign n18136 = ~n18120 & ~n18135;
  assign n18137 = ~n8506 & ~n18136;
  assign n18138 = n8506 & ~n18120;
  assign n18139 = ~n18135 & n18138;
  assign n18140 = n8506 & n18136;
  assign n18141 = ~n17460 & ~n17476;
  assign n18142 = ~n17885 & n18141;
  assign n18143 = ~n34553 & ~n18142;
  assign n18144 = n34553 & ~n17476;
  assign n18145 = ~n17460 & n18144;
  assign n18146 = n34553 & n18142;
  assign n18147 = ~n17885 & n18145;
  assign n18148 = ~n18143 & ~n34642;
  assign n18149 = ~n34641 & ~n18148;
  assign n18150 = ~n18137 & ~n18149;
  assign n18151 = ~n7975 & ~n18150;
  assign n18152 = n7975 & ~n18137;
  assign n18153 = ~n18149 & n18152;
  assign n18154 = ~n34554 & ~n17482;
  assign n18155 = ~n17482 & ~n17885;
  assign n18156 = ~n34554 & n18155;
  assign n18157 = ~n17885 & n18154;
  assign n18158 = n17275 & ~n34643;
  assign n18159 = n17481 & n18155;
  assign n18160 = n17275 & ~n34554;
  assign n18161 = ~n17482 & n18160;
  assign n18162 = ~n17885 & n18161;
  assign n18163 = ~n17275 & ~n34643;
  assign n18164 = ~n18162 & ~n18163;
  assign n18165 = ~n18158 & ~n18159;
  assign n18166 = ~n18153 & ~n34644;
  assign n18167 = ~n18151 & ~n18166;
  assign n18168 = ~n7512 & ~n18167;
  assign n18169 = n7512 & ~n18151;
  assign n18170 = ~n18166 & n18169;
  assign n18171 = n7512 & n18167;
  assign n18172 = ~n17484 & ~n17495;
  assign n18173 = ~n17495 & ~n17885;
  assign n18174 = ~n17484 & n18173;
  assign n18175 = ~n17885 & n18172;
  assign n18176 = n17492 & ~n34646;
  assign n18177 = n17493 & n18173;
  assign n18178 = ~n17492 & n34646;
  assign n18179 = n17492 & ~n17495;
  assign n18180 = ~n17484 & n18179;
  assign n18181 = ~n17885 & n18180;
  assign n18182 = ~n17492 & ~n34646;
  assign n18183 = ~n18181 & ~n18182;
  assign n18184 = ~n18176 & ~n34647;
  assign n18185 = ~n34645 & ~n34648;
  assign n18186 = ~n18168 & ~n18185;
  assign n18187 = ~n7015 & ~n18186;
  assign n18188 = n7015 & ~n18168;
  assign n18189 = ~n18185 & n18188;
  assign n18190 = ~n34556 & ~n17501;
  assign n18191 = ~n17501 & ~n17885;
  assign n18192 = ~n34556 & n18191;
  assign n18193 = ~n17885 & n18190;
  assign n18194 = n17267 & ~n34649;
  assign n18195 = n17500 & n18191;
  assign n18196 = n17267 & ~n34556;
  assign n18197 = ~n17501 & n18196;
  assign n18198 = ~n17885 & n18197;
  assign n18199 = ~n17267 & ~n34649;
  assign n18200 = ~n18198 & ~n18199;
  assign n18201 = ~n18194 & ~n18195;
  assign n18202 = ~n18189 & ~n34650;
  assign n18203 = ~n18187 & ~n18202;
  assign n18204 = ~n6579 & ~n18203;
  assign n18205 = n6579 & ~n18187;
  assign n18206 = ~n18202 & n18205;
  assign n18207 = n6579 & n18203;
  assign n18208 = ~n17503 & ~n17519;
  assign n18209 = ~n17885 & n18208;
  assign n18210 = ~n34559 & n18209;
  assign n18211 = n34559 & ~n18209;
  assign n18212 = n34559 & ~n17519;
  assign n18213 = ~n17503 & n18212;
  assign n18214 = n34559 & n18209;
  assign n18215 = ~n17885 & n18213;
  assign n18216 = ~n34559 & ~n18209;
  assign n18217 = ~n34652 & ~n18216;
  assign n18218 = ~n18210 & ~n18211;
  assign n18219 = ~n34651 & ~n34653;
  assign n18220 = ~n18204 & ~n18219;
  assign n18221 = ~n6117 & ~n18220;
  assign n18222 = n6117 & ~n18204;
  assign n18223 = ~n18219 & n18222;
  assign n18224 = ~n34560 & ~n17525;
  assign n18225 = ~n17525 & ~n17885;
  assign n18226 = ~n34560 & n18225;
  assign n18227 = ~n17885 & n18224;
  assign n18228 = n17259 & ~n34654;
  assign n18229 = n17524 & n18225;
  assign n18230 = n17259 & ~n34560;
  assign n18231 = ~n17525 & n18230;
  assign n18232 = ~n17885 & n18231;
  assign n18233 = ~n17259 & ~n34654;
  assign n18234 = ~n18232 & ~n18233;
  assign n18235 = ~n18228 & ~n18229;
  assign n18236 = ~n18223 & ~n34655;
  assign n18237 = ~n18221 & ~n18236;
  assign n18238 = ~n5708 & ~n18237;
  assign n18239 = n5708 & ~n18221;
  assign n18240 = ~n18236 & n18239;
  assign n18241 = n5708 & n18237;
  assign n18242 = ~n17527 & ~n17541;
  assign n18243 = ~n17541 & ~n17885;
  assign n18244 = ~n17527 & n18243;
  assign n18245 = ~n17885 & n18242;
  assign n18246 = n34562 & ~n34657;
  assign n18247 = n17539 & n18243;
  assign n18248 = ~n34562 & n34657;
  assign n18249 = n34562 & ~n17541;
  assign n18250 = ~n17527 & n18249;
  assign n18251 = ~n17885 & n18250;
  assign n18252 = ~n34562 & ~n34657;
  assign n18253 = ~n18251 & ~n18252;
  assign n18254 = ~n18246 & ~n34658;
  assign n18255 = ~n34656 & ~n34659;
  assign n18256 = ~n18238 & ~n18255;
  assign n18257 = ~n5278 & ~n18256;
  assign n18258 = n5278 & ~n18238;
  assign n18259 = ~n18255 & n18258;
  assign n18260 = ~n34563 & ~n17547;
  assign n18261 = ~n17547 & ~n17885;
  assign n18262 = ~n34563 & n18261;
  assign n18263 = ~n17885 & n18260;
  assign n18264 = n17251 & ~n34660;
  assign n18265 = n17546 & n18261;
  assign n18266 = n17251 & ~n34563;
  assign n18267 = ~n17547 & n18266;
  assign n18268 = ~n17885 & n18267;
  assign n18269 = ~n17251 & ~n34660;
  assign n18270 = ~n18268 & ~n18269;
  assign n18271 = ~n18264 & ~n18265;
  assign n18272 = ~n18259 & ~n34661;
  assign n18273 = ~n18257 & ~n18272;
  assign n18274 = ~n4903 & ~n18273;
  assign n18275 = ~n17549 & ~n17565;
  assign n18276 = ~n17885 & n18275;
  assign n18277 = ~n34566 & ~n18276;
  assign n18278 = n34566 & ~n17565;
  assign n18279 = ~n17549 & n18278;
  assign n18280 = n34566 & n18276;
  assign n18281 = ~n17885 & n18279;
  assign n18282 = ~n18277 & ~n34662;
  assign n18283 = n4903 & ~n18257;
  assign n18284 = ~n18272 & n18283;
  assign n18285 = n4903 & n18273;
  assign n18286 = ~n18282 & ~n34663;
  assign n18287 = ~n18274 & ~n18286;
  assign n18288 = ~n4508 & ~n18287;
  assign n18289 = n4508 & ~n18274;
  assign n18290 = ~n18286 & n18289;
  assign n18291 = ~n34567 & ~n17571;
  assign n18292 = ~n17571 & ~n17885;
  assign n18293 = ~n34567 & n18292;
  assign n18294 = ~n17885 & n18291;
  assign n18295 = n17243 & ~n34664;
  assign n18296 = n17570 & n18292;
  assign n18297 = n17243 & ~n34567;
  assign n18298 = ~n17571 & n18297;
  assign n18299 = ~n17885 & n18298;
  assign n18300 = ~n17243 & ~n34664;
  assign n18301 = ~n18299 & ~n18300;
  assign n18302 = ~n18295 & ~n18296;
  assign n18303 = ~n18290 & ~n34665;
  assign n18304 = ~n18288 & ~n18303;
  assign n18305 = ~n4155 & ~n18304;
  assign n18306 = n4155 & ~n18288;
  assign n18307 = ~n18303 & n18306;
  assign n18308 = n4155 & n18304;
  assign n18309 = ~n17573 & ~n17576;
  assign n18310 = ~n17576 & ~n17885;
  assign n18311 = ~n17573 & n18310;
  assign n18312 = ~n17885 & n18309;
  assign n18313 = n17235 & ~n34667;
  assign n18314 = n17574 & n18310;
  assign n18315 = n17235 & ~n17576;
  assign n18316 = ~n17573 & n18315;
  assign n18317 = ~n17885 & n18316;
  assign n18318 = ~n17235 & ~n34667;
  assign n18319 = ~n18317 & ~n18318;
  assign n18320 = ~n18313 & ~n18314;
  assign n18321 = ~n34666 & ~n34668;
  assign n18322 = ~n18305 & ~n18321;
  assign n18323 = ~n3788 & ~n18322;
  assign n18324 = n3788 & ~n18305;
  assign n18325 = ~n18321 & n18324;
  assign n18326 = ~n34568 & ~n17582;
  assign n18327 = ~n17582 & ~n17885;
  assign n18328 = ~n34568 & n18327;
  assign n18329 = ~n17885 & n18326;
  assign n18330 = n17227 & ~n34669;
  assign n18331 = n17581 & n18327;
  assign n18332 = n17227 & ~n34568;
  assign n18333 = ~n17582 & n18332;
  assign n18334 = ~n17885 & n18333;
  assign n18335 = ~n17227 & ~n34669;
  assign n18336 = ~n18334 & ~n18335;
  assign n18337 = ~n18330 & ~n18331;
  assign n18338 = ~n18325 & ~n34670;
  assign n18339 = ~n18323 & ~n18338;
  assign n18340 = ~n3473 & ~n18339;
  assign n18341 = ~n17584 & ~n17599;
  assign n18342 = ~n17885 & n18341;
  assign n18343 = ~n34570 & ~n18342;
  assign n18344 = n34570 & ~n17599;
  assign n18345 = ~n17584 & n18344;
  assign n18346 = n34570 & n18342;
  assign n18347 = ~n17885 & n18345;
  assign n18348 = ~n18343 & ~n34671;
  assign n18349 = n3473 & ~n18323;
  assign n18350 = ~n18338 & n18349;
  assign n18351 = n3473 & n18339;
  assign n18352 = ~n18348 & ~n34672;
  assign n18353 = ~n18340 & ~n18352;
  assign n18354 = ~n3140 & ~n18353;
  assign n18355 = n3140 & ~n18340;
  assign n18356 = ~n18352 & n18355;
  assign n18357 = ~n34571 & ~n17605;
  assign n18358 = ~n17605 & ~n17885;
  assign n18359 = ~n34571 & n18358;
  assign n18360 = ~n17885 & n18357;
  assign n18361 = n17219 & ~n34673;
  assign n18362 = n17604 & n18358;
  assign n18363 = n17219 & ~n34571;
  assign n18364 = ~n17605 & n18363;
  assign n18365 = ~n17885 & n18364;
  assign n18366 = ~n17219 & ~n34673;
  assign n18367 = ~n18365 & ~n18366;
  assign n18368 = ~n18361 & ~n18362;
  assign n18369 = ~n18356 & ~n34674;
  assign n18370 = ~n18354 & ~n18369;
  assign n18371 = ~n2855 & ~n18370;
  assign n18372 = n2855 & ~n18354;
  assign n18373 = ~n18369 & n18372;
  assign n18374 = n2855 & n18370;
  assign n18375 = ~n17607 & ~n17610;
  assign n18376 = ~n17610 & ~n17885;
  assign n18377 = ~n17607 & n18376;
  assign n18378 = ~n17885 & n18375;
  assign n18379 = n17211 & ~n34676;
  assign n18380 = n17608 & n18376;
  assign n18381 = n17211 & ~n17610;
  assign n18382 = ~n17607 & n18381;
  assign n18383 = ~n17885 & n18382;
  assign n18384 = ~n17211 & ~n34676;
  assign n18385 = ~n18383 & ~n18384;
  assign n18386 = ~n18379 & ~n18380;
  assign n18387 = ~n34675 & ~n34677;
  assign n18388 = ~n18371 & ~n18387;
  assign n18389 = ~n2556 & ~n18388;
  assign n18390 = n2556 & ~n18371;
  assign n18391 = ~n18387 & n18390;
  assign n18392 = n17203 & ~n34572;
  assign n18393 = ~n17616 & n18392;
  assign n18394 = ~n34572 & ~n17616;
  assign n18395 = ~n17885 & n18394;
  assign n18396 = n17203 & n18395;
  assign n18397 = ~n17885 & n18393;
  assign n18398 = ~n17203 & ~n18395;
  assign n18399 = ~n34678 & ~n18398;
  assign n18400 = ~n18391 & ~n18399;
  assign n18401 = ~n18389 & ~n18400;
  assign n18402 = ~n2301 & ~n18401;
  assign n18403 = n2301 & ~n18389;
  assign n18404 = ~n18400 & n18403;
  assign n18405 = n2301 & n18401;
  assign n18406 = ~n17618 & ~n17620;
  assign n18407 = ~n17885 & n18406;
  assign n18408 = ~n34574 & n18407;
  assign n18409 = n34574 & ~n18407;
  assign n18410 = ~n17618 & n34574;
  assign n18411 = ~n17620 & n18410;
  assign n18412 = n34574 & n18407;
  assign n18413 = ~n17885 & n18411;
  assign n18414 = ~n34574 & ~n18407;
  assign n18415 = ~n34680 & ~n18414;
  assign n18416 = ~n18408 & ~n18409;
  assign n18417 = ~n34679 & ~n34681;
  assign n18418 = ~n18402 & ~n18417;
  assign n18419 = ~n2038 & ~n18418;
  assign n18420 = n2038 & ~n18402;
  assign n18421 = ~n18417 & n18420;
  assign n18422 = ~n34607 & ~n18421;
  assign n18423 = ~n18419 & ~n18422;
  assign n18424 = ~n1812 & ~n18423;
  assign n18425 = ~n17640 & ~n17642;
  assign n18426 = ~n17885 & n18425;
  assign n18427 = ~n34577 & ~n18426;
  assign n18428 = ~n17640 & n34577;
  assign n18429 = ~n17642 & n18428;
  assign n18430 = n34577 & n18426;
  assign n18431 = ~n17885 & n18429;
  assign n18432 = ~n18427 & ~n34682;
  assign n18433 = n1812 & ~n18419;
  assign n18434 = ~n18422 & n18433;
  assign n18435 = n1812 & n18423;
  assign n18436 = ~n18432 & ~n34683;
  assign n18437 = ~n18424 & ~n18436;
  assign n18438 = ~n1582 & ~n18437;
  assign n18439 = n1582 & ~n18424;
  assign n18440 = ~n18436 & n18439;
  assign n18441 = ~n17657 & ~n34579;
  assign n18442 = ~n17657 & ~n17885;
  assign n18443 = ~n34579 & n18442;
  assign n18444 = ~n17885 & n18441;
  assign n18445 = n17665 & ~n34684;
  assign n18446 = n17669 & n18442;
  assign n18447 = n17665 & ~n34579;
  assign n18448 = ~n17657 & n18447;
  assign n18449 = ~n17885 & n18448;
  assign n18450 = ~n17665 & ~n34684;
  assign n18451 = ~n18449 & ~n18450;
  assign n18452 = ~n18445 & ~n18446;
  assign n18453 = ~n18440 & ~n34685;
  assign n18454 = ~n18438 & ~n18453;
  assign n18455 = ~n1388 & ~n18454;
  assign n18456 = ~n17671 & ~n17673;
  assign n18457 = ~n17885 & n18456;
  assign n18458 = ~n34581 & ~n18457;
  assign n18459 = ~n17671 & n34581;
  assign n18460 = ~n17673 & n18459;
  assign n18461 = n34581 & n18457;
  assign n18462 = ~n17885 & n18460;
  assign n18463 = ~n18458 & ~n34686;
  assign n18464 = n1388 & ~n18438;
  assign n18465 = ~n18453 & n18464;
  assign n18466 = n1388 & n18454;
  assign n18467 = ~n18463 & ~n34687;
  assign n18468 = ~n18455 & ~n18467;
  assign n18469 = ~n1192 & ~n18468;
  assign n18470 = n1192 & ~n18455;
  assign n18471 = ~n18467 & n18470;
  assign n18472 = ~n17688 & ~n34583;
  assign n18473 = ~n17688 & ~n17885;
  assign n18474 = ~n34583 & n18473;
  assign n18475 = ~n17885 & n18472;
  assign n18476 = n17696 & ~n34688;
  assign n18477 = n17700 & n18473;
  assign n18478 = n17696 & ~n34583;
  assign n18479 = ~n17688 & n18478;
  assign n18480 = ~n17885 & n18479;
  assign n18481 = ~n17696 & ~n34688;
  assign n18482 = ~n18480 & ~n18481;
  assign n18483 = ~n18476 & ~n18477;
  assign n18484 = ~n18471 & ~n34689;
  assign n18485 = ~n18469 & ~n18484;
  assign n18486 = ~n1028 & ~n18485;
  assign n18487 = n1028 & ~n18469;
  assign n18488 = ~n18484 & n18487;
  assign n18489 = n1028 & n18485;
  assign n18490 = ~n17702 & ~n17712;
  assign n18491 = ~n17702 & ~n17885;
  assign n18492 = ~n17712 & n18491;
  assign n18493 = ~n17885 & n18490;
  assign n18494 = n17710 & ~n34691;
  assign n18495 = n17713 & n18491;
  assign n18496 = ~n17702 & n17710;
  assign n18497 = ~n17712 & n18496;
  assign n18498 = ~n17885 & n18497;
  assign n18499 = ~n17710 & ~n34691;
  assign n18500 = ~n18498 & ~n18499;
  assign n18501 = ~n18494 & ~n18495;
  assign n18502 = ~n34690 & ~n34692;
  assign n18503 = ~n18486 & ~n18502;
  assign n18504 = ~n866 & ~n18503;
  assign n18505 = n866 & ~n18486;
  assign n18506 = ~n18502 & n18505;
  assign n18507 = ~n17715 & ~n34586;
  assign n18508 = ~n17715 & ~n17885;
  assign n18509 = ~n34586 & n18508;
  assign n18510 = ~n17885 & n18507;
  assign n18511 = n17723 & ~n34693;
  assign n18512 = n17727 & n18508;
  assign n18513 = n17723 & ~n34586;
  assign n18514 = ~n17715 & n18513;
  assign n18515 = ~n17885 & n18514;
  assign n18516 = ~n17723 & ~n34693;
  assign n18517 = ~n18515 & ~n18516;
  assign n18518 = ~n18511 & ~n18512;
  assign n18519 = ~n18506 & ~n34694;
  assign n18520 = ~n18504 & ~n18519;
  assign n18521 = ~n730 & ~n18520;
  assign n18522 = ~n17729 & ~n17731;
  assign n18523 = ~n17885 & n18522;
  assign n18524 = ~n34588 & ~n18523;
  assign n18525 = ~n17729 & n34588;
  assign n18526 = ~n17731 & n18525;
  assign n18527 = n34588 & n18523;
  assign n18528 = ~n17885 & n18526;
  assign n18529 = ~n18524 & ~n34695;
  assign n18530 = n730 & ~n18504;
  assign n18531 = ~n18519 & n18530;
  assign n18532 = n730 & n18520;
  assign n18533 = ~n18529 & ~n34696;
  assign n18534 = ~n18521 & ~n18533;
  assign n18535 = ~n602 & ~n18534;
  assign n18536 = n602 & ~n18521;
  assign n18537 = ~n18533 & n18536;
  assign n18538 = ~n17746 & ~n34590;
  assign n18539 = ~n17746 & ~n17885;
  assign n18540 = ~n34590 & n18539;
  assign n18541 = ~n17885 & n18538;
  assign n18542 = n17754 & ~n34697;
  assign n18543 = n17758 & n18539;
  assign n18544 = n17754 & ~n34590;
  assign n18545 = ~n17746 & n18544;
  assign n18546 = ~n17885 & n18545;
  assign n18547 = ~n17754 & ~n34697;
  assign n18548 = ~n18546 & ~n18547;
  assign n18549 = ~n18542 & ~n18543;
  assign n18550 = ~n18537 & ~n34698;
  assign n18551 = ~n18535 & ~n18550;
  assign n18552 = ~n497 & ~n18551;
  assign n18553 = n497 & ~n18535;
  assign n18554 = ~n18550 & n18553;
  assign n18555 = n497 & n18551;
  assign n18556 = ~n17760 & ~n17770;
  assign n18557 = ~n17760 & ~n17885;
  assign n18558 = ~n17770 & n18557;
  assign n18559 = ~n17885 & n18556;
  assign n18560 = n17768 & ~n34700;
  assign n18561 = n17771 & n18557;
  assign n18562 = ~n17760 & n17768;
  assign n18563 = ~n17770 & n18562;
  assign n18564 = ~n17885 & n18563;
  assign n18565 = ~n17768 & ~n34700;
  assign n18566 = ~n18564 & ~n18565;
  assign n18567 = ~n18560 & ~n18561;
  assign n18568 = ~n34699 & ~n34701;
  assign n18569 = ~n18552 & ~n18568;
  assign n18570 = ~n403 & ~n18569;
  assign n18571 = n403 & ~n18552;
  assign n18572 = ~n18568 & n18571;
  assign n18573 = ~n17773 & ~n34593;
  assign n18574 = ~n17773 & ~n17885;
  assign n18575 = ~n34593 & n18574;
  assign n18576 = ~n17885 & n18573;
  assign n18577 = n17781 & ~n34702;
  assign n18578 = n17785 & n18574;
  assign n18579 = n17781 & ~n34593;
  assign n18580 = ~n17773 & n18579;
  assign n18581 = ~n17885 & n18580;
  assign n18582 = ~n17781 & ~n34702;
  assign n18583 = ~n18581 & ~n18582;
  assign n18584 = ~n18577 & ~n18578;
  assign n18585 = ~n18572 & ~n34703;
  assign n18586 = ~n18570 & ~n18585;
  assign n18587 = ~n330 & ~n18586;
  assign n18588 = ~n17787 & ~n17789;
  assign n18589 = ~n17885 & n18588;
  assign n18590 = ~n34595 & ~n18589;
  assign n18591 = ~n17787 & n34595;
  assign n18592 = ~n17789 & n18591;
  assign n18593 = n34595 & n18589;
  assign n18594 = ~n17885 & n18592;
  assign n18595 = ~n18590 & ~n34704;
  assign n18596 = n330 & ~n18570;
  assign n18597 = ~n18585 & n18596;
  assign n18598 = n330 & n18586;
  assign n18599 = ~n18595 & ~n34705;
  assign n18600 = ~n18587 & ~n18599;
  assign n18601 = ~n271 & ~n18600;
  assign n18602 = n271 & ~n18587;
  assign n18603 = ~n18599 & n18602;
  assign n18604 = ~n17804 & ~n34597;
  assign n18605 = ~n17804 & ~n17885;
  assign n18606 = ~n34597 & n18605;
  assign n18607 = ~n17885 & n18604;
  assign n18608 = n17812 & ~n34706;
  assign n18609 = n17816 & n18605;
  assign n18610 = n17812 & ~n34597;
  assign n18611 = ~n17804 & n18610;
  assign n18612 = ~n17885 & n18611;
  assign n18613 = ~n17812 & ~n34706;
  assign n18614 = ~n18612 & ~n18613;
  assign n18615 = ~n18608 & ~n18609;
  assign n18616 = ~n18603 & ~n34707;
  assign n18617 = ~n18601 & ~n18616;
  assign n18618 = ~n217 & ~n18617;
  assign n18619 = n217 & ~n18601;
  assign n18620 = ~n18616 & n18619;
  assign n18621 = n217 & n18617;
  assign n18622 = ~n17818 & ~n17828;
  assign n18623 = ~n17818 & ~n17885;
  assign n18624 = ~n17828 & n18623;
  assign n18625 = ~n17885 & n18622;
  assign n18626 = n17826 & ~n34709;
  assign n18627 = n17829 & n18623;
  assign n18628 = ~n17818 & n17826;
  assign n18629 = ~n17828 & n18628;
  assign n18630 = ~n17885 & n18629;
  assign n18631 = ~n17826 & ~n34709;
  assign n18632 = ~n18630 & ~n18631;
  assign n18633 = ~n18626 & ~n18627;
  assign n18634 = ~n34708 & ~n34710;
  assign n18635 = ~n18618 & ~n18634;
  assign n18636 = ~n198 & ~n18635;
  assign n18637 = n198 & ~n18618;
  assign n18638 = ~n18634 & n18637;
  assign n18639 = ~n17831 & ~n34600;
  assign n18640 = ~n17831 & ~n17885;
  assign n18641 = ~n34600 & n18640;
  assign n18642 = ~n17885 & n18639;
  assign n18643 = n17839 & ~n34711;
  assign n18644 = n17843 & n18640;
  assign n18645 = n17839 & ~n34600;
  assign n18646 = ~n17831 & n18645;
  assign n18647 = ~n17885 & n18646;
  assign n18648 = ~n17839 & ~n34711;
  assign n18649 = ~n18647 & ~n18648;
  assign n18650 = ~n18643 & ~n18644;
  assign n18651 = ~n18638 & ~n34712;
  assign n18652 = ~n18636 & ~n18651;
  assign n18653 = ~n17845 & ~n17847;
  assign n18654 = ~n17885 & n18653;
  assign n18655 = ~n34602 & ~n18654;
  assign n18656 = ~n17845 & n34602;
  assign n18657 = ~n17847 & n18656;
  assign n18658 = n34602 & n18654;
  assign n18659 = ~n17885 & n18657;
  assign n18660 = ~n18655 & ~n34713;
  assign n18661 = ~n17861 & ~n17869;
  assign n18662 = ~n17869 & ~n17885;
  assign n18663 = ~n17861 & n18662;
  assign n18664 = ~n17885 & n18661;
  assign n18665 = ~n34605 & ~n34714;
  assign n18666 = ~n18660 & n18665;
  assign n18667 = ~n18652 & n18666;
  assign n18668 = n193 & ~n18667;
  assign n18669 = ~n18636 & n18660;
  assign n18670 = ~n18651 & n18669;
  assign n18671 = n18652 & n18660;
  assign n18672 = n17861 & ~n18662;
  assign n18673 = ~n193 & ~n18661;
  assign n18674 = ~n18672 & n18673;
  assign n18675 = ~n34715 & ~n18674;
  assign n18676 = ~n18668 & n18675;
  assign n18677 = ~n18419 & ~n18421;
  assign n18678 = ~n18676 & n18677;
  assign n18679 = ~n34607 & ~n18678;
  assign n18680 = n34607 & ~n18421;
  assign n18681 = ~n18419 & n18680;
  assign n18682 = n34607 & n18678;
  assign n18683 = ~n18676 & n18681;
  assign n18684 = ~n18679 & ~n34716;
  assign n18685 = ~n18389 & ~n18391;
  assign n18686 = ~n18676 & n18685;
  assign n18687 = ~n18399 & ~n18686;
  assign n18688 = ~n18391 & n18399;
  assign n18689 = ~n18389 & n18688;
  assign n18690 = n18399 & n18686;
  assign n18691 = ~n18676 & n18689;
  assign n18692 = ~n18687 & ~n34717;
  assign n18693 = ~n18371 & ~n34675;
  assign n18694 = ~n18676 & n18693;
  assign n18695 = ~n34677 & ~n18694;
  assign n18696 = ~n18371 & n34677;
  assign n18697 = ~n34675 & n18696;
  assign n18698 = n34677 & n18694;
  assign n18699 = ~n18676 & n18697;
  assign n18700 = ~n18695 & ~n34718;
  assign n18701 = ~n18354 & ~n18356;
  assign n18702 = ~n18676 & n18701;
  assign n18703 = ~n34674 & ~n18702;
  assign n18704 = ~n18356 & n34674;
  assign n18705 = ~n18354 & n18704;
  assign n18706 = n34674 & n18702;
  assign n18707 = ~n18676 & n18705;
  assign n18708 = ~n18703 & ~n34719;
  assign n18709 = ~n18323 & ~n18325;
  assign n18710 = ~n18676 & n18709;
  assign n18711 = ~n34670 & ~n18710;
  assign n18712 = ~n18325 & n34670;
  assign n18713 = ~n18323 & n18712;
  assign n18714 = n34670 & n18710;
  assign n18715 = ~n18676 & n18713;
  assign n18716 = ~n18711 & ~n34720;
  assign n18717 = ~n18305 & ~n34666;
  assign n18718 = ~n18676 & n18717;
  assign n18719 = ~n34668 & ~n18718;
  assign n18720 = ~n18305 & n34668;
  assign n18721 = ~n34666 & n18720;
  assign n18722 = n34668 & n18718;
  assign n18723 = ~n18676 & n18721;
  assign n18724 = ~n18719 & ~n34721;
  assign n18725 = ~n18288 & ~n18290;
  assign n18726 = ~n18676 & n18725;
  assign n18727 = ~n34665 & ~n18726;
  assign n18728 = ~n18290 & n34665;
  assign n18729 = ~n18288 & n18728;
  assign n18730 = n34665 & n18726;
  assign n18731 = ~n18676 & n18729;
  assign n18732 = ~n18727 & ~n34722;
  assign n18733 = ~n18257 & ~n18259;
  assign n18734 = ~n18676 & n18733;
  assign n18735 = ~n34661 & ~n18734;
  assign n18736 = ~n18259 & n34661;
  assign n18737 = ~n18257 & n18736;
  assign n18738 = n34661 & n18734;
  assign n18739 = ~n18676 & n18737;
  assign n18740 = ~n18735 & ~n34723;
  assign n18741 = ~n18238 & ~n34656;
  assign n18742 = ~n18676 & n18741;
  assign n18743 = ~n34659 & ~n18742;
  assign n18744 = ~n18238 & n34659;
  assign n18745 = ~n34656 & n18744;
  assign n18746 = n34659 & n18742;
  assign n18747 = ~n18676 & n18745;
  assign n18748 = ~n18743 & ~n34724;
  assign n18749 = ~n18221 & ~n18223;
  assign n18750 = ~n18676 & n18749;
  assign n18751 = ~n34655 & ~n18750;
  assign n18752 = ~n18223 & n34655;
  assign n18753 = ~n18221 & n18752;
  assign n18754 = n34655 & n18750;
  assign n18755 = ~n18676 & n18753;
  assign n18756 = ~n18751 & ~n34725;
  assign n18757 = ~n18187 & ~n18189;
  assign n18758 = ~n18676 & n18757;
  assign n18759 = ~n34650 & ~n18758;
  assign n18760 = ~n18189 & n34650;
  assign n18761 = ~n18187 & n18760;
  assign n18762 = n34650 & n18758;
  assign n18763 = ~n18676 & n18761;
  assign n18764 = ~n18759 & ~n34726;
  assign n18765 = ~n18151 & ~n18153;
  assign n18766 = ~n18676 & n18765;
  assign n18767 = ~n34644 & ~n18766;
  assign n18768 = ~n18153 & n34644;
  assign n18769 = ~n18151 & n18768;
  assign n18770 = n34644 & n18766;
  assign n18771 = ~n18676 & n18769;
  assign n18772 = ~n18767 & ~n34727;
  assign n18773 = ~n18120 & ~n18122;
  assign n18774 = ~n18676 & n18773;
  assign n18775 = ~n34640 & ~n18774;
  assign n18776 = ~n18122 & n34640;
  assign n18777 = ~n18120 & n18776;
  assign n18778 = n34640 & n18774;
  assign n18779 = ~n18676 & n18777;
  assign n18780 = ~n18775 & ~n34728;
  assign n18781 = ~n18084 & ~n18086;
  assign n18782 = ~n18676 & n18781;
  assign n18783 = ~n34634 & ~n18782;
  assign n18784 = ~n18086 & n34634;
  assign n18785 = ~n18084 & n18784;
  assign n18786 = n34634 & n18782;
  assign n18787 = ~n18676 & n18785;
  assign n18788 = ~n18783 & ~n34729;
  assign n18789 = ~n18050 & ~n18052;
  assign n18790 = ~n18676 & n18789;
  assign n18791 = ~n34629 & ~n18790;
  assign n18792 = ~n18052 & n34629;
  assign n18793 = ~n18050 & n18792;
  assign n18794 = n34629 & n18790;
  assign n18795 = ~n18676 & n18793;
  assign n18796 = ~n18791 & ~n34730;
  assign n18797 = ~n18016 & ~n18018;
  assign n18798 = ~n18676 & n18797;
  assign n18799 = ~n34624 & ~n18798;
  assign n18800 = ~n18018 & n34624;
  assign n18801 = ~n18016 & n18800;
  assign n18802 = n34624 & n18798;
  assign n18803 = ~n18676 & n18801;
  assign n18804 = ~n18799 & ~n34731;
  assign n18805 = ~n17983 & ~n17985;
  assign n18806 = ~n18676 & n18805;
  assign n18807 = ~n34620 & ~n18806;
  assign n18808 = ~n17985 & n34620;
  assign n18809 = ~n17983 & n18808;
  assign n18810 = n34620 & n18806;
  assign n18811 = ~n18676 & n18809;
  assign n18812 = ~n18807 & ~n34732;
  assign n18813 = ~n17949 & ~n17951;
  assign n18814 = ~n18676 & n18813;
  assign n18815 = ~n34615 & ~n18814;
  assign n18816 = ~n17951 & n34615;
  assign n18817 = ~n17949 & n18816;
  assign n18818 = n34615 & n18814;
  assign n18819 = ~n18676 & n18817;
  assign n18820 = ~n18815 & ~n34733;
  assign n18821 = ~n17922 & ~n17924;
  assign n18822 = ~n18676 & n18821;
  assign n18823 = ~n17933 & ~n18822;
  assign n18824 = ~n17924 & n17933;
  assign n18825 = ~n17922 & n18824;
  assign n18826 = n17933 & n18822;
  assign n18827 = ~n18676 & n18825;
  assign n18828 = ~n18823 & ~n34734;
  assign n18829 = ~pi30  & ~n18676;
  assign n18830 = ~pi31  & n18829;
  assign n18831 = n17899 & ~n18676;
  assign n18832 = ~n17885 & ~n18674;
  assign n18833 = ~n34715 & n18832;
  assign n18834 = ~n18668 & n18833;
  assign n18835 = ~n34735 & ~n18834;
  assign n18836 = pi32  & ~n18835;
  assign n18837 = ~pi32  & ~n18834;
  assign n18838 = ~pi32  & n18835;
  assign n18839 = ~n34735 & n18837;
  assign n18840 = ~n18836 & ~n34736;
  assign n18841 = pi30  & ~n18676;
  assign n18842 = ~pi28  & ~pi29 ;
  assign n18843 = ~pi30  & n18842;
  assign n18844 = ~n17168 & ~n34609;
  assign n18845 = ~n17169 & n18844;
  assign n18846 = ~n17185 & n18845;
  assign n18847 = ~n34516 & n18846;
  assign n18848 = n34514 & n17187;
  assign n18849 = ~n17179 & n18847;
  assign n18850 = ~n18843 & ~n34737;
  assign n18851 = ~n17883 & n18850;
  assign n18852 = ~n34605 & n18851;
  assign n18853 = ~n17877 & n18852;
  assign n18854 = ~n18841 & ~n18843;
  assign n18855 = n17885 & n18854;
  assign n18856 = ~n18841 & n18853;
  assign n18857 = pi31  & ~n18829;
  assign n18858 = ~n34735 & ~n18857;
  assign n18859 = ~n34738 & n18858;
  assign n18860 = ~n17885 & ~n18854;
  assign n18861 = n17187 & ~n18860;
  assign n18862 = ~n18859 & ~n18860;
  assign n18863 = n17187 & n18862;
  assign n18864 = ~n18859 & n18861;
  assign n18865 = ~n18840 & ~n34739;
  assign n18866 = ~n17187 & ~n18862;
  assign n18867 = n16428 & ~n18866;
  assign n18868 = ~n18865 & n18867;
  assign n18869 = ~n17902 & ~n34610;
  assign n18870 = ~n18676 & n18869;
  assign n18871 = n17907 & ~n18870;
  assign n18872 = ~n17907 & n18869;
  assign n18873 = ~n17907 & n18870;
  assign n18874 = ~n18676 & n18872;
  assign n18875 = ~n18871 & ~n34740;
  assign n18876 = ~n18868 & ~n18875;
  assign n18877 = ~n18865 & ~n18866;
  assign n18878 = ~n16428 & ~n18877;
  assign n18879 = n15760 & ~n18878;
  assign n18880 = ~n18876 & ~n18878;
  assign n18881 = n15760 & n18880;
  assign n18882 = ~n18876 & n18879;
  assign n18883 = ~n18828 & ~n34741;
  assign n18884 = ~n15760 & ~n18880;
  assign n18885 = n15033 & ~n18884;
  assign n18886 = ~n18883 & n18885;
  assign n18887 = ~n17936 & ~n34612;
  assign n18888 = ~n18676 & n18887;
  assign n18889 = n17946 & ~n18888;
  assign n18890 = ~n17946 & n18888;
  assign n18891 = ~n17936 & n17946;
  assign n18892 = ~n34612 & n18891;
  assign n18893 = n17946 & n18888;
  assign n18894 = ~n18676 & n18892;
  assign n18895 = ~n17946 & ~n18888;
  assign n18896 = ~n34742 & ~n18895;
  assign n18897 = ~n18889 & ~n18890;
  assign n18898 = ~n18886 & ~n34743;
  assign n18899 = ~n18883 & ~n18884;
  assign n18900 = ~n15033 & ~n18899;
  assign n18901 = n14394 & ~n18900;
  assign n18902 = ~n18898 & ~n18900;
  assign n18903 = n14394 & n18902;
  assign n18904 = ~n18898 & n18901;
  assign n18905 = ~n18820 & ~n34744;
  assign n18906 = ~n14394 & ~n18902;
  assign n18907 = n13704 & ~n18906;
  assign n18908 = ~n18905 & n18907;
  assign n18909 = ~n17966 & ~n34616;
  assign n18910 = ~n18676 & n18909;
  assign n18911 = ~n34618 & n18910;
  assign n18912 = n34618 & ~n18910;
  assign n18913 = ~n17966 & n34618;
  assign n18914 = ~n34616 & n18913;
  assign n18915 = ~n18676 & n18914;
  assign n18916 = ~n34618 & ~n18910;
  assign n18917 = ~n18915 & ~n18916;
  assign n18918 = ~n18911 & ~n18912;
  assign n18919 = ~n18908 & ~n34745;
  assign n18920 = ~n18905 & ~n18906;
  assign n18921 = ~n13704 & ~n18920;
  assign n18922 = n13099 & ~n18921;
  assign n18923 = ~n18919 & ~n18921;
  assign n18924 = n13099 & n18923;
  assign n18925 = ~n18919 & n18922;
  assign n18926 = ~n18812 & ~n34746;
  assign n18927 = ~n13099 & ~n18923;
  assign n18928 = n12442 & ~n18927;
  assign n18929 = ~n18926 & n18928;
  assign n18930 = ~n18000 & ~n34621;
  assign n18931 = ~n18676 & n18930;
  assign n18932 = ~n34622 & ~n18931;
  assign n18933 = ~n18000 & n34622;
  assign n18934 = ~n34621 & n18933;
  assign n18935 = n34622 & n18931;
  assign n18936 = ~n18676 & n18934;
  assign n18937 = n34622 & ~n18931;
  assign n18938 = ~n34622 & n18931;
  assign n18939 = ~n18937 & ~n18938;
  assign n18940 = ~n18932 & ~n34747;
  assign n18941 = ~n18929 & n34748;
  assign n18942 = ~n18926 & ~n18927;
  assign n18943 = ~n12442 & ~n18942;
  assign n18944 = n11858 & ~n18943;
  assign n18945 = ~n18941 & ~n18943;
  assign n18946 = n11858 & n18945;
  assign n18947 = ~n18941 & n18944;
  assign n18948 = ~n18804 & ~n34749;
  assign n18949 = ~n11858 & ~n18945;
  assign n18950 = n11229 & ~n18949;
  assign n18951 = ~n18948 & n18950;
  assign n18952 = ~n18033 & ~n34625;
  assign n18953 = ~n18676 & n18952;
  assign n18954 = n34627 & ~n18953;
  assign n18955 = ~n18033 & ~n34627;
  assign n18956 = ~n34625 & n18955;
  assign n18957 = ~n34627 & n18953;
  assign n18958 = ~n18676 & n18956;
  assign n18959 = n34627 & n18953;
  assign n18960 = ~n34627 & ~n18953;
  assign n18961 = ~n18959 & ~n18960;
  assign n18962 = ~n18954 & ~n34750;
  assign n18963 = ~n18951 & n34751;
  assign n18964 = ~n18948 & ~n18949;
  assign n18965 = ~n11229 & ~n18964;
  assign n18966 = n10681 & ~n18965;
  assign n18967 = ~n18963 & ~n18965;
  assign n18968 = n10681 & n18967;
  assign n18969 = ~n18963 & n18966;
  assign n18970 = ~n18796 & ~n34752;
  assign n18971 = ~n10681 & ~n18967;
  assign n18972 = n10086 & ~n18971;
  assign n18973 = ~n18970 & n18972;
  assign n18974 = ~n18067 & ~n34630;
  assign n18975 = ~n18067 & ~n18676;
  assign n18976 = ~n34630 & n18975;
  assign n18977 = ~n18676 & n18974;
  assign n18978 = ~n34632 & ~n34753;
  assign n18979 = n18082 & n18975;
  assign n18980 = n34632 & n34753;
  assign n18981 = ~n18067 & ~n34632;
  assign n18982 = ~n34630 & n18981;
  assign n18983 = ~n18676 & n18982;
  assign n18984 = n34632 & ~n34753;
  assign n18985 = ~n18983 & ~n18984;
  assign n18986 = ~n18978 & ~n34754;
  assign n18987 = ~n18973 & ~n34755;
  assign n18988 = ~n18970 & ~n18971;
  assign n18989 = ~n10086 & ~n18988;
  assign n18990 = n9565 & ~n18989;
  assign n18991 = ~n18987 & ~n18989;
  assign n18992 = n9565 & n18991;
  assign n18993 = ~n18987 & n18990;
  assign n18994 = ~n18788 & ~n34756;
  assign n18995 = ~n9565 & ~n18991;
  assign n18996 = n8998 & ~n18995;
  assign n18997 = ~n18994 & n18996;
  assign n18998 = ~n18101 & ~n34635;
  assign n18999 = ~n18676 & n18998;
  assign n19000 = ~n34638 & ~n18999;
  assign n19001 = ~n18101 & n34638;
  assign n19002 = ~n34635 & n19001;
  assign n19003 = n34638 & n18999;
  assign n19004 = ~n18676 & n19002;
  assign n19005 = ~n19000 & ~n34757;
  assign n19006 = ~n18997 & ~n19005;
  assign n19007 = ~n18994 & ~n18995;
  assign n19008 = ~n8998 & ~n19007;
  assign n19009 = n8506 & ~n19008;
  assign n19010 = ~n19006 & ~n19008;
  assign n19011 = n8506 & n19010;
  assign n19012 = ~n19006 & n19009;
  assign n19013 = ~n18780 & ~n34758;
  assign n19014 = ~n8506 & ~n19010;
  assign n19015 = n7975 & ~n19014;
  assign n19016 = ~n19013 & n19015;
  assign n19017 = ~n18137 & ~n34641;
  assign n19018 = ~n18137 & ~n18676;
  assign n19019 = ~n34641 & n19018;
  assign n19020 = ~n18676 & n19017;
  assign n19021 = n18148 & ~n34759;
  assign n19022 = n18149 & n19018;
  assign n19023 = ~n18148 & n34759;
  assign n19024 = ~n18137 & n18148;
  assign n19025 = ~n34641 & n19024;
  assign n19026 = ~n18676 & n19025;
  assign n19027 = ~n18148 & ~n34759;
  assign n19028 = ~n19026 & ~n19027;
  assign n19029 = ~n19021 & ~n34760;
  assign n19030 = ~n19016 & ~n34761;
  assign n19031 = ~n19013 & ~n19014;
  assign n19032 = ~n7975 & ~n19031;
  assign n19033 = n7512 & ~n19032;
  assign n19034 = ~n19030 & ~n19032;
  assign n19035 = n7512 & n19034;
  assign n19036 = ~n19030 & n19033;
  assign n19037 = ~n18772 & ~n34762;
  assign n19038 = ~n7512 & ~n19034;
  assign n19039 = n7015 & ~n19038;
  assign n19040 = ~n19037 & n19039;
  assign n19041 = ~n18168 & ~n34645;
  assign n19042 = ~n18676 & n19041;
  assign n19043 = ~n34648 & n19042;
  assign n19044 = n34648 & ~n19042;
  assign n19045 = ~n18168 & n34648;
  assign n19046 = ~n34645 & n19045;
  assign n19047 = n34648 & n19042;
  assign n19048 = ~n18676 & n19046;
  assign n19049 = ~n34648 & ~n19042;
  assign n19050 = ~n34763 & ~n19049;
  assign n19051 = ~n19043 & ~n19044;
  assign n19052 = ~n19040 & ~n34764;
  assign n19053 = ~n19037 & ~n19038;
  assign n19054 = ~n7015 & ~n19053;
  assign n19055 = n6579 & ~n19054;
  assign n19056 = ~n19052 & ~n19054;
  assign n19057 = n6579 & n19056;
  assign n19058 = ~n19052 & n19055;
  assign n19059 = ~n18764 & ~n34765;
  assign n19060 = ~n6579 & ~n19056;
  assign n19061 = n6117 & ~n19060;
  assign n19062 = ~n19059 & n19061;
  assign n19063 = ~n18204 & ~n34651;
  assign n19064 = ~n18204 & ~n18676;
  assign n19065 = ~n34651 & n19064;
  assign n19066 = ~n18676 & n19063;
  assign n19067 = n34653 & ~n34766;
  assign n19068 = n18219 & n19064;
  assign n19069 = ~n34653 & n34766;
  assign n19070 = ~n18204 & n34653;
  assign n19071 = ~n34651 & n19070;
  assign n19072 = ~n18676 & n19071;
  assign n19073 = ~n34653 & ~n34766;
  assign n19074 = ~n19072 & ~n19073;
  assign n19075 = ~n19067 & ~n34767;
  assign n19076 = ~n19062 & ~n34768;
  assign n19077 = ~n19059 & ~n19060;
  assign n19078 = ~n6117 & ~n19077;
  assign n19079 = n5708 & ~n19078;
  assign n19080 = ~n19076 & ~n19078;
  assign n19081 = n5708 & n19080;
  assign n19082 = ~n19076 & n19079;
  assign n19083 = ~n18756 & ~n34769;
  assign n19084 = ~n5708 & ~n19080;
  assign n19085 = n5278 & ~n19084;
  assign n19086 = ~n19083 & n19085;
  assign n19087 = ~n18748 & ~n19086;
  assign n19088 = ~n19083 & ~n19084;
  assign n19089 = ~n5278 & ~n19088;
  assign n19090 = n4903 & ~n19089;
  assign n19091 = ~n19087 & ~n19089;
  assign n19092 = n4903 & n19091;
  assign n19093 = ~n19087 & n19090;
  assign n19094 = ~n18740 & ~n34770;
  assign n19095 = ~n4903 & ~n19091;
  assign n19096 = n4508 & ~n19095;
  assign n19097 = ~n19094 & n19096;
  assign n19098 = ~n18274 & ~n34663;
  assign n19099 = ~n18274 & ~n18676;
  assign n19100 = ~n34663 & n19099;
  assign n19101 = ~n18676 & n19098;
  assign n19102 = n18282 & ~n34771;
  assign n19103 = n18286 & n19099;
  assign n19104 = ~n18274 & n18282;
  assign n19105 = ~n34663 & n19104;
  assign n19106 = ~n18676 & n19105;
  assign n19107 = ~n18282 & ~n34771;
  assign n19108 = ~n19106 & ~n19107;
  assign n19109 = ~n19102 & ~n19103;
  assign n19110 = ~n19097 & ~n34772;
  assign n19111 = ~n19094 & ~n19095;
  assign n19112 = ~n4508 & ~n19111;
  assign n19113 = n4155 & ~n19112;
  assign n19114 = ~n19110 & ~n19112;
  assign n19115 = n4155 & n19114;
  assign n19116 = ~n19110 & n19113;
  assign n19117 = ~n18732 & ~n34773;
  assign n19118 = ~n4155 & ~n19114;
  assign n19119 = n3788 & ~n19118;
  assign n19120 = ~n19117 & n19119;
  assign n19121 = ~n18724 & ~n19120;
  assign n19122 = ~n19117 & ~n19118;
  assign n19123 = ~n3788 & ~n19122;
  assign n19124 = n3473 & ~n19123;
  assign n19125 = ~n19121 & ~n19123;
  assign n19126 = n3473 & n19125;
  assign n19127 = ~n19121 & n19124;
  assign n19128 = ~n18716 & ~n34774;
  assign n19129 = ~n3473 & ~n19125;
  assign n19130 = n3140 & ~n19129;
  assign n19131 = ~n19128 & n19130;
  assign n19132 = ~n18340 & ~n34672;
  assign n19133 = ~n18340 & ~n18676;
  assign n19134 = ~n34672 & n19133;
  assign n19135 = ~n18676 & n19132;
  assign n19136 = n18348 & ~n34775;
  assign n19137 = n18352 & n19133;
  assign n19138 = ~n18340 & n18348;
  assign n19139 = ~n34672 & n19138;
  assign n19140 = ~n18676 & n19139;
  assign n19141 = ~n18348 & ~n34775;
  assign n19142 = ~n19140 & ~n19141;
  assign n19143 = ~n19136 & ~n19137;
  assign n19144 = ~n19131 & ~n34776;
  assign n19145 = ~n19128 & ~n19129;
  assign n19146 = ~n3140 & ~n19145;
  assign n19147 = n2855 & ~n19146;
  assign n19148 = ~n19144 & ~n19146;
  assign n19149 = n2855 & n19148;
  assign n19150 = ~n19144 & n19147;
  assign n19151 = ~n18708 & ~n34777;
  assign n19152 = ~n2855 & ~n19148;
  assign n19153 = n2556 & ~n19152;
  assign n19154 = ~n19151 & n19153;
  assign n19155 = ~n18700 & ~n19154;
  assign n19156 = ~n19151 & ~n19152;
  assign n19157 = ~n2556 & ~n19156;
  assign n19158 = n2301 & ~n19157;
  assign n19159 = ~n19155 & ~n19157;
  assign n19160 = n2301 & n19159;
  assign n19161 = ~n19155 & n19158;
  assign n19162 = ~n18692 & ~n34778;
  assign n19163 = ~n2301 & ~n19159;
  assign n19164 = ~n19162 & ~n19163;
  assign n19165 = ~n2038 & ~n19164;
  assign n19166 = n2038 & ~n19163;
  assign n19167 = ~n19162 & n19166;
  assign n19168 = ~n18402 & ~n34679;
  assign n19169 = ~n18676 & n19168;
  assign n19170 = ~n34681 & ~n19169;
  assign n19171 = ~n18402 & n34681;
  assign n19172 = ~n34679 & n19171;
  assign n19173 = n34681 & n19169;
  assign n19174 = ~n18676 & n19172;
  assign n19175 = n34681 & ~n19169;
  assign n19176 = ~n34681 & n19169;
  assign n19177 = ~n19175 & ~n19176;
  assign n19178 = ~n19170 & ~n34779;
  assign n19179 = ~n19167 & n34780;
  assign n19180 = ~n19165 & ~n19179;
  assign n19181 = ~n1812 & ~n19180;
  assign n19182 = n1812 & ~n19165;
  assign n19183 = n1812 & n19180;
  assign n19184 = ~n19179 & n19182;
  assign n19185 = ~n18684 & ~n34781;
  assign n19186 = ~n19181 & ~n19185;
  assign n19187 = ~n1582 & ~n19186;
  assign n19188 = n1582 & ~n19181;
  assign n19189 = ~n19185 & n19188;
  assign n19190 = ~n18424 & ~n34683;
  assign n19191 = ~n18424 & ~n18676;
  assign n19192 = ~n34683 & n19191;
  assign n19193 = ~n18676 & n19190;
  assign n19194 = n18432 & ~n34782;
  assign n19195 = n18436 & n19191;
  assign n19196 = ~n18424 & n18432;
  assign n19197 = ~n34683 & n19196;
  assign n19198 = ~n18676 & n19197;
  assign n19199 = ~n18432 & ~n34782;
  assign n19200 = ~n19198 & ~n19199;
  assign n19201 = ~n19194 & ~n19195;
  assign n19202 = ~n19189 & ~n34783;
  assign n19203 = ~n19187 & ~n19202;
  assign n19204 = ~n1388 & ~n19203;
  assign n19205 = ~n18438 & ~n18440;
  assign n19206 = ~n18676 & n19205;
  assign n19207 = ~n34685 & ~n19206;
  assign n19208 = ~n18440 & n34685;
  assign n19209 = ~n18438 & n19208;
  assign n19210 = n34685 & n19206;
  assign n19211 = ~n18676 & n19209;
  assign n19212 = ~n19207 & ~n34784;
  assign n19213 = n1388 & ~n19187;
  assign n19214 = n1388 & n19203;
  assign n19215 = ~n19202 & n19213;
  assign n19216 = ~n19212 & ~n34785;
  assign n19217 = ~n19204 & ~n19216;
  assign n19218 = ~n1192 & ~n19217;
  assign n19219 = n1192 & ~n19204;
  assign n19220 = ~n19216 & n19219;
  assign n19221 = ~n18455 & ~n34687;
  assign n19222 = ~n18455 & ~n18676;
  assign n19223 = ~n34687 & n19222;
  assign n19224 = ~n18676 & n19221;
  assign n19225 = n18463 & ~n34786;
  assign n19226 = n18467 & n19222;
  assign n19227 = ~n18455 & n18463;
  assign n19228 = ~n34687 & n19227;
  assign n19229 = ~n18676 & n19228;
  assign n19230 = ~n18463 & ~n34786;
  assign n19231 = ~n19229 & ~n19230;
  assign n19232 = ~n19225 & ~n19226;
  assign n19233 = ~n19220 & ~n34787;
  assign n19234 = ~n19218 & ~n19233;
  assign n19235 = ~n1028 & ~n19234;
  assign n19236 = ~n18469 & ~n18471;
  assign n19237 = ~n18676 & n19236;
  assign n19238 = ~n34689 & ~n19237;
  assign n19239 = ~n18471 & n34689;
  assign n19240 = ~n18469 & n19239;
  assign n19241 = n34689 & n19237;
  assign n19242 = ~n18676 & n19240;
  assign n19243 = ~n19238 & ~n34788;
  assign n19244 = n1028 & ~n19218;
  assign n19245 = n1028 & n19234;
  assign n19246 = ~n19233 & n19244;
  assign n19247 = ~n19243 & ~n34789;
  assign n19248 = ~n19235 & ~n19247;
  assign n19249 = ~n866 & ~n19248;
  assign n19250 = ~n18486 & ~n34690;
  assign n19251 = ~n18676 & n19250;
  assign n19252 = ~n34692 & ~n19251;
  assign n19253 = ~n18486 & n34692;
  assign n19254 = ~n34690 & n19253;
  assign n19255 = n34692 & n19251;
  assign n19256 = ~n18676 & n19254;
  assign n19257 = ~n19252 & ~n34790;
  assign n19258 = n866 & ~n19235;
  assign n19259 = ~n19247 & n19258;
  assign n19260 = ~n19257 & ~n19259;
  assign n19261 = ~n19249 & ~n19260;
  assign n19262 = ~n730 & ~n19261;
  assign n19263 = ~n18504 & ~n18506;
  assign n19264 = ~n18676 & n19263;
  assign n19265 = ~n34694 & ~n19264;
  assign n19266 = ~n18506 & n34694;
  assign n19267 = ~n18504 & n19266;
  assign n19268 = n34694 & n19264;
  assign n19269 = ~n18676 & n19267;
  assign n19270 = ~n19265 & ~n34791;
  assign n19271 = n730 & ~n19249;
  assign n19272 = n730 & n19261;
  assign n19273 = ~n19260 & n19271;
  assign n19274 = ~n19270 & ~n34792;
  assign n19275 = ~n19262 & ~n19274;
  assign n19276 = ~n602 & ~n19275;
  assign n19277 = n602 & ~n19262;
  assign n19278 = ~n19274 & n19277;
  assign n19279 = ~n18521 & ~n34696;
  assign n19280 = ~n18521 & ~n18676;
  assign n19281 = ~n34696 & n19280;
  assign n19282 = ~n18676 & n19279;
  assign n19283 = n18529 & ~n34793;
  assign n19284 = n18533 & n19280;
  assign n19285 = ~n18521 & n18529;
  assign n19286 = ~n34696 & n19285;
  assign n19287 = ~n18676 & n19286;
  assign n19288 = ~n18529 & ~n34793;
  assign n19289 = ~n19287 & ~n19288;
  assign n19290 = ~n19283 & ~n19284;
  assign n19291 = ~n19278 & ~n34794;
  assign n19292 = ~n19276 & ~n19291;
  assign n19293 = ~n497 & ~n19292;
  assign n19294 = ~n18535 & ~n18537;
  assign n19295 = ~n18676 & n19294;
  assign n19296 = ~n34698 & ~n19295;
  assign n19297 = ~n18537 & n34698;
  assign n19298 = ~n18535 & n19297;
  assign n19299 = n34698 & n19295;
  assign n19300 = ~n18676 & n19298;
  assign n19301 = ~n19296 & ~n34795;
  assign n19302 = n497 & ~n19276;
  assign n19303 = n497 & n19292;
  assign n19304 = ~n19291 & n19302;
  assign n19305 = ~n19301 & ~n34796;
  assign n19306 = ~n19293 & ~n19305;
  assign n19307 = ~n403 & ~n19306;
  assign n19308 = ~n18552 & ~n34699;
  assign n19309 = ~n18676 & n19308;
  assign n19310 = ~n34701 & ~n19309;
  assign n19311 = ~n18552 & n34701;
  assign n19312 = ~n34699 & n19311;
  assign n19313 = n34701 & n19309;
  assign n19314 = ~n18676 & n19312;
  assign n19315 = ~n19310 & ~n34797;
  assign n19316 = n403 & ~n19293;
  assign n19317 = ~n19305 & n19316;
  assign n19318 = ~n19315 & ~n19317;
  assign n19319 = ~n19307 & ~n19318;
  assign n19320 = ~n330 & ~n19319;
  assign n19321 = ~n18570 & ~n18572;
  assign n19322 = ~n18676 & n19321;
  assign n19323 = ~n34703 & ~n19322;
  assign n19324 = ~n18572 & n34703;
  assign n19325 = ~n18570 & n19324;
  assign n19326 = n34703 & n19322;
  assign n19327 = ~n18676 & n19325;
  assign n19328 = ~n19323 & ~n34798;
  assign n19329 = n330 & ~n19307;
  assign n19330 = n330 & n19319;
  assign n19331 = ~n19318 & n19329;
  assign n19332 = ~n19328 & ~n34799;
  assign n19333 = ~n19320 & ~n19332;
  assign n19334 = ~n271 & ~n19333;
  assign n19335 = n271 & ~n19320;
  assign n19336 = ~n19332 & n19335;
  assign n19337 = ~n18587 & ~n34705;
  assign n19338 = ~n18587 & ~n18676;
  assign n19339 = ~n34705 & n19338;
  assign n19340 = ~n18676 & n19337;
  assign n19341 = n18595 & ~n34800;
  assign n19342 = n18599 & n19338;
  assign n19343 = ~n18587 & n18595;
  assign n19344 = ~n34705 & n19343;
  assign n19345 = ~n18676 & n19344;
  assign n19346 = ~n18595 & ~n34800;
  assign n19347 = ~n19345 & ~n19346;
  assign n19348 = ~n19341 & ~n19342;
  assign n19349 = ~n19336 & ~n34801;
  assign n19350 = ~n19334 & ~n19349;
  assign n19351 = ~n217 & ~n19350;
  assign n19352 = ~n18601 & ~n18603;
  assign n19353 = ~n18676 & n19352;
  assign n19354 = ~n34707 & ~n19353;
  assign n19355 = ~n18603 & n34707;
  assign n19356 = ~n18601 & n19355;
  assign n19357 = n34707 & n19353;
  assign n19358 = ~n18676 & n19356;
  assign n19359 = ~n19354 & ~n34802;
  assign n19360 = n217 & ~n19334;
  assign n19361 = n217 & n19350;
  assign n19362 = ~n19349 & n19360;
  assign n19363 = ~n19359 & ~n34803;
  assign n19364 = ~n19351 & ~n19363;
  assign n19365 = ~n198 & ~n19364;
  assign n19366 = ~n18618 & ~n34708;
  assign n19367 = ~n18676 & n19366;
  assign n19368 = ~n34710 & ~n19367;
  assign n19369 = ~n18618 & n34710;
  assign n19370 = ~n34708 & n19369;
  assign n19371 = n34710 & n19367;
  assign n19372 = ~n18676 & n19370;
  assign n19373 = ~n19368 & ~n34804;
  assign n19374 = n198 & ~n19351;
  assign n19375 = ~n19363 & n19374;
  assign n19376 = ~n19373 & ~n19375;
  assign n19377 = ~n19365 & ~n19376;
  assign n19378 = ~n18636 & ~n18638;
  assign n19379 = ~n18676 & n19378;
  assign n19380 = ~n34712 & ~n19379;
  assign n19381 = ~n18638 & n34712;
  assign n19382 = ~n18636 & n19381;
  assign n19383 = n34712 & n19379;
  assign n19384 = ~n18676 & n19382;
  assign n19385 = ~n19380 & ~n34805;
  assign n19386 = ~n18652 & ~n18660;
  assign n19387 = ~n18660 & ~n18676;
  assign n19388 = ~n18652 & n19387;
  assign n19389 = ~n18676 & n19386;
  assign n19390 = ~n34715 & ~n34806;
  assign n19391 = ~n19385 & n19390;
  assign n19392 = ~n19377 & n19391;
  assign n19393 = n193 & ~n19392;
  assign n19394 = ~n19365 & n19385;
  assign n19395 = n19377 & n19385;
  assign n19396 = ~n19376 & n19394;
  assign n19397 = n18652 & ~n19387;
  assign n19398 = ~n193 & ~n19386;
  assign n19399 = ~n19397 & n19398;
  assign n19400 = ~n34807 & ~n19399;
  assign n19401 = ~n19393 & n19400;
  assign n19402 = ~n19181 & ~n34781;
  assign n19403 = ~n19181 & ~n19401;
  assign n19404 = ~n34781 & n19403;
  assign n19405 = ~n19401 & n19402;
  assign n19406 = n18684 & ~n34808;
  assign n19407 = n19185 & n19403;
  assign n19408 = n18684 & ~n34781;
  assign n19409 = ~n19181 & n19408;
  assign n19410 = ~n19401 & n19409;
  assign n19411 = ~n18684 & ~n34808;
  assign n19412 = ~n19410 & ~n19411;
  assign n19413 = ~n19406 & ~n19407;
  assign n19414 = pi28  & ~n19401;
  assign n19415 = ~pi26  & ~pi27 ;
  assign n19416 = ~pi28  & n19415;
  assign n19417 = ~n19414 & ~n19416;
  assign n19418 = ~n18676 & ~n19417;
  assign n19419 = ~pi28  & ~n19401;
  assign n19420 = pi29  & ~n19419;
  assign n19421 = ~pi29  & n19419;
  assign n19422 = n18842 & ~n19401;
  assign n19423 = ~n19420 & ~n34810;
  assign n19424 = ~n34603 & ~n34737;
  assign n19425 = ~n17864 & n19424;
  assign n19426 = ~n17883 & n19425;
  assign n19427 = ~n34605 & n19426;
  assign n19428 = n17869 & n17885;
  assign n19429 = ~n17877 & n19427;
  assign n19430 = ~n19416 & ~n34811;
  assign n19431 = ~n18674 & n19430;
  assign n19432 = ~n34715 & n19431;
  assign n19433 = ~n18668 & n19432;
  assign n19434 = n18676 & n19417;
  assign n19435 = ~n19414 & n19433;
  assign n19436 = n19423 & ~n34812;
  assign n19437 = ~n19418 & ~n19436;
  assign n19438 = ~n17885 & ~n19437;
  assign n19439 = n17885 & ~n19418;
  assign n19440 = ~n19436 & n19439;
  assign n19441 = ~n18676 & ~n19399;
  assign n19442 = ~n34807 & n19441;
  assign n19443 = ~n19393 & n19442;
  assign n19444 = ~n34810 & ~n19443;
  assign n19445 = pi30  & ~n19444;
  assign n19446 = ~pi30  & ~n19443;
  assign n19447 = ~pi30  & n19444;
  assign n19448 = ~n34810 & n19446;
  assign n19449 = ~n19445 & ~n34813;
  assign n19450 = ~n19440 & ~n19449;
  assign n19451 = ~n19438 & ~n19450;
  assign n19452 = ~n17187 & ~n19451;
  assign n19453 = n17187 & ~n19438;
  assign n19454 = ~n19450 & n19453;
  assign n19455 = n17187 & n19451;
  assign n19456 = ~n34738 & ~n18860;
  assign n19457 = ~n19401 & n19456;
  assign n19458 = n18858 & ~n19457;
  assign n19459 = ~n18858 & n19456;
  assign n19460 = ~n18858 & n19457;
  assign n19461 = ~n19401 & n19459;
  assign n19462 = ~n19458 & ~n34815;
  assign n19463 = ~n34814 & ~n19462;
  assign n19464 = ~n19452 & ~n19463;
  assign n19465 = ~n16428 & ~n19464;
  assign n19466 = n16428 & ~n19452;
  assign n19467 = ~n19463 & n19466;
  assign n19468 = ~n34739 & ~n18866;
  assign n19469 = ~n18866 & ~n19401;
  assign n19470 = ~n34739 & n19469;
  assign n19471 = ~n19401 & n19468;
  assign n19472 = n18840 & ~n34816;
  assign n19473 = n18865 & n19469;
  assign n19474 = n18840 & ~n34739;
  assign n19475 = ~n18866 & n19474;
  assign n19476 = ~n19401 & n19475;
  assign n19477 = ~n18840 & ~n34816;
  assign n19478 = ~n19476 & ~n19477;
  assign n19479 = ~n19472 & ~n19473;
  assign n19480 = ~n19467 & ~n34817;
  assign n19481 = ~n19465 & ~n19480;
  assign n19482 = ~n15760 & ~n19481;
  assign n19483 = n15760 & ~n19465;
  assign n19484 = ~n19480 & n19483;
  assign n19485 = n15760 & n19481;
  assign n19486 = ~n18868 & ~n18878;
  assign n19487 = ~n19401 & n19486;
  assign n19488 = n18875 & ~n19487;
  assign n19489 = ~n18875 & n19487;
  assign n19490 = n18875 & ~n18878;
  assign n19491 = ~n18868 & n19490;
  assign n19492 = n18875 & n19487;
  assign n19493 = ~n19401 & n19491;
  assign n19494 = ~n18875 & ~n19487;
  assign n19495 = ~n34819 & ~n19494;
  assign n19496 = ~n19488 & ~n19489;
  assign n19497 = ~n34818 & ~n34820;
  assign n19498 = ~n19482 & ~n19497;
  assign n19499 = ~n15033 & ~n19498;
  assign n19500 = n15033 & ~n19482;
  assign n19501 = ~n19497 & n19500;
  assign n19502 = ~n34741 & ~n18884;
  assign n19503 = ~n18884 & ~n19401;
  assign n19504 = ~n34741 & n19503;
  assign n19505 = ~n19401 & n19502;
  assign n19506 = n18828 & ~n34821;
  assign n19507 = n18883 & n19503;
  assign n19508 = n18828 & ~n34741;
  assign n19509 = ~n18884 & n19508;
  assign n19510 = ~n19401 & n19509;
  assign n19511 = ~n18828 & ~n34821;
  assign n19512 = ~n19510 & ~n19511;
  assign n19513 = ~n19506 & ~n19507;
  assign n19514 = ~n19501 & ~n34822;
  assign n19515 = ~n19499 & ~n19514;
  assign n19516 = ~n14394 & ~n19515;
  assign n19517 = n14394 & ~n19499;
  assign n19518 = ~n19514 & n19517;
  assign n19519 = n14394 & n19515;
  assign n19520 = ~n18886 & ~n18900;
  assign n19521 = ~n19401 & n19520;
  assign n19522 = ~n34743 & n19521;
  assign n19523 = n34743 & ~n19521;
  assign n19524 = n34743 & ~n18900;
  assign n19525 = ~n18886 & n19524;
  assign n19526 = ~n19401 & n19525;
  assign n19527 = ~n34743 & ~n19521;
  assign n19528 = ~n19526 & ~n19527;
  assign n19529 = ~n19522 & ~n19523;
  assign n19530 = ~n34823 & ~n34824;
  assign n19531 = ~n19516 & ~n19530;
  assign n19532 = ~n13704 & ~n19531;
  assign n19533 = n13704 & ~n19516;
  assign n19534 = ~n19530 & n19533;
  assign n19535 = ~n34744 & ~n18906;
  assign n19536 = ~n18906 & ~n19401;
  assign n19537 = ~n34744 & n19536;
  assign n19538 = ~n19401 & n19535;
  assign n19539 = n18820 & ~n34825;
  assign n19540 = n18905 & n19536;
  assign n19541 = n18820 & ~n34744;
  assign n19542 = ~n18906 & n19541;
  assign n19543 = ~n19401 & n19542;
  assign n19544 = ~n18820 & ~n34825;
  assign n19545 = ~n19543 & ~n19544;
  assign n19546 = ~n19539 & ~n19540;
  assign n19547 = ~n19534 & ~n34826;
  assign n19548 = ~n19532 & ~n19547;
  assign n19549 = ~n13099 & ~n19548;
  assign n19550 = n13099 & ~n19532;
  assign n19551 = ~n19547 & n19550;
  assign n19552 = n13099 & n19548;
  assign n19553 = ~n18908 & ~n18921;
  assign n19554 = ~n19401 & n19553;
  assign n19555 = ~n34745 & ~n19554;
  assign n19556 = n34745 & ~n18921;
  assign n19557 = ~n18908 & n19556;
  assign n19558 = n34745 & n19554;
  assign n19559 = ~n19401 & n19557;
  assign n19560 = n34745 & ~n19554;
  assign n19561 = ~n34745 & n19554;
  assign n19562 = ~n19560 & ~n19561;
  assign n19563 = ~n19555 & ~n34828;
  assign n19564 = ~n34827 & n34829;
  assign n19565 = ~n19549 & ~n19564;
  assign n19566 = ~n12442 & ~n19565;
  assign n19567 = n12442 & ~n19549;
  assign n19568 = ~n19564 & n19567;
  assign n19569 = ~n34746 & ~n18927;
  assign n19570 = ~n18927 & ~n19401;
  assign n19571 = ~n34746 & n19570;
  assign n19572 = ~n19401 & n19569;
  assign n19573 = n18812 & ~n34830;
  assign n19574 = n18926 & n19570;
  assign n19575 = n18812 & ~n34746;
  assign n19576 = ~n18927 & n19575;
  assign n19577 = ~n19401 & n19576;
  assign n19578 = ~n18812 & ~n34830;
  assign n19579 = ~n19577 & ~n19578;
  assign n19580 = ~n19573 & ~n19574;
  assign n19581 = ~n19568 & ~n34831;
  assign n19582 = ~n19566 & ~n19581;
  assign n19583 = ~n11858 & ~n19582;
  assign n19584 = n11858 & ~n19566;
  assign n19585 = ~n19581 & n19584;
  assign n19586 = n11858 & n19582;
  assign n19587 = ~n18929 & ~n18943;
  assign n19588 = ~n19401 & n19587;
  assign n19589 = n34748 & ~n19588;
  assign n19590 = ~n34748 & ~n18943;
  assign n19591 = ~n18929 & n19590;
  assign n19592 = ~n34748 & n19588;
  assign n19593 = ~n19401 & n19591;
  assign n19594 = n34748 & n19588;
  assign n19595 = ~n34748 & ~n19588;
  assign n19596 = ~n19594 & ~n19595;
  assign n19597 = ~n19589 & ~n34833;
  assign n19598 = ~n34832 & n34834;
  assign n19599 = ~n19583 & ~n19598;
  assign n19600 = ~n11229 & ~n19599;
  assign n19601 = n11229 & ~n19583;
  assign n19602 = ~n19598 & n19601;
  assign n19603 = ~n34749 & ~n18949;
  assign n19604 = ~n18949 & ~n19401;
  assign n19605 = ~n34749 & n19604;
  assign n19606 = ~n19401 & n19603;
  assign n19607 = n18804 & ~n34835;
  assign n19608 = n18948 & n19604;
  assign n19609 = n18804 & ~n34749;
  assign n19610 = ~n18949 & n19609;
  assign n19611 = ~n19401 & n19610;
  assign n19612 = ~n18804 & ~n34835;
  assign n19613 = ~n19611 & ~n19612;
  assign n19614 = ~n19607 & ~n19608;
  assign n19615 = ~n19602 & ~n34836;
  assign n19616 = ~n19600 & ~n19615;
  assign n19617 = ~n10681 & ~n19616;
  assign n19618 = n10681 & ~n19600;
  assign n19619 = ~n19615 & n19618;
  assign n19620 = n10681 & n19616;
  assign n19621 = ~n18951 & ~n18965;
  assign n19622 = ~n18965 & ~n19401;
  assign n19623 = ~n18951 & n19622;
  assign n19624 = ~n19401 & n19621;
  assign n19625 = ~n34751 & ~n34838;
  assign n19626 = n18963 & n19622;
  assign n19627 = n34751 & n34838;
  assign n19628 = ~n34751 & ~n18965;
  assign n19629 = ~n18951 & n19628;
  assign n19630 = ~n19401 & n19629;
  assign n19631 = n34751 & ~n34838;
  assign n19632 = ~n19630 & ~n19631;
  assign n19633 = ~n19625 & ~n34839;
  assign n19634 = ~n34837 & ~n34840;
  assign n19635 = ~n19617 & ~n19634;
  assign n19636 = ~n10086 & ~n19635;
  assign n19637 = n10086 & ~n19617;
  assign n19638 = ~n19634 & n19637;
  assign n19639 = ~n34752 & ~n18971;
  assign n19640 = ~n18971 & ~n19401;
  assign n19641 = ~n34752 & n19640;
  assign n19642 = ~n19401 & n19639;
  assign n19643 = n18796 & ~n34841;
  assign n19644 = n18970 & n19640;
  assign n19645 = n18796 & ~n34752;
  assign n19646 = ~n18971 & n19645;
  assign n19647 = ~n19401 & n19646;
  assign n19648 = ~n18796 & ~n34841;
  assign n19649 = ~n19647 & ~n19648;
  assign n19650 = ~n19643 & ~n19644;
  assign n19651 = ~n19638 & ~n34842;
  assign n19652 = ~n19636 & ~n19651;
  assign n19653 = ~n9565 & ~n19652;
  assign n19654 = n9565 & ~n19636;
  assign n19655 = ~n19651 & n19654;
  assign n19656 = n9565 & n19652;
  assign n19657 = ~n18973 & ~n18989;
  assign n19658 = ~n19401 & n19657;
  assign n19659 = ~n34755 & ~n19658;
  assign n19660 = n34755 & ~n18989;
  assign n19661 = ~n18973 & n19660;
  assign n19662 = n34755 & n19658;
  assign n19663 = ~n19401 & n19661;
  assign n19664 = ~n19659 & ~n34844;
  assign n19665 = ~n34843 & ~n19664;
  assign n19666 = ~n19653 & ~n19665;
  assign n19667 = ~n8998 & ~n19666;
  assign n19668 = n8998 & ~n19653;
  assign n19669 = ~n19665 & n19668;
  assign n19670 = ~n34756 & ~n18995;
  assign n19671 = ~n18995 & ~n19401;
  assign n19672 = ~n34756 & n19671;
  assign n19673 = ~n19401 & n19670;
  assign n19674 = n18788 & ~n34845;
  assign n19675 = n18994 & n19671;
  assign n19676 = n18788 & ~n34756;
  assign n19677 = ~n18995 & n19676;
  assign n19678 = ~n19401 & n19677;
  assign n19679 = ~n18788 & ~n34845;
  assign n19680 = ~n19678 & ~n19679;
  assign n19681 = ~n19674 & ~n19675;
  assign n19682 = ~n19669 & ~n34846;
  assign n19683 = ~n19667 & ~n19682;
  assign n19684 = ~n8506 & ~n19683;
  assign n19685 = n8506 & ~n19667;
  assign n19686 = ~n19682 & n19685;
  assign n19687 = n8506 & n19683;
  assign n19688 = ~n18997 & ~n19008;
  assign n19689 = ~n19008 & ~n19401;
  assign n19690 = ~n18997 & n19689;
  assign n19691 = ~n19401 & n19688;
  assign n19692 = n19005 & ~n34848;
  assign n19693 = n19006 & n19689;
  assign n19694 = ~n19005 & n34848;
  assign n19695 = n19005 & ~n19008;
  assign n19696 = ~n18997 & n19695;
  assign n19697 = ~n19401 & n19696;
  assign n19698 = ~n19005 & ~n34848;
  assign n19699 = ~n19697 & ~n19698;
  assign n19700 = ~n19692 & ~n34849;
  assign n19701 = ~n34847 & ~n34850;
  assign n19702 = ~n19684 & ~n19701;
  assign n19703 = ~n7975 & ~n19702;
  assign n19704 = n7975 & ~n19684;
  assign n19705 = ~n19701 & n19704;
  assign n19706 = ~n34758 & ~n19014;
  assign n19707 = ~n19014 & ~n19401;
  assign n19708 = ~n34758 & n19707;
  assign n19709 = ~n19401 & n19706;
  assign n19710 = n18780 & ~n34851;
  assign n19711 = n19013 & n19707;
  assign n19712 = n18780 & ~n34758;
  assign n19713 = ~n19014 & n19712;
  assign n19714 = ~n19401 & n19713;
  assign n19715 = ~n18780 & ~n34851;
  assign n19716 = ~n19714 & ~n19715;
  assign n19717 = ~n19710 & ~n19711;
  assign n19718 = ~n19705 & ~n34852;
  assign n19719 = ~n19703 & ~n19718;
  assign n19720 = ~n7512 & ~n19719;
  assign n19721 = n7512 & ~n19703;
  assign n19722 = ~n19718 & n19721;
  assign n19723 = n7512 & n19719;
  assign n19724 = ~n19016 & ~n19032;
  assign n19725 = ~n19401 & n19724;
  assign n19726 = ~n34761 & n19725;
  assign n19727 = n34761 & ~n19725;
  assign n19728 = n34761 & ~n19032;
  assign n19729 = ~n19016 & n19728;
  assign n19730 = n34761 & n19725;
  assign n19731 = ~n19401 & n19729;
  assign n19732 = ~n34761 & ~n19725;
  assign n19733 = ~n34854 & ~n19732;
  assign n19734 = ~n19726 & ~n19727;
  assign n19735 = ~n34853 & ~n34855;
  assign n19736 = ~n19720 & ~n19735;
  assign n19737 = ~n7015 & ~n19736;
  assign n19738 = n7015 & ~n19720;
  assign n19739 = ~n19735 & n19738;
  assign n19740 = ~n34762 & ~n19038;
  assign n19741 = ~n19038 & ~n19401;
  assign n19742 = ~n34762 & n19741;
  assign n19743 = ~n19401 & n19740;
  assign n19744 = n18772 & ~n34856;
  assign n19745 = n19037 & n19741;
  assign n19746 = n18772 & ~n34762;
  assign n19747 = ~n19038 & n19746;
  assign n19748 = ~n19401 & n19747;
  assign n19749 = ~n18772 & ~n34856;
  assign n19750 = ~n19748 & ~n19749;
  assign n19751 = ~n19744 & ~n19745;
  assign n19752 = ~n19739 & ~n34857;
  assign n19753 = ~n19737 & ~n19752;
  assign n19754 = ~n6579 & ~n19753;
  assign n19755 = n6579 & ~n19737;
  assign n19756 = ~n19752 & n19755;
  assign n19757 = n6579 & n19753;
  assign n19758 = ~n19040 & ~n19054;
  assign n19759 = ~n19054 & ~n19401;
  assign n19760 = ~n19040 & n19759;
  assign n19761 = ~n19401 & n19758;
  assign n19762 = n34764 & ~n34859;
  assign n19763 = n19052 & n19759;
  assign n19764 = ~n34764 & n34859;
  assign n19765 = n34764 & ~n19054;
  assign n19766 = ~n19040 & n19765;
  assign n19767 = ~n19401 & n19766;
  assign n19768 = ~n34764 & ~n34859;
  assign n19769 = ~n19767 & ~n19768;
  assign n19770 = ~n19762 & ~n34860;
  assign n19771 = ~n34858 & ~n34861;
  assign n19772 = ~n19754 & ~n19771;
  assign n19773 = ~n6117 & ~n19772;
  assign n19774 = n6117 & ~n19754;
  assign n19775 = ~n19771 & n19774;
  assign n19776 = ~n34765 & ~n19060;
  assign n19777 = ~n19060 & ~n19401;
  assign n19778 = ~n34765 & n19777;
  assign n19779 = ~n19401 & n19776;
  assign n19780 = n18764 & ~n34862;
  assign n19781 = n19059 & n19777;
  assign n19782 = n18764 & ~n34765;
  assign n19783 = ~n19060 & n19782;
  assign n19784 = ~n19401 & n19783;
  assign n19785 = ~n18764 & ~n34862;
  assign n19786 = ~n19784 & ~n19785;
  assign n19787 = ~n19780 & ~n19781;
  assign n19788 = ~n19775 & ~n34863;
  assign n19789 = ~n19773 & ~n19788;
  assign n19790 = ~n5708 & ~n19789;
  assign n19791 = ~n19062 & ~n19078;
  assign n19792 = ~n19401 & n19791;
  assign n19793 = ~n34768 & ~n19792;
  assign n19794 = n34768 & ~n19078;
  assign n19795 = ~n19062 & n19794;
  assign n19796 = n34768 & n19792;
  assign n19797 = ~n19401 & n19795;
  assign n19798 = ~n19793 & ~n34864;
  assign n19799 = n5708 & ~n19773;
  assign n19800 = ~n19788 & n19799;
  assign n19801 = n5708 & n19789;
  assign n19802 = ~n19798 & ~n34865;
  assign n19803 = ~n19790 & ~n19802;
  assign n19804 = ~n5278 & ~n19803;
  assign n19805 = n5278 & ~n19790;
  assign n19806 = ~n19802 & n19805;
  assign n19807 = ~n34769 & ~n19084;
  assign n19808 = ~n19084 & ~n19401;
  assign n19809 = ~n34769 & n19808;
  assign n19810 = ~n19401 & n19807;
  assign n19811 = n18756 & ~n34866;
  assign n19812 = n19083 & n19808;
  assign n19813 = n18756 & ~n34769;
  assign n19814 = ~n19084 & n19813;
  assign n19815 = ~n19401 & n19814;
  assign n19816 = ~n18756 & ~n34866;
  assign n19817 = ~n19815 & ~n19816;
  assign n19818 = ~n19811 & ~n19812;
  assign n19819 = ~n19806 & ~n34867;
  assign n19820 = ~n19804 & ~n19819;
  assign n19821 = ~n4903 & ~n19820;
  assign n19822 = n4903 & ~n19804;
  assign n19823 = ~n19819 & n19822;
  assign n19824 = n4903 & n19820;
  assign n19825 = ~n19086 & ~n19089;
  assign n19826 = ~n19089 & ~n19401;
  assign n19827 = ~n19086 & n19826;
  assign n19828 = ~n19401 & n19825;
  assign n19829 = n18748 & ~n34869;
  assign n19830 = n19087 & n19826;
  assign n19831 = n18748 & ~n19089;
  assign n19832 = ~n19086 & n19831;
  assign n19833 = ~n19401 & n19832;
  assign n19834 = ~n18748 & ~n34869;
  assign n19835 = ~n19833 & ~n19834;
  assign n19836 = ~n19829 & ~n19830;
  assign n19837 = ~n34868 & ~n34870;
  assign n19838 = ~n19821 & ~n19837;
  assign n19839 = ~n4508 & ~n19838;
  assign n19840 = n4508 & ~n19821;
  assign n19841 = ~n19837 & n19840;
  assign n19842 = ~n34770 & ~n19095;
  assign n19843 = ~n19095 & ~n19401;
  assign n19844 = ~n34770 & n19843;
  assign n19845 = ~n19401 & n19842;
  assign n19846 = n18740 & ~n34871;
  assign n19847 = n19094 & n19843;
  assign n19848 = n18740 & ~n34770;
  assign n19849 = ~n19095 & n19848;
  assign n19850 = ~n19401 & n19849;
  assign n19851 = ~n18740 & ~n34871;
  assign n19852 = ~n19850 & ~n19851;
  assign n19853 = ~n19846 & ~n19847;
  assign n19854 = ~n19841 & ~n34872;
  assign n19855 = ~n19839 & ~n19854;
  assign n19856 = ~n4155 & ~n19855;
  assign n19857 = ~n19097 & ~n19112;
  assign n19858 = ~n19401 & n19857;
  assign n19859 = ~n34772 & ~n19858;
  assign n19860 = n34772 & ~n19112;
  assign n19861 = ~n19097 & n19860;
  assign n19862 = n34772 & n19858;
  assign n19863 = ~n19401 & n19861;
  assign n19864 = ~n19859 & ~n34873;
  assign n19865 = n4155 & ~n19839;
  assign n19866 = ~n19854 & n19865;
  assign n19867 = n4155 & n19855;
  assign n19868 = ~n19864 & ~n34874;
  assign n19869 = ~n19856 & ~n19868;
  assign n19870 = ~n3788 & ~n19869;
  assign n19871 = n3788 & ~n19856;
  assign n19872 = ~n19868 & n19871;
  assign n19873 = ~n34773 & ~n19118;
  assign n19874 = ~n19118 & ~n19401;
  assign n19875 = ~n34773 & n19874;
  assign n19876 = ~n19401 & n19873;
  assign n19877 = n18732 & ~n34875;
  assign n19878 = n19117 & n19874;
  assign n19879 = n18732 & ~n34773;
  assign n19880 = ~n19118 & n19879;
  assign n19881 = ~n19401 & n19880;
  assign n19882 = ~n18732 & ~n34875;
  assign n19883 = ~n19881 & ~n19882;
  assign n19884 = ~n19877 & ~n19878;
  assign n19885 = ~n19872 & ~n34876;
  assign n19886 = ~n19870 & ~n19885;
  assign n19887 = ~n3473 & ~n19886;
  assign n19888 = n3473 & ~n19870;
  assign n19889 = ~n19885 & n19888;
  assign n19890 = n3473 & n19886;
  assign n19891 = ~n19120 & ~n19123;
  assign n19892 = ~n19123 & ~n19401;
  assign n19893 = ~n19120 & n19892;
  assign n19894 = ~n19401 & n19891;
  assign n19895 = n18724 & ~n34878;
  assign n19896 = n19121 & n19892;
  assign n19897 = n18724 & ~n19123;
  assign n19898 = ~n19120 & n19897;
  assign n19899 = ~n19401 & n19898;
  assign n19900 = ~n18724 & ~n34878;
  assign n19901 = ~n19899 & ~n19900;
  assign n19902 = ~n19895 & ~n19896;
  assign n19903 = ~n34877 & ~n34879;
  assign n19904 = ~n19887 & ~n19903;
  assign n19905 = ~n3140 & ~n19904;
  assign n19906 = n3140 & ~n19887;
  assign n19907 = ~n19903 & n19906;
  assign n19908 = ~n34774 & ~n19129;
  assign n19909 = ~n19129 & ~n19401;
  assign n19910 = ~n34774 & n19909;
  assign n19911 = ~n19401 & n19908;
  assign n19912 = n18716 & ~n34880;
  assign n19913 = n19128 & n19909;
  assign n19914 = n18716 & ~n34774;
  assign n19915 = ~n19129 & n19914;
  assign n19916 = ~n19401 & n19915;
  assign n19917 = ~n18716 & ~n34880;
  assign n19918 = ~n19916 & ~n19917;
  assign n19919 = ~n19912 & ~n19913;
  assign n19920 = ~n19907 & ~n34881;
  assign n19921 = ~n19905 & ~n19920;
  assign n19922 = ~n2855 & ~n19921;
  assign n19923 = ~n19131 & ~n19146;
  assign n19924 = ~n19401 & n19923;
  assign n19925 = ~n34776 & ~n19924;
  assign n19926 = n34776 & ~n19146;
  assign n19927 = ~n19131 & n19926;
  assign n19928 = n34776 & n19924;
  assign n19929 = ~n19401 & n19927;
  assign n19930 = ~n19925 & ~n34882;
  assign n19931 = n2855 & ~n19905;
  assign n19932 = ~n19920 & n19931;
  assign n19933 = n2855 & n19921;
  assign n19934 = ~n19930 & ~n34883;
  assign n19935 = ~n19922 & ~n19934;
  assign n19936 = ~n2556 & ~n19935;
  assign n19937 = n2556 & ~n19922;
  assign n19938 = ~n19934 & n19937;
  assign n19939 = ~n34777 & ~n19152;
  assign n19940 = ~n19152 & ~n19401;
  assign n19941 = ~n34777 & n19940;
  assign n19942 = ~n19401 & n19939;
  assign n19943 = n18708 & ~n34884;
  assign n19944 = n19151 & n19940;
  assign n19945 = n18708 & ~n34777;
  assign n19946 = ~n19152 & n19945;
  assign n19947 = ~n19401 & n19946;
  assign n19948 = ~n18708 & ~n34884;
  assign n19949 = ~n19947 & ~n19948;
  assign n19950 = ~n19943 & ~n19944;
  assign n19951 = ~n19938 & ~n34885;
  assign n19952 = ~n19936 & ~n19951;
  assign n19953 = ~n2301 & ~n19952;
  assign n19954 = n2301 & ~n19936;
  assign n19955 = ~n19951 & n19954;
  assign n19956 = n2301 & n19952;
  assign n19957 = ~n19154 & ~n19157;
  assign n19958 = ~n19157 & ~n19401;
  assign n19959 = ~n19154 & n19958;
  assign n19960 = ~n19401 & n19957;
  assign n19961 = n18700 & ~n34887;
  assign n19962 = n19155 & n19958;
  assign n19963 = n18700 & ~n19157;
  assign n19964 = ~n19154 & n19963;
  assign n19965 = ~n19401 & n19964;
  assign n19966 = ~n18700 & ~n34887;
  assign n19967 = ~n19965 & ~n19966;
  assign n19968 = ~n19961 & ~n19962;
  assign n19969 = ~n34886 & ~n34888;
  assign n19970 = ~n19953 & ~n19969;
  assign n19971 = ~n2038 & ~n19970;
  assign n19972 = n2038 & ~n19953;
  assign n19973 = ~n19969 & n19972;
  assign n19974 = ~n34778 & ~n19163;
  assign n19975 = ~n19401 & n19974;
  assign n19976 = n18692 & ~n19975;
  assign n19977 = ~n18692 & n19975;
  assign n19978 = n18692 & ~n34778;
  assign n19979 = ~n19163 & n19978;
  assign n19980 = ~n19401 & n19979;
  assign n19981 = ~n18692 & ~n19975;
  assign n19982 = ~n19980 & ~n19981;
  assign n19983 = ~n19976 & ~n19977;
  assign n19984 = ~n19973 & ~n34889;
  assign n19985 = ~n19971 & ~n19984;
  assign n19986 = ~n1812 & ~n19985;
  assign n19987 = ~n19165 & ~n19167;
  assign n19988 = ~n19401 & n19987;
  assign n19989 = n34780 & ~n19988;
  assign n19990 = ~n19165 & ~n34780;
  assign n19991 = ~n19167 & n19990;
  assign n19992 = ~n34780 & n19988;
  assign n19993 = ~n19401 & n19991;
  assign n19994 = n34780 & n19988;
  assign n19995 = ~n34780 & ~n19988;
  assign n19996 = ~n19994 & ~n19995;
  assign n19997 = ~n19989 & ~n34890;
  assign n19998 = n1812 & ~n19971;
  assign n19999 = ~n19984 & n19998;
  assign n20000 = n1812 & n19985;
  assign n20001 = n34891 & ~n34892;
  assign n20002 = ~n19986 & ~n20001;
  assign n20003 = ~n1582 & ~n20002;
  assign n20004 = n1582 & ~n19986;
  assign n20005 = ~n20001 & n20004;
  assign n20006 = ~n34809 & ~n20005;
  assign n20007 = ~n20003 & ~n20006;
  assign n20008 = ~n1388 & ~n20007;
  assign n20009 = ~n19187 & ~n19189;
  assign n20010 = ~n19401 & n20009;
  assign n20011 = ~n34783 & ~n20010;
  assign n20012 = ~n19187 & n34783;
  assign n20013 = ~n19189 & n20012;
  assign n20014 = n34783 & n20010;
  assign n20015 = ~n19401 & n20013;
  assign n20016 = ~n20011 & ~n34893;
  assign n20017 = n1388 & ~n20003;
  assign n20018 = ~n20006 & n20017;
  assign n20019 = n1388 & n20007;
  assign n20020 = ~n20016 & ~n34894;
  assign n20021 = ~n20008 & ~n20020;
  assign n20022 = ~n1192 & ~n20021;
  assign n20023 = n1192 & ~n20008;
  assign n20024 = ~n20020 & n20023;
  assign n20025 = ~n19204 & ~n34785;
  assign n20026 = ~n19204 & ~n19401;
  assign n20027 = ~n34785 & n20026;
  assign n20028 = ~n19401 & n20025;
  assign n20029 = n19212 & ~n34895;
  assign n20030 = n19216 & n20026;
  assign n20031 = n19212 & ~n34785;
  assign n20032 = ~n19204 & n20031;
  assign n20033 = ~n19401 & n20032;
  assign n20034 = ~n19212 & ~n34895;
  assign n20035 = ~n20033 & ~n20034;
  assign n20036 = ~n20029 & ~n20030;
  assign n20037 = ~n20024 & ~n34896;
  assign n20038 = ~n20022 & ~n20037;
  assign n20039 = ~n1028 & ~n20038;
  assign n20040 = ~n19218 & ~n19220;
  assign n20041 = ~n19401 & n20040;
  assign n20042 = ~n34787 & ~n20041;
  assign n20043 = ~n19218 & n34787;
  assign n20044 = ~n19220 & n20043;
  assign n20045 = n34787 & n20041;
  assign n20046 = ~n19401 & n20044;
  assign n20047 = ~n20042 & ~n34897;
  assign n20048 = n1028 & ~n20022;
  assign n20049 = ~n20037 & n20048;
  assign n20050 = n1028 & n20038;
  assign n20051 = ~n20047 & ~n34898;
  assign n20052 = ~n20039 & ~n20051;
  assign n20053 = ~n866 & ~n20052;
  assign n20054 = n866 & ~n20039;
  assign n20055 = ~n20051 & n20054;
  assign n20056 = ~n19235 & ~n34789;
  assign n20057 = ~n19235 & ~n19401;
  assign n20058 = ~n34789 & n20057;
  assign n20059 = ~n19401 & n20056;
  assign n20060 = n19243 & ~n34899;
  assign n20061 = n19247 & n20057;
  assign n20062 = n19243 & ~n34789;
  assign n20063 = ~n19235 & n20062;
  assign n20064 = ~n19401 & n20063;
  assign n20065 = ~n19243 & ~n34899;
  assign n20066 = ~n20064 & ~n20065;
  assign n20067 = ~n20060 & ~n20061;
  assign n20068 = ~n20055 & ~n34900;
  assign n20069 = ~n20053 & ~n20068;
  assign n20070 = ~n730 & ~n20069;
  assign n20071 = n730 & ~n20053;
  assign n20072 = ~n20068 & n20071;
  assign n20073 = n730 & n20069;
  assign n20074 = ~n19249 & ~n19259;
  assign n20075 = ~n19249 & ~n19401;
  assign n20076 = ~n19259 & n20075;
  assign n20077 = ~n19401 & n20074;
  assign n20078 = n19257 & ~n34902;
  assign n20079 = n19260 & n20075;
  assign n20080 = ~n19249 & n19257;
  assign n20081 = ~n19259 & n20080;
  assign n20082 = ~n19401 & n20081;
  assign n20083 = ~n19257 & ~n34902;
  assign n20084 = ~n20082 & ~n20083;
  assign n20085 = ~n20078 & ~n20079;
  assign n20086 = ~n34901 & ~n34903;
  assign n20087 = ~n20070 & ~n20086;
  assign n20088 = ~n602 & ~n20087;
  assign n20089 = n602 & ~n20070;
  assign n20090 = ~n20086 & n20089;
  assign n20091 = ~n19262 & ~n34792;
  assign n20092 = ~n19262 & ~n19401;
  assign n20093 = ~n34792 & n20092;
  assign n20094 = ~n19401 & n20091;
  assign n20095 = n19270 & ~n34904;
  assign n20096 = n19274 & n20092;
  assign n20097 = n19270 & ~n34792;
  assign n20098 = ~n19262 & n20097;
  assign n20099 = ~n19401 & n20098;
  assign n20100 = ~n19270 & ~n34904;
  assign n20101 = ~n20099 & ~n20100;
  assign n20102 = ~n20095 & ~n20096;
  assign n20103 = ~n20090 & ~n34905;
  assign n20104 = ~n20088 & ~n20103;
  assign n20105 = ~n497 & ~n20104;
  assign n20106 = ~n19276 & ~n19278;
  assign n20107 = ~n19401 & n20106;
  assign n20108 = ~n34794 & ~n20107;
  assign n20109 = ~n19276 & n34794;
  assign n20110 = ~n19278 & n20109;
  assign n20111 = n34794 & n20107;
  assign n20112 = ~n19401 & n20110;
  assign n20113 = ~n20108 & ~n34906;
  assign n20114 = n497 & ~n20088;
  assign n20115 = ~n20103 & n20114;
  assign n20116 = n497 & n20104;
  assign n20117 = ~n20113 & ~n34907;
  assign n20118 = ~n20105 & ~n20117;
  assign n20119 = ~n403 & ~n20118;
  assign n20120 = n403 & ~n20105;
  assign n20121 = ~n20117 & n20120;
  assign n20122 = ~n19293 & ~n34796;
  assign n20123 = ~n19293 & ~n19401;
  assign n20124 = ~n34796 & n20123;
  assign n20125 = ~n19401 & n20122;
  assign n20126 = n19301 & ~n34908;
  assign n20127 = n19305 & n20123;
  assign n20128 = n19301 & ~n34796;
  assign n20129 = ~n19293 & n20128;
  assign n20130 = ~n19401 & n20129;
  assign n20131 = ~n19301 & ~n34908;
  assign n20132 = ~n20130 & ~n20131;
  assign n20133 = ~n20126 & ~n20127;
  assign n20134 = ~n20121 & ~n34909;
  assign n20135 = ~n20119 & ~n20134;
  assign n20136 = ~n330 & ~n20135;
  assign n20137 = n330 & ~n20119;
  assign n20138 = ~n20134 & n20137;
  assign n20139 = n330 & n20135;
  assign n20140 = ~n19307 & ~n19317;
  assign n20141 = ~n19307 & ~n19401;
  assign n20142 = ~n19317 & n20141;
  assign n20143 = ~n19401 & n20140;
  assign n20144 = n19315 & ~n34911;
  assign n20145 = n19318 & n20141;
  assign n20146 = ~n19307 & n19315;
  assign n20147 = ~n19317 & n20146;
  assign n20148 = ~n19401 & n20147;
  assign n20149 = ~n19315 & ~n34911;
  assign n20150 = ~n20148 & ~n20149;
  assign n20151 = ~n20144 & ~n20145;
  assign n20152 = ~n34910 & ~n34912;
  assign n20153 = ~n20136 & ~n20152;
  assign n20154 = ~n271 & ~n20153;
  assign n20155 = n271 & ~n20136;
  assign n20156 = ~n20152 & n20155;
  assign n20157 = ~n19320 & ~n34799;
  assign n20158 = ~n19320 & ~n19401;
  assign n20159 = ~n34799 & n20158;
  assign n20160 = ~n19401 & n20157;
  assign n20161 = n19328 & ~n34913;
  assign n20162 = n19332 & n20158;
  assign n20163 = n19328 & ~n34799;
  assign n20164 = ~n19320 & n20163;
  assign n20165 = ~n19401 & n20164;
  assign n20166 = ~n19328 & ~n34913;
  assign n20167 = ~n20165 & ~n20166;
  assign n20168 = ~n20161 & ~n20162;
  assign n20169 = ~n20156 & ~n34914;
  assign n20170 = ~n20154 & ~n20169;
  assign n20171 = ~n217 & ~n20170;
  assign n20172 = ~n19334 & ~n19336;
  assign n20173 = ~n19401 & n20172;
  assign n20174 = ~n34801 & ~n20173;
  assign n20175 = ~n19334 & n34801;
  assign n20176 = ~n19336 & n20175;
  assign n20177 = n34801 & n20173;
  assign n20178 = ~n19401 & n20176;
  assign n20179 = ~n20174 & ~n34915;
  assign n20180 = n217 & ~n20154;
  assign n20181 = ~n20169 & n20180;
  assign n20182 = n217 & n20170;
  assign n20183 = ~n20179 & ~n34916;
  assign n20184 = ~n20171 & ~n20183;
  assign n20185 = ~n198 & ~n20184;
  assign n20186 = n198 & ~n20171;
  assign n20187 = ~n20183 & n20186;
  assign n20188 = ~n19351 & ~n34803;
  assign n20189 = ~n19351 & ~n19401;
  assign n20190 = ~n34803 & n20189;
  assign n20191 = ~n19401 & n20188;
  assign n20192 = n19359 & ~n34917;
  assign n20193 = n19363 & n20189;
  assign n20194 = n19359 & ~n34803;
  assign n20195 = ~n19351 & n20194;
  assign n20196 = ~n19401 & n20195;
  assign n20197 = ~n19359 & ~n34917;
  assign n20198 = ~n20196 & ~n20197;
  assign n20199 = ~n20192 & ~n20193;
  assign n20200 = ~n20187 & ~n34918;
  assign n20201 = ~n20185 & ~n20200;
  assign n20202 = ~n19365 & ~n19375;
  assign n20203 = ~n19365 & ~n19401;
  assign n20204 = ~n19375 & n20203;
  assign n20205 = ~n19401 & n20202;
  assign n20206 = n19373 & ~n34919;
  assign n20207 = n19376 & n20203;
  assign n20208 = ~n19365 & n19373;
  assign n20209 = ~n19375 & n20208;
  assign n20210 = ~n19401 & n20209;
  assign n20211 = ~n19373 & ~n34919;
  assign n20212 = ~n20210 & ~n20211;
  assign n20213 = ~n20206 & ~n20207;
  assign n20214 = ~n19377 & ~n19385;
  assign n20215 = ~n19385 & ~n19401;
  assign n20216 = ~n19377 & n20215;
  assign n20217 = ~n19401 & n20214;
  assign n20218 = ~n34807 & ~n34921;
  assign n20219 = ~n34920 & n20218;
  assign n20220 = ~n20201 & n20219;
  assign n20221 = n193 & ~n20220;
  assign n20222 = ~n20185 & n34920;
  assign n20223 = ~n20200 & n20222;
  assign n20224 = n20201 & n34920;
  assign n20225 = n19377 & ~n20215;
  assign n20226 = ~n193 & ~n20214;
  assign n20227 = ~n20225 & n20226;
  assign n20228 = ~n34922 & ~n20227;
  assign n20229 = ~n20221 & n20228;
  assign n20230 = ~n20003 & ~n20005;
  assign n20231 = ~n20229 & n20230;
  assign n20232 = ~n34809 & ~n20231;
  assign n20233 = n34809 & ~n20005;
  assign n20234 = ~n20003 & n20233;
  assign n20235 = n34809 & n20231;
  assign n20236 = ~n20229 & n20234;
  assign n20237 = ~n20232 & ~n34923;
  assign n20238 = ~n19953 & ~n34886;
  assign n20239 = ~n20229 & n20238;
  assign n20240 = ~n34888 & ~n20239;
  assign n20241 = ~n19953 & n34888;
  assign n20242 = ~n34886 & n20241;
  assign n20243 = n34888 & n20239;
  assign n20244 = ~n20229 & n20242;
  assign n20245 = ~n20240 & ~n34924;
  assign n20246 = ~n19936 & ~n19938;
  assign n20247 = ~n20229 & n20246;
  assign n20248 = ~n34885 & ~n20247;
  assign n20249 = ~n19938 & n34885;
  assign n20250 = ~n19936 & n20249;
  assign n20251 = n34885 & n20247;
  assign n20252 = ~n20229 & n20250;
  assign n20253 = ~n20248 & ~n34925;
  assign n20254 = ~n19905 & ~n19907;
  assign n20255 = ~n20229 & n20254;
  assign n20256 = ~n34881 & ~n20255;
  assign n20257 = ~n19907 & n34881;
  assign n20258 = ~n19905 & n20257;
  assign n20259 = n34881 & n20255;
  assign n20260 = ~n20229 & n20258;
  assign n20261 = ~n20256 & ~n34926;
  assign n20262 = ~n19887 & ~n34877;
  assign n20263 = ~n20229 & n20262;
  assign n20264 = ~n34879 & ~n20263;
  assign n20265 = ~n19887 & n34879;
  assign n20266 = ~n34877 & n20265;
  assign n20267 = n34879 & n20263;
  assign n20268 = ~n20229 & n20266;
  assign n20269 = ~n20264 & ~n34927;
  assign n20270 = ~n19870 & ~n19872;
  assign n20271 = ~n20229 & n20270;
  assign n20272 = ~n34876 & ~n20271;
  assign n20273 = ~n19872 & n34876;
  assign n20274 = ~n19870 & n20273;
  assign n20275 = n34876 & n20271;
  assign n20276 = ~n20229 & n20274;
  assign n20277 = ~n20272 & ~n34928;
  assign n20278 = ~n19839 & ~n19841;
  assign n20279 = ~n20229 & n20278;
  assign n20280 = ~n34872 & ~n20279;
  assign n20281 = ~n19841 & n34872;
  assign n20282 = ~n19839 & n20281;
  assign n20283 = n34872 & n20279;
  assign n20284 = ~n20229 & n20282;
  assign n20285 = ~n20280 & ~n34929;
  assign n20286 = ~n19821 & ~n34868;
  assign n20287 = ~n20229 & n20286;
  assign n20288 = ~n34870 & ~n20287;
  assign n20289 = ~n19821 & n34870;
  assign n20290 = ~n34868 & n20289;
  assign n20291 = n34870 & n20287;
  assign n20292 = ~n20229 & n20290;
  assign n20293 = ~n20288 & ~n34930;
  assign n20294 = ~n19804 & ~n19806;
  assign n20295 = ~n20229 & n20294;
  assign n20296 = ~n34867 & ~n20295;
  assign n20297 = ~n19806 & n34867;
  assign n20298 = ~n19804 & n20297;
  assign n20299 = n34867 & n20295;
  assign n20300 = ~n20229 & n20298;
  assign n20301 = ~n20296 & ~n34931;
  assign n20302 = ~n19773 & ~n19775;
  assign n20303 = ~n20229 & n20302;
  assign n20304 = ~n34863 & ~n20303;
  assign n20305 = ~n19775 & n34863;
  assign n20306 = ~n19773 & n20305;
  assign n20307 = n34863 & n20303;
  assign n20308 = ~n20229 & n20306;
  assign n20309 = ~n20304 & ~n34932;
  assign n20310 = ~n19754 & ~n34858;
  assign n20311 = ~n20229 & n20310;
  assign n20312 = ~n34861 & ~n20311;
  assign n20313 = ~n19754 & n34861;
  assign n20314 = ~n34858 & n20313;
  assign n20315 = n34861 & n20311;
  assign n20316 = ~n20229 & n20314;
  assign n20317 = ~n20312 & ~n34933;
  assign n20318 = ~n19737 & ~n19739;
  assign n20319 = ~n20229 & n20318;
  assign n20320 = ~n34857 & ~n20319;
  assign n20321 = ~n19739 & n34857;
  assign n20322 = ~n19737 & n20321;
  assign n20323 = n34857 & n20319;
  assign n20324 = ~n20229 & n20322;
  assign n20325 = ~n20320 & ~n34934;
  assign n20326 = ~n19703 & ~n19705;
  assign n20327 = ~n20229 & n20326;
  assign n20328 = ~n34852 & ~n20327;
  assign n20329 = ~n19705 & n34852;
  assign n20330 = ~n19703 & n20329;
  assign n20331 = n34852 & n20327;
  assign n20332 = ~n20229 & n20330;
  assign n20333 = ~n20328 & ~n34935;
  assign n20334 = ~n19667 & ~n19669;
  assign n20335 = ~n20229 & n20334;
  assign n20336 = ~n34846 & ~n20335;
  assign n20337 = ~n19669 & n34846;
  assign n20338 = ~n19667 & n20337;
  assign n20339 = n34846 & n20335;
  assign n20340 = ~n20229 & n20338;
  assign n20341 = ~n20336 & ~n34936;
  assign n20342 = ~n19636 & ~n19638;
  assign n20343 = ~n20229 & n20342;
  assign n20344 = ~n34842 & ~n20343;
  assign n20345 = ~n19638 & n34842;
  assign n20346 = ~n19636 & n20345;
  assign n20347 = n34842 & n20343;
  assign n20348 = ~n20229 & n20346;
  assign n20349 = ~n20344 & ~n34937;
  assign n20350 = ~n19600 & ~n19602;
  assign n20351 = ~n20229 & n20350;
  assign n20352 = ~n34836 & ~n20351;
  assign n20353 = ~n19602 & n34836;
  assign n20354 = ~n19600 & n20353;
  assign n20355 = n34836 & n20351;
  assign n20356 = ~n20229 & n20354;
  assign n20357 = ~n20352 & ~n34938;
  assign n20358 = ~n19566 & ~n19568;
  assign n20359 = ~n20229 & n20358;
  assign n20360 = ~n34831 & ~n20359;
  assign n20361 = ~n19568 & n34831;
  assign n20362 = ~n19566 & n20361;
  assign n20363 = n34831 & n20359;
  assign n20364 = ~n20229 & n20362;
  assign n20365 = ~n20360 & ~n34939;
  assign n20366 = ~n19532 & ~n19534;
  assign n20367 = ~n20229 & n20366;
  assign n20368 = ~n34826 & ~n20367;
  assign n20369 = ~n19534 & n34826;
  assign n20370 = ~n19532 & n20369;
  assign n20371 = n34826 & n20367;
  assign n20372 = ~n20229 & n20370;
  assign n20373 = ~n20368 & ~n34940;
  assign n20374 = ~n19499 & ~n19501;
  assign n20375 = ~n20229 & n20374;
  assign n20376 = ~n34822 & ~n20375;
  assign n20377 = ~n19501 & n34822;
  assign n20378 = ~n19499 & n20377;
  assign n20379 = n34822 & n20375;
  assign n20380 = ~n20229 & n20378;
  assign n20381 = ~n20376 & ~n34941;
  assign n20382 = ~n19465 & ~n19467;
  assign n20383 = ~n20229 & n20382;
  assign n20384 = ~n34817 & ~n20383;
  assign n20385 = ~n19467 & n34817;
  assign n20386 = ~n19465 & n20385;
  assign n20387 = n34817 & n20383;
  assign n20388 = ~n20229 & n20386;
  assign n20389 = ~n20384 & ~n34942;
  assign n20390 = ~n19438 & ~n19440;
  assign n20391 = ~n20229 & n20390;
  assign n20392 = ~n19449 & ~n20391;
  assign n20393 = ~n19440 & n19449;
  assign n20394 = ~n19438 & n20393;
  assign n20395 = n19449 & n20391;
  assign n20396 = ~n20229 & n20394;
  assign n20397 = ~n20392 & ~n34943;
  assign n20398 = ~pi26  & ~n20229;
  assign n20399 = ~pi27  & n20398;
  assign n20400 = n19415 & ~n20229;
  assign n20401 = ~n19401 & ~n20227;
  assign n20402 = ~n34922 & n20401;
  assign n20403 = ~n20221 & n20402;
  assign n20404 = ~n34944 & ~n20403;
  assign n20405 = pi28  & ~n20404;
  assign n20406 = ~pi28  & ~n20403;
  assign n20407 = ~pi28  & n20404;
  assign n20408 = ~n34944 & n20406;
  assign n20409 = ~n20405 & ~n34945;
  assign n20410 = pi26  & ~n20229;
  assign n20411 = ~pi24  & ~pi25 ;
  assign n20412 = ~pi26  & n20411;
  assign n20413 = ~n34713 & ~n34811;
  assign n20414 = ~n18655 & n20413;
  assign n20415 = ~n18674 & n20414;
  assign n20416 = ~n34715 & n20415;
  assign n20417 = n18660 & n18676;
  assign n20418 = ~n18668 & n20416;
  assign n20419 = ~n20412 & ~n34946;
  assign n20420 = ~n19399 & n20419;
  assign n20421 = ~n34807 & n20420;
  assign n20422 = ~n19393 & n20421;
  assign n20423 = ~n20410 & ~n20412;
  assign n20424 = n19401 & n20423;
  assign n20425 = ~n20410 & n20422;
  assign n20426 = pi27  & ~n20398;
  assign n20427 = ~n34944 & ~n20426;
  assign n20428 = ~n34947 & n20427;
  assign n20429 = ~n19401 & ~n20423;
  assign n20430 = n18676 & ~n20429;
  assign n20431 = ~n20428 & ~n20429;
  assign n20432 = n18676 & n20431;
  assign n20433 = ~n20428 & n20430;
  assign n20434 = ~n20409 & ~n34948;
  assign n20435 = ~n18676 & ~n20431;
  assign n20436 = n17885 & ~n20435;
  assign n20437 = ~n20434 & n20436;
  assign n20438 = ~n19418 & ~n34812;
  assign n20439 = ~n20229 & n20438;
  assign n20440 = n19423 & ~n20439;
  assign n20441 = ~n19423 & n20438;
  assign n20442 = ~n19423 & n20439;
  assign n20443 = ~n20229 & n20441;
  assign n20444 = ~n20440 & ~n34949;
  assign n20445 = ~n20437 & ~n20444;
  assign n20446 = ~n20434 & ~n20435;
  assign n20447 = ~n17885 & ~n20446;
  assign n20448 = n17187 & ~n20447;
  assign n20449 = ~n20445 & ~n20447;
  assign n20450 = n17187 & n20449;
  assign n20451 = ~n20445 & n20448;
  assign n20452 = ~n20397 & ~n34950;
  assign n20453 = ~n17187 & ~n20449;
  assign n20454 = n16428 & ~n20453;
  assign n20455 = ~n20452 & n20454;
  assign n20456 = ~n19452 & ~n34814;
  assign n20457 = ~n20229 & n20456;
  assign n20458 = n19462 & ~n20457;
  assign n20459 = ~n19462 & n20457;
  assign n20460 = ~n19452 & n19462;
  assign n20461 = ~n34814 & n20460;
  assign n20462 = n19462 & n20457;
  assign n20463 = ~n20229 & n20461;
  assign n20464 = ~n19462 & ~n20457;
  assign n20465 = ~n34951 & ~n20464;
  assign n20466 = ~n20458 & ~n20459;
  assign n20467 = ~n20455 & ~n34952;
  assign n20468 = ~n20452 & ~n20453;
  assign n20469 = ~n16428 & ~n20468;
  assign n20470 = n15760 & ~n20469;
  assign n20471 = ~n20467 & ~n20469;
  assign n20472 = n15760 & n20471;
  assign n20473 = ~n20467 & n20470;
  assign n20474 = ~n20389 & ~n34953;
  assign n20475 = ~n15760 & ~n20471;
  assign n20476 = n15033 & ~n20475;
  assign n20477 = ~n20474 & n20476;
  assign n20478 = ~n19482 & ~n34818;
  assign n20479 = ~n20229 & n20478;
  assign n20480 = ~n34820 & n20479;
  assign n20481 = n34820 & ~n20479;
  assign n20482 = ~n19482 & n34820;
  assign n20483 = ~n34818 & n20482;
  assign n20484 = ~n20229 & n20483;
  assign n20485 = ~n34820 & ~n20479;
  assign n20486 = ~n20484 & ~n20485;
  assign n20487 = ~n20480 & ~n20481;
  assign n20488 = ~n20477 & ~n34954;
  assign n20489 = ~n20474 & ~n20475;
  assign n20490 = ~n15033 & ~n20489;
  assign n20491 = n14394 & ~n20490;
  assign n20492 = ~n20488 & ~n20490;
  assign n20493 = n14394 & n20492;
  assign n20494 = ~n20488 & n20491;
  assign n20495 = ~n20381 & ~n34955;
  assign n20496 = ~n14394 & ~n20492;
  assign n20497 = n13704 & ~n20496;
  assign n20498 = ~n20495 & n20497;
  assign n20499 = ~n19516 & ~n34823;
  assign n20500 = ~n20229 & n20499;
  assign n20501 = ~n34824 & ~n20500;
  assign n20502 = ~n19516 & n34824;
  assign n20503 = ~n34823 & n20502;
  assign n20504 = n34824 & n20500;
  assign n20505 = ~n20229 & n20503;
  assign n20506 = n34824 & ~n20500;
  assign n20507 = ~n34824 & n20500;
  assign n20508 = ~n20506 & ~n20507;
  assign n20509 = ~n20501 & ~n34956;
  assign n20510 = ~n20498 & n34957;
  assign n20511 = ~n20495 & ~n20496;
  assign n20512 = ~n13704 & ~n20511;
  assign n20513 = n13099 & ~n20512;
  assign n20514 = ~n20510 & ~n20512;
  assign n20515 = n13099 & n20514;
  assign n20516 = ~n20510 & n20513;
  assign n20517 = ~n20373 & ~n34958;
  assign n20518 = ~n13099 & ~n20514;
  assign n20519 = n12442 & ~n20518;
  assign n20520 = ~n20517 & n20519;
  assign n20521 = ~n19549 & ~n34827;
  assign n20522 = ~n20229 & n20521;
  assign n20523 = n34829 & ~n20522;
  assign n20524 = ~n19549 & ~n34829;
  assign n20525 = ~n34827 & n20524;
  assign n20526 = ~n34829 & n20522;
  assign n20527 = ~n20229 & n20525;
  assign n20528 = n34829 & n20522;
  assign n20529 = ~n34829 & ~n20522;
  assign n20530 = ~n20528 & ~n20529;
  assign n20531 = ~n20523 & ~n34959;
  assign n20532 = ~n20520 & n34960;
  assign n20533 = ~n20517 & ~n20518;
  assign n20534 = ~n12442 & ~n20533;
  assign n20535 = n11858 & ~n20534;
  assign n20536 = ~n20532 & ~n20534;
  assign n20537 = n11858 & n20536;
  assign n20538 = ~n20532 & n20535;
  assign n20539 = ~n20365 & ~n34961;
  assign n20540 = ~n11858 & ~n20536;
  assign n20541 = n11229 & ~n20540;
  assign n20542 = ~n20539 & n20541;
  assign n20543 = ~n19583 & ~n34832;
  assign n20544 = ~n19583 & ~n20229;
  assign n20545 = ~n34832 & n20544;
  assign n20546 = ~n20229 & n20543;
  assign n20547 = ~n34834 & ~n34962;
  assign n20548 = n19598 & n20544;
  assign n20549 = n34834 & n34962;
  assign n20550 = ~n19583 & ~n34834;
  assign n20551 = ~n34832 & n20550;
  assign n20552 = ~n20229 & n20551;
  assign n20553 = n34834 & ~n34962;
  assign n20554 = ~n20552 & ~n20553;
  assign n20555 = ~n20547 & ~n34963;
  assign n20556 = ~n20542 & ~n34964;
  assign n20557 = ~n20539 & ~n20540;
  assign n20558 = ~n11229 & ~n20557;
  assign n20559 = n10681 & ~n20558;
  assign n20560 = ~n20556 & ~n20558;
  assign n20561 = n10681 & n20560;
  assign n20562 = ~n20556 & n20559;
  assign n20563 = ~n20357 & ~n34965;
  assign n20564 = ~n10681 & ~n20560;
  assign n20565 = n10086 & ~n20564;
  assign n20566 = ~n20563 & n20565;
  assign n20567 = ~n19617 & ~n34837;
  assign n20568 = ~n20229 & n20567;
  assign n20569 = ~n34840 & ~n20568;
  assign n20570 = ~n19617 & n34840;
  assign n20571 = ~n34837 & n20570;
  assign n20572 = n34840 & n20568;
  assign n20573 = ~n20229 & n20571;
  assign n20574 = ~n20569 & ~n34966;
  assign n20575 = ~n20566 & ~n20574;
  assign n20576 = ~n20563 & ~n20564;
  assign n20577 = ~n10086 & ~n20576;
  assign n20578 = n9565 & ~n20577;
  assign n20579 = ~n20575 & ~n20577;
  assign n20580 = n9565 & n20579;
  assign n20581 = ~n20575 & n20578;
  assign n20582 = ~n20349 & ~n34967;
  assign n20583 = ~n9565 & ~n20579;
  assign n20584 = n8998 & ~n20583;
  assign n20585 = ~n20582 & n20584;
  assign n20586 = ~n19653 & ~n34843;
  assign n20587 = ~n19653 & ~n20229;
  assign n20588 = ~n34843 & n20587;
  assign n20589 = ~n20229 & n20586;
  assign n20590 = n19664 & ~n34968;
  assign n20591 = n19665 & n20587;
  assign n20592 = ~n19664 & n34968;
  assign n20593 = ~n19653 & n19664;
  assign n20594 = ~n34843 & n20593;
  assign n20595 = ~n20229 & n20594;
  assign n20596 = ~n19664 & ~n34968;
  assign n20597 = ~n20595 & ~n20596;
  assign n20598 = ~n20590 & ~n34969;
  assign n20599 = ~n20585 & ~n34970;
  assign n20600 = ~n20582 & ~n20583;
  assign n20601 = ~n8998 & ~n20600;
  assign n20602 = n8506 & ~n20601;
  assign n20603 = ~n20599 & ~n20601;
  assign n20604 = n8506 & n20603;
  assign n20605 = ~n20599 & n20602;
  assign n20606 = ~n20341 & ~n34971;
  assign n20607 = ~n8506 & ~n20603;
  assign n20608 = n7975 & ~n20607;
  assign n20609 = ~n20606 & n20608;
  assign n20610 = ~n19684 & ~n34847;
  assign n20611 = ~n20229 & n20610;
  assign n20612 = ~n34850 & n20611;
  assign n20613 = n34850 & ~n20611;
  assign n20614 = ~n19684 & n34850;
  assign n20615 = ~n34847 & n20614;
  assign n20616 = n34850 & n20611;
  assign n20617 = ~n20229 & n20615;
  assign n20618 = ~n34850 & ~n20611;
  assign n20619 = ~n34972 & ~n20618;
  assign n20620 = ~n20612 & ~n20613;
  assign n20621 = ~n20609 & ~n34973;
  assign n20622 = ~n20606 & ~n20607;
  assign n20623 = ~n7975 & ~n20622;
  assign n20624 = n7512 & ~n20623;
  assign n20625 = ~n20621 & ~n20623;
  assign n20626 = n7512 & n20625;
  assign n20627 = ~n20621 & n20624;
  assign n20628 = ~n20333 & ~n34974;
  assign n20629 = ~n7512 & ~n20625;
  assign n20630 = n7015 & ~n20629;
  assign n20631 = ~n20628 & n20630;
  assign n20632 = ~n19720 & ~n34853;
  assign n20633 = ~n19720 & ~n20229;
  assign n20634 = ~n34853 & n20633;
  assign n20635 = ~n20229 & n20632;
  assign n20636 = n34855 & ~n34975;
  assign n20637 = n19735 & n20633;
  assign n20638 = ~n34855 & n34975;
  assign n20639 = ~n19720 & n34855;
  assign n20640 = ~n34853 & n20639;
  assign n20641 = ~n20229 & n20640;
  assign n20642 = ~n34855 & ~n34975;
  assign n20643 = ~n20641 & ~n20642;
  assign n20644 = ~n20636 & ~n34976;
  assign n20645 = ~n20631 & ~n34977;
  assign n20646 = ~n20628 & ~n20629;
  assign n20647 = ~n7015 & ~n20646;
  assign n20648 = n6579 & ~n20647;
  assign n20649 = ~n20645 & ~n20647;
  assign n20650 = n6579 & n20649;
  assign n20651 = ~n20645 & n20648;
  assign n20652 = ~n20325 & ~n34978;
  assign n20653 = ~n6579 & ~n20649;
  assign n20654 = n6117 & ~n20653;
  assign n20655 = ~n20652 & n20654;
  assign n20656 = ~n20317 & ~n20655;
  assign n20657 = ~n20652 & ~n20653;
  assign n20658 = ~n6117 & ~n20657;
  assign n20659 = n5708 & ~n20658;
  assign n20660 = ~n20656 & ~n20658;
  assign n20661 = n5708 & n20660;
  assign n20662 = ~n20656 & n20659;
  assign n20663 = ~n20309 & ~n34979;
  assign n20664 = ~n5708 & ~n20660;
  assign n20665 = n5278 & ~n20664;
  assign n20666 = ~n20663 & n20665;
  assign n20667 = ~n19790 & ~n34865;
  assign n20668 = ~n19790 & ~n20229;
  assign n20669 = ~n34865 & n20668;
  assign n20670 = ~n20229 & n20667;
  assign n20671 = n19798 & ~n34980;
  assign n20672 = n19802 & n20668;
  assign n20673 = ~n19790 & n19798;
  assign n20674 = ~n34865 & n20673;
  assign n20675 = ~n20229 & n20674;
  assign n20676 = ~n19798 & ~n34980;
  assign n20677 = ~n20675 & ~n20676;
  assign n20678 = ~n20671 & ~n20672;
  assign n20679 = ~n20666 & ~n34981;
  assign n20680 = ~n20663 & ~n20664;
  assign n20681 = ~n5278 & ~n20680;
  assign n20682 = n4903 & ~n20681;
  assign n20683 = ~n20679 & ~n20681;
  assign n20684 = n4903 & n20683;
  assign n20685 = ~n20679 & n20682;
  assign n20686 = ~n20301 & ~n34982;
  assign n20687 = ~n4903 & ~n20683;
  assign n20688 = n4508 & ~n20687;
  assign n20689 = ~n20686 & n20688;
  assign n20690 = ~n20293 & ~n20689;
  assign n20691 = ~n20686 & ~n20687;
  assign n20692 = ~n4508 & ~n20691;
  assign n20693 = n4155 & ~n20692;
  assign n20694 = ~n20690 & ~n20692;
  assign n20695 = n4155 & n20694;
  assign n20696 = ~n20690 & n20693;
  assign n20697 = ~n20285 & ~n34983;
  assign n20698 = ~n4155 & ~n20694;
  assign n20699 = n3788 & ~n20698;
  assign n20700 = ~n20697 & n20699;
  assign n20701 = ~n19856 & ~n34874;
  assign n20702 = ~n19856 & ~n20229;
  assign n20703 = ~n34874 & n20702;
  assign n20704 = ~n20229 & n20701;
  assign n20705 = n19864 & ~n34984;
  assign n20706 = n19868 & n20702;
  assign n20707 = ~n19856 & n19864;
  assign n20708 = ~n34874 & n20707;
  assign n20709 = ~n20229 & n20708;
  assign n20710 = ~n19864 & ~n34984;
  assign n20711 = ~n20709 & ~n20710;
  assign n20712 = ~n20705 & ~n20706;
  assign n20713 = ~n20700 & ~n34985;
  assign n20714 = ~n20697 & ~n20698;
  assign n20715 = ~n3788 & ~n20714;
  assign n20716 = n3473 & ~n20715;
  assign n20717 = ~n20713 & ~n20715;
  assign n20718 = n3473 & n20717;
  assign n20719 = ~n20713 & n20716;
  assign n20720 = ~n20277 & ~n34986;
  assign n20721 = ~n3473 & ~n20717;
  assign n20722 = n3140 & ~n20721;
  assign n20723 = ~n20720 & n20722;
  assign n20724 = ~n20269 & ~n20723;
  assign n20725 = ~n20720 & ~n20721;
  assign n20726 = ~n3140 & ~n20725;
  assign n20727 = n2855 & ~n20726;
  assign n20728 = ~n20724 & ~n20726;
  assign n20729 = n2855 & n20728;
  assign n20730 = ~n20724 & n20727;
  assign n20731 = ~n20261 & ~n34987;
  assign n20732 = ~n2855 & ~n20728;
  assign n20733 = n2556 & ~n20732;
  assign n20734 = ~n20731 & n20733;
  assign n20735 = ~n19922 & ~n34883;
  assign n20736 = ~n19922 & ~n20229;
  assign n20737 = ~n34883 & n20736;
  assign n20738 = ~n20229 & n20735;
  assign n20739 = n19930 & ~n34988;
  assign n20740 = n19934 & n20736;
  assign n20741 = ~n19922 & n19930;
  assign n20742 = ~n34883 & n20741;
  assign n20743 = ~n20229 & n20742;
  assign n20744 = ~n19930 & ~n34988;
  assign n20745 = ~n20743 & ~n20744;
  assign n20746 = ~n20739 & ~n20740;
  assign n20747 = ~n20734 & ~n34989;
  assign n20748 = ~n20731 & ~n20732;
  assign n20749 = ~n2556 & ~n20748;
  assign n20750 = n2301 & ~n20749;
  assign n20751 = ~n20747 & ~n20749;
  assign n20752 = n2301 & n20751;
  assign n20753 = ~n20747 & n20750;
  assign n20754 = ~n20253 & ~n34990;
  assign n20755 = ~n2301 & ~n20751;
  assign n20756 = n2038 & ~n20755;
  assign n20757 = ~n20754 & n20756;
  assign n20758 = ~n20245 & ~n20757;
  assign n20759 = ~n20754 & ~n20755;
  assign n20760 = ~n2038 & ~n20759;
  assign n20761 = n1812 & ~n20760;
  assign n20762 = ~n20758 & ~n20760;
  assign n20763 = n1812 & n20762;
  assign n20764 = ~n20758 & n20761;
  assign n20765 = ~n19971 & ~n19973;
  assign n20766 = ~n20229 & n20765;
  assign n20767 = ~n34889 & n20766;
  assign n20768 = n34889 & ~n20766;
  assign n20769 = ~n19973 & n34889;
  assign n20770 = ~n19971 & n20769;
  assign n20771 = ~n20229 & n20770;
  assign n20772 = ~n34889 & ~n20766;
  assign n20773 = ~n20771 & ~n20772;
  assign n20774 = ~n20767 & ~n20768;
  assign n20775 = ~n34991 & ~n34992;
  assign n20776 = ~n1812 & ~n20762;
  assign n20777 = ~n20775 & ~n20776;
  assign n20778 = ~n1582 & ~n20777;
  assign n20779 = n1582 & ~n20776;
  assign n20780 = ~n20775 & n20779;
  assign n20781 = ~n19986 & ~n34892;
  assign n20782 = ~n20229 & n20781;
  assign n20783 = ~n34891 & ~n20782;
  assign n20784 = n34891 & n20782;
  assign n20785 = ~n19986 & ~n34891;
  assign n20786 = ~n34892 & n20785;
  assign n20787 = ~n20229 & n20786;
  assign n20788 = n34891 & ~n20782;
  assign n20789 = ~n20787 & ~n20788;
  assign n20790 = ~n20783 & ~n20784;
  assign n20791 = ~n20780 & ~n34993;
  assign n20792 = ~n20778 & ~n20791;
  assign n20793 = ~n1388 & ~n20792;
  assign n20794 = n1388 & ~n20778;
  assign n20795 = n1388 & n20792;
  assign n20796 = ~n20791 & n20794;
  assign n20797 = ~n20237 & ~n34994;
  assign n20798 = ~n20793 & ~n20797;
  assign n20799 = ~n1192 & ~n20798;
  assign n20800 = n1192 & ~n20793;
  assign n20801 = ~n20797 & n20800;
  assign n20802 = ~n20008 & ~n34894;
  assign n20803 = ~n20008 & ~n20229;
  assign n20804 = ~n34894 & n20803;
  assign n20805 = ~n20229 & n20802;
  assign n20806 = n20016 & ~n34995;
  assign n20807 = n20020 & n20803;
  assign n20808 = ~n20008 & n20016;
  assign n20809 = ~n34894 & n20808;
  assign n20810 = ~n20229 & n20809;
  assign n20811 = ~n20016 & ~n34995;
  assign n20812 = ~n20810 & ~n20811;
  assign n20813 = ~n20806 & ~n20807;
  assign n20814 = ~n20801 & ~n34996;
  assign n20815 = ~n20799 & ~n20814;
  assign n20816 = ~n1028 & ~n20815;
  assign n20817 = ~n20022 & ~n20024;
  assign n20818 = ~n20229 & n20817;
  assign n20819 = ~n34896 & ~n20818;
  assign n20820 = ~n20024 & n34896;
  assign n20821 = ~n20022 & n20820;
  assign n20822 = n34896 & n20818;
  assign n20823 = ~n20229 & n20821;
  assign n20824 = ~n20819 & ~n34997;
  assign n20825 = n1028 & ~n20799;
  assign n20826 = n1028 & n20815;
  assign n20827 = ~n20814 & n20825;
  assign n20828 = ~n20824 & ~n34998;
  assign n20829 = ~n20816 & ~n20828;
  assign n20830 = ~n866 & ~n20829;
  assign n20831 = n866 & ~n20816;
  assign n20832 = ~n20828 & n20831;
  assign n20833 = ~n20039 & ~n34898;
  assign n20834 = ~n20039 & ~n20229;
  assign n20835 = ~n34898 & n20834;
  assign n20836 = ~n20229 & n20833;
  assign n20837 = n20047 & ~n34999;
  assign n20838 = n20051 & n20834;
  assign n20839 = ~n20039 & n20047;
  assign n20840 = ~n34898 & n20839;
  assign n20841 = ~n20229 & n20840;
  assign n20842 = ~n20047 & ~n34999;
  assign n20843 = ~n20841 & ~n20842;
  assign n20844 = ~n20837 & ~n20838;
  assign n20845 = ~n20832 & ~n35000;
  assign n20846 = ~n20830 & ~n20845;
  assign n20847 = ~n730 & ~n20846;
  assign n20848 = ~n20053 & ~n20055;
  assign n20849 = ~n20229 & n20848;
  assign n20850 = ~n34900 & ~n20849;
  assign n20851 = ~n20055 & n34900;
  assign n20852 = ~n20053 & n20851;
  assign n20853 = n34900 & n20849;
  assign n20854 = ~n20229 & n20852;
  assign n20855 = ~n20850 & ~n35001;
  assign n20856 = n730 & ~n20830;
  assign n20857 = n730 & n20846;
  assign n20858 = ~n20845 & n20856;
  assign n20859 = ~n20855 & ~n35002;
  assign n20860 = ~n20847 & ~n20859;
  assign n20861 = ~n602 & ~n20860;
  assign n20862 = ~n20070 & ~n34901;
  assign n20863 = ~n20229 & n20862;
  assign n20864 = ~n34903 & ~n20863;
  assign n20865 = ~n20070 & n34903;
  assign n20866 = ~n34901 & n20865;
  assign n20867 = n34903 & n20863;
  assign n20868 = ~n20229 & n20866;
  assign n20869 = ~n20864 & ~n35003;
  assign n20870 = n602 & ~n20847;
  assign n20871 = ~n20859 & n20870;
  assign n20872 = ~n20869 & ~n20871;
  assign n20873 = ~n20861 & ~n20872;
  assign n20874 = ~n497 & ~n20873;
  assign n20875 = ~n20088 & ~n20090;
  assign n20876 = ~n20229 & n20875;
  assign n20877 = ~n34905 & ~n20876;
  assign n20878 = ~n20090 & n34905;
  assign n20879 = ~n20088 & n20878;
  assign n20880 = n34905 & n20876;
  assign n20881 = ~n20229 & n20879;
  assign n20882 = ~n20877 & ~n35004;
  assign n20883 = n497 & ~n20861;
  assign n20884 = n497 & n20873;
  assign n20885 = ~n20872 & n20883;
  assign n20886 = ~n20882 & ~n35005;
  assign n20887 = ~n20874 & ~n20886;
  assign n20888 = ~n403 & ~n20887;
  assign n20889 = n403 & ~n20874;
  assign n20890 = ~n20886 & n20889;
  assign n20891 = ~n20105 & ~n34907;
  assign n20892 = ~n20105 & ~n20229;
  assign n20893 = ~n34907 & n20892;
  assign n20894 = ~n20229 & n20891;
  assign n20895 = n20113 & ~n35006;
  assign n20896 = n20117 & n20892;
  assign n20897 = ~n20105 & n20113;
  assign n20898 = ~n34907 & n20897;
  assign n20899 = ~n20229 & n20898;
  assign n20900 = ~n20113 & ~n35006;
  assign n20901 = ~n20899 & ~n20900;
  assign n20902 = ~n20895 & ~n20896;
  assign n20903 = ~n20890 & ~n35007;
  assign n20904 = ~n20888 & ~n20903;
  assign n20905 = ~n330 & ~n20904;
  assign n20906 = ~n20119 & ~n20121;
  assign n20907 = ~n20229 & n20906;
  assign n20908 = ~n34909 & ~n20907;
  assign n20909 = ~n20121 & n34909;
  assign n20910 = ~n20119 & n20909;
  assign n20911 = n34909 & n20907;
  assign n20912 = ~n20229 & n20910;
  assign n20913 = ~n20908 & ~n35008;
  assign n20914 = n330 & ~n20888;
  assign n20915 = n330 & n20904;
  assign n20916 = ~n20903 & n20914;
  assign n20917 = ~n20913 & ~n35009;
  assign n20918 = ~n20905 & ~n20917;
  assign n20919 = ~n271 & ~n20918;
  assign n20920 = ~n20136 & ~n34910;
  assign n20921 = ~n20229 & n20920;
  assign n20922 = ~n34912 & ~n20921;
  assign n20923 = ~n20136 & n34912;
  assign n20924 = ~n34910 & n20923;
  assign n20925 = n34912 & n20921;
  assign n20926 = ~n20229 & n20924;
  assign n20927 = ~n20922 & ~n35010;
  assign n20928 = n271 & ~n20905;
  assign n20929 = ~n20917 & n20928;
  assign n20930 = ~n20927 & ~n20929;
  assign n20931 = ~n20919 & ~n20930;
  assign n20932 = ~n217 & ~n20931;
  assign n20933 = ~n20154 & ~n20156;
  assign n20934 = ~n20229 & n20933;
  assign n20935 = ~n34914 & ~n20934;
  assign n20936 = ~n20156 & n34914;
  assign n20937 = ~n20154 & n20936;
  assign n20938 = n34914 & n20934;
  assign n20939 = ~n20229 & n20937;
  assign n20940 = ~n20935 & ~n35011;
  assign n20941 = n217 & ~n20919;
  assign n20942 = n217 & n20931;
  assign n20943 = ~n20930 & n20941;
  assign n20944 = ~n20940 & ~n35012;
  assign n20945 = ~n20932 & ~n20944;
  assign n20946 = ~n198 & ~n20945;
  assign n20947 = n198 & ~n20932;
  assign n20948 = ~n20944 & n20947;
  assign n20949 = ~n20171 & ~n34916;
  assign n20950 = ~n20171 & ~n20229;
  assign n20951 = ~n34916 & n20950;
  assign n20952 = ~n20229 & n20949;
  assign n20953 = n20179 & ~n35013;
  assign n20954 = n20183 & n20950;
  assign n20955 = ~n20171 & n20179;
  assign n20956 = ~n34916 & n20955;
  assign n20957 = ~n20229 & n20956;
  assign n20958 = ~n20179 & ~n35013;
  assign n20959 = ~n20957 & ~n20958;
  assign n20960 = ~n20953 & ~n20954;
  assign n20961 = ~n20948 & ~n35014;
  assign n20962 = ~n20946 & ~n20961;
  assign n20963 = ~n20185 & ~n20187;
  assign n20964 = ~n20229 & n20963;
  assign n20965 = ~n34918 & ~n20964;
  assign n20966 = ~n20187 & n34918;
  assign n20967 = ~n20185 & n20966;
  assign n20968 = n34918 & n20964;
  assign n20969 = ~n20229 & n20967;
  assign n20970 = ~n20965 & ~n35015;
  assign n20971 = ~n20201 & ~n34920;
  assign n20972 = ~n34920 & ~n20229;
  assign n20973 = ~n20201 & n20972;
  assign n20974 = ~n20229 & n20971;
  assign n20975 = ~n34922 & ~n35016;
  assign n20976 = ~n20970 & n20975;
  assign n20977 = ~n20962 & n20976;
  assign n20978 = n193 & ~n20977;
  assign n20979 = ~n20946 & n20970;
  assign n20980 = n20962 & n20970;
  assign n20981 = ~n20961 & n20979;
  assign n20982 = n20201 & ~n20972;
  assign n20983 = ~n193 & ~n20971;
  assign n20984 = ~n20982 & n20983;
  assign n20985 = ~n35017 & ~n20984;
  assign n20986 = ~n20978 & n20985;
  assign n20987 = ~n20793 & ~n34994;
  assign n20988 = ~n20793 & ~n20986;
  assign n20989 = ~n34994 & n20988;
  assign n20990 = ~n20986 & n20987;
  assign n20991 = n20237 & ~n35018;
  assign n20992 = n20797 & n20988;
  assign n20993 = n20237 & ~n34994;
  assign n20994 = ~n20793 & n20993;
  assign n20995 = ~n20986 & n20994;
  assign n20996 = ~n20237 & ~n35018;
  assign n20997 = ~n20995 & ~n20996;
  assign n20998 = ~n20991 & ~n20992;
  assign n20999 = pi24  & ~n20986;
  assign n21000 = ~pi22  & ~pi23 ;
  assign n21001 = ~pi24  & n21000;
  assign n21002 = ~n20999 & ~n21001;
  assign n21003 = ~n20229 & ~n21002;
  assign n21004 = ~pi24  & ~n20986;
  assign n21005 = pi25  & ~n21004;
  assign n21006 = ~pi25  & n21004;
  assign n21007 = n20411 & ~n20986;
  assign n21008 = ~n21005 & ~n35020;
  assign n21009 = ~n34805 & ~n34946;
  assign n21010 = ~n19380 & n21009;
  assign n21011 = ~n19399 & n21010;
  assign n21012 = ~n34807 & n21011;
  assign n21013 = n19385 & n19401;
  assign n21014 = ~n19393 & n21012;
  assign n21015 = ~n21001 & ~n35021;
  assign n21016 = ~n20227 & n21015;
  assign n21017 = ~n34922 & n21016;
  assign n21018 = ~n20221 & n21017;
  assign n21019 = n20229 & n21002;
  assign n21020 = ~n20999 & n21018;
  assign n21021 = n21008 & ~n35022;
  assign n21022 = ~n21003 & ~n21021;
  assign n21023 = ~n19401 & ~n21022;
  assign n21024 = n19401 & ~n21003;
  assign n21025 = ~n21021 & n21024;
  assign n21026 = ~n20229 & ~n20984;
  assign n21027 = ~n35017 & n21026;
  assign n21028 = ~n20978 & n21027;
  assign n21029 = ~n35020 & ~n21028;
  assign n21030 = pi26  & ~n21029;
  assign n21031 = ~pi26  & ~n21028;
  assign n21032 = ~pi26  & n21029;
  assign n21033 = ~n35020 & n21031;
  assign n21034 = ~n21030 & ~n35023;
  assign n21035 = ~n21025 & ~n21034;
  assign n21036 = ~n21023 & ~n21035;
  assign n21037 = ~n18676 & ~n21036;
  assign n21038 = n18676 & ~n21023;
  assign n21039 = ~n21035 & n21038;
  assign n21040 = n18676 & n21036;
  assign n21041 = ~n34947 & ~n20429;
  assign n21042 = ~n20986 & n21041;
  assign n21043 = n20427 & ~n21042;
  assign n21044 = ~n20427 & n21041;
  assign n21045 = ~n20427 & n21042;
  assign n21046 = ~n20986 & n21044;
  assign n21047 = ~n21043 & ~n35025;
  assign n21048 = ~n35024 & ~n21047;
  assign n21049 = ~n21037 & ~n21048;
  assign n21050 = ~n17885 & ~n21049;
  assign n21051 = n17885 & ~n21037;
  assign n21052 = ~n21048 & n21051;
  assign n21053 = ~n34948 & ~n20435;
  assign n21054 = ~n20435 & ~n20986;
  assign n21055 = ~n34948 & n21054;
  assign n21056 = ~n20986 & n21053;
  assign n21057 = n20409 & ~n35026;
  assign n21058 = n20434 & n21054;
  assign n21059 = n20409 & ~n34948;
  assign n21060 = ~n20435 & n21059;
  assign n21061 = ~n20986 & n21060;
  assign n21062 = ~n20409 & ~n35026;
  assign n21063 = ~n21061 & ~n21062;
  assign n21064 = ~n21057 & ~n21058;
  assign n21065 = ~n21052 & ~n35027;
  assign n21066 = ~n21050 & ~n21065;
  assign n21067 = ~n17187 & ~n21066;
  assign n21068 = n17187 & ~n21050;
  assign n21069 = ~n21065 & n21068;
  assign n21070 = n17187 & n21066;
  assign n21071 = ~n20437 & ~n20447;
  assign n21072 = ~n20986 & n21071;
  assign n21073 = n20444 & ~n21072;
  assign n21074 = ~n20444 & n21072;
  assign n21075 = n20444 & ~n20447;
  assign n21076 = ~n20437 & n21075;
  assign n21077 = n20444 & n21072;
  assign n21078 = ~n20986 & n21076;
  assign n21079 = ~n20444 & ~n21072;
  assign n21080 = ~n35029 & ~n21079;
  assign n21081 = ~n21073 & ~n21074;
  assign n21082 = ~n35028 & ~n35030;
  assign n21083 = ~n21067 & ~n21082;
  assign n21084 = ~n16428 & ~n21083;
  assign n21085 = n16428 & ~n21067;
  assign n21086 = ~n21082 & n21085;
  assign n21087 = ~n34950 & ~n20453;
  assign n21088 = ~n20453 & ~n20986;
  assign n21089 = ~n34950 & n21088;
  assign n21090 = ~n20986 & n21087;
  assign n21091 = n20397 & ~n35031;
  assign n21092 = n20452 & n21088;
  assign n21093 = n20397 & ~n34950;
  assign n21094 = ~n20453 & n21093;
  assign n21095 = ~n20986 & n21094;
  assign n21096 = ~n20397 & ~n35031;
  assign n21097 = ~n21095 & ~n21096;
  assign n21098 = ~n21091 & ~n21092;
  assign n21099 = ~n21086 & ~n35032;
  assign n21100 = ~n21084 & ~n21099;
  assign n21101 = ~n15760 & ~n21100;
  assign n21102 = n15760 & ~n21084;
  assign n21103 = ~n21099 & n21102;
  assign n21104 = n15760 & n21100;
  assign n21105 = ~n20455 & ~n20469;
  assign n21106 = ~n20986 & n21105;
  assign n21107 = ~n34952 & n21106;
  assign n21108 = n34952 & ~n21106;
  assign n21109 = n34952 & ~n20469;
  assign n21110 = ~n20455 & n21109;
  assign n21111 = ~n20986 & n21110;
  assign n21112 = ~n34952 & ~n21106;
  assign n21113 = ~n21111 & ~n21112;
  assign n21114 = ~n21107 & ~n21108;
  assign n21115 = ~n35033 & ~n35034;
  assign n21116 = ~n21101 & ~n21115;
  assign n21117 = ~n15033 & ~n21116;
  assign n21118 = n15033 & ~n21101;
  assign n21119 = ~n21115 & n21118;
  assign n21120 = ~n34953 & ~n20475;
  assign n21121 = ~n20475 & ~n20986;
  assign n21122 = ~n34953 & n21121;
  assign n21123 = ~n20986 & n21120;
  assign n21124 = n20389 & ~n35035;
  assign n21125 = n20474 & n21121;
  assign n21126 = n20389 & ~n34953;
  assign n21127 = ~n20475 & n21126;
  assign n21128 = ~n20986 & n21127;
  assign n21129 = ~n20389 & ~n35035;
  assign n21130 = ~n21128 & ~n21129;
  assign n21131 = ~n21124 & ~n21125;
  assign n21132 = ~n21119 & ~n35036;
  assign n21133 = ~n21117 & ~n21132;
  assign n21134 = ~n14394 & ~n21133;
  assign n21135 = n14394 & ~n21117;
  assign n21136 = ~n21132 & n21135;
  assign n21137 = n14394 & n21133;
  assign n21138 = ~n20477 & ~n20490;
  assign n21139 = ~n20986 & n21138;
  assign n21140 = ~n34954 & ~n21139;
  assign n21141 = n34954 & ~n20490;
  assign n21142 = ~n20477 & n21141;
  assign n21143 = n34954 & n21139;
  assign n21144 = ~n20986 & n21142;
  assign n21145 = n34954 & ~n21139;
  assign n21146 = ~n34954 & n21139;
  assign n21147 = ~n21145 & ~n21146;
  assign n21148 = ~n21140 & ~n35038;
  assign n21149 = ~n35037 & n35039;
  assign n21150 = ~n21134 & ~n21149;
  assign n21151 = ~n13704 & ~n21150;
  assign n21152 = n13704 & ~n21134;
  assign n21153 = ~n21149 & n21152;
  assign n21154 = ~n34955 & ~n20496;
  assign n21155 = ~n20496 & ~n20986;
  assign n21156 = ~n34955 & n21155;
  assign n21157 = ~n20986 & n21154;
  assign n21158 = n20381 & ~n35040;
  assign n21159 = n20495 & n21155;
  assign n21160 = n20381 & ~n34955;
  assign n21161 = ~n20496 & n21160;
  assign n21162 = ~n20986 & n21161;
  assign n21163 = ~n20381 & ~n35040;
  assign n21164 = ~n21162 & ~n21163;
  assign n21165 = ~n21158 & ~n21159;
  assign n21166 = ~n21153 & ~n35041;
  assign n21167 = ~n21151 & ~n21166;
  assign n21168 = ~n13099 & ~n21167;
  assign n21169 = n13099 & ~n21151;
  assign n21170 = ~n21166 & n21169;
  assign n21171 = n13099 & n21167;
  assign n21172 = ~n20498 & ~n20512;
  assign n21173 = ~n20986 & n21172;
  assign n21174 = n34957 & ~n21173;
  assign n21175 = ~n34957 & ~n20512;
  assign n21176 = ~n20498 & n21175;
  assign n21177 = ~n34957 & n21173;
  assign n21178 = ~n20986 & n21176;
  assign n21179 = n34957 & n21173;
  assign n21180 = ~n34957 & ~n21173;
  assign n21181 = ~n21179 & ~n21180;
  assign n21182 = ~n21174 & ~n35043;
  assign n21183 = ~n35042 & n35044;
  assign n21184 = ~n21168 & ~n21183;
  assign n21185 = ~n12442 & ~n21184;
  assign n21186 = n12442 & ~n21168;
  assign n21187 = ~n21183 & n21186;
  assign n21188 = ~n34958 & ~n20518;
  assign n21189 = ~n20518 & ~n20986;
  assign n21190 = ~n34958 & n21189;
  assign n21191 = ~n20986 & n21188;
  assign n21192 = n20373 & ~n35045;
  assign n21193 = n20517 & n21189;
  assign n21194 = n20373 & ~n34958;
  assign n21195 = ~n20518 & n21194;
  assign n21196 = ~n20986 & n21195;
  assign n21197 = ~n20373 & ~n35045;
  assign n21198 = ~n21196 & ~n21197;
  assign n21199 = ~n21192 & ~n21193;
  assign n21200 = ~n21187 & ~n35046;
  assign n21201 = ~n21185 & ~n21200;
  assign n21202 = ~n11858 & ~n21201;
  assign n21203 = n11858 & ~n21185;
  assign n21204 = ~n21200 & n21203;
  assign n21205 = n11858 & n21201;
  assign n21206 = ~n20520 & ~n20534;
  assign n21207 = ~n20534 & ~n20986;
  assign n21208 = ~n20520 & n21207;
  assign n21209 = ~n20986 & n21206;
  assign n21210 = ~n34960 & ~n35048;
  assign n21211 = n20532 & n21207;
  assign n21212 = n34960 & n35048;
  assign n21213 = ~n34960 & ~n20534;
  assign n21214 = ~n20520 & n21213;
  assign n21215 = ~n20986 & n21214;
  assign n21216 = n34960 & ~n35048;
  assign n21217 = ~n21215 & ~n21216;
  assign n21218 = ~n21210 & ~n35049;
  assign n21219 = ~n35047 & ~n35050;
  assign n21220 = ~n21202 & ~n21219;
  assign n21221 = ~n11229 & ~n21220;
  assign n21222 = n11229 & ~n21202;
  assign n21223 = ~n21219 & n21222;
  assign n21224 = ~n34961 & ~n20540;
  assign n21225 = ~n20540 & ~n20986;
  assign n21226 = ~n34961 & n21225;
  assign n21227 = ~n20986 & n21224;
  assign n21228 = n20365 & ~n35051;
  assign n21229 = n20539 & n21225;
  assign n21230 = n20365 & ~n34961;
  assign n21231 = ~n20540 & n21230;
  assign n21232 = ~n20986 & n21231;
  assign n21233 = ~n20365 & ~n35051;
  assign n21234 = ~n21232 & ~n21233;
  assign n21235 = ~n21228 & ~n21229;
  assign n21236 = ~n21223 & ~n35052;
  assign n21237 = ~n21221 & ~n21236;
  assign n21238 = ~n10681 & ~n21237;
  assign n21239 = n10681 & ~n21221;
  assign n21240 = ~n21236 & n21239;
  assign n21241 = n10681 & n21237;
  assign n21242 = ~n20542 & ~n20558;
  assign n21243 = ~n20986 & n21242;
  assign n21244 = ~n34964 & ~n21243;
  assign n21245 = n34964 & ~n20558;
  assign n21246 = ~n20542 & n21245;
  assign n21247 = n34964 & n21243;
  assign n21248 = ~n20986 & n21246;
  assign n21249 = ~n21244 & ~n35054;
  assign n21250 = ~n35053 & ~n21249;
  assign n21251 = ~n21238 & ~n21250;
  assign n21252 = ~n10086 & ~n21251;
  assign n21253 = n10086 & ~n21238;
  assign n21254 = ~n21250 & n21253;
  assign n21255 = ~n34965 & ~n20564;
  assign n21256 = ~n20564 & ~n20986;
  assign n21257 = ~n34965 & n21256;
  assign n21258 = ~n20986 & n21255;
  assign n21259 = n20357 & ~n35055;
  assign n21260 = n20563 & n21256;
  assign n21261 = n20357 & ~n34965;
  assign n21262 = ~n20564 & n21261;
  assign n21263 = ~n20986 & n21262;
  assign n21264 = ~n20357 & ~n35055;
  assign n21265 = ~n21263 & ~n21264;
  assign n21266 = ~n21259 & ~n21260;
  assign n21267 = ~n21254 & ~n35056;
  assign n21268 = ~n21252 & ~n21267;
  assign n21269 = ~n9565 & ~n21268;
  assign n21270 = n9565 & ~n21252;
  assign n21271 = ~n21267 & n21270;
  assign n21272 = n9565 & n21268;
  assign n21273 = ~n20566 & ~n20577;
  assign n21274 = ~n20577 & ~n20986;
  assign n21275 = ~n20566 & n21274;
  assign n21276 = ~n20986 & n21273;
  assign n21277 = n20574 & ~n35058;
  assign n21278 = n20575 & n21274;
  assign n21279 = ~n20574 & n35058;
  assign n21280 = n20574 & ~n20577;
  assign n21281 = ~n20566 & n21280;
  assign n21282 = ~n20986 & n21281;
  assign n21283 = ~n20574 & ~n35058;
  assign n21284 = ~n21282 & ~n21283;
  assign n21285 = ~n21277 & ~n35059;
  assign n21286 = ~n35057 & ~n35060;
  assign n21287 = ~n21269 & ~n21286;
  assign n21288 = ~n8998 & ~n21287;
  assign n21289 = n8998 & ~n21269;
  assign n21290 = ~n21286 & n21289;
  assign n21291 = ~n34967 & ~n20583;
  assign n21292 = ~n20583 & ~n20986;
  assign n21293 = ~n34967 & n21292;
  assign n21294 = ~n20986 & n21291;
  assign n21295 = n20349 & ~n35061;
  assign n21296 = n20582 & n21292;
  assign n21297 = n20349 & ~n34967;
  assign n21298 = ~n20583 & n21297;
  assign n21299 = ~n20986 & n21298;
  assign n21300 = ~n20349 & ~n35061;
  assign n21301 = ~n21299 & ~n21300;
  assign n21302 = ~n21295 & ~n21296;
  assign n21303 = ~n21290 & ~n35062;
  assign n21304 = ~n21288 & ~n21303;
  assign n21305 = ~n8506 & ~n21304;
  assign n21306 = n8506 & ~n21288;
  assign n21307 = ~n21303 & n21306;
  assign n21308 = n8506 & n21304;
  assign n21309 = ~n20585 & ~n20601;
  assign n21310 = ~n20986 & n21309;
  assign n21311 = ~n34970 & n21310;
  assign n21312 = n34970 & ~n21310;
  assign n21313 = n34970 & ~n20601;
  assign n21314 = ~n20585 & n21313;
  assign n21315 = n34970 & n21310;
  assign n21316 = ~n20986 & n21314;
  assign n21317 = ~n34970 & ~n21310;
  assign n21318 = ~n35064 & ~n21317;
  assign n21319 = ~n21311 & ~n21312;
  assign n21320 = ~n35063 & ~n35065;
  assign n21321 = ~n21305 & ~n21320;
  assign n21322 = ~n7975 & ~n21321;
  assign n21323 = n7975 & ~n21305;
  assign n21324 = ~n21320 & n21323;
  assign n21325 = ~n34971 & ~n20607;
  assign n21326 = ~n20607 & ~n20986;
  assign n21327 = ~n34971 & n21326;
  assign n21328 = ~n20986 & n21325;
  assign n21329 = n20341 & ~n35066;
  assign n21330 = n20606 & n21326;
  assign n21331 = n20341 & ~n34971;
  assign n21332 = ~n20607 & n21331;
  assign n21333 = ~n20986 & n21332;
  assign n21334 = ~n20341 & ~n35066;
  assign n21335 = ~n21333 & ~n21334;
  assign n21336 = ~n21329 & ~n21330;
  assign n21337 = ~n21324 & ~n35067;
  assign n21338 = ~n21322 & ~n21337;
  assign n21339 = ~n7512 & ~n21338;
  assign n21340 = n7512 & ~n21322;
  assign n21341 = ~n21337 & n21340;
  assign n21342 = n7512 & n21338;
  assign n21343 = ~n20609 & ~n20623;
  assign n21344 = ~n20623 & ~n20986;
  assign n21345 = ~n20609 & n21344;
  assign n21346 = ~n20986 & n21343;
  assign n21347 = n34973 & ~n35069;
  assign n21348 = n20621 & n21344;
  assign n21349 = ~n34973 & n35069;
  assign n21350 = n34973 & ~n20623;
  assign n21351 = ~n20609 & n21350;
  assign n21352 = ~n20986 & n21351;
  assign n21353 = ~n34973 & ~n35069;
  assign n21354 = ~n21352 & ~n21353;
  assign n21355 = ~n21347 & ~n35070;
  assign n21356 = ~n35068 & ~n35071;
  assign n21357 = ~n21339 & ~n21356;
  assign n21358 = ~n7015 & ~n21357;
  assign n21359 = n7015 & ~n21339;
  assign n21360 = ~n21356 & n21359;
  assign n21361 = ~n34974 & ~n20629;
  assign n21362 = ~n20629 & ~n20986;
  assign n21363 = ~n34974 & n21362;
  assign n21364 = ~n20986 & n21361;
  assign n21365 = n20333 & ~n35072;
  assign n21366 = n20628 & n21362;
  assign n21367 = n20333 & ~n34974;
  assign n21368 = ~n20629 & n21367;
  assign n21369 = ~n20986 & n21368;
  assign n21370 = ~n20333 & ~n35072;
  assign n21371 = ~n21369 & ~n21370;
  assign n21372 = ~n21365 & ~n21366;
  assign n21373 = ~n21360 & ~n35073;
  assign n21374 = ~n21358 & ~n21373;
  assign n21375 = ~n6579 & ~n21374;
  assign n21376 = ~n20631 & ~n20647;
  assign n21377 = ~n20986 & n21376;
  assign n21378 = ~n34977 & ~n21377;
  assign n21379 = n34977 & ~n20647;
  assign n21380 = ~n20631 & n21379;
  assign n21381 = n34977 & n21377;
  assign n21382 = ~n20986 & n21380;
  assign n21383 = ~n21378 & ~n35074;
  assign n21384 = n6579 & ~n21358;
  assign n21385 = ~n21373 & n21384;
  assign n21386 = n6579 & n21374;
  assign n21387 = ~n21383 & ~n35075;
  assign n21388 = ~n21375 & ~n21387;
  assign n21389 = ~n6117 & ~n21388;
  assign n21390 = n6117 & ~n21375;
  assign n21391 = ~n21387 & n21390;
  assign n21392 = ~n34978 & ~n20653;
  assign n21393 = ~n20653 & ~n20986;
  assign n21394 = ~n34978 & n21393;
  assign n21395 = ~n20986 & n21392;
  assign n21396 = n20325 & ~n35076;
  assign n21397 = n20652 & n21393;
  assign n21398 = n20325 & ~n34978;
  assign n21399 = ~n20653 & n21398;
  assign n21400 = ~n20986 & n21399;
  assign n21401 = ~n20325 & ~n35076;
  assign n21402 = ~n21400 & ~n21401;
  assign n21403 = ~n21396 & ~n21397;
  assign n21404 = ~n21391 & ~n35077;
  assign n21405 = ~n21389 & ~n21404;
  assign n21406 = ~n5708 & ~n21405;
  assign n21407 = n5708 & ~n21389;
  assign n21408 = ~n21404 & n21407;
  assign n21409 = n5708 & n21405;
  assign n21410 = ~n20655 & ~n20658;
  assign n21411 = ~n20658 & ~n20986;
  assign n21412 = ~n20655 & n21411;
  assign n21413 = ~n20986 & n21410;
  assign n21414 = n20317 & ~n35079;
  assign n21415 = n20656 & n21411;
  assign n21416 = n20317 & ~n20658;
  assign n21417 = ~n20655 & n21416;
  assign n21418 = ~n20986 & n21417;
  assign n21419 = ~n20317 & ~n35079;
  assign n21420 = ~n21418 & ~n21419;
  assign n21421 = ~n21414 & ~n21415;
  assign n21422 = ~n35078 & ~n35080;
  assign n21423 = ~n21406 & ~n21422;
  assign n21424 = ~n5278 & ~n21423;
  assign n21425 = n5278 & ~n21406;
  assign n21426 = ~n21422 & n21425;
  assign n21427 = ~n34979 & ~n20664;
  assign n21428 = ~n20664 & ~n20986;
  assign n21429 = ~n34979 & n21428;
  assign n21430 = ~n20986 & n21427;
  assign n21431 = n20309 & ~n35081;
  assign n21432 = n20663 & n21428;
  assign n21433 = n20309 & ~n34979;
  assign n21434 = ~n20664 & n21433;
  assign n21435 = ~n20986 & n21434;
  assign n21436 = ~n20309 & ~n35081;
  assign n21437 = ~n21435 & ~n21436;
  assign n21438 = ~n21431 & ~n21432;
  assign n21439 = ~n21426 & ~n35082;
  assign n21440 = ~n21424 & ~n21439;
  assign n21441 = ~n4903 & ~n21440;
  assign n21442 = ~n20666 & ~n20681;
  assign n21443 = ~n20986 & n21442;
  assign n21444 = ~n34981 & ~n21443;
  assign n21445 = n34981 & ~n20681;
  assign n21446 = ~n20666 & n21445;
  assign n21447 = n34981 & n21443;
  assign n21448 = ~n20986 & n21446;
  assign n21449 = ~n21444 & ~n35083;
  assign n21450 = n4903 & ~n21424;
  assign n21451 = ~n21439 & n21450;
  assign n21452 = n4903 & n21440;
  assign n21453 = ~n21449 & ~n35084;
  assign n21454 = ~n21441 & ~n21453;
  assign n21455 = ~n4508 & ~n21454;
  assign n21456 = n4508 & ~n21441;
  assign n21457 = ~n21453 & n21456;
  assign n21458 = ~n34982 & ~n20687;
  assign n21459 = ~n20687 & ~n20986;
  assign n21460 = ~n34982 & n21459;
  assign n21461 = ~n20986 & n21458;
  assign n21462 = n20301 & ~n35085;
  assign n21463 = n20686 & n21459;
  assign n21464 = n20301 & ~n34982;
  assign n21465 = ~n20687 & n21464;
  assign n21466 = ~n20986 & n21465;
  assign n21467 = ~n20301 & ~n35085;
  assign n21468 = ~n21466 & ~n21467;
  assign n21469 = ~n21462 & ~n21463;
  assign n21470 = ~n21457 & ~n35086;
  assign n21471 = ~n21455 & ~n21470;
  assign n21472 = ~n4155 & ~n21471;
  assign n21473 = n4155 & ~n21455;
  assign n21474 = ~n21470 & n21473;
  assign n21475 = n4155 & n21471;
  assign n21476 = ~n20689 & ~n20692;
  assign n21477 = ~n20692 & ~n20986;
  assign n21478 = ~n20689 & n21477;
  assign n21479 = ~n20986 & n21476;
  assign n21480 = n20293 & ~n35088;
  assign n21481 = n20690 & n21477;
  assign n21482 = n20293 & ~n20692;
  assign n21483 = ~n20689 & n21482;
  assign n21484 = ~n20986 & n21483;
  assign n21485 = ~n20293 & ~n35088;
  assign n21486 = ~n21484 & ~n21485;
  assign n21487 = ~n21480 & ~n21481;
  assign n21488 = ~n35087 & ~n35089;
  assign n21489 = ~n21472 & ~n21488;
  assign n21490 = ~n3788 & ~n21489;
  assign n21491 = n3788 & ~n21472;
  assign n21492 = ~n21488 & n21491;
  assign n21493 = ~n34983 & ~n20698;
  assign n21494 = ~n20698 & ~n20986;
  assign n21495 = ~n34983 & n21494;
  assign n21496 = ~n20986 & n21493;
  assign n21497 = n20285 & ~n35090;
  assign n21498 = n20697 & n21494;
  assign n21499 = n20285 & ~n34983;
  assign n21500 = ~n20698 & n21499;
  assign n21501 = ~n20986 & n21500;
  assign n21502 = ~n20285 & ~n35090;
  assign n21503 = ~n21501 & ~n21502;
  assign n21504 = ~n21497 & ~n21498;
  assign n21505 = ~n21492 & ~n35091;
  assign n21506 = ~n21490 & ~n21505;
  assign n21507 = ~n3473 & ~n21506;
  assign n21508 = ~n20700 & ~n20715;
  assign n21509 = ~n20986 & n21508;
  assign n21510 = ~n34985 & ~n21509;
  assign n21511 = n34985 & ~n20715;
  assign n21512 = ~n20700 & n21511;
  assign n21513 = n34985 & n21509;
  assign n21514 = ~n20986 & n21512;
  assign n21515 = ~n21510 & ~n35092;
  assign n21516 = n3473 & ~n21490;
  assign n21517 = ~n21505 & n21516;
  assign n21518 = n3473 & n21506;
  assign n21519 = ~n21515 & ~n35093;
  assign n21520 = ~n21507 & ~n21519;
  assign n21521 = ~n3140 & ~n21520;
  assign n21522 = n3140 & ~n21507;
  assign n21523 = ~n21519 & n21522;
  assign n21524 = ~n34986 & ~n20721;
  assign n21525 = ~n20721 & ~n20986;
  assign n21526 = ~n34986 & n21525;
  assign n21527 = ~n20986 & n21524;
  assign n21528 = n20277 & ~n35094;
  assign n21529 = n20720 & n21525;
  assign n21530 = n20277 & ~n34986;
  assign n21531 = ~n20721 & n21530;
  assign n21532 = ~n20986 & n21531;
  assign n21533 = ~n20277 & ~n35094;
  assign n21534 = ~n21532 & ~n21533;
  assign n21535 = ~n21528 & ~n21529;
  assign n21536 = ~n21523 & ~n35095;
  assign n21537 = ~n21521 & ~n21536;
  assign n21538 = ~n2855 & ~n21537;
  assign n21539 = n2855 & ~n21521;
  assign n21540 = ~n21536 & n21539;
  assign n21541 = n2855 & n21537;
  assign n21542 = ~n20723 & ~n20726;
  assign n21543 = ~n20726 & ~n20986;
  assign n21544 = ~n20723 & n21543;
  assign n21545 = ~n20986 & n21542;
  assign n21546 = n20269 & ~n35097;
  assign n21547 = n20724 & n21543;
  assign n21548 = n20269 & ~n20726;
  assign n21549 = ~n20723 & n21548;
  assign n21550 = ~n20986 & n21549;
  assign n21551 = ~n20269 & ~n35097;
  assign n21552 = ~n21550 & ~n21551;
  assign n21553 = ~n21546 & ~n21547;
  assign n21554 = ~n35096 & ~n35098;
  assign n21555 = ~n21538 & ~n21554;
  assign n21556 = ~n2556 & ~n21555;
  assign n21557 = n2556 & ~n21538;
  assign n21558 = ~n21554 & n21557;
  assign n21559 = ~n34987 & ~n20732;
  assign n21560 = ~n20732 & ~n20986;
  assign n21561 = ~n34987 & n21560;
  assign n21562 = ~n20986 & n21559;
  assign n21563 = n20261 & ~n35099;
  assign n21564 = n20731 & n21560;
  assign n21565 = n20261 & ~n34987;
  assign n21566 = ~n20732 & n21565;
  assign n21567 = ~n20986 & n21566;
  assign n21568 = ~n20261 & ~n35099;
  assign n21569 = ~n21567 & ~n21568;
  assign n21570 = ~n21563 & ~n21564;
  assign n21571 = ~n21558 & ~n35100;
  assign n21572 = ~n21556 & ~n21571;
  assign n21573 = ~n2301 & ~n21572;
  assign n21574 = ~n20734 & ~n20749;
  assign n21575 = ~n20986 & n21574;
  assign n21576 = ~n34989 & ~n21575;
  assign n21577 = n34989 & ~n20749;
  assign n21578 = ~n20734 & n21577;
  assign n21579 = n34989 & n21575;
  assign n21580 = ~n20986 & n21578;
  assign n21581 = ~n21576 & ~n35101;
  assign n21582 = n2301 & ~n21556;
  assign n21583 = ~n21571 & n21582;
  assign n21584 = n2301 & n21572;
  assign n21585 = ~n21581 & ~n35102;
  assign n21586 = ~n21573 & ~n21585;
  assign n21587 = ~n2038 & ~n21586;
  assign n21588 = n2038 & ~n21573;
  assign n21589 = ~n21585 & n21588;
  assign n21590 = ~n34990 & ~n20755;
  assign n21591 = ~n20755 & ~n20986;
  assign n21592 = ~n34990 & n21591;
  assign n21593 = ~n20986 & n21590;
  assign n21594 = n20253 & ~n35103;
  assign n21595 = n20754 & n21591;
  assign n21596 = n20253 & ~n34990;
  assign n21597 = ~n20755 & n21596;
  assign n21598 = ~n20986 & n21597;
  assign n21599 = ~n20253 & ~n35103;
  assign n21600 = ~n21598 & ~n21599;
  assign n21601 = ~n21594 & ~n21595;
  assign n21602 = ~n21589 & ~n35104;
  assign n21603 = ~n21587 & ~n21602;
  assign n21604 = ~n1812 & ~n21603;
  assign n21605 = n1812 & ~n21587;
  assign n21606 = ~n21602 & n21605;
  assign n21607 = n1812 & n21603;
  assign n21608 = ~n20757 & ~n20760;
  assign n21609 = ~n20760 & ~n20986;
  assign n21610 = ~n20757 & n21609;
  assign n21611 = ~n20986 & n21608;
  assign n21612 = n20245 & ~n35106;
  assign n21613 = n20758 & n21609;
  assign n21614 = n20245 & ~n20760;
  assign n21615 = ~n20757 & n21614;
  assign n21616 = ~n20986 & n21615;
  assign n21617 = ~n20245 & ~n35106;
  assign n21618 = ~n21616 & ~n21617;
  assign n21619 = ~n21612 & ~n21613;
  assign n21620 = ~n35105 & ~n35107;
  assign n21621 = ~n21604 & ~n21620;
  assign n21622 = ~n1582 & ~n21621;
  assign n21623 = n1582 & ~n21604;
  assign n21624 = ~n21620 & n21623;
  assign n21625 = ~n34991 & ~n20776;
  assign n21626 = ~n20986 & n21625;
  assign n21627 = ~n34992 & n21626;
  assign n21628 = n34992 & ~n21626;
  assign n21629 = ~n34991 & n34992;
  assign n21630 = ~n20776 & n21629;
  assign n21631 = ~n20986 & n21630;
  assign n21632 = ~n34992 & ~n21626;
  assign n21633 = ~n21631 & ~n21632;
  assign n21634 = ~n21627 & ~n21628;
  assign n21635 = ~n21624 & ~n35108;
  assign n21636 = ~n21622 & ~n21635;
  assign n21637 = ~n1388 & ~n21636;
  assign n21638 = n1388 & ~n21622;
  assign n21639 = ~n21635 & n21638;
  assign n21640 = n1388 & n21636;
  assign n21641 = ~n20778 & ~n20780;
  assign n21642 = ~n20986 & n21641;
  assign n21643 = ~n34993 & ~n21642;
  assign n21644 = ~n20778 & n34993;
  assign n21645 = ~n20780 & n21644;
  assign n21646 = n34993 & n21642;
  assign n21647 = ~n20986 & n21645;
  assign n21648 = ~n21643 & ~n35110;
  assign n21649 = ~n35109 & ~n21648;
  assign n21650 = ~n21637 & ~n21649;
  assign n21651 = ~n1192 & ~n21650;
  assign n21652 = n1192 & ~n21637;
  assign n21653 = ~n21649 & n21652;
  assign n21654 = ~n35019 & ~n21653;
  assign n21655 = ~n21651 & ~n21654;
  assign n21656 = ~n1028 & ~n21655;
  assign n21657 = ~n20799 & ~n20801;
  assign n21658 = ~n20986 & n21657;
  assign n21659 = ~n34996 & ~n21658;
  assign n21660 = ~n20799 & n34996;
  assign n21661 = ~n20801 & n21660;
  assign n21662 = n34996 & n21658;
  assign n21663 = ~n20986 & n21661;
  assign n21664 = ~n21659 & ~n35111;
  assign n21665 = n1028 & ~n21651;
  assign n21666 = ~n21654 & n21665;
  assign n21667 = n1028 & n21655;
  assign n21668 = ~n21664 & ~n35112;
  assign n21669 = ~n21656 & ~n21668;
  assign n21670 = ~n866 & ~n21669;
  assign n21671 = n866 & ~n21656;
  assign n21672 = ~n21668 & n21671;
  assign n21673 = ~n20816 & ~n34998;
  assign n21674 = ~n20816 & ~n20986;
  assign n21675 = ~n34998 & n21674;
  assign n21676 = ~n20986 & n21673;
  assign n21677 = n20824 & ~n35113;
  assign n21678 = n20828 & n21674;
  assign n21679 = n20824 & ~n34998;
  assign n21680 = ~n20816 & n21679;
  assign n21681 = ~n20986 & n21680;
  assign n21682 = ~n20824 & ~n35113;
  assign n21683 = ~n21681 & ~n21682;
  assign n21684 = ~n21677 & ~n21678;
  assign n21685 = ~n21672 & ~n35114;
  assign n21686 = ~n21670 & ~n21685;
  assign n21687 = ~n730 & ~n21686;
  assign n21688 = ~n20830 & ~n20832;
  assign n21689 = ~n20986 & n21688;
  assign n21690 = ~n35000 & ~n21689;
  assign n21691 = ~n20830 & n35000;
  assign n21692 = ~n20832 & n21691;
  assign n21693 = n35000 & n21689;
  assign n21694 = ~n20986 & n21692;
  assign n21695 = ~n21690 & ~n35115;
  assign n21696 = n730 & ~n21670;
  assign n21697 = ~n21685 & n21696;
  assign n21698 = n730 & n21686;
  assign n21699 = ~n21695 & ~n35116;
  assign n21700 = ~n21687 & ~n21699;
  assign n21701 = ~n602 & ~n21700;
  assign n21702 = n602 & ~n21687;
  assign n21703 = ~n21699 & n21702;
  assign n21704 = ~n20847 & ~n35002;
  assign n21705 = ~n20847 & ~n20986;
  assign n21706 = ~n35002 & n21705;
  assign n21707 = ~n20986 & n21704;
  assign n21708 = n20855 & ~n35117;
  assign n21709 = n20859 & n21705;
  assign n21710 = n20855 & ~n35002;
  assign n21711 = ~n20847 & n21710;
  assign n21712 = ~n20986 & n21711;
  assign n21713 = ~n20855 & ~n35117;
  assign n21714 = ~n21712 & ~n21713;
  assign n21715 = ~n21708 & ~n21709;
  assign n21716 = ~n21703 & ~n35118;
  assign n21717 = ~n21701 & ~n21716;
  assign n21718 = ~n497 & ~n21717;
  assign n21719 = n497 & ~n21701;
  assign n21720 = ~n21716 & n21719;
  assign n21721 = n497 & n21717;
  assign n21722 = ~n20861 & ~n20871;
  assign n21723 = ~n20861 & ~n20986;
  assign n21724 = ~n20871 & n21723;
  assign n21725 = ~n20986 & n21722;
  assign n21726 = n20869 & ~n35120;
  assign n21727 = n20872 & n21723;
  assign n21728 = ~n20861 & n20869;
  assign n21729 = ~n20871 & n21728;
  assign n21730 = ~n20986 & n21729;
  assign n21731 = ~n20869 & ~n35120;
  assign n21732 = ~n21730 & ~n21731;
  assign n21733 = ~n21726 & ~n21727;
  assign n21734 = ~n35119 & ~n35121;
  assign n21735 = ~n21718 & ~n21734;
  assign n21736 = ~n403 & ~n21735;
  assign n21737 = n403 & ~n21718;
  assign n21738 = ~n21734 & n21737;
  assign n21739 = ~n20874 & ~n35005;
  assign n21740 = ~n20874 & ~n20986;
  assign n21741 = ~n35005 & n21740;
  assign n21742 = ~n20986 & n21739;
  assign n21743 = n20882 & ~n35122;
  assign n21744 = n20886 & n21740;
  assign n21745 = n20882 & ~n35005;
  assign n21746 = ~n20874 & n21745;
  assign n21747 = ~n20986 & n21746;
  assign n21748 = ~n20882 & ~n35122;
  assign n21749 = ~n21747 & ~n21748;
  assign n21750 = ~n21743 & ~n21744;
  assign n21751 = ~n21738 & ~n35123;
  assign n21752 = ~n21736 & ~n21751;
  assign n21753 = ~n330 & ~n21752;
  assign n21754 = ~n20888 & ~n20890;
  assign n21755 = ~n20986 & n21754;
  assign n21756 = ~n35007 & ~n21755;
  assign n21757 = ~n20888 & n35007;
  assign n21758 = ~n20890 & n21757;
  assign n21759 = n35007 & n21755;
  assign n21760 = ~n20986 & n21758;
  assign n21761 = ~n21756 & ~n35124;
  assign n21762 = n330 & ~n21736;
  assign n21763 = ~n21751 & n21762;
  assign n21764 = n330 & n21752;
  assign n21765 = ~n21761 & ~n35125;
  assign n21766 = ~n21753 & ~n21765;
  assign n21767 = ~n271 & ~n21766;
  assign n21768 = n271 & ~n21753;
  assign n21769 = ~n21765 & n21768;
  assign n21770 = ~n20905 & ~n35009;
  assign n21771 = ~n20905 & ~n20986;
  assign n21772 = ~n35009 & n21771;
  assign n21773 = ~n20986 & n21770;
  assign n21774 = n20913 & ~n35126;
  assign n21775 = n20917 & n21771;
  assign n21776 = n20913 & ~n35009;
  assign n21777 = ~n20905 & n21776;
  assign n21778 = ~n20986 & n21777;
  assign n21779 = ~n20913 & ~n35126;
  assign n21780 = ~n21778 & ~n21779;
  assign n21781 = ~n21774 & ~n21775;
  assign n21782 = ~n21769 & ~n35127;
  assign n21783 = ~n21767 & ~n21782;
  assign n21784 = ~n217 & ~n21783;
  assign n21785 = n217 & ~n21767;
  assign n21786 = ~n21782 & n21785;
  assign n21787 = n217 & n21783;
  assign n21788 = ~n20919 & ~n20929;
  assign n21789 = ~n20919 & ~n20986;
  assign n21790 = ~n20929 & n21789;
  assign n21791 = ~n20986 & n21788;
  assign n21792 = n20927 & ~n35129;
  assign n21793 = n20930 & n21789;
  assign n21794 = ~n20919 & n20927;
  assign n21795 = ~n20929 & n21794;
  assign n21796 = ~n20986 & n21795;
  assign n21797 = ~n20927 & ~n35129;
  assign n21798 = ~n21796 & ~n21797;
  assign n21799 = ~n21792 & ~n21793;
  assign n21800 = ~n35128 & ~n35130;
  assign n21801 = ~n21784 & ~n21800;
  assign n21802 = ~n198 & ~n21801;
  assign n21803 = n198 & ~n21784;
  assign n21804 = ~n21800 & n21803;
  assign n21805 = ~n20932 & ~n35012;
  assign n21806 = ~n20932 & ~n20986;
  assign n21807 = ~n35012 & n21806;
  assign n21808 = ~n20986 & n21805;
  assign n21809 = n20940 & ~n35131;
  assign n21810 = n20944 & n21806;
  assign n21811 = n20940 & ~n35012;
  assign n21812 = ~n20932 & n21811;
  assign n21813 = ~n20986 & n21812;
  assign n21814 = ~n20940 & ~n35131;
  assign n21815 = ~n21813 & ~n21814;
  assign n21816 = ~n21809 & ~n21810;
  assign n21817 = ~n21804 & ~n35132;
  assign n21818 = ~n21802 & ~n21817;
  assign n21819 = ~n20946 & ~n20948;
  assign n21820 = ~n20986 & n21819;
  assign n21821 = ~n35014 & ~n21820;
  assign n21822 = ~n20946 & n35014;
  assign n21823 = ~n20948 & n21822;
  assign n21824 = n35014 & n21820;
  assign n21825 = ~n20986 & n21823;
  assign n21826 = ~n21821 & ~n35133;
  assign n21827 = ~n20962 & ~n20970;
  assign n21828 = ~n20970 & ~n20986;
  assign n21829 = ~n20962 & n21828;
  assign n21830 = ~n20986 & n21827;
  assign n21831 = ~n35017 & ~n35134;
  assign n21832 = ~n21826 & n21831;
  assign n21833 = ~n21818 & n21832;
  assign n21834 = n193 & ~n21833;
  assign n21835 = ~n21802 & n21826;
  assign n21836 = ~n21817 & n21835;
  assign n21837 = n21818 & n21826;
  assign n21838 = n20962 & ~n21828;
  assign n21839 = ~n193 & ~n21827;
  assign n21840 = ~n21838 & n21839;
  assign n21841 = ~n35135 & ~n21840;
  assign n21842 = ~n21834 & n21841;
  assign n21843 = ~n21651 & ~n21653;
  assign n21844 = ~n21842 & n21843;
  assign n21845 = ~n35019 & ~n21844;
  assign n21846 = n35019 & ~n21653;
  assign n21847 = ~n21651 & n21846;
  assign n21848 = n35019 & n21844;
  assign n21849 = ~n21842 & n21847;
  assign n21850 = ~n21845 & ~n35136;
  assign n21851 = ~n21622 & ~n21624;
  assign n21852 = ~n21842 & n21851;
  assign n21853 = ~n35108 & ~n21852;
  assign n21854 = ~n21624 & n35108;
  assign n21855 = ~n21622 & n21854;
  assign n21856 = n35108 & n21852;
  assign n21857 = ~n21842 & n21855;
  assign n21858 = ~n21853 & ~n35137;
  assign n21859 = ~n21604 & ~n35105;
  assign n21860 = ~n21842 & n21859;
  assign n21861 = ~n35107 & ~n21860;
  assign n21862 = ~n21604 & n35107;
  assign n21863 = ~n35105 & n21862;
  assign n21864 = n35107 & n21860;
  assign n21865 = ~n21842 & n21863;
  assign n21866 = ~n21861 & ~n35138;
  assign n21867 = ~n21587 & ~n21589;
  assign n21868 = ~n21842 & n21867;
  assign n21869 = ~n35104 & ~n21868;
  assign n21870 = ~n21589 & n35104;
  assign n21871 = ~n21587 & n21870;
  assign n21872 = n35104 & n21868;
  assign n21873 = ~n21842 & n21871;
  assign n21874 = ~n21869 & ~n35139;
  assign n21875 = ~n21556 & ~n21558;
  assign n21876 = ~n21842 & n21875;
  assign n21877 = ~n35100 & ~n21876;
  assign n21878 = ~n21558 & n35100;
  assign n21879 = ~n21556 & n21878;
  assign n21880 = n35100 & n21876;
  assign n21881 = ~n21842 & n21879;
  assign n21882 = ~n21877 & ~n35140;
  assign n21883 = ~n21538 & ~n35096;
  assign n21884 = ~n21842 & n21883;
  assign n21885 = ~n35098 & ~n21884;
  assign n21886 = ~n21538 & n35098;
  assign n21887 = ~n35096 & n21886;
  assign n21888 = n35098 & n21884;
  assign n21889 = ~n21842 & n21887;
  assign n21890 = ~n21885 & ~n35141;
  assign n21891 = ~n21521 & ~n21523;
  assign n21892 = ~n21842 & n21891;
  assign n21893 = ~n35095 & ~n21892;
  assign n21894 = ~n21523 & n35095;
  assign n21895 = ~n21521 & n21894;
  assign n21896 = n35095 & n21892;
  assign n21897 = ~n21842 & n21895;
  assign n21898 = ~n21893 & ~n35142;
  assign n21899 = ~n21490 & ~n21492;
  assign n21900 = ~n21842 & n21899;
  assign n21901 = ~n35091 & ~n21900;
  assign n21902 = ~n21492 & n35091;
  assign n21903 = ~n21490 & n21902;
  assign n21904 = n35091 & n21900;
  assign n21905 = ~n21842 & n21903;
  assign n21906 = ~n21901 & ~n35143;
  assign n21907 = ~n21472 & ~n35087;
  assign n21908 = ~n21842 & n21907;
  assign n21909 = ~n35089 & ~n21908;
  assign n21910 = ~n21472 & n35089;
  assign n21911 = ~n35087 & n21910;
  assign n21912 = n35089 & n21908;
  assign n21913 = ~n21842 & n21911;
  assign n21914 = ~n21909 & ~n35144;
  assign n21915 = ~n21455 & ~n21457;
  assign n21916 = ~n21842 & n21915;
  assign n21917 = ~n35086 & ~n21916;
  assign n21918 = ~n21457 & n35086;
  assign n21919 = ~n21455 & n21918;
  assign n21920 = n35086 & n21916;
  assign n21921 = ~n21842 & n21919;
  assign n21922 = ~n21917 & ~n35145;
  assign n21923 = ~n21424 & ~n21426;
  assign n21924 = ~n21842 & n21923;
  assign n21925 = ~n35082 & ~n21924;
  assign n21926 = ~n21426 & n35082;
  assign n21927 = ~n21424 & n21926;
  assign n21928 = n35082 & n21924;
  assign n21929 = ~n21842 & n21927;
  assign n21930 = ~n21925 & ~n35146;
  assign n21931 = ~n21406 & ~n35078;
  assign n21932 = ~n21842 & n21931;
  assign n21933 = ~n35080 & ~n21932;
  assign n21934 = ~n21406 & n35080;
  assign n21935 = ~n35078 & n21934;
  assign n21936 = n35080 & n21932;
  assign n21937 = ~n21842 & n21935;
  assign n21938 = ~n21933 & ~n35147;
  assign n21939 = ~n21389 & ~n21391;
  assign n21940 = ~n21842 & n21939;
  assign n21941 = ~n35077 & ~n21940;
  assign n21942 = ~n21391 & n35077;
  assign n21943 = ~n21389 & n21942;
  assign n21944 = n35077 & n21940;
  assign n21945 = ~n21842 & n21943;
  assign n21946 = ~n21941 & ~n35148;
  assign n21947 = ~n21358 & ~n21360;
  assign n21948 = ~n21842 & n21947;
  assign n21949 = ~n35073 & ~n21948;
  assign n21950 = ~n21360 & n35073;
  assign n21951 = ~n21358 & n21950;
  assign n21952 = n35073 & n21948;
  assign n21953 = ~n21842 & n21951;
  assign n21954 = ~n21949 & ~n35149;
  assign n21955 = ~n21339 & ~n35068;
  assign n21956 = ~n21842 & n21955;
  assign n21957 = ~n35071 & ~n21956;
  assign n21958 = ~n21339 & n35071;
  assign n21959 = ~n35068 & n21958;
  assign n21960 = n35071 & n21956;
  assign n21961 = ~n21842 & n21959;
  assign n21962 = ~n21957 & ~n35150;
  assign n21963 = ~n21322 & ~n21324;
  assign n21964 = ~n21842 & n21963;
  assign n21965 = ~n35067 & ~n21964;
  assign n21966 = ~n21324 & n35067;
  assign n21967 = ~n21322 & n21966;
  assign n21968 = n35067 & n21964;
  assign n21969 = ~n21842 & n21967;
  assign n21970 = ~n21965 & ~n35151;
  assign n21971 = ~n21288 & ~n21290;
  assign n21972 = ~n21842 & n21971;
  assign n21973 = ~n35062 & ~n21972;
  assign n21974 = ~n21290 & n35062;
  assign n21975 = ~n21288 & n21974;
  assign n21976 = n35062 & n21972;
  assign n21977 = ~n21842 & n21975;
  assign n21978 = ~n21973 & ~n35152;
  assign n21979 = ~n21252 & ~n21254;
  assign n21980 = ~n21842 & n21979;
  assign n21981 = ~n35056 & ~n21980;
  assign n21982 = ~n21254 & n35056;
  assign n21983 = ~n21252 & n21982;
  assign n21984 = n35056 & n21980;
  assign n21985 = ~n21842 & n21983;
  assign n21986 = ~n21981 & ~n35153;
  assign n21987 = ~n21221 & ~n21223;
  assign n21988 = ~n21842 & n21987;
  assign n21989 = ~n35052 & ~n21988;
  assign n21990 = ~n21223 & n35052;
  assign n21991 = ~n21221 & n21990;
  assign n21992 = n35052 & n21988;
  assign n21993 = ~n21842 & n21991;
  assign n21994 = ~n21989 & ~n35154;
  assign n21995 = ~n21185 & ~n21187;
  assign n21996 = ~n21842 & n21995;
  assign n21997 = ~n35046 & ~n21996;
  assign n21998 = ~n21187 & n35046;
  assign n21999 = ~n21185 & n21998;
  assign n22000 = n35046 & n21996;
  assign n22001 = ~n21842 & n21999;
  assign n22002 = ~n21997 & ~n35155;
  assign n22003 = ~n21151 & ~n21153;
  assign n22004 = ~n21842 & n22003;
  assign n22005 = ~n35041 & ~n22004;
  assign n22006 = ~n21153 & n35041;
  assign n22007 = ~n21151 & n22006;
  assign n22008 = n35041 & n22004;
  assign n22009 = ~n21842 & n22007;
  assign n22010 = ~n22005 & ~n35156;
  assign n22011 = ~n21117 & ~n21119;
  assign n22012 = ~n21842 & n22011;
  assign n22013 = ~n35036 & ~n22012;
  assign n22014 = ~n21119 & n35036;
  assign n22015 = ~n21117 & n22014;
  assign n22016 = n35036 & n22012;
  assign n22017 = ~n21842 & n22015;
  assign n22018 = ~n22013 & ~n35157;
  assign n22019 = ~n21084 & ~n21086;
  assign n22020 = ~n21842 & n22019;
  assign n22021 = ~n35032 & ~n22020;
  assign n22022 = ~n21086 & n35032;
  assign n22023 = ~n21084 & n22022;
  assign n22024 = n35032 & n22020;
  assign n22025 = ~n21842 & n22023;
  assign n22026 = ~n22021 & ~n35158;
  assign n22027 = ~n21050 & ~n21052;
  assign n22028 = ~n21842 & n22027;
  assign n22029 = ~n35027 & ~n22028;
  assign n22030 = ~n21052 & n35027;
  assign n22031 = ~n21050 & n22030;
  assign n22032 = n35027 & n22028;
  assign n22033 = ~n21842 & n22031;
  assign n22034 = ~n22029 & ~n35159;
  assign n22035 = ~n21023 & ~n21025;
  assign n22036 = ~n21842 & n22035;
  assign n22037 = ~n21034 & ~n22036;
  assign n22038 = ~n21025 & n21034;
  assign n22039 = ~n21023 & n22038;
  assign n22040 = n21034 & n22036;
  assign n22041 = ~n21842 & n22039;
  assign n22042 = ~n22037 & ~n35160;
  assign n22043 = ~pi22  & ~n21842;
  assign n22044 = ~pi23  & n22043;
  assign n22045 = n21000 & ~n21842;
  assign n22046 = ~n20986 & ~n21840;
  assign n22047 = ~n35135 & n22046;
  assign n22048 = ~n21834 & n22047;
  assign n22049 = ~n35161 & ~n22048;
  assign n22050 = pi24  & ~n22049;
  assign n22051 = ~pi24  & ~n22048;
  assign n22052 = ~pi24  & n22049;
  assign n22053 = ~n35161 & n22051;
  assign n22054 = ~n22050 & ~n35162;
  assign n22055 = pi22  & ~n21842;
  assign n22056 = ~pi20  & ~pi21 ;
  assign n22057 = ~pi22  & n22056;
  assign n22058 = ~n20210 & ~n35021;
  assign n22059 = ~n20211 & n22058;
  assign n22060 = ~n20227 & n22059;
  assign n22061 = ~n34922 & n22060;
  assign n22062 = n34920 & n20229;
  assign n22063 = ~n20221 & n22061;
  assign n22064 = ~n22057 & ~n35163;
  assign n22065 = ~n20984 & n22064;
  assign n22066 = ~n35017 & n22065;
  assign n22067 = ~n20978 & n22066;
  assign n22068 = ~n22055 & ~n22057;
  assign n22069 = n20986 & n22068;
  assign n22070 = ~n22055 & n22067;
  assign n22071 = pi23  & ~n22043;
  assign n22072 = ~n35161 & ~n22071;
  assign n22073 = ~n35164 & n22072;
  assign n22074 = ~n20986 & ~n22068;
  assign n22075 = n20229 & ~n22074;
  assign n22076 = ~n22073 & ~n22074;
  assign n22077 = n20229 & n22076;
  assign n22078 = ~n22073 & n22075;
  assign n22079 = ~n22054 & ~n35165;
  assign n22080 = ~n20229 & ~n22076;
  assign n22081 = n19401 & ~n22080;
  assign n22082 = ~n22079 & n22081;
  assign n22083 = ~n21003 & ~n35022;
  assign n22084 = ~n21842 & n22083;
  assign n22085 = n21008 & ~n22084;
  assign n22086 = ~n21008 & n22083;
  assign n22087 = ~n21008 & n22084;
  assign n22088 = ~n21842 & n22086;
  assign n22089 = ~n22085 & ~n35166;
  assign n22090 = ~n22082 & ~n22089;
  assign n22091 = ~n22079 & ~n22080;
  assign n22092 = ~n19401 & ~n22091;
  assign n22093 = n18676 & ~n22092;
  assign n22094 = ~n22090 & ~n22092;
  assign n22095 = n18676 & n22094;
  assign n22096 = ~n22090 & n22093;
  assign n22097 = ~n22042 & ~n35167;
  assign n22098 = ~n18676 & ~n22094;
  assign n22099 = n17885 & ~n22098;
  assign n22100 = ~n22097 & n22099;
  assign n22101 = ~n21037 & ~n35024;
  assign n22102 = ~n21842 & n22101;
  assign n22103 = n21047 & ~n22102;
  assign n22104 = ~n21047 & n22102;
  assign n22105 = ~n21037 & n21047;
  assign n22106 = ~n35024 & n22105;
  assign n22107 = n21047 & n22102;
  assign n22108 = ~n21842 & n22106;
  assign n22109 = ~n21047 & ~n22102;
  assign n22110 = ~n35168 & ~n22109;
  assign n22111 = ~n22103 & ~n22104;
  assign n22112 = ~n22100 & ~n35169;
  assign n22113 = ~n22097 & ~n22098;
  assign n22114 = ~n17885 & ~n22113;
  assign n22115 = n17187 & ~n22114;
  assign n22116 = ~n22112 & ~n22114;
  assign n22117 = n17187 & n22116;
  assign n22118 = ~n22112 & n22115;
  assign n22119 = ~n22034 & ~n35170;
  assign n22120 = ~n17187 & ~n22116;
  assign n22121 = n16428 & ~n22120;
  assign n22122 = ~n22119 & n22121;
  assign n22123 = ~n21067 & ~n35028;
  assign n22124 = ~n21842 & n22123;
  assign n22125 = ~n35030 & n22124;
  assign n22126 = n35030 & ~n22124;
  assign n22127 = ~n21067 & n35030;
  assign n22128 = ~n35028 & n22127;
  assign n22129 = ~n21842 & n22128;
  assign n22130 = ~n35030 & ~n22124;
  assign n22131 = ~n22129 & ~n22130;
  assign n22132 = ~n22125 & ~n22126;
  assign n22133 = ~n22122 & ~n35171;
  assign n22134 = ~n22119 & ~n22120;
  assign n22135 = ~n16428 & ~n22134;
  assign n22136 = n15760 & ~n22135;
  assign n22137 = ~n22133 & ~n22135;
  assign n22138 = n15760 & n22137;
  assign n22139 = ~n22133 & n22136;
  assign n22140 = ~n22026 & ~n35172;
  assign n22141 = ~n15760 & ~n22137;
  assign n22142 = n15033 & ~n22141;
  assign n22143 = ~n22140 & n22142;
  assign n22144 = ~n21101 & ~n35033;
  assign n22145 = ~n21842 & n22144;
  assign n22146 = ~n35034 & ~n22145;
  assign n22147 = ~n21101 & n35034;
  assign n22148 = ~n35033 & n22147;
  assign n22149 = n35034 & n22145;
  assign n22150 = ~n21842 & n22148;
  assign n22151 = n35034 & ~n22145;
  assign n22152 = ~n35034 & n22145;
  assign n22153 = ~n22151 & ~n22152;
  assign n22154 = ~n22146 & ~n35173;
  assign n22155 = ~n22143 & n35174;
  assign n22156 = ~n22140 & ~n22141;
  assign n22157 = ~n15033 & ~n22156;
  assign n22158 = n14394 & ~n22157;
  assign n22159 = ~n22155 & ~n22157;
  assign n22160 = n14394 & n22159;
  assign n22161 = ~n22155 & n22158;
  assign n22162 = ~n22018 & ~n35175;
  assign n22163 = ~n14394 & ~n22159;
  assign n22164 = n13704 & ~n22163;
  assign n22165 = ~n22162 & n22164;
  assign n22166 = ~n21134 & ~n35037;
  assign n22167 = ~n21842 & n22166;
  assign n22168 = n35039 & ~n22167;
  assign n22169 = ~n21134 & ~n35039;
  assign n22170 = ~n35037 & n22169;
  assign n22171 = ~n35039 & n22167;
  assign n22172 = ~n21842 & n22170;
  assign n22173 = n35039 & n22167;
  assign n22174 = ~n35039 & ~n22167;
  assign n22175 = ~n22173 & ~n22174;
  assign n22176 = ~n22168 & ~n35176;
  assign n22177 = ~n22165 & n35177;
  assign n22178 = ~n22162 & ~n22163;
  assign n22179 = ~n13704 & ~n22178;
  assign n22180 = n13099 & ~n22179;
  assign n22181 = ~n22177 & ~n22179;
  assign n22182 = n13099 & n22181;
  assign n22183 = ~n22177 & n22180;
  assign n22184 = ~n22010 & ~n35178;
  assign n22185 = ~n13099 & ~n22181;
  assign n22186 = n12442 & ~n22185;
  assign n22187 = ~n22184 & n22186;
  assign n22188 = ~n21168 & ~n35042;
  assign n22189 = ~n21168 & ~n21842;
  assign n22190 = ~n35042 & n22189;
  assign n22191 = ~n21842 & n22188;
  assign n22192 = ~n35044 & ~n35179;
  assign n22193 = n21183 & n22189;
  assign n22194 = n35044 & n35179;
  assign n22195 = ~n21168 & ~n35044;
  assign n22196 = ~n35042 & n22195;
  assign n22197 = ~n21842 & n22196;
  assign n22198 = n35044 & ~n35179;
  assign n22199 = ~n22197 & ~n22198;
  assign n22200 = ~n22192 & ~n35180;
  assign n22201 = ~n22187 & ~n35181;
  assign n22202 = ~n22184 & ~n22185;
  assign n22203 = ~n12442 & ~n22202;
  assign n22204 = n11858 & ~n22203;
  assign n22205 = ~n22201 & ~n22203;
  assign n22206 = n11858 & n22205;
  assign n22207 = ~n22201 & n22204;
  assign n22208 = ~n22002 & ~n35182;
  assign n22209 = ~n11858 & ~n22205;
  assign n22210 = n11229 & ~n22209;
  assign n22211 = ~n22208 & n22210;
  assign n22212 = ~n21202 & ~n35047;
  assign n22213 = ~n21842 & n22212;
  assign n22214 = ~n35050 & ~n22213;
  assign n22215 = ~n21202 & n35050;
  assign n22216 = ~n35047 & n22215;
  assign n22217 = n35050 & n22213;
  assign n22218 = ~n21842 & n22216;
  assign n22219 = ~n22214 & ~n35183;
  assign n22220 = ~n22211 & ~n22219;
  assign n22221 = ~n22208 & ~n22209;
  assign n22222 = ~n11229 & ~n22221;
  assign n22223 = n10681 & ~n22222;
  assign n22224 = ~n22220 & ~n22222;
  assign n22225 = n10681 & n22224;
  assign n22226 = ~n22220 & n22223;
  assign n22227 = ~n21994 & ~n35184;
  assign n22228 = ~n10681 & ~n22224;
  assign n22229 = n10086 & ~n22228;
  assign n22230 = ~n22227 & n22229;
  assign n22231 = ~n21238 & ~n35053;
  assign n22232 = ~n21238 & ~n21842;
  assign n22233 = ~n35053 & n22232;
  assign n22234 = ~n21842 & n22231;
  assign n22235 = n21249 & ~n35185;
  assign n22236 = n21250 & n22232;
  assign n22237 = ~n21249 & n35185;
  assign n22238 = ~n21238 & n21249;
  assign n22239 = ~n35053 & n22238;
  assign n22240 = ~n21842 & n22239;
  assign n22241 = ~n21249 & ~n35185;
  assign n22242 = ~n22240 & ~n22241;
  assign n22243 = ~n22235 & ~n35186;
  assign n22244 = ~n22230 & ~n35187;
  assign n22245 = ~n22227 & ~n22228;
  assign n22246 = ~n10086 & ~n22245;
  assign n22247 = n9565 & ~n22246;
  assign n22248 = ~n22244 & ~n22246;
  assign n22249 = n9565 & n22248;
  assign n22250 = ~n22244 & n22247;
  assign n22251 = ~n21986 & ~n35188;
  assign n22252 = ~n9565 & ~n22248;
  assign n22253 = n8998 & ~n22252;
  assign n22254 = ~n22251 & n22253;
  assign n22255 = ~n21269 & ~n35057;
  assign n22256 = ~n21842 & n22255;
  assign n22257 = ~n35060 & n22256;
  assign n22258 = n35060 & ~n22256;
  assign n22259 = ~n21269 & n35060;
  assign n22260 = ~n35057 & n22259;
  assign n22261 = n35060 & n22256;
  assign n22262 = ~n21842 & n22260;
  assign n22263 = ~n35060 & ~n22256;
  assign n22264 = ~n35189 & ~n22263;
  assign n22265 = ~n22257 & ~n22258;
  assign n22266 = ~n22254 & ~n35190;
  assign n22267 = ~n22251 & ~n22252;
  assign n22268 = ~n8998 & ~n22267;
  assign n22269 = n8506 & ~n22268;
  assign n22270 = ~n22266 & ~n22268;
  assign n22271 = n8506 & n22270;
  assign n22272 = ~n22266 & n22269;
  assign n22273 = ~n21978 & ~n35191;
  assign n22274 = ~n8506 & ~n22270;
  assign n22275 = n7975 & ~n22274;
  assign n22276 = ~n22273 & n22275;
  assign n22277 = ~n21305 & ~n35063;
  assign n22278 = ~n21305 & ~n21842;
  assign n22279 = ~n35063 & n22278;
  assign n22280 = ~n21842 & n22277;
  assign n22281 = n35065 & ~n35192;
  assign n22282 = n21320 & n22278;
  assign n22283 = ~n35065 & n35192;
  assign n22284 = ~n21305 & n35065;
  assign n22285 = ~n35063 & n22284;
  assign n22286 = ~n21842 & n22285;
  assign n22287 = ~n35065 & ~n35192;
  assign n22288 = ~n22286 & ~n22287;
  assign n22289 = ~n22281 & ~n35193;
  assign n22290 = ~n22276 & ~n35194;
  assign n22291 = ~n22273 & ~n22274;
  assign n22292 = ~n7975 & ~n22291;
  assign n22293 = n7512 & ~n22292;
  assign n22294 = ~n22290 & ~n22292;
  assign n22295 = n7512 & n22294;
  assign n22296 = ~n22290 & n22293;
  assign n22297 = ~n21970 & ~n35195;
  assign n22298 = ~n7512 & ~n22294;
  assign n22299 = n7015 & ~n22298;
  assign n22300 = ~n22297 & n22299;
  assign n22301 = ~n21962 & ~n22300;
  assign n22302 = ~n22297 & ~n22298;
  assign n22303 = ~n7015 & ~n22302;
  assign n22304 = n6579 & ~n22303;
  assign n22305 = ~n22301 & ~n22303;
  assign n22306 = n6579 & n22305;
  assign n22307 = ~n22301 & n22304;
  assign n22308 = ~n21954 & ~n35196;
  assign n22309 = ~n6579 & ~n22305;
  assign n22310 = n6117 & ~n22309;
  assign n22311 = ~n22308 & n22310;
  assign n22312 = ~n21375 & ~n35075;
  assign n22313 = ~n21375 & ~n21842;
  assign n22314 = ~n35075 & n22313;
  assign n22315 = ~n21842 & n22312;
  assign n22316 = n21383 & ~n35197;
  assign n22317 = n21387 & n22313;
  assign n22318 = ~n21375 & n21383;
  assign n22319 = ~n35075 & n22318;
  assign n22320 = ~n21842 & n22319;
  assign n22321 = ~n21383 & ~n35197;
  assign n22322 = ~n22320 & ~n22321;
  assign n22323 = ~n22316 & ~n22317;
  assign n22324 = ~n22311 & ~n35198;
  assign n22325 = ~n22308 & ~n22309;
  assign n22326 = ~n6117 & ~n22325;
  assign n22327 = n5708 & ~n22326;
  assign n22328 = ~n22324 & ~n22326;
  assign n22329 = n5708 & n22328;
  assign n22330 = ~n22324 & n22327;
  assign n22331 = ~n21946 & ~n35199;
  assign n22332 = ~n5708 & ~n22328;
  assign n22333 = n5278 & ~n22332;
  assign n22334 = ~n22331 & n22333;
  assign n22335 = ~n21938 & ~n22334;
  assign n22336 = ~n22331 & ~n22332;
  assign n22337 = ~n5278 & ~n22336;
  assign n22338 = n4903 & ~n22337;
  assign n22339 = ~n22335 & ~n22337;
  assign n22340 = n4903 & n22339;
  assign n22341 = ~n22335 & n22338;
  assign n22342 = ~n21930 & ~n35200;
  assign n22343 = ~n4903 & ~n22339;
  assign n22344 = n4508 & ~n22343;
  assign n22345 = ~n22342 & n22344;
  assign n22346 = ~n21441 & ~n35084;
  assign n22347 = ~n21441 & ~n21842;
  assign n22348 = ~n35084 & n22347;
  assign n22349 = ~n21842 & n22346;
  assign n22350 = n21449 & ~n35201;
  assign n22351 = n21453 & n22347;
  assign n22352 = ~n21441 & n21449;
  assign n22353 = ~n35084 & n22352;
  assign n22354 = ~n21842 & n22353;
  assign n22355 = ~n21449 & ~n35201;
  assign n22356 = ~n22354 & ~n22355;
  assign n22357 = ~n22350 & ~n22351;
  assign n22358 = ~n22345 & ~n35202;
  assign n22359 = ~n22342 & ~n22343;
  assign n22360 = ~n4508 & ~n22359;
  assign n22361 = n4155 & ~n22360;
  assign n22362 = ~n22358 & ~n22360;
  assign n22363 = n4155 & n22362;
  assign n22364 = ~n22358 & n22361;
  assign n22365 = ~n21922 & ~n35203;
  assign n22366 = ~n4155 & ~n22362;
  assign n22367 = n3788 & ~n22366;
  assign n22368 = ~n22365 & n22367;
  assign n22369 = ~n21914 & ~n22368;
  assign n22370 = ~n22365 & ~n22366;
  assign n22371 = ~n3788 & ~n22370;
  assign n22372 = n3473 & ~n22371;
  assign n22373 = ~n22369 & ~n22371;
  assign n22374 = n3473 & n22373;
  assign n22375 = ~n22369 & n22372;
  assign n22376 = ~n21906 & ~n35204;
  assign n22377 = ~n3473 & ~n22373;
  assign n22378 = n3140 & ~n22377;
  assign n22379 = ~n22376 & n22378;
  assign n22380 = ~n21507 & ~n35093;
  assign n22381 = ~n21507 & ~n21842;
  assign n22382 = ~n35093 & n22381;
  assign n22383 = ~n21842 & n22380;
  assign n22384 = n21515 & ~n35205;
  assign n22385 = n21519 & n22381;
  assign n22386 = ~n21507 & n21515;
  assign n22387 = ~n35093 & n22386;
  assign n22388 = ~n21842 & n22387;
  assign n22389 = ~n21515 & ~n35205;
  assign n22390 = ~n22388 & ~n22389;
  assign n22391 = ~n22384 & ~n22385;
  assign n22392 = ~n22379 & ~n35206;
  assign n22393 = ~n22376 & ~n22377;
  assign n22394 = ~n3140 & ~n22393;
  assign n22395 = n2855 & ~n22394;
  assign n22396 = ~n22392 & ~n22394;
  assign n22397 = n2855 & n22396;
  assign n22398 = ~n22392 & n22395;
  assign n22399 = ~n21898 & ~n35207;
  assign n22400 = ~n2855 & ~n22396;
  assign n22401 = n2556 & ~n22400;
  assign n22402 = ~n22399 & n22401;
  assign n22403 = ~n21890 & ~n22402;
  assign n22404 = ~n22399 & ~n22400;
  assign n22405 = ~n2556 & ~n22404;
  assign n22406 = n2301 & ~n22405;
  assign n22407 = ~n22403 & ~n22405;
  assign n22408 = n2301 & n22407;
  assign n22409 = ~n22403 & n22406;
  assign n22410 = ~n21882 & ~n35208;
  assign n22411 = ~n2301 & ~n22407;
  assign n22412 = n2038 & ~n22411;
  assign n22413 = ~n22410 & n22412;
  assign n22414 = ~n21573 & ~n35102;
  assign n22415 = ~n21573 & ~n21842;
  assign n22416 = ~n35102 & n22415;
  assign n22417 = ~n21842 & n22414;
  assign n22418 = n21581 & ~n35209;
  assign n22419 = n21585 & n22415;
  assign n22420 = ~n21573 & n21581;
  assign n22421 = ~n35102 & n22420;
  assign n22422 = ~n21842 & n22421;
  assign n22423 = ~n21581 & ~n35209;
  assign n22424 = ~n22422 & ~n22423;
  assign n22425 = ~n22418 & ~n22419;
  assign n22426 = ~n22413 & ~n35210;
  assign n22427 = ~n22410 & ~n22411;
  assign n22428 = ~n2038 & ~n22427;
  assign n22429 = n1812 & ~n22428;
  assign n22430 = ~n22426 & ~n22428;
  assign n22431 = n1812 & n22430;
  assign n22432 = ~n22426 & n22429;
  assign n22433 = ~n21874 & ~n35211;
  assign n22434 = ~n1812 & ~n22430;
  assign n22435 = n1582 & ~n22434;
  assign n22436 = ~n22433 & n22435;
  assign n22437 = ~n21866 & ~n22436;
  assign n22438 = ~n22433 & ~n22434;
  assign n22439 = ~n1582 & ~n22438;
  assign n22440 = n1388 & ~n22439;
  assign n22441 = ~n22437 & ~n22439;
  assign n22442 = n1388 & n22441;
  assign n22443 = ~n22437 & n22440;
  assign n22444 = ~n21858 & ~n35212;
  assign n22445 = ~n1388 & ~n22441;
  assign n22446 = ~n22444 & ~n22445;
  assign n22447 = ~n1192 & ~n22446;
  assign n22448 = n1192 & ~n22445;
  assign n22449 = ~n22444 & n22448;
  assign n22450 = ~n21637 & ~n35109;
  assign n22451 = ~n21842 & n22450;
  assign n22452 = n21648 & ~n22451;
  assign n22453 = ~n21648 & n22451;
  assign n22454 = ~n21637 & n21648;
  assign n22455 = ~n35109 & n22454;
  assign n22456 = n21648 & n22451;
  assign n22457 = ~n21842 & n22455;
  assign n22458 = ~n21648 & ~n22451;
  assign n22459 = ~n35213 & ~n22458;
  assign n22460 = ~n22452 & ~n22453;
  assign n22461 = ~n22449 & ~n35214;
  assign n22462 = ~n22447 & ~n22461;
  assign n22463 = ~n1028 & ~n22462;
  assign n22464 = n1028 & ~n22447;
  assign n22465 = n1028 & n22462;
  assign n22466 = ~n22461 & n22464;
  assign n22467 = ~n21850 & ~n35215;
  assign n22468 = ~n22463 & ~n22467;
  assign n22469 = ~n866 & ~n22468;
  assign n22470 = n866 & ~n22463;
  assign n22471 = ~n22467 & n22470;
  assign n22472 = ~n21656 & ~n35112;
  assign n22473 = ~n21656 & ~n21842;
  assign n22474 = ~n35112 & n22473;
  assign n22475 = ~n21842 & n22472;
  assign n22476 = n21664 & ~n35216;
  assign n22477 = n21668 & n22473;
  assign n22478 = ~n21656 & n21664;
  assign n22479 = ~n35112 & n22478;
  assign n22480 = ~n21842 & n22479;
  assign n22481 = ~n21664 & ~n35216;
  assign n22482 = ~n22480 & ~n22481;
  assign n22483 = ~n22476 & ~n22477;
  assign n22484 = ~n22471 & ~n35217;
  assign n22485 = ~n22469 & ~n22484;
  assign n22486 = ~n730 & ~n22485;
  assign n22487 = ~n21670 & ~n21672;
  assign n22488 = ~n21842 & n22487;
  assign n22489 = ~n35114 & ~n22488;
  assign n22490 = ~n21672 & n35114;
  assign n22491 = ~n21670 & n22490;
  assign n22492 = n35114 & n22488;
  assign n22493 = ~n21842 & n22491;
  assign n22494 = ~n22489 & ~n35218;
  assign n22495 = n730 & ~n22469;
  assign n22496 = n730 & n22485;
  assign n22497 = ~n22484 & n22495;
  assign n22498 = ~n22494 & ~n35219;
  assign n22499 = ~n22486 & ~n22498;
  assign n22500 = ~n602 & ~n22499;
  assign n22501 = n602 & ~n22486;
  assign n22502 = ~n22498 & n22501;
  assign n22503 = ~n21687 & ~n35116;
  assign n22504 = ~n21687 & ~n21842;
  assign n22505 = ~n35116 & n22504;
  assign n22506 = ~n21842 & n22503;
  assign n22507 = n21695 & ~n35220;
  assign n22508 = n21699 & n22504;
  assign n22509 = ~n21687 & n21695;
  assign n22510 = ~n35116 & n22509;
  assign n22511 = ~n21842 & n22510;
  assign n22512 = ~n21695 & ~n35220;
  assign n22513 = ~n22511 & ~n22512;
  assign n22514 = ~n22507 & ~n22508;
  assign n22515 = ~n22502 & ~n35221;
  assign n22516 = ~n22500 & ~n22515;
  assign n22517 = ~n497 & ~n22516;
  assign n22518 = ~n21701 & ~n21703;
  assign n22519 = ~n21842 & n22518;
  assign n22520 = ~n35118 & ~n22519;
  assign n22521 = ~n21703 & n35118;
  assign n22522 = ~n21701 & n22521;
  assign n22523 = n35118 & n22519;
  assign n22524 = ~n21842 & n22522;
  assign n22525 = ~n22520 & ~n35222;
  assign n22526 = n497 & ~n22500;
  assign n22527 = n497 & n22516;
  assign n22528 = ~n22515 & n22526;
  assign n22529 = ~n22525 & ~n35223;
  assign n22530 = ~n22517 & ~n22529;
  assign n22531 = ~n403 & ~n22530;
  assign n22532 = ~n21718 & ~n35119;
  assign n22533 = ~n21842 & n22532;
  assign n22534 = ~n35121 & ~n22533;
  assign n22535 = ~n21718 & n35121;
  assign n22536 = ~n35119 & n22535;
  assign n22537 = n35121 & n22533;
  assign n22538 = ~n21842 & n22536;
  assign n22539 = ~n22534 & ~n35224;
  assign n22540 = n403 & ~n22517;
  assign n22541 = ~n22529 & n22540;
  assign n22542 = ~n22539 & ~n22541;
  assign n22543 = ~n22531 & ~n22542;
  assign n22544 = ~n330 & ~n22543;
  assign n22545 = ~n21736 & ~n21738;
  assign n22546 = ~n21842 & n22545;
  assign n22547 = ~n35123 & ~n22546;
  assign n22548 = ~n21738 & n35123;
  assign n22549 = ~n21736 & n22548;
  assign n22550 = n35123 & n22546;
  assign n22551 = ~n21842 & n22549;
  assign n22552 = ~n22547 & ~n35225;
  assign n22553 = n330 & ~n22531;
  assign n22554 = n330 & n22543;
  assign n22555 = ~n22542 & n22553;
  assign n22556 = ~n22552 & ~n35226;
  assign n22557 = ~n22544 & ~n22556;
  assign n22558 = ~n271 & ~n22557;
  assign n22559 = n271 & ~n22544;
  assign n22560 = ~n22556 & n22559;
  assign n22561 = ~n21753 & ~n35125;
  assign n22562 = ~n21753 & ~n21842;
  assign n22563 = ~n35125 & n22562;
  assign n22564 = ~n21842 & n22561;
  assign n22565 = n21761 & ~n35227;
  assign n22566 = n21765 & n22562;
  assign n22567 = ~n21753 & n21761;
  assign n22568 = ~n35125 & n22567;
  assign n22569 = ~n21842 & n22568;
  assign n22570 = ~n21761 & ~n35227;
  assign n22571 = ~n22569 & ~n22570;
  assign n22572 = ~n22565 & ~n22566;
  assign n22573 = ~n22560 & ~n35228;
  assign n22574 = ~n22558 & ~n22573;
  assign n22575 = ~n217 & ~n22574;
  assign n22576 = ~n21767 & ~n21769;
  assign n22577 = ~n21842 & n22576;
  assign n22578 = ~n35127 & ~n22577;
  assign n22579 = ~n21769 & n35127;
  assign n22580 = ~n21767 & n22579;
  assign n22581 = n35127 & n22577;
  assign n22582 = ~n21842 & n22580;
  assign n22583 = ~n22578 & ~n35229;
  assign n22584 = n217 & ~n22558;
  assign n22585 = n217 & n22574;
  assign n22586 = ~n22573 & n22584;
  assign n22587 = ~n22583 & ~n35230;
  assign n22588 = ~n22575 & ~n22587;
  assign n22589 = ~n198 & ~n22588;
  assign n22590 = ~n21784 & ~n35128;
  assign n22591 = ~n21842 & n22590;
  assign n22592 = ~n35130 & ~n22591;
  assign n22593 = ~n21784 & n35130;
  assign n22594 = ~n35128 & n22593;
  assign n22595 = n35130 & n22591;
  assign n22596 = ~n21842 & n22594;
  assign n22597 = ~n22592 & ~n35231;
  assign n22598 = n198 & ~n22575;
  assign n22599 = ~n22587 & n22598;
  assign n22600 = ~n22597 & ~n22599;
  assign n22601 = ~n22589 & ~n22600;
  assign n22602 = ~n21802 & ~n21804;
  assign n22603 = ~n21842 & n22602;
  assign n22604 = ~n35132 & ~n22603;
  assign n22605 = ~n21804 & n35132;
  assign n22606 = ~n21802 & n22605;
  assign n22607 = n35132 & n22603;
  assign n22608 = ~n21842 & n22606;
  assign n22609 = ~n22604 & ~n35232;
  assign n22610 = ~n21818 & ~n21826;
  assign n22611 = ~n21826 & ~n21842;
  assign n22612 = ~n21818 & n22611;
  assign n22613 = ~n21842 & n22610;
  assign n22614 = ~n35135 & ~n35233;
  assign n22615 = ~n22609 & n22614;
  assign n22616 = ~n22601 & n22615;
  assign n22617 = n193 & ~n22616;
  assign n22618 = ~n22589 & n22609;
  assign n22619 = n22601 & n22609;
  assign n22620 = ~n22600 & n22618;
  assign n22621 = n21818 & ~n22611;
  assign n22622 = ~n193 & ~n22610;
  assign n22623 = ~n22621 & n22622;
  assign n22624 = ~n35234 & ~n22623;
  assign n22625 = ~n22617 & n22624;
  assign n22626 = ~n22463 & ~n35215;
  assign n22627 = ~n22463 & ~n22625;
  assign n22628 = ~n35215 & n22627;
  assign n22629 = ~n22625 & n22626;
  assign n22630 = n21850 & ~n35235;
  assign n22631 = n22467 & n22627;
  assign n22632 = n21850 & ~n35215;
  assign n22633 = ~n22463 & n22632;
  assign n22634 = ~n22625 & n22633;
  assign n22635 = ~n21850 & ~n35235;
  assign n22636 = ~n22634 & ~n22635;
  assign n22637 = ~n22630 & ~n22631;
  assign n22638 = pi20  & ~n22625;
  assign n22639 = ~pi18  & ~pi19 ;
  assign n22640 = ~pi20  & n22639;
  assign n22641 = ~n22638 & ~n22640;
  assign n22642 = ~n21842 & ~n22641;
  assign n22643 = ~pi20  & ~n22625;
  assign n22644 = pi21  & ~n22643;
  assign n22645 = ~pi21  & n22643;
  assign n22646 = n22056 & ~n22625;
  assign n22647 = ~n22644 & ~n35237;
  assign n22648 = ~n35015 & ~n35163;
  assign n22649 = ~n20965 & n22648;
  assign n22650 = ~n20984 & n22649;
  assign n22651 = ~n35017 & n22650;
  assign n22652 = n20970 & n20986;
  assign n22653 = ~n20978 & n22651;
  assign n22654 = ~n22640 & ~n35238;
  assign n22655 = ~n21840 & n22654;
  assign n22656 = ~n35135 & n22655;
  assign n22657 = ~n21834 & n22656;
  assign n22658 = n21842 & n22641;
  assign n22659 = ~n22638 & n22657;
  assign n22660 = n22647 & ~n35239;
  assign n22661 = ~n22642 & ~n22660;
  assign n22662 = ~n20986 & ~n22661;
  assign n22663 = n20986 & ~n22642;
  assign n22664 = ~n22660 & n22663;
  assign n22665 = ~n21842 & ~n22623;
  assign n22666 = ~n35234 & n22665;
  assign n22667 = ~n22617 & n22666;
  assign n22668 = ~n35237 & ~n22667;
  assign n22669 = pi22  & ~n22668;
  assign n22670 = ~pi22  & ~n22667;
  assign n22671 = ~pi22  & n22668;
  assign n22672 = ~n35237 & n22670;
  assign n22673 = ~n22669 & ~n35240;
  assign n22674 = ~n22664 & ~n22673;
  assign n22675 = ~n22662 & ~n22674;
  assign n22676 = ~n20229 & ~n22675;
  assign n22677 = n20229 & ~n22662;
  assign n22678 = ~n22674 & n22677;
  assign n22679 = n20229 & n22675;
  assign n22680 = ~n35164 & ~n22074;
  assign n22681 = ~n22625 & n22680;
  assign n22682 = n22072 & ~n22681;
  assign n22683 = ~n22072 & n22680;
  assign n22684 = ~n22072 & n22681;
  assign n22685 = ~n22625 & n22683;
  assign n22686 = ~n22682 & ~n35242;
  assign n22687 = ~n35241 & ~n22686;
  assign n22688 = ~n22676 & ~n22687;
  assign n22689 = ~n19401 & ~n22688;
  assign n22690 = n19401 & ~n22676;
  assign n22691 = ~n22687 & n22690;
  assign n22692 = ~n35165 & ~n22080;
  assign n22693 = ~n22080 & ~n22625;
  assign n22694 = ~n35165 & n22693;
  assign n22695 = ~n22625 & n22692;
  assign n22696 = n22054 & ~n35243;
  assign n22697 = n22079 & n22693;
  assign n22698 = n22054 & ~n35165;
  assign n22699 = ~n22080 & n22698;
  assign n22700 = ~n22625 & n22699;
  assign n22701 = ~n22054 & ~n35243;
  assign n22702 = ~n22700 & ~n22701;
  assign n22703 = ~n22696 & ~n22697;
  assign n22704 = ~n22691 & ~n35244;
  assign n22705 = ~n22689 & ~n22704;
  assign n22706 = ~n18676 & ~n22705;
  assign n22707 = n18676 & ~n22689;
  assign n22708 = ~n22704 & n22707;
  assign n22709 = n18676 & n22705;
  assign n22710 = ~n22082 & ~n22092;
  assign n22711 = ~n22625 & n22710;
  assign n22712 = n22089 & ~n22711;
  assign n22713 = ~n22089 & n22711;
  assign n22714 = n22089 & ~n22092;
  assign n22715 = ~n22082 & n22714;
  assign n22716 = n22089 & n22711;
  assign n22717 = ~n22625 & n22715;
  assign n22718 = ~n22089 & ~n22711;
  assign n22719 = ~n35246 & ~n22718;
  assign n22720 = ~n22712 & ~n22713;
  assign n22721 = ~n35245 & ~n35247;
  assign n22722 = ~n22706 & ~n22721;
  assign n22723 = ~n17885 & ~n22722;
  assign n22724 = n17885 & ~n22706;
  assign n22725 = ~n22721 & n22724;
  assign n22726 = ~n35167 & ~n22098;
  assign n22727 = ~n22098 & ~n22625;
  assign n22728 = ~n35167 & n22727;
  assign n22729 = ~n22625 & n22726;
  assign n22730 = n22042 & ~n35248;
  assign n22731 = n22097 & n22727;
  assign n22732 = n22042 & ~n35167;
  assign n22733 = ~n22098 & n22732;
  assign n22734 = ~n22625 & n22733;
  assign n22735 = ~n22042 & ~n35248;
  assign n22736 = ~n22734 & ~n22735;
  assign n22737 = ~n22730 & ~n22731;
  assign n22738 = ~n22725 & ~n35249;
  assign n22739 = ~n22723 & ~n22738;
  assign n22740 = ~n17187 & ~n22739;
  assign n22741 = n17187 & ~n22723;
  assign n22742 = ~n22738 & n22741;
  assign n22743 = n17187 & n22739;
  assign n22744 = ~n22100 & ~n22114;
  assign n22745 = ~n22625 & n22744;
  assign n22746 = ~n35169 & n22745;
  assign n22747 = n35169 & ~n22745;
  assign n22748 = n35169 & ~n22114;
  assign n22749 = ~n22100 & n22748;
  assign n22750 = ~n22625 & n22749;
  assign n22751 = ~n35169 & ~n22745;
  assign n22752 = ~n22750 & ~n22751;
  assign n22753 = ~n22746 & ~n22747;
  assign n22754 = ~n35250 & ~n35251;
  assign n22755 = ~n22740 & ~n22754;
  assign n22756 = ~n16428 & ~n22755;
  assign n22757 = n16428 & ~n22740;
  assign n22758 = ~n22754 & n22757;
  assign n22759 = ~n35170 & ~n22120;
  assign n22760 = ~n22120 & ~n22625;
  assign n22761 = ~n35170 & n22760;
  assign n22762 = ~n22625 & n22759;
  assign n22763 = n22034 & ~n35252;
  assign n22764 = n22119 & n22760;
  assign n22765 = n22034 & ~n35170;
  assign n22766 = ~n22120 & n22765;
  assign n22767 = ~n22625 & n22766;
  assign n22768 = ~n22034 & ~n35252;
  assign n22769 = ~n22767 & ~n22768;
  assign n22770 = ~n22763 & ~n22764;
  assign n22771 = ~n22758 & ~n35253;
  assign n22772 = ~n22756 & ~n22771;
  assign n22773 = ~n15760 & ~n22772;
  assign n22774 = n15760 & ~n22756;
  assign n22775 = ~n22771 & n22774;
  assign n22776 = n15760 & n22772;
  assign n22777 = ~n22122 & ~n22135;
  assign n22778 = ~n22625 & n22777;
  assign n22779 = ~n35171 & ~n22778;
  assign n22780 = n35171 & ~n22135;
  assign n22781 = ~n22122 & n22780;
  assign n22782 = n35171 & n22778;
  assign n22783 = ~n22625 & n22781;
  assign n22784 = n35171 & ~n22778;
  assign n22785 = ~n35171 & n22778;
  assign n22786 = ~n22784 & ~n22785;
  assign n22787 = ~n22779 & ~n35255;
  assign n22788 = ~n35254 & n35256;
  assign n22789 = ~n22773 & ~n22788;
  assign n22790 = ~n15033 & ~n22789;
  assign n22791 = n15033 & ~n22773;
  assign n22792 = ~n22788 & n22791;
  assign n22793 = ~n35172 & ~n22141;
  assign n22794 = ~n22141 & ~n22625;
  assign n22795 = ~n35172 & n22794;
  assign n22796 = ~n22625 & n22793;
  assign n22797 = n22026 & ~n35257;
  assign n22798 = n22140 & n22794;
  assign n22799 = n22026 & ~n35172;
  assign n22800 = ~n22141 & n22799;
  assign n22801 = ~n22625 & n22800;
  assign n22802 = ~n22026 & ~n35257;
  assign n22803 = ~n22801 & ~n22802;
  assign n22804 = ~n22797 & ~n22798;
  assign n22805 = ~n22792 & ~n35258;
  assign n22806 = ~n22790 & ~n22805;
  assign n22807 = ~n14394 & ~n22806;
  assign n22808 = n14394 & ~n22790;
  assign n22809 = ~n22805 & n22808;
  assign n22810 = n14394 & n22806;
  assign n22811 = ~n22143 & ~n22157;
  assign n22812 = ~n22625 & n22811;
  assign n22813 = n35174 & ~n22812;
  assign n22814 = ~n35174 & ~n22157;
  assign n22815 = ~n22143 & n22814;
  assign n22816 = ~n35174 & n22812;
  assign n22817 = ~n22625 & n22815;
  assign n22818 = n35174 & n22812;
  assign n22819 = ~n35174 & ~n22812;
  assign n22820 = ~n22818 & ~n22819;
  assign n22821 = ~n22813 & ~n35260;
  assign n22822 = ~n35259 & n35261;
  assign n22823 = ~n22807 & ~n22822;
  assign n22824 = ~n13704 & ~n22823;
  assign n22825 = n13704 & ~n22807;
  assign n22826 = ~n22822 & n22825;
  assign n22827 = ~n35175 & ~n22163;
  assign n22828 = ~n22163 & ~n22625;
  assign n22829 = ~n35175 & n22828;
  assign n22830 = ~n22625 & n22827;
  assign n22831 = n22018 & ~n35262;
  assign n22832 = n22162 & n22828;
  assign n22833 = n22018 & ~n35175;
  assign n22834 = ~n22163 & n22833;
  assign n22835 = ~n22625 & n22834;
  assign n22836 = ~n22018 & ~n35262;
  assign n22837 = ~n22835 & ~n22836;
  assign n22838 = ~n22831 & ~n22832;
  assign n22839 = ~n22826 & ~n35263;
  assign n22840 = ~n22824 & ~n22839;
  assign n22841 = ~n13099 & ~n22840;
  assign n22842 = n13099 & ~n22824;
  assign n22843 = ~n22839 & n22842;
  assign n22844 = n13099 & n22840;
  assign n22845 = ~n22165 & ~n22179;
  assign n22846 = ~n22179 & ~n22625;
  assign n22847 = ~n22165 & n22846;
  assign n22848 = ~n22625 & n22845;
  assign n22849 = ~n35177 & ~n35265;
  assign n22850 = n22177 & n22846;
  assign n22851 = n35177 & n35265;
  assign n22852 = ~n35177 & ~n22179;
  assign n22853 = ~n22165 & n22852;
  assign n22854 = ~n22625 & n22853;
  assign n22855 = n35177 & ~n35265;
  assign n22856 = ~n22854 & ~n22855;
  assign n22857 = ~n22849 & ~n35266;
  assign n22858 = ~n35264 & ~n35267;
  assign n22859 = ~n22841 & ~n22858;
  assign n22860 = ~n12442 & ~n22859;
  assign n22861 = n12442 & ~n22841;
  assign n22862 = ~n22858 & n22861;
  assign n22863 = ~n35178 & ~n22185;
  assign n22864 = ~n22185 & ~n22625;
  assign n22865 = ~n35178 & n22864;
  assign n22866 = ~n22625 & n22863;
  assign n22867 = n22010 & ~n35268;
  assign n22868 = n22184 & n22864;
  assign n22869 = n22010 & ~n35178;
  assign n22870 = ~n22185 & n22869;
  assign n22871 = ~n22625 & n22870;
  assign n22872 = ~n22010 & ~n35268;
  assign n22873 = ~n22871 & ~n22872;
  assign n22874 = ~n22867 & ~n22868;
  assign n22875 = ~n22862 & ~n35269;
  assign n22876 = ~n22860 & ~n22875;
  assign n22877 = ~n11858 & ~n22876;
  assign n22878 = n11858 & ~n22860;
  assign n22879 = ~n22875 & n22878;
  assign n22880 = n11858 & n22876;
  assign n22881 = ~n22187 & ~n22203;
  assign n22882 = ~n22625 & n22881;
  assign n22883 = ~n35181 & ~n22882;
  assign n22884 = n35181 & ~n22203;
  assign n22885 = ~n22187 & n22884;
  assign n22886 = n35181 & n22882;
  assign n22887 = ~n22625 & n22885;
  assign n22888 = ~n22883 & ~n35271;
  assign n22889 = ~n35270 & ~n22888;
  assign n22890 = ~n22877 & ~n22889;
  assign n22891 = ~n11229 & ~n22890;
  assign n22892 = n11229 & ~n22877;
  assign n22893 = ~n22889 & n22892;
  assign n22894 = ~n35182 & ~n22209;
  assign n22895 = ~n22209 & ~n22625;
  assign n22896 = ~n35182 & n22895;
  assign n22897 = ~n22625 & n22894;
  assign n22898 = n22002 & ~n35272;
  assign n22899 = n22208 & n22895;
  assign n22900 = n22002 & ~n35182;
  assign n22901 = ~n22209 & n22900;
  assign n22902 = ~n22625 & n22901;
  assign n22903 = ~n22002 & ~n35272;
  assign n22904 = ~n22902 & ~n22903;
  assign n22905 = ~n22898 & ~n22899;
  assign n22906 = ~n22893 & ~n35273;
  assign n22907 = ~n22891 & ~n22906;
  assign n22908 = ~n10681 & ~n22907;
  assign n22909 = n10681 & ~n22891;
  assign n22910 = ~n22906 & n22909;
  assign n22911 = n10681 & n22907;
  assign n22912 = ~n22211 & ~n22222;
  assign n22913 = ~n22222 & ~n22625;
  assign n22914 = ~n22211 & n22913;
  assign n22915 = ~n22625 & n22912;
  assign n22916 = n22219 & ~n35275;
  assign n22917 = n22220 & n22913;
  assign n22918 = ~n22219 & n35275;
  assign n22919 = n22219 & ~n22222;
  assign n22920 = ~n22211 & n22919;
  assign n22921 = ~n22625 & n22920;
  assign n22922 = ~n22219 & ~n35275;
  assign n22923 = ~n22921 & ~n22922;
  assign n22924 = ~n22916 & ~n35276;
  assign n22925 = ~n35274 & ~n35277;
  assign n22926 = ~n22908 & ~n22925;
  assign n22927 = ~n10086 & ~n22926;
  assign n22928 = n10086 & ~n22908;
  assign n22929 = ~n22925 & n22928;
  assign n22930 = ~n35184 & ~n22228;
  assign n22931 = ~n22228 & ~n22625;
  assign n22932 = ~n35184 & n22931;
  assign n22933 = ~n22625 & n22930;
  assign n22934 = n21994 & ~n35278;
  assign n22935 = n22227 & n22931;
  assign n22936 = n21994 & ~n35184;
  assign n22937 = ~n22228 & n22936;
  assign n22938 = ~n22625 & n22937;
  assign n22939 = ~n21994 & ~n35278;
  assign n22940 = ~n22938 & ~n22939;
  assign n22941 = ~n22934 & ~n22935;
  assign n22942 = ~n22929 & ~n35279;
  assign n22943 = ~n22927 & ~n22942;
  assign n22944 = ~n9565 & ~n22943;
  assign n22945 = n9565 & ~n22927;
  assign n22946 = ~n22942 & n22945;
  assign n22947 = n9565 & n22943;
  assign n22948 = ~n22230 & ~n22246;
  assign n22949 = ~n22625 & n22948;
  assign n22950 = ~n35187 & n22949;
  assign n22951 = n35187 & ~n22949;
  assign n22952 = n35187 & ~n22246;
  assign n22953 = ~n22230 & n22952;
  assign n22954 = n35187 & n22949;
  assign n22955 = ~n22625 & n22953;
  assign n22956 = ~n35187 & ~n22949;
  assign n22957 = ~n35281 & ~n22956;
  assign n22958 = ~n22950 & ~n22951;
  assign n22959 = ~n35280 & ~n35282;
  assign n22960 = ~n22944 & ~n22959;
  assign n22961 = ~n8998 & ~n22960;
  assign n22962 = n8998 & ~n22944;
  assign n22963 = ~n22959 & n22962;
  assign n22964 = ~n35188 & ~n22252;
  assign n22965 = ~n22252 & ~n22625;
  assign n22966 = ~n35188 & n22965;
  assign n22967 = ~n22625 & n22964;
  assign n22968 = n21986 & ~n35283;
  assign n22969 = n22251 & n22965;
  assign n22970 = n21986 & ~n35188;
  assign n22971 = ~n22252 & n22970;
  assign n22972 = ~n22625 & n22971;
  assign n22973 = ~n21986 & ~n35283;
  assign n22974 = ~n22972 & ~n22973;
  assign n22975 = ~n22968 & ~n22969;
  assign n22976 = ~n22963 & ~n35284;
  assign n22977 = ~n22961 & ~n22976;
  assign n22978 = ~n8506 & ~n22977;
  assign n22979 = n8506 & ~n22961;
  assign n22980 = ~n22976 & n22979;
  assign n22981 = n8506 & n22977;
  assign n22982 = ~n22254 & ~n22268;
  assign n22983 = ~n22268 & ~n22625;
  assign n22984 = ~n22254 & n22983;
  assign n22985 = ~n22625 & n22982;
  assign n22986 = n35190 & ~n35286;
  assign n22987 = n22266 & n22983;
  assign n22988 = ~n35190 & n35286;
  assign n22989 = n35190 & ~n22268;
  assign n22990 = ~n22254 & n22989;
  assign n22991 = ~n22625 & n22990;
  assign n22992 = ~n35190 & ~n35286;
  assign n22993 = ~n22991 & ~n22992;
  assign n22994 = ~n22986 & ~n35287;
  assign n22995 = ~n35285 & ~n35288;
  assign n22996 = ~n22978 & ~n22995;
  assign n22997 = ~n7975 & ~n22996;
  assign n22998 = n7975 & ~n22978;
  assign n22999 = ~n22995 & n22998;
  assign n23000 = ~n35191 & ~n22274;
  assign n23001 = ~n22274 & ~n22625;
  assign n23002 = ~n35191 & n23001;
  assign n23003 = ~n22625 & n23000;
  assign n23004 = n21978 & ~n35289;
  assign n23005 = n22273 & n23001;
  assign n23006 = n21978 & ~n35191;
  assign n23007 = ~n22274 & n23006;
  assign n23008 = ~n22625 & n23007;
  assign n23009 = ~n21978 & ~n35289;
  assign n23010 = ~n23008 & ~n23009;
  assign n23011 = ~n23004 & ~n23005;
  assign n23012 = ~n22999 & ~n35290;
  assign n23013 = ~n22997 & ~n23012;
  assign n23014 = ~n7512 & ~n23013;
  assign n23015 = ~n22276 & ~n22292;
  assign n23016 = ~n22625 & n23015;
  assign n23017 = ~n35194 & ~n23016;
  assign n23018 = n35194 & ~n22292;
  assign n23019 = ~n22276 & n23018;
  assign n23020 = n35194 & n23016;
  assign n23021 = ~n22625 & n23019;
  assign n23022 = ~n23017 & ~n35291;
  assign n23023 = n7512 & ~n22997;
  assign n23024 = ~n23012 & n23023;
  assign n23025 = n7512 & n23013;
  assign n23026 = ~n23022 & ~n35292;
  assign n23027 = ~n23014 & ~n23026;
  assign n23028 = ~n7015 & ~n23027;
  assign n23029 = n7015 & ~n23014;
  assign n23030 = ~n23026 & n23029;
  assign n23031 = ~n35195 & ~n22298;
  assign n23032 = ~n22298 & ~n22625;
  assign n23033 = ~n35195 & n23032;
  assign n23034 = ~n22625 & n23031;
  assign n23035 = n21970 & ~n35293;
  assign n23036 = n22297 & n23032;
  assign n23037 = n21970 & ~n35195;
  assign n23038 = ~n22298 & n23037;
  assign n23039 = ~n22625 & n23038;
  assign n23040 = ~n21970 & ~n35293;
  assign n23041 = ~n23039 & ~n23040;
  assign n23042 = ~n23035 & ~n23036;
  assign n23043 = ~n23030 & ~n35294;
  assign n23044 = ~n23028 & ~n23043;
  assign n23045 = ~n6579 & ~n23044;
  assign n23046 = n6579 & ~n23028;
  assign n23047 = ~n23043 & n23046;
  assign n23048 = n6579 & n23044;
  assign n23049 = ~n22300 & ~n22303;
  assign n23050 = ~n22303 & ~n22625;
  assign n23051 = ~n22300 & n23050;
  assign n23052 = ~n22625 & n23049;
  assign n23053 = n21962 & ~n35296;
  assign n23054 = n22301 & n23050;
  assign n23055 = n21962 & ~n22303;
  assign n23056 = ~n22300 & n23055;
  assign n23057 = ~n22625 & n23056;
  assign n23058 = ~n21962 & ~n35296;
  assign n23059 = ~n23057 & ~n23058;
  assign n23060 = ~n23053 & ~n23054;
  assign n23061 = ~n35295 & ~n35297;
  assign n23062 = ~n23045 & ~n23061;
  assign n23063 = ~n6117 & ~n23062;
  assign n23064 = n6117 & ~n23045;
  assign n23065 = ~n23061 & n23064;
  assign n23066 = ~n35196 & ~n22309;
  assign n23067 = ~n22309 & ~n22625;
  assign n23068 = ~n35196 & n23067;
  assign n23069 = ~n22625 & n23066;
  assign n23070 = n21954 & ~n35298;
  assign n23071 = n22308 & n23067;
  assign n23072 = n21954 & ~n35196;
  assign n23073 = ~n22309 & n23072;
  assign n23074 = ~n22625 & n23073;
  assign n23075 = ~n21954 & ~n35298;
  assign n23076 = ~n23074 & ~n23075;
  assign n23077 = ~n23070 & ~n23071;
  assign n23078 = ~n23065 & ~n35299;
  assign n23079 = ~n23063 & ~n23078;
  assign n23080 = ~n5708 & ~n23079;
  assign n23081 = ~n22311 & ~n22326;
  assign n23082 = ~n22625 & n23081;
  assign n23083 = ~n35198 & ~n23082;
  assign n23084 = n35198 & ~n22326;
  assign n23085 = ~n22311 & n23084;
  assign n23086 = n35198 & n23082;
  assign n23087 = ~n22625 & n23085;
  assign n23088 = ~n23083 & ~n35300;
  assign n23089 = n5708 & ~n23063;
  assign n23090 = ~n23078 & n23089;
  assign n23091 = n5708 & n23079;
  assign n23092 = ~n23088 & ~n35301;
  assign n23093 = ~n23080 & ~n23092;
  assign n23094 = ~n5278 & ~n23093;
  assign n23095 = n5278 & ~n23080;
  assign n23096 = ~n23092 & n23095;
  assign n23097 = ~n35199 & ~n22332;
  assign n23098 = ~n22332 & ~n22625;
  assign n23099 = ~n35199 & n23098;
  assign n23100 = ~n22625 & n23097;
  assign n23101 = n21946 & ~n35302;
  assign n23102 = n22331 & n23098;
  assign n23103 = n21946 & ~n35199;
  assign n23104 = ~n22332 & n23103;
  assign n23105 = ~n22625 & n23104;
  assign n23106 = ~n21946 & ~n35302;
  assign n23107 = ~n23105 & ~n23106;
  assign n23108 = ~n23101 & ~n23102;
  assign n23109 = ~n23096 & ~n35303;
  assign n23110 = ~n23094 & ~n23109;
  assign n23111 = ~n4903 & ~n23110;
  assign n23112 = n4903 & ~n23094;
  assign n23113 = ~n23109 & n23112;
  assign n23114 = n4903 & n23110;
  assign n23115 = ~n22334 & ~n22337;
  assign n23116 = ~n22337 & ~n22625;
  assign n23117 = ~n22334 & n23116;
  assign n23118 = ~n22625 & n23115;
  assign n23119 = n21938 & ~n35305;
  assign n23120 = n22335 & n23116;
  assign n23121 = n21938 & ~n22337;
  assign n23122 = ~n22334 & n23121;
  assign n23123 = ~n22625 & n23122;
  assign n23124 = ~n21938 & ~n35305;
  assign n23125 = ~n23123 & ~n23124;
  assign n23126 = ~n23119 & ~n23120;
  assign n23127 = ~n35304 & ~n35306;
  assign n23128 = ~n23111 & ~n23127;
  assign n23129 = ~n4508 & ~n23128;
  assign n23130 = n4508 & ~n23111;
  assign n23131 = ~n23127 & n23130;
  assign n23132 = ~n35200 & ~n22343;
  assign n23133 = ~n22343 & ~n22625;
  assign n23134 = ~n35200 & n23133;
  assign n23135 = ~n22625 & n23132;
  assign n23136 = n21930 & ~n35307;
  assign n23137 = n22342 & n23133;
  assign n23138 = n21930 & ~n35200;
  assign n23139 = ~n22343 & n23138;
  assign n23140 = ~n22625 & n23139;
  assign n23141 = ~n21930 & ~n35307;
  assign n23142 = ~n23140 & ~n23141;
  assign n23143 = ~n23136 & ~n23137;
  assign n23144 = ~n23131 & ~n35308;
  assign n23145 = ~n23129 & ~n23144;
  assign n23146 = ~n4155 & ~n23145;
  assign n23147 = ~n22345 & ~n22360;
  assign n23148 = ~n22625 & n23147;
  assign n23149 = ~n35202 & ~n23148;
  assign n23150 = n35202 & ~n22360;
  assign n23151 = ~n22345 & n23150;
  assign n23152 = n35202 & n23148;
  assign n23153 = ~n22625 & n23151;
  assign n23154 = ~n23149 & ~n35309;
  assign n23155 = n4155 & ~n23129;
  assign n23156 = ~n23144 & n23155;
  assign n23157 = n4155 & n23145;
  assign n23158 = ~n23154 & ~n35310;
  assign n23159 = ~n23146 & ~n23158;
  assign n23160 = ~n3788 & ~n23159;
  assign n23161 = n3788 & ~n23146;
  assign n23162 = ~n23158 & n23161;
  assign n23163 = ~n35203 & ~n22366;
  assign n23164 = ~n22366 & ~n22625;
  assign n23165 = ~n35203 & n23164;
  assign n23166 = ~n22625 & n23163;
  assign n23167 = n21922 & ~n35311;
  assign n23168 = n22365 & n23164;
  assign n23169 = n21922 & ~n35203;
  assign n23170 = ~n22366 & n23169;
  assign n23171 = ~n22625 & n23170;
  assign n23172 = ~n21922 & ~n35311;
  assign n23173 = ~n23171 & ~n23172;
  assign n23174 = ~n23167 & ~n23168;
  assign n23175 = ~n23162 & ~n35312;
  assign n23176 = ~n23160 & ~n23175;
  assign n23177 = ~n3473 & ~n23176;
  assign n23178 = n3473 & ~n23160;
  assign n23179 = ~n23175 & n23178;
  assign n23180 = n3473 & n23176;
  assign n23181 = ~n22368 & ~n22371;
  assign n23182 = ~n22371 & ~n22625;
  assign n23183 = ~n22368 & n23182;
  assign n23184 = ~n22625 & n23181;
  assign n23185 = n21914 & ~n35314;
  assign n23186 = n22369 & n23182;
  assign n23187 = n21914 & ~n22371;
  assign n23188 = ~n22368 & n23187;
  assign n23189 = ~n22625 & n23188;
  assign n23190 = ~n21914 & ~n35314;
  assign n23191 = ~n23189 & ~n23190;
  assign n23192 = ~n23185 & ~n23186;
  assign n23193 = ~n35313 & ~n35315;
  assign n23194 = ~n23177 & ~n23193;
  assign n23195 = ~n3140 & ~n23194;
  assign n23196 = n3140 & ~n23177;
  assign n23197 = ~n23193 & n23196;
  assign n23198 = ~n35204 & ~n22377;
  assign n23199 = ~n22377 & ~n22625;
  assign n23200 = ~n35204 & n23199;
  assign n23201 = ~n22625 & n23198;
  assign n23202 = n21906 & ~n35316;
  assign n23203 = n22376 & n23199;
  assign n23204 = n21906 & ~n35204;
  assign n23205 = ~n22377 & n23204;
  assign n23206 = ~n22625 & n23205;
  assign n23207 = ~n21906 & ~n35316;
  assign n23208 = ~n23206 & ~n23207;
  assign n23209 = ~n23202 & ~n23203;
  assign n23210 = ~n23197 & ~n35317;
  assign n23211 = ~n23195 & ~n23210;
  assign n23212 = ~n2855 & ~n23211;
  assign n23213 = ~n22379 & ~n22394;
  assign n23214 = ~n22625 & n23213;
  assign n23215 = ~n35206 & ~n23214;
  assign n23216 = n35206 & ~n22394;
  assign n23217 = ~n22379 & n23216;
  assign n23218 = n35206 & n23214;
  assign n23219 = ~n22625 & n23217;
  assign n23220 = ~n23215 & ~n35318;
  assign n23221 = n2855 & ~n23195;
  assign n23222 = ~n23210 & n23221;
  assign n23223 = n2855 & n23211;
  assign n23224 = ~n23220 & ~n35319;
  assign n23225 = ~n23212 & ~n23224;
  assign n23226 = ~n2556 & ~n23225;
  assign n23227 = n2556 & ~n23212;
  assign n23228 = ~n23224 & n23227;
  assign n23229 = ~n35207 & ~n22400;
  assign n23230 = ~n22400 & ~n22625;
  assign n23231 = ~n35207 & n23230;
  assign n23232 = ~n22625 & n23229;
  assign n23233 = n21898 & ~n35320;
  assign n23234 = n22399 & n23230;
  assign n23235 = n21898 & ~n35207;
  assign n23236 = ~n22400 & n23235;
  assign n23237 = ~n22625 & n23236;
  assign n23238 = ~n21898 & ~n35320;
  assign n23239 = ~n23237 & ~n23238;
  assign n23240 = ~n23233 & ~n23234;
  assign n23241 = ~n23228 & ~n35321;
  assign n23242 = ~n23226 & ~n23241;
  assign n23243 = ~n2301 & ~n23242;
  assign n23244 = n2301 & ~n23226;
  assign n23245 = ~n23241 & n23244;
  assign n23246 = n2301 & n23242;
  assign n23247 = ~n22402 & ~n22405;
  assign n23248 = ~n22405 & ~n22625;
  assign n23249 = ~n22402 & n23248;
  assign n23250 = ~n22625 & n23247;
  assign n23251 = n21890 & ~n35323;
  assign n23252 = n22403 & n23248;
  assign n23253 = n21890 & ~n22405;
  assign n23254 = ~n22402 & n23253;
  assign n23255 = ~n22625 & n23254;
  assign n23256 = ~n21890 & ~n35323;
  assign n23257 = ~n23255 & ~n23256;
  assign n23258 = ~n23251 & ~n23252;
  assign n23259 = ~n35322 & ~n35324;
  assign n23260 = ~n23243 & ~n23259;
  assign n23261 = ~n2038 & ~n23260;
  assign n23262 = n2038 & ~n23243;
  assign n23263 = ~n23259 & n23262;
  assign n23264 = ~n35208 & ~n22411;
  assign n23265 = ~n22411 & ~n22625;
  assign n23266 = ~n35208 & n23265;
  assign n23267 = ~n22625 & n23264;
  assign n23268 = n21882 & ~n35325;
  assign n23269 = n22410 & n23265;
  assign n23270 = n21882 & ~n35208;
  assign n23271 = ~n22411 & n23270;
  assign n23272 = ~n22625 & n23271;
  assign n23273 = ~n21882 & ~n35325;
  assign n23274 = ~n23272 & ~n23273;
  assign n23275 = ~n23268 & ~n23269;
  assign n23276 = ~n23263 & ~n35326;
  assign n23277 = ~n23261 & ~n23276;
  assign n23278 = ~n1812 & ~n23277;
  assign n23279 = ~n22413 & ~n22428;
  assign n23280 = ~n22625 & n23279;
  assign n23281 = ~n35210 & ~n23280;
  assign n23282 = n35210 & ~n22428;
  assign n23283 = ~n22413 & n23282;
  assign n23284 = n35210 & n23280;
  assign n23285 = ~n22625 & n23283;
  assign n23286 = ~n23281 & ~n35327;
  assign n23287 = n1812 & ~n23261;
  assign n23288 = ~n23276 & n23287;
  assign n23289 = n1812 & n23277;
  assign n23290 = ~n23286 & ~n35328;
  assign n23291 = ~n23278 & ~n23290;
  assign n23292 = ~n1582 & ~n23291;
  assign n23293 = n1582 & ~n23278;
  assign n23294 = ~n23290 & n23293;
  assign n23295 = ~n35211 & ~n22434;
  assign n23296 = ~n22434 & ~n22625;
  assign n23297 = ~n35211 & n23296;
  assign n23298 = ~n22625 & n23295;
  assign n23299 = n21874 & ~n35329;
  assign n23300 = n22433 & n23296;
  assign n23301 = n21874 & ~n35211;
  assign n23302 = ~n22434 & n23301;
  assign n23303 = ~n22625 & n23302;
  assign n23304 = ~n21874 & ~n35329;
  assign n23305 = ~n23303 & ~n23304;
  assign n23306 = ~n23299 & ~n23300;
  assign n23307 = ~n23294 & ~n35330;
  assign n23308 = ~n23292 & ~n23307;
  assign n23309 = ~n1388 & ~n23308;
  assign n23310 = n1388 & ~n23292;
  assign n23311 = ~n23307 & n23310;
  assign n23312 = n1388 & n23308;
  assign n23313 = ~n22436 & ~n22439;
  assign n23314 = ~n22439 & ~n22625;
  assign n23315 = ~n22436 & n23314;
  assign n23316 = ~n22625 & n23313;
  assign n23317 = n21866 & ~n35332;
  assign n23318 = n22437 & n23314;
  assign n23319 = n21866 & ~n22439;
  assign n23320 = ~n22436 & n23319;
  assign n23321 = ~n22625 & n23320;
  assign n23322 = ~n21866 & ~n35332;
  assign n23323 = ~n23321 & ~n23322;
  assign n23324 = ~n23317 & ~n23318;
  assign n23325 = ~n35331 & ~n35333;
  assign n23326 = ~n23309 & ~n23325;
  assign n23327 = ~n1192 & ~n23326;
  assign n23328 = n1192 & ~n23309;
  assign n23329 = ~n23325 & n23328;
  assign n23330 = n21858 & ~n35212;
  assign n23331 = ~n22445 & n23330;
  assign n23332 = ~n35212 & ~n22445;
  assign n23333 = ~n22625 & n23332;
  assign n23334 = n21858 & n23333;
  assign n23335 = ~n22625 & n23331;
  assign n23336 = ~n21858 & ~n23333;
  assign n23337 = ~n35334 & ~n23336;
  assign n23338 = ~n23329 & ~n23337;
  assign n23339 = ~n23327 & ~n23338;
  assign n23340 = ~n1028 & ~n23339;
  assign n23341 = n1028 & ~n23327;
  assign n23342 = ~n23338 & n23341;
  assign n23343 = n1028 & n23339;
  assign n23344 = ~n22447 & ~n22449;
  assign n23345 = ~n22625 & n23344;
  assign n23346 = ~n35214 & n23345;
  assign n23347 = n35214 & ~n23345;
  assign n23348 = ~n22447 & n35214;
  assign n23349 = ~n22449 & n23348;
  assign n23350 = n35214 & n23345;
  assign n23351 = ~n22625 & n23349;
  assign n23352 = ~n35214 & ~n23345;
  assign n23353 = ~n35336 & ~n23352;
  assign n23354 = ~n23346 & ~n23347;
  assign n23355 = ~n35335 & ~n35337;
  assign n23356 = ~n23340 & ~n23355;
  assign n23357 = ~n866 & ~n23356;
  assign n23358 = n866 & ~n23340;
  assign n23359 = ~n23355 & n23358;
  assign n23360 = ~n35236 & ~n23359;
  assign n23361 = ~n23357 & ~n23360;
  assign n23362 = ~n730 & ~n23361;
  assign n23363 = ~n22469 & ~n22471;
  assign n23364 = ~n22625 & n23363;
  assign n23365 = ~n35217 & ~n23364;
  assign n23366 = ~n22469 & n35217;
  assign n23367 = ~n22471 & n23366;
  assign n23368 = n35217 & n23364;
  assign n23369 = ~n22625 & n23367;
  assign n23370 = ~n23365 & ~n35338;
  assign n23371 = n730 & ~n23357;
  assign n23372 = ~n23360 & n23371;
  assign n23373 = n730 & n23361;
  assign n23374 = ~n23370 & ~n35339;
  assign n23375 = ~n23362 & ~n23374;
  assign n23376 = ~n602 & ~n23375;
  assign n23377 = n602 & ~n23362;
  assign n23378 = ~n23374 & n23377;
  assign n23379 = ~n22486 & ~n35219;
  assign n23380 = ~n22486 & ~n22625;
  assign n23381 = ~n35219 & n23380;
  assign n23382 = ~n22625 & n23379;
  assign n23383 = n22494 & ~n35340;
  assign n23384 = n22498 & n23380;
  assign n23385 = n22494 & ~n35219;
  assign n23386 = ~n22486 & n23385;
  assign n23387 = ~n22625 & n23386;
  assign n23388 = ~n22494 & ~n35340;
  assign n23389 = ~n23387 & ~n23388;
  assign n23390 = ~n23383 & ~n23384;
  assign n23391 = ~n23378 & ~n35341;
  assign n23392 = ~n23376 & ~n23391;
  assign n23393 = ~n497 & ~n23392;
  assign n23394 = ~n22500 & ~n22502;
  assign n23395 = ~n22625 & n23394;
  assign n23396 = ~n35221 & ~n23395;
  assign n23397 = ~n22500 & n35221;
  assign n23398 = ~n22502 & n23397;
  assign n23399 = n35221 & n23395;
  assign n23400 = ~n22625 & n23398;
  assign n23401 = ~n23396 & ~n35342;
  assign n23402 = n497 & ~n23376;
  assign n23403 = ~n23391 & n23402;
  assign n23404 = n497 & n23392;
  assign n23405 = ~n23401 & ~n35343;
  assign n23406 = ~n23393 & ~n23405;
  assign n23407 = ~n403 & ~n23406;
  assign n23408 = n403 & ~n23393;
  assign n23409 = ~n23405 & n23408;
  assign n23410 = ~n22517 & ~n35223;
  assign n23411 = ~n22517 & ~n22625;
  assign n23412 = ~n35223 & n23411;
  assign n23413 = ~n22625 & n23410;
  assign n23414 = n22525 & ~n35344;
  assign n23415 = n22529 & n23411;
  assign n23416 = n22525 & ~n35223;
  assign n23417 = ~n22517 & n23416;
  assign n23418 = ~n22625 & n23417;
  assign n23419 = ~n22525 & ~n35344;
  assign n23420 = ~n23418 & ~n23419;
  assign n23421 = ~n23414 & ~n23415;
  assign n23422 = ~n23409 & ~n35345;
  assign n23423 = ~n23407 & ~n23422;
  assign n23424 = ~n330 & ~n23423;
  assign n23425 = n330 & ~n23407;
  assign n23426 = ~n23422 & n23425;
  assign n23427 = n330 & n23423;
  assign n23428 = ~n22531 & ~n22541;
  assign n23429 = ~n22531 & ~n22625;
  assign n23430 = ~n22541 & n23429;
  assign n23431 = ~n22625 & n23428;
  assign n23432 = n22539 & ~n35347;
  assign n23433 = n22542 & n23429;
  assign n23434 = ~n22531 & n22539;
  assign n23435 = ~n22541 & n23434;
  assign n23436 = ~n22625 & n23435;
  assign n23437 = ~n22539 & ~n35347;
  assign n23438 = ~n23436 & ~n23437;
  assign n23439 = ~n23432 & ~n23433;
  assign n23440 = ~n35346 & ~n35348;
  assign n23441 = ~n23424 & ~n23440;
  assign n23442 = ~n271 & ~n23441;
  assign n23443 = n271 & ~n23424;
  assign n23444 = ~n23440 & n23443;
  assign n23445 = ~n22544 & ~n35226;
  assign n23446 = ~n22544 & ~n22625;
  assign n23447 = ~n35226 & n23446;
  assign n23448 = ~n22625 & n23445;
  assign n23449 = n22552 & ~n35349;
  assign n23450 = n22556 & n23446;
  assign n23451 = n22552 & ~n35226;
  assign n23452 = ~n22544 & n23451;
  assign n23453 = ~n22625 & n23452;
  assign n23454 = ~n22552 & ~n35349;
  assign n23455 = ~n23453 & ~n23454;
  assign n23456 = ~n23449 & ~n23450;
  assign n23457 = ~n23444 & ~n35350;
  assign n23458 = ~n23442 & ~n23457;
  assign n23459 = ~n217 & ~n23458;
  assign n23460 = ~n22558 & ~n22560;
  assign n23461 = ~n22625 & n23460;
  assign n23462 = ~n35228 & ~n23461;
  assign n23463 = ~n22558 & n35228;
  assign n23464 = ~n22560 & n23463;
  assign n23465 = n35228 & n23461;
  assign n23466 = ~n22625 & n23464;
  assign n23467 = ~n23462 & ~n35351;
  assign n23468 = n217 & ~n23442;
  assign n23469 = ~n23457 & n23468;
  assign n23470 = n217 & n23458;
  assign n23471 = ~n23467 & ~n35352;
  assign n23472 = ~n23459 & ~n23471;
  assign n23473 = ~n198 & ~n23472;
  assign n23474 = n198 & ~n23459;
  assign n23475 = ~n23471 & n23474;
  assign n23476 = ~n22575 & ~n35230;
  assign n23477 = ~n22575 & ~n22625;
  assign n23478 = ~n35230 & n23477;
  assign n23479 = ~n22625 & n23476;
  assign n23480 = n22583 & ~n35353;
  assign n23481 = n22587 & n23477;
  assign n23482 = n22583 & ~n35230;
  assign n23483 = ~n22575 & n23482;
  assign n23484 = ~n22625 & n23483;
  assign n23485 = ~n22583 & ~n35353;
  assign n23486 = ~n23484 & ~n23485;
  assign n23487 = ~n23480 & ~n23481;
  assign n23488 = ~n23475 & ~n35354;
  assign n23489 = ~n23473 & ~n23488;
  assign n23490 = ~n22589 & ~n22599;
  assign n23491 = ~n22589 & ~n22625;
  assign n23492 = ~n22599 & n23491;
  assign n23493 = ~n22625 & n23490;
  assign n23494 = n22597 & ~n35355;
  assign n23495 = n22600 & n23491;
  assign n23496 = ~n22589 & n22597;
  assign n23497 = ~n22599 & n23496;
  assign n23498 = ~n22625 & n23497;
  assign n23499 = ~n22597 & ~n35355;
  assign n23500 = ~n23498 & ~n23499;
  assign n23501 = ~n23494 & ~n23495;
  assign n23502 = ~n22601 & ~n22609;
  assign n23503 = ~n22609 & ~n22625;
  assign n23504 = ~n22601 & n23503;
  assign n23505 = ~n22625 & n23502;
  assign n23506 = ~n35234 & ~n35357;
  assign n23507 = ~n35356 & n23506;
  assign n23508 = ~n23489 & n23507;
  assign n23509 = n193 & ~n23508;
  assign n23510 = ~n23473 & n35356;
  assign n23511 = ~n23488 & n23510;
  assign n23512 = n23489 & n35356;
  assign n23513 = n22601 & ~n23503;
  assign n23514 = ~n193 & ~n23502;
  assign n23515 = ~n23513 & n23514;
  assign n23516 = ~n35358 & ~n23515;
  assign n23517 = ~n23509 & n23516;
  assign n23518 = ~n23357 & ~n23359;
  assign n23519 = ~n23517 & n23518;
  assign n23520 = ~n35236 & ~n23519;
  assign n23521 = n35236 & ~n23359;
  assign n23522 = ~n23357 & n23521;
  assign n23523 = n35236 & n23519;
  assign n23524 = ~n23517 & n23522;
  assign n23525 = ~n23520 & ~n35359;
  assign n23526 = ~n23327 & ~n23329;
  assign n23527 = ~n23517 & n23526;
  assign n23528 = ~n23337 & ~n23527;
  assign n23529 = ~n23329 & n23337;
  assign n23530 = ~n23327 & n23529;
  assign n23531 = n23337 & n23527;
  assign n23532 = ~n23517 & n23530;
  assign n23533 = ~n23528 & ~n35360;
  assign n23534 = ~n23309 & ~n35331;
  assign n23535 = ~n23517 & n23534;
  assign n23536 = ~n35333 & ~n23535;
  assign n23537 = ~n23309 & n35333;
  assign n23538 = ~n35331 & n23537;
  assign n23539 = n35333 & n23535;
  assign n23540 = ~n23517 & n23538;
  assign n23541 = ~n23536 & ~n35361;
  assign n23542 = ~n23292 & ~n23294;
  assign n23543 = ~n23517 & n23542;
  assign n23544 = ~n35330 & ~n23543;
  assign n23545 = ~n23294 & n35330;
  assign n23546 = ~n23292 & n23545;
  assign n23547 = n35330 & n23543;
  assign n23548 = ~n23517 & n23546;
  assign n23549 = ~n23544 & ~n35362;
  assign n23550 = ~n23261 & ~n23263;
  assign n23551 = ~n23517 & n23550;
  assign n23552 = ~n35326 & ~n23551;
  assign n23553 = ~n23263 & n35326;
  assign n23554 = ~n23261 & n23553;
  assign n23555 = n35326 & n23551;
  assign n23556 = ~n23517 & n23554;
  assign n23557 = ~n23552 & ~n35363;
  assign n23558 = ~n23243 & ~n35322;
  assign n23559 = ~n23517 & n23558;
  assign n23560 = ~n35324 & ~n23559;
  assign n23561 = ~n23243 & n35324;
  assign n23562 = ~n35322 & n23561;
  assign n23563 = n35324 & n23559;
  assign n23564 = ~n23517 & n23562;
  assign n23565 = ~n23560 & ~n35364;
  assign n23566 = ~n23226 & ~n23228;
  assign n23567 = ~n23517 & n23566;
  assign n23568 = ~n35321 & ~n23567;
  assign n23569 = ~n23228 & n35321;
  assign n23570 = ~n23226 & n23569;
  assign n23571 = n35321 & n23567;
  assign n23572 = ~n23517 & n23570;
  assign n23573 = ~n23568 & ~n35365;
  assign n23574 = ~n23195 & ~n23197;
  assign n23575 = ~n23517 & n23574;
  assign n23576 = ~n35317 & ~n23575;
  assign n23577 = ~n23197 & n35317;
  assign n23578 = ~n23195 & n23577;
  assign n23579 = n35317 & n23575;
  assign n23580 = ~n23517 & n23578;
  assign n23581 = ~n23576 & ~n35366;
  assign n23582 = ~n23177 & ~n35313;
  assign n23583 = ~n23517 & n23582;
  assign n23584 = ~n35315 & ~n23583;
  assign n23585 = ~n23177 & n35315;
  assign n23586 = ~n35313 & n23585;
  assign n23587 = n35315 & n23583;
  assign n23588 = ~n23517 & n23586;
  assign n23589 = ~n23584 & ~n35367;
  assign n23590 = ~n23160 & ~n23162;
  assign n23591 = ~n23517 & n23590;
  assign n23592 = ~n35312 & ~n23591;
  assign n23593 = ~n23162 & n35312;
  assign n23594 = ~n23160 & n23593;
  assign n23595 = n35312 & n23591;
  assign n23596 = ~n23517 & n23594;
  assign n23597 = ~n23592 & ~n35368;
  assign n23598 = ~n23129 & ~n23131;
  assign n23599 = ~n23517 & n23598;
  assign n23600 = ~n35308 & ~n23599;
  assign n23601 = ~n23131 & n35308;
  assign n23602 = ~n23129 & n23601;
  assign n23603 = n35308 & n23599;
  assign n23604 = ~n23517 & n23602;
  assign n23605 = ~n23600 & ~n35369;
  assign n23606 = ~n23111 & ~n35304;
  assign n23607 = ~n23517 & n23606;
  assign n23608 = ~n35306 & ~n23607;
  assign n23609 = ~n23111 & n35306;
  assign n23610 = ~n35304 & n23609;
  assign n23611 = n35306 & n23607;
  assign n23612 = ~n23517 & n23610;
  assign n23613 = ~n23608 & ~n35370;
  assign n23614 = ~n23094 & ~n23096;
  assign n23615 = ~n23517 & n23614;
  assign n23616 = ~n35303 & ~n23615;
  assign n23617 = ~n23096 & n35303;
  assign n23618 = ~n23094 & n23617;
  assign n23619 = n35303 & n23615;
  assign n23620 = ~n23517 & n23618;
  assign n23621 = ~n23616 & ~n35371;
  assign n23622 = ~n23063 & ~n23065;
  assign n23623 = ~n23517 & n23622;
  assign n23624 = ~n35299 & ~n23623;
  assign n23625 = ~n23065 & n35299;
  assign n23626 = ~n23063 & n23625;
  assign n23627 = n35299 & n23623;
  assign n23628 = ~n23517 & n23626;
  assign n23629 = ~n23624 & ~n35372;
  assign n23630 = ~n23045 & ~n35295;
  assign n23631 = ~n23517 & n23630;
  assign n23632 = ~n35297 & ~n23631;
  assign n23633 = ~n23045 & n35297;
  assign n23634 = ~n35295 & n23633;
  assign n23635 = n35297 & n23631;
  assign n23636 = ~n23517 & n23634;
  assign n23637 = ~n23632 & ~n35373;
  assign n23638 = ~n23028 & ~n23030;
  assign n23639 = ~n23517 & n23638;
  assign n23640 = ~n35294 & ~n23639;
  assign n23641 = ~n23030 & n35294;
  assign n23642 = ~n23028 & n23641;
  assign n23643 = n35294 & n23639;
  assign n23644 = ~n23517 & n23642;
  assign n23645 = ~n23640 & ~n35374;
  assign n23646 = ~n22997 & ~n22999;
  assign n23647 = ~n23517 & n23646;
  assign n23648 = ~n35290 & ~n23647;
  assign n23649 = ~n22999 & n35290;
  assign n23650 = ~n22997 & n23649;
  assign n23651 = n35290 & n23647;
  assign n23652 = ~n23517 & n23650;
  assign n23653 = ~n23648 & ~n35375;
  assign n23654 = ~n22978 & ~n35285;
  assign n23655 = ~n23517 & n23654;
  assign n23656 = ~n35288 & ~n23655;
  assign n23657 = ~n22978 & n35288;
  assign n23658 = ~n35285 & n23657;
  assign n23659 = n35288 & n23655;
  assign n23660 = ~n23517 & n23658;
  assign n23661 = ~n23656 & ~n35376;
  assign n23662 = ~n22961 & ~n22963;
  assign n23663 = ~n23517 & n23662;
  assign n23664 = ~n35284 & ~n23663;
  assign n23665 = ~n22963 & n35284;
  assign n23666 = ~n22961 & n23665;
  assign n23667 = n35284 & n23663;
  assign n23668 = ~n23517 & n23666;
  assign n23669 = ~n23664 & ~n35377;
  assign n23670 = ~n22927 & ~n22929;
  assign n23671 = ~n23517 & n23670;
  assign n23672 = ~n35279 & ~n23671;
  assign n23673 = ~n22929 & n35279;
  assign n23674 = ~n22927 & n23673;
  assign n23675 = n35279 & n23671;
  assign n23676 = ~n23517 & n23674;
  assign n23677 = ~n23672 & ~n35378;
  assign n23678 = ~n22891 & ~n22893;
  assign n23679 = ~n23517 & n23678;
  assign n23680 = ~n35273 & ~n23679;
  assign n23681 = ~n22893 & n35273;
  assign n23682 = ~n22891 & n23681;
  assign n23683 = n35273 & n23679;
  assign n23684 = ~n23517 & n23682;
  assign n23685 = ~n23680 & ~n35379;
  assign n23686 = ~n22860 & ~n22862;
  assign n23687 = ~n23517 & n23686;
  assign n23688 = ~n35269 & ~n23687;
  assign n23689 = ~n22862 & n35269;
  assign n23690 = ~n22860 & n23689;
  assign n23691 = n35269 & n23687;
  assign n23692 = ~n23517 & n23690;
  assign n23693 = ~n23688 & ~n35380;
  assign n23694 = ~n22824 & ~n22826;
  assign n23695 = ~n23517 & n23694;
  assign n23696 = ~n35263 & ~n23695;
  assign n23697 = ~n22826 & n35263;
  assign n23698 = ~n22824 & n23697;
  assign n23699 = n35263 & n23695;
  assign n23700 = ~n23517 & n23698;
  assign n23701 = ~n23696 & ~n35381;
  assign n23702 = ~n22790 & ~n22792;
  assign n23703 = ~n23517 & n23702;
  assign n23704 = ~n35258 & ~n23703;
  assign n23705 = ~n22792 & n35258;
  assign n23706 = ~n22790 & n23705;
  assign n23707 = n35258 & n23703;
  assign n23708 = ~n23517 & n23706;
  assign n23709 = ~n23704 & ~n35382;
  assign n23710 = ~n22756 & ~n22758;
  assign n23711 = ~n23517 & n23710;
  assign n23712 = ~n35253 & ~n23711;
  assign n23713 = ~n22758 & n35253;
  assign n23714 = ~n22756 & n23713;
  assign n23715 = n35253 & n23711;
  assign n23716 = ~n23517 & n23714;
  assign n23717 = ~n23712 & ~n35383;
  assign n23718 = ~n22723 & ~n22725;
  assign n23719 = ~n23517 & n23718;
  assign n23720 = ~n35249 & ~n23719;
  assign n23721 = ~n22725 & n35249;
  assign n23722 = ~n22723 & n23721;
  assign n23723 = n35249 & n23719;
  assign n23724 = ~n23517 & n23722;
  assign n23725 = ~n23720 & ~n35384;
  assign n23726 = ~n22689 & ~n22691;
  assign n23727 = ~n23517 & n23726;
  assign n23728 = ~n35244 & ~n23727;
  assign n23729 = ~n22691 & n35244;
  assign n23730 = ~n22689 & n23729;
  assign n23731 = n35244 & n23727;
  assign n23732 = ~n23517 & n23730;
  assign n23733 = ~n23728 & ~n35385;
  assign n23734 = ~n22662 & ~n22664;
  assign n23735 = ~n23517 & n23734;
  assign n23736 = ~n22673 & ~n23735;
  assign n23737 = ~n22664 & n22673;
  assign n23738 = ~n22662 & n23737;
  assign n23739 = n22673 & n23735;
  assign n23740 = ~n23517 & n23738;
  assign n23741 = ~n23736 & ~n35386;
  assign n23742 = ~pi18  & ~n23517;
  assign n23743 = ~pi19  & n23742;
  assign n23744 = n22639 & ~n23517;
  assign n23745 = ~n22625 & ~n23515;
  assign n23746 = ~n35358 & n23745;
  assign n23747 = ~n23509 & n23746;
  assign n23748 = ~n35387 & ~n23747;
  assign n23749 = pi20  & ~n23748;
  assign n23750 = ~pi20  & ~n23747;
  assign n23751 = ~pi20  & n23748;
  assign n23752 = ~n35387 & n23750;
  assign n23753 = ~n23749 & ~n35388;
  assign n23754 = pi18  & ~n23517;
  assign n23755 = ~pi16  & ~pi17 ;
  assign n23756 = ~pi18  & n23755;
  assign n23757 = ~n35133 & ~n35238;
  assign n23758 = ~n21821 & n23757;
  assign n23759 = ~n21840 & n23758;
  assign n23760 = ~n35135 & n23759;
  assign n23761 = n21826 & n21842;
  assign n23762 = ~n21834 & n23760;
  assign n23763 = ~n23756 & ~n35389;
  assign n23764 = ~n22623 & n23763;
  assign n23765 = ~n35234 & n23764;
  assign n23766 = ~n22617 & n23765;
  assign n23767 = ~n23754 & ~n23756;
  assign n23768 = n22625 & n23767;
  assign n23769 = ~n23754 & n23766;
  assign n23770 = pi19  & ~n23742;
  assign n23771 = ~n35387 & ~n23770;
  assign n23772 = ~n35390 & n23771;
  assign n23773 = ~n22625 & ~n23767;
  assign n23774 = n21842 & ~n23773;
  assign n23775 = ~n23772 & ~n23773;
  assign n23776 = n21842 & n23775;
  assign n23777 = ~n23772 & n23774;
  assign n23778 = ~n23753 & ~n35391;
  assign n23779 = ~n21842 & ~n23775;
  assign n23780 = n20986 & ~n23779;
  assign n23781 = ~n23778 & n23780;
  assign n23782 = ~n22642 & ~n35239;
  assign n23783 = ~n23517 & n23782;
  assign n23784 = n22647 & ~n23783;
  assign n23785 = ~n22647 & n23782;
  assign n23786 = ~n22647 & n23783;
  assign n23787 = ~n23517 & n23785;
  assign n23788 = ~n23784 & ~n35392;
  assign n23789 = ~n23781 & ~n23788;
  assign n23790 = ~n23778 & ~n23779;
  assign n23791 = ~n20986 & ~n23790;
  assign n23792 = n20229 & ~n23791;
  assign n23793 = ~n23789 & ~n23791;
  assign n23794 = n20229 & n23793;
  assign n23795 = ~n23789 & n23792;
  assign n23796 = ~n23741 & ~n35393;
  assign n23797 = ~n20229 & ~n23793;
  assign n23798 = n19401 & ~n23797;
  assign n23799 = ~n23796 & n23798;
  assign n23800 = ~n22676 & ~n35241;
  assign n23801 = ~n23517 & n23800;
  assign n23802 = n22686 & ~n23801;
  assign n23803 = ~n22686 & n23801;
  assign n23804 = ~n22676 & n22686;
  assign n23805 = ~n35241 & n23804;
  assign n23806 = n22686 & n23801;
  assign n23807 = ~n23517 & n23805;
  assign n23808 = ~n22686 & ~n23801;
  assign n23809 = ~n35394 & ~n23808;
  assign n23810 = ~n23802 & ~n23803;
  assign n23811 = ~n23799 & ~n35395;
  assign n23812 = ~n23796 & ~n23797;
  assign n23813 = ~n19401 & ~n23812;
  assign n23814 = n18676 & ~n23813;
  assign n23815 = ~n23811 & ~n23813;
  assign n23816 = n18676 & n23815;
  assign n23817 = ~n23811 & n23814;
  assign n23818 = ~n23733 & ~n35396;
  assign n23819 = ~n18676 & ~n23815;
  assign n23820 = n17885 & ~n23819;
  assign n23821 = ~n23818 & n23820;
  assign n23822 = ~n22706 & ~n35245;
  assign n23823 = ~n23517 & n23822;
  assign n23824 = ~n35247 & n23823;
  assign n23825 = n35247 & ~n23823;
  assign n23826 = ~n22706 & n35247;
  assign n23827 = ~n35245 & n23826;
  assign n23828 = ~n23517 & n23827;
  assign n23829 = ~n35247 & ~n23823;
  assign n23830 = ~n23828 & ~n23829;
  assign n23831 = ~n23824 & ~n23825;
  assign n23832 = ~n23821 & ~n35397;
  assign n23833 = ~n23818 & ~n23819;
  assign n23834 = ~n17885 & ~n23833;
  assign n23835 = n17187 & ~n23834;
  assign n23836 = ~n23832 & ~n23834;
  assign n23837 = n17187 & n23836;
  assign n23838 = ~n23832 & n23835;
  assign n23839 = ~n23725 & ~n35398;
  assign n23840 = ~n17187 & ~n23836;
  assign n23841 = n16428 & ~n23840;
  assign n23842 = ~n23839 & n23841;
  assign n23843 = ~n22740 & ~n35250;
  assign n23844 = ~n23517 & n23843;
  assign n23845 = ~n35251 & ~n23844;
  assign n23846 = ~n22740 & n35251;
  assign n23847 = ~n35250 & n23846;
  assign n23848 = n35251 & n23844;
  assign n23849 = ~n23517 & n23847;
  assign n23850 = n35251 & ~n23844;
  assign n23851 = ~n35251 & n23844;
  assign n23852 = ~n23850 & ~n23851;
  assign n23853 = ~n23845 & ~n35399;
  assign n23854 = ~n23842 & n35400;
  assign n23855 = ~n23839 & ~n23840;
  assign n23856 = ~n16428 & ~n23855;
  assign n23857 = n15760 & ~n23856;
  assign n23858 = ~n23854 & ~n23856;
  assign n23859 = n15760 & n23858;
  assign n23860 = ~n23854 & n23857;
  assign n23861 = ~n23717 & ~n35401;
  assign n23862 = ~n15760 & ~n23858;
  assign n23863 = n15033 & ~n23862;
  assign n23864 = ~n23861 & n23863;
  assign n23865 = ~n22773 & ~n35254;
  assign n23866 = ~n23517 & n23865;
  assign n23867 = n35256 & ~n23866;
  assign n23868 = ~n22773 & ~n35256;
  assign n23869 = ~n35254 & n23868;
  assign n23870 = ~n35256 & n23866;
  assign n23871 = ~n23517 & n23869;
  assign n23872 = n35256 & n23866;
  assign n23873 = ~n35256 & ~n23866;
  assign n23874 = ~n23872 & ~n23873;
  assign n23875 = ~n23867 & ~n35402;
  assign n23876 = ~n23864 & n35403;
  assign n23877 = ~n23861 & ~n23862;
  assign n23878 = ~n15033 & ~n23877;
  assign n23879 = n14394 & ~n23878;
  assign n23880 = ~n23876 & ~n23878;
  assign n23881 = n14394 & n23880;
  assign n23882 = ~n23876 & n23879;
  assign n23883 = ~n23709 & ~n35404;
  assign n23884 = ~n14394 & ~n23880;
  assign n23885 = n13704 & ~n23884;
  assign n23886 = ~n23883 & n23885;
  assign n23887 = ~n22807 & ~n35259;
  assign n23888 = ~n22807 & ~n23517;
  assign n23889 = ~n35259 & n23888;
  assign n23890 = ~n23517 & n23887;
  assign n23891 = ~n35261 & ~n35405;
  assign n23892 = n22822 & n23888;
  assign n23893 = n35261 & n35405;
  assign n23894 = ~n22807 & ~n35261;
  assign n23895 = ~n35259 & n23894;
  assign n23896 = ~n23517 & n23895;
  assign n23897 = n35261 & ~n35405;
  assign n23898 = ~n23896 & ~n23897;
  assign n23899 = ~n23891 & ~n35406;
  assign n23900 = ~n23886 & ~n35407;
  assign n23901 = ~n23883 & ~n23884;
  assign n23902 = ~n13704 & ~n23901;
  assign n23903 = n13099 & ~n23902;
  assign n23904 = ~n23900 & ~n23902;
  assign n23905 = n13099 & n23904;
  assign n23906 = ~n23900 & n23903;
  assign n23907 = ~n23701 & ~n35408;
  assign n23908 = ~n13099 & ~n23904;
  assign n23909 = n12442 & ~n23908;
  assign n23910 = ~n23907 & n23909;
  assign n23911 = ~n22841 & ~n35264;
  assign n23912 = ~n23517 & n23911;
  assign n23913 = ~n35267 & ~n23912;
  assign n23914 = ~n22841 & n35267;
  assign n23915 = ~n35264 & n23914;
  assign n23916 = n35267 & n23912;
  assign n23917 = ~n23517 & n23915;
  assign n23918 = ~n23913 & ~n35409;
  assign n23919 = ~n23910 & ~n23918;
  assign n23920 = ~n23907 & ~n23908;
  assign n23921 = ~n12442 & ~n23920;
  assign n23922 = n11858 & ~n23921;
  assign n23923 = ~n23919 & ~n23921;
  assign n23924 = n11858 & n23923;
  assign n23925 = ~n23919 & n23922;
  assign n23926 = ~n23693 & ~n35410;
  assign n23927 = ~n11858 & ~n23923;
  assign n23928 = n11229 & ~n23927;
  assign n23929 = ~n23926 & n23928;
  assign n23930 = ~n22877 & ~n35270;
  assign n23931 = ~n22877 & ~n23517;
  assign n23932 = ~n35270 & n23931;
  assign n23933 = ~n23517 & n23930;
  assign n23934 = n22888 & ~n35411;
  assign n23935 = n22889 & n23931;
  assign n23936 = ~n22888 & n35411;
  assign n23937 = ~n22877 & n22888;
  assign n23938 = ~n35270 & n23937;
  assign n23939 = ~n23517 & n23938;
  assign n23940 = ~n22888 & ~n35411;
  assign n23941 = ~n23939 & ~n23940;
  assign n23942 = ~n23934 & ~n35412;
  assign n23943 = ~n23929 & ~n35413;
  assign n23944 = ~n23926 & ~n23927;
  assign n23945 = ~n11229 & ~n23944;
  assign n23946 = n10681 & ~n23945;
  assign n23947 = ~n23943 & ~n23945;
  assign n23948 = n10681 & n23947;
  assign n23949 = ~n23943 & n23946;
  assign n23950 = ~n23685 & ~n35414;
  assign n23951 = ~n10681 & ~n23947;
  assign n23952 = n10086 & ~n23951;
  assign n23953 = ~n23950 & n23952;
  assign n23954 = ~n22908 & ~n35274;
  assign n23955 = ~n23517 & n23954;
  assign n23956 = ~n35277 & n23955;
  assign n23957 = n35277 & ~n23955;
  assign n23958 = ~n22908 & n35277;
  assign n23959 = ~n35274 & n23958;
  assign n23960 = n35277 & n23955;
  assign n23961 = ~n23517 & n23959;
  assign n23962 = ~n35277 & ~n23955;
  assign n23963 = ~n35415 & ~n23962;
  assign n23964 = ~n23956 & ~n23957;
  assign n23965 = ~n23953 & ~n35416;
  assign n23966 = ~n23950 & ~n23951;
  assign n23967 = ~n10086 & ~n23966;
  assign n23968 = n9565 & ~n23967;
  assign n23969 = ~n23965 & ~n23967;
  assign n23970 = n9565 & n23969;
  assign n23971 = ~n23965 & n23968;
  assign n23972 = ~n23677 & ~n35417;
  assign n23973 = ~n9565 & ~n23969;
  assign n23974 = n8998 & ~n23973;
  assign n23975 = ~n23972 & n23974;
  assign n23976 = ~n22944 & ~n35280;
  assign n23977 = ~n22944 & ~n23517;
  assign n23978 = ~n35280 & n23977;
  assign n23979 = ~n23517 & n23976;
  assign n23980 = n35282 & ~n35418;
  assign n23981 = n22959 & n23977;
  assign n23982 = ~n35282 & n35418;
  assign n23983 = ~n22944 & n35282;
  assign n23984 = ~n35280 & n23983;
  assign n23985 = ~n23517 & n23984;
  assign n23986 = ~n35282 & ~n35418;
  assign n23987 = ~n23985 & ~n23986;
  assign n23988 = ~n23980 & ~n35419;
  assign n23989 = ~n23975 & ~n35420;
  assign n23990 = ~n23972 & ~n23973;
  assign n23991 = ~n8998 & ~n23990;
  assign n23992 = n8506 & ~n23991;
  assign n23993 = ~n23989 & ~n23991;
  assign n23994 = n8506 & n23993;
  assign n23995 = ~n23989 & n23992;
  assign n23996 = ~n23669 & ~n35421;
  assign n23997 = ~n8506 & ~n23993;
  assign n23998 = n7975 & ~n23997;
  assign n23999 = ~n23996 & n23998;
  assign n24000 = ~n23661 & ~n23999;
  assign n24001 = ~n23996 & ~n23997;
  assign n24002 = ~n7975 & ~n24001;
  assign n24003 = n7512 & ~n24002;
  assign n24004 = ~n24000 & ~n24002;
  assign n24005 = n7512 & n24004;
  assign n24006 = ~n24000 & n24003;
  assign n24007 = ~n23653 & ~n35422;
  assign n24008 = ~n7512 & ~n24004;
  assign n24009 = n7015 & ~n24008;
  assign n24010 = ~n24007 & n24009;
  assign n24011 = ~n23014 & ~n35292;
  assign n24012 = ~n23014 & ~n23517;
  assign n24013 = ~n35292 & n24012;
  assign n24014 = ~n23517 & n24011;
  assign n24015 = n23022 & ~n35423;
  assign n24016 = n23026 & n24012;
  assign n24017 = ~n23014 & n23022;
  assign n24018 = ~n35292 & n24017;
  assign n24019 = ~n23517 & n24018;
  assign n24020 = ~n23022 & ~n35423;
  assign n24021 = ~n24019 & ~n24020;
  assign n24022 = ~n24015 & ~n24016;
  assign n24023 = ~n24010 & ~n35424;
  assign n24024 = ~n24007 & ~n24008;
  assign n24025 = ~n7015 & ~n24024;
  assign n24026 = n6579 & ~n24025;
  assign n24027 = ~n24023 & ~n24025;
  assign n24028 = n6579 & n24027;
  assign n24029 = ~n24023 & n24026;
  assign n24030 = ~n23645 & ~n35425;
  assign n24031 = ~n6579 & ~n24027;
  assign n24032 = n6117 & ~n24031;
  assign n24033 = ~n24030 & n24032;
  assign n24034 = ~n23637 & ~n24033;
  assign n24035 = ~n24030 & ~n24031;
  assign n24036 = ~n6117 & ~n24035;
  assign n24037 = n5708 & ~n24036;
  assign n24038 = ~n24034 & ~n24036;
  assign n24039 = n5708 & n24038;
  assign n24040 = ~n24034 & n24037;
  assign n24041 = ~n23629 & ~n35426;
  assign n24042 = ~n5708 & ~n24038;
  assign n24043 = n5278 & ~n24042;
  assign n24044 = ~n24041 & n24043;
  assign n24045 = ~n23080 & ~n35301;
  assign n24046 = ~n23080 & ~n23517;
  assign n24047 = ~n35301 & n24046;
  assign n24048 = ~n23517 & n24045;
  assign n24049 = n23088 & ~n35427;
  assign n24050 = n23092 & n24046;
  assign n24051 = ~n23080 & n23088;
  assign n24052 = ~n35301 & n24051;
  assign n24053 = ~n23517 & n24052;
  assign n24054 = ~n23088 & ~n35427;
  assign n24055 = ~n24053 & ~n24054;
  assign n24056 = ~n24049 & ~n24050;
  assign n24057 = ~n24044 & ~n35428;
  assign n24058 = ~n24041 & ~n24042;
  assign n24059 = ~n5278 & ~n24058;
  assign n24060 = n4903 & ~n24059;
  assign n24061 = ~n24057 & ~n24059;
  assign n24062 = n4903 & n24061;
  assign n24063 = ~n24057 & n24060;
  assign n24064 = ~n23621 & ~n35429;
  assign n24065 = ~n4903 & ~n24061;
  assign n24066 = n4508 & ~n24065;
  assign n24067 = ~n24064 & n24066;
  assign n24068 = ~n23613 & ~n24067;
  assign n24069 = ~n24064 & ~n24065;
  assign n24070 = ~n4508 & ~n24069;
  assign n24071 = n4155 & ~n24070;
  assign n24072 = ~n24068 & ~n24070;
  assign n24073 = n4155 & n24072;
  assign n24074 = ~n24068 & n24071;
  assign n24075 = ~n23605 & ~n35430;
  assign n24076 = ~n4155 & ~n24072;
  assign n24077 = n3788 & ~n24076;
  assign n24078 = ~n24075 & n24077;
  assign n24079 = ~n23146 & ~n35310;
  assign n24080 = ~n23146 & ~n23517;
  assign n24081 = ~n35310 & n24080;
  assign n24082 = ~n23517 & n24079;
  assign n24083 = n23154 & ~n35431;
  assign n24084 = n23158 & n24080;
  assign n24085 = ~n23146 & n23154;
  assign n24086 = ~n35310 & n24085;
  assign n24087 = ~n23517 & n24086;
  assign n24088 = ~n23154 & ~n35431;
  assign n24089 = ~n24087 & ~n24088;
  assign n24090 = ~n24083 & ~n24084;
  assign n24091 = ~n24078 & ~n35432;
  assign n24092 = ~n24075 & ~n24076;
  assign n24093 = ~n3788 & ~n24092;
  assign n24094 = n3473 & ~n24093;
  assign n24095 = ~n24091 & ~n24093;
  assign n24096 = n3473 & n24095;
  assign n24097 = ~n24091 & n24094;
  assign n24098 = ~n23597 & ~n35433;
  assign n24099 = ~n3473 & ~n24095;
  assign n24100 = n3140 & ~n24099;
  assign n24101 = ~n24098 & n24100;
  assign n24102 = ~n23589 & ~n24101;
  assign n24103 = ~n24098 & ~n24099;
  assign n24104 = ~n3140 & ~n24103;
  assign n24105 = n2855 & ~n24104;
  assign n24106 = ~n24102 & ~n24104;
  assign n24107 = n2855 & n24106;
  assign n24108 = ~n24102 & n24105;
  assign n24109 = ~n23581 & ~n35434;
  assign n24110 = ~n2855 & ~n24106;
  assign n24111 = n2556 & ~n24110;
  assign n24112 = ~n24109 & n24111;
  assign n24113 = ~n23212 & ~n35319;
  assign n24114 = ~n23212 & ~n23517;
  assign n24115 = ~n35319 & n24114;
  assign n24116 = ~n23517 & n24113;
  assign n24117 = n23220 & ~n35435;
  assign n24118 = n23224 & n24114;
  assign n24119 = ~n23212 & n23220;
  assign n24120 = ~n35319 & n24119;
  assign n24121 = ~n23517 & n24120;
  assign n24122 = ~n23220 & ~n35435;
  assign n24123 = ~n24121 & ~n24122;
  assign n24124 = ~n24117 & ~n24118;
  assign n24125 = ~n24112 & ~n35436;
  assign n24126 = ~n24109 & ~n24110;
  assign n24127 = ~n2556 & ~n24126;
  assign n24128 = n2301 & ~n24127;
  assign n24129 = ~n24125 & ~n24127;
  assign n24130 = n2301 & n24129;
  assign n24131 = ~n24125 & n24128;
  assign n24132 = ~n23573 & ~n35437;
  assign n24133 = ~n2301 & ~n24129;
  assign n24134 = n2038 & ~n24133;
  assign n24135 = ~n24132 & n24134;
  assign n24136 = ~n23565 & ~n24135;
  assign n24137 = ~n24132 & ~n24133;
  assign n24138 = ~n2038 & ~n24137;
  assign n24139 = n1812 & ~n24138;
  assign n24140 = ~n24136 & ~n24138;
  assign n24141 = n1812 & n24140;
  assign n24142 = ~n24136 & n24139;
  assign n24143 = ~n23557 & ~n35438;
  assign n24144 = ~n1812 & ~n24140;
  assign n24145 = n1582 & ~n24144;
  assign n24146 = ~n24143 & n24145;
  assign n24147 = ~n23278 & ~n35328;
  assign n24148 = ~n23278 & ~n23517;
  assign n24149 = ~n35328 & n24148;
  assign n24150 = ~n23517 & n24147;
  assign n24151 = n23286 & ~n35439;
  assign n24152 = n23290 & n24148;
  assign n24153 = ~n23278 & n23286;
  assign n24154 = ~n35328 & n24153;
  assign n24155 = ~n23517 & n24154;
  assign n24156 = ~n23286 & ~n35439;
  assign n24157 = ~n24155 & ~n24156;
  assign n24158 = ~n24151 & ~n24152;
  assign n24159 = ~n24146 & ~n35440;
  assign n24160 = ~n24143 & ~n24144;
  assign n24161 = ~n1582 & ~n24160;
  assign n24162 = n1388 & ~n24161;
  assign n24163 = ~n24159 & ~n24161;
  assign n24164 = n1388 & n24163;
  assign n24165 = ~n24159 & n24162;
  assign n24166 = ~n23549 & ~n35441;
  assign n24167 = ~n1388 & ~n24163;
  assign n24168 = n1192 & ~n24167;
  assign n24169 = ~n24166 & n24168;
  assign n24170 = ~n23541 & ~n24169;
  assign n24171 = ~n24166 & ~n24167;
  assign n24172 = ~n1192 & ~n24171;
  assign n24173 = n1028 & ~n24172;
  assign n24174 = ~n24170 & ~n24172;
  assign n24175 = n1028 & n24174;
  assign n24176 = ~n24170 & n24173;
  assign n24177 = ~n23533 & ~n35442;
  assign n24178 = ~n1028 & ~n24174;
  assign n24179 = ~n24177 & ~n24178;
  assign n24180 = ~n866 & ~n24179;
  assign n24181 = n866 & ~n24178;
  assign n24182 = ~n24177 & n24181;
  assign n24183 = ~n23340 & ~n35335;
  assign n24184 = ~n23517 & n24183;
  assign n24185 = ~n35337 & ~n24184;
  assign n24186 = ~n23340 & n35337;
  assign n24187 = ~n35335 & n24186;
  assign n24188 = n35337 & n24184;
  assign n24189 = ~n23517 & n24187;
  assign n24190 = n35337 & ~n24184;
  assign n24191 = ~n35337 & n24184;
  assign n24192 = ~n24190 & ~n24191;
  assign n24193 = ~n24185 & ~n35443;
  assign n24194 = ~n24182 & n35444;
  assign n24195 = ~n24180 & ~n24194;
  assign n24196 = ~n730 & ~n24195;
  assign n24197 = n730 & ~n24180;
  assign n24198 = n730 & n24195;
  assign n24199 = ~n24194 & n24197;
  assign n24200 = ~n23525 & ~n35445;
  assign n24201 = ~n24196 & ~n24200;
  assign n24202 = ~n602 & ~n24201;
  assign n24203 = n602 & ~n24196;
  assign n24204 = ~n24200 & n24203;
  assign n24205 = ~n23362 & ~n35339;
  assign n24206 = ~n23362 & ~n23517;
  assign n24207 = ~n35339 & n24206;
  assign n24208 = ~n23517 & n24205;
  assign n24209 = n23370 & ~n35446;
  assign n24210 = n23374 & n24206;
  assign n24211 = ~n23362 & n23370;
  assign n24212 = ~n35339 & n24211;
  assign n24213 = ~n23517 & n24212;
  assign n24214 = ~n23370 & ~n35446;
  assign n24215 = ~n24213 & ~n24214;
  assign n24216 = ~n24209 & ~n24210;
  assign n24217 = ~n24204 & ~n35447;
  assign n24218 = ~n24202 & ~n24217;
  assign n24219 = ~n497 & ~n24218;
  assign n24220 = ~n23376 & ~n23378;
  assign n24221 = ~n23517 & n24220;
  assign n24222 = ~n35341 & ~n24221;
  assign n24223 = ~n23378 & n35341;
  assign n24224 = ~n23376 & n24223;
  assign n24225 = n35341 & n24221;
  assign n24226 = ~n23517 & n24224;
  assign n24227 = ~n24222 & ~n35448;
  assign n24228 = n497 & ~n24202;
  assign n24229 = n497 & n24218;
  assign n24230 = ~n24217 & n24228;
  assign n24231 = ~n24227 & ~n35449;
  assign n24232 = ~n24219 & ~n24231;
  assign n24233 = ~n403 & ~n24232;
  assign n24234 = n403 & ~n24219;
  assign n24235 = ~n24231 & n24234;
  assign n24236 = ~n23393 & ~n35343;
  assign n24237 = ~n23393 & ~n23517;
  assign n24238 = ~n35343 & n24237;
  assign n24239 = ~n23517 & n24236;
  assign n24240 = n23401 & ~n35450;
  assign n24241 = n23405 & n24237;
  assign n24242 = ~n23393 & n23401;
  assign n24243 = ~n35343 & n24242;
  assign n24244 = ~n23517 & n24243;
  assign n24245 = ~n23401 & ~n35450;
  assign n24246 = ~n24244 & ~n24245;
  assign n24247 = ~n24240 & ~n24241;
  assign n24248 = ~n24235 & ~n35451;
  assign n24249 = ~n24233 & ~n24248;
  assign n24250 = ~n330 & ~n24249;
  assign n24251 = ~n23407 & ~n23409;
  assign n24252 = ~n23517 & n24251;
  assign n24253 = ~n35345 & ~n24252;
  assign n24254 = ~n23409 & n35345;
  assign n24255 = ~n23407 & n24254;
  assign n24256 = n35345 & n24252;
  assign n24257 = ~n23517 & n24255;
  assign n24258 = ~n24253 & ~n35452;
  assign n24259 = n330 & ~n24233;
  assign n24260 = n330 & n24249;
  assign n24261 = ~n24248 & n24259;
  assign n24262 = ~n24258 & ~n35453;
  assign n24263 = ~n24250 & ~n24262;
  assign n24264 = ~n271 & ~n24263;
  assign n24265 = ~n23424 & ~n35346;
  assign n24266 = ~n23517 & n24265;
  assign n24267 = ~n35348 & ~n24266;
  assign n24268 = ~n23424 & n35348;
  assign n24269 = ~n35346 & n24268;
  assign n24270 = n35348 & n24266;
  assign n24271 = ~n23517 & n24269;
  assign n24272 = ~n24267 & ~n35454;
  assign n24273 = n271 & ~n24250;
  assign n24274 = ~n24262 & n24273;
  assign n24275 = ~n24272 & ~n24274;
  assign n24276 = ~n24264 & ~n24275;
  assign n24277 = ~n217 & ~n24276;
  assign n24278 = ~n23442 & ~n23444;
  assign n24279 = ~n23517 & n24278;
  assign n24280 = ~n35350 & ~n24279;
  assign n24281 = ~n23444 & n35350;
  assign n24282 = ~n23442 & n24281;
  assign n24283 = n35350 & n24279;
  assign n24284 = ~n23517 & n24282;
  assign n24285 = ~n24280 & ~n35455;
  assign n24286 = n217 & ~n24264;
  assign n24287 = n217 & n24276;
  assign n24288 = ~n24275 & n24286;
  assign n24289 = ~n24285 & ~n35456;
  assign n24290 = ~n24277 & ~n24289;
  assign n24291 = ~n198 & ~n24290;
  assign n24292 = n198 & ~n24277;
  assign n24293 = ~n24289 & n24292;
  assign n24294 = ~n23459 & ~n35352;
  assign n24295 = ~n23459 & ~n23517;
  assign n24296 = ~n35352 & n24295;
  assign n24297 = ~n23517 & n24294;
  assign n24298 = n23467 & ~n35457;
  assign n24299 = n23471 & n24295;
  assign n24300 = ~n23459 & n23467;
  assign n24301 = ~n35352 & n24300;
  assign n24302 = ~n23517 & n24301;
  assign n24303 = ~n23467 & ~n35457;
  assign n24304 = ~n24302 & ~n24303;
  assign n24305 = ~n24298 & ~n24299;
  assign n24306 = ~n24293 & ~n35458;
  assign n24307 = ~n24291 & ~n24306;
  assign n24308 = ~n23473 & ~n23475;
  assign n24309 = ~n23517 & n24308;
  assign n24310 = ~n35354 & ~n24309;
  assign n24311 = ~n23475 & n35354;
  assign n24312 = ~n23473 & n24311;
  assign n24313 = n35354 & n24309;
  assign n24314 = ~n23517 & n24312;
  assign n24315 = ~n24310 & ~n35459;
  assign n24316 = ~n23489 & ~n35356;
  assign n24317 = ~n35356 & ~n23517;
  assign n24318 = ~n23489 & n24317;
  assign n24319 = ~n23517 & n24316;
  assign n24320 = ~n35358 & ~n35460;
  assign n24321 = ~n24315 & n24320;
  assign n24322 = ~n24307 & n24321;
  assign n24323 = n193 & ~n24322;
  assign n24324 = ~n24291 & n24315;
  assign n24325 = n24307 & n24315;
  assign n24326 = ~n24306 & n24324;
  assign n24327 = n23489 & ~n24317;
  assign n24328 = ~n193 & ~n24316;
  assign n24329 = ~n24327 & n24328;
  assign n24330 = ~n35461 & ~n24329;
  assign n24331 = ~n24323 & n24330;
  assign n24332 = ~n24196 & ~n35445;
  assign n24333 = ~n24196 & ~n24331;
  assign n24334 = ~n35445 & n24333;
  assign n24335 = ~n24331 & n24332;
  assign n24336 = n23525 & ~n35462;
  assign n24337 = n24200 & n24333;
  assign n24338 = n23525 & ~n35445;
  assign n24339 = ~n24196 & n24338;
  assign n24340 = ~n24331 & n24339;
  assign n24341 = ~n23525 & ~n35462;
  assign n24342 = ~n24340 & ~n24341;
  assign n24343 = ~n24336 & ~n24337;
  assign n24344 = pi16  & ~n24331;
  assign n24345 = ~pi14  & ~pi15 ;
  assign n24346 = ~pi16  & n24345;
  assign n24347 = ~n24344 & ~n24346;
  assign n24348 = ~n23517 & ~n24347;
  assign n24349 = ~pi16  & ~n24331;
  assign n24350 = pi17  & ~n24349;
  assign n24351 = ~pi17  & n24349;
  assign n24352 = n23755 & ~n24331;
  assign n24353 = ~n24350 & ~n35464;
  assign n24354 = ~n35232 & ~n35389;
  assign n24355 = ~n22604 & n24354;
  assign n24356 = ~n22623 & n24355;
  assign n24357 = ~n35234 & n24356;
  assign n24358 = n22609 & n22625;
  assign n24359 = ~n22617 & n24357;
  assign n24360 = ~n24346 & ~n35465;
  assign n24361 = ~n23515 & n24360;
  assign n24362 = ~n35358 & n24361;
  assign n24363 = ~n23509 & n24362;
  assign n24364 = n23517 & n24347;
  assign n24365 = ~n24344 & n24363;
  assign n24366 = n24353 & ~n35466;
  assign n24367 = ~n24348 & ~n24366;
  assign n24368 = ~n22625 & ~n24367;
  assign n24369 = n22625 & ~n24348;
  assign n24370 = ~n24366 & n24369;
  assign n24371 = ~n23517 & ~n24329;
  assign n24372 = ~n35461 & n24371;
  assign n24373 = ~n24323 & n24372;
  assign n24374 = ~n35464 & ~n24373;
  assign n24375 = pi18  & ~n24374;
  assign n24376 = ~pi18  & ~n24373;
  assign n24377 = ~pi18  & n24374;
  assign n24378 = ~n35464 & n24376;
  assign n24379 = ~n24375 & ~n35467;
  assign n24380 = ~n24370 & ~n24379;
  assign n24381 = ~n24368 & ~n24380;
  assign n24382 = ~n21842 & ~n24381;
  assign n24383 = n21842 & ~n24368;
  assign n24384 = ~n24380 & n24383;
  assign n24385 = n21842 & n24381;
  assign n24386 = ~n35390 & ~n23773;
  assign n24387 = ~n24331 & n24386;
  assign n24388 = n23771 & ~n24387;
  assign n24389 = ~n23771 & n24386;
  assign n24390 = ~n23771 & n24387;
  assign n24391 = ~n24331 & n24389;
  assign n24392 = ~n24388 & ~n35469;
  assign n24393 = ~n35468 & ~n24392;
  assign n24394 = ~n24382 & ~n24393;
  assign n24395 = ~n20986 & ~n24394;
  assign n24396 = n20986 & ~n24382;
  assign n24397 = ~n24393 & n24396;
  assign n24398 = ~n35391 & ~n23779;
  assign n24399 = ~n23779 & ~n24331;
  assign n24400 = ~n35391 & n24399;
  assign n24401 = ~n24331 & n24398;
  assign n24402 = n23753 & ~n35470;
  assign n24403 = n23778 & n24399;
  assign n24404 = n23753 & ~n35391;
  assign n24405 = ~n23779 & n24404;
  assign n24406 = ~n24331 & n24405;
  assign n24407 = ~n23753 & ~n35470;
  assign n24408 = ~n24406 & ~n24407;
  assign n24409 = ~n24402 & ~n24403;
  assign n24410 = ~n24397 & ~n35471;
  assign n24411 = ~n24395 & ~n24410;
  assign n24412 = ~n20229 & ~n24411;
  assign n24413 = n20229 & ~n24395;
  assign n24414 = ~n24410 & n24413;
  assign n24415 = n20229 & n24411;
  assign n24416 = ~n23781 & ~n23791;
  assign n24417 = ~n24331 & n24416;
  assign n24418 = n23788 & ~n24417;
  assign n24419 = ~n23788 & n24417;
  assign n24420 = n23788 & ~n23791;
  assign n24421 = ~n23781 & n24420;
  assign n24422 = n23788 & n24417;
  assign n24423 = ~n24331 & n24421;
  assign n24424 = ~n23788 & ~n24417;
  assign n24425 = ~n35473 & ~n24424;
  assign n24426 = ~n24418 & ~n24419;
  assign n24427 = ~n35472 & ~n35474;
  assign n24428 = ~n24412 & ~n24427;
  assign n24429 = ~n19401 & ~n24428;
  assign n24430 = n19401 & ~n24412;
  assign n24431 = ~n24427 & n24430;
  assign n24432 = ~n35393 & ~n23797;
  assign n24433 = ~n23797 & ~n24331;
  assign n24434 = ~n35393 & n24433;
  assign n24435 = ~n24331 & n24432;
  assign n24436 = n23741 & ~n35475;
  assign n24437 = n23796 & n24433;
  assign n24438 = n23741 & ~n35393;
  assign n24439 = ~n23797 & n24438;
  assign n24440 = ~n24331 & n24439;
  assign n24441 = ~n23741 & ~n35475;
  assign n24442 = ~n24440 & ~n24441;
  assign n24443 = ~n24436 & ~n24437;
  assign n24444 = ~n24431 & ~n35476;
  assign n24445 = ~n24429 & ~n24444;
  assign n24446 = ~n18676 & ~n24445;
  assign n24447 = n18676 & ~n24429;
  assign n24448 = ~n24444 & n24447;
  assign n24449 = n18676 & n24445;
  assign n24450 = ~n23799 & ~n23813;
  assign n24451 = ~n24331 & n24450;
  assign n24452 = ~n35395 & n24451;
  assign n24453 = n35395 & ~n24451;
  assign n24454 = n35395 & ~n23813;
  assign n24455 = ~n23799 & n24454;
  assign n24456 = ~n24331 & n24455;
  assign n24457 = ~n35395 & ~n24451;
  assign n24458 = ~n24456 & ~n24457;
  assign n24459 = ~n24452 & ~n24453;
  assign n24460 = ~n35477 & ~n35478;
  assign n24461 = ~n24446 & ~n24460;
  assign n24462 = ~n17885 & ~n24461;
  assign n24463 = n17885 & ~n24446;
  assign n24464 = ~n24460 & n24463;
  assign n24465 = ~n35396 & ~n23819;
  assign n24466 = ~n23819 & ~n24331;
  assign n24467 = ~n35396 & n24466;
  assign n24468 = ~n24331 & n24465;
  assign n24469 = n23733 & ~n35479;
  assign n24470 = n23818 & n24466;
  assign n24471 = n23733 & ~n35396;
  assign n24472 = ~n23819 & n24471;
  assign n24473 = ~n24331 & n24472;
  assign n24474 = ~n23733 & ~n35479;
  assign n24475 = ~n24473 & ~n24474;
  assign n24476 = ~n24469 & ~n24470;
  assign n24477 = ~n24464 & ~n35480;
  assign n24478 = ~n24462 & ~n24477;
  assign n24479 = ~n17187 & ~n24478;
  assign n24480 = n17187 & ~n24462;
  assign n24481 = ~n24477 & n24480;
  assign n24482 = n17187 & n24478;
  assign n24483 = ~n23821 & ~n23834;
  assign n24484 = ~n24331 & n24483;
  assign n24485 = ~n35397 & ~n24484;
  assign n24486 = n35397 & ~n23834;
  assign n24487 = ~n23821 & n24486;
  assign n24488 = n35397 & n24484;
  assign n24489 = ~n24331 & n24487;
  assign n24490 = n35397 & ~n24484;
  assign n24491 = ~n35397 & n24484;
  assign n24492 = ~n24490 & ~n24491;
  assign n24493 = ~n24485 & ~n35482;
  assign n24494 = ~n35481 & n35483;
  assign n24495 = ~n24479 & ~n24494;
  assign n24496 = ~n16428 & ~n24495;
  assign n24497 = n16428 & ~n24479;
  assign n24498 = ~n24494 & n24497;
  assign n24499 = ~n35398 & ~n23840;
  assign n24500 = ~n23840 & ~n24331;
  assign n24501 = ~n35398 & n24500;
  assign n24502 = ~n24331 & n24499;
  assign n24503 = n23725 & ~n35484;
  assign n24504 = n23839 & n24500;
  assign n24505 = n23725 & ~n35398;
  assign n24506 = ~n23840 & n24505;
  assign n24507 = ~n24331 & n24506;
  assign n24508 = ~n23725 & ~n35484;
  assign n24509 = ~n24507 & ~n24508;
  assign n24510 = ~n24503 & ~n24504;
  assign n24511 = ~n24498 & ~n35485;
  assign n24512 = ~n24496 & ~n24511;
  assign n24513 = ~n15760 & ~n24512;
  assign n24514 = n15760 & ~n24496;
  assign n24515 = ~n24511 & n24514;
  assign n24516 = n15760 & n24512;
  assign n24517 = ~n23842 & ~n23856;
  assign n24518 = ~n24331 & n24517;
  assign n24519 = n35400 & ~n24518;
  assign n24520 = ~n35400 & ~n23856;
  assign n24521 = ~n23842 & n24520;
  assign n24522 = ~n35400 & n24518;
  assign n24523 = ~n24331 & n24521;
  assign n24524 = n35400 & n24518;
  assign n24525 = ~n35400 & ~n24518;
  assign n24526 = ~n24524 & ~n24525;
  assign n24527 = ~n24519 & ~n35487;
  assign n24528 = ~n35486 & n35488;
  assign n24529 = ~n24513 & ~n24528;
  assign n24530 = ~n15033 & ~n24529;
  assign n24531 = n15033 & ~n24513;
  assign n24532 = ~n24528 & n24531;
  assign n24533 = ~n35401 & ~n23862;
  assign n24534 = ~n23862 & ~n24331;
  assign n24535 = ~n35401 & n24534;
  assign n24536 = ~n24331 & n24533;
  assign n24537 = n23717 & ~n35489;
  assign n24538 = n23861 & n24534;
  assign n24539 = n23717 & ~n35401;
  assign n24540 = ~n23862 & n24539;
  assign n24541 = ~n24331 & n24540;
  assign n24542 = ~n23717 & ~n35489;
  assign n24543 = ~n24541 & ~n24542;
  assign n24544 = ~n24537 & ~n24538;
  assign n24545 = ~n24532 & ~n35490;
  assign n24546 = ~n24530 & ~n24545;
  assign n24547 = ~n14394 & ~n24546;
  assign n24548 = n14394 & ~n24530;
  assign n24549 = ~n24545 & n24548;
  assign n24550 = n14394 & n24546;
  assign n24551 = ~n23864 & ~n23878;
  assign n24552 = ~n23878 & ~n24331;
  assign n24553 = ~n23864 & n24552;
  assign n24554 = ~n24331 & n24551;
  assign n24555 = ~n35403 & ~n35492;
  assign n24556 = n23876 & n24552;
  assign n24557 = n35403 & n35492;
  assign n24558 = ~n35403 & ~n23878;
  assign n24559 = ~n23864 & n24558;
  assign n24560 = ~n24331 & n24559;
  assign n24561 = n35403 & ~n35492;
  assign n24562 = ~n24560 & ~n24561;
  assign n24563 = ~n24555 & ~n35493;
  assign n24564 = ~n35491 & ~n35494;
  assign n24565 = ~n24547 & ~n24564;
  assign n24566 = ~n13704 & ~n24565;
  assign n24567 = n13704 & ~n24547;
  assign n24568 = ~n24564 & n24567;
  assign n24569 = ~n35404 & ~n23884;
  assign n24570 = ~n23884 & ~n24331;
  assign n24571 = ~n35404 & n24570;
  assign n24572 = ~n24331 & n24569;
  assign n24573 = n23709 & ~n35495;
  assign n24574 = n23883 & n24570;
  assign n24575 = n23709 & ~n35404;
  assign n24576 = ~n23884 & n24575;
  assign n24577 = ~n24331 & n24576;
  assign n24578 = ~n23709 & ~n35495;
  assign n24579 = ~n24577 & ~n24578;
  assign n24580 = ~n24573 & ~n24574;
  assign n24581 = ~n24568 & ~n35496;
  assign n24582 = ~n24566 & ~n24581;
  assign n24583 = ~n13099 & ~n24582;
  assign n24584 = n13099 & ~n24566;
  assign n24585 = ~n24581 & n24584;
  assign n24586 = n13099 & n24582;
  assign n24587 = ~n23886 & ~n23902;
  assign n24588 = ~n24331 & n24587;
  assign n24589 = ~n35407 & ~n24588;
  assign n24590 = n35407 & ~n23902;
  assign n24591 = ~n23886 & n24590;
  assign n24592 = n35407 & n24588;
  assign n24593 = ~n24331 & n24591;
  assign n24594 = ~n24589 & ~n35498;
  assign n24595 = ~n35497 & ~n24594;
  assign n24596 = ~n24583 & ~n24595;
  assign n24597 = ~n12442 & ~n24596;
  assign n24598 = n12442 & ~n24583;
  assign n24599 = ~n24595 & n24598;
  assign n24600 = ~n35408 & ~n23908;
  assign n24601 = ~n23908 & ~n24331;
  assign n24602 = ~n35408 & n24601;
  assign n24603 = ~n24331 & n24600;
  assign n24604 = n23701 & ~n35499;
  assign n24605 = n23907 & n24601;
  assign n24606 = n23701 & ~n35408;
  assign n24607 = ~n23908 & n24606;
  assign n24608 = ~n24331 & n24607;
  assign n24609 = ~n23701 & ~n35499;
  assign n24610 = ~n24608 & ~n24609;
  assign n24611 = ~n24604 & ~n24605;
  assign n24612 = ~n24599 & ~n35500;
  assign n24613 = ~n24597 & ~n24612;
  assign n24614 = ~n11858 & ~n24613;
  assign n24615 = n11858 & ~n24597;
  assign n24616 = ~n24612 & n24615;
  assign n24617 = n11858 & n24613;
  assign n24618 = ~n23910 & ~n23921;
  assign n24619 = ~n23921 & ~n24331;
  assign n24620 = ~n23910 & n24619;
  assign n24621 = ~n24331 & n24618;
  assign n24622 = n23918 & ~n35502;
  assign n24623 = n23919 & n24619;
  assign n24624 = ~n23918 & n35502;
  assign n24625 = n23918 & ~n23921;
  assign n24626 = ~n23910 & n24625;
  assign n24627 = ~n24331 & n24626;
  assign n24628 = ~n23918 & ~n35502;
  assign n24629 = ~n24627 & ~n24628;
  assign n24630 = ~n24622 & ~n35503;
  assign n24631 = ~n35501 & ~n35504;
  assign n24632 = ~n24614 & ~n24631;
  assign n24633 = ~n11229 & ~n24632;
  assign n24634 = n11229 & ~n24614;
  assign n24635 = ~n24631 & n24634;
  assign n24636 = ~n35410 & ~n23927;
  assign n24637 = ~n23927 & ~n24331;
  assign n24638 = ~n35410 & n24637;
  assign n24639 = ~n24331 & n24636;
  assign n24640 = n23693 & ~n35505;
  assign n24641 = n23926 & n24637;
  assign n24642 = n23693 & ~n35410;
  assign n24643 = ~n23927 & n24642;
  assign n24644 = ~n24331 & n24643;
  assign n24645 = ~n23693 & ~n35505;
  assign n24646 = ~n24644 & ~n24645;
  assign n24647 = ~n24640 & ~n24641;
  assign n24648 = ~n24635 & ~n35506;
  assign n24649 = ~n24633 & ~n24648;
  assign n24650 = ~n10681 & ~n24649;
  assign n24651 = n10681 & ~n24633;
  assign n24652 = ~n24648 & n24651;
  assign n24653 = n10681 & n24649;
  assign n24654 = ~n23929 & ~n23945;
  assign n24655 = ~n24331 & n24654;
  assign n24656 = ~n35413 & n24655;
  assign n24657 = n35413 & ~n24655;
  assign n24658 = n35413 & ~n23945;
  assign n24659 = ~n23929 & n24658;
  assign n24660 = n35413 & n24655;
  assign n24661 = ~n24331 & n24659;
  assign n24662 = ~n35413 & ~n24655;
  assign n24663 = ~n35508 & ~n24662;
  assign n24664 = ~n24656 & ~n24657;
  assign n24665 = ~n35507 & ~n35509;
  assign n24666 = ~n24650 & ~n24665;
  assign n24667 = ~n10086 & ~n24666;
  assign n24668 = n10086 & ~n24650;
  assign n24669 = ~n24665 & n24668;
  assign n24670 = ~n35414 & ~n23951;
  assign n24671 = ~n23951 & ~n24331;
  assign n24672 = ~n35414 & n24671;
  assign n24673 = ~n24331 & n24670;
  assign n24674 = n23685 & ~n35510;
  assign n24675 = n23950 & n24671;
  assign n24676 = n23685 & ~n35414;
  assign n24677 = ~n23951 & n24676;
  assign n24678 = ~n24331 & n24677;
  assign n24679 = ~n23685 & ~n35510;
  assign n24680 = ~n24678 & ~n24679;
  assign n24681 = ~n24674 & ~n24675;
  assign n24682 = ~n24669 & ~n35511;
  assign n24683 = ~n24667 & ~n24682;
  assign n24684 = ~n9565 & ~n24683;
  assign n24685 = n9565 & ~n24667;
  assign n24686 = ~n24682 & n24685;
  assign n24687 = n9565 & n24683;
  assign n24688 = ~n23953 & ~n23967;
  assign n24689 = ~n23967 & ~n24331;
  assign n24690 = ~n23953 & n24689;
  assign n24691 = ~n24331 & n24688;
  assign n24692 = n35416 & ~n35513;
  assign n24693 = n23965 & n24689;
  assign n24694 = ~n35416 & n35513;
  assign n24695 = n35416 & ~n23967;
  assign n24696 = ~n23953 & n24695;
  assign n24697 = ~n24331 & n24696;
  assign n24698 = ~n35416 & ~n35513;
  assign n24699 = ~n24697 & ~n24698;
  assign n24700 = ~n24692 & ~n35514;
  assign n24701 = ~n35512 & ~n35515;
  assign n24702 = ~n24684 & ~n24701;
  assign n24703 = ~n8998 & ~n24702;
  assign n24704 = n8998 & ~n24684;
  assign n24705 = ~n24701 & n24704;
  assign n24706 = ~n35417 & ~n23973;
  assign n24707 = ~n23973 & ~n24331;
  assign n24708 = ~n35417 & n24707;
  assign n24709 = ~n24331 & n24706;
  assign n24710 = n23677 & ~n35516;
  assign n24711 = n23972 & n24707;
  assign n24712 = n23677 & ~n35417;
  assign n24713 = ~n23973 & n24712;
  assign n24714 = ~n24331 & n24713;
  assign n24715 = ~n23677 & ~n35516;
  assign n24716 = ~n24714 & ~n24715;
  assign n24717 = ~n24710 & ~n24711;
  assign n24718 = ~n24705 & ~n35517;
  assign n24719 = ~n24703 & ~n24718;
  assign n24720 = ~n8506 & ~n24719;
  assign n24721 = ~n23975 & ~n23991;
  assign n24722 = ~n24331 & n24721;
  assign n24723 = ~n35420 & ~n24722;
  assign n24724 = n35420 & ~n23991;
  assign n24725 = ~n23975 & n24724;
  assign n24726 = n35420 & n24722;
  assign n24727 = ~n24331 & n24725;
  assign n24728 = ~n24723 & ~n35518;
  assign n24729 = n8506 & ~n24703;
  assign n24730 = ~n24718 & n24729;
  assign n24731 = n8506 & n24719;
  assign n24732 = ~n24728 & ~n35519;
  assign n24733 = ~n24720 & ~n24732;
  assign n24734 = ~n7975 & ~n24733;
  assign n24735 = n7975 & ~n24720;
  assign n24736 = ~n24732 & n24735;
  assign n24737 = ~n35421 & ~n23997;
  assign n24738 = ~n23997 & ~n24331;
  assign n24739 = ~n35421 & n24738;
  assign n24740 = ~n24331 & n24737;
  assign n24741 = n23669 & ~n35520;
  assign n24742 = n23996 & n24738;
  assign n24743 = n23669 & ~n35421;
  assign n24744 = ~n23997 & n24743;
  assign n24745 = ~n24331 & n24744;
  assign n24746 = ~n23669 & ~n35520;
  assign n24747 = ~n24745 & ~n24746;
  assign n24748 = ~n24741 & ~n24742;
  assign n24749 = ~n24736 & ~n35521;
  assign n24750 = ~n24734 & ~n24749;
  assign n24751 = ~n7512 & ~n24750;
  assign n24752 = n7512 & ~n24734;
  assign n24753 = ~n24749 & n24752;
  assign n24754 = n7512 & n24750;
  assign n24755 = ~n23999 & ~n24002;
  assign n24756 = ~n24002 & ~n24331;
  assign n24757 = ~n23999 & n24756;
  assign n24758 = ~n24331 & n24755;
  assign n24759 = n23661 & ~n35523;
  assign n24760 = n24000 & n24756;
  assign n24761 = n23661 & ~n24002;
  assign n24762 = ~n23999 & n24761;
  assign n24763 = ~n24331 & n24762;
  assign n24764 = ~n23661 & ~n35523;
  assign n24765 = ~n24763 & ~n24764;
  assign n24766 = ~n24759 & ~n24760;
  assign n24767 = ~n35522 & ~n35524;
  assign n24768 = ~n24751 & ~n24767;
  assign n24769 = ~n7015 & ~n24768;
  assign n24770 = n7015 & ~n24751;
  assign n24771 = ~n24767 & n24770;
  assign n24772 = ~n35422 & ~n24008;
  assign n24773 = ~n24008 & ~n24331;
  assign n24774 = ~n35422 & n24773;
  assign n24775 = ~n24331 & n24772;
  assign n24776 = n23653 & ~n35525;
  assign n24777 = n24007 & n24773;
  assign n24778 = n23653 & ~n35422;
  assign n24779 = ~n24008 & n24778;
  assign n24780 = ~n24331 & n24779;
  assign n24781 = ~n23653 & ~n35525;
  assign n24782 = ~n24780 & ~n24781;
  assign n24783 = ~n24776 & ~n24777;
  assign n24784 = ~n24771 & ~n35526;
  assign n24785 = ~n24769 & ~n24784;
  assign n24786 = ~n6579 & ~n24785;
  assign n24787 = ~n24010 & ~n24025;
  assign n24788 = ~n24331 & n24787;
  assign n24789 = ~n35424 & ~n24788;
  assign n24790 = n35424 & ~n24025;
  assign n24791 = ~n24010 & n24790;
  assign n24792 = n35424 & n24788;
  assign n24793 = ~n24331 & n24791;
  assign n24794 = ~n24789 & ~n35527;
  assign n24795 = n6579 & ~n24769;
  assign n24796 = ~n24784 & n24795;
  assign n24797 = n6579 & n24785;
  assign n24798 = ~n24794 & ~n35528;
  assign n24799 = ~n24786 & ~n24798;
  assign n24800 = ~n6117 & ~n24799;
  assign n24801 = n6117 & ~n24786;
  assign n24802 = ~n24798 & n24801;
  assign n24803 = ~n35425 & ~n24031;
  assign n24804 = ~n24031 & ~n24331;
  assign n24805 = ~n35425 & n24804;
  assign n24806 = ~n24331 & n24803;
  assign n24807 = n23645 & ~n35529;
  assign n24808 = n24030 & n24804;
  assign n24809 = n23645 & ~n35425;
  assign n24810 = ~n24031 & n24809;
  assign n24811 = ~n24331 & n24810;
  assign n24812 = ~n23645 & ~n35529;
  assign n24813 = ~n24811 & ~n24812;
  assign n24814 = ~n24807 & ~n24808;
  assign n24815 = ~n24802 & ~n35530;
  assign n24816 = ~n24800 & ~n24815;
  assign n24817 = ~n5708 & ~n24816;
  assign n24818 = n5708 & ~n24800;
  assign n24819 = ~n24815 & n24818;
  assign n24820 = n5708 & n24816;
  assign n24821 = ~n24033 & ~n24036;
  assign n24822 = ~n24036 & ~n24331;
  assign n24823 = ~n24033 & n24822;
  assign n24824 = ~n24331 & n24821;
  assign n24825 = n23637 & ~n35532;
  assign n24826 = n24034 & n24822;
  assign n24827 = n23637 & ~n24036;
  assign n24828 = ~n24033 & n24827;
  assign n24829 = ~n24331 & n24828;
  assign n24830 = ~n23637 & ~n35532;
  assign n24831 = ~n24829 & ~n24830;
  assign n24832 = ~n24825 & ~n24826;
  assign n24833 = ~n35531 & ~n35533;
  assign n24834 = ~n24817 & ~n24833;
  assign n24835 = ~n5278 & ~n24834;
  assign n24836 = n5278 & ~n24817;
  assign n24837 = ~n24833 & n24836;
  assign n24838 = ~n35426 & ~n24042;
  assign n24839 = ~n24042 & ~n24331;
  assign n24840 = ~n35426 & n24839;
  assign n24841 = ~n24331 & n24838;
  assign n24842 = n23629 & ~n35534;
  assign n24843 = n24041 & n24839;
  assign n24844 = n23629 & ~n35426;
  assign n24845 = ~n24042 & n24844;
  assign n24846 = ~n24331 & n24845;
  assign n24847 = ~n23629 & ~n35534;
  assign n24848 = ~n24846 & ~n24847;
  assign n24849 = ~n24842 & ~n24843;
  assign n24850 = ~n24837 & ~n35535;
  assign n24851 = ~n24835 & ~n24850;
  assign n24852 = ~n4903 & ~n24851;
  assign n24853 = ~n24044 & ~n24059;
  assign n24854 = ~n24331 & n24853;
  assign n24855 = ~n35428 & ~n24854;
  assign n24856 = n35428 & ~n24059;
  assign n24857 = ~n24044 & n24856;
  assign n24858 = n35428 & n24854;
  assign n24859 = ~n24331 & n24857;
  assign n24860 = ~n24855 & ~n35536;
  assign n24861 = n4903 & ~n24835;
  assign n24862 = ~n24850 & n24861;
  assign n24863 = n4903 & n24851;
  assign n24864 = ~n24860 & ~n35537;
  assign n24865 = ~n24852 & ~n24864;
  assign n24866 = ~n4508 & ~n24865;
  assign n24867 = n4508 & ~n24852;
  assign n24868 = ~n24864 & n24867;
  assign n24869 = ~n35429 & ~n24065;
  assign n24870 = ~n24065 & ~n24331;
  assign n24871 = ~n35429 & n24870;
  assign n24872 = ~n24331 & n24869;
  assign n24873 = n23621 & ~n35538;
  assign n24874 = n24064 & n24870;
  assign n24875 = n23621 & ~n35429;
  assign n24876 = ~n24065 & n24875;
  assign n24877 = ~n24331 & n24876;
  assign n24878 = ~n23621 & ~n35538;
  assign n24879 = ~n24877 & ~n24878;
  assign n24880 = ~n24873 & ~n24874;
  assign n24881 = ~n24868 & ~n35539;
  assign n24882 = ~n24866 & ~n24881;
  assign n24883 = ~n4155 & ~n24882;
  assign n24884 = n4155 & ~n24866;
  assign n24885 = ~n24881 & n24884;
  assign n24886 = n4155 & n24882;
  assign n24887 = ~n24067 & ~n24070;
  assign n24888 = ~n24070 & ~n24331;
  assign n24889 = ~n24067 & n24888;
  assign n24890 = ~n24331 & n24887;
  assign n24891 = n23613 & ~n35541;
  assign n24892 = n24068 & n24888;
  assign n24893 = n23613 & ~n24070;
  assign n24894 = ~n24067 & n24893;
  assign n24895 = ~n24331 & n24894;
  assign n24896 = ~n23613 & ~n35541;
  assign n24897 = ~n24895 & ~n24896;
  assign n24898 = ~n24891 & ~n24892;
  assign n24899 = ~n35540 & ~n35542;
  assign n24900 = ~n24883 & ~n24899;
  assign n24901 = ~n3788 & ~n24900;
  assign n24902 = n3788 & ~n24883;
  assign n24903 = ~n24899 & n24902;
  assign n24904 = ~n35430 & ~n24076;
  assign n24905 = ~n24076 & ~n24331;
  assign n24906 = ~n35430 & n24905;
  assign n24907 = ~n24331 & n24904;
  assign n24908 = n23605 & ~n35543;
  assign n24909 = n24075 & n24905;
  assign n24910 = n23605 & ~n35430;
  assign n24911 = ~n24076 & n24910;
  assign n24912 = ~n24331 & n24911;
  assign n24913 = ~n23605 & ~n35543;
  assign n24914 = ~n24912 & ~n24913;
  assign n24915 = ~n24908 & ~n24909;
  assign n24916 = ~n24903 & ~n35544;
  assign n24917 = ~n24901 & ~n24916;
  assign n24918 = ~n3473 & ~n24917;
  assign n24919 = ~n24078 & ~n24093;
  assign n24920 = ~n24331 & n24919;
  assign n24921 = ~n35432 & ~n24920;
  assign n24922 = n35432 & ~n24093;
  assign n24923 = ~n24078 & n24922;
  assign n24924 = n35432 & n24920;
  assign n24925 = ~n24331 & n24923;
  assign n24926 = ~n24921 & ~n35545;
  assign n24927 = n3473 & ~n24901;
  assign n24928 = ~n24916 & n24927;
  assign n24929 = n3473 & n24917;
  assign n24930 = ~n24926 & ~n35546;
  assign n24931 = ~n24918 & ~n24930;
  assign n24932 = ~n3140 & ~n24931;
  assign n24933 = n3140 & ~n24918;
  assign n24934 = ~n24930 & n24933;
  assign n24935 = ~n35433 & ~n24099;
  assign n24936 = ~n24099 & ~n24331;
  assign n24937 = ~n35433 & n24936;
  assign n24938 = ~n24331 & n24935;
  assign n24939 = n23597 & ~n35547;
  assign n24940 = n24098 & n24936;
  assign n24941 = n23597 & ~n35433;
  assign n24942 = ~n24099 & n24941;
  assign n24943 = ~n24331 & n24942;
  assign n24944 = ~n23597 & ~n35547;
  assign n24945 = ~n24943 & ~n24944;
  assign n24946 = ~n24939 & ~n24940;
  assign n24947 = ~n24934 & ~n35548;
  assign n24948 = ~n24932 & ~n24947;
  assign n24949 = ~n2855 & ~n24948;
  assign n24950 = n2855 & ~n24932;
  assign n24951 = ~n24947 & n24950;
  assign n24952 = n2855 & n24948;
  assign n24953 = ~n24101 & ~n24104;
  assign n24954 = ~n24104 & ~n24331;
  assign n24955 = ~n24101 & n24954;
  assign n24956 = ~n24331 & n24953;
  assign n24957 = n23589 & ~n35550;
  assign n24958 = n24102 & n24954;
  assign n24959 = n23589 & ~n24104;
  assign n24960 = ~n24101 & n24959;
  assign n24961 = ~n24331 & n24960;
  assign n24962 = ~n23589 & ~n35550;
  assign n24963 = ~n24961 & ~n24962;
  assign n24964 = ~n24957 & ~n24958;
  assign n24965 = ~n35549 & ~n35551;
  assign n24966 = ~n24949 & ~n24965;
  assign n24967 = ~n2556 & ~n24966;
  assign n24968 = n2556 & ~n24949;
  assign n24969 = ~n24965 & n24968;
  assign n24970 = ~n35434 & ~n24110;
  assign n24971 = ~n24110 & ~n24331;
  assign n24972 = ~n35434 & n24971;
  assign n24973 = ~n24331 & n24970;
  assign n24974 = n23581 & ~n35552;
  assign n24975 = n24109 & n24971;
  assign n24976 = n23581 & ~n35434;
  assign n24977 = ~n24110 & n24976;
  assign n24978 = ~n24331 & n24977;
  assign n24979 = ~n23581 & ~n35552;
  assign n24980 = ~n24978 & ~n24979;
  assign n24981 = ~n24974 & ~n24975;
  assign n24982 = ~n24969 & ~n35553;
  assign n24983 = ~n24967 & ~n24982;
  assign n24984 = ~n2301 & ~n24983;
  assign n24985 = ~n24112 & ~n24127;
  assign n24986 = ~n24331 & n24985;
  assign n24987 = ~n35436 & ~n24986;
  assign n24988 = n35436 & ~n24127;
  assign n24989 = ~n24112 & n24988;
  assign n24990 = n35436 & n24986;
  assign n24991 = ~n24331 & n24989;
  assign n24992 = ~n24987 & ~n35554;
  assign n24993 = n2301 & ~n24967;
  assign n24994 = ~n24982 & n24993;
  assign n24995 = n2301 & n24983;
  assign n24996 = ~n24992 & ~n35555;
  assign n24997 = ~n24984 & ~n24996;
  assign n24998 = ~n2038 & ~n24997;
  assign n24999 = n2038 & ~n24984;
  assign n25000 = ~n24996 & n24999;
  assign n25001 = ~n35437 & ~n24133;
  assign n25002 = ~n24133 & ~n24331;
  assign n25003 = ~n35437 & n25002;
  assign n25004 = ~n24331 & n25001;
  assign n25005 = n23573 & ~n35556;
  assign n25006 = n24132 & n25002;
  assign n25007 = n23573 & ~n35437;
  assign n25008 = ~n24133 & n25007;
  assign n25009 = ~n24331 & n25008;
  assign n25010 = ~n23573 & ~n35556;
  assign n25011 = ~n25009 & ~n25010;
  assign n25012 = ~n25005 & ~n25006;
  assign n25013 = ~n25000 & ~n35557;
  assign n25014 = ~n24998 & ~n25013;
  assign n25015 = ~n1812 & ~n25014;
  assign n25016 = n1812 & ~n24998;
  assign n25017 = ~n25013 & n25016;
  assign n25018 = n1812 & n25014;
  assign n25019 = ~n24135 & ~n24138;
  assign n25020 = ~n24138 & ~n24331;
  assign n25021 = ~n24135 & n25020;
  assign n25022 = ~n24331 & n25019;
  assign n25023 = n23565 & ~n35559;
  assign n25024 = n24136 & n25020;
  assign n25025 = n23565 & ~n24138;
  assign n25026 = ~n24135 & n25025;
  assign n25027 = ~n24331 & n25026;
  assign n25028 = ~n23565 & ~n35559;
  assign n25029 = ~n25027 & ~n25028;
  assign n25030 = ~n25023 & ~n25024;
  assign n25031 = ~n35558 & ~n35560;
  assign n25032 = ~n25015 & ~n25031;
  assign n25033 = ~n1582 & ~n25032;
  assign n25034 = n1582 & ~n25015;
  assign n25035 = ~n25031 & n25034;
  assign n25036 = ~n35438 & ~n24144;
  assign n25037 = ~n24144 & ~n24331;
  assign n25038 = ~n35438 & n25037;
  assign n25039 = ~n24331 & n25036;
  assign n25040 = n23557 & ~n35561;
  assign n25041 = n24143 & n25037;
  assign n25042 = n23557 & ~n35438;
  assign n25043 = ~n24144 & n25042;
  assign n25044 = ~n24331 & n25043;
  assign n25045 = ~n23557 & ~n35561;
  assign n25046 = ~n25044 & ~n25045;
  assign n25047 = ~n25040 & ~n25041;
  assign n25048 = ~n25035 & ~n35562;
  assign n25049 = ~n25033 & ~n25048;
  assign n25050 = ~n1388 & ~n25049;
  assign n25051 = ~n24146 & ~n24161;
  assign n25052 = ~n24331 & n25051;
  assign n25053 = ~n35440 & ~n25052;
  assign n25054 = n35440 & ~n24161;
  assign n25055 = ~n24146 & n25054;
  assign n25056 = n35440 & n25052;
  assign n25057 = ~n24331 & n25055;
  assign n25058 = ~n25053 & ~n35563;
  assign n25059 = n1388 & ~n25033;
  assign n25060 = ~n25048 & n25059;
  assign n25061 = n1388 & n25049;
  assign n25062 = ~n25058 & ~n35564;
  assign n25063 = ~n25050 & ~n25062;
  assign n25064 = ~n1192 & ~n25063;
  assign n25065 = n1192 & ~n25050;
  assign n25066 = ~n25062 & n25065;
  assign n25067 = ~n35441 & ~n24167;
  assign n25068 = ~n24167 & ~n24331;
  assign n25069 = ~n35441 & n25068;
  assign n25070 = ~n24331 & n25067;
  assign n25071 = n23549 & ~n35565;
  assign n25072 = n24166 & n25068;
  assign n25073 = n23549 & ~n35441;
  assign n25074 = ~n24167 & n25073;
  assign n25075 = ~n24331 & n25074;
  assign n25076 = ~n23549 & ~n35565;
  assign n25077 = ~n25075 & ~n25076;
  assign n25078 = ~n25071 & ~n25072;
  assign n25079 = ~n25066 & ~n35566;
  assign n25080 = ~n25064 & ~n25079;
  assign n25081 = ~n1028 & ~n25080;
  assign n25082 = n1028 & ~n25064;
  assign n25083 = ~n25079 & n25082;
  assign n25084 = n1028 & n25080;
  assign n25085 = ~n24169 & ~n24172;
  assign n25086 = ~n24172 & ~n24331;
  assign n25087 = ~n24169 & n25086;
  assign n25088 = ~n24331 & n25085;
  assign n25089 = n23541 & ~n35568;
  assign n25090 = n24170 & n25086;
  assign n25091 = n23541 & ~n24172;
  assign n25092 = ~n24169 & n25091;
  assign n25093 = ~n24331 & n25092;
  assign n25094 = ~n23541 & ~n35568;
  assign n25095 = ~n25093 & ~n25094;
  assign n25096 = ~n25089 & ~n25090;
  assign n25097 = ~n35567 & ~n35569;
  assign n25098 = ~n25081 & ~n25097;
  assign n25099 = ~n866 & ~n25098;
  assign n25100 = n866 & ~n25081;
  assign n25101 = ~n25097 & n25100;
  assign n25102 = ~n35442 & ~n24178;
  assign n25103 = ~n24331 & n25102;
  assign n25104 = n23533 & ~n25103;
  assign n25105 = ~n23533 & n25103;
  assign n25106 = n23533 & ~n35442;
  assign n25107 = ~n24178 & n25106;
  assign n25108 = ~n24331 & n25107;
  assign n25109 = ~n23533 & ~n25103;
  assign n25110 = ~n25108 & ~n25109;
  assign n25111 = ~n25104 & ~n25105;
  assign n25112 = ~n25101 & ~n35570;
  assign n25113 = ~n25099 & ~n25112;
  assign n25114 = ~n730 & ~n25113;
  assign n25115 = ~n24180 & ~n24182;
  assign n25116 = ~n24331 & n25115;
  assign n25117 = n35444 & ~n25116;
  assign n25118 = ~n24180 & ~n35444;
  assign n25119 = ~n24182 & n25118;
  assign n25120 = ~n35444 & n25116;
  assign n25121 = ~n24331 & n25119;
  assign n25122 = n35444 & n25116;
  assign n25123 = ~n35444 & ~n25116;
  assign n25124 = ~n25122 & ~n25123;
  assign n25125 = ~n25117 & ~n35571;
  assign n25126 = n730 & ~n25099;
  assign n25127 = ~n25112 & n25126;
  assign n25128 = n730 & n25113;
  assign n25129 = n35572 & ~n35573;
  assign n25130 = ~n25114 & ~n25129;
  assign n25131 = ~n602 & ~n25130;
  assign n25132 = n602 & ~n25114;
  assign n25133 = ~n25129 & n25132;
  assign n25134 = ~n35463 & ~n25133;
  assign n25135 = ~n25131 & ~n25134;
  assign n25136 = ~n497 & ~n25135;
  assign n25137 = ~n24202 & ~n24204;
  assign n25138 = ~n24331 & n25137;
  assign n25139 = ~n35447 & ~n25138;
  assign n25140 = ~n24202 & n35447;
  assign n25141 = ~n24204 & n25140;
  assign n25142 = n35447 & n25138;
  assign n25143 = ~n24331 & n25141;
  assign n25144 = ~n25139 & ~n35574;
  assign n25145 = n497 & ~n25131;
  assign n25146 = ~n25134 & n25145;
  assign n25147 = n497 & n25135;
  assign n25148 = ~n25144 & ~n35575;
  assign n25149 = ~n25136 & ~n25148;
  assign n25150 = ~n403 & ~n25149;
  assign n25151 = n403 & ~n25136;
  assign n25152 = ~n25148 & n25151;
  assign n25153 = ~n24219 & ~n35449;
  assign n25154 = ~n24219 & ~n24331;
  assign n25155 = ~n35449 & n25154;
  assign n25156 = ~n24331 & n25153;
  assign n25157 = n24227 & ~n35576;
  assign n25158 = n24231 & n25154;
  assign n25159 = n24227 & ~n35449;
  assign n25160 = ~n24219 & n25159;
  assign n25161 = ~n24331 & n25160;
  assign n25162 = ~n24227 & ~n35576;
  assign n25163 = ~n25161 & ~n25162;
  assign n25164 = ~n25157 & ~n25158;
  assign n25165 = ~n25152 & ~n35577;
  assign n25166 = ~n25150 & ~n25165;
  assign n25167 = ~n330 & ~n25166;
  assign n25168 = ~n24233 & ~n24235;
  assign n25169 = ~n24331 & n25168;
  assign n25170 = ~n35451 & ~n25169;
  assign n25171 = ~n24233 & n35451;
  assign n25172 = ~n24235 & n25171;
  assign n25173 = n35451 & n25169;
  assign n25174 = ~n24331 & n25172;
  assign n25175 = ~n25170 & ~n35578;
  assign n25176 = n330 & ~n25150;
  assign n25177 = ~n25165 & n25176;
  assign n25178 = n330 & n25166;
  assign n25179 = ~n25175 & ~n35579;
  assign n25180 = ~n25167 & ~n25179;
  assign n25181 = ~n271 & ~n25180;
  assign n25182 = n271 & ~n25167;
  assign n25183 = ~n25179 & n25182;
  assign n25184 = ~n24250 & ~n35453;
  assign n25185 = ~n24250 & ~n24331;
  assign n25186 = ~n35453 & n25185;
  assign n25187 = ~n24331 & n25184;
  assign n25188 = n24258 & ~n35580;
  assign n25189 = n24262 & n25185;
  assign n25190 = n24258 & ~n35453;
  assign n25191 = ~n24250 & n25190;
  assign n25192 = ~n24331 & n25191;
  assign n25193 = ~n24258 & ~n35580;
  assign n25194 = ~n25192 & ~n25193;
  assign n25195 = ~n25188 & ~n25189;
  assign n25196 = ~n25183 & ~n35581;
  assign n25197 = ~n25181 & ~n25196;
  assign n25198 = ~n217 & ~n25197;
  assign n25199 = n217 & ~n25181;
  assign n25200 = ~n25196 & n25199;
  assign n25201 = n217 & n25197;
  assign n25202 = ~n24264 & ~n24274;
  assign n25203 = ~n24264 & ~n24331;
  assign n25204 = ~n24274 & n25203;
  assign n25205 = ~n24331 & n25202;
  assign n25206 = n24272 & ~n35583;
  assign n25207 = n24275 & n25203;
  assign n25208 = ~n24264 & n24272;
  assign n25209 = ~n24274 & n25208;
  assign n25210 = ~n24331 & n25209;
  assign n25211 = ~n24272 & ~n35583;
  assign n25212 = ~n25210 & ~n25211;
  assign n25213 = ~n25206 & ~n25207;
  assign n25214 = ~n35582 & ~n35584;
  assign n25215 = ~n25198 & ~n25214;
  assign n25216 = ~n198 & ~n25215;
  assign n25217 = n198 & ~n25198;
  assign n25218 = ~n25214 & n25217;
  assign n25219 = ~n24277 & ~n35456;
  assign n25220 = ~n24277 & ~n24331;
  assign n25221 = ~n35456 & n25220;
  assign n25222 = ~n24331 & n25219;
  assign n25223 = n24285 & ~n35585;
  assign n25224 = n24289 & n25220;
  assign n25225 = n24285 & ~n35456;
  assign n25226 = ~n24277 & n25225;
  assign n25227 = ~n24331 & n25226;
  assign n25228 = ~n24285 & ~n35585;
  assign n25229 = ~n25227 & ~n25228;
  assign n25230 = ~n25223 & ~n25224;
  assign n25231 = ~n25218 & ~n35586;
  assign n25232 = ~n25216 & ~n25231;
  assign n25233 = ~n24291 & ~n24293;
  assign n25234 = ~n24331 & n25233;
  assign n25235 = ~n35458 & ~n25234;
  assign n25236 = ~n24291 & n35458;
  assign n25237 = ~n24293 & n25236;
  assign n25238 = n35458 & n25234;
  assign n25239 = ~n24331 & n25237;
  assign n25240 = ~n25235 & ~n35587;
  assign n25241 = ~n24307 & ~n24315;
  assign n25242 = ~n24315 & ~n24331;
  assign n25243 = ~n24307 & n25242;
  assign n25244 = ~n24331 & n25241;
  assign n25245 = ~n35461 & ~n35588;
  assign n25246 = ~n25240 & n25245;
  assign n25247 = ~n25232 & n25246;
  assign n25248 = n193 & ~n25247;
  assign n25249 = ~n25216 & n25240;
  assign n25250 = ~n25231 & n25249;
  assign n25251 = n25232 & n25240;
  assign n25252 = n24307 & ~n25242;
  assign n25253 = ~n193 & ~n25241;
  assign n25254 = ~n25252 & n25253;
  assign n25255 = ~n35589 & ~n25254;
  assign n25256 = ~n25248 & n25255;
  assign n25257 = ~n25131 & ~n25133;
  assign n25258 = ~n25256 & n25257;
  assign n25259 = ~n35463 & ~n25258;
  assign n25260 = n35463 & ~n25133;
  assign n25261 = ~n25131 & n25260;
  assign n25262 = n35463 & n25258;
  assign n25263 = ~n25256 & n25261;
  assign n25264 = ~n25259 & ~n35590;
  assign n25265 = ~n25081 & ~n35567;
  assign n25266 = ~n25256 & n25265;
  assign n25267 = ~n35569 & ~n25266;
  assign n25268 = ~n25081 & n35569;
  assign n25269 = ~n35567 & n25268;
  assign n25270 = n35569 & n25266;
  assign n25271 = ~n25256 & n25269;
  assign n25272 = ~n25267 & ~n35591;
  assign n25273 = ~n25064 & ~n25066;
  assign n25274 = ~n25256 & n25273;
  assign n25275 = ~n35566 & ~n25274;
  assign n25276 = ~n25066 & n35566;
  assign n25277 = ~n25064 & n25276;
  assign n25278 = n35566 & n25274;
  assign n25279 = ~n25256 & n25277;
  assign n25280 = ~n25275 & ~n35592;
  assign n25281 = ~n25033 & ~n25035;
  assign n25282 = ~n25256 & n25281;
  assign n25283 = ~n35562 & ~n25282;
  assign n25284 = ~n25035 & n35562;
  assign n25285 = ~n25033 & n25284;
  assign n25286 = n35562 & n25282;
  assign n25287 = ~n25256 & n25285;
  assign n25288 = ~n25283 & ~n35593;
  assign n25289 = ~n25015 & ~n35558;
  assign n25290 = ~n25256 & n25289;
  assign n25291 = ~n35560 & ~n25290;
  assign n25292 = ~n25015 & n35560;
  assign n25293 = ~n35558 & n25292;
  assign n25294 = n35560 & n25290;
  assign n25295 = ~n25256 & n25293;
  assign n25296 = ~n25291 & ~n35594;
  assign n25297 = ~n24998 & ~n25000;
  assign n25298 = ~n25256 & n25297;
  assign n25299 = ~n35557 & ~n25298;
  assign n25300 = ~n25000 & n35557;
  assign n25301 = ~n24998 & n25300;
  assign n25302 = n35557 & n25298;
  assign n25303 = ~n25256 & n25301;
  assign n25304 = ~n25299 & ~n35595;
  assign n25305 = ~n24967 & ~n24969;
  assign n25306 = ~n25256 & n25305;
  assign n25307 = ~n35553 & ~n25306;
  assign n25308 = ~n24969 & n35553;
  assign n25309 = ~n24967 & n25308;
  assign n25310 = n35553 & n25306;
  assign n25311 = ~n25256 & n25309;
  assign n25312 = ~n25307 & ~n35596;
  assign n25313 = ~n24949 & ~n35549;
  assign n25314 = ~n25256 & n25313;
  assign n25315 = ~n35551 & ~n25314;
  assign n25316 = ~n24949 & n35551;
  assign n25317 = ~n35549 & n25316;
  assign n25318 = n35551 & n25314;
  assign n25319 = ~n25256 & n25317;
  assign n25320 = ~n25315 & ~n35597;
  assign n25321 = ~n24932 & ~n24934;
  assign n25322 = ~n25256 & n25321;
  assign n25323 = ~n35548 & ~n25322;
  assign n25324 = ~n24934 & n35548;
  assign n25325 = ~n24932 & n25324;
  assign n25326 = n35548 & n25322;
  assign n25327 = ~n25256 & n25325;
  assign n25328 = ~n25323 & ~n35598;
  assign n25329 = ~n24901 & ~n24903;
  assign n25330 = ~n25256 & n25329;
  assign n25331 = ~n35544 & ~n25330;
  assign n25332 = ~n24903 & n35544;
  assign n25333 = ~n24901 & n25332;
  assign n25334 = n35544 & n25330;
  assign n25335 = ~n25256 & n25333;
  assign n25336 = ~n25331 & ~n35599;
  assign n25337 = ~n24883 & ~n35540;
  assign n25338 = ~n25256 & n25337;
  assign n25339 = ~n35542 & ~n25338;
  assign n25340 = ~n24883 & n35542;
  assign n25341 = ~n35540 & n25340;
  assign n25342 = n35542 & n25338;
  assign n25343 = ~n25256 & n25341;
  assign n25344 = ~n25339 & ~n35600;
  assign n25345 = ~n24866 & ~n24868;
  assign n25346 = ~n25256 & n25345;
  assign n25347 = ~n35539 & ~n25346;
  assign n25348 = ~n24868 & n35539;
  assign n25349 = ~n24866 & n25348;
  assign n25350 = n35539 & n25346;
  assign n25351 = ~n25256 & n25349;
  assign n25352 = ~n25347 & ~n35601;
  assign n25353 = ~n24835 & ~n24837;
  assign n25354 = ~n25256 & n25353;
  assign n25355 = ~n35535 & ~n25354;
  assign n25356 = ~n24837 & n35535;
  assign n25357 = ~n24835 & n25356;
  assign n25358 = n35535 & n25354;
  assign n25359 = ~n25256 & n25357;
  assign n25360 = ~n25355 & ~n35602;
  assign n25361 = ~n24817 & ~n35531;
  assign n25362 = ~n25256 & n25361;
  assign n25363 = ~n35533 & ~n25362;
  assign n25364 = ~n24817 & n35533;
  assign n25365 = ~n35531 & n25364;
  assign n25366 = n35533 & n25362;
  assign n25367 = ~n25256 & n25365;
  assign n25368 = ~n25363 & ~n35603;
  assign n25369 = ~n24800 & ~n24802;
  assign n25370 = ~n25256 & n25369;
  assign n25371 = ~n35530 & ~n25370;
  assign n25372 = ~n24802 & n35530;
  assign n25373 = ~n24800 & n25372;
  assign n25374 = n35530 & n25370;
  assign n25375 = ~n25256 & n25373;
  assign n25376 = ~n25371 & ~n35604;
  assign n25377 = ~n24769 & ~n24771;
  assign n25378 = ~n25256 & n25377;
  assign n25379 = ~n35526 & ~n25378;
  assign n25380 = ~n24771 & n35526;
  assign n25381 = ~n24769 & n25380;
  assign n25382 = n35526 & n25378;
  assign n25383 = ~n25256 & n25381;
  assign n25384 = ~n25379 & ~n35605;
  assign n25385 = ~n24751 & ~n35522;
  assign n25386 = ~n25256 & n25385;
  assign n25387 = ~n35524 & ~n25386;
  assign n25388 = ~n24751 & n35524;
  assign n25389 = ~n35522 & n25388;
  assign n25390 = n35524 & n25386;
  assign n25391 = ~n25256 & n25389;
  assign n25392 = ~n25387 & ~n35606;
  assign n25393 = ~n24734 & ~n24736;
  assign n25394 = ~n25256 & n25393;
  assign n25395 = ~n35521 & ~n25394;
  assign n25396 = ~n24736 & n35521;
  assign n25397 = ~n24734 & n25396;
  assign n25398 = n35521 & n25394;
  assign n25399 = ~n25256 & n25397;
  assign n25400 = ~n25395 & ~n35607;
  assign n25401 = ~n24703 & ~n24705;
  assign n25402 = ~n25256 & n25401;
  assign n25403 = ~n35517 & ~n25402;
  assign n25404 = ~n24705 & n35517;
  assign n25405 = ~n24703 & n25404;
  assign n25406 = n35517 & n25402;
  assign n25407 = ~n25256 & n25405;
  assign n25408 = ~n25403 & ~n35608;
  assign n25409 = ~n24684 & ~n35512;
  assign n25410 = ~n25256 & n25409;
  assign n25411 = ~n35515 & ~n25410;
  assign n25412 = ~n24684 & n35515;
  assign n25413 = ~n35512 & n25412;
  assign n25414 = n35515 & n25410;
  assign n25415 = ~n25256 & n25413;
  assign n25416 = ~n25411 & ~n35609;
  assign n25417 = ~n24667 & ~n24669;
  assign n25418 = ~n25256 & n25417;
  assign n25419 = ~n35511 & ~n25418;
  assign n25420 = ~n24669 & n35511;
  assign n25421 = ~n24667 & n25420;
  assign n25422 = n35511 & n25418;
  assign n25423 = ~n25256 & n25421;
  assign n25424 = ~n25419 & ~n35610;
  assign n25425 = ~n24633 & ~n24635;
  assign n25426 = ~n25256 & n25425;
  assign n25427 = ~n35506 & ~n25426;
  assign n25428 = ~n24635 & n35506;
  assign n25429 = ~n24633 & n25428;
  assign n25430 = n35506 & n25426;
  assign n25431 = ~n25256 & n25429;
  assign n25432 = ~n25427 & ~n35611;
  assign n25433 = ~n24597 & ~n24599;
  assign n25434 = ~n25256 & n25433;
  assign n25435 = ~n35500 & ~n25434;
  assign n25436 = ~n24599 & n35500;
  assign n25437 = ~n24597 & n25436;
  assign n25438 = n35500 & n25434;
  assign n25439 = ~n25256 & n25437;
  assign n25440 = ~n25435 & ~n35612;
  assign n25441 = ~n24566 & ~n24568;
  assign n25442 = ~n25256 & n25441;
  assign n25443 = ~n35496 & ~n25442;
  assign n25444 = ~n24568 & n35496;
  assign n25445 = ~n24566 & n25444;
  assign n25446 = n35496 & n25442;
  assign n25447 = ~n25256 & n25445;
  assign n25448 = ~n25443 & ~n35613;
  assign n25449 = ~n24530 & ~n24532;
  assign n25450 = ~n25256 & n25449;
  assign n25451 = ~n35490 & ~n25450;
  assign n25452 = ~n24532 & n35490;
  assign n25453 = ~n24530 & n25452;
  assign n25454 = n35490 & n25450;
  assign n25455 = ~n25256 & n25453;
  assign n25456 = ~n25451 & ~n35614;
  assign n25457 = ~n24496 & ~n24498;
  assign n25458 = ~n25256 & n25457;
  assign n25459 = ~n35485 & ~n25458;
  assign n25460 = ~n24498 & n35485;
  assign n25461 = ~n24496 & n25460;
  assign n25462 = n35485 & n25458;
  assign n25463 = ~n25256 & n25461;
  assign n25464 = ~n25459 & ~n35615;
  assign n25465 = ~n24462 & ~n24464;
  assign n25466 = ~n25256 & n25465;
  assign n25467 = ~n35480 & ~n25466;
  assign n25468 = ~n24464 & n35480;
  assign n25469 = ~n24462 & n25468;
  assign n25470 = n35480 & n25466;
  assign n25471 = ~n25256 & n25469;
  assign n25472 = ~n25467 & ~n35616;
  assign n25473 = ~n24429 & ~n24431;
  assign n25474 = ~n25256 & n25473;
  assign n25475 = ~n35476 & ~n25474;
  assign n25476 = ~n24431 & n35476;
  assign n25477 = ~n24429 & n25476;
  assign n25478 = n35476 & n25474;
  assign n25479 = ~n25256 & n25477;
  assign n25480 = ~n25475 & ~n35617;
  assign n25481 = ~n24395 & ~n24397;
  assign n25482 = ~n25256 & n25481;
  assign n25483 = ~n35471 & ~n25482;
  assign n25484 = ~n24397 & n35471;
  assign n25485 = ~n24395 & n25484;
  assign n25486 = n35471 & n25482;
  assign n25487 = ~n25256 & n25485;
  assign n25488 = ~n25483 & ~n35618;
  assign n25489 = ~n24368 & ~n24370;
  assign n25490 = ~n25256 & n25489;
  assign n25491 = ~n24379 & ~n25490;
  assign n25492 = ~n24370 & n24379;
  assign n25493 = ~n24368 & n25492;
  assign n25494 = n24379 & n25490;
  assign n25495 = ~n25256 & n25493;
  assign n25496 = ~n25491 & ~n35619;
  assign n25497 = ~pi14  & ~n25256;
  assign n25498 = ~pi15  & n25497;
  assign n25499 = n24345 & ~n25256;
  assign n25500 = ~n24331 & ~n25254;
  assign n25501 = ~n35589 & n25500;
  assign n25502 = ~n25248 & n25501;
  assign n25503 = ~n35620 & ~n25502;
  assign n25504 = pi16  & ~n25503;
  assign n25505 = ~pi16  & ~n25502;
  assign n25506 = ~pi16  & n25503;
  assign n25507 = ~n35620 & n25505;
  assign n25508 = ~n25504 & ~n35621;
  assign n25509 = pi14  & ~n25256;
  assign n25510 = ~pi12  & ~pi13 ;
  assign n25511 = ~pi14  & n25510;
  assign n25512 = ~n23498 & ~n35465;
  assign n25513 = ~n23499 & n25512;
  assign n25514 = ~n23515 & n25513;
  assign n25515 = ~n35358 & n25514;
  assign n25516 = n35356 & n23517;
  assign n25517 = ~n23509 & n25515;
  assign n25518 = ~n25511 & ~n35622;
  assign n25519 = ~n24329 & n25518;
  assign n25520 = ~n35461 & n25519;
  assign n25521 = ~n24323 & n25520;
  assign n25522 = ~n25509 & ~n25511;
  assign n25523 = n24331 & n25522;
  assign n25524 = ~n25509 & n25521;
  assign n25525 = pi15  & ~n25497;
  assign n25526 = ~n35620 & ~n25525;
  assign n25527 = ~n35623 & n25526;
  assign n25528 = ~n24331 & ~n25522;
  assign n25529 = n23517 & ~n25528;
  assign n25530 = ~n25527 & ~n25528;
  assign n25531 = n23517 & n25530;
  assign n25532 = ~n25527 & n25529;
  assign n25533 = ~n25508 & ~n35624;
  assign n25534 = ~n23517 & ~n25530;
  assign n25535 = n22625 & ~n25534;
  assign n25536 = ~n25533 & n25535;
  assign n25537 = ~n24348 & ~n35466;
  assign n25538 = ~n25256 & n25537;
  assign n25539 = n24353 & ~n25538;
  assign n25540 = ~n24353 & n25537;
  assign n25541 = ~n24353 & n25538;
  assign n25542 = ~n25256 & n25540;
  assign n25543 = ~n25539 & ~n35625;
  assign n25544 = ~n25536 & ~n25543;
  assign n25545 = ~n25533 & ~n25534;
  assign n25546 = ~n22625 & ~n25545;
  assign n25547 = n21842 & ~n25546;
  assign n25548 = ~n25544 & ~n25546;
  assign n25549 = n21842 & n25548;
  assign n25550 = ~n25544 & n25547;
  assign n25551 = ~n25496 & ~n35626;
  assign n25552 = ~n21842 & ~n25548;
  assign n25553 = n20986 & ~n25552;
  assign n25554 = ~n25551 & n25553;
  assign n25555 = ~n24382 & ~n35468;
  assign n25556 = ~n25256 & n25555;
  assign n25557 = n24392 & ~n25556;
  assign n25558 = ~n24392 & n25556;
  assign n25559 = ~n24382 & n24392;
  assign n25560 = ~n35468 & n25559;
  assign n25561 = n24392 & n25556;
  assign n25562 = ~n25256 & n25560;
  assign n25563 = ~n24392 & ~n25556;
  assign n25564 = ~n35627 & ~n25563;
  assign n25565 = ~n25557 & ~n25558;
  assign n25566 = ~n25554 & ~n35628;
  assign n25567 = ~n25551 & ~n25552;
  assign n25568 = ~n20986 & ~n25567;
  assign n25569 = n20229 & ~n25568;
  assign n25570 = ~n25566 & ~n25568;
  assign n25571 = n20229 & n25570;
  assign n25572 = ~n25566 & n25569;
  assign n25573 = ~n25488 & ~n35629;
  assign n25574 = ~n20229 & ~n25570;
  assign n25575 = n19401 & ~n25574;
  assign n25576 = ~n25573 & n25575;
  assign n25577 = ~n24412 & ~n35472;
  assign n25578 = ~n25256 & n25577;
  assign n25579 = ~n35474 & n25578;
  assign n25580 = n35474 & ~n25578;
  assign n25581 = ~n24412 & n35474;
  assign n25582 = ~n35472 & n25581;
  assign n25583 = ~n25256 & n25582;
  assign n25584 = ~n35474 & ~n25578;
  assign n25585 = ~n25583 & ~n25584;
  assign n25586 = ~n25579 & ~n25580;
  assign n25587 = ~n25576 & ~n35630;
  assign n25588 = ~n25573 & ~n25574;
  assign n25589 = ~n19401 & ~n25588;
  assign n25590 = n18676 & ~n25589;
  assign n25591 = ~n25587 & ~n25589;
  assign n25592 = n18676 & n25591;
  assign n25593 = ~n25587 & n25590;
  assign n25594 = ~n25480 & ~n35631;
  assign n25595 = ~n18676 & ~n25591;
  assign n25596 = n17885 & ~n25595;
  assign n25597 = ~n25594 & n25596;
  assign n25598 = ~n24446 & ~n35477;
  assign n25599 = ~n25256 & n25598;
  assign n25600 = ~n35478 & ~n25599;
  assign n25601 = ~n24446 & n35478;
  assign n25602 = ~n35477 & n25601;
  assign n25603 = n35478 & n25599;
  assign n25604 = ~n25256 & n25602;
  assign n25605 = n35478 & ~n25599;
  assign n25606 = ~n35478 & n25599;
  assign n25607 = ~n25605 & ~n25606;
  assign n25608 = ~n25600 & ~n35632;
  assign n25609 = ~n25597 & n35633;
  assign n25610 = ~n25594 & ~n25595;
  assign n25611 = ~n17885 & ~n25610;
  assign n25612 = n17187 & ~n25611;
  assign n25613 = ~n25609 & ~n25611;
  assign n25614 = n17187 & n25613;
  assign n25615 = ~n25609 & n25612;
  assign n25616 = ~n25472 & ~n35634;
  assign n25617 = ~n17187 & ~n25613;
  assign n25618 = n16428 & ~n25617;
  assign n25619 = ~n25616 & n25618;
  assign n25620 = ~n24479 & ~n35481;
  assign n25621 = ~n25256 & n25620;
  assign n25622 = n35483 & ~n25621;
  assign n25623 = ~n24479 & ~n35483;
  assign n25624 = ~n35481 & n25623;
  assign n25625 = ~n35483 & n25621;
  assign n25626 = ~n25256 & n25624;
  assign n25627 = n35483 & n25621;
  assign n25628 = ~n35483 & ~n25621;
  assign n25629 = ~n25627 & ~n25628;
  assign n25630 = ~n25622 & ~n35635;
  assign n25631 = ~n25619 & n35636;
  assign n25632 = ~n25616 & ~n25617;
  assign n25633 = ~n16428 & ~n25632;
  assign n25634 = n15760 & ~n25633;
  assign n25635 = ~n25631 & ~n25633;
  assign n25636 = n15760 & n25635;
  assign n25637 = ~n25631 & n25634;
  assign n25638 = ~n25464 & ~n35637;
  assign n25639 = ~n15760 & ~n25635;
  assign n25640 = n15033 & ~n25639;
  assign n25641 = ~n25638 & n25640;
  assign n25642 = ~n24513 & ~n35486;
  assign n25643 = ~n24513 & ~n25256;
  assign n25644 = ~n35486 & n25643;
  assign n25645 = ~n25256 & n25642;
  assign n25646 = ~n35488 & ~n35638;
  assign n25647 = n24528 & n25643;
  assign n25648 = n35488 & n35638;
  assign n25649 = ~n24513 & ~n35488;
  assign n25650 = ~n35486 & n25649;
  assign n25651 = ~n25256 & n25650;
  assign n25652 = n35488 & ~n35638;
  assign n25653 = ~n25651 & ~n25652;
  assign n25654 = ~n25646 & ~n35639;
  assign n25655 = ~n25641 & ~n35640;
  assign n25656 = ~n25638 & ~n25639;
  assign n25657 = ~n15033 & ~n25656;
  assign n25658 = n14394 & ~n25657;
  assign n25659 = ~n25655 & ~n25657;
  assign n25660 = n14394 & n25659;
  assign n25661 = ~n25655 & n25658;
  assign n25662 = ~n25456 & ~n35641;
  assign n25663 = ~n14394 & ~n25659;
  assign n25664 = n13704 & ~n25663;
  assign n25665 = ~n25662 & n25664;
  assign n25666 = ~n24547 & ~n35491;
  assign n25667 = ~n25256 & n25666;
  assign n25668 = ~n35494 & ~n25667;
  assign n25669 = ~n24547 & n35494;
  assign n25670 = ~n35491 & n25669;
  assign n25671 = n35494 & n25667;
  assign n25672 = ~n25256 & n25670;
  assign n25673 = ~n25668 & ~n35642;
  assign n25674 = ~n25665 & ~n25673;
  assign n25675 = ~n25662 & ~n25663;
  assign n25676 = ~n13704 & ~n25675;
  assign n25677 = n13099 & ~n25676;
  assign n25678 = ~n25674 & ~n25676;
  assign n25679 = n13099 & n25678;
  assign n25680 = ~n25674 & n25677;
  assign n25681 = ~n25448 & ~n35643;
  assign n25682 = ~n13099 & ~n25678;
  assign n25683 = n12442 & ~n25682;
  assign n25684 = ~n25681 & n25683;
  assign n25685 = ~n24583 & ~n35497;
  assign n25686 = ~n24583 & ~n25256;
  assign n25687 = ~n35497 & n25686;
  assign n25688 = ~n25256 & n25685;
  assign n25689 = n24594 & ~n35644;
  assign n25690 = n24595 & n25686;
  assign n25691 = ~n24594 & n35644;
  assign n25692 = ~n24583 & n24594;
  assign n25693 = ~n35497 & n25692;
  assign n25694 = ~n25256 & n25693;
  assign n25695 = ~n24594 & ~n35644;
  assign n25696 = ~n25694 & ~n25695;
  assign n25697 = ~n25689 & ~n35645;
  assign n25698 = ~n25684 & ~n35646;
  assign n25699 = ~n25681 & ~n25682;
  assign n25700 = ~n12442 & ~n25699;
  assign n25701 = n11858 & ~n25700;
  assign n25702 = ~n25698 & ~n25700;
  assign n25703 = n11858 & n25702;
  assign n25704 = ~n25698 & n25701;
  assign n25705 = ~n25440 & ~n35647;
  assign n25706 = ~n11858 & ~n25702;
  assign n25707 = n11229 & ~n25706;
  assign n25708 = ~n25705 & n25707;
  assign n25709 = ~n24614 & ~n35501;
  assign n25710 = ~n25256 & n25709;
  assign n25711 = ~n35504 & n25710;
  assign n25712 = n35504 & ~n25710;
  assign n25713 = ~n24614 & n35504;
  assign n25714 = ~n35501 & n25713;
  assign n25715 = n35504 & n25710;
  assign n25716 = ~n25256 & n25714;
  assign n25717 = ~n35504 & ~n25710;
  assign n25718 = ~n35648 & ~n25717;
  assign n25719 = ~n25711 & ~n25712;
  assign n25720 = ~n25708 & ~n35649;
  assign n25721 = ~n25705 & ~n25706;
  assign n25722 = ~n11229 & ~n25721;
  assign n25723 = n10681 & ~n25722;
  assign n25724 = ~n25720 & ~n25722;
  assign n25725 = n10681 & n25724;
  assign n25726 = ~n25720 & n25723;
  assign n25727 = ~n25432 & ~n35650;
  assign n25728 = ~n10681 & ~n25724;
  assign n25729 = n10086 & ~n25728;
  assign n25730 = ~n25727 & n25729;
  assign n25731 = ~n24650 & ~n35507;
  assign n25732 = ~n24650 & ~n25256;
  assign n25733 = ~n35507 & n25732;
  assign n25734 = ~n25256 & n25731;
  assign n25735 = n35509 & ~n35651;
  assign n25736 = n24665 & n25732;
  assign n25737 = ~n35509 & n35651;
  assign n25738 = ~n24650 & n35509;
  assign n25739 = ~n35507 & n25738;
  assign n25740 = ~n25256 & n25739;
  assign n25741 = ~n35509 & ~n35651;
  assign n25742 = ~n25740 & ~n25741;
  assign n25743 = ~n25735 & ~n35652;
  assign n25744 = ~n25730 & ~n35653;
  assign n25745 = ~n25727 & ~n25728;
  assign n25746 = ~n10086 & ~n25745;
  assign n25747 = n9565 & ~n25746;
  assign n25748 = ~n25744 & ~n25746;
  assign n25749 = n9565 & n25748;
  assign n25750 = ~n25744 & n25747;
  assign n25751 = ~n25424 & ~n35654;
  assign n25752 = ~n9565 & ~n25748;
  assign n25753 = n8998 & ~n25752;
  assign n25754 = ~n25751 & n25753;
  assign n25755 = ~n25416 & ~n25754;
  assign n25756 = ~n25751 & ~n25752;
  assign n25757 = ~n8998 & ~n25756;
  assign n25758 = n8506 & ~n25757;
  assign n25759 = ~n25755 & ~n25757;
  assign n25760 = n8506 & n25759;
  assign n25761 = ~n25755 & n25758;
  assign n25762 = ~n25408 & ~n35655;
  assign n25763 = ~n8506 & ~n25759;
  assign n25764 = n7975 & ~n25763;
  assign n25765 = ~n25762 & n25764;
  assign n25766 = ~n24720 & ~n35519;
  assign n25767 = ~n24720 & ~n25256;
  assign n25768 = ~n35519 & n25767;
  assign n25769 = ~n25256 & n25766;
  assign n25770 = n24728 & ~n35656;
  assign n25771 = n24732 & n25767;
  assign n25772 = ~n24720 & n24728;
  assign n25773 = ~n35519 & n25772;
  assign n25774 = ~n25256 & n25773;
  assign n25775 = ~n24728 & ~n35656;
  assign n25776 = ~n25774 & ~n25775;
  assign n25777 = ~n25770 & ~n25771;
  assign n25778 = ~n25765 & ~n35657;
  assign n25779 = ~n25762 & ~n25763;
  assign n25780 = ~n7975 & ~n25779;
  assign n25781 = n7512 & ~n25780;
  assign n25782 = ~n25778 & ~n25780;
  assign n25783 = n7512 & n25782;
  assign n25784 = ~n25778 & n25781;
  assign n25785 = ~n25400 & ~n35658;
  assign n25786 = ~n7512 & ~n25782;
  assign n25787 = n7015 & ~n25786;
  assign n25788 = ~n25785 & n25787;
  assign n25789 = ~n25392 & ~n25788;
  assign n25790 = ~n25785 & ~n25786;
  assign n25791 = ~n7015 & ~n25790;
  assign n25792 = n6579 & ~n25791;
  assign n25793 = ~n25789 & ~n25791;
  assign n25794 = n6579 & n25793;
  assign n25795 = ~n25789 & n25792;
  assign n25796 = ~n25384 & ~n35659;
  assign n25797 = ~n6579 & ~n25793;
  assign n25798 = n6117 & ~n25797;
  assign n25799 = ~n25796 & n25798;
  assign n25800 = ~n24786 & ~n35528;
  assign n25801 = ~n24786 & ~n25256;
  assign n25802 = ~n35528 & n25801;
  assign n25803 = ~n25256 & n25800;
  assign n25804 = n24794 & ~n35660;
  assign n25805 = n24798 & n25801;
  assign n25806 = ~n24786 & n24794;
  assign n25807 = ~n35528 & n25806;
  assign n25808 = ~n25256 & n25807;
  assign n25809 = ~n24794 & ~n35660;
  assign n25810 = ~n25808 & ~n25809;
  assign n25811 = ~n25804 & ~n25805;
  assign n25812 = ~n25799 & ~n35661;
  assign n25813 = ~n25796 & ~n25797;
  assign n25814 = ~n6117 & ~n25813;
  assign n25815 = n5708 & ~n25814;
  assign n25816 = ~n25812 & ~n25814;
  assign n25817 = n5708 & n25816;
  assign n25818 = ~n25812 & n25815;
  assign n25819 = ~n25376 & ~n35662;
  assign n25820 = ~n5708 & ~n25816;
  assign n25821 = n5278 & ~n25820;
  assign n25822 = ~n25819 & n25821;
  assign n25823 = ~n25368 & ~n25822;
  assign n25824 = ~n25819 & ~n25820;
  assign n25825 = ~n5278 & ~n25824;
  assign n25826 = n4903 & ~n25825;
  assign n25827 = ~n25823 & ~n25825;
  assign n25828 = n4903 & n25827;
  assign n25829 = ~n25823 & n25826;
  assign n25830 = ~n25360 & ~n35663;
  assign n25831 = ~n4903 & ~n25827;
  assign n25832 = n4508 & ~n25831;
  assign n25833 = ~n25830 & n25832;
  assign n25834 = ~n24852 & ~n35537;
  assign n25835 = ~n24852 & ~n25256;
  assign n25836 = ~n35537 & n25835;
  assign n25837 = ~n25256 & n25834;
  assign n25838 = n24860 & ~n35664;
  assign n25839 = n24864 & n25835;
  assign n25840 = ~n24852 & n24860;
  assign n25841 = ~n35537 & n25840;
  assign n25842 = ~n25256 & n25841;
  assign n25843 = ~n24860 & ~n35664;
  assign n25844 = ~n25842 & ~n25843;
  assign n25845 = ~n25838 & ~n25839;
  assign n25846 = ~n25833 & ~n35665;
  assign n25847 = ~n25830 & ~n25831;
  assign n25848 = ~n4508 & ~n25847;
  assign n25849 = n4155 & ~n25848;
  assign n25850 = ~n25846 & ~n25848;
  assign n25851 = n4155 & n25850;
  assign n25852 = ~n25846 & n25849;
  assign n25853 = ~n25352 & ~n35666;
  assign n25854 = ~n4155 & ~n25850;
  assign n25855 = n3788 & ~n25854;
  assign n25856 = ~n25853 & n25855;
  assign n25857 = ~n25344 & ~n25856;
  assign n25858 = ~n25853 & ~n25854;
  assign n25859 = ~n3788 & ~n25858;
  assign n25860 = n3473 & ~n25859;
  assign n25861 = ~n25857 & ~n25859;
  assign n25862 = n3473 & n25861;
  assign n25863 = ~n25857 & n25860;
  assign n25864 = ~n25336 & ~n35667;
  assign n25865 = ~n3473 & ~n25861;
  assign n25866 = n3140 & ~n25865;
  assign n25867 = ~n25864 & n25866;
  assign n25868 = ~n24918 & ~n35546;
  assign n25869 = ~n24918 & ~n25256;
  assign n25870 = ~n35546 & n25869;
  assign n25871 = ~n25256 & n25868;
  assign n25872 = n24926 & ~n35668;
  assign n25873 = n24930 & n25869;
  assign n25874 = ~n24918 & n24926;
  assign n25875 = ~n35546 & n25874;
  assign n25876 = ~n25256 & n25875;
  assign n25877 = ~n24926 & ~n35668;
  assign n25878 = ~n25876 & ~n25877;
  assign n25879 = ~n25872 & ~n25873;
  assign n25880 = ~n25867 & ~n35669;
  assign n25881 = ~n25864 & ~n25865;
  assign n25882 = ~n3140 & ~n25881;
  assign n25883 = n2855 & ~n25882;
  assign n25884 = ~n25880 & ~n25882;
  assign n25885 = n2855 & n25884;
  assign n25886 = ~n25880 & n25883;
  assign n25887 = ~n25328 & ~n35670;
  assign n25888 = ~n2855 & ~n25884;
  assign n25889 = n2556 & ~n25888;
  assign n25890 = ~n25887 & n25889;
  assign n25891 = ~n25320 & ~n25890;
  assign n25892 = ~n25887 & ~n25888;
  assign n25893 = ~n2556 & ~n25892;
  assign n25894 = n2301 & ~n25893;
  assign n25895 = ~n25891 & ~n25893;
  assign n25896 = n2301 & n25895;
  assign n25897 = ~n25891 & n25894;
  assign n25898 = ~n25312 & ~n35671;
  assign n25899 = ~n2301 & ~n25895;
  assign n25900 = n2038 & ~n25899;
  assign n25901 = ~n25898 & n25900;
  assign n25902 = ~n24984 & ~n35555;
  assign n25903 = ~n24984 & ~n25256;
  assign n25904 = ~n35555 & n25903;
  assign n25905 = ~n25256 & n25902;
  assign n25906 = n24992 & ~n35672;
  assign n25907 = n24996 & n25903;
  assign n25908 = ~n24984 & n24992;
  assign n25909 = ~n35555 & n25908;
  assign n25910 = ~n25256 & n25909;
  assign n25911 = ~n24992 & ~n35672;
  assign n25912 = ~n25910 & ~n25911;
  assign n25913 = ~n25906 & ~n25907;
  assign n25914 = ~n25901 & ~n35673;
  assign n25915 = ~n25898 & ~n25899;
  assign n25916 = ~n2038 & ~n25915;
  assign n25917 = n1812 & ~n25916;
  assign n25918 = ~n25914 & ~n25916;
  assign n25919 = n1812 & n25918;
  assign n25920 = ~n25914 & n25917;
  assign n25921 = ~n25304 & ~n35674;
  assign n25922 = ~n1812 & ~n25918;
  assign n25923 = n1582 & ~n25922;
  assign n25924 = ~n25921 & n25923;
  assign n25925 = ~n25296 & ~n25924;
  assign n25926 = ~n25921 & ~n25922;
  assign n25927 = ~n1582 & ~n25926;
  assign n25928 = n1388 & ~n25927;
  assign n25929 = ~n25925 & ~n25927;
  assign n25930 = n1388 & n25929;
  assign n25931 = ~n25925 & n25928;
  assign n25932 = ~n25288 & ~n35675;
  assign n25933 = ~n1388 & ~n25929;
  assign n25934 = n1192 & ~n25933;
  assign n25935 = ~n25932 & n25934;
  assign n25936 = ~n25050 & ~n35564;
  assign n25937 = ~n25050 & ~n25256;
  assign n25938 = ~n35564 & n25937;
  assign n25939 = ~n25256 & n25936;
  assign n25940 = n25058 & ~n35676;
  assign n25941 = n25062 & n25937;
  assign n25942 = ~n25050 & n25058;
  assign n25943 = ~n35564 & n25942;
  assign n25944 = ~n25256 & n25943;
  assign n25945 = ~n25058 & ~n35676;
  assign n25946 = ~n25944 & ~n25945;
  assign n25947 = ~n25940 & ~n25941;
  assign n25948 = ~n25935 & ~n35677;
  assign n25949 = ~n25932 & ~n25933;
  assign n25950 = ~n1192 & ~n25949;
  assign n25951 = n1028 & ~n25950;
  assign n25952 = ~n25948 & ~n25950;
  assign n25953 = n1028 & n25952;
  assign n25954 = ~n25948 & n25951;
  assign n25955 = ~n25280 & ~n35678;
  assign n25956 = ~n1028 & ~n25952;
  assign n25957 = n866 & ~n25956;
  assign n25958 = ~n25955 & n25957;
  assign n25959 = ~n25272 & ~n25958;
  assign n25960 = ~n25955 & ~n25956;
  assign n25961 = ~n866 & ~n25960;
  assign n25962 = n730 & ~n25961;
  assign n25963 = ~n25959 & ~n25961;
  assign n25964 = n730 & n25963;
  assign n25965 = ~n25959 & n25962;
  assign n25966 = ~n25099 & ~n25101;
  assign n25967 = ~n25256 & n25966;
  assign n25968 = ~n35570 & n25967;
  assign n25969 = n35570 & ~n25967;
  assign n25970 = ~n25101 & n35570;
  assign n25971 = ~n25099 & n25970;
  assign n25972 = ~n25256 & n25971;
  assign n25973 = ~n35570 & ~n25967;
  assign n25974 = ~n25972 & ~n25973;
  assign n25975 = ~n25968 & ~n25969;
  assign n25976 = ~n35679 & ~n35680;
  assign n25977 = ~n730 & ~n25963;
  assign n25978 = ~n25976 & ~n25977;
  assign n25979 = ~n602 & ~n25978;
  assign n25980 = n602 & ~n25977;
  assign n25981 = ~n25976 & n25980;
  assign n25982 = ~n25114 & ~n35573;
  assign n25983 = ~n25256 & n25982;
  assign n25984 = ~n35572 & ~n25983;
  assign n25985 = n35572 & n25983;
  assign n25986 = ~n25114 & ~n35572;
  assign n25987 = ~n35573 & n25986;
  assign n25988 = ~n25256 & n25987;
  assign n25989 = n35572 & ~n25983;
  assign n25990 = ~n25988 & ~n25989;
  assign n25991 = ~n25984 & ~n25985;
  assign n25992 = ~n25981 & ~n35681;
  assign n25993 = ~n25979 & ~n25992;
  assign n25994 = ~n497 & ~n25993;
  assign n25995 = n497 & ~n25979;
  assign n25996 = n497 & n25993;
  assign n25997 = ~n25992 & n25995;
  assign n25998 = ~n25264 & ~n35682;
  assign n25999 = ~n25994 & ~n25998;
  assign n26000 = ~n403 & ~n25999;
  assign n26001 = n403 & ~n25994;
  assign n26002 = ~n25998 & n26001;
  assign n26003 = ~n25136 & ~n35575;
  assign n26004 = ~n25136 & ~n25256;
  assign n26005 = ~n35575 & n26004;
  assign n26006 = ~n25256 & n26003;
  assign n26007 = n25144 & ~n35683;
  assign n26008 = n25148 & n26004;
  assign n26009 = ~n25136 & n25144;
  assign n26010 = ~n35575 & n26009;
  assign n26011 = ~n25256 & n26010;
  assign n26012 = ~n25144 & ~n35683;
  assign n26013 = ~n26011 & ~n26012;
  assign n26014 = ~n26007 & ~n26008;
  assign n26015 = ~n26002 & ~n35684;
  assign n26016 = ~n26000 & ~n26015;
  assign n26017 = ~n330 & ~n26016;
  assign n26018 = ~n25150 & ~n25152;
  assign n26019 = ~n25256 & n26018;
  assign n26020 = ~n35577 & ~n26019;
  assign n26021 = ~n25152 & n35577;
  assign n26022 = ~n25150 & n26021;
  assign n26023 = n35577 & n26019;
  assign n26024 = ~n25256 & n26022;
  assign n26025 = ~n26020 & ~n35685;
  assign n26026 = n330 & ~n26000;
  assign n26027 = n330 & n26016;
  assign n26028 = ~n26015 & n26026;
  assign n26029 = ~n26025 & ~n35686;
  assign n26030 = ~n26017 & ~n26029;
  assign n26031 = ~n271 & ~n26030;
  assign n26032 = n271 & ~n26017;
  assign n26033 = ~n26029 & n26032;
  assign n26034 = ~n25167 & ~n35579;
  assign n26035 = ~n25167 & ~n25256;
  assign n26036 = ~n35579 & n26035;
  assign n26037 = ~n25256 & n26034;
  assign n26038 = n25175 & ~n35687;
  assign n26039 = n25179 & n26035;
  assign n26040 = ~n25167 & n25175;
  assign n26041 = ~n35579 & n26040;
  assign n26042 = ~n25256 & n26041;
  assign n26043 = ~n25175 & ~n35687;
  assign n26044 = ~n26042 & ~n26043;
  assign n26045 = ~n26038 & ~n26039;
  assign n26046 = ~n26033 & ~n35688;
  assign n26047 = ~n26031 & ~n26046;
  assign n26048 = ~n217 & ~n26047;
  assign n26049 = ~n25181 & ~n25183;
  assign n26050 = ~n25256 & n26049;
  assign n26051 = ~n35581 & ~n26050;
  assign n26052 = ~n25183 & n35581;
  assign n26053 = ~n25181 & n26052;
  assign n26054 = n35581 & n26050;
  assign n26055 = ~n25256 & n26053;
  assign n26056 = ~n26051 & ~n35689;
  assign n26057 = n217 & ~n26031;
  assign n26058 = n217 & n26047;
  assign n26059 = ~n26046 & n26057;
  assign n26060 = ~n26056 & ~n35690;
  assign n26061 = ~n26048 & ~n26060;
  assign n26062 = ~n198 & ~n26061;
  assign n26063 = ~n25198 & ~n35582;
  assign n26064 = ~n25256 & n26063;
  assign n26065 = ~n35584 & ~n26064;
  assign n26066 = ~n25198 & n35584;
  assign n26067 = ~n35582 & n26066;
  assign n26068 = n35584 & n26064;
  assign n26069 = ~n25256 & n26067;
  assign n26070 = ~n26065 & ~n35691;
  assign n26071 = n198 & ~n26048;
  assign n26072 = ~n26060 & n26071;
  assign n26073 = ~n26070 & ~n26072;
  assign n26074 = ~n26062 & ~n26073;
  assign n26075 = ~n25216 & ~n25218;
  assign n26076 = ~n25256 & n26075;
  assign n26077 = ~n35586 & ~n26076;
  assign n26078 = ~n25218 & n35586;
  assign n26079 = ~n25216 & n26078;
  assign n26080 = n35586 & n26076;
  assign n26081 = ~n25256 & n26079;
  assign n26082 = ~n26077 & ~n35692;
  assign n26083 = ~n25232 & ~n25240;
  assign n26084 = ~n25240 & ~n25256;
  assign n26085 = ~n25232 & n26084;
  assign n26086 = ~n25256 & n26083;
  assign n26087 = ~n35589 & ~n35693;
  assign n26088 = ~n26082 & n26087;
  assign n26089 = ~n26074 & n26088;
  assign n26090 = n193 & ~n26089;
  assign n26091 = ~n26062 & n26082;
  assign n26092 = n26074 & n26082;
  assign n26093 = ~n26073 & n26091;
  assign n26094 = n25232 & ~n26084;
  assign n26095 = ~n193 & ~n26083;
  assign n26096 = ~n26094 & n26095;
  assign n26097 = ~n35694 & ~n26096;
  assign n26098 = ~n26090 & n26097;
  assign n26099 = ~n25994 & ~n35682;
  assign n26100 = ~n25994 & ~n26098;
  assign n26101 = ~n35682 & n26100;
  assign n26102 = ~n26098 & n26099;
  assign n26103 = n25264 & ~n35695;
  assign n26104 = n25998 & n26100;
  assign n26105 = n25264 & ~n35682;
  assign n26106 = ~n25994 & n26105;
  assign n26107 = ~n26098 & n26106;
  assign n26108 = ~n25264 & ~n35695;
  assign n26109 = ~n26107 & ~n26108;
  assign n26110 = ~n26103 & ~n26104;
  assign n26111 = pi12  & ~n26098;
  assign n26112 = ~pi10  & ~pi11 ;
  assign n26113 = ~pi12  & n26112;
  assign n26114 = ~n26111 & ~n26113;
  assign n26115 = ~n25256 & ~n26114;
  assign n26116 = ~pi12  & ~n26098;
  assign n26117 = pi13  & ~n26116;
  assign n26118 = ~pi13  & n26116;
  assign n26119 = n25510 & ~n26098;
  assign n26120 = ~n26117 & ~n35697;
  assign n26121 = ~n35459 & ~n35622;
  assign n26122 = ~n24310 & n26121;
  assign n26123 = ~n24329 & n26122;
  assign n26124 = ~n35461 & n26123;
  assign n26125 = n24315 & n24331;
  assign n26126 = ~n24323 & n26124;
  assign n26127 = ~n26113 & ~n35698;
  assign n26128 = ~n25254 & n26127;
  assign n26129 = ~n35589 & n26128;
  assign n26130 = ~n25248 & n26129;
  assign n26131 = n25256 & n26114;
  assign n26132 = ~n26111 & n26130;
  assign n26133 = n26120 & ~n35699;
  assign n26134 = ~n26115 & ~n26133;
  assign n26135 = ~n24331 & ~n26134;
  assign n26136 = n24331 & ~n26115;
  assign n26137 = ~n26133 & n26136;
  assign n26138 = ~n25256 & ~n26096;
  assign n26139 = ~n35694 & n26138;
  assign n26140 = ~n26090 & n26139;
  assign n26141 = ~n35697 & ~n26140;
  assign n26142 = pi14  & ~n26141;
  assign n26143 = ~pi14  & ~n26140;
  assign n26144 = ~pi14  & n26141;
  assign n26145 = ~n35697 & n26143;
  assign n26146 = ~n26142 & ~n35700;
  assign n26147 = ~n26137 & ~n26146;
  assign n26148 = ~n26135 & ~n26147;
  assign n26149 = ~n23517 & ~n26148;
  assign n26150 = n23517 & ~n26135;
  assign n26151 = ~n26147 & n26150;
  assign n26152 = n23517 & n26148;
  assign n26153 = ~n35623 & ~n25528;
  assign n26154 = ~n26098 & n26153;
  assign n26155 = n25526 & ~n26154;
  assign n26156 = ~n25526 & n26153;
  assign n26157 = ~n25526 & n26154;
  assign n26158 = ~n26098 & n26156;
  assign n26159 = ~n26155 & ~n35702;
  assign n26160 = ~n35701 & ~n26159;
  assign n26161 = ~n26149 & ~n26160;
  assign n26162 = ~n22625 & ~n26161;
  assign n26163 = n22625 & ~n26149;
  assign n26164 = ~n26160 & n26163;
  assign n26165 = ~n35624 & ~n25534;
  assign n26166 = ~n25534 & ~n26098;
  assign n26167 = ~n35624 & n26166;
  assign n26168 = ~n26098 & n26165;
  assign n26169 = n25508 & ~n35703;
  assign n26170 = n25533 & n26166;
  assign n26171 = n25508 & ~n35624;
  assign n26172 = ~n25534 & n26171;
  assign n26173 = ~n26098 & n26172;
  assign n26174 = ~n25508 & ~n35703;
  assign n26175 = ~n26173 & ~n26174;
  assign n26176 = ~n26169 & ~n26170;
  assign n26177 = ~n26164 & ~n35704;
  assign n26178 = ~n26162 & ~n26177;
  assign n26179 = ~n21842 & ~n26178;
  assign n26180 = n21842 & ~n26162;
  assign n26181 = ~n26177 & n26180;
  assign n26182 = n21842 & n26178;
  assign n26183 = ~n25536 & ~n25546;
  assign n26184 = ~n26098 & n26183;
  assign n26185 = n25543 & ~n26184;
  assign n26186 = ~n25543 & n26184;
  assign n26187 = n25543 & ~n25546;
  assign n26188 = ~n25536 & n26187;
  assign n26189 = n25543 & n26184;
  assign n26190 = ~n26098 & n26188;
  assign n26191 = ~n25543 & ~n26184;
  assign n26192 = ~n35706 & ~n26191;
  assign n26193 = ~n26185 & ~n26186;
  assign n26194 = ~n35705 & ~n35707;
  assign n26195 = ~n26179 & ~n26194;
  assign n26196 = ~n20986 & ~n26195;
  assign n26197 = n20986 & ~n26179;
  assign n26198 = ~n26194 & n26197;
  assign n26199 = ~n35626 & ~n25552;
  assign n26200 = ~n25552 & ~n26098;
  assign n26201 = ~n35626 & n26200;
  assign n26202 = ~n26098 & n26199;
  assign n26203 = n25496 & ~n35708;
  assign n26204 = n25551 & n26200;
  assign n26205 = n25496 & ~n35626;
  assign n26206 = ~n25552 & n26205;
  assign n26207 = ~n26098 & n26206;
  assign n26208 = ~n25496 & ~n35708;
  assign n26209 = ~n26207 & ~n26208;
  assign n26210 = ~n26203 & ~n26204;
  assign n26211 = ~n26198 & ~n35709;
  assign n26212 = ~n26196 & ~n26211;
  assign n26213 = ~n20229 & ~n26212;
  assign n26214 = n20229 & ~n26196;
  assign n26215 = ~n26211 & n26214;
  assign n26216 = n20229 & n26212;
  assign n26217 = ~n25554 & ~n25568;
  assign n26218 = ~n26098 & n26217;
  assign n26219 = ~n35628 & n26218;
  assign n26220 = n35628 & ~n26218;
  assign n26221 = n35628 & ~n25568;
  assign n26222 = ~n25554 & n26221;
  assign n26223 = ~n26098 & n26222;
  assign n26224 = ~n35628 & ~n26218;
  assign n26225 = ~n26223 & ~n26224;
  assign n26226 = ~n26219 & ~n26220;
  assign n26227 = ~n35710 & ~n35711;
  assign n26228 = ~n26213 & ~n26227;
  assign n26229 = ~n19401 & ~n26228;
  assign n26230 = n19401 & ~n26213;
  assign n26231 = ~n26227 & n26230;
  assign n26232 = ~n35629 & ~n25574;
  assign n26233 = ~n25574 & ~n26098;
  assign n26234 = ~n35629 & n26233;
  assign n26235 = ~n26098 & n26232;
  assign n26236 = n25488 & ~n35712;
  assign n26237 = n25573 & n26233;
  assign n26238 = n25488 & ~n35629;
  assign n26239 = ~n25574 & n26238;
  assign n26240 = ~n26098 & n26239;
  assign n26241 = ~n25488 & ~n35712;
  assign n26242 = ~n26240 & ~n26241;
  assign n26243 = ~n26236 & ~n26237;
  assign n26244 = ~n26231 & ~n35713;
  assign n26245 = ~n26229 & ~n26244;
  assign n26246 = ~n18676 & ~n26245;
  assign n26247 = n18676 & ~n26229;
  assign n26248 = ~n26244 & n26247;
  assign n26249 = n18676 & n26245;
  assign n26250 = ~n25576 & ~n25589;
  assign n26251 = ~n26098 & n26250;
  assign n26252 = ~n35630 & ~n26251;
  assign n26253 = n35630 & ~n25589;
  assign n26254 = ~n25576 & n26253;
  assign n26255 = n35630 & n26251;
  assign n26256 = ~n26098 & n26254;
  assign n26257 = n35630 & ~n26251;
  assign n26258 = ~n35630 & n26251;
  assign n26259 = ~n26257 & ~n26258;
  assign n26260 = ~n26252 & ~n35715;
  assign n26261 = ~n35714 & n35716;
  assign n26262 = ~n26246 & ~n26261;
  assign n26263 = ~n17885 & ~n26262;
  assign n26264 = n17885 & ~n26246;
  assign n26265 = ~n26261 & n26264;
  assign n26266 = ~n35631 & ~n25595;
  assign n26267 = ~n25595 & ~n26098;
  assign n26268 = ~n35631 & n26267;
  assign n26269 = ~n26098 & n26266;
  assign n26270 = n25480 & ~n35717;
  assign n26271 = n25594 & n26267;
  assign n26272 = n25480 & ~n35631;
  assign n26273 = ~n25595 & n26272;
  assign n26274 = ~n26098 & n26273;
  assign n26275 = ~n25480 & ~n35717;
  assign n26276 = ~n26274 & ~n26275;
  assign n26277 = ~n26270 & ~n26271;
  assign n26278 = ~n26265 & ~n35718;
  assign n26279 = ~n26263 & ~n26278;
  assign n26280 = ~n17187 & ~n26279;
  assign n26281 = n17187 & ~n26263;
  assign n26282 = ~n26278 & n26281;
  assign n26283 = n17187 & n26279;
  assign n26284 = ~n25597 & ~n25611;
  assign n26285 = ~n26098 & n26284;
  assign n26286 = n35633 & ~n26285;
  assign n26287 = ~n35633 & ~n25611;
  assign n26288 = ~n25597 & n26287;
  assign n26289 = ~n35633 & n26285;
  assign n26290 = ~n26098 & n26288;
  assign n26291 = n35633 & n26285;
  assign n26292 = ~n35633 & ~n26285;
  assign n26293 = ~n26291 & ~n26292;
  assign n26294 = ~n26286 & ~n35720;
  assign n26295 = ~n35719 & n35721;
  assign n26296 = ~n26280 & ~n26295;
  assign n26297 = ~n16428 & ~n26296;
  assign n26298 = n16428 & ~n26280;
  assign n26299 = ~n26295 & n26298;
  assign n26300 = ~n35634 & ~n25617;
  assign n26301 = ~n25617 & ~n26098;
  assign n26302 = ~n35634 & n26301;
  assign n26303 = ~n26098 & n26300;
  assign n26304 = n25472 & ~n35722;
  assign n26305 = n25616 & n26301;
  assign n26306 = n25472 & ~n35634;
  assign n26307 = ~n25617 & n26306;
  assign n26308 = ~n26098 & n26307;
  assign n26309 = ~n25472 & ~n35722;
  assign n26310 = ~n26308 & ~n26309;
  assign n26311 = ~n26304 & ~n26305;
  assign n26312 = ~n26299 & ~n35723;
  assign n26313 = ~n26297 & ~n26312;
  assign n26314 = ~n15760 & ~n26313;
  assign n26315 = n15760 & ~n26297;
  assign n26316 = ~n26312 & n26315;
  assign n26317 = n15760 & n26313;
  assign n26318 = ~n25619 & ~n25633;
  assign n26319 = ~n25633 & ~n26098;
  assign n26320 = ~n25619 & n26319;
  assign n26321 = ~n26098 & n26318;
  assign n26322 = ~n35636 & ~n35725;
  assign n26323 = n25631 & n26319;
  assign n26324 = n35636 & n35725;
  assign n26325 = ~n35636 & ~n25633;
  assign n26326 = ~n25619 & n26325;
  assign n26327 = ~n26098 & n26326;
  assign n26328 = n35636 & ~n35725;
  assign n26329 = ~n26327 & ~n26328;
  assign n26330 = ~n26322 & ~n35726;
  assign n26331 = ~n35724 & ~n35727;
  assign n26332 = ~n26314 & ~n26331;
  assign n26333 = ~n15033 & ~n26332;
  assign n26334 = n15033 & ~n26314;
  assign n26335 = ~n26331 & n26334;
  assign n26336 = ~n35637 & ~n25639;
  assign n26337 = ~n25639 & ~n26098;
  assign n26338 = ~n35637 & n26337;
  assign n26339 = ~n26098 & n26336;
  assign n26340 = n25464 & ~n35728;
  assign n26341 = n25638 & n26337;
  assign n26342 = n25464 & ~n35637;
  assign n26343 = ~n25639 & n26342;
  assign n26344 = ~n26098 & n26343;
  assign n26345 = ~n25464 & ~n35728;
  assign n26346 = ~n26344 & ~n26345;
  assign n26347 = ~n26340 & ~n26341;
  assign n26348 = ~n26335 & ~n35729;
  assign n26349 = ~n26333 & ~n26348;
  assign n26350 = ~n14394 & ~n26349;
  assign n26351 = n14394 & ~n26333;
  assign n26352 = ~n26348 & n26351;
  assign n26353 = n14394 & n26349;
  assign n26354 = ~n25641 & ~n25657;
  assign n26355 = ~n26098 & n26354;
  assign n26356 = ~n35640 & ~n26355;
  assign n26357 = n35640 & ~n25657;
  assign n26358 = ~n25641 & n26357;
  assign n26359 = n35640 & n26355;
  assign n26360 = ~n26098 & n26358;
  assign n26361 = ~n26356 & ~n35731;
  assign n26362 = ~n35730 & ~n26361;
  assign n26363 = ~n26350 & ~n26362;
  assign n26364 = ~n13704 & ~n26363;
  assign n26365 = n13704 & ~n26350;
  assign n26366 = ~n26362 & n26365;
  assign n26367 = ~n35641 & ~n25663;
  assign n26368 = ~n25663 & ~n26098;
  assign n26369 = ~n35641 & n26368;
  assign n26370 = ~n26098 & n26367;
  assign n26371 = n25456 & ~n35732;
  assign n26372 = n25662 & n26368;
  assign n26373 = n25456 & ~n35641;
  assign n26374 = ~n25663 & n26373;
  assign n26375 = ~n26098 & n26374;
  assign n26376 = ~n25456 & ~n35732;
  assign n26377 = ~n26375 & ~n26376;
  assign n26378 = ~n26371 & ~n26372;
  assign n26379 = ~n26366 & ~n35733;
  assign n26380 = ~n26364 & ~n26379;
  assign n26381 = ~n13099 & ~n26380;
  assign n26382 = n13099 & ~n26364;
  assign n26383 = ~n26379 & n26382;
  assign n26384 = n13099 & n26380;
  assign n26385 = ~n25665 & ~n25676;
  assign n26386 = ~n25676 & ~n26098;
  assign n26387 = ~n25665 & n26386;
  assign n26388 = ~n26098 & n26385;
  assign n26389 = n25673 & ~n35735;
  assign n26390 = n25674 & n26386;
  assign n26391 = ~n25673 & n35735;
  assign n26392 = n25673 & ~n25676;
  assign n26393 = ~n25665 & n26392;
  assign n26394 = ~n26098 & n26393;
  assign n26395 = ~n25673 & ~n35735;
  assign n26396 = ~n26394 & ~n26395;
  assign n26397 = ~n26389 & ~n35736;
  assign n26398 = ~n35734 & ~n35737;
  assign n26399 = ~n26381 & ~n26398;
  assign n26400 = ~n12442 & ~n26399;
  assign n26401 = n12442 & ~n26381;
  assign n26402 = ~n26398 & n26401;
  assign n26403 = ~n35643 & ~n25682;
  assign n26404 = ~n25682 & ~n26098;
  assign n26405 = ~n35643 & n26404;
  assign n26406 = ~n26098 & n26403;
  assign n26407 = n25448 & ~n35738;
  assign n26408 = n25681 & n26404;
  assign n26409 = n25448 & ~n35643;
  assign n26410 = ~n25682 & n26409;
  assign n26411 = ~n26098 & n26410;
  assign n26412 = ~n25448 & ~n35738;
  assign n26413 = ~n26411 & ~n26412;
  assign n26414 = ~n26407 & ~n26408;
  assign n26415 = ~n26402 & ~n35739;
  assign n26416 = ~n26400 & ~n26415;
  assign n26417 = ~n11858 & ~n26416;
  assign n26418 = n11858 & ~n26400;
  assign n26419 = ~n26415 & n26418;
  assign n26420 = n11858 & n26416;
  assign n26421 = ~n25684 & ~n25700;
  assign n26422 = ~n26098 & n26421;
  assign n26423 = ~n35646 & n26422;
  assign n26424 = n35646 & ~n26422;
  assign n26425 = n35646 & ~n25700;
  assign n26426 = ~n25684 & n26425;
  assign n26427 = n35646 & n26422;
  assign n26428 = ~n26098 & n26426;
  assign n26429 = ~n35646 & ~n26422;
  assign n26430 = ~n35741 & ~n26429;
  assign n26431 = ~n26423 & ~n26424;
  assign n26432 = ~n35740 & ~n35742;
  assign n26433 = ~n26417 & ~n26432;
  assign n26434 = ~n11229 & ~n26433;
  assign n26435 = n11229 & ~n26417;
  assign n26436 = ~n26432 & n26435;
  assign n26437 = ~n35647 & ~n25706;
  assign n26438 = ~n25706 & ~n26098;
  assign n26439 = ~n35647 & n26438;
  assign n26440 = ~n26098 & n26437;
  assign n26441 = n25440 & ~n35743;
  assign n26442 = n25705 & n26438;
  assign n26443 = n25440 & ~n35647;
  assign n26444 = ~n25706 & n26443;
  assign n26445 = ~n26098 & n26444;
  assign n26446 = ~n25440 & ~n35743;
  assign n26447 = ~n26445 & ~n26446;
  assign n26448 = ~n26441 & ~n26442;
  assign n26449 = ~n26436 & ~n35744;
  assign n26450 = ~n26434 & ~n26449;
  assign n26451 = ~n10681 & ~n26450;
  assign n26452 = n10681 & ~n26434;
  assign n26453 = ~n26449 & n26452;
  assign n26454 = n10681 & n26450;
  assign n26455 = ~n25708 & ~n25722;
  assign n26456 = ~n25722 & ~n26098;
  assign n26457 = ~n25708 & n26456;
  assign n26458 = ~n26098 & n26455;
  assign n26459 = n35649 & ~n35746;
  assign n26460 = n25720 & n26456;
  assign n26461 = ~n35649 & n35746;
  assign n26462 = n35649 & ~n25722;
  assign n26463 = ~n25708 & n26462;
  assign n26464 = ~n26098 & n26463;
  assign n26465 = ~n35649 & ~n35746;
  assign n26466 = ~n26464 & ~n26465;
  assign n26467 = ~n26459 & ~n35747;
  assign n26468 = ~n35745 & ~n35748;
  assign n26469 = ~n26451 & ~n26468;
  assign n26470 = ~n10086 & ~n26469;
  assign n26471 = n10086 & ~n26451;
  assign n26472 = ~n26468 & n26471;
  assign n26473 = ~n35650 & ~n25728;
  assign n26474 = ~n25728 & ~n26098;
  assign n26475 = ~n35650 & n26474;
  assign n26476 = ~n26098 & n26473;
  assign n26477 = n25432 & ~n35749;
  assign n26478 = n25727 & n26474;
  assign n26479 = n25432 & ~n35650;
  assign n26480 = ~n25728 & n26479;
  assign n26481 = ~n26098 & n26480;
  assign n26482 = ~n25432 & ~n35749;
  assign n26483 = ~n26481 & ~n26482;
  assign n26484 = ~n26477 & ~n26478;
  assign n26485 = ~n26472 & ~n35750;
  assign n26486 = ~n26470 & ~n26485;
  assign n26487 = ~n9565 & ~n26486;
  assign n26488 = ~n25730 & ~n25746;
  assign n26489 = ~n26098 & n26488;
  assign n26490 = ~n35653 & ~n26489;
  assign n26491 = n35653 & ~n25746;
  assign n26492 = ~n25730 & n26491;
  assign n26493 = n35653 & n26489;
  assign n26494 = ~n26098 & n26492;
  assign n26495 = ~n26490 & ~n35751;
  assign n26496 = n9565 & ~n26470;
  assign n26497 = ~n26485 & n26496;
  assign n26498 = n9565 & n26486;
  assign n26499 = ~n26495 & ~n35752;
  assign n26500 = ~n26487 & ~n26499;
  assign n26501 = ~n8998 & ~n26500;
  assign n26502 = n8998 & ~n26487;
  assign n26503 = ~n26499 & n26502;
  assign n26504 = ~n35654 & ~n25752;
  assign n26505 = ~n25752 & ~n26098;
  assign n26506 = ~n35654 & n26505;
  assign n26507 = ~n26098 & n26504;
  assign n26508 = n25424 & ~n35753;
  assign n26509 = n25751 & n26505;
  assign n26510 = n25424 & ~n35654;
  assign n26511 = ~n25752 & n26510;
  assign n26512 = ~n26098 & n26511;
  assign n26513 = ~n25424 & ~n35753;
  assign n26514 = ~n26512 & ~n26513;
  assign n26515 = ~n26508 & ~n26509;
  assign n26516 = ~n26503 & ~n35754;
  assign n26517 = ~n26501 & ~n26516;
  assign n26518 = ~n8506 & ~n26517;
  assign n26519 = n8506 & ~n26501;
  assign n26520 = ~n26516 & n26519;
  assign n26521 = n8506 & n26517;
  assign n26522 = ~n25754 & ~n25757;
  assign n26523 = ~n25757 & ~n26098;
  assign n26524 = ~n25754 & n26523;
  assign n26525 = ~n26098 & n26522;
  assign n26526 = n25416 & ~n35756;
  assign n26527 = n25755 & n26523;
  assign n26528 = n25416 & ~n25757;
  assign n26529 = ~n25754 & n26528;
  assign n26530 = ~n26098 & n26529;
  assign n26531 = ~n25416 & ~n35756;
  assign n26532 = ~n26530 & ~n26531;
  assign n26533 = ~n26526 & ~n26527;
  assign n26534 = ~n35755 & ~n35757;
  assign n26535 = ~n26518 & ~n26534;
  assign n26536 = ~n7975 & ~n26535;
  assign n26537 = n7975 & ~n26518;
  assign n26538 = ~n26534 & n26537;
  assign n26539 = ~n35655 & ~n25763;
  assign n26540 = ~n25763 & ~n26098;
  assign n26541 = ~n35655 & n26540;
  assign n26542 = ~n26098 & n26539;
  assign n26543 = n25408 & ~n35758;
  assign n26544 = n25762 & n26540;
  assign n26545 = n25408 & ~n35655;
  assign n26546 = ~n25763 & n26545;
  assign n26547 = ~n26098 & n26546;
  assign n26548 = ~n25408 & ~n35758;
  assign n26549 = ~n26547 & ~n26548;
  assign n26550 = ~n26543 & ~n26544;
  assign n26551 = ~n26538 & ~n35759;
  assign n26552 = ~n26536 & ~n26551;
  assign n26553 = ~n7512 & ~n26552;
  assign n26554 = ~n25765 & ~n25780;
  assign n26555 = ~n26098 & n26554;
  assign n26556 = ~n35657 & ~n26555;
  assign n26557 = n35657 & ~n25780;
  assign n26558 = ~n25765 & n26557;
  assign n26559 = n35657 & n26555;
  assign n26560 = ~n26098 & n26558;
  assign n26561 = ~n26556 & ~n35760;
  assign n26562 = n7512 & ~n26536;
  assign n26563 = ~n26551 & n26562;
  assign n26564 = n7512 & n26552;
  assign n26565 = ~n26561 & ~n35761;
  assign n26566 = ~n26553 & ~n26565;
  assign n26567 = ~n7015 & ~n26566;
  assign n26568 = n7015 & ~n26553;
  assign n26569 = ~n26565 & n26568;
  assign n26570 = ~n35658 & ~n25786;
  assign n26571 = ~n25786 & ~n26098;
  assign n26572 = ~n35658 & n26571;
  assign n26573 = ~n26098 & n26570;
  assign n26574 = n25400 & ~n35762;
  assign n26575 = n25785 & n26571;
  assign n26576 = n25400 & ~n35658;
  assign n26577 = ~n25786 & n26576;
  assign n26578 = ~n26098 & n26577;
  assign n26579 = ~n25400 & ~n35762;
  assign n26580 = ~n26578 & ~n26579;
  assign n26581 = ~n26574 & ~n26575;
  assign n26582 = ~n26569 & ~n35763;
  assign n26583 = ~n26567 & ~n26582;
  assign n26584 = ~n6579 & ~n26583;
  assign n26585 = n6579 & ~n26567;
  assign n26586 = ~n26582 & n26585;
  assign n26587 = n6579 & n26583;
  assign n26588 = ~n25788 & ~n25791;
  assign n26589 = ~n25791 & ~n26098;
  assign n26590 = ~n25788 & n26589;
  assign n26591 = ~n26098 & n26588;
  assign n26592 = n25392 & ~n35765;
  assign n26593 = n25789 & n26589;
  assign n26594 = n25392 & ~n25791;
  assign n26595 = ~n25788 & n26594;
  assign n26596 = ~n26098 & n26595;
  assign n26597 = ~n25392 & ~n35765;
  assign n26598 = ~n26596 & ~n26597;
  assign n26599 = ~n26592 & ~n26593;
  assign n26600 = ~n35764 & ~n35766;
  assign n26601 = ~n26584 & ~n26600;
  assign n26602 = ~n6117 & ~n26601;
  assign n26603 = n6117 & ~n26584;
  assign n26604 = ~n26600 & n26603;
  assign n26605 = ~n35659 & ~n25797;
  assign n26606 = ~n25797 & ~n26098;
  assign n26607 = ~n35659 & n26606;
  assign n26608 = ~n26098 & n26605;
  assign n26609 = n25384 & ~n35767;
  assign n26610 = n25796 & n26606;
  assign n26611 = n25384 & ~n35659;
  assign n26612 = ~n25797 & n26611;
  assign n26613 = ~n26098 & n26612;
  assign n26614 = ~n25384 & ~n35767;
  assign n26615 = ~n26613 & ~n26614;
  assign n26616 = ~n26609 & ~n26610;
  assign n26617 = ~n26604 & ~n35768;
  assign n26618 = ~n26602 & ~n26617;
  assign n26619 = ~n5708 & ~n26618;
  assign n26620 = ~n25799 & ~n25814;
  assign n26621 = ~n26098 & n26620;
  assign n26622 = ~n35661 & ~n26621;
  assign n26623 = n35661 & ~n25814;
  assign n26624 = ~n25799 & n26623;
  assign n26625 = n35661 & n26621;
  assign n26626 = ~n26098 & n26624;
  assign n26627 = ~n26622 & ~n35769;
  assign n26628 = n5708 & ~n26602;
  assign n26629 = ~n26617 & n26628;
  assign n26630 = n5708 & n26618;
  assign n26631 = ~n26627 & ~n35770;
  assign n26632 = ~n26619 & ~n26631;
  assign n26633 = ~n5278 & ~n26632;
  assign n26634 = n5278 & ~n26619;
  assign n26635 = ~n26631 & n26634;
  assign n26636 = ~n35662 & ~n25820;
  assign n26637 = ~n25820 & ~n26098;
  assign n26638 = ~n35662 & n26637;
  assign n26639 = ~n26098 & n26636;
  assign n26640 = n25376 & ~n35771;
  assign n26641 = n25819 & n26637;
  assign n26642 = n25376 & ~n35662;
  assign n26643 = ~n25820 & n26642;
  assign n26644 = ~n26098 & n26643;
  assign n26645 = ~n25376 & ~n35771;
  assign n26646 = ~n26644 & ~n26645;
  assign n26647 = ~n26640 & ~n26641;
  assign n26648 = ~n26635 & ~n35772;
  assign n26649 = ~n26633 & ~n26648;
  assign n26650 = ~n4903 & ~n26649;
  assign n26651 = n4903 & ~n26633;
  assign n26652 = ~n26648 & n26651;
  assign n26653 = n4903 & n26649;
  assign n26654 = ~n25822 & ~n25825;
  assign n26655 = ~n25825 & ~n26098;
  assign n26656 = ~n25822 & n26655;
  assign n26657 = ~n26098 & n26654;
  assign n26658 = n25368 & ~n35774;
  assign n26659 = n25823 & n26655;
  assign n26660 = n25368 & ~n25825;
  assign n26661 = ~n25822 & n26660;
  assign n26662 = ~n26098 & n26661;
  assign n26663 = ~n25368 & ~n35774;
  assign n26664 = ~n26662 & ~n26663;
  assign n26665 = ~n26658 & ~n26659;
  assign n26666 = ~n35773 & ~n35775;
  assign n26667 = ~n26650 & ~n26666;
  assign n26668 = ~n4508 & ~n26667;
  assign n26669 = n4508 & ~n26650;
  assign n26670 = ~n26666 & n26669;
  assign n26671 = ~n35663 & ~n25831;
  assign n26672 = ~n25831 & ~n26098;
  assign n26673 = ~n35663 & n26672;
  assign n26674 = ~n26098 & n26671;
  assign n26675 = n25360 & ~n35776;
  assign n26676 = n25830 & n26672;
  assign n26677 = n25360 & ~n35663;
  assign n26678 = ~n25831 & n26677;
  assign n26679 = ~n26098 & n26678;
  assign n26680 = ~n25360 & ~n35776;
  assign n26681 = ~n26679 & ~n26680;
  assign n26682 = ~n26675 & ~n26676;
  assign n26683 = ~n26670 & ~n35777;
  assign n26684 = ~n26668 & ~n26683;
  assign n26685 = ~n4155 & ~n26684;
  assign n26686 = ~n25833 & ~n25848;
  assign n26687 = ~n26098 & n26686;
  assign n26688 = ~n35665 & ~n26687;
  assign n26689 = n35665 & ~n25848;
  assign n26690 = ~n25833 & n26689;
  assign n26691 = n35665 & n26687;
  assign n26692 = ~n26098 & n26690;
  assign n26693 = ~n26688 & ~n35778;
  assign n26694 = n4155 & ~n26668;
  assign n26695 = ~n26683 & n26694;
  assign n26696 = n4155 & n26684;
  assign n26697 = ~n26693 & ~n35779;
  assign n26698 = ~n26685 & ~n26697;
  assign n26699 = ~n3788 & ~n26698;
  assign n26700 = n3788 & ~n26685;
  assign n26701 = ~n26697 & n26700;
  assign n26702 = ~n35666 & ~n25854;
  assign n26703 = ~n25854 & ~n26098;
  assign n26704 = ~n35666 & n26703;
  assign n26705 = ~n26098 & n26702;
  assign n26706 = n25352 & ~n35780;
  assign n26707 = n25853 & n26703;
  assign n26708 = n25352 & ~n35666;
  assign n26709 = ~n25854 & n26708;
  assign n26710 = ~n26098 & n26709;
  assign n26711 = ~n25352 & ~n35780;
  assign n26712 = ~n26710 & ~n26711;
  assign n26713 = ~n26706 & ~n26707;
  assign n26714 = ~n26701 & ~n35781;
  assign n26715 = ~n26699 & ~n26714;
  assign n26716 = ~n3473 & ~n26715;
  assign n26717 = n3473 & ~n26699;
  assign n26718 = ~n26714 & n26717;
  assign n26719 = n3473 & n26715;
  assign n26720 = ~n25856 & ~n25859;
  assign n26721 = ~n25859 & ~n26098;
  assign n26722 = ~n25856 & n26721;
  assign n26723 = ~n26098 & n26720;
  assign n26724 = n25344 & ~n35783;
  assign n26725 = n25857 & n26721;
  assign n26726 = n25344 & ~n25859;
  assign n26727 = ~n25856 & n26726;
  assign n26728 = ~n26098 & n26727;
  assign n26729 = ~n25344 & ~n35783;
  assign n26730 = ~n26728 & ~n26729;
  assign n26731 = ~n26724 & ~n26725;
  assign n26732 = ~n35782 & ~n35784;
  assign n26733 = ~n26716 & ~n26732;
  assign n26734 = ~n3140 & ~n26733;
  assign n26735 = n3140 & ~n26716;
  assign n26736 = ~n26732 & n26735;
  assign n26737 = ~n35667 & ~n25865;
  assign n26738 = ~n25865 & ~n26098;
  assign n26739 = ~n35667 & n26738;
  assign n26740 = ~n26098 & n26737;
  assign n26741 = n25336 & ~n35785;
  assign n26742 = n25864 & n26738;
  assign n26743 = n25336 & ~n35667;
  assign n26744 = ~n25865 & n26743;
  assign n26745 = ~n26098 & n26744;
  assign n26746 = ~n25336 & ~n35785;
  assign n26747 = ~n26745 & ~n26746;
  assign n26748 = ~n26741 & ~n26742;
  assign n26749 = ~n26736 & ~n35786;
  assign n26750 = ~n26734 & ~n26749;
  assign n26751 = ~n2855 & ~n26750;
  assign n26752 = ~n25867 & ~n25882;
  assign n26753 = ~n26098 & n26752;
  assign n26754 = ~n35669 & ~n26753;
  assign n26755 = n35669 & ~n25882;
  assign n26756 = ~n25867 & n26755;
  assign n26757 = n35669 & n26753;
  assign n26758 = ~n26098 & n26756;
  assign n26759 = ~n26754 & ~n35787;
  assign n26760 = n2855 & ~n26734;
  assign n26761 = ~n26749 & n26760;
  assign n26762 = n2855 & n26750;
  assign n26763 = ~n26759 & ~n35788;
  assign n26764 = ~n26751 & ~n26763;
  assign n26765 = ~n2556 & ~n26764;
  assign n26766 = n2556 & ~n26751;
  assign n26767 = ~n26763 & n26766;
  assign n26768 = ~n35670 & ~n25888;
  assign n26769 = ~n25888 & ~n26098;
  assign n26770 = ~n35670 & n26769;
  assign n26771 = ~n26098 & n26768;
  assign n26772 = n25328 & ~n35789;
  assign n26773 = n25887 & n26769;
  assign n26774 = n25328 & ~n35670;
  assign n26775 = ~n25888 & n26774;
  assign n26776 = ~n26098 & n26775;
  assign n26777 = ~n25328 & ~n35789;
  assign n26778 = ~n26776 & ~n26777;
  assign n26779 = ~n26772 & ~n26773;
  assign n26780 = ~n26767 & ~n35790;
  assign n26781 = ~n26765 & ~n26780;
  assign n26782 = ~n2301 & ~n26781;
  assign n26783 = n2301 & ~n26765;
  assign n26784 = ~n26780 & n26783;
  assign n26785 = n2301 & n26781;
  assign n26786 = ~n25890 & ~n25893;
  assign n26787 = ~n25893 & ~n26098;
  assign n26788 = ~n25890 & n26787;
  assign n26789 = ~n26098 & n26786;
  assign n26790 = n25320 & ~n35792;
  assign n26791 = n25891 & n26787;
  assign n26792 = n25320 & ~n25893;
  assign n26793 = ~n25890 & n26792;
  assign n26794 = ~n26098 & n26793;
  assign n26795 = ~n25320 & ~n35792;
  assign n26796 = ~n26794 & ~n26795;
  assign n26797 = ~n26790 & ~n26791;
  assign n26798 = ~n35791 & ~n35793;
  assign n26799 = ~n26782 & ~n26798;
  assign n26800 = ~n2038 & ~n26799;
  assign n26801 = n2038 & ~n26782;
  assign n26802 = ~n26798 & n26801;
  assign n26803 = ~n35671 & ~n25899;
  assign n26804 = ~n25899 & ~n26098;
  assign n26805 = ~n35671 & n26804;
  assign n26806 = ~n26098 & n26803;
  assign n26807 = n25312 & ~n35794;
  assign n26808 = n25898 & n26804;
  assign n26809 = n25312 & ~n35671;
  assign n26810 = ~n25899 & n26809;
  assign n26811 = ~n26098 & n26810;
  assign n26812 = ~n25312 & ~n35794;
  assign n26813 = ~n26811 & ~n26812;
  assign n26814 = ~n26807 & ~n26808;
  assign n26815 = ~n26802 & ~n35795;
  assign n26816 = ~n26800 & ~n26815;
  assign n26817 = ~n1812 & ~n26816;
  assign n26818 = ~n25901 & ~n25916;
  assign n26819 = ~n26098 & n26818;
  assign n26820 = ~n35673 & ~n26819;
  assign n26821 = n35673 & ~n25916;
  assign n26822 = ~n25901 & n26821;
  assign n26823 = n35673 & n26819;
  assign n26824 = ~n26098 & n26822;
  assign n26825 = ~n26820 & ~n35796;
  assign n26826 = n1812 & ~n26800;
  assign n26827 = ~n26815 & n26826;
  assign n26828 = n1812 & n26816;
  assign n26829 = ~n26825 & ~n35797;
  assign n26830 = ~n26817 & ~n26829;
  assign n26831 = ~n1582 & ~n26830;
  assign n26832 = n1582 & ~n26817;
  assign n26833 = ~n26829 & n26832;
  assign n26834 = ~n35674 & ~n25922;
  assign n26835 = ~n25922 & ~n26098;
  assign n26836 = ~n35674 & n26835;
  assign n26837 = ~n26098 & n26834;
  assign n26838 = n25304 & ~n35798;
  assign n26839 = n25921 & n26835;
  assign n26840 = n25304 & ~n35674;
  assign n26841 = ~n25922 & n26840;
  assign n26842 = ~n26098 & n26841;
  assign n26843 = ~n25304 & ~n35798;
  assign n26844 = ~n26842 & ~n26843;
  assign n26845 = ~n26838 & ~n26839;
  assign n26846 = ~n26833 & ~n35799;
  assign n26847 = ~n26831 & ~n26846;
  assign n26848 = ~n1388 & ~n26847;
  assign n26849 = n1388 & ~n26831;
  assign n26850 = ~n26846 & n26849;
  assign n26851 = n1388 & n26847;
  assign n26852 = ~n25924 & ~n25927;
  assign n26853 = ~n25927 & ~n26098;
  assign n26854 = ~n25924 & n26853;
  assign n26855 = ~n26098 & n26852;
  assign n26856 = n25296 & ~n35801;
  assign n26857 = n25925 & n26853;
  assign n26858 = n25296 & ~n25927;
  assign n26859 = ~n25924 & n26858;
  assign n26860 = ~n26098 & n26859;
  assign n26861 = ~n25296 & ~n35801;
  assign n26862 = ~n26860 & ~n26861;
  assign n26863 = ~n26856 & ~n26857;
  assign n26864 = ~n35800 & ~n35802;
  assign n26865 = ~n26848 & ~n26864;
  assign n26866 = ~n1192 & ~n26865;
  assign n26867 = n1192 & ~n26848;
  assign n26868 = ~n26864 & n26867;
  assign n26869 = ~n35675 & ~n25933;
  assign n26870 = ~n25933 & ~n26098;
  assign n26871 = ~n35675 & n26870;
  assign n26872 = ~n26098 & n26869;
  assign n26873 = n25288 & ~n35803;
  assign n26874 = n25932 & n26870;
  assign n26875 = n25288 & ~n35675;
  assign n26876 = ~n25933 & n26875;
  assign n26877 = ~n26098 & n26876;
  assign n26878 = ~n25288 & ~n35803;
  assign n26879 = ~n26877 & ~n26878;
  assign n26880 = ~n26873 & ~n26874;
  assign n26881 = ~n26868 & ~n35804;
  assign n26882 = ~n26866 & ~n26881;
  assign n26883 = ~n1028 & ~n26882;
  assign n26884 = ~n25935 & ~n25950;
  assign n26885 = ~n26098 & n26884;
  assign n26886 = ~n35677 & ~n26885;
  assign n26887 = n35677 & ~n25950;
  assign n26888 = ~n25935 & n26887;
  assign n26889 = n35677 & n26885;
  assign n26890 = ~n26098 & n26888;
  assign n26891 = ~n26886 & ~n35805;
  assign n26892 = n1028 & ~n26866;
  assign n26893 = ~n26881 & n26892;
  assign n26894 = n1028 & n26882;
  assign n26895 = ~n26891 & ~n35806;
  assign n26896 = ~n26883 & ~n26895;
  assign n26897 = ~n866 & ~n26896;
  assign n26898 = n866 & ~n26883;
  assign n26899 = ~n26895 & n26898;
  assign n26900 = ~n35678 & ~n25956;
  assign n26901 = ~n25956 & ~n26098;
  assign n26902 = ~n35678 & n26901;
  assign n26903 = ~n26098 & n26900;
  assign n26904 = n25280 & ~n35807;
  assign n26905 = n25955 & n26901;
  assign n26906 = n25280 & ~n35678;
  assign n26907 = ~n25956 & n26906;
  assign n26908 = ~n26098 & n26907;
  assign n26909 = ~n25280 & ~n35807;
  assign n26910 = ~n26908 & ~n26909;
  assign n26911 = ~n26904 & ~n26905;
  assign n26912 = ~n26899 & ~n35808;
  assign n26913 = ~n26897 & ~n26912;
  assign n26914 = ~n730 & ~n26913;
  assign n26915 = n730 & ~n26897;
  assign n26916 = ~n26912 & n26915;
  assign n26917 = n730 & n26913;
  assign n26918 = ~n25958 & ~n25961;
  assign n26919 = ~n25961 & ~n26098;
  assign n26920 = ~n25958 & n26919;
  assign n26921 = ~n26098 & n26918;
  assign n26922 = n25272 & ~n35810;
  assign n26923 = n25959 & n26919;
  assign n26924 = n25272 & ~n25961;
  assign n26925 = ~n25958 & n26924;
  assign n26926 = ~n26098 & n26925;
  assign n26927 = ~n25272 & ~n35810;
  assign n26928 = ~n26926 & ~n26927;
  assign n26929 = ~n26922 & ~n26923;
  assign n26930 = ~n35809 & ~n35811;
  assign n26931 = ~n26914 & ~n26930;
  assign n26932 = ~n602 & ~n26931;
  assign n26933 = n602 & ~n26914;
  assign n26934 = ~n26930 & n26933;
  assign n26935 = ~n35679 & ~n25977;
  assign n26936 = ~n26098 & n26935;
  assign n26937 = ~n35680 & n26936;
  assign n26938 = n35680 & ~n26936;
  assign n26939 = ~n35679 & n35680;
  assign n26940 = ~n25977 & n26939;
  assign n26941 = ~n26098 & n26940;
  assign n26942 = ~n35680 & ~n26936;
  assign n26943 = ~n26941 & ~n26942;
  assign n26944 = ~n26937 & ~n26938;
  assign n26945 = ~n26934 & ~n35812;
  assign n26946 = ~n26932 & ~n26945;
  assign n26947 = ~n497 & ~n26946;
  assign n26948 = n497 & ~n26932;
  assign n26949 = ~n26945 & n26948;
  assign n26950 = n497 & n26946;
  assign n26951 = ~n25979 & ~n25981;
  assign n26952 = ~n26098 & n26951;
  assign n26953 = ~n35681 & ~n26952;
  assign n26954 = ~n25979 & n35681;
  assign n26955 = ~n25981 & n26954;
  assign n26956 = n35681 & n26952;
  assign n26957 = ~n26098 & n26955;
  assign n26958 = ~n26953 & ~n35814;
  assign n26959 = ~n35813 & ~n26958;
  assign n26960 = ~n26947 & ~n26959;
  assign n26961 = ~n403 & ~n26960;
  assign n26962 = n403 & ~n26947;
  assign n26963 = ~n26959 & n26962;
  assign n26964 = ~n35696 & ~n26963;
  assign n26965 = ~n26961 & ~n26964;
  assign n26966 = ~n330 & ~n26965;
  assign n26967 = ~n26000 & ~n26002;
  assign n26968 = ~n26098 & n26967;
  assign n26969 = ~n35684 & ~n26968;
  assign n26970 = ~n26000 & n35684;
  assign n26971 = ~n26002 & n26970;
  assign n26972 = n35684 & n26968;
  assign n26973 = ~n26098 & n26971;
  assign n26974 = ~n26969 & ~n35815;
  assign n26975 = n330 & ~n26961;
  assign n26976 = ~n26964 & n26975;
  assign n26977 = n330 & n26965;
  assign n26978 = ~n26974 & ~n35816;
  assign n26979 = ~n26966 & ~n26978;
  assign n26980 = ~n271 & ~n26979;
  assign n26981 = n271 & ~n26966;
  assign n26982 = ~n26978 & n26981;
  assign n26983 = ~n26017 & ~n35686;
  assign n26984 = ~n26017 & ~n26098;
  assign n26985 = ~n35686 & n26984;
  assign n26986 = ~n26098 & n26983;
  assign n26987 = n26025 & ~n35817;
  assign n26988 = n26029 & n26984;
  assign n26989 = n26025 & ~n35686;
  assign n26990 = ~n26017 & n26989;
  assign n26991 = ~n26098 & n26990;
  assign n26992 = ~n26025 & ~n35817;
  assign n26993 = ~n26991 & ~n26992;
  assign n26994 = ~n26987 & ~n26988;
  assign n26995 = ~n26982 & ~n35818;
  assign n26996 = ~n26980 & ~n26995;
  assign n26997 = ~n217 & ~n26996;
  assign n26998 = ~n26031 & ~n26033;
  assign n26999 = ~n26098 & n26998;
  assign n27000 = ~n35688 & ~n26999;
  assign n27001 = ~n26031 & n35688;
  assign n27002 = ~n26033 & n27001;
  assign n27003 = n35688 & n26999;
  assign n27004 = ~n26098 & n27002;
  assign n27005 = ~n27000 & ~n35819;
  assign n27006 = n217 & ~n26980;
  assign n27007 = ~n26995 & n27006;
  assign n27008 = n217 & n26996;
  assign n27009 = ~n27005 & ~n35820;
  assign n27010 = ~n26997 & ~n27009;
  assign n27011 = ~n198 & ~n27010;
  assign n27012 = n198 & ~n26997;
  assign n27013 = ~n27009 & n27012;
  assign n27014 = ~n26048 & ~n35690;
  assign n27015 = ~n26048 & ~n26098;
  assign n27016 = ~n35690 & n27015;
  assign n27017 = ~n26098 & n27014;
  assign n27018 = n26056 & ~n35821;
  assign n27019 = n26060 & n27015;
  assign n27020 = n26056 & ~n35690;
  assign n27021 = ~n26048 & n27020;
  assign n27022 = ~n26098 & n27021;
  assign n27023 = ~n26056 & ~n35821;
  assign n27024 = ~n27022 & ~n27023;
  assign n27025 = ~n27018 & ~n27019;
  assign n27026 = ~n27013 & ~n35822;
  assign n27027 = ~n27011 & ~n27026;
  assign n27028 = ~n26062 & ~n26072;
  assign n27029 = ~n26062 & ~n26098;
  assign n27030 = ~n26072 & n27029;
  assign n27031 = ~n26098 & n27028;
  assign n27032 = n26070 & ~n35823;
  assign n27033 = n26073 & n27029;
  assign n27034 = ~n26062 & n26070;
  assign n27035 = ~n26072 & n27034;
  assign n27036 = ~n26098 & n27035;
  assign n27037 = ~n26070 & ~n35823;
  assign n27038 = ~n27036 & ~n27037;
  assign n27039 = ~n27032 & ~n27033;
  assign n27040 = ~n26074 & ~n26082;
  assign n27041 = ~n26082 & ~n26098;
  assign n27042 = ~n26074 & n27041;
  assign n27043 = ~n26098 & n27040;
  assign n27044 = ~n35694 & ~n35825;
  assign n27045 = ~n35824 & n27044;
  assign n27046 = ~n27027 & n27045;
  assign n27047 = n193 & ~n27046;
  assign n27048 = ~n27011 & n35824;
  assign n27049 = ~n27026 & n27048;
  assign n27050 = n27027 & n35824;
  assign n27051 = n26074 & ~n27041;
  assign n27052 = ~n193 & ~n27040;
  assign n27053 = ~n27051 & n27052;
  assign n27054 = ~n35826 & ~n27053;
  assign n27055 = ~n27047 & n27054;
  assign n27056 = ~n26961 & ~n26963;
  assign n27057 = ~n27055 & n27056;
  assign n27058 = ~n35696 & ~n27057;
  assign n27059 = n35696 & ~n26963;
  assign n27060 = ~n26961 & n27059;
  assign n27061 = n35696 & n27057;
  assign n27062 = ~n27055 & n27060;
  assign n27063 = ~n27058 & ~n35827;
  assign n27064 = ~n26932 & ~n26934;
  assign n27065 = ~n27055 & n27064;
  assign n27066 = ~n35812 & ~n27065;
  assign n27067 = ~n26934 & n35812;
  assign n27068 = ~n26932 & n27067;
  assign n27069 = n35812 & n27065;
  assign n27070 = ~n27055 & n27068;
  assign n27071 = ~n27066 & ~n35828;
  assign n27072 = ~n26914 & ~n35809;
  assign n27073 = ~n27055 & n27072;
  assign n27074 = ~n35811 & ~n27073;
  assign n27075 = ~n26914 & n35811;
  assign n27076 = ~n35809 & n27075;
  assign n27077 = n35811 & n27073;
  assign n27078 = ~n27055 & n27076;
  assign n27079 = ~n27074 & ~n35829;
  assign n27080 = ~n26897 & ~n26899;
  assign n27081 = ~n27055 & n27080;
  assign n27082 = ~n35808 & ~n27081;
  assign n27083 = ~n26899 & n35808;
  assign n27084 = ~n26897 & n27083;
  assign n27085 = n35808 & n27081;
  assign n27086 = ~n27055 & n27084;
  assign n27087 = ~n27082 & ~n35830;
  assign n27088 = ~n26866 & ~n26868;
  assign n27089 = ~n27055 & n27088;
  assign n27090 = ~n35804 & ~n27089;
  assign n27091 = ~n26868 & n35804;
  assign n27092 = ~n26866 & n27091;
  assign n27093 = n35804 & n27089;
  assign n27094 = ~n27055 & n27092;
  assign n27095 = ~n27090 & ~n35831;
  assign n27096 = ~n26848 & ~n35800;
  assign n27097 = ~n27055 & n27096;
  assign n27098 = ~n35802 & ~n27097;
  assign n27099 = ~n26848 & n35802;
  assign n27100 = ~n35800 & n27099;
  assign n27101 = n35802 & n27097;
  assign n27102 = ~n27055 & n27100;
  assign n27103 = ~n27098 & ~n35832;
  assign n27104 = ~n26831 & ~n26833;
  assign n27105 = ~n27055 & n27104;
  assign n27106 = ~n35799 & ~n27105;
  assign n27107 = ~n26833 & n35799;
  assign n27108 = ~n26831 & n27107;
  assign n27109 = n35799 & n27105;
  assign n27110 = ~n27055 & n27108;
  assign n27111 = ~n27106 & ~n35833;
  assign n27112 = ~n26800 & ~n26802;
  assign n27113 = ~n27055 & n27112;
  assign n27114 = ~n35795 & ~n27113;
  assign n27115 = ~n26802 & n35795;
  assign n27116 = ~n26800 & n27115;
  assign n27117 = n35795 & n27113;
  assign n27118 = ~n27055 & n27116;
  assign n27119 = ~n27114 & ~n35834;
  assign n27120 = ~n26782 & ~n35791;
  assign n27121 = ~n27055 & n27120;
  assign n27122 = ~n35793 & ~n27121;
  assign n27123 = ~n26782 & n35793;
  assign n27124 = ~n35791 & n27123;
  assign n27125 = n35793 & n27121;
  assign n27126 = ~n27055 & n27124;
  assign n27127 = ~n27122 & ~n35835;
  assign n27128 = ~n26765 & ~n26767;
  assign n27129 = ~n27055 & n27128;
  assign n27130 = ~n35790 & ~n27129;
  assign n27131 = ~n26767 & n35790;
  assign n27132 = ~n26765 & n27131;
  assign n27133 = n35790 & n27129;
  assign n27134 = ~n27055 & n27132;
  assign n27135 = ~n27130 & ~n35836;
  assign n27136 = ~n26734 & ~n26736;
  assign n27137 = ~n27055 & n27136;
  assign n27138 = ~n35786 & ~n27137;
  assign n27139 = ~n26736 & n35786;
  assign n27140 = ~n26734 & n27139;
  assign n27141 = n35786 & n27137;
  assign n27142 = ~n27055 & n27140;
  assign n27143 = ~n27138 & ~n35837;
  assign n27144 = ~n26716 & ~n35782;
  assign n27145 = ~n27055 & n27144;
  assign n27146 = ~n35784 & ~n27145;
  assign n27147 = ~n26716 & n35784;
  assign n27148 = ~n35782 & n27147;
  assign n27149 = n35784 & n27145;
  assign n27150 = ~n27055 & n27148;
  assign n27151 = ~n27146 & ~n35838;
  assign n27152 = ~n26699 & ~n26701;
  assign n27153 = ~n27055 & n27152;
  assign n27154 = ~n35781 & ~n27153;
  assign n27155 = ~n26701 & n35781;
  assign n27156 = ~n26699 & n27155;
  assign n27157 = n35781 & n27153;
  assign n27158 = ~n27055 & n27156;
  assign n27159 = ~n27154 & ~n35839;
  assign n27160 = ~n26668 & ~n26670;
  assign n27161 = ~n27055 & n27160;
  assign n27162 = ~n35777 & ~n27161;
  assign n27163 = ~n26670 & n35777;
  assign n27164 = ~n26668 & n27163;
  assign n27165 = n35777 & n27161;
  assign n27166 = ~n27055 & n27164;
  assign n27167 = ~n27162 & ~n35840;
  assign n27168 = ~n26650 & ~n35773;
  assign n27169 = ~n27055 & n27168;
  assign n27170 = ~n35775 & ~n27169;
  assign n27171 = ~n26650 & n35775;
  assign n27172 = ~n35773 & n27171;
  assign n27173 = n35775 & n27169;
  assign n27174 = ~n27055 & n27172;
  assign n27175 = ~n27170 & ~n35841;
  assign n27176 = ~n26633 & ~n26635;
  assign n27177 = ~n27055 & n27176;
  assign n27178 = ~n35772 & ~n27177;
  assign n27179 = ~n26635 & n35772;
  assign n27180 = ~n26633 & n27179;
  assign n27181 = n35772 & n27177;
  assign n27182 = ~n27055 & n27180;
  assign n27183 = ~n27178 & ~n35842;
  assign n27184 = ~n26602 & ~n26604;
  assign n27185 = ~n27055 & n27184;
  assign n27186 = ~n35768 & ~n27185;
  assign n27187 = ~n26604 & n35768;
  assign n27188 = ~n26602 & n27187;
  assign n27189 = n35768 & n27185;
  assign n27190 = ~n27055 & n27188;
  assign n27191 = ~n27186 & ~n35843;
  assign n27192 = ~n26584 & ~n35764;
  assign n27193 = ~n27055 & n27192;
  assign n27194 = ~n35766 & ~n27193;
  assign n27195 = ~n26584 & n35766;
  assign n27196 = ~n35764 & n27195;
  assign n27197 = n35766 & n27193;
  assign n27198 = ~n27055 & n27196;
  assign n27199 = ~n27194 & ~n35844;
  assign n27200 = ~n26567 & ~n26569;
  assign n27201 = ~n27055 & n27200;
  assign n27202 = ~n35763 & ~n27201;
  assign n27203 = ~n26569 & n35763;
  assign n27204 = ~n26567 & n27203;
  assign n27205 = n35763 & n27201;
  assign n27206 = ~n27055 & n27204;
  assign n27207 = ~n27202 & ~n35845;
  assign n27208 = ~n26536 & ~n26538;
  assign n27209 = ~n27055 & n27208;
  assign n27210 = ~n35759 & ~n27209;
  assign n27211 = ~n26538 & n35759;
  assign n27212 = ~n26536 & n27211;
  assign n27213 = n35759 & n27209;
  assign n27214 = ~n27055 & n27212;
  assign n27215 = ~n27210 & ~n35846;
  assign n27216 = ~n26518 & ~n35755;
  assign n27217 = ~n27055 & n27216;
  assign n27218 = ~n35757 & ~n27217;
  assign n27219 = ~n26518 & n35757;
  assign n27220 = ~n35755 & n27219;
  assign n27221 = n35757 & n27217;
  assign n27222 = ~n27055 & n27220;
  assign n27223 = ~n27218 & ~n35847;
  assign n27224 = ~n26501 & ~n26503;
  assign n27225 = ~n27055 & n27224;
  assign n27226 = ~n35754 & ~n27225;
  assign n27227 = ~n26503 & n35754;
  assign n27228 = ~n26501 & n27227;
  assign n27229 = n35754 & n27225;
  assign n27230 = ~n27055 & n27228;
  assign n27231 = ~n27226 & ~n35848;
  assign n27232 = ~n26470 & ~n26472;
  assign n27233 = ~n27055 & n27232;
  assign n27234 = ~n35750 & ~n27233;
  assign n27235 = ~n26472 & n35750;
  assign n27236 = ~n26470 & n27235;
  assign n27237 = n35750 & n27233;
  assign n27238 = ~n27055 & n27236;
  assign n27239 = ~n27234 & ~n35849;
  assign n27240 = ~n26451 & ~n35745;
  assign n27241 = ~n27055 & n27240;
  assign n27242 = ~n35748 & ~n27241;
  assign n27243 = ~n26451 & n35748;
  assign n27244 = ~n35745 & n27243;
  assign n27245 = n35748 & n27241;
  assign n27246 = ~n27055 & n27244;
  assign n27247 = ~n27242 & ~n35850;
  assign n27248 = ~n26434 & ~n26436;
  assign n27249 = ~n27055 & n27248;
  assign n27250 = ~n35744 & ~n27249;
  assign n27251 = ~n26436 & n35744;
  assign n27252 = ~n26434 & n27251;
  assign n27253 = n35744 & n27249;
  assign n27254 = ~n27055 & n27252;
  assign n27255 = ~n27250 & ~n35851;
  assign n27256 = ~n26400 & ~n26402;
  assign n27257 = ~n27055 & n27256;
  assign n27258 = ~n35739 & ~n27257;
  assign n27259 = ~n26402 & n35739;
  assign n27260 = ~n26400 & n27259;
  assign n27261 = n35739 & n27257;
  assign n27262 = ~n27055 & n27260;
  assign n27263 = ~n27258 & ~n35852;
  assign n27264 = ~n26364 & ~n26366;
  assign n27265 = ~n27055 & n27264;
  assign n27266 = ~n35733 & ~n27265;
  assign n27267 = ~n26366 & n35733;
  assign n27268 = ~n26364 & n27267;
  assign n27269 = n35733 & n27265;
  assign n27270 = ~n27055 & n27268;
  assign n27271 = ~n27266 & ~n35853;
  assign n27272 = ~n26333 & ~n26335;
  assign n27273 = ~n27055 & n27272;
  assign n27274 = ~n35729 & ~n27273;
  assign n27275 = ~n26335 & n35729;
  assign n27276 = ~n26333 & n27275;
  assign n27277 = n35729 & n27273;
  assign n27278 = ~n27055 & n27276;
  assign n27279 = ~n27274 & ~n35854;
  assign n27280 = ~n26297 & ~n26299;
  assign n27281 = ~n27055 & n27280;
  assign n27282 = ~n35723 & ~n27281;
  assign n27283 = ~n26299 & n35723;
  assign n27284 = ~n26297 & n27283;
  assign n27285 = n35723 & n27281;
  assign n27286 = ~n27055 & n27284;
  assign n27287 = ~n27282 & ~n35855;
  assign n27288 = ~n26263 & ~n26265;
  assign n27289 = ~n27055 & n27288;
  assign n27290 = ~n35718 & ~n27289;
  assign n27291 = ~n26265 & n35718;
  assign n27292 = ~n26263 & n27291;
  assign n27293 = n35718 & n27289;
  assign n27294 = ~n27055 & n27292;
  assign n27295 = ~n27290 & ~n35856;
  assign n27296 = ~n26229 & ~n26231;
  assign n27297 = ~n27055 & n27296;
  assign n27298 = ~n35713 & ~n27297;
  assign n27299 = ~n26231 & n35713;
  assign n27300 = ~n26229 & n27299;
  assign n27301 = n35713 & n27297;
  assign n27302 = ~n27055 & n27300;
  assign n27303 = ~n27298 & ~n35857;
  assign n27304 = ~n26196 & ~n26198;
  assign n27305 = ~n27055 & n27304;
  assign n27306 = ~n35709 & ~n27305;
  assign n27307 = ~n26198 & n35709;
  assign n27308 = ~n26196 & n27307;
  assign n27309 = n35709 & n27305;
  assign n27310 = ~n27055 & n27308;
  assign n27311 = ~n27306 & ~n35858;
  assign n27312 = ~n26162 & ~n26164;
  assign n27313 = ~n27055 & n27312;
  assign n27314 = ~n35704 & ~n27313;
  assign n27315 = ~n26164 & n35704;
  assign n27316 = ~n26162 & n27315;
  assign n27317 = n35704 & n27313;
  assign n27318 = ~n27055 & n27316;
  assign n27319 = ~n27314 & ~n35859;
  assign n27320 = ~n26135 & ~n26137;
  assign n27321 = ~n27055 & n27320;
  assign n27322 = ~n26146 & ~n27321;
  assign n27323 = ~n26137 & n26146;
  assign n27324 = ~n26135 & n27323;
  assign n27325 = n26146 & n27321;
  assign n27326 = ~n27055 & n27324;
  assign n27327 = ~n27322 & ~n35860;
  assign n27328 = ~pi10  & ~n27055;
  assign n27329 = ~pi11  & n27328;
  assign n27330 = n26112 & ~n27055;
  assign n27331 = ~n26098 & ~n27053;
  assign n27332 = ~n35826 & n27331;
  assign n27333 = ~n26098 & n27055;
  assign n27334 = ~n27047 & n27332;
  assign n27335 = ~n35861 & ~n35862;
  assign n27336 = pi12  & ~n27335;
  assign n27337 = ~pi12  & ~n35862;
  assign n27338 = ~pi12  & n27335;
  assign n27339 = ~n35861 & n27337;
  assign n27340 = ~n27336 & ~n35863;
  assign n27341 = pi10  & ~n27055;
  assign n27342 = ~pi8  & ~pi9 ;
  assign n27343 = ~pi10  & n27342;
  assign n27344 = ~n35587 & ~n35698;
  assign n27345 = ~n25235 & n27344;
  assign n27346 = ~n25254 & n27345;
  assign n27347 = ~n35589 & n27346;
  assign n27348 = n25240 & n25256;
  assign n27349 = ~n25248 & n27347;
  assign n27350 = ~n27343 & ~n35864;
  assign n27351 = ~n26096 & n27350;
  assign n27352 = ~n35694 & n27351;
  assign n27353 = ~n26090 & n27352;
  assign n27354 = ~pi10  & ~n27342;
  assign n27355 = pi10  & n27055;
  assign n27356 = ~n27354 & ~n27355;
  assign n27357 = ~n27341 & ~n27343;
  assign n27358 = n26098 & ~n35865;
  assign n27359 = ~n27341 & n27353;
  assign n27360 = pi11  & ~n27328;
  assign n27361 = ~n35861 & ~n27360;
  assign n27362 = ~n35866 & n27361;
  assign n27363 = ~n26098 & n35865;
  assign n27364 = n25256 & ~n27363;
  assign n27365 = ~n27362 & ~n27363;
  assign n27366 = n25256 & n27365;
  assign n27367 = ~n27362 & n27364;
  assign n27368 = ~n27340 & ~n35867;
  assign n27369 = ~n25256 & ~n27365;
  assign n27370 = n24331 & ~n27369;
  assign n27371 = ~n27368 & n27370;
  assign n27372 = ~n26115 & ~n35699;
  assign n27373 = ~n27055 & n27372;
  assign n27374 = n26120 & ~n27373;
  assign n27375 = ~n26120 & n27372;
  assign n27376 = ~n26120 & n27373;
  assign n27377 = ~n27055 & n27375;
  assign n27378 = ~n27374 & ~n35868;
  assign n27379 = ~n27371 & ~n27378;
  assign n27380 = ~n27368 & ~n27369;
  assign n27381 = ~n24331 & ~n27380;
  assign n27382 = n23517 & ~n27381;
  assign n27383 = ~n27379 & ~n27381;
  assign n27384 = n23517 & n27383;
  assign n27385 = ~n27379 & n27382;
  assign n27386 = ~n27327 & ~n35869;
  assign n27387 = ~n23517 & ~n27383;
  assign n27388 = n22625 & ~n27387;
  assign n27389 = ~n27386 & n27388;
  assign n27390 = ~n26149 & ~n35701;
  assign n27391 = ~n27055 & n27390;
  assign n27392 = n26159 & ~n27391;
  assign n27393 = ~n26159 & n27391;
  assign n27394 = ~n26149 & n26159;
  assign n27395 = ~n35701 & n27394;
  assign n27396 = n26159 & n27391;
  assign n27397 = ~n27055 & n27395;
  assign n27398 = ~n26159 & ~n27391;
  assign n27399 = ~n35870 & ~n27398;
  assign n27400 = ~n27392 & ~n27393;
  assign n27401 = ~n27389 & ~n35871;
  assign n27402 = ~n27386 & ~n27387;
  assign n27403 = ~n22625 & ~n27402;
  assign n27404 = n21842 & ~n27403;
  assign n27405 = ~n27401 & ~n27403;
  assign n27406 = n21842 & n27405;
  assign n27407 = ~n27401 & n27404;
  assign n27408 = ~n27319 & ~n35872;
  assign n27409 = ~n21842 & ~n27405;
  assign n27410 = n20986 & ~n27409;
  assign n27411 = ~n27408 & n27410;
  assign n27412 = ~n26179 & ~n35705;
  assign n27413 = ~n27055 & n27412;
  assign n27414 = ~n35707 & n27413;
  assign n27415 = n35707 & ~n27413;
  assign n27416 = ~n26179 & n35707;
  assign n27417 = ~n35705 & n27416;
  assign n27418 = ~n27055 & n27417;
  assign n27419 = ~n35707 & ~n27413;
  assign n27420 = ~n27418 & ~n27419;
  assign n27421 = ~n27414 & ~n27415;
  assign n27422 = ~n27411 & ~n35873;
  assign n27423 = ~n27408 & ~n27409;
  assign n27424 = ~n20986 & ~n27423;
  assign n27425 = n20229 & ~n27424;
  assign n27426 = ~n27422 & ~n27424;
  assign n27427 = n20229 & n27426;
  assign n27428 = ~n27422 & n27425;
  assign n27429 = ~n27311 & ~n35874;
  assign n27430 = ~n20229 & ~n27426;
  assign n27431 = n19401 & ~n27430;
  assign n27432 = ~n27429 & n27431;
  assign n27433 = ~n26213 & ~n35710;
  assign n27434 = ~n27055 & n27433;
  assign n27435 = ~n35711 & ~n27434;
  assign n27436 = ~n26213 & n35711;
  assign n27437 = ~n35710 & n27436;
  assign n27438 = n35711 & n27434;
  assign n27439 = ~n27055 & n27437;
  assign n27440 = n35711 & ~n27434;
  assign n27441 = ~n35711 & n27434;
  assign n27442 = ~n27440 & ~n27441;
  assign n27443 = ~n27435 & ~n35875;
  assign n27444 = ~n27432 & n35876;
  assign n27445 = ~n27429 & ~n27430;
  assign n27446 = ~n19401 & ~n27445;
  assign n27447 = n18676 & ~n27446;
  assign n27448 = ~n27444 & ~n27446;
  assign n27449 = n18676 & n27448;
  assign n27450 = ~n27444 & n27447;
  assign n27451 = ~n27303 & ~n35877;
  assign n27452 = ~n18676 & ~n27448;
  assign n27453 = n17885 & ~n27452;
  assign n27454 = ~n27451 & n27453;
  assign n27455 = ~n26246 & ~n35714;
  assign n27456 = ~n27055 & n27455;
  assign n27457 = n35716 & ~n27456;
  assign n27458 = ~n26246 & ~n35716;
  assign n27459 = ~n35714 & n27458;
  assign n27460 = ~n35716 & n27456;
  assign n27461 = ~n27055 & n27459;
  assign n27462 = n35716 & n27456;
  assign n27463 = ~n35716 & ~n27456;
  assign n27464 = ~n27462 & ~n27463;
  assign n27465 = ~n27457 & ~n35878;
  assign n27466 = ~n27454 & n35879;
  assign n27467 = ~n27451 & ~n27452;
  assign n27468 = ~n17885 & ~n27467;
  assign n27469 = n17187 & ~n27468;
  assign n27470 = ~n27466 & ~n27468;
  assign n27471 = n17187 & n27470;
  assign n27472 = ~n27466 & n27469;
  assign n27473 = ~n27295 & ~n35880;
  assign n27474 = ~n17187 & ~n27470;
  assign n27475 = n16428 & ~n27474;
  assign n27476 = ~n27473 & n27475;
  assign n27477 = ~n26280 & ~n35719;
  assign n27478 = ~n26280 & ~n27055;
  assign n27479 = ~n35719 & n27478;
  assign n27480 = ~n27055 & n27477;
  assign n27481 = ~n35721 & ~n35881;
  assign n27482 = n26295 & n27478;
  assign n27483 = n35721 & n35881;
  assign n27484 = ~n26280 & ~n35721;
  assign n27485 = ~n35719 & n27484;
  assign n27486 = ~n27055 & n27485;
  assign n27487 = n35721 & ~n35881;
  assign n27488 = ~n27486 & ~n27487;
  assign n27489 = ~n27481 & ~n35882;
  assign n27490 = ~n27476 & ~n35883;
  assign n27491 = ~n27473 & ~n27474;
  assign n27492 = ~n16428 & ~n27491;
  assign n27493 = n15760 & ~n27492;
  assign n27494 = ~n27490 & ~n27492;
  assign n27495 = n15760 & n27494;
  assign n27496 = ~n27490 & n27493;
  assign n27497 = ~n27287 & ~n35884;
  assign n27498 = ~n15760 & ~n27494;
  assign n27499 = n15033 & ~n27498;
  assign n27500 = ~n27497 & n27499;
  assign n27501 = ~n26314 & ~n35724;
  assign n27502 = ~n27055 & n27501;
  assign n27503 = ~n35727 & ~n27502;
  assign n27504 = ~n26314 & n35727;
  assign n27505 = ~n35724 & n27504;
  assign n27506 = n35727 & n27502;
  assign n27507 = ~n27055 & n27505;
  assign n27508 = ~n27503 & ~n35885;
  assign n27509 = ~n27500 & ~n27508;
  assign n27510 = ~n27497 & ~n27498;
  assign n27511 = ~n15033 & ~n27510;
  assign n27512 = n14394 & ~n27511;
  assign n27513 = ~n27509 & ~n27511;
  assign n27514 = n14394 & n27513;
  assign n27515 = ~n27509 & n27512;
  assign n27516 = ~n27279 & ~n35886;
  assign n27517 = ~n14394 & ~n27513;
  assign n27518 = n13704 & ~n27517;
  assign n27519 = ~n27516 & n27518;
  assign n27520 = ~n26350 & ~n35730;
  assign n27521 = ~n26350 & ~n27055;
  assign n27522 = ~n35730 & n27521;
  assign n27523 = ~n27055 & n27520;
  assign n27524 = n26361 & ~n35887;
  assign n27525 = n26362 & n27521;
  assign n27526 = ~n26361 & n35887;
  assign n27527 = ~n26350 & n26361;
  assign n27528 = ~n35730 & n27527;
  assign n27529 = ~n27055 & n27528;
  assign n27530 = ~n26361 & ~n35887;
  assign n27531 = ~n27529 & ~n27530;
  assign n27532 = ~n27524 & ~n35888;
  assign n27533 = ~n27519 & ~n35889;
  assign n27534 = ~n27516 & ~n27517;
  assign n27535 = ~n13704 & ~n27534;
  assign n27536 = n13099 & ~n27535;
  assign n27537 = ~n27533 & ~n27535;
  assign n27538 = n13099 & n27537;
  assign n27539 = ~n27533 & n27536;
  assign n27540 = ~n27271 & ~n35890;
  assign n27541 = ~n13099 & ~n27537;
  assign n27542 = n12442 & ~n27541;
  assign n27543 = ~n27540 & n27542;
  assign n27544 = ~n26381 & ~n35734;
  assign n27545 = ~n27055 & n27544;
  assign n27546 = ~n35737 & n27545;
  assign n27547 = n35737 & ~n27545;
  assign n27548 = ~n26381 & n35737;
  assign n27549 = ~n35734 & n27548;
  assign n27550 = n35737 & n27545;
  assign n27551 = ~n27055 & n27549;
  assign n27552 = ~n35737 & ~n27545;
  assign n27553 = ~n35891 & ~n27552;
  assign n27554 = ~n27546 & ~n27547;
  assign n27555 = ~n27543 & ~n35892;
  assign n27556 = ~n27540 & ~n27541;
  assign n27557 = ~n12442 & ~n27556;
  assign n27558 = n11858 & ~n27557;
  assign n27559 = ~n27555 & ~n27557;
  assign n27560 = n11858 & n27559;
  assign n27561 = ~n27555 & n27558;
  assign n27562 = ~n27263 & ~n35893;
  assign n27563 = ~n11858 & ~n27559;
  assign n27564 = n11229 & ~n27563;
  assign n27565 = ~n27562 & n27564;
  assign n27566 = ~n26417 & ~n35740;
  assign n27567 = ~n26417 & ~n27055;
  assign n27568 = ~n35740 & n27567;
  assign n27569 = ~n27055 & n27566;
  assign n27570 = n35742 & ~n35894;
  assign n27571 = n26432 & n27567;
  assign n27572 = ~n35742 & n35894;
  assign n27573 = ~n26417 & n35742;
  assign n27574 = ~n35740 & n27573;
  assign n27575 = ~n27055 & n27574;
  assign n27576 = ~n35742 & ~n35894;
  assign n27577 = ~n27575 & ~n27576;
  assign n27578 = ~n27570 & ~n35895;
  assign n27579 = ~n27565 & ~n35896;
  assign n27580 = ~n27562 & ~n27563;
  assign n27581 = ~n11229 & ~n27580;
  assign n27582 = n10681 & ~n27581;
  assign n27583 = ~n27579 & ~n27581;
  assign n27584 = n10681 & n27583;
  assign n27585 = ~n27579 & n27582;
  assign n27586 = ~n27255 & ~n35897;
  assign n27587 = ~n10681 & ~n27583;
  assign n27588 = n10086 & ~n27587;
  assign n27589 = ~n27586 & n27588;
  assign n27590 = ~n27247 & ~n27589;
  assign n27591 = ~n27586 & ~n27587;
  assign n27592 = ~n10086 & ~n27591;
  assign n27593 = n9565 & ~n27592;
  assign n27594 = ~n27590 & ~n27592;
  assign n27595 = n9565 & n27594;
  assign n27596 = ~n27590 & n27593;
  assign n27597 = ~n27239 & ~n35898;
  assign n27598 = ~n9565 & ~n27594;
  assign n27599 = n8998 & ~n27598;
  assign n27600 = ~n27597 & n27599;
  assign n27601 = ~n26487 & ~n35752;
  assign n27602 = ~n26487 & ~n27055;
  assign n27603 = ~n35752 & n27602;
  assign n27604 = ~n27055 & n27601;
  assign n27605 = n26495 & ~n35899;
  assign n27606 = n26499 & n27602;
  assign n27607 = ~n26487 & n26495;
  assign n27608 = ~n35752 & n27607;
  assign n27609 = ~n27055 & n27608;
  assign n27610 = ~n26495 & ~n35899;
  assign n27611 = ~n27609 & ~n27610;
  assign n27612 = ~n27605 & ~n27606;
  assign n27613 = ~n27600 & ~n35900;
  assign n27614 = ~n27597 & ~n27598;
  assign n27615 = ~n8998 & ~n27614;
  assign n27616 = n8506 & ~n27615;
  assign n27617 = ~n27613 & ~n27615;
  assign n27618 = n8506 & n27617;
  assign n27619 = ~n27613 & n27616;
  assign n27620 = ~n27231 & ~n35901;
  assign n27621 = ~n8506 & ~n27617;
  assign n27622 = n7975 & ~n27621;
  assign n27623 = ~n27620 & n27622;
  assign n27624 = ~n27223 & ~n27623;
  assign n27625 = ~n27620 & ~n27621;
  assign n27626 = ~n7975 & ~n27625;
  assign n27627 = n7512 & ~n27626;
  assign n27628 = ~n27624 & ~n27626;
  assign n27629 = n7512 & n27628;
  assign n27630 = ~n27624 & n27627;
  assign n27631 = ~n27215 & ~n35902;
  assign n27632 = ~n7512 & ~n27628;
  assign n27633 = n7015 & ~n27632;
  assign n27634 = ~n27631 & n27633;
  assign n27635 = ~n26553 & ~n35761;
  assign n27636 = ~n26553 & ~n27055;
  assign n27637 = ~n35761 & n27636;
  assign n27638 = ~n27055 & n27635;
  assign n27639 = n26561 & ~n35903;
  assign n27640 = n26565 & n27636;
  assign n27641 = ~n26553 & n26561;
  assign n27642 = ~n35761 & n27641;
  assign n27643 = ~n27055 & n27642;
  assign n27644 = ~n26561 & ~n35903;
  assign n27645 = ~n27643 & ~n27644;
  assign n27646 = ~n27639 & ~n27640;
  assign n27647 = ~n27634 & ~n35904;
  assign n27648 = ~n27631 & ~n27632;
  assign n27649 = ~n7015 & ~n27648;
  assign n27650 = n6579 & ~n27649;
  assign n27651 = ~n27647 & ~n27649;
  assign n27652 = n6579 & n27651;
  assign n27653 = ~n27647 & n27650;
  assign n27654 = ~n27207 & ~n35905;
  assign n27655 = ~n6579 & ~n27651;
  assign n27656 = n6117 & ~n27655;
  assign n27657 = ~n27654 & n27656;
  assign n27658 = ~n27199 & ~n27657;
  assign n27659 = ~n27654 & ~n27655;
  assign n27660 = ~n6117 & ~n27659;
  assign n27661 = n5708 & ~n27660;
  assign n27662 = ~n27658 & ~n27660;
  assign n27663 = n5708 & n27662;
  assign n27664 = ~n27658 & n27661;
  assign n27665 = ~n27191 & ~n35906;
  assign n27666 = ~n5708 & ~n27662;
  assign n27667 = n5278 & ~n27666;
  assign n27668 = ~n27665 & n27667;
  assign n27669 = ~n26619 & ~n35770;
  assign n27670 = ~n26619 & ~n27055;
  assign n27671 = ~n35770 & n27670;
  assign n27672 = ~n27055 & n27669;
  assign n27673 = n26627 & ~n35907;
  assign n27674 = n26631 & n27670;
  assign n27675 = ~n26619 & n26627;
  assign n27676 = ~n35770 & n27675;
  assign n27677 = ~n27055 & n27676;
  assign n27678 = ~n26627 & ~n35907;
  assign n27679 = ~n27677 & ~n27678;
  assign n27680 = ~n27673 & ~n27674;
  assign n27681 = ~n27668 & ~n35908;
  assign n27682 = ~n27665 & ~n27666;
  assign n27683 = ~n5278 & ~n27682;
  assign n27684 = n4903 & ~n27683;
  assign n27685 = ~n27681 & ~n27683;
  assign n27686 = n4903 & n27685;
  assign n27687 = ~n27681 & n27684;
  assign n27688 = ~n27183 & ~n35909;
  assign n27689 = ~n4903 & ~n27685;
  assign n27690 = n4508 & ~n27689;
  assign n27691 = ~n27688 & n27690;
  assign n27692 = ~n27175 & ~n27691;
  assign n27693 = ~n27688 & ~n27689;
  assign n27694 = ~n4508 & ~n27693;
  assign n27695 = n4155 & ~n27694;
  assign n27696 = ~n27692 & ~n27694;
  assign n27697 = n4155 & n27696;
  assign n27698 = ~n27692 & n27695;
  assign n27699 = ~n27167 & ~n35910;
  assign n27700 = ~n4155 & ~n27696;
  assign n27701 = n3788 & ~n27700;
  assign n27702 = ~n27699 & n27701;
  assign n27703 = ~n26685 & ~n35779;
  assign n27704 = ~n26685 & ~n27055;
  assign n27705 = ~n35779 & n27704;
  assign n27706 = ~n27055 & n27703;
  assign n27707 = n26693 & ~n35911;
  assign n27708 = n26697 & n27704;
  assign n27709 = ~n26685 & n26693;
  assign n27710 = ~n35779 & n27709;
  assign n27711 = ~n27055 & n27710;
  assign n27712 = ~n26693 & ~n35911;
  assign n27713 = ~n27711 & ~n27712;
  assign n27714 = ~n27707 & ~n27708;
  assign n27715 = ~n27702 & ~n35912;
  assign n27716 = ~n27699 & ~n27700;
  assign n27717 = ~n3788 & ~n27716;
  assign n27718 = n3473 & ~n27717;
  assign n27719 = ~n27715 & ~n27717;
  assign n27720 = n3473 & n27719;
  assign n27721 = ~n27715 & n27718;
  assign n27722 = ~n27159 & ~n35913;
  assign n27723 = ~n3473 & ~n27719;
  assign n27724 = n3140 & ~n27723;
  assign n27725 = ~n27722 & n27724;
  assign n27726 = ~n27151 & ~n27725;
  assign n27727 = ~n27722 & ~n27723;
  assign n27728 = ~n3140 & ~n27727;
  assign n27729 = n2855 & ~n27728;
  assign n27730 = ~n27726 & ~n27728;
  assign n27731 = n2855 & n27730;
  assign n27732 = ~n27726 & n27729;
  assign n27733 = ~n27143 & ~n35914;
  assign n27734 = ~n2855 & ~n27730;
  assign n27735 = n2556 & ~n27734;
  assign n27736 = ~n27733 & n27735;
  assign n27737 = ~n26751 & ~n35788;
  assign n27738 = ~n26751 & ~n27055;
  assign n27739 = ~n35788 & n27738;
  assign n27740 = ~n27055 & n27737;
  assign n27741 = n26759 & ~n35915;
  assign n27742 = n26763 & n27738;
  assign n27743 = ~n26751 & n26759;
  assign n27744 = ~n35788 & n27743;
  assign n27745 = ~n27055 & n27744;
  assign n27746 = ~n26759 & ~n35915;
  assign n27747 = ~n27745 & ~n27746;
  assign n27748 = ~n27741 & ~n27742;
  assign n27749 = ~n27736 & ~n35916;
  assign n27750 = ~n27733 & ~n27734;
  assign n27751 = ~n2556 & ~n27750;
  assign n27752 = n2301 & ~n27751;
  assign n27753 = ~n27749 & ~n27751;
  assign n27754 = n2301 & n27753;
  assign n27755 = ~n27749 & n27752;
  assign n27756 = ~n27135 & ~n35917;
  assign n27757 = ~n2301 & ~n27753;
  assign n27758 = n2038 & ~n27757;
  assign n27759 = ~n27756 & n27758;
  assign n27760 = ~n27127 & ~n27759;
  assign n27761 = ~n27756 & ~n27757;
  assign n27762 = ~n2038 & ~n27761;
  assign n27763 = n1812 & ~n27762;
  assign n27764 = ~n27760 & ~n27762;
  assign n27765 = n1812 & n27764;
  assign n27766 = ~n27760 & n27763;
  assign n27767 = ~n27119 & ~n35918;
  assign n27768 = ~n1812 & ~n27764;
  assign n27769 = n1582 & ~n27768;
  assign n27770 = ~n27767 & n27769;
  assign n27771 = ~n26817 & ~n35797;
  assign n27772 = ~n26817 & ~n27055;
  assign n27773 = ~n35797 & n27772;
  assign n27774 = ~n27055 & n27771;
  assign n27775 = n26825 & ~n35919;
  assign n27776 = n26829 & n27772;
  assign n27777 = ~n26817 & n26825;
  assign n27778 = ~n35797 & n27777;
  assign n27779 = ~n27055 & n27778;
  assign n27780 = ~n26825 & ~n35919;
  assign n27781 = ~n27779 & ~n27780;
  assign n27782 = ~n27775 & ~n27776;
  assign n27783 = ~n27770 & ~n35920;
  assign n27784 = ~n27767 & ~n27768;
  assign n27785 = ~n1582 & ~n27784;
  assign n27786 = n1388 & ~n27785;
  assign n27787 = ~n27783 & ~n27785;
  assign n27788 = n1388 & n27787;
  assign n27789 = ~n27783 & n27786;
  assign n27790 = ~n27111 & ~n35921;
  assign n27791 = ~n1388 & ~n27787;
  assign n27792 = n1192 & ~n27791;
  assign n27793 = ~n27790 & n27792;
  assign n27794 = ~n27103 & ~n27793;
  assign n27795 = ~n27790 & ~n27791;
  assign n27796 = ~n1192 & ~n27795;
  assign n27797 = n1028 & ~n27796;
  assign n27798 = ~n27794 & ~n27796;
  assign n27799 = n1028 & n27798;
  assign n27800 = ~n27794 & n27797;
  assign n27801 = ~n27095 & ~n35922;
  assign n27802 = ~n1028 & ~n27798;
  assign n27803 = n866 & ~n27802;
  assign n27804 = ~n27801 & n27803;
  assign n27805 = ~n26883 & ~n35806;
  assign n27806 = ~n26883 & ~n27055;
  assign n27807 = ~n35806 & n27806;
  assign n27808 = ~n27055 & n27805;
  assign n27809 = n26891 & ~n35923;
  assign n27810 = n26895 & n27806;
  assign n27811 = ~n26883 & n26891;
  assign n27812 = ~n35806 & n27811;
  assign n27813 = ~n27055 & n27812;
  assign n27814 = ~n26891 & ~n35923;
  assign n27815 = ~n27813 & ~n27814;
  assign n27816 = ~n27809 & ~n27810;
  assign n27817 = ~n27804 & ~n35924;
  assign n27818 = ~n27801 & ~n27802;
  assign n27819 = ~n866 & ~n27818;
  assign n27820 = n730 & ~n27819;
  assign n27821 = ~n27817 & ~n27819;
  assign n27822 = n730 & n27821;
  assign n27823 = ~n27817 & n27820;
  assign n27824 = ~n27087 & ~n35925;
  assign n27825 = ~n730 & ~n27821;
  assign n27826 = n602 & ~n27825;
  assign n27827 = ~n27824 & n27826;
  assign n27828 = ~n27079 & ~n27827;
  assign n27829 = ~n27824 & ~n27825;
  assign n27830 = ~n602 & ~n27829;
  assign n27831 = n497 & ~n27830;
  assign n27832 = ~n27828 & ~n27830;
  assign n27833 = n497 & n27832;
  assign n27834 = ~n27828 & n27831;
  assign n27835 = ~n27071 & ~n35926;
  assign n27836 = ~n497 & ~n27832;
  assign n27837 = ~n27835 & ~n27836;
  assign n27838 = ~n403 & ~n27837;
  assign n27839 = n403 & ~n27836;
  assign n27840 = ~n27835 & n27839;
  assign n27841 = ~n26947 & ~n35813;
  assign n27842 = ~n27055 & n27841;
  assign n27843 = n26958 & ~n27842;
  assign n27844 = ~n26958 & n27842;
  assign n27845 = ~n26947 & n26958;
  assign n27846 = ~n35813 & n27845;
  assign n27847 = n26958 & n27842;
  assign n27848 = ~n27055 & n27846;
  assign n27849 = ~n26958 & ~n27842;
  assign n27850 = ~n35927 & ~n27849;
  assign n27851 = ~n27843 & ~n27844;
  assign n27852 = ~n27840 & ~n35928;
  assign n27853 = ~n27838 & ~n27852;
  assign n27854 = ~n330 & ~n27853;
  assign n27855 = n330 & ~n27838;
  assign n27856 = n330 & n27853;
  assign n27857 = ~n27852 & n27855;
  assign n27858 = ~n27063 & ~n35929;
  assign n27859 = ~n27854 & ~n27858;
  assign n27860 = ~n271 & ~n27859;
  assign n27861 = n271 & ~n27854;
  assign n27862 = ~n27858 & n27861;
  assign n27863 = ~n26966 & ~n35816;
  assign n27864 = ~n26966 & ~n27055;
  assign n27865 = ~n35816 & n27864;
  assign n27866 = ~n27055 & n27863;
  assign n27867 = n26974 & ~n35930;
  assign n27868 = n26978 & n27864;
  assign n27869 = ~n26966 & n26974;
  assign n27870 = ~n35816 & n27869;
  assign n27871 = ~n27055 & n27870;
  assign n27872 = ~n26974 & ~n35930;
  assign n27873 = ~n27871 & ~n27872;
  assign n27874 = ~n27867 & ~n27868;
  assign n27875 = ~n27862 & ~n35931;
  assign n27876 = ~n27860 & ~n27875;
  assign n27877 = ~n217 & ~n27876;
  assign n27878 = ~n26980 & ~n26982;
  assign n27879 = ~n27055 & n27878;
  assign n27880 = ~n35818 & ~n27879;
  assign n27881 = ~n26982 & n35818;
  assign n27882 = ~n26980 & n27881;
  assign n27883 = n35818 & n27879;
  assign n27884 = ~n27055 & n27882;
  assign n27885 = ~n27880 & ~n35932;
  assign n27886 = n217 & ~n27860;
  assign n27887 = n217 & n27876;
  assign n27888 = ~n27875 & n27886;
  assign n27889 = ~n27885 & ~n35933;
  assign n27890 = ~n27877 & ~n27889;
  assign n27891 = ~n198 & ~n27890;
  assign n27892 = n198 & ~n27877;
  assign n27893 = ~n27889 & n27892;
  assign n27894 = ~n26997 & ~n35820;
  assign n27895 = ~n26997 & ~n27055;
  assign n27896 = ~n35820 & n27895;
  assign n27897 = ~n27055 & n27894;
  assign n27898 = n27005 & ~n35934;
  assign n27899 = n27009 & n27895;
  assign n27900 = ~n26997 & n27005;
  assign n27901 = ~n35820 & n27900;
  assign n27902 = ~n27055 & n27901;
  assign n27903 = ~n27005 & ~n35934;
  assign n27904 = ~n27902 & ~n27903;
  assign n27905 = ~n27898 & ~n27899;
  assign n27906 = ~n27893 & ~n35935;
  assign n27907 = ~n27891 & ~n27906;
  assign n27908 = ~n27011 & ~n27013;
  assign n27909 = ~n27055 & n27908;
  assign n27910 = ~n35822 & ~n27909;
  assign n27911 = ~n27013 & n35822;
  assign n27912 = ~n27011 & n27911;
  assign n27913 = n35822 & n27909;
  assign n27914 = ~n27055 & n27912;
  assign n27915 = ~n27910 & ~n35936;
  assign n27916 = ~n27027 & ~n35824;
  assign n27917 = ~n35824 & ~n27055;
  assign n27918 = ~n27027 & n27917;
  assign n27919 = ~n27055 & n27916;
  assign n27920 = ~n35826 & ~n35937;
  assign n27921 = ~n27915 & n27920;
  assign n27922 = ~n27907 & n27921;
  assign n27923 = n193 & ~n27922;
  assign n27924 = ~n27891 & n27915;
  assign n27925 = n27907 & n27915;
  assign n27926 = ~n27906 & n27924;
  assign n27927 = n27027 & ~n27917;
  assign n27928 = ~n193 & ~n27916;
  assign n27929 = ~n27927 & n27928;
  assign n27930 = ~n35938 & ~n27929;
  assign n27931 = ~n27923 & n27930;
  assign n27932 = ~n27854 & ~n35929;
  assign n27933 = ~n27854 & ~n27931;
  assign n27934 = ~n35929 & n27933;
  assign n27935 = ~n27931 & n27932;
  assign n27936 = n27063 & ~n35939;
  assign n27937 = n27858 & n27933;
  assign n27938 = n27063 & ~n35929;
  assign n27939 = ~n27854 & n27938;
  assign n27940 = ~n27931 & n27939;
  assign n27941 = ~n27063 & ~n35939;
  assign n27942 = ~n27940 & ~n27941;
  assign n27943 = ~n27936 & ~n27937;
  assign n27944 = pi8  & ~n27931;
  assign n27945 = ~pi6  & ~pi7 ;
  assign n27946 = ~pi8  & n27945;
  assign n27947 = ~pi8  & ~n27945;
  assign n27948 = pi8  & n27931;
  assign n27949 = ~n27947 & ~n27948;
  assign n27950 = ~n27944 & ~n27946;
  assign n27951 = ~n27055 & n35941;
  assign n27952 = ~pi8  & ~n27931;
  assign n27953 = pi9  & ~n27952;
  assign n27954 = ~pi9  & n27952;
  assign n27955 = n27342 & ~n27931;
  assign n27956 = ~n27953 & ~n35942;
  assign n27957 = ~n27053 & ~n27946;
  assign n27958 = ~n35826 & n27957;
  assign n27959 = ~n27047 & n27958;
  assign n27960 = n27055 & ~n35941;
  assign n27961 = ~n27944 & n27959;
  assign n27962 = n27956 & ~n35943;
  assign n27963 = ~n27951 & ~n27962;
  assign n27964 = ~n26098 & ~n27963;
  assign n27965 = n26098 & ~n27951;
  assign n27966 = ~n27962 & n27965;
  assign n27967 = ~n27055 & ~n27929;
  assign n27968 = ~n35938 & n27967;
  assign n27969 = ~n27055 & n27931;
  assign n27970 = ~n27923 & n27968;
  assign n27971 = ~n35942 & ~n35944;
  assign n27972 = pi10  & ~n27971;
  assign n27973 = ~pi10  & ~n35944;
  assign n27974 = ~pi10  & n27971;
  assign n27975 = ~n35942 & n27973;
  assign n27976 = ~n27972 & ~n35945;
  assign n27977 = ~n27966 & ~n27976;
  assign n27978 = ~n27964 & ~n27977;
  assign n27979 = ~n25256 & ~n27978;
  assign n27980 = n25256 & ~n27964;
  assign n27981 = ~n27977 & n27980;
  assign n27982 = n25256 & n27978;
  assign n27983 = ~n35866 & ~n27363;
  assign n27984 = ~n27931 & n27983;
  assign n27985 = n27361 & ~n27984;
  assign n27986 = ~n27361 & n27983;
  assign n27987 = ~n27361 & n27984;
  assign n27988 = ~n27931 & n27986;
  assign n27989 = ~n27985 & ~n35947;
  assign n27990 = ~n35946 & ~n27989;
  assign n27991 = ~n27979 & ~n27990;
  assign n27992 = ~n24331 & ~n27991;
  assign n27993 = n24331 & ~n27979;
  assign n27994 = ~n27990 & n27993;
  assign n27995 = ~n35867 & ~n27369;
  assign n27996 = ~n27369 & ~n27931;
  assign n27997 = ~n35867 & n27996;
  assign n27998 = ~n27931 & n27995;
  assign n27999 = n27340 & ~n35948;
  assign n28000 = n27368 & n27996;
  assign n28001 = n27340 & ~n35867;
  assign n28002 = ~n27369 & n28001;
  assign n28003 = ~n27931 & n28002;
  assign n28004 = ~n27340 & ~n35948;
  assign n28005 = ~n28003 & ~n28004;
  assign n28006 = ~n27999 & ~n28000;
  assign n28007 = ~n27994 & ~n35949;
  assign n28008 = ~n27992 & ~n28007;
  assign n28009 = ~n23517 & ~n28008;
  assign n28010 = n23517 & ~n27992;
  assign n28011 = ~n28007 & n28010;
  assign n28012 = n23517 & n28008;
  assign n28013 = ~n27371 & ~n27381;
  assign n28014 = ~n27931 & n28013;
  assign n28015 = n27378 & ~n28014;
  assign n28016 = ~n27378 & n28014;
  assign n28017 = n27378 & ~n27381;
  assign n28018 = ~n27371 & n28017;
  assign n28019 = n27378 & n28014;
  assign n28020 = ~n27931 & n28018;
  assign n28021 = ~n27378 & ~n28014;
  assign n28022 = ~n35951 & ~n28021;
  assign n28023 = ~n28015 & ~n28016;
  assign n28024 = ~n35950 & ~n35952;
  assign n28025 = ~n28009 & ~n28024;
  assign n28026 = ~n22625 & ~n28025;
  assign n28027 = n22625 & ~n28009;
  assign n28028 = ~n28024 & n28027;
  assign n28029 = ~n35869 & ~n27387;
  assign n28030 = ~n27387 & ~n27931;
  assign n28031 = ~n35869 & n28030;
  assign n28032 = ~n27931 & n28029;
  assign n28033 = n27327 & ~n35953;
  assign n28034 = n27386 & n28030;
  assign n28035 = n27327 & ~n35869;
  assign n28036 = ~n27387 & n28035;
  assign n28037 = ~n27931 & n28036;
  assign n28038 = ~n27327 & ~n35953;
  assign n28039 = ~n28037 & ~n28038;
  assign n28040 = ~n28033 & ~n28034;
  assign n28041 = ~n28028 & ~n35954;
  assign n28042 = ~n28026 & ~n28041;
  assign n28043 = ~n21842 & ~n28042;
  assign n28044 = n21842 & ~n28026;
  assign n28045 = ~n28041 & n28044;
  assign n28046 = n21842 & n28042;
  assign n28047 = ~n27389 & ~n27403;
  assign n28048 = ~n27931 & n28047;
  assign n28049 = ~n35871 & n28048;
  assign n28050 = n35871 & ~n28048;
  assign n28051 = n35871 & ~n27403;
  assign n28052 = ~n27389 & n28051;
  assign n28053 = ~n27931 & n28052;
  assign n28054 = ~n35871 & ~n28048;
  assign n28055 = ~n28053 & ~n28054;
  assign n28056 = ~n28049 & ~n28050;
  assign n28057 = ~n35955 & ~n35956;
  assign n28058 = ~n28043 & ~n28057;
  assign n28059 = ~n20986 & ~n28058;
  assign n28060 = n20986 & ~n28043;
  assign n28061 = ~n28057 & n28060;
  assign n28062 = ~n35872 & ~n27409;
  assign n28063 = ~n27409 & ~n27931;
  assign n28064 = ~n35872 & n28063;
  assign n28065 = ~n27931 & n28062;
  assign n28066 = n27319 & ~n35957;
  assign n28067 = n27408 & n28063;
  assign n28068 = n27319 & ~n35872;
  assign n28069 = ~n27409 & n28068;
  assign n28070 = ~n27931 & n28069;
  assign n28071 = ~n27319 & ~n35957;
  assign n28072 = ~n28070 & ~n28071;
  assign n28073 = ~n28066 & ~n28067;
  assign n28074 = ~n28061 & ~n35958;
  assign n28075 = ~n28059 & ~n28074;
  assign n28076 = ~n20229 & ~n28075;
  assign n28077 = n20229 & ~n28059;
  assign n28078 = ~n28074 & n28077;
  assign n28079 = n20229 & n28075;
  assign n28080 = ~n27411 & ~n27424;
  assign n28081 = ~n27931 & n28080;
  assign n28082 = ~n35873 & ~n28081;
  assign n28083 = n35873 & ~n27424;
  assign n28084 = ~n27411 & n28083;
  assign n28085 = n35873 & n28081;
  assign n28086 = ~n27931 & n28084;
  assign n28087 = n35873 & ~n28081;
  assign n28088 = ~n35873 & n28081;
  assign n28089 = ~n28087 & ~n28088;
  assign n28090 = ~n28082 & ~n35960;
  assign n28091 = ~n35959 & n35961;
  assign n28092 = ~n28076 & ~n28091;
  assign n28093 = ~n19401 & ~n28092;
  assign n28094 = n19401 & ~n28076;
  assign n28095 = ~n28091 & n28094;
  assign n28096 = ~n35874 & ~n27430;
  assign n28097 = ~n27430 & ~n27931;
  assign n28098 = ~n35874 & n28097;
  assign n28099 = ~n27931 & n28096;
  assign n28100 = n27311 & ~n35962;
  assign n28101 = n27429 & n28097;
  assign n28102 = n27311 & ~n35874;
  assign n28103 = ~n27430 & n28102;
  assign n28104 = ~n27931 & n28103;
  assign n28105 = ~n27311 & ~n35962;
  assign n28106 = ~n28104 & ~n28105;
  assign n28107 = ~n28100 & ~n28101;
  assign n28108 = ~n28095 & ~n35963;
  assign n28109 = ~n28093 & ~n28108;
  assign n28110 = ~n18676 & ~n28109;
  assign n28111 = n18676 & ~n28093;
  assign n28112 = ~n28108 & n28111;
  assign n28113 = n18676 & n28109;
  assign n28114 = ~n27432 & ~n27446;
  assign n28115 = ~n27931 & n28114;
  assign n28116 = n35876 & ~n28115;
  assign n28117 = ~n35876 & ~n27446;
  assign n28118 = ~n27432 & n28117;
  assign n28119 = ~n35876 & n28115;
  assign n28120 = ~n27931 & n28118;
  assign n28121 = n35876 & n28115;
  assign n28122 = ~n35876 & ~n28115;
  assign n28123 = ~n28121 & ~n28122;
  assign n28124 = ~n28116 & ~n35965;
  assign n28125 = ~n35964 & n35966;
  assign n28126 = ~n28110 & ~n28125;
  assign n28127 = ~n17885 & ~n28126;
  assign n28128 = n17885 & ~n28110;
  assign n28129 = ~n28125 & n28128;
  assign n28130 = ~n35877 & ~n27452;
  assign n28131 = ~n27452 & ~n27931;
  assign n28132 = ~n35877 & n28131;
  assign n28133 = ~n27931 & n28130;
  assign n28134 = n27303 & ~n35967;
  assign n28135 = n27451 & n28131;
  assign n28136 = n27303 & ~n35877;
  assign n28137 = ~n27452 & n28136;
  assign n28138 = ~n27931 & n28137;
  assign n28139 = ~n27303 & ~n35967;
  assign n28140 = ~n28138 & ~n28139;
  assign n28141 = ~n28134 & ~n28135;
  assign n28142 = ~n28129 & ~n35968;
  assign n28143 = ~n28127 & ~n28142;
  assign n28144 = ~n17187 & ~n28143;
  assign n28145 = n17187 & ~n28127;
  assign n28146 = ~n28142 & n28145;
  assign n28147 = n17187 & n28143;
  assign n28148 = ~n27454 & ~n27468;
  assign n28149 = ~n27468 & ~n27931;
  assign n28150 = ~n27454 & n28149;
  assign n28151 = ~n27931 & n28148;
  assign n28152 = ~n35879 & ~n35970;
  assign n28153 = n27466 & n28149;
  assign n28154 = n35879 & n35970;
  assign n28155 = ~n35879 & ~n27468;
  assign n28156 = ~n27454 & n28155;
  assign n28157 = ~n27931 & n28156;
  assign n28158 = n35879 & ~n35970;
  assign n28159 = ~n28157 & ~n28158;
  assign n28160 = ~n28152 & ~n35971;
  assign n28161 = ~n35969 & ~n35972;
  assign n28162 = ~n28144 & ~n28161;
  assign n28163 = ~n16428 & ~n28162;
  assign n28164 = n16428 & ~n28144;
  assign n28165 = ~n28161 & n28164;
  assign n28166 = ~n35880 & ~n27474;
  assign n28167 = ~n27474 & ~n27931;
  assign n28168 = ~n35880 & n28167;
  assign n28169 = ~n27931 & n28166;
  assign n28170 = n27295 & ~n35973;
  assign n28171 = n27473 & n28167;
  assign n28172 = n27295 & ~n35880;
  assign n28173 = ~n27474 & n28172;
  assign n28174 = ~n27931 & n28173;
  assign n28175 = ~n27295 & ~n35973;
  assign n28176 = ~n28174 & ~n28175;
  assign n28177 = ~n28170 & ~n28171;
  assign n28178 = ~n28165 & ~n35974;
  assign n28179 = ~n28163 & ~n28178;
  assign n28180 = ~n15760 & ~n28179;
  assign n28181 = n15760 & ~n28163;
  assign n28182 = ~n28178 & n28181;
  assign n28183 = n15760 & n28179;
  assign n28184 = ~n27476 & ~n27492;
  assign n28185 = ~n27931 & n28184;
  assign n28186 = ~n35883 & ~n28185;
  assign n28187 = n35883 & ~n27492;
  assign n28188 = ~n27476 & n28187;
  assign n28189 = n35883 & n28185;
  assign n28190 = ~n27931 & n28188;
  assign n28191 = ~n28186 & ~n35976;
  assign n28192 = ~n35975 & ~n28191;
  assign n28193 = ~n28180 & ~n28192;
  assign n28194 = ~n15033 & ~n28193;
  assign n28195 = n15033 & ~n28180;
  assign n28196 = ~n28192 & n28195;
  assign n28197 = ~n35884 & ~n27498;
  assign n28198 = ~n27498 & ~n27931;
  assign n28199 = ~n35884 & n28198;
  assign n28200 = ~n27931 & n28197;
  assign n28201 = n27287 & ~n35977;
  assign n28202 = n27497 & n28198;
  assign n28203 = n27287 & ~n35884;
  assign n28204 = ~n27498 & n28203;
  assign n28205 = ~n27931 & n28204;
  assign n28206 = ~n27287 & ~n35977;
  assign n28207 = ~n28205 & ~n28206;
  assign n28208 = ~n28201 & ~n28202;
  assign n28209 = ~n28196 & ~n35978;
  assign n28210 = ~n28194 & ~n28209;
  assign n28211 = ~n14394 & ~n28210;
  assign n28212 = n14394 & ~n28194;
  assign n28213 = ~n28209 & n28212;
  assign n28214 = n14394 & n28210;
  assign n28215 = ~n27500 & ~n27511;
  assign n28216 = ~n27511 & ~n27931;
  assign n28217 = ~n27500 & n28216;
  assign n28218 = ~n27931 & n28215;
  assign n28219 = n27508 & ~n35980;
  assign n28220 = n27509 & n28216;
  assign n28221 = ~n27508 & n35980;
  assign n28222 = n27508 & ~n27511;
  assign n28223 = ~n27500 & n28222;
  assign n28224 = ~n27931 & n28223;
  assign n28225 = ~n27508 & ~n35980;
  assign n28226 = ~n28224 & ~n28225;
  assign n28227 = ~n28219 & ~n35981;
  assign n28228 = ~n35979 & ~n35982;
  assign n28229 = ~n28211 & ~n28228;
  assign n28230 = ~n13704 & ~n28229;
  assign n28231 = n13704 & ~n28211;
  assign n28232 = ~n28228 & n28231;
  assign n28233 = ~n35886 & ~n27517;
  assign n28234 = ~n27517 & ~n27931;
  assign n28235 = ~n35886 & n28234;
  assign n28236 = ~n27931 & n28233;
  assign n28237 = n27279 & ~n35983;
  assign n28238 = n27516 & n28234;
  assign n28239 = n27279 & ~n35886;
  assign n28240 = ~n27517 & n28239;
  assign n28241 = ~n27931 & n28240;
  assign n28242 = ~n27279 & ~n35983;
  assign n28243 = ~n28241 & ~n28242;
  assign n28244 = ~n28237 & ~n28238;
  assign n28245 = ~n28232 & ~n35984;
  assign n28246 = ~n28230 & ~n28245;
  assign n28247 = ~n13099 & ~n28246;
  assign n28248 = n13099 & ~n28230;
  assign n28249 = ~n28245 & n28248;
  assign n28250 = n13099 & n28246;
  assign n28251 = ~n27519 & ~n27535;
  assign n28252 = ~n27931 & n28251;
  assign n28253 = ~n35889 & n28252;
  assign n28254 = n35889 & ~n28252;
  assign n28255 = n35889 & ~n27535;
  assign n28256 = ~n27519 & n28255;
  assign n28257 = n35889 & n28252;
  assign n28258 = ~n27931 & n28256;
  assign n28259 = ~n35889 & ~n28252;
  assign n28260 = ~n35986 & ~n28259;
  assign n28261 = ~n28253 & ~n28254;
  assign n28262 = ~n35985 & ~n35987;
  assign n28263 = ~n28247 & ~n28262;
  assign n28264 = ~n12442 & ~n28263;
  assign n28265 = n12442 & ~n28247;
  assign n28266 = ~n28262 & n28265;
  assign n28267 = ~n35890 & ~n27541;
  assign n28268 = ~n27541 & ~n27931;
  assign n28269 = ~n35890 & n28268;
  assign n28270 = ~n27931 & n28267;
  assign n28271 = n27271 & ~n35988;
  assign n28272 = n27540 & n28268;
  assign n28273 = n27271 & ~n35890;
  assign n28274 = ~n27541 & n28273;
  assign n28275 = ~n27931 & n28274;
  assign n28276 = ~n27271 & ~n35988;
  assign n28277 = ~n28275 & ~n28276;
  assign n28278 = ~n28271 & ~n28272;
  assign n28279 = ~n28266 & ~n35989;
  assign n28280 = ~n28264 & ~n28279;
  assign n28281 = ~n11858 & ~n28280;
  assign n28282 = n11858 & ~n28264;
  assign n28283 = ~n28279 & n28282;
  assign n28284 = n11858 & n28280;
  assign n28285 = ~n27543 & ~n27557;
  assign n28286 = ~n27557 & ~n27931;
  assign n28287 = ~n27543 & n28286;
  assign n28288 = ~n27931 & n28285;
  assign n28289 = n35892 & ~n35991;
  assign n28290 = n27555 & n28286;
  assign n28291 = ~n35892 & n35991;
  assign n28292 = n35892 & ~n27557;
  assign n28293 = ~n27543 & n28292;
  assign n28294 = ~n27931 & n28293;
  assign n28295 = ~n35892 & ~n35991;
  assign n28296 = ~n28294 & ~n28295;
  assign n28297 = ~n28289 & ~n35992;
  assign n28298 = ~n35990 & ~n35993;
  assign n28299 = ~n28281 & ~n28298;
  assign n28300 = ~n11229 & ~n28299;
  assign n28301 = n11229 & ~n28281;
  assign n28302 = ~n28298 & n28301;
  assign n28303 = ~n35893 & ~n27563;
  assign n28304 = ~n27563 & ~n27931;
  assign n28305 = ~n35893 & n28304;
  assign n28306 = ~n27931 & n28303;
  assign n28307 = n27263 & ~n35994;
  assign n28308 = n27562 & n28304;
  assign n28309 = n27263 & ~n35893;
  assign n28310 = ~n27563 & n28309;
  assign n28311 = ~n27931 & n28310;
  assign n28312 = ~n27263 & ~n35994;
  assign n28313 = ~n28311 & ~n28312;
  assign n28314 = ~n28307 & ~n28308;
  assign n28315 = ~n28302 & ~n35995;
  assign n28316 = ~n28300 & ~n28315;
  assign n28317 = ~n10681 & ~n28316;
  assign n28318 = ~n27565 & ~n27581;
  assign n28319 = ~n27931 & n28318;
  assign n28320 = ~n35896 & ~n28319;
  assign n28321 = n35896 & ~n27581;
  assign n28322 = ~n27565 & n28321;
  assign n28323 = n35896 & n28319;
  assign n28324 = ~n27931 & n28322;
  assign n28325 = ~n28320 & ~n35996;
  assign n28326 = n10681 & ~n28300;
  assign n28327 = ~n28315 & n28326;
  assign n28328 = n10681 & n28316;
  assign n28329 = ~n28325 & ~n35997;
  assign n28330 = ~n28317 & ~n28329;
  assign n28331 = ~n10086 & ~n28330;
  assign n28332 = n10086 & ~n28317;
  assign n28333 = ~n28329 & n28332;
  assign n28334 = ~n35897 & ~n27587;
  assign n28335 = ~n27587 & ~n27931;
  assign n28336 = ~n35897 & n28335;
  assign n28337 = ~n27931 & n28334;
  assign n28338 = n27255 & ~n35998;
  assign n28339 = n27586 & n28335;
  assign n28340 = n27255 & ~n35897;
  assign n28341 = ~n27587 & n28340;
  assign n28342 = ~n27931 & n28341;
  assign n28343 = ~n27255 & ~n35998;
  assign n28344 = ~n28342 & ~n28343;
  assign n28345 = ~n28338 & ~n28339;
  assign n28346 = ~n28333 & ~n35999;
  assign n28347 = ~n28331 & ~n28346;
  assign n28348 = ~n9565 & ~n28347;
  assign n28349 = n9565 & ~n28331;
  assign n28350 = ~n28346 & n28349;
  assign n28351 = n9565 & n28347;
  assign n28352 = ~n27589 & ~n27592;
  assign n28353 = ~n27592 & ~n27931;
  assign n28354 = ~n27589 & n28353;
  assign n28355 = ~n27931 & n28352;
  assign n28356 = n27247 & ~n36001;
  assign n28357 = n27590 & n28353;
  assign n28358 = n27247 & ~n27592;
  assign n28359 = ~n27589 & n28358;
  assign n28360 = ~n27931 & n28359;
  assign n28361 = ~n27247 & ~n36001;
  assign n28362 = ~n28360 & ~n28361;
  assign n28363 = ~n28356 & ~n28357;
  assign n28364 = ~n36000 & ~n36002;
  assign n28365 = ~n28348 & ~n28364;
  assign n28366 = ~n8998 & ~n28365;
  assign n28367 = n8998 & ~n28348;
  assign n28368 = ~n28364 & n28367;
  assign n28369 = ~n35898 & ~n27598;
  assign n28370 = ~n27598 & ~n27931;
  assign n28371 = ~n35898 & n28370;
  assign n28372 = ~n27931 & n28369;
  assign n28373 = n27239 & ~n36003;
  assign n28374 = n27597 & n28370;
  assign n28375 = n27239 & ~n35898;
  assign n28376 = ~n27598 & n28375;
  assign n28377 = ~n27931 & n28376;
  assign n28378 = ~n27239 & ~n36003;
  assign n28379 = ~n28377 & ~n28378;
  assign n28380 = ~n28373 & ~n28374;
  assign n28381 = ~n28368 & ~n36004;
  assign n28382 = ~n28366 & ~n28381;
  assign n28383 = ~n8506 & ~n28382;
  assign n28384 = ~n27600 & ~n27615;
  assign n28385 = ~n27931 & n28384;
  assign n28386 = ~n35900 & ~n28385;
  assign n28387 = n35900 & ~n27615;
  assign n28388 = ~n27600 & n28387;
  assign n28389 = n35900 & n28385;
  assign n28390 = ~n27931 & n28388;
  assign n28391 = ~n28386 & ~n36005;
  assign n28392 = n8506 & ~n28366;
  assign n28393 = ~n28381 & n28392;
  assign n28394 = n8506 & n28382;
  assign n28395 = ~n28391 & ~n36006;
  assign n28396 = ~n28383 & ~n28395;
  assign n28397 = ~n7975 & ~n28396;
  assign n28398 = n7975 & ~n28383;
  assign n28399 = ~n28395 & n28398;
  assign n28400 = ~n35901 & ~n27621;
  assign n28401 = ~n27621 & ~n27931;
  assign n28402 = ~n35901 & n28401;
  assign n28403 = ~n27931 & n28400;
  assign n28404 = n27231 & ~n36007;
  assign n28405 = n27620 & n28401;
  assign n28406 = n27231 & ~n35901;
  assign n28407 = ~n27621 & n28406;
  assign n28408 = ~n27931 & n28407;
  assign n28409 = ~n27231 & ~n36007;
  assign n28410 = ~n28408 & ~n28409;
  assign n28411 = ~n28404 & ~n28405;
  assign n28412 = ~n28399 & ~n36008;
  assign n28413 = ~n28397 & ~n28412;
  assign n28414 = ~n7512 & ~n28413;
  assign n28415 = n7512 & ~n28397;
  assign n28416 = ~n28412 & n28415;
  assign n28417 = n7512 & n28413;
  assign n28418 = ~n27623 & ~n27626;
  assign n28419 = ~n27626 & ~n27931;
  assign n28420 = ~n27623 & n28419;
  assign n28421 = ~n27931 & n28418;
  assign n28422 = n27223 & ~n36010;
  assign n28423 = n27624 & n28419;
  assign n28424 = n27223 & ~n27626;
  assign n28425 = ~n27623 & n28424;
  assign n28426 = ~n27931 & n28425;
  assign n28427 = ~n27223 & ~n36010;
  assign n28428 = ~n28426 & ~n28427;
  assign n28429 = ~n28422 & ~n28423;
  assign n28430 = ~n36009 & ~n36011;
  assign n28431 = ~n28414 & ~n28430;
  assign n28432 = ~n7015 & ~n28431;
  assign n28433 = n7015 & ~n28414;
  assign n28434 = ~n28430 & n28433;
  assign n28435 = ~n35902 & ~n27632;
  assign n28436 = ~n27632 & ~n27931;
  assign n28437 = ~n35902 & n28436;
  assign n28438 = ~n27931 & n28435;
  assign n28439 = n27215 & ~n36012;
  assign n28440 = n27631 & n28436;
  assign n28441 = n27215 & ~n35902;
  assign n28442 = ~n27632 & n28441;
  assign n28443 = ~n27931 & n28442;
  assign n28444 = ~n27215 & ~n36012;
  assign n28445 = ~n28443 & ~n28444;
  assign n28446 = ~n28439 & ~n28440;
  assign n28447 = ~n28434 & ~n36013;
  assign n28448 = ~n28432 & ~n28447;
  assign n28449 = ~n6579 & ~n28448;
  assign n28450 = ~n27634 & ~n27649;
  assign n28451 = ~n27931 & n28450;
  assign n28452 = ~n35904 & ~n28451;
  assign n28453 = n35904 & ~n27649;
  assign n28454 = ~n27634 & n28453;
  assign n28455 = n35904 & n28451;
  assign n28456 = ~n27931 & n28454;
  assign n28457 = ~n28452 & ~n36014;
  assign n28458 = n6579 & ~n28432;
  assign n28459 = ~n28447 & n28458;
  assign n28460 = n6579 & n28448;
  assign n28461 = ~n28457 & ~n36015;
  assign n28462 = ~n28449 & ~n28461;
  assign n28463 = ~n6117 & ~n28462;
  assign n28464 = n6117 & ~n28449;
  assign n28465 = ~n28461 & n28464;
  assign n28466 = ~n35905 & ~n27655;
  assign n28467 = ~n27655 & ~n27931;
  assign n28468 = ~n35905 & n28467;
  assign n28469 = ~n27931 & n28466;
  assign n28470 = n27207 & ~n36016;
  assign n28471 = n27654 & n28467;
  assign n28472 = n27207 & ~n35905;
  assign n28473 = ~n27655 & n28472;
  assign n28474 = ~n27931 & n28473;
  assign n28475 = ~n27207 & ~n36016;
  assign n28476 = ~n28474 & ~n28475;
  assign n28477 = ~n28470 & ~n28471;
  assign n28478 = ~n28465 & ~n36017;
  assign n28479 = ~n28463 & ~n28478;
  assign n28480 = ~n5708 & ~n28479;
  assign n28481 = n5708 & ~n28463;
  assign n28482 = ~n28478 & n28481;
  assign n28483 = n5708 & n28479;
  assign n28484 = ~n27657 & ~n27660;
  assign n28485 = ~n27660 & ~n27931;
  assign n28486 = ~n27657 & n28485;
  assign n28487 = ~n27931 & n28484;
  assign n28488 = n27199 & ~n36019;
  assign n28489 = n27658 & n28485;
  assign n28490 = n27199 & ~n27660;
  assign n28491 = ~n27657 & n28490;
  assign n28492 = ~n27931 & n28491;
  assign n28493 = ~n27199 & ~n36019;
  assign n28494 = ~n28492 & ~n28493;
  assign n28495 = ~n28488 & ~n28489;
  assign n28496 = ~n36018 & ~n36020;
  assign n28497 = ~n28480 & ~n28496;
  assign n28498 = ~n5278 & ~n28497;
  assign n28499 = n5278 & ~n28480;
  assign n28500 = ~n28496 & n28499;
  assign n28501 = ~n35906 & ~n27666;
  assign n28502 = ~n27666 & ~n27931;
  assign n28503 = ~n35906 & n28502;
  assign n28504 = ~n27931 & n28501;
  assign n28505 = n27191 & ~n36021;
  assign n28506 = n27665 & n28502;
  assign n28507 = n27191 & ~n35906;
  assign n28508 = ~n27666 & n28507;
  assign n28509 = ~n27931 & n28508;
  assign n28510 = ~n27191 & ~n36021;
  assign n28511 = ~n28509 & ~n28510;
  assign n28512 = ~n28505 & ~n28506;
  assign n28513 = ~n28500 & ~n36022;
  assign n28514 = ~n28498 & ~n28513;
  assign n28515 = ~n4903 & ~n28514;
  assign n28516 = ~n27668 & ~n27683;
  assign n28517 = ~n27931 & n28516;
  assign n28518 = ~n35908 & ~n28517;
  assign n28519 = n35908 & ~n27683;
  assign n28520 = ~n27668 & n28519;
  assign n28521 = n35908 & n28517;
  assign n28522 = ~n27931 & n28520;
  assign n28523 = ~n28518 & ~n36023;
  assign n28524 = n4903 & ~n28498;
  assign n28525 = ~n28513 & n28524;
  assign n28526 = n4903 & n28514;
  assign n28527 = ~n28523 & ~n36024;
  assign n28528 = ~n28515 & ~n28527;
  assign n28529 = ~n4508 & ~n28528;
  assign n28530 = n4508 & ~n28515;
  assign n28531 = ~n28527 & n28530;
  assign n28532 = ~n35909 & ~n27689;
  assign n28533 = ~n27689 & ~n27931;
  assign n28534 = ~n35909 & n28533;
  assign n28535 = ~n27931 & n28532;
  assign n28536 = n27183 & ~n36025;
  assign n28537 = n27688 & n28533;
  assign n28538 = n27183 & ~n35909;
  assign n28539 = ~n27689 & n28538;
  assign n28540 = ~n27931 & n28539;
  assign n28541 = ~n27183 & ~n36025;
  assign n28542 = ~n28540 & ~n28541;
  assign n28543 = ~n28536 & ~n28537;
  assign n28544 = ~n28531 & ~n36026;
  assign n28545 = ~n28529 & ~n28544;
  assign n28546 = ~n4155 & ~n28545;
  assign n28547 = n4155 & ~n28529;
  assign n28548 = ~n28544 & n28547;
  assign n28549 = n4155 & n28545;
  assign n28550 = ~n27691 & ~n27694;
  assign n28551 = ~n27694 & ~n27931;
  assign n28552 = ~n27691 & n28551;
  assign n28553 = ~n27931 & n28550;
  assign n28554 = n27175 & ~n36028;
  assign n28555 = n27692 & n28551;
  assign n28556 = n27175 & ~n27694;
  assign n28557 = ~n27691 & n28556;
  assign n28558 = ~n27931 & n28557;
  assign n28559 = ~n27175 & ~n36028;
  assign n28560 = ~n28558 & ~n28559;
  assign n28561 = ~n28554 & ~n28555;
  assign n28562 = ~n36027 & ~n36029;
  assign n28563 = ~n28546 & ~n28562;
  assign n28564 = ~n3788 & ~n28563;
  assign n28565 = n3788 & ~n28546;
  assign n28566 = ~n28562 & n28565;
  assign n28567 = ~n35910 & ~n27700;
  assign n28568 = ~n27700 & ~n27931;
  assign n28569 = ~n35910 & n28568;
  assign n28570 = ~n27931 & n28567;
  assign n28571 = n27167 & ~n36030;
  assign n28572 = n27699 & n28568;
  assign n28573 = n27167 & ~n35910;
  assign n28574 = ~n27700 & n28573;
  assign n28575 = ~n27931 & n28574;
  assign n28576 = ~n27167 & ~n36030;
  assign n28577 = ~n28575 & ~n28576;
  assign n28578 = ~n28571 & ~n28572;
  assign n28579 = ~n28566 & ~n36031;
  assign n28580 = ~n28564 & ~n28579;
  assign n28581 = ~n3473 & ~n28580;
  assign n28582 = ~n27702 & ~n27717;
  assign n28583 = ~n27931 & n28582;
  assign n28584 = ~n35912 & ~n28583;
  assign n28585 = n35912 & ~n27717;
  assign n28586 = ~n27702 & n28585;
  assign n28587 = n35912 & n28583;
  assign n28588 = ~n27931 & n28586;
  assign n28589 = ~n28584 & ~n36032;
  assign n28590 = n3473 & ~n28564;
  assign n28591 = ~n28579 & n28590;
  assign n28592 = n3473 & n28580;
  assign n28593 = ~n28589 & ~n36033;
  assign n28594 = ~n28581 & ~n28593;
  assign n28595 = ~n3140 & ~n28594;
  assign n28596 = n3140 & ~n28581;
  assign n28597 = ~n28593 & n28596;
  assign n28598 = ~n35913 & ~n27723;
  assign n28599 = ~n27723 & ~n27931;
  assign n28600 = ~n35913 & n28599;
  assign n28601 = ~n27931 & n28598;
  assign n28602 = n27159 & ~n36034;
  assign n28603 = n27722 & n28599;
  assign n28604 = n27159 & ~n35913;
  assign n28605 = ~n27723 & n28604;
  assign n28606 = ~n27931 & n28605;
  assign n28607 = ~n27159 & ~n36034;
  assign n28608 = ~n28606 & ~n28607;
  assign n28609 = ~n28602 & ~n28603;
  assign n28610 = ~n28597 & ~n36035;
  assign n28611 = ~n28595 & ~n28610;
  assign n28612 = ~n2855 & ~n28611;
  assign n28613 = n2855 & ~n28595;
  assign n28614 = ~n28610 & n28613;
  assign n28615 = n2855 & n28611;
  assign n28616 = ~n27725 & ~n27728;
  assign n28617 = ~n27728 & ~n27931;
  assign n28618 = ~n27725 & n28617;
  assign n28619 = ~n27931 & n28616;
  assign n28620 = n27151 & ~n36037;
  assign n28621 = n27726 & n28617;
  assign n28622 = n27151 & ~n27728;
  assign n28623 = ~n27725 & n28622;
  assign n28624 = ~n27931 & n28623;
  assign n28625 = ~n27151 & ~n36037;
  assign n28626 = ~n28624 & ~n28625;
  assign n28627 = ~n28620 & ~n28621;
  assign n28628 = ~n36036 & ~n36038;
  assign n28629 = ~n28612 & ~n28628;
  assign n28630 = ~n2556 & ~n28629;
  assign n28631 = n2556 & ~n28612;
  assign n28632 = ~n28628 & n28631;
  assign n28633 = ~n35914 & ~n27734;
  assign n28634 = ~n27734 & ~n27931;
  assign n28635 = ~n35914 & n28634;
  assign n28636 = ~n27931 & n28633;
  assign n28637 = n27143 & ~n36039;
  assign n28638 = n27733 & n28634;
  assign n28639 = n27143 & ~n35914;
  assign n28640 = ~n27734 & n28639;
  assign n28641 = ~n27931 & n28640;
  assign n28642 = ~n27143 & ~n36039;
  assign n28643 = ~n28641 & ~n28642;
  assign n28644 = ~n28637 & ~n28638;
  assign n28645 = ~n28632 & ~n36040;
  assign n28646 = ~n28630 & ~n28645;
  assign n28647 = ~n2301 & ~n28646;
  assign n28648 = ~n27736 & ~n27751;
  assign n28649 = ~n27931 & n28648;
  assign n28650 = ~n35916 & ~n28649;
  assign n28651 = n35916 & ~n27751;
  assign n28652 = ~n27736 & n28651;
  assign n28653 = n35916 & n28649;
  assign n28654 = ~n27931 & n28652;
  assign n28655 = ~n28650 & ~n36041;
  assign n28656 = n2301 & ~n28630;
  assign n28657 = ~n28645 & n28656;
  assign n28658 = n2301 & n28646;
  assign n28659 = ~n28655 & ~n36042;
  assign n28660 = ~n28647 & ~n28659;
  assign n28661 = ~n2038 & ~n28660;
  assign n28662 = n2038 & ~n28647;
  assign n28663 = ~n28659 & n28662;
  assign n28664 = ~n35917 & ~n27757;
  assign n28665 = ~n27757 & ~n27931;
  assign n28666 = ~n35917 & n28665;
  assign n28667 = ~n27931 & n28664;
  assign n28668 = n27135 & ~n36043;
  assign n28669 = n27756 & n28665;
  assign n28670 = n27135 & ~n35917;
  assign n28671 = ~n27757 & n28670;
  assign n28672 = ~n27931 & n28671;
  assign n28673 = ~n27135 & ~n36043;
  assign n28674 = ~n28672 & ~n28673;
  assign n28675 = ~n28668 & ~n28669;
  assign n28676 = ~n28663 & ~n36044;
  assign n28677 = ~n28661 & ~n28676;
  assign n28678 = ~n1812 & ~n28677;
  assign n28679 = n1812 & ~n28661;
  assign n28680 = ~n28676 & n28679;
  assign n28681 = n1812 & n28677;
  assign n28682 = ~n27759 & ~n27762;
  assign n28683 = ~n27762 & ~n27931;
  assign n28684 = ~n27759 & n28683;
  assign n28685 = ~n27931 & n28682;
  assign n28686 = n27127 & ~n36046;
  assign n28687 = n27760 & n28683;
  assign n28688 = n27127 & ~n27762;
  assign n28689 = ~n27759 & n28688;
  assign n28690 = ~n27931 & n28689;
  assign n28691 = ~n27127 & ~n36046;
  assign n28692 = ~n28690 & ~n28691;
  assign n28693 = ~n28686 & ~n28687;
  assign n28694 = ~n36045 & ~n36047;
  assign n28695 = ~n28678 & ~n28694;
  assign n28696 = ~n1582 & ~n28695;
  assign n28697 = n1582 & ~n28678;
  assign n28698 = ~n28694 & n28697;
  assign n28699 = ~n35918 & ~n27768;
  assign n28700 = ~n27768 & ~n27931;
  assign n28701 = ~n35918 & n28700;
  assign n28702 = ~n27931 & n28699;
  assign n28703 = n27119 & ~n36048;
  assign n28704 = n27767 & n28700;
  assign n28705 = n27119 & ~n35918;
  assign n28706 = ~n27768 & n28705;
  assign n28707 = ~n27931 & n28706;
  assign n28708 = ~n27119 & ~n36048;
  assign n28709 = ~n28707 & ~n28708;
  assign n28710 = ~n28703 & ~n28704;
  assign n28711 = ~n28698 & ~n36049;
  assign n28712 = ~n28696 & ~n28711;
  assign n28713 = ~n1388 & ~n28712;
  assign n28714 = ~n27770 & ~n27785;
  assign n28715 = ~n27931 & n28714;
  assign n28716 = ~n35920 & ~n28715;
  assign n28717 = n35920 & ~n27785;
  assign n28718 = ~n27770 & n28717;
  assign n28719 = n35920 & n28715;
  assign n28720 = ~n27931 & n28718;
  assign n28721 = ~n28716 & ~n36050;
  assign n28722 = n1388 & ~n28696;
  assign n28723 = ~n28711 & n28722;
  assign n28724 = n1388 & n28712;
  assign n28725 = ~n28721 & ~n36051;
  assign n28726 = ~n28713 & ~n28725;
  assign n28727 = ~n1192 & ~n28726;
  assign n28728 = n1192 & ~n28713;
  assign n28729 = ~n28725 & n28728;
  assign n28730 = ~n35921 & ~n27791;
  assign n28731 = ~n27791 & ~n27931;
  assign n28732 = ~n35921 & n28731;
  assign n28733 = ~n27931 & n28730;
  assign n28734 = n27111 & ~n36052;
  assign n28735 = n27790 & n28731;
  assign n28736 = n27111 & ~n35921;
  assign n28737 = ~n27791 & n28736;
  assign n28738 = ~n27931 & n28737;
  assign n28739 = ~n27111 & ~n36052;
  assign n28740 = ~n28738 & ~n28739;
  assign n28741 = ~n28734 & ~n28735;
  assign n28742 = ~n28729 & ~n36053;
  assign n28743 = ~n28727 & ~n28742;
  assign n28744 = ~n1028 & ~n28743;
  assign n28745 = n1028 & ~n28727;
  assign n28746 = ~n28742 & n28745;
  assign n28747 = n1028 & n28743;
  assign n28748 = ~n27793 & ~n27796;
  assign n28749 = ~n27796 & ~n27931;
  assign n28750 = ~n27793 & n28749;
  assign n28751 = ~n27931 & n28748;
  assign n28752 = n27103 & ~n36055;
  assign n28753 = n27794 & n28749;
  assign n28754 = n27103 & ~n27796;
  assign n28755 = ~n27793 & n28754;
  assign n28756 = ~n27931 & n28755;
  assign n28757 = ~n27103 & ~n36055;
  assign n28758 = ~n28756 & ~n28757;
  assign n28759 = ~n28752 & ~n28753;
  assign n28760 = ~n36054 & ~n36056;
  assign n28761 = ~n28744 & ~n28760;
  assign n28762 = ~n866 & ~n28761;
  assign n28763 = n866 & ~n28744;
  assign n28764 = ~n28760 & n28763;
  assign n28765 = ~n35922 & ~n27802;
  assign n28766 = ~n27802 & ~n27931;
  assign n28767 = ~n35922 & n28766;
  assign n28768 = ~n27931 & n28765;
  assign n28769 = n27095 & ~n36057;
  assign n28770 = n27801 & n28766;
  assign n28771 = n27095 & ~n35922;
  assign n28772 = ~n27802 & n28771;
  assign n28773 = ~n27931 & n28772;
  assign n28774 = ~n27095 & ~n36057;
  assign n28775 = ~n28773 & ~n28774;
  assign n28776 = ~n28769 & ~n28770;
  assign n28777 = ~n28764 & ~n36058;
  assign n28778 = ~n28762 & ~n28777;
  assign n28779 = ~n730 & ~n28778;
  assign n28780 = ~n27804 & ~n27819;
  assign n28781 = ~n27931 & n28780;
  assign n28782 = ~n35924 & ~n28781;
  assign n28783 = n35924 & ~n27819;
  assign n28784 = ~n27804 & n28783;
  assign n28785 = n35924 & n28781;
  assign n28786 = ~n27931 & n28784;
  assign n28787 = ~n28782 & ~n36059;
  assign n28788 = n730 & ~n28762;
  assign n28789 = ~n28777 & n28788;
  assign n28790 = n730 & n28778;
  assign n28791 = ~n28787 & ~n36060;
  assign n28792 = ~n28779 & ~n28791;
  assign n28793 = ~n602 & ~n28792;
  assign n28794 = n602 & ~n28779;
  assign n28795 = ~n28791 & n28794;
  assign n28796 = ~n35925 & ~n27825;
  assign n28797 = ~n27825 & ~n27931;
  assign n28798 = ~n35925 & n28797;
  assign n28799 = ~n27931 & n28796;
  assign n28800 = n27087 & ~n36061;
  assign n28801 = n27824 & n28797;
  assign n28802 = n27087 & ~n35925;
  assign n28803 = ~n27825 & n28802;
  assign n28804 = ~n27931 & n28803;
  assign n28805 = ~n27087 & ~n36061;
  assign n28806 = ~n28804 & ~n28805;
  assign n28807 = ~n28800 & ~n28801;
  assign n28808 = ~n28795 & ~n36062;
  assign n28809 = ~n28793 & ~n28808;
  assign n28810 = ~n497 & ~n28809;
  assign n28811 = n497 & ~n28793;
  assign n28812 = ~n28808 & n28811;
  assign n28813 = n497 & n28809;
  assign n28814 = ~n27827 & ~n27830;
  assign n28815 = ~n27830 & ~n27931;
  assign n28816 = ~n27827 & n28815;
  assign n28817 = ~n27931 & n28814;
  assign n28818 = n27079 & ~n36064;
  assign n28819 = n27828 & n28815;
  assign n28820 = n27079 & ~n27830;
  assign n28821 = ~n27827 & n28820;
  assign n28822 = ~n27931 & n28821;
  assign n28823 = ~n27079 & ~n36064;
  assign n28824 = ~n28822 & ~n28823;
  assign n28825 = ~n28818 & ~n28819;
  assign n28826 = ~n36063 & ~n36065;
  assign n28827 = ~n28810 & ~n28826;
  assign n28828 = ~n403 & ~n28827;
  assign n28829 = n403 & ~n28810;
  assign n28830 = ~n28826 & n28829;
  assign n28831 = n27071 & ~n35926;
  assign n28832 = ~n27836 & n28831;
  assign n28833 = ~n35926 & ~n27836;
  assign n28834 = ~n27931 & n28833;
  assign n28835 = n27071 & n28834;
  assign n28836 = ~n27931 & n28832;
  assign n28837 = ~n27071 & ~n28834;
  assign n28838 = ~n36066 & ~n28837;
  assign n28839 = ~n28830 & ~n28838;
  assign n28840 = ~n28828 & ~n28839;
  assign n28841 = ~n330 & ~n28840;
  assign n28842 = n330 & ~n28828;
  assign n28843 = ~n28839 & n28842;
  assign n28844 = n330 & n28840;
  assign n28845 = ~n27838 & ~n27840;
  assign n28846 = ~n27931 & n28845;
  assign n28847 = ~n35928 & n28846;
  assign n28848 = n35928 & ~n28846;
  assign n28849 = ~n27838 & n35928;
  assign n28850 = ~n27840 & n28849;
  assign n28851 = n35928 & n28846;
  assign n28852 = ~n27931 & n28850;
  assign n28853 = ~n35928 & ~n28846;
  assign n28854 = ~n36068 & ~n28853;
  assign n28855 = ~n28847 & ~n28848;
  assign n28856 = ~n36067 & ~n36069;
  assign n28857 = ~n28841 & ~n28856;
  assign n28858 = ~n271 & ~n28857;
  assign n28859 = n271 & ~n28841;
  assign n28860 = ~n28856 & n28859;
  assign n28861 = ~n35940 & ~n28860;
  assign n28862 = ~n28858 & ~n28861;
  assign n28863 = ~n217 & ~n28862;
  assign n28864 = ~n27860 & ~n27862;
  assign n28865 = ~n27931 & n28864;
  assign n28866 = ~n35931 & ~n28865;
  assign n28867 = ~n27860 & n35931;
  assign n28868 = ~n27862 & n28867;
  assign n28869 = n35931 & n28865;
  assign n28870 = ~n27931 & n28868;
  assign n28871 = ~n28866 & ~n36070;
  assign n28872 = n217 & ~n28858;
  assign n28873 = ~n28861 & n28872;
  assign n28874 = n217 & n28862;
  assign n28875 = ~n28871 & ~n36071;
  assign n28876 = ~n28863 & ~n28875;
  assign n28877 = ~n198 & ~n28876;
  assign n28878 = n198 & ~n28863;
  assign n28879 = ~n28875 & n28878;
  assign n28880 = ~n27877 & ~n35933;
  assign n28881 = ~n27877 & ~n27931;
  assign n28882 = ~n35933 & n28881;
  assign n28883 = ~n27931 & n28880;
  assign n28884 = n27885 & ~n36072;
  assign n28885 = n27889 & n28881;
  assign n28886 = n27885 & ~n35933;
  assign n28887 = ~n27877 & n28886;
  assign n28888 = ~n27931 & n28887;
  assign n28889 = ~n27885 & ~n36072;
  assign n28890 = ~n28888 & ~n28889;
  assign n28891 = ~n28884 & ~n28885;
  assign n28892 = ~n28879 & ~n36073;
  assign n28893 = ~n28877 & ~n28892;
  assign n28894 = ~n27891 & ~n27893;
  assign n28895 = ~n27931 & n28894;
  assign n28896 = ~n35935 & ~n28895;
  assign n28897 = ~n27891 & n35935;
  assign n28898 = ~n27893 & n28897;
  assign n28899 = n35935 & n28895;
  assign n28900 = ~n27931 & n28898;
  assign n28901 = ~n28896 & ~n36074;
  assign n28902 = ~n27907 & ~n27915;
  assign n28903 = ~n27915 & ~n27931;
  assign n28904 = ~n27907 & n28903;
  assign n28905 = ~n27931 & n28902;
  assign n28906 = ~n35938 & ~n36075;
  assign n28907 = ~n28901 & n28906;
  assign n28908 = ~n28893 & n28907;
  assign n28909 = n193 & ~n28908;
  assign n28910 = ~n28877 & n28901;
  assign n28911 = ~n28892 & n28910;
  assign n28912 = n28893 & n28901;
  assign n28913 = n27907 & ~n28903;
  assign n28914 = ~n193 & ~n28902;
  assign n28915 = ~n28913 & n28914;
  assign n28916 = ~n36076 & ~n28915;
  assign n28917 = ~n28909 & n28916;
  assign n28918 = ~n28858 & ~n28860;
  assign n28919 = ~n28917 & n28918;
  assign n28920 = ~n35940 & ~n28919;
  assign n28921 = n35940 & ~n28860;
  assign n28922 = ~n28858 & n28921;
  assign n28923 = n35940 & n28919;
  assign n28924 = ~n28917 & n28922;
  assign n28925 = ~n28920 & ~n36077;
  assign n28926 = ~n28828 & ~n28830;
  assign n28927 = ~n28917 & n28926;
  assign n28928 = ~n28838 & ~n28927;
  assign n28929 = ~n28830 & n28838;
  assign n28930 = ~n28828 & n28929;
  assign n28931 = n28838 & n28927;
  assign n28932 = ~n28917 & n28930;
  assign n28933 = ~n28928 & ~n36078;
  assign n28934 = ~n28810 & ~n36063;
  assign n28935 = ~n28917 & n28934;
  assign n28936 = ~n36065 & ~n28935;
  assign n28937 = ~n28810 & n36065;
  assign n28938 = ~n36063 & n28937;
  assign n28939 = n36065 & n28935;
  assign n28940 = ~n28917 & n28938;
  assign n28941 = ~n28936 & ~n36079;
  assign n28942 = ~n28793 & ~n28795;
  assign n28943 = ~n28917 & n28942;
  assign n28944 = ~n36062 & ~n28943;
  assign n28945 = ~n28795 & n36062;
  assign n28946 = ~n28793 & n28945;
  assign n28947 = n36062 & n28943;
  assign n28948 = ~n28917 & n28946;
  assign n28949 = ~n28944 & ~n36080;
  assign n28950 = ~n28762 & ~n28764;
  assign n28951 = ~n28917 & n28950;
  assign n28952 = ~n36058 & ~n28951;
  assign n28953 = ~n28764 & n36058;
  assign n28954 = ~n28762 & n28953;
  assign n28955 = n36058 & n28951;
  assign n28956 = ~n28917 & n28954;
  assign n28957 = ~n28952 & ~n36081;
  assign n28958 = ~n28744 & ~n36054;
  assign n28959 = ~n28917 & n28958;
  assign n28960 = ~n36056 & ~n28959;
  assign n28961 = ~n28744 & n36056;
  assign n28962 = ~n36054 & n28961;
  assign n28963 = n36056 & n28959;
  assign n28964 = ~n28917 & n28962;
  assign n28965 = ~n28960 & ~n36082;
  assign n28966 = ~n28727 & ~n28729;
  assign n28967 = ~n28917 & n28966;
  assign n28968 = ~n36053 & ~n28967;
  assign n28969 = ~n28729 & n36053;
  assign n28970 = ~n28727 & n28969;
  assign n28971 = n36053 & n28967;
  assign n28972 = ~n28917 & n28970;
  assign n28973 = ~n28968 & ~n36083;
  assign n28974 = ~n28696 & ~n28698;
  assign n28975 = ~n28917 & n28974;
  assign n28976 = ~n36049 & ~n28975;
  assign n28977 = ~n28698 & n36049;
  assign n28978 = ~n28696 & n28977;
  assign n28979 = n36049 & n28975;
  assign n28980 = ~n28917 & n28978;
  assign n28981 = ~n28976 & ~n36084;
  assign n28982 = ~n28678 & ~n36045;
  assign n28983 = ~n28917 & n28982;
  assign n28984 = ~n36047 & ~n28983;
  assign n28985 = ~n28678 & n36047;
  assign n28986 = ~n36045 & n28985;
  assign n28987 = n36047 & n28983;
  assign n28988 = ~n28917 & n28986;
  assign n28989 = ~n28984 & ~n36085;
  assign n28990 = ~n28661 & ~n28663;
  assign n28991 = ~n28917 & n28990;
  assign n28992 = ~n36044 & ~n28991;
  assign n28993 = ~n28663 & n36044;
  assign n28994 = ~n28661 & n28993;
  assign n28995 = n36044 & n28991;
  assign n28996 = ~n28917 & n28994;
  assign n28997 = ~n28992 & ~n36086;
  assign n28998 = ~n28630 & ~n28632;
  assign n28999 = ~n28917 & n28998;
  assign n29000 = ~n36040 & ~n28999;
  assign n29001 = ~n28632 & n36040;
  assign n29002 = ~n28630 & n29001;
  assign n29003 = n36040 & n28999;
  assign n29004 = ~n28917 & n29002;
  assign n29005 = ~n29000 & ~n36087;
  assign n29006 = ~n28612 & ~n36036;
  assign n29007 = ~n28917 & n29006;
  assign n29008 = ~n36038 & ~n29007;
  assign n29009 = ~n28612 & n36038;
  assign n29010 = ~n36036 & n29009;
  assign n29011 = n36038 & n29007;
  assign n29012 = ~n28917 & n29010;
  assign n29013 = ~n29008 & ~n36088;
  assign n29014 = ~n28595 & ~n28597;
  assign n29015 = ~n28917 & n29014;
  assign n29016 = ~n36035 & ~n29015;
  assign n29017 = ~n28597 & n36035;
  assign n29018 = ~n28595 & n29017;
  assign n29019 = n36035 & n29015;
  assign n29020 = ~n28917 & n29018;
  assign n29021 = ~n29016 & ~n36089;
  assign n29022 = ~n28564 & ~n28566;
  assign n29023 = ~n28917 & n29022;
  assign n29024 = ~n36031 & ~n29023;
  assign n29025 = ~n28566 & n36031;
  assign n29026 = ~n28564 & n29025;
  assign n29027 = n36031 & n29023;
  assign n29028 = ~n28917 & n29026;
  assign n29029 = ~n29024 & ~n36090;
  assign n29030 = ~n28546 & ~n36027;
  assign n29031 = ~n28917 & n29030;
  assign n29032 = ~n36029 & ~n29031;
  assign n29033 = ~n28546 & n36029;
  assign n29034 = ~n36027 & n29033;
  assign n29035 = n36029 & n29031;
  assign n29036 = ~n28917 & n29034;
  assign n29037 = ~n29032 & ~n36091;
  assign n29038 = ~n28529 & ~n28531;
  assign n29039 = ~n28917 & n29038;
  assign n29040 = ~n36026 & ~n29039;
  assign n29041 = ~n28531 & n36026;
  assign n29042 = ~n28529 & n29041;
  assign n29043 = n36026 & n29039;
  assign n29044 = ~n28917 & n29042;
  assign n29045 = ~n29040 & ~n36092;
  assign n29046 = ~n28498 & ~n28500;
  assign n29047 = ~n28917 & n29046;
  assign n29048 = ~n36022 & ~n29047;
  assign n29049 = ~n28500 & n36022;
  assign n29050 = ~n28498 & n29049;
  assign n29051 = n36022 & n29047;
  assign n29052 = ~n28917 & n29050;
  assign n29053 = ~n29048 & ~n36093;
  assign n29054 = ~n28480 & ~n36018;
  assign n29055 = ~n28917 & n29054;
  assign n29056 = ~n36020 & ~n29055;
  assign n29057 = ~n28480 & n36020;
  assign n29058 = ~n36018 & n29057;
  assign n29059 = n36020 & n29055;
  assign n29060 = ~n28917 & n29058;
  assign n29061 = ~n29056 & ~n36094;
  assign n29062 = ~n28463 & ~n28465;
  assign n29063 = ~n28917 & n29062;
  assign n29064 = ~n36017 & ~n29063;
  assign n29065 = ~n28465 & n36017;
  assign n29066 = ~n28463 & n29065;
  assign n29067 = n36017 & n29063;
  assign n29068 = ~n28917 & n29066;
  assign n29069 = ~n29064 & ~n36095;
  assign n29070 = ~n28432 & ~n28434;
  assign n29071 = ~n28917 & n29070;
  assign n29072 = ~n36013 & ~n29071;
  assign n29073 = ~n28434 & n36013;
  assign n29074 = ~n28432 & n29073;
  assign n29075 = n36013 & n29071;
  assign n29076 = ~n28917 & n29074;
  assign n29077 = ~n29072 & ~n36096;
  assign n29078 = ~n28414 & ~n36009;
  assign n29079 = ~n28917 & n29078;
  assign n29080 = ~n36011 & ~n29079;
  assign n29081 = ~n28414 & n36011;
  assign n29082 = ~n36009 & n29081;
  assign n29083 = n36011 & n29079;
  assign n29084 = ~n28917 & n29082;
  assign n29085 = ~n29080 & ~n36097;
  assign n29086 = ~n28397 & ~n28399;
  assign n29087 = ~n28917 & n29086;
  assign n29088 = ~n36008 & ~n29087;
  assign n29089 = ~n28399 & n36008;
  assign n29090 = ~n28397 & n29089;
  assign n29091 = n36008 & n29087;
  assign n29092 = ~n28917 & n29090;
  assign n29093 = ~n29088 & ~n36098;
  assign n29094 = ~n28366 & ~n28368;
  assign n29095 = ~n28917 & n29094;
  assign n29096 = ~n36004 & ~n29095;
  assign n29097 = ~n28368 & n36004;
  assign n29098 = ~n28366 & n29097;
  assign n29099 = n36004 & n29095;
  assign n29100 = ~n28917 & n29098;
  assign n29101 = ~n29096 & ~n36099;
  assign n29102 = ~n28348 & ~n36000;
  assign n29103 = ~n28917 & n29102;
  assign n29104 = ~n36002 & ~n29103;
  assign n29105 = ~n28348 & n36002;
  assign n29106 = ~n36000 & n29105;
  assign n29107 = n36002 & n29103;
  assign n29108 = ~n28917 & n29106;
  assign n29109 = ~n29104 & ~n36100;
  assign n29110 = ~n28331 & ~n28333;
  assign n29111 = ~n28917 & n29110;
  assign n29112 = ~n35999 & ~n29111;
  assign n29113 = ~n28333 & n35999;
  assign n29114 = ~n28331 & n29113;
  assign n29115 = n35999 & n29111;
  assign n29116 = ~n28917 & n29114;
  assign n29117 = ~n29112 & ~n36101;
  assign n29118 = ~n28300 & ~n28302;
  assign n29119 = ~n28917 & n29118;
  assign n29120 = ~n35995 & ~n29119;
  assign n29121 = ~n28302 & n35995;
  assign n29122 = ~n28300 & n29121;
  assign n29123 = n35995 & n29119;
  assign n29124 = ~n28917 & n29122;
  assign n29125 = ~n29120 & ~n36102;
  assign n29126 = ~n28281 & ~n35990;
  assign n29127 = ~n28917 & n29126;
  assign n29128 = ~n35993 & ~n29127;
  assign n29129 = ~n28281 & n35993;
  assign n29130 = ~n35990 & n29129;
  assign n29131 = n35993 & n29127;
  assign n29132 = ~n28917 & n29130;
  assign n29133 = ~n29128 & ~n36103;
  assign n29134 = ~n28264 & ~n28266;
  assign n29135 = ~n28917 & n29134;
  assign n29136 = ~n35989 & ~n29135;
  assign n29137 = ~n28266 & n35989;
  assign n29138 = ~n28264 & n29137;
  assign n29139 = n35989 & n29135;
  assign n29140 = ~n28917 & n29138;
  assign n29141 = ~n29136 & ~n36104;
  assign n29142 = ~n28230 & ~n28232;
  assign n29143 = ~n28917 & n29142;
  assign n29144 = ~n35984 & ~n29143;
  assign n29145 = ~n28232 & n35984;
  assign n29146 = ~n28230 & n29145;
  assign n29147 = n35984 & n29143;
  assign n29148 = ~n28917 & n29146;
  assign n29149 = ~n29144 & ~n36105;
  assign n29150 = ~n28194 & ~n28196;
  assign n29151 = ~n28917 & n29150;
  assign n29152 = ~n35978 & ~n29151;
  assign n29153 = ~n28196 & n35978;
  assign n29154 = ~n28194 & n29153;
  assign n29155 = n35978 & n29151;
  assign n29156 = ~n28917 & n29154;
  assign n29157 = ~n29152 & ~n36106;
  assign n29158 = ~n28163 & ~n28165;
  assign n29159 = ~n28917 & n29158;
  assign n29160 = ~n35974 & ~n29159;
  assign n29161 = ~n28165 & n35974;
  assign n29162 = ~n28163 & n29161;
  assign n29163 = n35974 & n29159;
  assign n29164 = ~n28917 & n29162;
  assign n29165 = ~n29160 & ~n36107;
  assign n29166 = ~n28127 & ~n28129;
  assign n29167 = ~n28917 & n29166;
  assign n29168 = ~n35968 & ~n29167;
  assign n29169 = ~n28129 & n35968;
  assign n29170 = ~n28127 & n29169;
  assign n29171 = n35968 & n29167;
  assign n29172 = ~n28917 & n29170;
  assign n29173 = ~n29168 & ~n36108;
  assign n29174 = ~n28093 & ~n28095;
  assign n29175 = ~n28917 & n29174;
  assign n29176 = ~n35963 & ~n29175;
  assign n29177 = ~n28095 & n35963;
  assign n29178 = ~n28093 & n29177;
  assign n29179 = n35963 & n29175;
  assign n29180 = ~n28917 & n29178;
  assign n29181 = ~n29176 & ~n36109;
  assign n29182 = ~n28059 & ~n28061;
  assign n29183 = ~n28917 & n29182;
  assign n29184 = ~n35958 & ~n29183;
  assign n29185 = ~n28061 & n35958;
  assign n29186 = ~n28059 & n29185;
  assign n29187 = n35958 & n29183;
  assign n29188 = ~n28917 & n29186;
  assign n29189 = ~n29184 & ~n36110;
  assign n29190 = ~n28026 & ~n28028;
  assign n29191 = ~n28917 & n29190;
  assign n29192 = ~n35954 & ~n29191;
  assign n29193 = ~n28028 & n35954;
  assign n29194 = ~n28026 & n29193;
  assign n29195 = n35954 & n29191;
  assign n29196 = ~n28917 & n29194;
  assign n29197 = ~n29192 & ~n36111;
  assign n29198 = ~n27992 & ~n27994;
  assign n29199 = ~n28917 & n29198;
  assign n29200 = ~n35949 & ~n29199;
  assign n29201 = ~n27994 & n35949;
  assign n29202 = ~n27992 & n29201;
  assign n29203 = n35949 & n29199;
  assign n29204 = ~n28917 & n29202;
  assign n29205 = ~n29200 & ~n36112;
  assign n29206 = ~n27964 & ~n27966;
  assign n29207 = ~n28917 & n29206;
  assign n29208 = ~n27976 & ~n29207;
  assign n29209 = ~n27966 & n27976;
  assign n29210 = ~n27964 & n29209;
  assign n29211 = n27976 & n29207;
  assign n29212 = ~n28917 & n29210;
  assign n29213 = ~n29208 & ~n36113;
  assign n29214 = ~pi6  & ~n28917;
  assign n29215 = ~pi7  & n29214;
  assign n29216 = n27945 & ~n28917;
  assign n29217 = ~n27931 & ~n28915;
  assign n29218 = ~n36076 & n29217;
  assign n29219 = ~n27931 & n28917;
  assign n29220 = ~n28909 & n29218;
  assign n29221 = ~n36114 & ~n36115;
  assign n29222 = pi8  & ~n29221;
  assign n29223 = ~pi8  & ~n36115;
  assign n29224 = ~pi8  & n29221;
  assign n29225 = ~n36114 & n29223;
  assign n29226 = ~n29222 & ~n36116;
  assign n29227 = pi6  & ~n28917;
  assign n29228 = ~pi4  & ~pi5 ;
  assign n29229 = ~pi6  & n29228;
  assign n29230 = ~n27929 & ~n29229;
  assign n29231 = ~n35938 & n29230;
  assign n29232 = ~n27923 & n29231;
  assign n29233 = ~pi6  & ~n29228;
  assign n29234 = pi6  & n28917;
  assign n29235 = ~n29233 & ~n29234;
  assign n29236 = ~n29227 & ~n29229;
  assign n29237 = n27931 & ~n36117;
  assign n29238 = ~n29227 & n29232;
  assign n29239 = pi7  & ~n29214;
  assign n29240 = ~n36114 & ~n29239;
  assign n29241 = ~n36118 & n29240;
  assign n29242 = ~n27931 & n36117;
  assign n29243 = n27055 & ~n29242;
  assign n29244 = ~n29241 & ~n29242;
  assign n29245 = n27055 & n29244;
  assign n29246 = ~n29241 & n29243;
  assign n29247 = ~n29226 & ~n36119;
  assign n29248 = ~n27055 & ~n29244;
  assign n29249 = n26098 & ~n29248;
  assign n29250 = ~n29247 & n29249;
  assign n29251 = ~n27951 & ~n35943;
  assign n29252 = ~n28917 & n29251;
  assign n29253 = n27956 & ~n29252;
  assign n29254 = ~n27956 & n29251;
  assign n29255 = ~n27956 & n29252;
  assign n29256 = ~n28917 & n29254;
  assign n29257 = ~n29253 & ~n36120;
  assign n29258 = ~n29250 & ~n29257;
  assign n29259 = ~n29247 & ~n29248;
  assign n29260 = ~n26098 & ~n29259;
  assign n29261 = n25256 & ~n29260;
  assign n29262 = ~n29258 & ~n29260;
  assign n29263 = n25256 & n29262;
  assign n29264 = ~n29258 & n29261;
  assign n29265 = ~n29213 & ~n36121;
  assign n29266 = ~n25256 & ~n29262;
  assign n29267 = n24331 & ~n29266;
  assign n29268 = ~n29265 & n29267;
  assign n29269 = ~n27979 & ~n35946;
  assign n29270 = ~n28917 & n29269;
  assign n29271 = n27989 & ~n29270;
  assign n29272 = ~n27989 & n29270;
  assign n29273 = ~n27979 & n27989;
  assign n29274 = ~n35946 & n29273;
  assign n29275 = n27989 & n29270;
  assign n29276 = ~n28917 & n29274;
  assign n29277 = ~n27989 & ~n29270;
  assign n29278 = ~n36122 & ~n29277;
  assign n29279 = ~n29271 & ~n29272;
  assign n29280 = ~n29268 & ~n36123;
  assign n29281 = ~n29265 & ~n29266;
  assign n29282 = ~n24331 & ~n29281;
  assign n29283 = n23517 & ~n29282;
  assign n29284 = ~n29280 & ~n29282;
  assign n29285 = n23517 & n29284;
  assign n29286 = ~n29280 & n29283;
  assign n29287 = ~n29205 & ~n36124;
  assign n29288 = ~n23517 & ~n29284;
  assign n29289 = n22625 & ~n29288;
  assign n29290 = ~n29287 & n29289;
  assign n29291 = ~n28009 & ~n35950;
  assign n29292 = ~n28917 & n29291;
  assign n29293 = ~n35952 & n29292;
  assign n29294 = n35952 & ~n29292;
  assign n29295 = ~n28009 & n35952;
  assign n29296 = ~n35950 & n29295;
  assign n29297 = ~n28917 & n29296;
  assign n29298 = ~n35952 & ~n29292;
  assign n29299 = ~n29297 & ~n29298;
  assign n29300 = ~n29293 & ~n29294;
  assign n29301 = ~n29290 & ~n36125;
  assign n29302 = ~n29287 & ~n29288;
  assign n29303 = ~n22625 & ~n29302;
  assign n29304 = n21842 & ~n29303;
  assign n29305 = ~n29301 & ~n29303;
  assign n29306 = n21842 & n29305;
  assign n29307 = ~n29301 & n29304;
  assign n29308 = ~n29197 & ~n36126;
  assign n29309 = ~n21842 & ~n29305;
  assign n29310 = n20986 & ~n29309;
  assign n29311 = ~n29308 & n29310;
  assign n29312 = ~n28043 & ~n35955;
  assign n29313 = ~n28917 & n29312;
  assign n29314 = ~n35956 & ~n29313;
  assign n29315 = ~n28043 & n35956;
  assign n29316 = ~n35955 & n29315;
  assign n29317 = n35956 & n29313;
  assign n29318 = ~n28917 & n29316;
  assign n29319 = n35956 & ~n29313;
  assign n29320 = ~n35956 & n29313;
  assign n29321 = ~n29319 & ~n29320;
  assign n29322 = ~n29314 & ~n36127;
  assign n29323 = ~n29311 & n36128;
  assign n29324 = ~n29308 & ~n29309;
  assign n29325 = ~n20986 & ~n29324;
  assign n29326 = n20229 & ~n29325;
  assign n29327 = ~n29323 & ~n29325;
  assign n29328 = n20229 & n29327;
  assign n29329 = ~n29323 & n29326;
  assign n29330 = ~n29189 & ~n36129;
  assign n29331 = ~n20229 & ~n29327;
  assign n29332 = n19401 & ~n29331;
  assign n29333 = ~n29330 & n29332;
  assign n29334 = ~n28076 & ~n35959;
  assign n29335 = ~n28917 & n29334;
  assign n29336 = n35961 & ~n29335;
  assign n29337 = ~n28076 & ~n35961;
  assign n29338 = ~n35959 & n29337;
  assign n29339 = ~n35961 & n29335;
  assign n29340 = ~n28917 & n29338;
  assign n29341 = n35961 & n29335;
  assign n29342 = ~n35961 & ~n29335;
  assign n29343 = ~n29341 & ~n29342;
  assign n29344 = ~n29336 & ~n36130;
  assign n29345 = ~n29333 & n36131;
  assign n29346 = ~n29330 & ~n29331;
  assign n29347 = ~n19401 & ~n29346;
  assign n29348 = n18676 & ~n29347;
  assign n29349 = ~n29345 & ~n29347;
  assign n29350 = n18676 & n29349;
  assign n29351 = ~n29345 & n29348;
  assign n29352 = ~n29181 & ~n36132;
  assign n29353 = ~n18676 & ~n29349;
  assign n29354 = n17885 & ~n29353;
  assign n29355 = ~n29352 & n29354;
  assign n29356 = ~n28110 & ~n35964;
  assign n29357 = ~n28110 & ~n28917;
  assign n29358 = ~n35964 & n29357;
  assign n29359 = ~n28917 & n29356;
  assign n29360 = ~n35966 & ~n36133;
  assign n29361 = n28125 & n29357;
  assign n29362 = n35966 & n36133;
  assign n29363 = ~n28110 & ~n35966;
  assign n29364 = ~n35964 & n29363;
  assign n29365 = ~n28917 & n29364;
  assign n29366 = n35966 & ~n36133;
  assign n29367 = ~n29365 & ~n29366;
  assign n29368 = ~n29360 & ~n36134;
  assign n29369 = ~n29355 & ~n36135;
  assign n29370 = ~n29352 & ~n29353;
  assign n29371 = ~n17885 & ~n29370;
  assign n29372 = n17187 & ~n29371;
  assign n29373 = ~n29369 & ~n29371;
  assign n29374 = n17187 & n29373;
  assign n29375 = ~n29369 & n29372;
  assign n29376 = ~n29173 & ~n36136;
  assign n29377 = ~n17187 & ~n29373;
  assign n29378 = n16428 & ~n29377;
  assign n29379 = ~n29376 & n29378;
  assign n29380 = ~n28144 & ~n35969;
  assign n29381 = ~n28917 & n29380;
  assign n29382 = ~n35972 & ~n29381;
  assign n29383 = ~n28144 & n35972;
  assign n29384 = ~n35969 & n29383;
  assign n29385 = n35972 & n29381;
  assign n29386 = ~n28917 & n29384;
  assign n29387 = ~n29382 & ~n36137;
  assign n29388 = ~n29379 & ~n29387;
  assign n29389 = ~n29376 & ~n29377;
  assign n29390 = ~n16428 & ~n29389;
  assign n29391 = n15760 & ~n29390;
  assign n29392 = ~n29388 & ~n29390;
  assign n29393 = n15760 & n29392;
  assign n29394 = ~n29388 & n29391;
  assign n29395 = ~n29165 & ~n36138;
  assign n29396 = ~n15760 & ~n29392;
  assign n29397 = n15033 & ~n29396;
  assign n29398 = ~n29395 & n29397;
  assign n29399 = ~n28180 & ~n35975;
  assign n29400 = ~n28180 & ~n28917;
  assign n29401 = ~n35975 & n29400;
  assign n29402 = ~n28917 & n29399;
  assign n29403 = n28191 & ~n36139;
  assign n29404 = n28192 & n29400;
  assign n29405 = ~n28191 & n36139;
  assign n29406 = ~n28180 & n28191;
  assign n29407 = ~n35975 & n29406;
  assign n29408 = ~n28917 & n29407;
  assign n29409 = ~n28191 & ~n36139;
  assign n29410 = ~n29408 & ~n29409;
  assign n29411 = ~n29403 & ~n36140;
  assign n29412 = ~n29398 & ~n36141;
  assign n29413 = ~n29395 & ~n29396;
  assign n29414 = ~n15033 & ~n29413;
  assign n29415 = n14394 & ~n29414;
  assign n29416 = ~n29412 & ~n29414;
  assign n29417 = n14394 & n29416;
  assign n29418 = ~n29412 & n29415;
  assign n29419 = ~n29157 & ~n36142;
  assign n29420 = ~n14394 & ~n29416;
  assign n29421 = n13704 & ~n29420;
  assign n29422 = ~n29419 & n29421;
  assign n29423 = ~n28211 & ~n35979;
  assign n29424 = ~n28917 & n29423;
  assign n29425 = ~n35982 & n29424;
  assign n29426 = n35982 & ~n29424;
  assign n29427 = ~n28211 & n35982;
  assign n29428 = ~n35979 & n29427;
  assign n29429 = n35982 & n29424;
  assign n29430 = ~n28917 & n29428;
  assign n29431 = ~n35982 & ~n29424;
  assign n29432 = ~n36143 & ~n29431;
  assign n29433 = ~n29425 & ~n29426;
  assign n29434 = ~n29422 & ~n36144;
  assign n29435 = ~n29419 & ~n29420;
  assign n29436 = ~n13704 & ~n29435;
  assign n29437 = n13099 & ~n29436;
  assign n29438 = ~n29434 & ~n29436;
  assign n29439 = n13099 & n29438;
  assign n29440 = ~n29434 & n29437;
  assign n29441 = ~n29149 & ~n36145;
  assign n29442 = ~n13099 & ~n29438;
  assign n29443 = n12442 & ~n29442;
  assign n29444 = ~n29441 & n29443;
  assign n29445 = ~n28247 & ~n35985;
  assign n29446 = ~n28247 & ~n28917;
  assign n29447 = ~n35985 & n29446;
  assign n29448 = ~n28917 & n29445;
  assign n29449 = n35987 & ~n36146;
  assign n29450 = n28262 & n29446;
  assign n29451 = ~n35987 & n36146;
  assign n29452 = ~n28247 & n35987;
  assign n29453 = ~n35985 & n29452;
  assign n29454 = ~n28917 & n29453;
  assign n29455 = ~n35987 & ~n36146;
  assign n29456 = ~n29454 & ~n29455;
  assign n29457 = ~n29449 & ~n36147;
  assign n29458 = ~n29444 & ~n36148;
  assign n29459 = ~n29441 & ~n29442;
  assign n29460 = ~n12442 & ~n29459;
  assign n29461 = n11858 & ~n29460;
  assign n29462 = ~n29458 & ~n29460;
  assign n29463 = n11858 & n29462;
  assign n29464 = ~n29458 & n29461;
  assign n29465 = ~n29141 & ~n36149;
  assign n29466 = ~n11858 & ~n29462;
  assign n29467 = n11229 & ~n29466;
  assign n29468 = ~n29465 & n29467;
  assign n29469 = ~n29133 & ~n29468;
  assign n29470 = ~n29465 & ~n29466;
  assign n29471 = ~n11229 & ~n29470;
  assign n29472 = n10681 & ~n29471;
  assign n29473 = ~n29469 & ~n29471;
  assign n29474 = n10681 & n29473;
  assign n29475 = ~n29469 & n29472;
  assign n29476 = ~n29125 & ~n36150;
  assign n29477 = ~n10681 & ~n29473;
  assign n29478 = n10086 & ~n29477;
  assign n29479 = ~n29476 & n29478;
  assign n29480 = ~n28317 & ~n35997;
  assign n29481 = ~n28317 & ~n28917;
  assign n29482 = ~n35997 & n29481;
  assign n29483 = ~n28917 & n29480;
  assign n29484 = n28325 & ~n36151;
  assign n29485 = n28329 & n29481;
  assign n29486 = ~n28317 & n28325;
  assign n29487 = ~n35997 & n29486;
  assign n29488 = ~n28917 & n29487;
  assign n29489 = ~n28325 & ~n36151;
  assign n29490 = ~n29488 & ~n29489;
  assign n29491 = ~n29484 & ~n29485;
  assign n29492 = ~n29479 & ~n36152;
  assign n29493 = ~n29476 & ~n29477;
  assign n29494 = ~n10086 & ~n29493;
  assign n29495 = n9565 & ~n29494;
  assign n29496 = ~n29492 & ~n29494;
  assign n29497 = n9565 & n29496;
  assign n29498 = ~n29492 & n29495;
  assign n29499 = ~n29117 & ~n36153;
  assign n29500 = ~n9565 & ~n29496;
  assign n29501 = n8998 & ~n29500;
  assign n29502 = ~n29499 & n29501;
  assign n29503 = ~n29109 & ~n29502;
  assign n29504 = ~n29499 & ~n29500;
  assign n29505 = ~n8998 & ~n29504;
  assign n29506 = n8506 & ~n29505;
  assign n29507 = ~n29503 & ~n29505;
  assign n29508 = n8506 & n29507;
  assign n29509 = ~n29503 & n29506;
  assign n29510 = ~n29101 & ~n36154;
  assign n29511 = ~n8506 & ~n29507;
  assign n29512 = n7975 & ~n29511;
  assign n29513 = ~n29510 & n29512;
  assign n29514 = ~n28383 & ~n36006;
  assign n29515 = ~n28383 & ~n28917;
  assign n29516 = ~n36006 & n29515;
  assign n29517 = ~n28917 & n29514;
  assign n29518 = n28391 & ~n36155;
  assign n29519 = n28395 & n29515;
  assign n29520 = ~n28383 & n28391;
  assign n29521 = ~n36006 & n29520;
  assign n29522 = ~n28917 & n29521;
  assign n29523 = ~n28391 & ~n36155;
  assign n29524 = ~n29522 & ~n29523;
  assign n29525 = ~n29518 & ~n29519;
  assign n29526 = ~n29513 & ~n36156;
  assign n29527 = ~n29510 & ~n29511;
  assign n29528 = ~n7975 & ~n29527;
  assign n29529 = n7512 & ~n29528;
  assign n29530 = ~n29526 & ~n29528;
  assign n29531 = n7512 & n29530;
  assign n29532 = ~n29526 & n29529;
  assign n29533 = ~n29093 & ~n36157;
  assign n29534 = ~n7512 & ~n29530;
  assign n29535 = n7015 & ~n29534;
  assign n29536 = ~n29533 & n29535;
  assign n29537 = ~n29085 & ~n29536;
  assign n29538 = ~n29533 & ~n29534;
  assign n29539 = ~n7015 & ~n29538;
  assign n29540 = n6579 & ~n29539;
  assign n29541 = ~n29537 & ~n29539;
  assign n29542 = n6579 & n29541;
  assign n29543 = ~n29537 & n29540;
  assign n29544 = ~n29077 & ~n36158;
  assign n29545 = ~n6579 & ~n29541;
  assign n29546 = n6117 & ~n29545;
  assign n29547 = ~n29544 & n29546;
  assign n29548 = ~n28449 & ~n36015;
  assign n29549 = ~n28449 & ~n28917;
  assign n29550 = ~n36015 & n29549;
  assign n29551 = ~n28917 & n29548;
  assign n29552 = n28457 & ~n36159;
  assign n29553 = n28461 & n29549;
  assign n29554 = ~n28449 & n28457;
  assign n29555 = ~n36015 & n29554;
  assign n29556 = ~n28917 & n29555;
  assign n29557 = ~n28457 & ~n36159;
  assign n29558 = ~n29556 & ~n29557;
  assign n29559 = ~n29552 & ~n29553;
  assign n29560 = ~n29547 & ~n36160;
  assign n29561 = ~n29544 & ~n29545;
  assign n29562 = ~n6117 & ~n29561;
  assign n29563 = n5708 & ~n29562;
  assign n29564 = ~n29560 & ~n29562;
  assign n29565 = n5708 & n29564;
  assign n29566 = ~n29560 & n29563;
  assign n29567 = ~n29069 & ~n36161;
  assign n29568 = ~n5708 & ~n29564;
  assign n29569 = n5278 & ~n29568;
  assign n29570 = ~n29567 & n29569;
  assign n29571 = ~n29061 & ~n29570;
  assign n29572 = ~n29567 & ~n29568;
  assign n29573 = ~n5278 & ~n29572;
  assign n29574 = n4903 & ~n29573;
  assign n29575 = ~n29571 & ~n29573;
  assign n29576 = n4903 & n29575;
  assign n29577 = ~n29571 & n29574;
  assign n29578 = ~n29053 & ~n36162;
  assign n29579 = ~n4903 & ~n29575;
  assign n29580 = n4508 & ~n29579;
  assign n29581 = ~n29578 & n29580;
  assign n29582 = ~n28515 & ~n36024;
  assign n29583 = ~n28515 & ~n28917;
  assign n29584 = ~n36024 & n29583;
  assign n29585 = ~n28917 & n29582;
  assign n29586 = n28523 & ~n36163;
  assign n29587 = n28527 & n29583;
  assign n29588 = ~n28515 & n28523;
  assign n29589 = ~n36024 & n29588;
  assign n29590 = ~n28917 & n29589;
  assign n29591 = ~n28523 & ~n36163;
  assign n29592 = ~n29590 & ~n29591;
  assign n29593 = ~n29586 & ~n29587;
  assign n29594 = ~n29581 & ~n36164;
  assign n29595 = ~n29578 & ~n29579;
  assign n29596 = ~n4508 & ~n29595;
  assign n29597 = n4155 & ~n29596;
  assign n29598 = ~n29594 & ~n29596;
  assign n29599 = n4155 & n29598;
  assign n29600 = ~n29594 & n29597;
  assign n29601 = ~n29045 & ~n36165;
  assign n29602 = ~n4155 & ~n29598;
  assign n29603 = n3788 & ~n29602;
  assign n29604 = ~n29601 & n29603;
  assign n29605 = ~n29037 & ~n29604;
  assign n29606 = ~n29601 & ~n29602;
  assign n29607 = ~n3788 & ~n29606;
  assign n29608 = n3473 & ~n29607;
  assign n29609 = ~n29605 & ~n29607;
  assign n29610 = n3473 & n29609;
  assign n29611 = ~n29605 & n29608;
  assign n29612 = ~n29029 & ~n36166;
  assign n29613 = ~n3473 & ~n29609;
  assign n29614 = n3140 & ~n29613;
  assign n29615 = ~n29612 & n29614;
  assign n29616 = ~n28581 & ~n36033;
  assign n29617 = ~n28581 & ~n28917;
  assign n29618 = ~n36033 & n29617;
  assign n29619 = ~n28917 & n29616;
  assign n29620 = n28589 & ~n36167;
  assign n29621 = n28593 & n29617;
  assign n29622 = ~n28581 & n28589;
  assign n29623 = ~n36033 & n29622;
  assign n29624 = ~n28917 & n29623;
  assign n29625 = ~n28589 & ~n36167;
  assign n29626 = ~n29624 & ~n29625;
  assign n29627 = ~n29620 & ~n29621;
  assign n29628 = ~n29615 & ~n36168;
  assign n29629 = ~n29612 & ~n29613;
  assign n29630 = ~n3140 & ~n29629;
  assign n29631 = n2855 & ~n29630;
  assign n29632 = ~n29628 & ~n29630;
  assign n29633 = n2855 & n29632;
  assign n29634 = ~n29628 & n29631;
  assign n29635 = ~n29021 & ~n36169;
  assign n29636 = ~n2855 & ~n29632;
  assign n29637 = n2556 & ~n29636;
  assign n29638 = ~n29635 & n29637;
  assign n29639 = ~n29013 & ~n29638;
  assign n29640 = ~n29635 & ~n29636;
  assign n29641 = ~n2556 & ~n29640;
  assign n29642 = n2301 & ~n29641;
  assign n29643 = ~n29639 & ~n29641;
  assign n29644 = n2301 & n29643;
  assign n29645 = ~n29639 & n29642;
  assign n29646 = ~n29005 & ~n36170;
  assign n29647 = ~n2301 & ~n29643;
  assign n29648 = n2038 & ~n29647;
  assign n29649 = ~n29646 & n29648;
  assign n29650 = ~n28647 & ~n36042;
  assign n29651 = ~n28647 & ~n28917;
  assign n29652 = ~n36042 & n29651;
  assign n29653 = ~n28917 & n29650;
  assign n29654 = n28655 & ~n36171;
  assign n29655 = n28659 & n29651;
  assign n29656 = ~n28647 & n28655;
  assign n29657 = ~n36042 & n29656;
  assign n29658 = ~n28917 & n29657;
  assign n29659 = ~n28655 & ~n36171;
  assign n29660 = ~n29658 & ~n29659;
  assign n29661 = ~n29654 & ~n29655;
  assign n29662 = ~n29649 & ~n36172;
  assign n29663 = ~n29646 & ~n29647;
  assign n29664 = ~n2038 & ~n29663;
  assign n29665 = n1812 & ~n29664;
  assign n29666 = ~n29662 & ~n29664;
  assign n29667 = n1812 & n29666;
  assign n29668 = ~n29662 & n29665;
  assign n29669 = ~n28997 & ~n36173;
  assign n29670 = ~n1812 & ~n29666;
  assign n29671 = n1582 & ~n29670;
  assign n29672 = ~n29669 & n29671;
  assign n29673 = ~n28989 & ~n29672;
  assign n29674 = ~n29669 & ~n29670;
  assign n29675 = ~n1582 & ~n29674;
  assign n29676 = n1388 & ~n29675;
  assign n29677 = ~n29673 & ~n29675;
  assign n29678 = n1388 & n29677;
  assign n29679 = ~n29673 & n29676;
  assign n29680 = ~n28981 & ~n36174;
  assign n29681 = ~n1388 & ~n29677;
  assign n29682 = n1192 & ~n29681;
  assign n29683 = ~n29680 & n29682;
  assign n29684 = ~n28713 & ~n36051;
  assign n29685 = ~n28713 & ~n28917;
  assign n29686 = ~n36051 & n29685;
  assign n29687 = ~n28917 & n29684;
  assign n29688 = n28721 & ~n36175;
  assign n29689 = n28725 & n29685;
  assign n29690 = ~n28713 & n28721;
  assign n29691 = ~n36051 & n29690;
  assign n29692 = ~n28917 & n29691;
  assign n29693 = ~n28721 & ~n36175;
  assign n29694 = ~n29692 & ~n29693;
  assign n29695 = ~n29688 & ~n29689;
  assign n29696 = ~n29683 & ~n36176;
  assign n29697 = ~n29680 & ~n29681;
  assign n29698 = ~n1192 & ~n29697;
  assign n29699 = n1028 & ~n29698;
  assign n29700 = ~n29696 & ~n29698;
  assign n29701 = n1028 & n29700;
  assign n29702 = ~n29696 & n29699;
  assign n29703 = ~n28973 & ~n36177;
  assign n29704 = ~n1028 & ~n29700;
  assign n29705 = n866 & ~n29704;
  assign n29706 = ~n29703 & n29705;
  assign n29707 = ~n28965 & ~n29706;
  assign n29708 = ~n29703 & ~n29704;
  assign n29709 = ~n866 & ~n29708;
  assign n29710 = n730 & ~n29709;
  assign n29711 = ~n29707 & ~n29709;
  assign n29712 = n730 & n29711;
  assign n29713 = ~n29707 & n29710;
  assign n29714 = ~n28957 & ~n36178;
  assign n29715 = ~n730 & ~n29711;
  assign n29716 = n602 & ~n29715;
  assign n29717 = ~n29714 & n29716;
  assign n29718 = ~n28779 & ~n36060;
  assign n29719 = ~n28779 & ~n28917;
  assign n29720 = ~n36060 & n29719;
  assign n29721 = ~n28917 & n29718;
  assign n29722 = n28787 & ~n36179;
  assign n29723 = n28791 & n29719;
  assign n29724 = ~n28779 & n28787;
  assign n29725 = ~n36060 & n29724;
  assign n29726 = ~n28917 & n29725;
  assign n29727 = ~n28787 & ~n36179;
  assign n29728 = ~n29726 & ~n29727;
  assign n29729 = ~n29722 & ~n29723;
  assign n29730 = ~n29717 & ~n36180;
  assign n29731 = ~n29714 & ~n29715;
  assign n29732 = ~n602 & ~n29731;
  assign n29733 = n497 & ~n29732;
  assign n29734 = ~n29730 & ~n29732;
  assign n29735 = n497 & n29734;
  assign n29736 = ~n29730 & n29733;
  assign n29737 = ~n28949 & ~n36181;
  assign n29738 = ~n497 & ~n29734;
  assign n29739 = n403 & ~n29738;
  assign n29740 = ~n29737 & n29739;
  assign n29741 = ~n28941 & ~n29740;
  assign n29742 = ~n29737 & ~n29738;
  assign n29743 = ~n403 & ~n29742;
  assign n29744 = n330 & ~n29743;
  assign n29745 = ~n29741 & ~n29743;
  assign n29746 = n330 & n29745;
  assign n29747 = ~n29741 & n29744;
  assign n29748 = ~n28933 & ~n36182;
  assign n29749 = ~n330 & ~n29745;
  assign n29750 = ~n29748 & ~n29749;
  assign n29751 = ~n271 & ~n29750;
  assign n29752 = n271 & ~n29749;
  assign n29753 = ~n29748 & n29752;
  assign n29754 = ~n28841 & ~n36067;
  assign n29755 = ~n28917 & n29754;
  assign n29756 = ~n36069 & ~n29755;
  assign n29757 = ~n28841 & n36069;
  assign n29758 = ~n36067 & n29757;
  assign n29759 = n36069 & n29755;
  assign n29760 = ~n28917 & n29758;
  assign n29761 = n36069 & ~n29755;
  assign n29762 = ~n36069 & n29755;
  assign n29763 = ~n29761 & ~n29762;
  assign n29764 = ~n29756 & ~n36183;
  assign n29765 = ~n29753 & n36184;
  assign n29766 = ~n29751 & ~n29765;
  assign n29767 = ~n217 & ~n29766;
  assign n29768 = n217 & ~n29751;
  assign n29769 = n217 & n29766;
  assign n29770 = ~n29765 & n29768;
  assign n29771 = ~n28925 & ~n36185;
  assign n29772 = ~n29767 & ~n29771;
  assign n29773 = ~n198 & ~n29772;
  assign n29774 = n198 & ~n29767;
  assign n29775 = ~n29771 & n29774;
  assign n29776 = ~n28863 & ~n36071;
  assign n29777 = ~n28863 & ~n28917;
  assign n29778 = ~n36071 & n29777;
  assign n29779 = ~n28917 & n29776;
  assign n29780 = n28871 & ~n36186;
  assign n29781 = n28875 & n29777;
  assign n29782 = ~n28863 & n28871;
  assign n29783 = ~n36071 & n29782;
  assign n29784 = ~n28917 & n29783;
  assign n29785 = ~n28871 & ~n36186;
  assign n29786 = ~n29784 & ~n29785;
  assign n29787 = ~n29780 & ~n29781;
  assign n29788 = ~n29775 & ~n36187;
  assign n29789 = ~n29773 & ~n29788;
  assign n29790 = ~n28877 & ~n28879;
  assign n29791 = ~n28917 & n29790;
  assign n29792 = ~n36073 & ~n29791;
  assign n29793 = ~n28879 & n36073;
  assign n29794 = ~n28877 & n29793;
  assign n29795 = n36073 & n29791;
  assign n29796 = ~n28917 & n29794;
  assign n29797 = ~n29792 & ~n36188;
  assign n29798 = ~n28893 & ~n28901;
  assign n29799 = ~n28901 & ~n28917;
  assign n29800 = ~n28893 & n29799;
  assign n29801 = ~n28917 & n29798;
  assign n29802 = ~n36076 & ~n36189;
  assign n29803 = ~n29797 & n29802;
  assign n29804 = ~n29789 & n29803;
  assign n29805 = n193 & ~n29804;
  assign n29806 = ~n29773 & n29797;
  assign n29807 = n29789 & n29797;
  assign n29808 = ~n29788 & n29806;
  assign n29809 = n28893 & ~n29799;
  assign n29810 = ~n193 & ~n29798;
  assign n29811 = ~n29809 & n29810;
  assign n29812 = ~n36190 & ~n29811;
  assign n29813 = ~n29805 & n29812;
  assign n29814 = ~n29767 & ~n36185;
  assign n29815 = ~n29767 & ~n29813;
  assign n29816 = ~n36185 & n29815;
  assign n29817 = ~n29813 & n29814;
  assign n29818 = n28925 & ~n36191;
  assign n29819 = n29771 & n29815;
  assign n29820 = n28925 & ~n36185;
  assign n29821 = ~n29767 & n29820;
  assign n29822 = ~n29813 & n29821;
  assign n29823 = ~n28925 & ~n36191;
  assign n29824 = ~n29822 & ~n29823;
  assign n29825 = ~n29818 & ~n29819;
  assign n29826 = pi4  & ~n29813;
  assign n29827 = ~pi2  & ~pi3 ;
  assign n29828 = ~pi4  & n29827;
  assign n29829 = ~pi4  & ~n29827;
  assign n29830 = pi4  & n29813;
  assign n29831 = ~n29829 & ~n29830;
  assign n29832 = ~n29826 & ~n29828;
  assign n29833 = ~n28917 & n36193;
  assign n29834 = ~pi4  & ~n29813;
  assign n29835 = pi5  & ~n29834;
  assign n29836 = ~pi5  & n29834;
  assign n29837 = n29228 & ~n29813;
  assign n29838 = ~n29835 & ~n36194;
  assign n29839 = ~n28915 & ~n29828;
  assign n29840 = ~n36076 & n29839;
  assign n29841 = ~n28909 & n29840;
  assign n29842 = n28917 & ~n36193;
  assign n29843 = ~n29826 & n29841;
  assign n29844 = n29838 & ~n36195;
  assign n29845 = ~n29833 & ~n29844;
  assign n29846 = ~n27931 & ~n29845;
  assign n29847 = n27931 & ~n29833;
  assign n29848 = ~n29844 & n29847;
  assign n29849 = ~n28917 & ~n29811;
  assign n29850 = ~n36190 & n29849;
  assign n29851 = ~n28917 & n29813;
  assign n29852 = ~n29805 & n29850;
  assign n29853 = ~n36194 & ~n36196;
  assign n29854 = pi6  & ~n29853;
  assign n29855 = ~pi6  & ~n36196;
  assign n29856 = ~pi6  & n29853;
  assign n29857 = ~n36194 & n29855;
  assign n29858 = ~n29854 & ~n36197;
  assign n29859 = ~n29848 & ~n29858;
  assign n29860 = ~n29846 & ~n29859;
  assign n29861 = ~n27055 & ~n29860;
  assign n29862 = n27055 & ~n29846;
  assign n29863 = ~n29859 & n29862;
  assign n29864 = n27055 & n29860;
  assign n29865 = ~n36118 & ~n29242;
  assign n29866 = ~n29813 & n29865;
  assign n29867 = n29240 & ~n29866;
  assign n29868 = ~n29240 & n29865;
  assign n29869 = ~n29240 & n29866;
  assign n29870 = ~n29813 & n29868;
  assign n29871 = ~n29867 & ~n36199;
  assign n29872 = ~n36198 & ~n29871;
  assign n29873 = ~n29861 & ~n29872;
  assign n29874 = ~n26098 & ~n29873;
  assign n29875 = n26098 & ~n29861;
  assign n29876 = ~n29872 & n29875;
  assign n29877 = ~n36119 & ~n29248;
  assign n29878 = ~n29248 & ~n29813;
  assign n29879 = ~n36119 & n29878;
  assign n29880 = ~n29813 & n29877;
  assign n29881 = n29226 & ~n36200;
  assign n29882 = n29247 & n29878;
  assign n29883 = n29226 & ~n36119;
  assign n29884 = ~n29248 & n29883;
  assign n29885 = ~n29813 & n29884;
  assign n29886 = ~n29226 & ~n36200;
  assign n29887 = ~n29885 & ~n29886;
  assign n29888 = ~n29881 & ~n29882;
  assign n29889 = ~n29876 & ~n36201;
  assign n29890 = ~n29874 & ~n29889;
  assign n29891 = ~n25256 & ~n29890;
  assign n29892 = n25256 & ~n29874;
  assign n29893 = ~n29889 & n29892;
  assign n29894 = n25256 & n29890;
  assign n29895 = ~n29250 & ~n29260;
  assign n29896 = ~n29813 & n29895;
  assign n29897 = n29257 & ~n29896;
  assign n29898 = ~n29257 & n29896;
  assign n29899 = n29257 & ~n29260;
  assign n29900 = ~n29250 & n29899;
  assign n29901 = n29257 & n29896;
  assign n29902 = ~n29813 & n29900;
  assign n29903 = ~n29257 & ~n29896;
  assign n29904 = ~n36203 & ~n29903;
  assign n29905 = ~n29897 & ~n29898;
  assign n29906 = ~n36202 & ~n36204;
  assign n29907 = ~n29891 & ~n29906;
  assign n29908 = ~n24331 & ~n29907;
  assign n29909 = n24331 & ~n29891;
  assign n29910 = ~n29906 & n29909;
  assign n29911 = ~n36121 & ~n29266;
  assign n29912 = ~n29266 & ~n29813;
  assign n29913 = ~n36121 & n29912;
  assign n29914 = ~n29813 & n29911;
  assign n29915 = n29213 & ~n36205;
  assign n29916 = n29265 & n29912;
  assign n29917 = n29213 & ~n36121;
  assign n29918 = ~n29266 & n29917;
  assign n29919 = ~n29813 & n29918;
  assign n29920 = ~n29213 & ~n36205;
  assign n29921 = ~n29919 & ~n29920;
  assign n29922 = ~n29915 & ~n29916;
  assign n29923 = ~n29910 & ~n36206;
  assign n29924 = ~n29908 & ~n29923;
  assign n29925 = ~n23517 & ~n29924;
  assign n29926 = n23517 & ~n29908;
  assign n29927 = ~n29923 & n29926;
  assign n29928 = n23517 & n29924;
  assign n29929 = ~n29268 & ~n29282;
  assign n29930 = ~n29813 & n29929;
  assign n29931 = ~n36123 & n29930;
  assign n29932 = n36123 & ~n29930;
  assign n29933 = n36123 & ~n29282;
  assign n29934 = ~n29268 & n29933;
  assign n29935 = ~n29813 & n29934;
  assign n29936 = ~n36123 & ~n29930;
  assign n29937 = ~n29935 & ~n29936;
  assign n29938 = ~n29931 & ~n29932;
  assign n29939 = ~n36207 & ~n36208;
  assign n29940 = ~n29925 & ~n29939;
  assign n29941 = ~n22625 & ~n29940;
  assign n29942 = n22625 & ~n29925;
  assign n29943 = ~n29939 & n29942;
  assign n29944 = ~n36124 & ~n29288;
  assign n29945 = ~n29288 & ~n29813;
  assign n29946 = ~n36124 & n29945;
  assign n29947 = ~n29813 & n29944;
  assign n29948 = n29205 & ~n36209;
  assign n29949 = n29287 & n29945;
  assign n29950 = n29205 & ~n36124;
  assign n29951 = ~n29288 & n29950;
  assign n29952 = ~n29813 & n29951;
  assign n29953 = ~n29205 & ~n36209;
  assign n29954 = ~n29952 & ~n29953;
  assign n29955 = ~n29948 & ~n29949;
  assign n29956 = ~n29943 & ~n36210;
  assign n29957 = ~n29941 & ~n29956;
  assign n29958 = ~n21842 & ~n29957;
  assign n29959 = n21842 & ~n29941;
  assign n29960 = ~n29956 & n29959;
  assign n29961 = n21842 & n29957;
  assign n29962 = ~n29290 & ~n29303;
  assign n29963 = ~n29813 & n29962;
  assign n29964 = ~n36125 & ~n29963;
  assign n29965 = n36125 & ~n29303;
  assign n29966 = ~n29290 & n29965;
  assign n29967 = n36125 & n29963;
  assign n29968 = ~n29813 & n29966;
  assign n29969 = n36125 & ~n29963;
  assign n29970 = ~n36125 & n29963;
  assign n29971 = ~n29969 & ~n29970;
  assign n29972 = ~n29964 & ~n36212;
  assign n29973 = ~n36211 & n36213;
  assign n29974 = ~n29958 & ~n29973;
  assign n29975 = ~n20986 & ~n29974;
  assign n29976 = n20986 & ~n29958;
  assign n29977 = ~n29973 & n29976;
  assign n29978 = ~n36126 & ~n29309;
  assign n29979 = ~n29309 & ~n29813;
  assign n29980 = ~n36126 & n29979;
  assign n29981 = ~n29813 & n29978;
  assign n29982 = n29197 & ~n36214;
  assign n29983 = n29308 & n29979;
  assign n29984 = n29197 & ~n36126;
  assign n29985 = ~n29309 & n29984;
  assign n29986 = ~n29813 & n29985;
  assign n29987 = ~n29197 & ~n36214;
  assign n29988 = ~n29986 & ~n29987;
  assign n29989 = ~n29982 & ~n29983;
  assign n29990 = ~n29977 & ~n36215;
  assign n29991 = ~n29975 & ~n29990;
  assign n29992 = ~n20229 & ~n29991;
  assign n29993 = n20229 & ~n29975;
  assign n29994 = ~n29990 & n29993;
  assign n29995 = n20229 & n29991;
  assign n29996 = ~n29311 & ~n29325;
  assign n29997 = ~n29813 & n29996;
  assign n29998 = n36128 & ~n29997;
  assign n29999 = ~n36128 & ~n29325;
  assign n30000 = ~n29311 & n29999;
  assign n30001 = ~n36128 & n29997;
  assign n30002 = ~n29813 & n30000;
  assign n30003 = n36128 & n29997;
  assign n30004 = ~n36128 & ~n29997;
  assign n30005 = ~n30003 & ~n30004;
  assign n30006 = ~n29998 & ~n36217;
  assign n30007 = ~n36216 & n36218;
  assign n30008 = ~n29992 & ~n30007;
  assign n30009 = ~n19401 & ~n30008;
  assign n30010 = n19401 & ~n29992;
  assign n30011 = ~n30007 & n30010;
  assign n30012 = ~n36129 & ~n29331;
  assign n30013 = ~n29331 & ~n29813;
  assign n30014 = ~n36129 & n30013;
  assign n30015 = ~n29813 & n30012;
  assign n30016 = n29189 & ~n36219;
  assign n30017 = n29330 & n30013;
  assign n30018 = n29189 & ~n36129;
  assign n30019 = ~n29331 & n30018;
  assign n30020 = ~n29813 & n30019;
  assign n30021 = ~n29189 & ~n36219;
  assign n30022 = ~n30020 & ~n30021;
  assign n30023 = ~n30016 & ~n30017;
  assign n30024 = ~n30011 & ~n36220;
  assign n30025 = ~n30009 & ~n30024;
  assign n30026 = ~n18676 & ~n30025;
  assign n30027 = n18676 & ~n30009;
  assign n30028 = ~n30024 & n30027;
  assign n30029 = n18676 & n30025;
  assign n30030 = ~n29333 & ~n29347;
  assign n30031 = ~n29347 & ~n29813;
  assign n30032 = ~n29333 & n30031;
  assign n30033 = ~n29813 & n30030;
  assign n30034 = ~n36131 & ~n36222;
  assign n30035 = n29345 & n30031;
  assign n30036 = n36131 & n36222;
  assign n30037 = ~n36131 & ~n29347;
  assign n30038 = ~n29333 & n30037;
  assign n30039 = ~n29813 & n30038;
  assign n30040 = n36131 & ~n36222;
  assign n30041 = ~n30039 & ~n30040;
  assign n30042 = ~n30034 & ~n36223;
  assign n30043 = ~n36221 & ~n36224;
  assign n30044 = ~n30026 & ~n30043;
  assign n30045 = ~n17885 & ~n30044;
  assign n30046 = n17885 & ~n30026;
  assign n30047 = ~n30043 & n30046;
  assign n30048 = ~n36132 & ~n29353;
  assign n30049 = ~n29353 & ~n29813;
  assign n30050 = ~n36132 & n30049;
  assign n30051 = ~n29813 & n30048;
  assign n30052 = n29181 & ~n36225;
  assign n30053 = n29352 & n30049;
  assign n30054 = n29181 & ~n36132;
  assign n30055 = ~n29353 & n30054;
  assign n30056 = ~n29813 & n30055;
  assign n30057 = ~n29181 & ~n36225;
  assign n30058 = ~n30056 & ~n30057;
  assign n30059 = ~n30052 & ~n30053;
  assign n30060 = ~n30047 & ~n36226;
  assign n30061 = ~n30045 & ~n30060;
  assign n30062 = ~n17187 & ~n30061;
  assign n30063 = n17187 & ~n30045;
  assign n30064 = ~n30060 & n30063;
  assign n30065 = n17187 & n30061;
  assign n30066 = ~n29355 & ~n29371;
  assign n30067 = ~n29813 & n30066;
  assign n30068 = ~n36135 & ~n30067;
  assign n30069 = n36135 & ~n29371;
  assign n30070 = ~n29355 & n30069;
  assign n30071 = n36135 & n30067;
  assign n30072 = ~n29813 & n30070;
  assign n30073 = ~n30068 & ~n36228;
  assign n30074 = ~n36227 & ~n30073;
  assign n30075 = ~n30062 & ~n30074;
  assign n30076 = ~n16428 & ~n30075;
  assign n30077 = n16428 & ~n30062;
  assign n30078 = ~n30074 & n30077;
  assign n30079 = ~n36136 & ~n29377;
  assign n30080 = ~n29377 & ~n29813;
  assign n30081 = ~n36136 & n30080;
  assign n30082 = ~n29813 & n30079;
  assign n30083 = n29173 & ~n36229;
  assign n30084 = n29376 & n30080;
  assign n30085 = n29173 & ~n36136;
  assign n30086 = ~n29377 & n30085;
  assign n30087 = ~n29813 & n30086;
  assign n30088 = ~n29173 & ~n36229;
  assign n30089 = ~n30087 & ~n30088;
  assign n30090 = ~n30083 & ~n30084;
  assign n30091 = ~n30078 & ~n36230;
  assign n30092 = ~n30076 & ~n30091;
  assign n30093 = ~n15760 & ~n30092;
  assign n30094 = n15760 & ~n30076;
  assign n30095 = ~n30091 & n30094;
  assign n30096 = n15760 & n30092;
  assign n30097 = ~n29379 & ~n29390;
  assign n30098 = ~n29390 & ~n29813;
  assign n30099 = ~n29379 & n30098;
  assign n30100 = ~n29813 & n30097;
  assign n30101 = n29387 & ~n36232;
  assign n30102 = n29388 & n30098;
  assign n30103 = ~n29387 & n36232;
  assign n30104 = n29387 & ~n29390;
  assign n30105 = ~n29379 & n30104;
  assign n30106 = ~n29813 & n30105;
  assign n30107 = ~n29387 & ~n36232;
  assign n30108 = ~n30106 & ~n30107;
  assign n30109 = ~n30101 & ~n36233;
  assign n30110 = ~n36231 & ~n36234;
  assign n30111 = ~n30093 & ~n30110;
  assign n30112 = ~n15033 & ~n30111;
  assign n30113 = n15033 & ~n30093;
  assign n30114 = ~n30110 & n30113;
  assign n30115 = ~n36138 & ~n29396;
  assign n30116 = ~n29396 & ~n29813;
  assign n30117 = ~n36138 & n30116;
  assign n30118 = ~n29813 & n30115;
  assign n30119 = n29165 & ~n36235;
  assign n30120 = n29395 & n30116;
  assign n30121 = n29165 & ~n36138;
  assign n30122 = ~n29396 & n30121;
  assign n30123 = ~n29813 & n30122;
  assign n30124 = ~n29165 & ~n36235;
  assign n30125 = ~n30123 & ~n30124;
  assign n30126 = ~n30119 & ~n30120;
  assign n30127 = ~n30114 & ~n36236;
  assign n30128 = ~n30112 & ~n30127;
  assign n30129 = ~n14394 & ~n30128;
  assign n30130 = n14394 & ~n30112;
  assign n30131 = ~n30127 & n30130;
  assign n30132 = n14394 & n30128;
  assign n30133 = ~n29398 & ~n29414;
  assign n30134 = ~n29813 & n30133;
  assign n30135 = ~n36141 & n30134;
  assign n30136 = n36141 & ~n30134;
  assign n30137 = n36141 & ~n29414;
  assign n30138 = ~n29398 & n30137;
  assign n30139 = n36141 & n30134;
  assign n30140 = ~n29813 & n30138;
  assign n30141 = ~n36141 & ~n30134;
  assign n30142 = ~n36238 & ~n30141;
  assign n30143 = ~n30135 & ~n30136;
  assign n30144 = ~n36237 & ~n36239;
  assign n30145 = ~n30129 & ~n30144;
  assign n30146 = ~n13704 & ~n30145;
  assign n30147 = n13704 & ~n30129;
  assign n30148 = ~n30144 & n30147;
  assign n30149 = ~n36142 & ~n29420;
  assign n30150 = ~n29420 & ~n29813;
  assign n30151 = ~n36142 & n30150;
  assign n30152 = ~n29813 & n30149;
  assign n30153 = n29157 & ~n36240;
  assign n30154 = n29419 & n30150;
  assign n30155 = n29157 & ~n36142;
  assign n30156 = ~n29420 & n30155;
  assign n30157 = ~n29813 & n30156;
  assign n30158 = ~n29157 & ~n36240;
  assign n30159 = ~n30157 & ~n30158;
  assign n30160 = ~n30153 & ~n30154;
  assign n30161 = ~n30148 & ~n36241;
  assign n30162 = ~n30146 & ~n30161;
  assign n30163 = ~n13099 & ~n30162;
  assign n30164 = n13099 & ~n30146;
  assign n30165 = ~n30161 & n30164;
  assign n30166 = n13099 & n30162;
  assign n30167 = ~n29422 & ~n29436;
  assign n30168 = ~n29436 & ~n29813;
  assign n30169 = ~n29422 & n30168;
  assign n30170 = ~n29813 & n30167;
  assign n30171 = n36144 & ~n36243;
  assign n30172 = n29434 & n30168;
  assign n30173 = ~n36144 & n36243;
  assign n30174 = n36144 & ~n29436;
  assign n30175 = ~n29422 & n30174;
  assign n30176 = ~n29813 & n30175;
  assign n30177 = ~n36144 & ~n36243;
  assign n30178 = ~n30176 & ~n30177;
  assign n30179 = ~n30171 & ~n36244;
  assign n30180 = ~n36242 & ~n36245;
  assign n30181 = ~n30163 & ~n30180;
  assign n30182 = ~n12442 & ~n30181;
  assign n30183 = n12442 & ~n30163;
  assign n30184 = ~n30180 & n30183;
  assign n30185 = ~n36145 & ~n29442;
  assign n30186 = ~n29442 & ~n29813;
  assign n30187 = ~n36145 & n30186;
  assign n30188 = ~n29813 & n30185;
  assign n30189 = n29149 & ~n36246;
  assign n30190 = n29441 & n30186;
  assign n30191 = n29149 & ~n36145;
  assign n30192 = ~n29442 & n30191;
  assign n30193 = ~n29813 & n30192;
  assign n30194 = ~n29149 & ~n36246;
  assign n30195 = ~n30193 & ~n30194;
  assign n30196 = ~n30189 & ~n30190;
  assign n30197 = ~n30184 & ~n36247;
  assign n30198 = ~n30182 & ~n30197;
  assign n30199 = ~n11858 & ~n30198;
  assign n30200 = ~n29444 & ~n29460;
  assign n30201 = ~n29813 & n30200;
  assign n30202 = ~n36148 & ~n30201;
  assign n30203 = n36148 & ~n29460;
  assign n30204 = ~n29444 & n30203;
  assign n30205 = n36148 & n30201;
  assign n30206 = ~n29813 & n30204;
  assign n30207 = ~n30202 & ~n36248;
  assign n30208 = n11858 & ~n30182;
  assign n30209 = ~n30197 & n30208;
  assign n30210 = n11858 & n30198;
  assign n30211 = ~n30207 & ~n36249;
  assign n30212 = ~n30199 & ~n30211;
  assign n30213 = ~n11229 & ~n30212;
  assign n30214 = n11229 & ~n30199;
  assign n30215 = ~n30211 & n30214;
  assign n30216 = ~n36149 & ~n29466;
  assign n30217 = ~n29466 & ~n29813;
  assign n30218 = ~n36149 & n30217;
  assign n30219 = ~n29813 & n30216;
  assign n30220 = n29141 & ~n36250;
  assign n30221 = n29465 & n30217;
  assign n30222 = n29141 & ~n36149;
  assign n30223 = ~n29466 & n30222;
  assign n30224 = ~n29813 & n30223;
  assign n30225 = ~n29141 & ~n36250;
  assign n30226 = ~n30224 & ~n30225;
  assign n30227 = ~n30220 & ~n30221;
  assign n30228 = ~n30215 & ~n36251;
  assign n30229 = ~n30213 & ~n30228;
  assign n30230 = ~n10681 & ~n30229;
  assign n30231 = n10681 & ~n30213;
  assign n30232 = ~n30228 & n30231;
  assign n30233 = n10681 & n30229;
  assign n30234 = ~n29468 & ~n29471;
  assign n30235 = ~n29471 & ~n29813;
  assign n30236 = ~n29468 & n30235;
  assign n30237 = ~n29813 & n30234;
  assign n30238 = n29133 & ~n36253;
  assign n30239 = n29469 & n30235;
  assign n30240 = n29133 & ~n29471;
  assign n30241 = ~n29468 & n30240;
  assign n30242 = ~n29813 & n30241;
  assign n30243 = ~n29133 & ~n36253;
  assign n30244 = ~n30242 & ~n30243;
  assign n30245 = ~n30238 & ~n30239;
  assign n30246 = ~n36252 & ~n36254;
  assign n30247 = ~n30230 & ~n30246;
  assign n30248 = ~n10086 & ~n30247;
  assign n30249 = n10086 & ~n30230;
  assign n30250 = ~n30246 & n30249;
  assign n30251 = ~n36150 & ~n29477;
  assign n30252 = ~n29477 & ~n29813;
  assign n30253 = ~n36150 & n30252;
  assign n30254 = ~n29813 & n30251;
  assign n30255 = n29125 & ~n36255;
  assign n30256 = n29476 & n30252;
  assign n30257 = n29125 & ~n36150;
  assign n30258 = ~n29477 & n30257;
  assign n30259 = ~n29813 & n30258;
  assign n30260 = ~n29125 & ~n36255;
  assign n30261 = ~n30259 & ~n30260;
  assign n30262 = ~n30255 & ~n30256;
  assign n30263 = ~n30250 & ~n36256;
  assign n30264 = ~n30248 & ~n30263;
  assign n30265 = ~n9565 & ~n30264;
  assign n30266 = ~n29479 & ~n29494;
  assign n30267 = ~n29813 & n30266;
  assign n30268 = ~n36152 & ~n30267;
  assign n30269 = n36152 & ~n29494;
  assign n30270 = ~n29479 & n30269;
  assign n30271 = n36152 & n30267;
  assign n30272 = ~n29813 & n30270;
  assign n30273 = ~n30268 & ~n36257;
  assign n30274 = n9565 & ~n30248;
  assign n30275 = ~n30263 & n30274;
  assign n30276 = n9565 & n30264;
  assign n30277 = ~n30273 & ~n36258;
  assign n30278 = ~n30265 & ~n30277;
  assign n30279 = ~n8998 & ~n30278;
  assign n30280 = n8998 & ~n30265;
  assign n30281 = ~n30277 & n30280;
  assign n30282 = ~n36153 & ~n29500;
  assign n30283 = ~n29500 & ~n29813;
  assign n30284 = ~n36153 & n30283;
  assign n30285 = ~n29813 & n30282;
  assign n30286 = n29117 & ~n36259;
  assign n30287 = n29499 & n30283;
  assign n30288 = n29117 & ~n36153;
  assign n30289 = ~n29500 & n30288;
  assign n30290 = ~n29813 & n30289;
  assign n30291 = ~n29117 & ~n36259;
  assign n30292 = ~n30290 & ~n30291;
  assign n30293 = ~n30286 & ~n30287;
  assign n30294 = ~n30281 & ~n36260;
  assign n30295 = ~n30279 & ~n30294;
  assign n30296 = ~n8506 & ~n30295;
  assign n30297 = n8506 & ~n30279;
  assign n30298 = ~n30294 & n30297;
  assign n30299 = n8506 & n30295;
  assign n30300 = ~n29502 & ~n29505;
  assign n30301 = ~n29505 & ~n29813;
  assign n30302 = ~n29502 & n30301;
  assign n30303 = ~n29813 & n30300;
  assign n30304 = n29109 & ~n36262;
  assign n30305 = n29503 & n30301;
  assign n30306 = n29109 & ~n29505;
  assign n30307 = ~n29502 & n30306;
  assign n30308 = ~n29813 & n30307;
  assign n30309 = ~n29109 & ~n36262;
  assign n30310 = ~n30308 & ~n30309;
  assign n30311 = ~n30304 & ~n30305;
  assign n30312 = ~n36261 & ~n36263;
  assign n30313 = ~n30296 & ~n30312;
  assign n30314 = ~n7975 & ~n30313;
  assign n30315 = n7975 & ~n30296;
  assign n30316 = ~n30312 & n30315;
  assign n30317 = ~n36154 & ~n29511;
  assign n30318 = ~n29511 & ~n29813;
  assign n30319 = ~n36154 & n30318;
  assign n30320 = ~n29813 & n30317;
  assign n30321 = n29101 & ~n36264;
  assign n30322 = n29510 & n30318;
  assign n30323 = n29101 & ~n36154;
  assign n30324 = ~n29511 & n30323;
  assign n30325 = ~n29813 & n30324;
  assign n30326 = ~n29101 & ~n36264;
  assign n30327 = ~n30325 & ~n30326;
  assign n30328 = ~n30321 & ~n30322;
  assign n30329 = ~n30316 & ~n36265;
  assign n30330 = ~n30314 & ~n30329;
  assign n30331 = ~n7512 & ~n30330;
  assign n30332 = ~n29513 & ~n29528;
  assign n30333 = ~n29813 & n30332;
  assign n30334 = ~n36156 & ~n30333;
  assign n30335 = n36156 & ~n29528;
  assign n30336 = ~n29513 & n30335;
  assign n30337 = n36156 & n30333;
  assign n30338 = ~n29813 & n30336;
  assign n30339 = ~n30334 & ~n36266;
  assign n30340 = n7512 & ~n30314;
  assign n30341 = ~n30329 & n30340;
  assign n30342 = n7512 & n30330;
  assign n30343 = ~n30339 & ~n36267;
  assign n30344 = ~n30331 & ~n30343;
  assign n30345 = ~n7015 & ~n30344;
  assign n30346 = n7015 & ~n30331;
  assign n30347 = ~n30343 & n30346;
  assign n30348 = ~n36157 & ~n29534;
  assign n30349 = ~n29534 & ~n29813;
  assign n30350 = ~n36157 & n30349;
  assign n30351 = ~n29813 & n30348;
  assign n30352 = n29093 & ~n36268;
  assign n30353 = n29533 & n30349;
  assign n30354 = n29093 & ~n36157;
  assign n30355 = ~n29534 & n30354;
  assign n30356 = ~n29813 & n30355;
  assign n30357 = ~n29093 & ~n36268;
  assign n30358 = ~n30356 & ~n30357;
  assign n30359 = ~n30352 & ~n30353;
  assign n30360 = ~n30347 & ~n36269;
  assign n30361 = ~n30345 & ~n30360;
  assign n30362 = ~n6579 & ~n30361;
  assign n30363 = n6579 & ~n30345;
  assign n30364 = ~n30360 & n30363;
  assign n30365 = n6579 & n30361;
  assign n30366 = ~n29536 & ~n29539;
  assign n30367 = ~n29539 & ~n29813;
  assign n30368 = ~n29536 & n30367;
  assign n30369 = ~n29813 & n30366;
  assign n30370 = n29085 & ~n36271;
  assign n30371 = n29537 & n30367;
  assign n30372 = n29085 & ~n29539;
  assign n30373 = ~n29536 & n30372;
  assign n30374 = ~n29813 & n30373;
  assign n30375 = ~n29085 & ~n36271;
  assign n30376 = ~n30374 & ~n30375;
  assign n30377 = ~n30370 & ~n30371;
  assign n30378 = ~n36270 & ~n36272;
  assign n30379 = ~n30362 & ~n30378;
  assign n30380 = ~n6117 & ~n30379;
  assign n30381 = n6117 & ~n30362;
  assign n30382 = ~n30378 & n30381;
  assign n30383 = ~n36158 & ~n29545;
  assign n30384 = ~n29545 & ~n29813;
  assign n30385 = ~n36158 & n30384;
  assign n30386 = ~n29813 & n30383;
  assign n30387 = n29077 & ~n36273;
  assign n30388 = n29544 & n30384;
  assign n30389 = n29077 & ~n36158;
  assign n30390 = ~n29545 & n30389;
  assign n30391 = ~n29813 & n30390;
  assign n30392 = ~n29077 & ~n36273;
  assign n30393 = ~n30391 & ~n30392;
  assign n30394 = ~n30387 & ~n30388;
  assign n30395 = ~n30382 & ~n36274;
  assign n30396 = ~n30380 & ~n30395;
  assign n30397 = ~n5708 & ~n30396;
  assign n30398 = ~n29547 & ~n29562;
  assign n30399 = ~n29813 & n30398;
  assign n30400 = ~n36160 & ~n30399;
  assign n30401 = n36160 & ~n29562;
  assign n30402 = ~n29547 & n30401;
  assign n30403 = n36160 & n30399;
  assign n30404 = ~n29813 & n30402;
  assign n30405 = ~n30400 & ~n36275;
  assign n30406 = n5708 & ~n30380;
  assign n30407 = ~n30395 & n30406;
  assign n30408 = n5708 & n30396;
  assign n30409 = ~n30405 & ~n36276;
  assign n30410 = ~n30397 & ~n30409;
  assign n30411 = ~n5278 & ~n30410;
  assign n30412 = n5278 & ~n30397;
  assign n30413 = ~n30409 & n30412;
  assign n30414 = ~n36161 & ~n29568;
  assign n30415 = ~n29568 & ~n29813;
  assign n30416 = ~n36161 & n30415;
  assign n30417 = ~n29813 & n30414;
  assign n30418 = n29069 & ~n36277;
  assign n30419 = n29567 & n30415;
  assign n30420 = n29069 & ~n36161;
  assign n30421 = ~n29568 & n30420;
  assign n30422 = ~n29813 & n30421;
  assign n30423 = ~n29069 & ~n36277;
  assign n30424 = ~n30422 & ~n30423;
  assign n30425 = ~n30418 & ~n30419;
  assign n30426 = ~n30413 & ~n36278;
  assign n30427 = ~n30411 & ~n30426;
  assign n30428 = ~n4903 & ~n30427;
  assign n30429 = n4903 & ~n30411;
  assign n30430 = ~n30426 & n30429;
  assign n30431 = n4903 & n30427;
  assign n30432 = ~n29570 & ~n29573;
  assign n30433 = ~n29573 & ~n29813;
  assign n30434 = ~n29570 & n30433;
  assign n30435 = ~n29813 & n30432;
  assign n30436 = n29061 & ~n36280;
  assign n30437 = n29571 & n30433;
  assign n30438 = n29061 & ~n29573;
  assign n30439 = ~n29570 & n30438;
  assign n30440 = ~n29813 & n30439;
  assign n30441 = ~n29061 & ~n36280;
  assign n30442 = ~n30440 & ~n30441;
  assign n30443 = ~n30436 & ~n30437;
  assign n30444 = ~n36279 & ~n36281;
  assign n30445 = ~n30428 & ~n30444;
  assign n30446 = ~n4508 & ~n30445;
  assign n30447 = n4508 & ~n30428;
  assign n30448 = ~n30444 & n30447;
  assign n30449 = ~n36162 & ~n29579;
  assign n30450 = ~n29579 & ~n29813;
  assign n30451 = ~n36162 & n30450;
  assign n30452 = ~n29813 & n30449;
  assign n30453 = n29053 & ~n36282;
  assign n30454 = n29578 & n30450;
  assign n30455 = n29053 & ~n36162;
  assign n30456 = ~n29579 & n30455;
  assign n30457 = ~n29813 & n30456;
  assign n30458 = ~n29053 & ~n36282;
  assign n30459 = ~n30457 & ~n30458;
  assign n30460 = ~n30453 & ~n30454;
  assign n30461 = ~n30448 & ~n36283;
  assign n30462 = ~n30446 & ~n30461;
  assign n30463 = ~n4155 & ~n30462;
  assign n30464 = ~n29581 & ~n29596;
  assign n30465 = ~n29813 & n30464;
  assign n30466 = ~n36164 & ~n30465;
  assign n30467 = n36164 & ~n29596;
  assign n30468 = ~n29581 & n30467;
  assign n30469 = n36164 & n30465;
  assign n30470 = ~n29813 & n30468;
  assign n30471 = ~n30466 & ~n36284;
  assign n30472 = n4155 & ~n30446;
  assign n30473 = ~n30461 & n30472;
  assign n30474 = n4155 & n30462;
  assign n30475 = ~n30471 & ~n36285;
  assign n30476 = ~n30463 & ~n30475;
  assign n30477 = ~n3788 & ~n30476;
  assign n30478 = n3788 & ~n30463;
  assign n30479 = ~n30475 & n30478;
  assign n30480 = ~n36165 & ~n29602;
  assign n30481 = ~n29602 & ~n29813;
  assign n30482 = ~n36165 & n30481;
  assign n30483 = ~n29813 & n30480;
  assign n30484 = n29045 & ~n36286;
  assign n30485 = n29601 & n30481;
  assign n30486 = n29045 & ~n36165;
  assign n30487 = ~n29602 & n30486;
  assign n30488 = ~n29813 & n30487;
  assign n30489 = ~n29045 & ~n36286;
  assign n30490 = ~n30488 & ~n30489;
  assign n30491 = ~n30484 & ~n30485;
  assign n30492 = ~n30479 & ~n36287;
  assign n30493 = ~n30477 & ~n30492;
  assign n30494 = ~n3473 & ~n30493;
  assign n30495 = n3473 & ~n30477;
  assign n30496 = ~n30492 & n30495;
  assign n30497 = n3473 & n30493;
  assign n30498 = ~n29604 & ~n29607;
  assign n30499 = ~n29607 & ~n29813;
  assign n30500 = ~n29604 & n30499;
  assign n30501 = ~n29813 & n30498;
  assign n30502 = n29037 & ~n36289;
  assign n30503 = n29605 & n30499;
  assign n30504 = n29037 & ~n29607;
  assign n30505 = ~n29604 & n30504;
  assign n30506 = ~n29813 & n30505;
  assign n30507 = ~n29037 & ~n36289;
  assign n30508 = ~n30506 & ~n30507;
  assign n30509 = ~n30502 & ~n30503;
  assign n30510 = ~n36288 & ~n36290;
  assign n30511 = ~n30494 & ~n30510;
  assign n30512 = ~n3140 & ~n30511;
  assign n30513 = n3140 & ~n30494;
  assign n30514 = ~n30510 & n30513;
  assign n30515 = ~n36166 & ~n29613;
  assign n30516 = ~n29613 & ~n29813;
  assign n30517 = ~n36166 & n30516;
  assign n30518 = ~n29813 & n30515;
  assign n30519 = n29029 & ~n36291;
  assign n30520 = n29612 & n30516;
  assign n30521 = n29029 & ~n36166;
  assign n30522 = ~n29613 & n30521;
  assign n30523 = ~n29813 & n30522;
  assign n30524 = ~n29029 & ~n36291;
  assign n30525 = ~n30523 & ~n30524;
  assign n30526 = ~n30519 & ~n30520;
  assign n30527 = ~n30514 & ~n36292;
  assign n30528 = ~n30512 & ~n30527;
  assign n30529 = ~n2855 & ~n30528;
  assign n30530 = ~n29615 & ~n29630;
  assign n30531 = ~n29813 & n30530;
  assign n30532 = ~n36168 & ~n30531;
  assign n30533 = n36168 & ~n29630;
  assign n30534 = ~n29615 & n30533;
  assign n30535 = n36168 & n30531;
  assign n30536 = ~n29813 & n30534;
  assign n30537 = ~n30532 & ~n36293;
  assign n30538 = n2855 & ~n30512;
  assign n30539 = ~n30527 & n30538;
  assign n30540 = n2855 & n30528;
  assign n30541 = ~n30537 & ~n36294;
  assign n30542 = ~n30529 & ~n30541;
  assign n30543 = ~n2556 & ~n30542;
  assign n30544 = n2556 & ~n30529;
  assign n30545 = ~n30541 & n30544;
  assign n30546 = ~n36169 & ~n29636;
  assign n30547 = ~n29636 & ~n29813;
  assign n30548 = ~n36169 & n30547;
  assign n30549 = ~n29813 & n30546;
  assign n30550 = n29021 & ~n36295;
  assign n30551 = n29635 & n30547;
  assign n30552 = n29021 & ~n36169;
  assign n30553 = ~n29636 & n30552;
  assign n30554 = ~n29813 & n30553;
  assign n30555 = ~n29021 & ~n36295;
  assign n30556 = ~n30554 & ~n30555;
  assign n30557 = ~n30550 & ~n30551;
  assign n30558 = ~n30545 & ~n36296;
  assign n30559 = ~n30543 & ~n30558;
  assign n30560 = ~n2301 & ~n30559;
  assign n30561 = n2301 & ~n30543;
  assign n30562 = ~n30558 & n30561;
  assign n30563 = n2301 & n30559;
  assign n30564 = ~n29638 & ~n29641;
  assign n30565 = ~n29641 & ~n29813;
  assign n30566 = ~n29638 & n30565;
  assign n30567 = ~n29813 & n30564;
  assign n30568 = n29013 & ~n36298;
  assign n30569 = n29639 & n30565;
  assign n30570 = n29013 & ~n29641;
  assign n30571 = ~n29638 & n30570;
  assign n30572 = ~n29813 & n30571;
  assign n30573 = ~n29013 & ~n36298;
  assign n30574 = ~n30572 & ~n30573;
  assign n30575 = ~n30568 & ~n30569;
  assign n30576 = ~n36297 & ~n36299;
  assign n30577 = ~n30560 & ~n30576;
  assign n30578 = ~n2038 & ~n30577;
  assign n30579 = n2038 & ~n30560;
  assign n30580 = ~n30576 & n30579;
  assign n30581 = ~n36170 & ~n29647;
  assign n30582 = ~n29647 & ~n29813;
  assign n30583 = ~n36170 & n30582;
  assign n30584 = ~n29813 & n30581;
  assign n30585 = n29005 & ~n36300;
  assign n30586 = n29646 & n30582;
  assign n30587 = n29005 & ~n36170;
  assign n30588 = ~n29647 & n30587;
  assign n30589 = ~n29813 & n30588;
  assign n30590 = ~n29005 & ~n36300;
  assign n30591 = ~n30589 & ~n30590;
  assign n30592 = ~n30585 & ~n30586;
  assign n30593 = ~n30580 & ~n36301;
  assign n30594 = ~n30578 & ~n30593;
  assign n30595 = ~n1812 & ~n30594;
  assign n30596 = ~n29649 & ~n29664;
  assign n30597 = ~n29813 & n30596;
  assign n30598 = ~n36172 & ~n30597;
  assign n30599 = n36172 & ~n29664;
  assign n30600 = ~n29649 & n30599;
  assign n30601 = n36172 & n30597;
  assign n30602 = ~n29813 & n30600;
  assign n30603 = ~n30598 & ~n36302;
  assign n30604 = n1812 & ~n30578;
  assign n30605 = ~n30593 & n30604;
  assign n30606 = n1812 & n30594;
  assign n30607 = ~n30603 & ~n36303;
  assign n30608 = ~n30595 & ~n30607;
  assign n30609 = ~n1582 & ~n30608;
  assign n30610 = n1582 & ~n30595;
  assign n30611 = ~n30607 & n30610;
  assign n30612 = ~n36173 & ~n29670;
  assign n30613 = ~n29670 & ~n29813;
  assign n30614 = ~n36173 & n30613;
  assign n30615 = ~n29813 & n30612;
  assign n30616 = n28997 & ~n36304;
  assign n30617 = n29669 & n30613;
  assign n30618 = n28997 & ~n36173;
  assign n30619 = ~n29670 & n30618;
  assign n30620 = ~n29813 & n30619;
  assign n30621 = ~n28997 & ~n36304;
  assign n30622 = ~n30620 & ~n30621;
  assign n30623 = ~n30616 & ~n30617;
  assign n30624 = ~n30611 & ~n36305;
  assign n30625 = ~n30609 & ~n30624;
  assign n30626 = ~n1388 & ~n30625;
  assign n30627 = n1388 & ~n30609;
  assign n30628 = ~n30624 & n30627;
  assign n30629 = n1388 & n30625;
  assign n30630 = ~n29672 & ~n29675;
  assign n30631 = ~n29675 & ~n29813;
  assign n30632 = ~n29672 & n30631;
  assign n30633 = ~n29813 & n30630;
  assign n30634 = n28989 & ~n36307;
  assign n30635 = n29673 & n30631;
  assign n30636 = n28989 & ~n29675;
  assign n30637 = ~n29672 & n30636;
  assign n30638 = ~n29813 & n30637;
  assign n30639 = ~n28989 & ~n36307;
  assign n30640 = ~n30638 & ~n30639;
  assign n30641 = ~n30634 & ~n30635;
  assign n30642 = ~n36306 & ~n36308;
  assign n30643 = ~n30626 & ~n30642;
  assign n30644 = ~n1192 & ~n30643;
  assign n30645 = n1192 & ~n30626;
  assign n30646 = ~n30642 & n30645;
  assign n30647 = ~n36174 & ~n29681;
  assign n30648 = ~n29681 & ~n29813;
  assign n30649 = ~n36174 & n30648;
  assign n30650 = ~n29813 & n30647;
  assign n30651 = n28981 & ~n36309;
  assign n30652 = n29680 & n30648;
  assign n30653 = n28981 & ~n36174;
  assign n30654 = ~n29681 & n30653;
  assign n30655 = ~n29813 & n30654;
  assign n30656 = ~n28981 & ~n36309;
  assign n30657 = ~n30655 & ~n30656;
  assign n30658 = ~n30651 & ~n30652;
  assign n30659 = ~n30646 & ~n36310;
  assign n30660 = ~n30644 & ~n30659;
  assign n30661 = ~n1028 & ~n30660;
  assign n30662 = ~n29683 & ~n29698;
  assign n30663 = ~n29813 & n30662;
  assign n30664 = ~n36176 & ~n30663;
  assign n30665 = n36176 & ~n29698;
  assign n30666 = ~n29683 & n30665;
  assign n30667 = n36176 & n30663;
  assign n30668 = ~n29813 & n30666;
  assign n30669 = ~n30664 & ~n36311;
  assign n30670 = n1028 & ~n30644;
  assign n30671 = ~n30659 & n30670;
  assign n30672 = n1028 & n30660;
  assign n30673 = ~n30669 & ~n36312;
  assign n30674 = ~n30661 & ~n30673;
  assign n30675 = ~n866 & ~n30674;
  assign n30676 = n866 & ~n30661;
  assign n30677 = ~n30673 & n30676;
  assign n30678 = ~n36177 & ~n29704;
  assign n30679 = ~n29704 & ~n29813;
  assign n30680 = ~n36177 & n30679;
  assign n30681 = ~n29813 & n30678;
  assign n30682 = n28973 & ~n36313;
  assign n30683 = n29703 & n30679;
  assign n30684 = n28973 & ~n36177;
  assign n30685 = ~n29704 & n30684;
  assign n30686 = ~n29813 & n30685;
  assign n30687 = ~n28973 & ~n36313;
  assign n30688 = ~n30686 & ~n30687;
  assign n30689 = ~n30682 & ~n30683;
  assign n30690 = ~n30677 & ~n36314;
  assign n30691 = ~n30675 & ~n30690;
  assign n30692 = ~n730 & ~n30691;
  assign n30693 = n730 & ~n30675;
  assign n30694 = ~n30690 & n30693;
  assign n30695 = n730 & n30691;
  assign n30696 = ~n29706 & ~n29709;
  assign n30697 = ~n29709 & ~n29813;
  assign n30698 = ~n29706 & n30697;
  assign n30699 = ~n29813 & n30696;
  assign n30700 = n28965 & ~n36316;
  assign n30701 = n29707 & n30697;
  assign n30702 = n28965 & ~n29709;
  assign n30703 = ~n29706 & n30702;
  assign n30704 = ~n29813 & n30703;
  assign n30705 = ~n28965 & ~n36316;
  assign n30706 = ~n30704 & ~n30705;
  assign n30707 = ~n30700 & ~n30701;
  assign n30708 = ~n36315 & ~n36317;
  assign n30709 = ~n30692 & ~n30708;
  assign n30710 = ~n602 & ~n30709;
  assign n30711 = n602 & ~n30692;
  assign n30712 = ~n30708 & n30711;
  assign n30713 = ~n36178 & ~n29715;
  assign n30714 = ~n29715 & ~n29813;
  assign n30715 = ~n36178 & n30714;
  assign n30716 = ~n29813 & n30713;
  assign n30717 = n28957 & ~n36318;
  assign n30718 = n29714 & n30714;
  assign n30719 = n28957 & ~n36178;
  assign n30720 = ~n29715 & n30719;
  assign n30721 = ~n29813 & n30720;
  assign n30722 = ~n28957 & ~n36318;
  assign n30723 = ~n30721 & ~n30722;
  assign n30724 = ~n30717 & ~n30718;
  assign n30725 = ~n30712 & ~n36319;
  assign n30726 = ~n30710 & ~n30725;
  assign n30727 = ~n497 & ~n30726;
  assign n30728 = ~n29717 & ~n29732;
  assign n30729 = ~n29813 & n30728;
  assign n30730 = ~n36180 & ~n30729;
  assign n30731 = n36180 & ~n29732;
  assign n30732 = ~n29717 & n30731;
  assign n30733 = n36180 & n30729;
  assign n30734 = ~n29813 & n30732;
  assign n30735 = ~n30730 & ~n36320;
  assign n30736 = n497 & ~n30710;
  assign n30737 = ~n30725 & n30736;
  assign n30738 = n497 & n30726;
  assign n30739 = ~n30735 & ~n36321;
  assign n30740 = ~n30727 & ~n30739;
  assign n30741 = ~n403 & ~n30740;
  assign n30742 = n403 & ~n30727;
  assign n30743 = ~n30739 & n30742;
  assign n30744 = ~n36181 & ~n29738;
  assign n30745 = ~n29738 & ~n29813;
  assign n30746 = ~n36181 & n30745;
  assign n30747 = ~n29813 & n30744;
  assign n30748 = n28949 & ~n36322;
  assign n30749 = n29737 & n30745;
  assign n30750 = n28949 & ~n36181;
  assign n30751 = ~n29738 & n30750;
  assign n30752 = ~n29813 & n30751;
  assign n30753 = ~n28949 & ~n36322;
  assign n30754 = ~n30752 & ~n30753;
  assign n30755 = ~n30748 & ~n30749;
  assign n30756 = ~n30743 & ~n36323;
  assign n30757 = ~n30741 & ~n30756;
  assign n30758 = ~n330 & ~n30757;
  assign n30759 = n330 & ~n30741;
  assign n30760 = ~n30756 & n30759;
  assign n30761 = n330 & n30757;
  assign n30762 = ~n29740 & ~n29743;
  assign n30763 = ~n29743 & ~n29813;
  assign n30764 = ~n29740 & n30763;
  assign n30765 = ~n29813 & n30762;
  assign n30766 = n28941 & ~n36325;
  assign n30767 = n29741 & n30763;
  assign n30768 = n28941 & ~n29743;
  assign n30769 = ~n29740 & n30768;
  assign n30770 = ~n29813 & n30769;
  assign n30771 = ~n28941 & ~n36325;
  assign n30772 = ~n30770 & ~n30771;
  assign n30773 = ~n30766 & ~n30767;
  assign n30774 = ~n36324 & ~n36326;
  assign n30775 = ~n30758 & ~n30774;
  assign n30776 = ~n271 & ~n30775;
  assign n30777 = n271 & ~n30758;
  assign n30778 = ~n30774 & n30777;
  assign n30779 = ~n36182 & ~n29749;
  assign n30780 = ~n29813 & n30779;
  assign n30781 = n28933 & ~n30780;
  assign n30782 = ~n28933 & n30780;
  assign n30783 = n28933 & ~n36182;
  assign n30784 = ~n29749 & n30783;
  assign n30785 = ~n29813 & n30784;
  assign n30786 = ~n28933 & ~n30780;
  assign n30787 = ~n30785 & ~n30786;
  assign n30788 = ~n30781 & ~n30782;
  assign n30789 = ~n30778 & ~n36327;
  assign n30790 = ~n30776 & ~n30789;
  assign n30791 = ~n217 & ~n30790;
  assign n30792 = ~n29751 & ~n29753;
  assign n30793 = ~n29813 & n30792;
  assign n30794 = n36184 & ~n30793;
  assign n30795 = ~n29751 & ~n36184;
  assign n30796 = ~n29753 & n30795;
  assign n30797 = ~n36184 & n30793;
  assign n30798 = ~n29813 & n30796;
  assign n30799 = n36184 & n30793;
  assign n30800 = ~n36184 & ~n30793;
  assign n30801 = ~n30799 & ~n30800;
  assign n30802 = ~n30794 & ~n36328;
  assign n30803 = n217 & ~n30776;
  assign n30804 = ~n30789 & n30803;
  assign n30805 = n217 & n30790;
  assign n30806 = n36329 & ~n36330;
  assign n30807 = ~n30791 & ~n30806;
  assign n30808 = ~n198 & ~n30807;
  assign n30809 = n198 & ~n30791;
  assign n30810 = ~n30806 & n30809;
  assign n30811 = ~n36192 & ~n30810;
  assign n30812 = ~n30808 & ~n30811;
  assign n30813 = ~n29773 & ~n29775;
  assign n30814 = ~n29813 & n30813;
  assign n30815 = ~n36187 & ~n30814;
  assign n30816 = ~n29773 & n36187;
  assign n30817 = ~n29775 & n30816;
  assign n30818 = n36187 & n30814;
  assign n30819 = ~n29813 & n30817;
  assign n30820 = ~n30815 & ~n36331;
  assign n30821 = ~n29789 & ~n29797;
  assign n30822 = ~n29797 & ~n29813;
  assign n30823 = ~n29789 & n30822;
  assign n30824 = ~n29813 & n30821;
  assign n30825 = ~n36190 & ~n36332;
  assign n30826 = ~n30820 & n30825;
  assign n30827 = ~n30812 & n30826;
  assign n30828 = n193 & ~n30827;
  assign n30829 = ~n30808 & n30820;
  assign n30830 = ~n30811 & n30829;
  assign n30831 = n30812 & n30820;
  assign n30832 = n29789 & ~n30822;
  assign n30833 = ~n193 & ~n30821;
  assign n30834 = ~n30832 & n30833;
  assign n30835 = ~n36333 & ~n30834;
  assign n30836 = ~n30828 & n30835;
  assign n30837 = ~n30808 & ~n30810;
  assign n30838 = ~n30836 & n30837;
  assign n30839 = ~n36192 & ~n30838;
  assign n30840 = n36192 & ~n30810;
  assign n30841 = ~n30808 & n30840;
  assign n30842 = n36192 & n30838;
  assign n30843 = ~n30836 & n30841;
  assign n30844 = ~n30839 & ~n36334;
  assign n30845 = ~n193 & ~n30844;
  assign n30846 = ~n30791 & ~n36330;
  assign n30847 = ~n30836 & n30846;
  assign n30848 = ~n36329 & ~n30847;
  assign n30849 = n36329 & n30847;
  assign n30850 = n36329 & ~n30847;
  assign n30851 = ~n30791 & ~n36329;
  assign n30852 = ~n36330 & n30851;
  assign n30853 = ~n30836 & n30852;
  assign n30854 = ~n30850 & ~n30853;
  assign n30855 = ~n30848 & ~n30849;
  assign n30856 = n198 & n36335;
  assign n30857 = ~n198 & ~n36335;
  assign n30858 = ~n30776 & ~n30778;
  assign n30859 = ~n30836 & n30858;
  assign n30860 = ~n36327 & n30859;
  assign n30861 = n36327 & ~n30859;
  assign n30862 = ~n36327 & ~n30859;
  assign n30863 = ~n30778 & n36327;
  assign n30864 = ~n30776 & n30863;
  assign n30865 = ~n30836 & n30864;
  assign n30866 = ~n30862 & ~n30865;
  assign n30867 = ~n30860 & ~n30861;
  assign n30868 = n217 & n36336;
  assign n30869 = ~n30692 & ~n36315;
  assign n30870 = ~n30836 & n30869;
  assign n30871 = ~n36317 & ~n30870;
  assign n30872 = ~n30692 & n36317;
  assign n30873 = ~n36315 & n30872;
  assign n30874 = n36317 & n30870;
  assign n30875 = ~n30836 & n30873;
  assign n30876 = ~n30871 & ~n36337;
  assign n30877 = ~n602 & ~n30876;
  assign n30878 = ~n30661 & ~n36312;
  assign n30879 = ~n30661 & ~n30836;
  assign n30880 = ~n36312 & n30879;
  assign n30881 = ~n30836 & n30878;
  assign n30882 = n30669 & ~n36338;
  assign n30883 = n30673 & n30879;
  assign n30884 = ~n30669 & ~n36338;
  assign n30885 = ~n30661 & n30669;
  assign n30886 = ~n36312 & n30885;
  assign n30887 = ~n30836 & n30886;
  assign n30888 = ~n30884 & ~n30887;
  assign n30889 = ~n30882 & ~n30883;
  assign n30890 = ~n866 & ~n36339;
  assign n30891 = ~n30626 & ~n36306;
  assign n30892 = ~n30836 & n30891;
  assign n30893 = ~n36308 & ~n30892;
  assign n30894 = ~n30626 & n36308;
  assign n30895 = ~n36306 & n30894;
  assign n30896 = n36308 & n30892;
  assign n30897 = ~n30836 & n30895;
  assign n30898 = ~n30893 & ~n36340;
  assign n30899 = ~n1192 & ~n30898;
  assign n30900 = ~n30595 & ~n36303;
  assign n30901 = ~n30595 & ~n30836;
  assign n30902 = ~n36303 & n30901;
  assign n30903 = ~n30836 & n30900;
  assign n30904 = n30603 & ~n36341;
  assign n30905 = n30607 & n30901;
  assign n30906 = ~n30603 & ~n36341;
  assign n30907 = ~n30595 & n30603;
  assign n30908 = ~n36303 & n30907;
  assign n30909 = ~n30836 & n30908;
  assign n30910 = ~n30906 & ~n30909;
  assign n30911 = ~n30904 & ~n30905;
  assign n30912 = ~n1582 & ~n36342;
  assign n30913 = ~n30560 & ~n36297;
  assign n30914 = ~n30836 & n30913;
  assign n30915 = ~n36299 & ~n30914;
  assign n30916 = ~n30560 & n36299;
  assign n30917 = ~n36297 & n30916;
  assign n30918 = n36299 & n30914;
  assign n30919 = ~n30836 & n30917;
  assign n30920 = ~n30915 & ~n36343;
  assign n30921 = ~n2038 & ~n30920;
  assign n30922 = ~n30529 & ~n36294;
  assign n30923 = ~n30529 & ~n30836;
  assign n30924 = ~n36294 & n30923;
  assign n30925 = ~n30836 & n30922;
  assign n30926 = n30537 & ~n36344;
  assign n30927 = n30541 & n30923;
  assign n30928 = ~n30537 & ~n36344;
  assign n30929 = ~n30529 & n30537;
  assign n30930 = ~n36294 & n30929;
  assign n30931 = ~n30836 & n30930;
  assign n30932 = ~n30928 & ~n30931;
  assign n30933 = ~n30926 & ~n30927;
  assign n30934 = ~n2556 & ~n36345;
  assign n30935 = ~n30494 & ~n36288;
  assign n30936 = ~n30836 & n30935;
  assign n30937 = ~n36290 & ~n30936;
  assign n30938 = ~n30494 & n36290;
  assign n30939 = ~n36288 & n30938;
  assign n30940 = n36290 & n30936;
  assign n30941 = ~n30836 & n30939;
  assign n30942 = ~n30937 & ~n36346;
  assign n30943 = ~n3140 & ~n30942;
  assign n30944 = ~n30463 & ~n36285;
  assign n30945 = ~n30463 & ~n30836;
  assign n30946 = ~n36285 & n30945;
  assign n30947 = ~n30836 & n30944;
  assign n30948 = n30471 & ~n36347;
  assign n30949 = n30475 & n30945;
  assign n30950 = ~n30471 & ~n36347;
  assign n30951 = ~n30463 & n30471;
  assign n30952 = ~n36285 & n30951;
  assign n30953 = ~n30836 & n30952;
  assign n30954 = ~n30950 & ~n30953;
  assign n30955 = ~n30948 & ~n30949;
  assign n30956 = ~n3788 & ~n36348;
  assign n30957 = ~n30428 & ~n36279;
  assign n30958 = ~n30836 & n30957;
  assign n30959 = ~n36281 & ~n30958;
  assign n30960 = ~n30428 & n36281;
  assign n30961 = ~n36279 & n30960;
  assign n30962 = n36281 & n30958;
  assign n30963 = ~n30836 & n30961;
  assign n30964 = ~n30959 & ~n36349;
  assign n30965 = ~n4508 & ~n30964;
  assign n30966 = ~n30397 & ~n36276;
  assign n30967 = ~n30397 & ~n30836;
  assign n30968 = ~n36276 & n30967;
  assign n30969 = ~n30836 & n30966;
  assign n30970 = n30405 & ~n36350;
  assign n30971 = n30409 & n30967;
  assign n30972 = ~n30405 & ~n36350;
  assign n30973 = ~n30397 & n30405;
  assign n30974 = ~n36276 & n30973;
  assign n30975 = ~n30836 & n30974;
  assign n30976 = ~n30972 & ~n30975;
  assign n30977 = ~n30970 & ~n30971;
  assign n30978 = ~n5278 & ~n36351;
  assign n30979 = ~n30362 & ~n36270;
  assign n30980 = ~n30836 & n30979;
  assign n30981 = ~n36272 & ~n30980;
  assign n30982 = ~n30362 & n36272;
  assign n30983 = ~n36270 & n30982;
  assign n30984 = n36272 & n30980;
  assign n30985 = ~n30836 & n30983;
  assign n30986 = ~n30981 & ~n36352;
  assign n30987 = ~n6117 & ~n30986;
  assign n30988 = ~n30331 & ~n36267;
  assign n30989 = ~n30331 & ~n30836;
  assign n30990 = ~n36267 & n30989;
  assign n30991 = ~n30836 & n30988;
  assign n30992 = n30339 & ~n36353;
  assign n30993 = n30343 & n30989;
  assign n30994 = ~n30339 & ~n36353;
  assign n30995 = ~n30331 & n30339;
  assign n30996 = ~n36267 & n30995;
  assign n30997 = ~n30836 & n30996;
  assign n30998 = ~n30994 & ~n30997;
  assign n30999 = ~n30992 & ~n30993;
  assign n31000 = ~n7015 & ~n36354;
  assign n31001 = ~n30296 & ~n36261;
  assign n31002 = ~n30836 & n31001;
  assign n31003 = ~n36263 & ~n31002;
  assign n31004 = ~n30296 & n36263;
  assign n31005 = ~n36261 & n31004;
  assign n31006 = n36263 & n31002;
  assign n31007 = ~n30836 & n31005;
  assign n31008 = ~n31003 & ~n36355;
  assign n31009 = ~n7975 & ~n31008;
  assign n31010 = ~n30265 & ~n36258;
  assign n31011 = ~n30265 & ~n30836;
  assign n31012 = ~n36258 & n31011;
  assign n31013 = ~n30836 & n31010;
  assign n31014 = n30273 & ~n36356;
  assign n31015 = n30277 & n31011;
  assign n31016 = ~n30273 & ~n36356;
  assign n31017 = ~n30265 & n30273;
  assign n31018 = ~n36258 & n31017;
  assign n31019 = ~n30836 & n31018;
  assign n31020 = ~n31016 & ~n31019;
  assign n31021 = ~n31014 & ~n31015;
  assign n31022 = ~n8998 & ~n36357;
  assign n31023 = ~n30230 & ~n36252;
  assign n31024 = ~n30836 & n31023;
  assign n31025 = ~n36254 & ~n31024;
  assign n31026 = ~n30230 & n36254;
  assign n31027 = ~n36252 & n31026;
  assign n31028 = n36254 & n31024;
  assign n31029 = ~n30836 & n31027;
  assign n31030 = ~n31025 & ~n36358;
  assign n31031 = ~n10086 & ~n31030;
  assign n31032 = ~n30199 & ~n36249;
  assign n31033 = ~n30199 & ~n30836;
  assign n31034 = ~n36249 & n31033;
  assign n31035 = ~n30836 & n31032;
  assign n31036 = n30207 & ~n36359;
  assign n31037 = n30211 & n31033;
  assign n31038 = ~n30207 & ~n36359;
  assign n31039 = ~n30199 & n30207;
  assign n31040 = ~n36249 & n31039;
  assign n31041 = ~n30836 & n31040;
  assign n31042 = ~n31038 & ~n31041;
  assign n31043 = ~n31036 & ~n31037;
  assign n31044 = ~n11229 & ~n36360;
  assign n31045 = ~n30163 & ~n36242;
  assign n31046 = ~n30836 & n31045;
  assign n31047 = ~n36245 & ~n31046;
  assign n31048 = ~n30163 & n36245;
  assign n31049 = ~n36242 & n31048;
  assign n31050 = n36245 & n31046;
  assign n31051 = ~n30836 & n31049;
  assign n31052 = ~n31047 & ~n36361;
  assign n31053 = ~n12442 & ~n31052;
  assign n31054 = ~n30129 & ~n36237;
  assign n31055 = ~n30129 & ~n30836;
  assign n31056 = ~n36237 & n31055;
  assign n31057 = ~n30836 & n31054;
  assign n31058 = n36239 & ~n36362;
  assign n31059 = n30144 & n31055;
  assign n31060 = ~n36239 & n36362;
  assign n31061 = ~n36239 & ~n36362;
  assign n31062 = ~n30129 & n36239;
  assign n31063 = ~n36237 & n31062;
  assign n31064 = ~n30836 & n31063;
  assign n31065 = ~n31061 & ~n31064;
  assign n31066 = ~n31058 & ~n36363;
  assign n31067 = ~n13704 & ~n36364;
  assign n31068 = ~n30093 & ~n36231;
  assign n31069 = ~n30836 & n31068;
  assign n31070 = ~n36234 & n31069;
  assign n31071 = n36234 & ~n31069;
  assign n31072 = ~n36234 & ~n31069;
  assign n31073 = ~n30093 & n36234;
  assign n31074 = ~n36231 & n31073;
  assign n31075 = n36234 & n31069;
  assign n31076 = ~n30836 & n31074;
  assign n31077 = ~n31072 & ~n36365;
  assign n31078 = ~n31070 & ~n31071;
  assign n31079 = ~n15033 & ~n36366;
  assign n31080 = ~n30062 & ~n36227;
  assign n31081 = ~n30062 & ~n30836;
  assign n31082 = ~n36227 & n31081;
  assign n31083 = ~n30836 & n31080;
  assign n31084 = n30073 & ~n36367;
  assign n31085 = n30074 & n31081;
  assign n31086 = ~n30073 & n36367;
  assign n31087 = ~n30073 & ~n36367;
  assign n31088 = ~n30062 & n30073;
  assign n31089 = ~n36227 & n31088;
  assign n31090 = ~n30836 & n31089;
  assign n31091 = ~n31087 & ~n31090;
  assign n31092 = ~n31084 & ~n36368;
  assign n31093 = ~n16428 & ~n36369;
  assign n31094 = ~n30026 & ~n36221;
  assign n31095 = ~n30836 & n31094;
  assign n31096 = ~n36224 & ~n31095;
  assign n31097 = ~n30026 & n36224;
  assign n31098 = ~n36221 & n31097;
  assign n31099 = n36224 & n31095;
  assign n31100 = ~n30836 & n31098;
  assign n31101 = ~n31096 & ~n36370;
  assign n31102 = ~n17885 & ~n31101;
  assign n31103 = ~n29992 & ~n36216;
  assign n31104 = ~n29992 & ~n30836;
  assign n31105 = ~n36216 & n31104;
  assign n31106 = ~n30836 & n31103;
  assign n31107 = ~n36218 & ~n36371;
  assign n31108 = n30007 & n31104;
  assign n31109 = n36218 & n36371;
  assign n31110 = n36218 & ~n36371;
  assign n31111 = ~n29992 & ~n36218;
  assign n31112 = ~n36216 & n31111;
  assign n31113 = ~n30836 & n31112;
  assign n31114 = ~n31110 & ~n31113;
  assign n31115 = ~n31107 & ~n36372;
  assign n31116 = ~n19401 & ~n36373;
  assign n31117 = ~n29958 & ~n36211;
  assign n31118 = ~n30836 & n31117;
  assign n31119 = n36213 & ~n31118;
  assign n31120 = ~n29958 & ~n36213;
  assign n31121 = ~n36211 & n31120;
  assign n31122 = ~n36213 & n31118;
  assign n31123 = ~n30836 & n31121;
  assign n31124 = n36213 & n31118;
  assign n31125 = ~n36213 & ~n31118;
  assign n31126 = ~n31124 & ~n31125;
  assign n31127 = ~n31119 & ~n36374;
  assign n31128 = ~n20986 & n36375;
  assign n31129 = ~n29925 & ~n36207;
  assign n31130 = ~n30836 & n31129;
  assign n31131 = ~n36208 & ~n31130;
  assign n31132 = ~n29925 & n36208;
  assign n31133 = ~n36207 & n31132;
  assign n31134 = n36208 & n31130;
  assign n31135 = ~n30836 & n31133;
  assign n31136 = n36208 & ~n31130;
  assign n31137 = ~n36208 & n31130;
  assign n31138 = ~n31136 & ~n31137;
  assign n31139 = ~n31131 & ~n36376;
  assign n31140 = ~n22625 & n36377;
  assign n31141 = ~n29891 & ~n36202;
  assign n31142 = ~n30836 & n31141;
  assign n31143 = ~n36204 & n31142;
  assign n31144 = n36204 & ~n31142;
  assign n31145 = ~n36204 & ~n31142;
  assign n31146 = ~n29891 & n36204;
  assign n31147 = ~n36202 & n31146;
  assign n31148 = ~n30836 & n31147;
  assign n31149 = ~n31145 & ~n31148;
  assign n31150 = ~n31143 & ~n31144;
  assign n31151 = ~n24331 & ~n36378;
  assign n31152 = ~n29861 & ~n36198;
  assign n31153 = ~n30836 & n31152;
  assign n31154 = n29871 & ~n31153;
  assign n31155 = ~n29871 & n31153;
  assign n31156 = ~n29861 & n29871;
  assign n31157 = ~n36198 & n31156;
  assign n31158 = n29871 & n31153;
  assign n31159 = ~n30836 & n31157;
  assign n31160 = ~n29871 & ~n31153;
  assign n31161 = ~n36379 & ~n31160;
  assign n31162 = ~n31154 & ~n31155;
  assign n31163 = n26098 & n36380;
  assign n31164 = ~n26098 & ~n36380;
  assign n31165 = ~n29846 & ~n29848;
  assign n31166 = ~n30836 & n31165;
  assign n31167 = ~n29858 & ~n31166;
  assign n31168 = ~n29848 & n29858;
  assign n31169 = ~n29846 & n31168;
  assign n31170 = n29858 & n31166;
  assign n31171 = ~n30836 & n31169;
  assign n31172 = ~n31167 & ~n36381;
  assign n31173 = n27055 & n31172;
  assign n31174 = ~pi0  & ~pi1 ;
  assign n31175 = ~pi2  & ~n31174;
  assign n31176 = pi2  & ~n30834;
  assign n31177 = ~n36333 & n31176;
  assign n31178 = pi2  & n30836;
  assign n31179 = ~n30828 & n31177;
  assign n31180 = ~n31175 & ~n36382;
  assign n31181 = n29813 & ~n31180;
  assign n31182 = ~pi2  & ~n30836;
  assign n31183 = ~pi3  & n31182;
  assign n31184 = n29827 & ~n30836;
  assign n31185 = pi3  & ~n31182;
  assign n31186 = ~n36383 & ~n31185;
  assign n31187 = ~n29813 & n31180;
  assign n31188 = ~n31186 & ~n31187;
  assign n31189 = n31180 & ~n36383;
  assign n31190 = n31180 & n31186;
  assign n31191 = ~n31185 & n31189;
  assign n31192 = ~n31180 & ~n31186;
  assign n31193 = ~n29813 & ~n31192;
  assign n31194 = ~n36384 & ~n31193;
  assign n31195 = n29813 & ~n36384;
  assign n31196 = ~n31192 & ~n31195;
  assign n31197 = ~n31181 & ~n31188;
  assign n31198 = ~n28917 & ~n36385;
  assign n31199 = ~n29813 & ~n30834;
  assign n31200 = ~n36333 & n31199;
  assign n31201 = ~n29813 & n30836;
  assign n31202 = ~n30828 & n31200;
  assign n31203 = ~n36383 & ~n36386;
  assign n31204 = pi4  & ~n31203;
  assign n31205 = ~pi4  & ~n36386;
  assign n31206 = ~pi4  & n31203;
  assign n31207 = ~n36383 & n31205;
  assign n31208 = ~n31204 & ~n36387;
  assign n31209 = ~n31198 & n31208;
  assign n31210 = ~n29833 & ~n36195;
  assign n31211 = ~n30836 & n31210;
  assign n31212 = n29838 & ~n31211;
  assign n31213 = ~n29838 & n31210;
  assign n31214 = ~n29838 & n31211;
  assign n31215 = ~n30836 & n31213;
  assign n31216 = ~n31212 & ~n36388;
  assign n31217 = n27931 & n31216;
  assign n31218 = n28917 & n36385;
  assign n31219 = ~n31217 & ~n31218;
  assign n31220 = ~n31209 & n31219;
  assign n31221 = ~n27931 & ~n31216;
  assign n31222 = ~n27055 & ~n31172;
  assign n31223 = ~n31221 & ~n31222;
  assign n31224 = ~n31220 & n31223;
  assign n31225 = ~n36385 & ~n31208;
  assign n31226 = n28917 & ~n31225;
  assign n31227 = n36385 & n31208;
  assign n31228 = ~n31216 & ~n31227;
  assign n31229 = ~n31226 & n31228;
  assign n31230 = n27931 & ~n31229;
  assign n31231 = ~n31209 & ~n31218;
  assign n31232 = ~n31226 & ~n31227;
  assign n31233 = n31216 & ~n36389;
  assign n31234 = ~n31172 & ~n31233;
  assign n31235 = ~n31172 & ~n31230;
  assign n31236 = ~n31233 & n31235;
  assign n31237 = ~n31230 & n31234;
  assign n31238 = n27055 & ~n36390;
  assign n31239 = ~n31221 & ~n36389;
  assign n31240 = ~n31217 & ~n31239;
  assign n31241 = ~n31230 & ~n31233;
  assign n31242 = ~n31220 & ~n31221;
  assign n31243 = n31172 & ~n36391;
  assign n31244 = ~n31238 & ~n31243;
  assign n31245 = ~n27055 & n36391;
  assign n31246 = n31172 & ~n31245;
  assign n31247 = n27055 & ~n36391;
  assign n31248 = ~n31246 & ~n31247;
  assign n31249 = ~n31173 & ~n31224;
  assign n31250 = ~n31164 & ~n36392;
  assign n31251 = ~n31163 & ~n31247;
  assign n31252 = ~n31246 & n31251;
  assign n31253 = ~n31164 & ~n31252;
  assign n31254 = ~n36380 & ~n31243;
  assign n31255 = ~n31238 & n31254;
  assign n31256 = n26098 & ~n31255;
  assign n31257 = n36380 & ~n36392;
  assign n31258 = ~n31256 & ~n31257;
  assign n31259 = ~n31163 & ~n31250;
  assign n31260 = ~n25256 & ~n36393;
  assign n31261 = ~n29874 & ~n29876;
  assign n31262 = ~n30836 & n31261;
  assign n31263 = ~n36201 & ~n31262;
  assign n31264 = ~n29876 & n36201;
  assign n31265 = ~n29874 & n31264;
  assign n31266 = n36201 & n31262;
  assign n31267 = ~n30836 & n31265;
  assign n31268 = ~n31263 & ~n36394;
  assign n31269 = ~n31260 & n31268;
  assign n31270 = n24331 & n36378;
  assign n31271 = n25256 & n36393;
  assign n31272 = ~n31270 & ~n31271;
  assign n31273 = ~n31269 & n31272;
  assign n31274 = n25256 & n31268;
  assign n31275 = ~n25256 & ~n31268;
  assign n31276 = n36393 & ~n31275;
  assign n31277 = ~n31257 & ~n31268;
  assign n31278 = ~n31256 & ~n31268;
  assign n31279 = ~n31257 & n31278;
  assign n31280 = ~n31256 & n31277;
  assign n31281 = n25256 & ~n36395;
  assign n31282 = n36393 & n31268;
  assign n31283 = ~n31281 & ~n31282;
  assign n31284 = ~n31269 & ~n31271;
  assign n31285 = ~n31274 & ~n31276;
  assign n31286 = ~n31151 & ~n36396;
  assign n31287 = ~n31270 & ~n31286;
  assign n31288 = ~n36378 & ~n31282;
  assign n31289 = ~n31281 & n31288;
  assign n31290 = n24331 & ~n31289;
  assign n31291 = n36378 & ~n36396;
  assign n31292 = ~n31290 & ~n31291;
  assign n31293 = ~n31151 & ~n31273;
  assign n31294 = ~n23517 & n36397;
  assign n31295 = ~n29908 & ~n29910;
  assign n31296 = ~n30836 & n31295;
  assign n31297 = ~n36206 & ~n31296;
  assign n31298 = ~n29910 & n36206;
  assign n31299 = ~n29908 & n31298;
  assign n31300 = n36206 & n31296;
  assign n31301 = ~n30836 & n31299;
  assign n31302 = ~n31297 & ~n36398;
  assign n31303 = ~n31294 & n31302;
  assign n31304 = n22625 & ~n36377;
  assign n31305 = n23517 & ~n36397;
  assign n31306 = ~n31304 & ~n31305;
  assign n31307 = ~n31303 & n31306;
  assign n31308 = n23517 & n31302;
  assign n31309 = ~n23517 & ~n31302;
  assign n31310 = ~n36397 & ~n31309;
  assign n31311 = ~n31291 & ~n31302;
  assign n31312 = ~n31290 & ~n31302;
  assign n31313 = ~n31291 & n31312;
  assign n31314 = ~n31290 & n31311;
  assign n31315 = n23517 & ~n36399;
  assign n31316 = ~n36397 & n31302;
  assign n31317 = ~n31315 & ~n31316;
  assign n31318 = ~n31303 & ~n31305;
  assign n31319 = ~n31308 & ~n31310;
  assign n31320 = ~n31140 & ~n36400;
  assign n31321 = ~n31304 & ~n31320;
  assign n31322 = n36377 & ~n31316;
  assign n31323 = ~n31315 & n31322;
  assign n31324 = n22625 & ~n31323;
  assign n31325 = ~n36377 & ~n36400;
  assign n31326 = ~n31324 & ~n31325;
  assign n31327 = ~n31140 & ~n31307;
  assign n31328 = ~n21842 & n36401;
  assign n31329 = ~n29941 & ~n29943;
  assign n31330 = ~n30836 & n31329;
  assign n31331 = ~n36210 & ~n31330;
  assign n31332 = ~n29943 & n36210;
  assign n31333 = ~n29941 & n31332;
  assign n31334 = n36210 & n31330;
  assign n31335 = ~n30836 & n31333;
  assign n31336 = ~n31331 & ~n36402;
  assign n31337 = ~n31328 & n31336;
  assign n31338 = n20986 & ~n36375;
  assign n31339 = n21842 & ~n36401;
  assign n31340 = ~n31338 & ~n31339;
  assign n31341 = ~n31337 & n31340;
  assign n31342 = n21842 & n31336;
  assign n31343 = ~n21842 & ~n31336;
  assign n31344 = ~n36401 & ~n31343;
  assign n31345 = ~n31325 & ~n31336;
  assign n31346 = ~n31324 & ~n31336;
  assign n31347 = ~n31325 & n31346;
  assign n31348 = ~n31324 & n31345;
  assign n31349 = n21842 & ~n36403;
  assign n31350 = ~n36401 & n31336;
  assign n31351 = ~n31349 & ~n31350;
  assign n31352 = ~n31337 & ~n31339;
  assign n31353 = ~n31342 & ~n31344;
  assign n31354 = ~n31128 & ~n36404;
  assign n31355 = ~n31338 & ~n31354;
  assign n31356 = n36375 & ~n31350;
  assign n31357 = ~n31349 & n31356;
  assign n31358 = n20986 & ~n31357;
  assign n31359 = ~n36375 & ~n36404;
  assign n31360 = ~n31358 & ~n31359;
  assign n31361 = ~n31128 & ~n31341;
  assign n31362 = ~n20229 & n36405;
  assign n31363 = ~n29975 & ~n29977;
  assign n31364 = ~n30836 & n31363;
  assign n31365 = ~n36215 & ~n31364;
  assign n31366 = ~n29977 & n36215;
  assign n31367 = ~n29975 & n31366;
  assign n31368 = n36215 & n31364;
  assign n31369 = ~n30836 & n31367;
  assign n31370 = ~n31365 & ~n36406;
  assign n31371 = ~n31362 & n31370;
  assign n31372 = n19401 & n36373;
  assign n31373 = n20229 & ~n36405;
  assign n31374 = ~n31372 & ~n31373;
  assign n31375 = ~n31371 & n31374;
  assign n31376 = n20229 & n31370;
  assign n31377 = ~n20229 & ~n31370;
  assign n31378 = ~n36405 & ~n31377;
  assign n31379 = ~n31359 & ~n31370;
  assign n31380 = ~n31358 & ~n31370;
  assign n31381 = ~n31359 & n31380;
  assign n31382 = ~n31358 & n31379;
  assign n31383 = n20229 & ~n36407;
  assign n31384 = ~n36405 & n31370;
  assign n31385 = ~n31383 & ~n31384;
  assign n31386 = ~n31371 & ~n31373;
  assign n31387 = ~n31376 & ~n31378;
  assign n31388 = ~n31116 & ~n36408;
  assign n31389 = ~n31372 & ~n31388;
  assign n31390 = ~n36373 & ~n31384;
  assign n31391 = ~n31383 & n31390;
  assign n31392 = n19401 & ~n31391;
  assign n31393 = n36373 & ~n36408;
  assign n31394 = ~n31392 & ~n31393;
  assign n31395 = ~n31116 & ~n31375;
  assign n31396 = ~n18676 & n36409;
  assign n31397 = ~n30009 & ~n30011;
  assign n31398 = ~n30836 & n31397;
  assign n31399 = ~n36220 & ~n31398;
  assign n31400 = ~n30011 & n36220;
  assign n31401 = ~n30009 & n31400;
  assign n31402 = n36220 & n31398;
  assign n31403 = ~n30836 & n31401;
  assign n31404 = ~n31399 & ~n36410;
  assign n31405 = ~n31396 & n31404;
  assign n31406 = n17885 & n31101;
  assign n31407 = n18676 & ~n36409;
  assign n31408 = ~n31406 & ~n31407;
  assign n31409 = ~n31405 & n31408;
  assign n31410 = n18676 & n31404;
  assign n31411 = ~n18676 & ~n31404;
  assign n31412 = ~n36409 & ~n31411;
  assign n31413 = ~n31393 & ~n31404;
  assign n31414 = ~n31392 & ~n31404;
  assign n31415 = ~n31393 & n31414;
  assign n31416 = ~n31392 & n31413;
  assign n31417 = n18676 & ~n36411;
  assign n31418 = ~n36409 & n31404;
  assign n31419 = ~n31417 & ~n31418;
  assign n31420 = ~n31405 & ~n31407;
  assign n31421 = ~n31410 & ~n31412;
  assign n31422 = ~n31102 & ~n36412;
  assign n31423 = ~n31406 & ~n31422;
  assign n31424 = ~n31101 & ~n31418;
  assign n31425 = ~n31417 & n31424;
  assign n31426 = n17885 & ~n31425;
  assign n31427 = n31101 & ~n36412;
  assign n31428 = ~n31426 & ~n31427;
  assign n31429 = ~n31102 & ~n31409;
  assign n31430 = ~n17187 & n36413;
  assign n31431 = ~n30045 & ~n30047;
  assign n31432 = ~n30836 & n31431;
  assign n31433 = ~n36226 & ~n31432;
  assign n31434 = ~n30047 & n36226;
  assign n31435 = ~n30045 & n31434;
  assign n31436 = n36226 & n31432;
  assign n31437 = ~n30836 & n31435;
  assign n31438 = ~n31433 & ~n36414;
  assign n31439 = ~n31430 & n31438;
  assign n31440 = n16428 & n36369;
  assign n31441 = n17187 & ~n36413;
  assign n31442 = ~n31440 & ~n31441;
  assign n31443 = ~n31439 & n31442;
  assign n31444 = n17187 & n31438;
  assign n31445 = ~n17187 & ~n31438;
  assign n31446 = ~n36413 & ~n31445;
  assign n31447 = ~n31427 & ~n31438;
  assign n31448 = ~n31426 & ~n31438;
  assign n31449 = ~n31427 & n31448;
  assign n31450 = ~n31426 & n31447;
  assign n31451 = n17187 & ~n36415;
  assign n31452 = ~n36413 & n31438;
  assign n31453 = ~n31451 & ~n31452;
  assign n31454 = ~n31439 & ~n31441;
  assign n31455 = ~n31444 & ~n31446;
  assign n31456 = ~n31093 & ~n36416;
  assign n31457 = ~n31440 & ~n31456;
  assign n31458 = ~n36369 & ~n31452;
  assign n31459 = ~n31451 & n31458;
  assign n31460 = n16428 & ~n31459;
  assign n31461 = n36369 & ~n36416;
  assign n31462 = ~n31460 & ~n31461;
  assign n31463 = ~n31093 & ~n31443;
  assign n31464 = ~n15760 & n36417;
  assign n31465 = ~n30076 & ~n30078;
  assign n31466 = ~n30836 & n31465;
  assign n31467 = ~n36230 & ~n31466;
  assign n31468 = ~n30078 & n36230;
  assign n31469 = ~n30076 & n31468;
  assign n31470 = n36230 & n31466;
  assign n31471 = ~n30836 & n31469;
  assign n31472 = ~n31467 & ~n36418;
  assign n31473 = ~n31464 & n31472;
  assign n31474 = n15033 & n36366;
  assign n31475 = n15760 & ~n36417;
  assign n31476 = ~n31474 & ~n31475;
  assign n31477 = ~n31473 & n31476;
  assign n31478 = n15760 & n31472;
  assign n31479 = ~n15760 & ~n31472;
  assign n31480 = ~n36417 & ~n31479;
  assign n31481 = ~n31461 & ~n31472;
  assign n31482 = ~n31460 & ~n31472;
  assign n31483 = ~n31461 & n31482;
  assign n31484 = ~n31460 & n31481;
  assign n31485 = n15760 & ~n36419;
  assign n31486 = ~n36417 & n31472;
  assign n31487 = ~n31485 & ~n31486;
  assign n31488 = ~n31473 & ~n31475;
  assign n31489 = ~n31478 & ~n31480;
  assign n31490 = ~n31079 & ~n36420;
  assign n31491 = ~n31474 & ~n31490;
  assign n31492 = ~n36366 & ~n31486;
  assign n31493 = ~n31485 & n31492;
  assign n31494 = n15033 & ~n31493;
  assign n31495 = n36366 & ~n36420;
  assign n31496 = ~n31494 & ~n31495;
  assign n31497 = ~n31079 & ~n31477;
  assign n31498 = ~n14394 & n36421;
  assign n31499 = ~n30112 & ~n30114;
  assign n31500 = ~n30836 & n31499;
  assign n31501 = ~n36236 & ~n31500;
  assign n31502 = ~n30114 & n36236;
  assign n31503 = ~n30112 & n31502;
  assign n31504 = n36236 & n31500;
  assign n31505 = ~n30836 & n31503;
  assign n31506 = ~n31501 & ~n36422;
  assign n31507 = ~n31498 & n31506;
  assign n31508 = n13704 & n36364;
  assign n31509 = n14394 & ~n36421;
  assign n31510 = ~n31508 & ~n31509;
  assign n31511 = ~n31507 & n31510;
  assign n31512 = n14394 & n31506;
  assign n31513 = ~n14394 & ~n31506;
  assign n31514 = ~n36421 & ~n31513;
  assign n31515 = ~n31495 & ~n31506;
  assign n31516 = ~n31494 & ~n31506;
  assign n31517 = ~n31495 & n31516;
  assign n31518 = ~n31494 & n31515;
  assign n31519 = n14394 & ~n36423;
  assign n31520 = ~n36421 & n31506;
  assign n31521 = ~n31519 & ~n31520;
  assign n31522 = ~n31507 & ~n31509;
  assign n31523 = ~n31512 & ~n31514;
  assign n31524 = ~n31067 & ~n36424;
  assign n31525 = ~n31508 & ~n31524;
  assign n31526 = ~n36364 & ~n31520;
  assign n31527 = ~n31519 & n31526;
  assign n31528 = n13704 & ~n31527;
  assign n31529 = n36364 & ~n36424;
  assign n31530 = ~n31528 & ~n31529;
  assign n31531 = ~n31067 & ~n31511;
  assign n31532 = ~n13099 & n36425;
  assign n31533 = ~n30146 & ~n30148;
  assign n31534 = ~n30836 & n31533;
  assign n31535 = ~n36241 & ~n31534;
  assign n31536 = ~n30148 & n36241;
  assign n31537 = ~n30146 & n31536;
  assign n31538 = n36241 & n31534;
  assign n31539 = ~n30836 & n31537;
  assign n31540 = ~n31535 & ~n36426;
  assign n31541 = ~n31532 & n31540;
  assign n31542 = n12442 & n31052;
  assign n31543 = n13099 & ~n36425;
  assign n31544 = ~n31542 & ~n31543;
  assign n31545 = ~n31541 & n31544;
  assign n31546 = n13099 & n31540;
  assign n31547 = ~n13099 & ~n31540;
  assign n31548 = ~n36425 & ~n31547;
  assign n31549 = ~n31529 & ~n31540;
  assign n31550 = ~n31528 & ~n31540;
  assign n31551 = ~n31529 & n31550;
  assign n31552 = ~n31528 & n31549;
  assign n31553 = n13099 & ~n36427;
  assign n31554 = ~n36425 & n31540;
  assign n31555 = ~n31553 & ~n31554;
  assign n31556 = ~n31541 & ~n31543;
  assign n31557 = ~n31546 & ~n31548;
  assign n31558 = ~n31053 & ~n36428;
  assign n31559 = ~n31542 & ~n31558;
  assign n31560 = ~n31052 & ~n31554;
  assign n31561 = ~n31553 & n31560;
  assign n31562 = n12442 & ~n31561;
  assign n31563 = n31052 & ~n36428;
  assign n31564 = ~n31562 & ~n31563;
  assign n31565 = ~n31053 & ~n31545;
  assign n31566 = ~n11858 & n36429;
  assign n31567 = ~n30182 & ~n30184;
  assign n31568 = ~n30836 & n31567;
  assign n31569 = ~n36247 & ~n31568;
  assign n31570 = ~n30184 & n36247;
  assign n31571 = ~n30182 & n31570;
  assign n31572 = n36247 & n31568;
  assign n31573 = ~n30836 & n31571;
  assign n31574 = ~n31569 & ~n36430;
  assign n31575 = ~n31566 & n31574;
  assign n31576 = n11229 & n36360;
  assign n31577 = n11858 & ~n36429;
  assign n31578 = ~n31576 & ~n31577;
  assign n31579 = ~n31575 & n31578;
  assign n31580 = n11858 & n31574;
  assign n31581 = ~n11858 & ~n31574;
  assign n31582 = ~n36429 & ~n31581;
  assign n31583 = ~n31563 & ~n31574;
  assign n31584 = ~n31562 & ~n31574;
  assign n31585 = ~n31563 & n31584;
  assign n31586 = ~n31562 & n31583;
  assign n31587 = n11858 & ~n36431;
  assign n31588 = ~n36429 & n31574;
  assign n31589 = ~n31587 & ~n31588;
  assign n31590 = ~n31575 & ~n31577;
  assign n31591 = ~n31580 & ~n31582;
  assign n31592 = ~n31044 & ~n36432;
  assign n31593 = ~n31576 & ~n31592;
  assign n31594 = ~n36360 & ~n31588;
  assign n31595 = ~n31587 & n31594;
  assign n31596 = n11229 & ~n31595;
  assign n31597 = n36360 & ~n36432;
  assign n31598 = ~n31596 & ~n31597;
  assign n31599 = ~n31044 & ~n31579;
  assign n31600 = ~n10681 & n36433;
  assign n31601 = ~n30213 & ~n30215;
  assign n31602 = ~n30836 & n31601;
  assign n31603 = ~n36251 & ~n31602;
  assign n31604 = ~n30215 & n36251;
  assign n31605 = ~n30213 & n31604;
  assign n31606 = n36251 & n31602;
  assign n31607 = ~n30836 & n31605;
  assign n31608 = ~n31603 & ~n36434;
  assign n31609 = ~n31600 & n31608;
  assign n31610 = n10086 & n31030;
  assign n31611 = n10681 & ~n36433;
  assign n31612 = ~n31610 & ~n31611;
  assign n31613 = ~n31609 & n31612;
  assign n31614 = n10681 & n31608;
  assign n31615 = ~n10681 & ~n31608;
  assign n31616 = ~n36433 & ~n31615;
  assign n31617 = ~n31597 & ~n31608;
  assign n31618 = ~n31596 & ~n31608;
  assign n31619 = ~n31597 & n31618;
  assign n31620 = ~n31596 & n31617;
  assign n31621 = n10681 & ~n36435;
  assign n31622 = ~n36433 & n31608;
  assign n31623 = ~n31621 & ~n31622;
  assign n31624 = ~n31609 & ~n31611;
  assign n31625 = ~n31614 & ~n31616;
  assign n31626 = ~n31031 & ~n36436;
  assign n31627 = ~n31610 & ~n31626;
  assign n31628 = ~n31030 & ~n31622;
  assign n31629 = ~n31621 & n31628;
  assign n31630 = n10086 & ~n31629;
  assign n31631 = n31030 & ~n36436;
  assign n31632 = ~n31630 & ~n31631;
  assign n31633 = ~n31031 & ~n31613;
  assign n31634 = ~n9565 & n36437;
  assign n31635 = ~n30248 & ~n30250;
  assign n31636 = ~n30836 & n31635;
  assign n31637 = ~n36256 & ~n31636;
  assign n31638 = ~n30250 & n36256;
  assign n31639 = ~n30248 & n31638;
  assign n31640 = n36256 & n31636;
  assign n31641 = ~n30836 & n31639;
  assign n31642 = ~n31637 & ~n36438;
  assign n31643 = ~n31634 & n31642;
  assign n31644 = n8998 & n36357;
  assign n31645 = n9565 & ~n36437;
  assign n31646 = ~n31644 & ~n31645;
  assign n31647 = ~n31643 & n31646;
  assign n31648 = n9565 & n31642;
  assign n31649 = ~n9565 & ~n31642;
  assign n31650 = ~n36437 & ~n31649;
  assign n31651 = ~n31631 & ~n31642;
  assign n31652 = ~n31630 & ~n31642;
  assign n31653 = ~n31631 & n31652;
  assign n31654 = ~n31630 & n31651;
  assign n31655 = n9565 & ~n36439;
  assign n31656 = ~n36437 & n31642;
  assign n31657 = ~n31655 & ~n31656;
  assign n31658 = ~n31643 & ~n31645;
  assign n31659 = ~n31648 & ~n31650;
  assign n31660 = ~n31022 & ~n36440;
  assign n31661 = ~n31644 & ~n31660;
  assign n31662 = ~n36357 & ~n31656;
  assign n31663 = ~n31655 & n31662;
  assign n31664 = n8998 & ~n31663;
  assign n31665 = n36357 & ~n36440;
  assign n31666 = ~n31664 & ~n31665;
  assign n31667 = ~n31022 & ~n31647;
  assign n31668 = ~n8506 & n36441;
  assign n31669 = ~n30279 & ~n30281;
  assign n31670 = ~n30836 & n31669;
  assign n31671 = ~n36260 & ~n31670;
  assign n31672 = ~n30281 & n36260;
  assign n31673 = ~n30279 & n31672;
  assign n31674 = n36260 & n31670;
  assign n31675 = ~n30836 & n31673;
  assign n31676 = ~n31671 & ~n36442;
  assign n31677 = ~n31668 & n31676;
  assign n31678 = n7975 & n31008;
  assign n31679 = n8506 & ~n36441;
  assign n31680 = ~n31678 & ~n31679;
  assign n31681 = ~n31677 & n31680;
  assign n31682 = n8506 & n31676;
  assign n31683 = ~n8506 & ~n31676;
  assign n31684 = ~n36441 & ~n31683;
  assign n31685 = ~n31665 & ~n31676;
  assign n31686 = ~n31664 & ~n31676;
  assign n31687 = ~n31665 & n31686;
  assign n31688 = ~n31664 & n31685;
  assign n31689 = n8506 & ~n36443;
  assign n31690 = ~n36441 & n31676;
  assign n31691 = ~n31689 & ~n31690;
  assign n31692 = ~n31677 & ~n31679;
  assign n31693 = ~n31682 & ~n31684;
  assign n31694 = ~n31009 & ~n36444;
  assign n31695 = ~n31678 & ~n31694;
  assign n31696 = ~n31008 & ~n31690;
  assign n31697 = ~n31689 & n31696;
  assign n31698 = n7975 & ~n31697;
  assign n31699 = n31008 & ~n36444;
  assign n31700 = ~n31698 & ~n31699;
  assign n31701 = ~n31009 & ~n31681;
  assign n31702 = ~n7512 & n36445;
  assign n31703 = ~n30314 & ~n30316;
  assign n31704 = ~n30836 & n31703;
  assign n31705 = ~n36265 & ~n31704;
  assign n31706 = ~n30316 & n36265;
  assign n31707 = ~n30314 & n31706;
  assign n31708 = n36265 & n31704;
  assign n31709 = ~n30836 & n31707;
  assign n31710 = ~n31705 & ~n36446;
  assign n31711 = ~n31702 & n31710;
  assign n31712 = n7015 & n36354;
  assign n31713 = n7512 & ~n36445;
  assign n31714 = ~n31712 & ~n31713;
  assign n31715 = ~n31711 & n31714;
  assign n31716 = n7512 & n31710;
  assign n31717 = ~n7512 & ~n31710;
  assign n31718 = ~n36445 & ~n31717;
  assign n31719 = ~n31699 & ~n31710;
  assign n31720 = ~n31698 & ~n31710;
  assign n31721 = ~n31699 & n31720;
  assign n31722 = ~n31698 & n31719;
  assign n31723 = n7512 & ~n36447;
  assign n31724 = ~n36445 & n31710;
  assign n31725 = ~n31723 & ~n31724;
  assign n31726 = ~n31711 & ~n31713;
  assign n31727 = ~n31716 & ~n31718;
  assign n31728 = ~n31000 & ~n36448;
  assign n31729 = ~n31712 & ~n31728;
  assign n31730 = ~n36354 & ~n31724;
  assign n31731 = ~n31723 & n31730;
  assign n31732 = n7015 & ~n31731;
  assign n31733 = n36354 & ~n36448;
  assign n31734 = ~n31732 & ~n31733;
  assign n31735 = ~n31000 & ~n31715;
  assign n31736 = ~n6579 & n36449;
  assign n31737 = ~n30345 & ~n30347;
  assign n31738 = ~n30836 & n31737;
  assign n31739 = ~n36269 & ~n31738;
  assign n31740 = ~n30347 & n36269;
  assign n31741 = ~n30345 & n31740;
  assign n31742 = n36269 & n31738;
  assign n31743 = ~n30836 & n31741;
  assign n31744 = ~n31739 & ~n36450;
  assign n31745 = ~n31736 & n31744;
  assign n31746 = n6117 & n30986;
  assign n31747 = n6579 & ~n36449;
  assign n31748 = ~n31746 & ~n31747;
  assign n31749 = ~n31745 & n31748;
  assign n31750 = n6579 & n31744;
  assign n31751 = ~n6579 & ~n31744;
  assign n31752 = ~n36449 & ~n31751;
  assign n31753 = ~n31733 & ~n31744;
  assign n31754 = ~n31732 & ~n31744;
  assign n31755 = ~n31733 & n31754;
  assign n31756 = ~n31732 & n31753;
  assign n31757 = n6579 & ~n36451;
  assign n31758 = ~n36449 & n31744;
  assign n31759 = ~n31757 & ~n31758;
  assign n31760 = ~n31745 & ~n31747;
  assign n31761 = ~n31750 & ~n31752;
  assign n31762 = ~n30987 & ~n36452;
  assign n31763 = ~n31746 & ~n31762;
  assign n31764 = ~n30986 & ~n31758;
  assign n31765 = ~n31757 & n31764;
  assign n31766 = n6117 & ~n31765;
  assign n31767 = n30986 & ~n36452;
  assign n31768 = ~n31766 & ~n31767;
  assign n31769 = ~n30987 & ~n31749;
  assign n31770 = ~n5708 & n36453;
  assign n31771 = ~n30380 & ~n30382;
  assign n31772 = ~n30836 & n31771;
  assign n31773 = ~n36274 & ~n31772;
  assign n31774 = ~n30382 & n36274;
  assign n31775 = ~n30380 & n31774;
  assign n31776 = n36274 & n31772;
  assign n31777 = ~n30836 & n31775;
  assign n31778 = ~n31773 & ~n36454;
  assign n31779 = ~n31770 & n31778;
  assign n31780 = n5278 & n36351;
  assign n31781 = n5708 & ~n36453;
  assign n31782 = ~n31780 & ~n31781;
  assign n31783 = ~n31779 & n31782;
  assign n31784 = n5708 & n31778;
  assign n31785 = ~n5708 & ~n31778;
  assign n31786 = ~n36453 & ~n31785;
  assign n31787 = ~n31767 & ~n31778;
  assign n31788 = ~n31766 & ~n31778;
  assign n31789 = ~n31767 & n31788;
  assign n31790 = ~n31766 & n31787;
  assign n31791 = n5708 & ~n36455;
  assign n31792 = ~n36453 & n31778;
  assign n31793 = ~n31791 & ~n31792;
  assign n31794 = ~n31779 & ~n31781;
  assign n31795 = ~n31784 & ~n31786;
  assign n31796 = ~n30978 & ~n36456;
  assign n31797 = ~n31780 & ~n31796;
  assign n31798 = ~n36351 & ~n31792;
  assign n31799 = ~n31791 & n31798;
  assign n31800 = n5278 & ~n31799;
  assign n31801 = n36351 & ~n36456;
  assign n31802 = ~n31800 & ~n31801;
  assign n31803 = ~n30978 & ~n31783;
  assign n31804 = ~n4903 & n36457;
  assign n31805 = ~n30411 & ~n30413;
  assign n31806 = ~n30836 & n31805;
  assign n31807 = ~n36278 & ~n31806;
  assign n31808 = ~n30413 & n36278;
  assign n31809 = ~n30411 & n31808;
  assign n31810 = n36278 & n31806;
  assign n31811 = ~n30836 & n31809;
  assign n31812 = ~n31807 & ~n36458;
  assign n31813 = ~n31804 & n31812;
  assign n31814 = n4508 & n30964;
  assign n31815 = n4903 & ~n36457;
  assign n31816 = ~n31814 & ~n31815;
  assign n31817 = ~n31813 & n31816;
  assign n31818 = n4903 & n31812;
  assign n31819 = ~n4903 & ~n31812;
  assign n31820 = ~n36457 & ~n31819;
  assign n31821 = ~n31801 & ~n31812;
  assign n31822 = ~n31800 & ~n31812;
  assign n31823 = ~n31801 & n31822;
  assign n31824 = ~n31800 & n31821;
  assign n31825 = n4903 & ~n36459;
  assign n31826 = ~n36457 & n31812;
  assign n31827 = ~n31825 & ~n31826;
  assign n31828 = ~n31813 & ~n31815;
  assign n31829 = ~n31818 & ~n31820;
  assign n31830 = ~n30965 & ~n36460;
  assign n31831 = ~n31814 & ~n31830;
  assign n31832 = ~n30964 & ~n31826;
  assign n31833 = ~n31825 & n31832;
  assign n31834 = n4508 & ~n31833;
  assign n31835 = n30964 & ~n36460;
  assign n31836 = ~n31834 & ~n31835;
  assign n31837 = ~n30965 & ~n31817;
  assign n31838 = ~n4155 & n36461;
  assign n31839 = ~n30446 & ~n30448;
  assign n31840 = ~n30836 & n31839;
  assign n31841 = ~n36283 & ~n31840;
  assign n31842 = ~n30448 & n36283;
  assign n31843 = ~n30446 & n31842;
  assign n31844 = n36283 & n31840;
  assign n31845 = ~n30836 & n31843;
  assign n31846 = ~n31841 & ~n36462;
  assign n31847 = ~n31838 & n31846;
  assign n31848 = n3788 & n36348;
  assign n31849 = n4155 & ~n36461;
  assign n31850 = ~n31848 & ~n31849;
  assign n31851 = ~n31847 & n31850;
  assign n31852 = n4155 & n31846;
  assign n31853 = ~n4155 & ~n31846;
  assign n31854 = ~n36461 & ~n31853;
  assign n31855 = ~n31835 & ~n31846;
  assign n31856 = ~n31834 & ~n31846;
  assign n31857 = ~n31835 & n31856;
  assign n31858 = ~n31834 & n31855;
  assign n31859 = n4155 & ~n36463;
  assign n31860 = ~n36461 & n31846;
  assign n31861 = ~n31859 & ~n31860;
  assign n31862 = ~n31847 & ~n31849;
  assign n31863 = ~n31852 & ~n31854;
  assign n31864 = ~n30956 & ~n36464;
  assign n31865 = ~n31848 & ~n31864;
  assign n31866 = ~n36348 & ~n31860;
  assign n31867 = ~n31859 & n31866;
  assign n31868 = n3788 & ~n31867;
  assign n31869 = n36348 & ~n36464;
  assign n31870 = ~n31868 & ~n31869;
  assign n31871 = ~n30956 & ~n31851;
  assign n31872 = ~n3473 & n36465;
  assign n31873 = ~n30477 & ~n30479;
  assign n31874 = ~n30836 & n31873;
  assign n31875 = ~n36287 & ~n31874;
  assign n31876 = ~n30479 & n36287;
  assign n31877 = ~n30477 & n31876;
  assign n31878 = n36287 & n31874;
  assign n31879 = ~n30836 & n31877;
  assign n31880 = ~n31875 & ~n36466;
  assign n31881 = ~n31872 & n31880;
  assign n31882 = n3140 & n30942;
  assign n31883 = n3473 & ~n36465;
  assign n31884 = ~n31882 & ~n31883;
  assign n31885 = ~n31881 & n31884;
  assign n31886 = n3473 & n31880;
  assign n31887 = ~n3473 & ~n31880;
  assign n31888 = ~n36465 & ~n31887;
  assign n31889 = ~n31869 & ~n31880;
  assign n31890 = ~n31868 & ~n31880;
  assign n31891 = ~n31869 & n31890;
  assign n31892 = ~n31868 & n31889;
  assign n31893 = n3473 & ~n36467;
  assign n31894 = ~n36465 & n31880;
  assign n31895 = ~n31893 & ~n31894;
  assign n31896 = ~n31881 & ~n31883;
  assign n31897 = ~n31886 & ~n31888;
  assign n31898 = ~n30943 & ~n36468;
  assign n31899 = ~n31882 & ~n31898;
  assign n31900 = ~n30942 & ~n31894;
  assign n31901 = ~n31893 & n31900;
  assign n31902 = n3140 & ~n31901;
  assign n31903 = n30942 & ~n36468;
  assign n31904 = ~n31902 & ~n31903;
  assign n31905 = ~n30943 & ~n31885;
  assign n31906 = ~n2855 & n36469;
  assign n31907 = ~n30512 & ~n30514;
  assign n31908 = ~n30836 & n31907;
  assign n31909 = ~n36292 & ~n31908;
  assign n31910 = ~n30514 & n36292;
  assign n31911 = ~n30512 & n31910;
  assign n31912 = n36292 & n31908;
  assign n31913 = ~n30836 & n31911;
  assign n31914 = ~n31909 & ~n36470;
  assign n31915 = ~n31906 & n31914;
  assign n31916 = n2556 & n36345;
  assign n31917 = n2855 & ~n36469;
  assign n31918 = ~n31916 & ~n31917;
  assign n31919 = ~n31915 & n31918;
  assign n31920 = n2855 & n31914;
  assign n31921 = ~n2855 & ~n31914;
  assign n31922 = ~n36469 & ~n31921;
  assign n31923 = ~n31903 & ~n31914;
  assign n31924 = ~n31902 & ~n31914;
  assign n31925 = ~n31903 & n31924;
  assign n31926 = ~n31902 & n31923;
  assign n31927 = n2855 & ~n36471;
  assign n31928 = ~n36469 & n31914;
  assign n31929 = ~n31927 & ~n31928;
  assign n31930 = ~n31915 & ~n31917;
  assign n31931 = ~n31920 & ~n31922;
  assign n31932 = ~n30934 & ~n36472;
  assign n31933 = ~n31916 & ~n31932;
  assign n31934 = ~n36345 & ~n31928;
  assign n31935 = ~n31927 & n31934;
  assign n31936 = n2556 & ~n31935;
  assign n31937 = n36345 & ~n36472;
  assign n31938 = ~n31936 & ~n31937;
  assign n31939 = ~n30934 & ~n31919;
  assign n31940 = ~n2301 & n36473;
  assign n31941 = ~n30543 & ~n30545;
  assign n31942 = ~n30836 & n31941;
  assign n31943 = ~n36296 & ~n31942;
  assign n31944 = ~n30545 & n36296;
  assign n31945 = ~n30543 & n31944;
  assign n31946 = n36296 & n31942;
  assign n31947 = ~n30836 & n31945;
  assign n31948 = ~n31943 & ~n36474;
  assign n31949 = ~n31940 & n31948;
  assign n31950 = n2038 & n30920;
  assign n31951 = n2301 & ~n36473;
  assign n31952 = ~n31950 & ~n31951;
  assign n31953 = ~n31949 & n31952;
  assign n31954 = n2301 & n31948;
  assign n31955 = ~n2301 & ~n31948;
  assign n31956 = ~n36473 & ~n31955;
  assign n31957 = ~n31937 & ~n31948;
  assign n31958 = ~n31936 & ~n31948;
  assign n31959 = ~n31937 & n31958;
  assign n31960 = ~n31936 & n31957;
  assign n31961 = n2301 & ~n36475;
  assign n31962 = ~n36473 & n31948;
  assign n31963 = ~n31961 & ~n31962;
  assign n31964 = ~n31949 & ~n31951;
  assign n31965 = ~n31954 & ~n31956;
  assign n31966 = ~n30921 & ~n36476;
  assign n31967 = ~n31950 & ~n31966;
  assign n31968 = ~n30920 & ~n31962;
  assign n31969 = ~n31961 & n31968;
  assign n31970 = n2038 & ~n31969;
  assign n31971 = n30920 & ~n36476;
  assign n31972 = ~n31970 & ~n31971;
  assign n31973 = ~n30921 & ~n31953;
  assign n31974 = ~n1812 & n36477;
  assign n31975 = ~n30578 & ~n30580;
  assign n31976 = ~n30836 & n31975;
  assign n31977 = ~n36301 & ~n31976;
  assign n31978 = ~n30580 & n36301;
  assign n31979 = ~n30578 & n31978;
  assign n31980 = n36301 & n31976;
  assign n31981 = ~n30836 & n31979;
  assign n31982 = ~n31977 & ~n36478;
  assign n31983 = ~n31974 & n31982;
  assign n31984 = n1582 & n36342;
  assign n31985 = n1812 & ~n36477;
  assign n31986 = ~n31984 & ~n31985;
  assign n31987 = ~n31983 & n31986;
  assign n31988 = n1812 & n31982;
  assign n31989 = ~n1812 & ~n31982;
  assign n31990 = ~n36477 & ~n31989;
  assign n31991 = ~n31971 & ~n31982;
  assign n31992 = ~n31970 & ~n31982;
  assign n31993 = ~n31971 & n31992;
  assign n31994 = ~n31970 & n31991;
  assign n31995 = n1812 & ~n36479;
  assign n31996 = ~n36477 & n31982;
  assign n31997 = ~n31995 & ~n31996;
  assign n31998 = ~n31983 & ~n31985;
  assign n31999 = ~n31988 & ~n31990;
  assign n32000 = ~n30912 & ~n36480;
  assign n32001 = ~n31984 & ~n32000;
  assign n32002 = ~n36342 & ~n31996;
  assign n32003 = ~n31995 & n32002;
  assign n32004 = n1582 & ~n32003;
  assign n32005 = n36342 & ~n36480;
  assign n32006 = ~n32004 & ~n32005;
  assign n32007 = ~n30912 & ~n31987;
  assign n32008 = ~n1388 & n36481;
  assign n32009 = ~n30609 & ~n30611;
  assign n32010 = ~n30836 & n32009;
  assign n32011 = ~n36305 & ~n32010;
  assign n32012 = ~n30611 & n36305;
  assign n32013 = ~n30609 & n32012;
  assign n32014 = n36305 & n32010;
  assign n32015 = ~n30836 & n32013;
  assign n32016 = ~n32011 & ~n36482;
  assign n32017 = ~n32008 & n32016;
  assign n32018 = n1192 & n30898;
  assign n32019 = n1388 & ~n36481;
  assign n32020 = ~n32018 & ~n32019;
  assign n32021 = ~n32017 & n32020;
  assign n32022 = n1388 & n32016;
  assign n32023 = ~n1388 & ~n32016;
  assign n32024 = ~n36481 & ~n32023;
  assign n32025 = ~n32005 & ~n32016;
  assign n32026 = ~n32004 & ~n32016;
  assign n32027 = ~n32005 & n32026;
  assign n32028 = ~n32004 & n32025;
  assign n32029 = n1388 & ~n36483;
  assign n32030 = ~n36481 & n32016;
  assign n32031 = ~n32029 & ~n32030;
  assign n32032 = ~n32017 & ~n32019;
  assign n32033 = ~n32022 & ~n32024;
  assign n32034 = ~n30899 & ~n36484;
  assign n32035 = ~n32018 & ~n32034;
  assign n32036 = ~n30898 & ~n32030;
  assign n32037 = ~n32029 & n32036;
  assign n32038 = n1192 & ~n32037;
  assign n32039 = n30898 & ~n36484;
  assign n32040 = ~n32038 & ~n32039;
  assign n32041 = ~n30899 & ~n32021;
  assign n32042 = ~n1028 & n36485;
  assign n32043 = ~n30644 & ~n30646;
  assign n32044 = ~n30836 & n32043;
  assign n32045 = ~n36310 & ~n32044;
  assign n32046 = ~n30646 & n36310;
  assign n32047 = ~n30644 & n32046;
  assign n32048 = n36310 & n32044;
  assign n32049 = ~n30836 & n32047;
  assign n32050 = ~n32045 & ~n36486;
  assign n32051 = ~n32042 & n32050;
  assign n32052 = n866 & n36339;
  assign n32053 = n1028 & ~n36485;
  assign n32054 = ~n32052 & ~n32053;
  assign n32055 = ~n32051 & n32054;
  assign n32056 = n1028 & n32050;
  assign n32057 = ~n1028 & ~n32050;
  assign n32058 = ~n36485 & ~n32057;
  assign n32059 = ~n32039 & ~n32050;
  assign n32060 = ~n32038 & ~n32050;
  assign n32061 = ~n32039 & n32060;
  assign n32062 = ~n32038 & n32059;
  assign n32063 = n1028 & ~n36487;
  assign n32064 = ~n36485 & n32050;
  assign n32065 = ~n32063 & ~n32064;
  assign n32066 = ~n32051 & ~n32053;
  assign n32067 = ~n32056 & ~n32058;
  assign n32068 = ~n30890 & ~n36488;
  assign n32069 = ~n32052 & ~n32068;
  assign n32070 = ~n36339 & ~n32064;
  assign n32071 = ~n32063 & n32070;
  assign n32072 = n866 & ~n32071;
  assign n32073 = n36339 & ~n36488;
  assign n32074 = ~n32072 & ~n32073;
  assign n32075 = ~n30890 & ~n32055;
  assign n32076 = ~n730 & n36489;
  assign n32077 = ~n30675 & ~n30677;
  assign n32078 = ~n30836 & n32077;
  assign n32079 = ~n36314 & ~n32078;
  assign n32080 = ~n30677 & n36314;
  assign n32081 = ~n30675 & n32080;
  assign n32082 = n36314 & n32078;
  assign n32083 = ~n30836 & n32081;
  assign n32084 = ~n32079 & ~n36490;
  assign n32085 = ~n32076 & n32084;
  assign n32086 = n602 & n30876;
  assign n32087 = n730 & ~n36489;
  assign n32088 = ~n32086 & ~n32087;
  assign n32089 = ~n32085 & n32088;
  assign n32090 = n730 & n32084;
  assign n32091 = ~n730 & ~n32084;
  assign n32092 = ~n36489 & ~n32091;
  assign n32093 = ~n32073 & ~n32084;
  assign n32094 = ~n32072 & ~n32084;
  assign n32095 = ~n32073 & n32094;
  assign n32096 = ~n32072 & n32093;
  assign n32097 = n730 & ~n36491;
  assign n32098 = ~n36489 & n32084;
  assign n32099 = ~n32097 & ~n32098;
  assign n32100 = ~n32085 & ~n32087;
  assign n32101 = ~n32090 & ~n32092;
  assign n32102 = ~n30877 & ~n36492;
  assign n32103 = ~n32086 & ~n32102;
  assign n32104 = ~n30876 & ~n32098;
  assign n32105 = ~n32097 & n32104;
  assign n32106 = n602 & ~n32105;
  assign n32107 = n30876 & ~n36492;
  assign n32108 = ~n32106 & ~n32107;
  assign n32109 = ~n30877 & ~n32089;
  assign n32110 = ~n497 & n36493;
  assign n32111 = ~n30710 & ~n30712;
  assign n32112 = ~n30836 & n32111;
  assign n32113 = ~n36319 & ~n32112;
  assign n32114 = ~n30712 & n36319;
  assign n32115 = ~n30710 & n32114;
  assign n32116 = n36319 & n32112;
  assign n32117 = ~n30836 & n32115;
  assign n32118 = ~n32113 & ~n36494;
  assign n32119 = ~n32110 & n32118;
  assign n32120 = ~n30727 & ~n36321;
  assign n32121 = ~n30727 & ~n30836;
  assign n32122 = ~n36321 & n32121;
  assign n32123 = ~n30836 & n32120;
  assign n32124 = n30735 & ~n36495;
  assign n32125 = n30739 & n32121;
  assign n32126 = ~n30735 & ~n36495;
  assign n32127 = ~n30727 & n30735;
  assign n32128 = ~n36321 & n32127;
  assign n32129 = ~n30836 & n32128;
  assign n32130 = ~n32126 & ~n32129;
  assign n32131 = ~n32124 & ~n32125;
  assign n32132 = n403 & n36496;
  assign n32133 = n497 & ~n36493;
  assign n32134 = ~n32132 & ~n32133;
  assign n32135 = ~n32119 & n32134;
  assign n32136 = ~n403 & ~n36496;
  assign n32137 = ~n30741 & ~n30743;
  assign n32138 = ~n30836 & n32137;
  assign n32139 = ~n36323 & ~n32138;
  assign n32140 = ~n30743 & n36323;
  assign n32141 = ~n30741 & n32140;
  assign n32142 = n36323 & n32138;
  assign n32143 = ~n30836 & n32141;
  assign n32144 = ~n32139 & ~n36497;
  assign n32145 = ~n330 & ~n32144;
  assign n32146 = ~n32136 & ~n32145;
  assign n32147 = n497 & n32118;
  assign n32148 = ~n497 & ~n32118;
  assign n32149 = ~n36493 & ~n32148;
  assign n32150 = ~n32107 & ~n32118;
  assign n32151 = ~n32106 & ~n32118;
  assign n32152 = ~n32107 & n32151;
  assign n32153 = ~n32106 & n32150;
  assign n32154 = n497 & ~n36498;
  assign n32155 = ~n36493 & n32118;
  assign n32156 = ~n32154 & ~n32155;
  assign n32157 = ~n32119 & ~n32133;
  assign n32158 = ~n32147 & ~n32149;
  assign n32159 = ~n32136 & ~n36499;
  assign n32160 = ~n36496 & ~n32155;
  assign n32161 = ~n32154 & n32160;
  assign n32162 = n403 & ~n32161;
  assign n32163 = n36496 & ~n36499;
  assign n32164 = ~n32162 & ~n32163;
  assign n32165 = ~n32132 & ~n32159;
  assign n32166 = ~n32145 & ~n36500;
  assign n32167 = ~n32135 & n32146;
  assign n32168 = n330 & n32144;
  assign n32169 = ~n30758 & ~n36324;
  assign n32170 = ~n30836 & n32169;
  assign n32171 = ~n36326 & ~n32170;
  assign n32172 = ~n30758 & n36326;
  assign n32173 = ~n36324 & n32172;
  assign n32174 = n36326 & n32170;
  assign n32175 = ~n30836 & n32173;
  assign n32176 = ~n32171 & ~n36502;
  assign n32177 = n271 & n32176;
  assign n32178 = ~n32168 & ~n32177;
  assign n32179 = ~n36501 & n32178;
  assign n32180 = ~n271 & ~n32176;
  assign n32181 = ~n217 & ~n36336;
  assign n32182 = ~n32180 & ~n32181;
  assign n32183 = ~n32179 & n32182;
  assign n32184 = ~n330 & n36500;
  assign n32185 = n32144 & ~n32184;
  assign n32186 = n330 & ~n36500;
  assign n32187 = ~n32144 & ~n32163;
  assign n32188 = ~n32144 & ~n32162;
  assign n32189 = ~n32163 & n32188;
  assign n32190 = ~n32162 & n32187;
  assign n32191 = n330 & ~n36503;
  assign n32192 = n32144 & ~n36500;
  assign n32193 = ~n32191 & ~n32192;
  assign n32194 = ~n32185 & ~n32186;
  assign n32195 = ~n32180 & ~n36504;
  assign n32196 = ~n32176 & ~n32192;
  assign n32197 = ~n32191 & n32196;
  assign n32198 = n271 & ~n32197;
  assign n32199 = n32176 & ~n36504;
  assign n32200 = ~n32198 & ~n32199;
  assign n32201 = ~n32177 & ~n32195;
  assign n32202 = ~n36336 & ~n32199;
  assign n32203 = ~n32198 & n32202;
  assign n32204 = ~n36336 & ~n32198;
  assign n32205 = ~n32199 & n32204;
  assign n32206 = ~n36336 & n36505;
  assign n32207 = n217 & ~n36506;
  assign n32208 = n36336 & ~n36505;
  assign n32209 = ~n32207 & ~n32208;
  assign n32210 = ~n30868 & ~n32183;
  assign n32211 = ~n30857 & ~n36507;
  assign n32212 = ~n36335 & ~n32208;
  assign n32213 = ~n32207 & n32212;
  assign n32214 = n198 & ~n32213;
  assign n32215 = n36335 & ~n36507;
  assign n32216 = ~n32214 & ~n32215;
  assign n32217 = ~n30856 & ~n32211;
  assign n32218 = ~n30845 & ~n36508;
  assign n32219 = ~n30820 & ~n30836;
  assign n32220 = n30812 & ~n32219;
  assign n32221 = ~n30812 & ~n30820;
  assign n32222 = ~n193 & ~n32221;
  assign n32223 = ~n32220 & n32222;
  assign n32224 = ~n30812 & n32219;
  assign n32225 = ~n30836 & n32221;
  assign n32226 = ~n36333 & ~n36509;
  assign n32227 = ~n30844 & n32226;
  assign n32228 = n193 & ~n32227;
  assign n32229 = ~n32223 & ~n32228;
  assign n32230 = ~n32215 & n32227;
  assign n32231 = ~n32214 & n32230;
  assign n32232 = ~n32214 & n32227;
  assign n32233 = ~n32215 & n32232;
  assign n32234 = n36508 & n32227;
  assign n32235 = n193 & ~n36510;
  assign n32236 = n30844 & ~n36508;
  assign n32237 = ~n32223 & ~n32236;
  assign n32238 = ~n32235 & n32237;
  assign n32239 = ~n32218 & n32229;
  assign n32240 = n201 | n202;
  assign n32241 = n214 | n215;
  assign n32242 = n225 | ~n226;
  assign n32243 = n227 | n228;
  assign n32244 = n231 | n232;
  assign n32245 = n237 | ~n238;
  assign n32246 = n241 | n242;
  assign n32247 = n246 | n247;
  assign n32248 = n251 | n252;
  assign n32249 = n253 | ~n254;
  assign n32250 = n257 | n258;
  assign n32251 = n269 | n265 | n268;
  assign n32252 = n279 | n280;
  assign n32253 = n285 | n286;
  assign n32254 = ~n294 | n292 | n293;
  assign n32255 = n300 | n301;
  assign n32256 = n309 | n310;
  assign n32257 = n318 | n319;
  assign n32258 = n327 | n328;
  assign n32259 = n338 | n339;
  assign n32260 = n344 | n345;
  assign n32261 = n348 | n349;
  assign n32262 = n359 | n360;
  assign n32263 = n363 | n364;
  assign n32264 = n374 | n375;
  assign n32265 = n376 | n377;
  assign n32266 = n386 | n387;
  assign n32267 = n396 | n397;
  assign n32268 = n411 | n412;
  assign n32269 = n423 | n424;
  assign n32270 = n436 | n437;
  assign n32271 = n443 | n444;
  assign n32272 = n449 | n450;
  assign n32273 = n459 | n460;
  assign n32274 = n467 | ~n468;
  assign n32275 = n477 | n478;
  assign n32276 = n480 | ~n481;
  assign n32277 = n484 | n485;
  assign n32278 = n491 | n492;
  assign n32279 = n507 | n508;
  assign n32280 = n513 | n514;
  assign n32281 = n517 | n518;
  assign n32282 = n529 | n530;
  assign n32283 = n533 | n534;
  assign n32284 = n544 | n545;
  assign n32285 = n555 | n556;
  assign n32286 = n559 | n560;
  assign n32287 = n572 | n573;
  assign n32288 = n575 | ~n576;
  assign n32289 = n584 | n585;
  assign n32290 = n589 | n590;
  assign n32291 = n596 | n597;
  assign n32292 = n610 | n611;
  assign n32293 = n617 | n618;
  assign n32294 = n623 | n624;
  assign n32295 = n636 | n637;
  assign n32296 = n643 | n644;
  assign n32297 = n649 | n650;
  assign n32298 = n659 | n660;
  assign n32299 = n667 | ~n668;
  assign n32300 = n673 | n674;
  assign n32301 = n681 | n682;
  assign n32302 = n684 | ~n685;
  assign n32303 = n693 | n694;
  assign n32304 = n701 | ~n702;
  assign n32305 = n713 | ~n714;
  assign n32306 = n717 | n718;
  assign n32307 = n724 | n725;
  assign n32308 = n740 | n741;
  assign n32309 = n746 | n747;
  assign n32310 = n750 | n751;
  assign n32311 = n762 | n763;
  assign n32312 = n766 | n767;
  assign n32313 = n777 | n778;
  assign n32314 = n779 | n780;
  assign n32315 = n790 | n791;
  assign n32316 = n794 | n795;
  assign n32317 = n807 | n808;
  assign n32318 = n810 | ~n811;
  assign n32319 = n820 | n821;
  assign n32320 = n824 | n825;
  assign n32321 = n839 | ~n840;
  assign n32322 = n848 | n849;
  assign n32323 = n853 | n854;
  assign n32324 = n860 | n861;
  assign n32325 = n874 | n875;
  assign n32326 = n881 | n882;
  assign n32327 = n887 | n888;
  assign n32328 = n900 | n901;
  assign n32329 = n907 | n908;
  assign n32330 = n913 | n914;
  assign n32331 = n923 | n924;
  assign n32332 = n931 | ~n932;
  assign n32333 = n937 | n938;
  assign n32334 = n945 | n946;
  assign n32335 = n948 | ~n949;
  assign n32336 = n957 | n958;
  assign n32337 = n965 | ~n966;
  assign n32338 = n971 | n972;
  assign n32339 = n981 | ~n982;
  assign n32340 = n990 | n991;
  assign n32341 = n998 | ~n999;
  assign n32342 = n1007 | n1008;
  assign n32343 = n1011 | ~n1012;
  assign n32344 = n1015 | n1016;
  assign n32345 = n1022 | n1023;
  assign n32346 = n1038 | n1039;
  assign n32347 = n1044 | n1045;
  assign n32348 = n1048 | n1049;
  assign n32349 = n1060 | n1061;
  assign n32350 = n1064 | n1065;
  assign n32351 = n1075 | n1076;
  assign n32352 = n1086 | n1087;
  assign n32353 = n1090 | n1091;
  assign n32354 = n1103 | n1104;
  assign n32355 = n1106 | ~n1107;
  assign n32356 = n1116 | n1117;
  assign n32357 = n1120 | n1121;
  assign n32358 = n1135 | ~n1136;
  assign n32359 = n1145 | n1146;
  assign n32360 = n1149 | n1150;
  assign n32361 = n1161 | n1162;
  assign n32362 = n1165 | ~n1166;
  assign n32363 = n1174 | n1175;
  assign n32364 = n1179 | n1180;
  assign n32365 = n1186 | n1187;
  assign n32366 = n1200 | n1201;
  assign n32367 = n1207 | n1208;
  assign n32368 = n1213 | n1214;
  assign n32369 = n1226 | n1227;
  assign n32370 = n1233 | n1234;
  assign n32371 = n1239 | n1240;
  assign n32372 = n1249 | n1250;
  assign n32373 = n1257 | ~n1258;
  assign n32374 = n1263 | n1264;
  assign n32375 = n1271 | n1272;
  assign n32376 = n1274 | ~n1275;
  assign n32377 = n1283 | n1284;
  assign n32378 = n1291 | ~n1292;
  assign n32379 = n1297 | n1298;
  assign n32380 = n1307 | ~n1308;
  assign n32381 = n1316 | n1317;
  assign n32382 = n1324 | ~n1325;
  assign n32383 = n1330 | n1331;
  assign n32384 = n1337 | n1338;
  assign n32385 = n1341 | ~n1342;
  assign n32386 = n1350 | n1351;
  assign n32387 = n1358 | ~n1359;
  assign n32388 = n1367 | n1368;
  assign n32389 = n1371 | ~n1372;
  assign n32390 = n1375 | n1376;
  assign n32391 = n1382 | n1383;
  assign n32392 = n1398 | n1399;
  assign n32393 = n1404 | n1405;
  assign n32394 = n1408 | n1409;
  assign n32395 = n1420 | n1421;
  assign n32396 = n1424 | n1425;
  assign n32397 = n1435 | n1436;
  assign n32398 = n1446 | n1447;
  assign n32399 = n1450 | n1451;
  assign n32400 = n1463 | n1464;
  assign n32401 = n1466 | ~n1467;
  assign n32402 = n1476 | n1477;
  assign n32403 = n1480 | n1481;
  assign n32404 = n1495 | ~n1496;
  assign n32405 = n1505 | n1506;
  assign n32406 = n1509 | n1510;
  assign n32407 = n1521 | n1522;
  assign n32408 = n1525 | ~n1526;
  assign n32409 = n1535 | n1536;
  assign n32410 = n1539 | n1540;
  assign n32411 = n1552 | n1553;
  assign n32412 = n1555 | ~n1556;
  assign n32413 = n1564 | n1565;
  assign n32414 = n1569 | n1570;
  assign n32415 = n1576 | n1577;
  assign n32416 = n1590 | n1591;
  assign n32417 = n1597 | n1598;
  assign n32418 = n1603 | n1604;
  assign n32419 = n1616 | n1617;
  assign n32420 = n1623 | n1624;
  assign n32421 = n1629 | n1630;
  assign n32422 = n1639 | n1640;
  assign n32423 = n1647 | ~n1648;
  assign n32424 = n1653 | n1654;
  assign n32425 = n1661 | n1662;
  assign n32426 = n1664 | ~n1665;
  assign n32427 = n1673 | n1674;
  assign n32428 = n1681 | ~n1682;
  assign n32429 = n1687 | n1688;
  assign n32430 = n1697 | ~n1698;
  assign n32431 = n1706 | n1707;
  assign n32432 = n1714 | ~n1715;
  assign n32433 = n1720 | n1721;
  assign n32434 = n1727 | n1728;
  assign n32435 = n1731 | ~n1732;
  assign n32436 = n1740 | n1741;
  assign n32437 = n1748 | ~n1749;
  assign n32438 = n1754 | n1755;
  assign n32439 = n1761 | n1762;
  assign n32440 = n1765 | ~n1766;
  assign n32441 = n1774 | n1775;
  assign n32442 = n1782 | ~n1783;
  assign n32443 = n1792 | n1793;
  assign n32444 = n1795 | ~n1796;
  assign n32445 = n1799 | n1800;
  assign n32446 = n1806 | n1807;
  assign n32447 = n1822 | n1823;
  assign n32448 = n1828 | n1829;
  assign n32449 = n1832 | n1833;
  assign n32450 = n1844 | n1845;
  assign n32451 = n1848 | n1849;
  assign n32452 = n1859 | n1860;
  assign n32453 = n1870 | n1871;
  assign n32454 = n1874 | n1875;
  assign n32455 = n1887 | n1888;
  assign n32456 = n1890 | ~n1891;
  assign n32457 = n1900 | n1901;
  assign n32458 = n1904 | n1905;
  assign n32459 = n1919 | ~n1920;
  assign n32460 = n1929 | n1930;
  assign n32461 = n1933 | n1934;
  assign n32462 = n1945 | n1946;
  assign n32463 = n1949 | ~n1950;
  assign n32464 = n1959 | n1960;
  assign n32465 = n1963 | n1964;
  assign n32466 = n1975 | n1976;
  assign n32467 = n1979 | ~n1980;
  assign n32468 = n1989 | n1990;
  assign n32469 = n1993 | n1994;
  assign n32470 = n2002 | n2003;
  assign n32471 = n2005 | n2006;
  assign n32472 = n2011 | ~n2012;
  assign n32473 = n2020 | n2021;
  assign n32474 = n2025 | n2026;
  assign n32475 = n2032 | n2033;
  assign n32476 = n2046 | n2047;
  assign n32477 = n2053 | n2054;
  assign n32478 = n2059 | n2060;
  assign n32479 = n2072 | n2073;
  assign n32480 = n2079 | n2080;
  assign n32481 = n2085 | n2086;
  assign n32482 = n2095 | n2096;
  assign n32483 = n2103 | ~n2104;
  assign n32484 = n2109 | n2110;
  assign n32485 = n2117 | n2118;
  assign n32486 = n2120 | ~n2121;
  assign n32487 = n2129 | n2130;
  assign n32488 = n2137 | ~n2138;
  assign n32489 = n2143 | n2144;
  assign n32490 = n2153 | ~n2154;
  assign n32491 = n2162 | n2163;
  assign n32492 = n2170 | ~n2171;
  assign n32493 = n2176 | n2177;
  assign n32494 = n2183 | n2184;
  assign n32495 = n2187 | ~n2188;
  assign n32496 = n2196 | n2197;
  assign n32497 = n2204 | ~n2205;
  assign n32498 = n2210 | n2211;
  assign n32499 = n2217 | n2218;
  assign n32500 = n2221 | ~n2222;
  assign n32501 = n2230 | n2231;
  assign n32502 = n2238 | ~n2239;
  assign n32503 = n2244 | n2245;
  assign n32504 = n2248 | n2249;
  assign n32505 = n2251 | n2252;
  assign n32506 = n2257 | ~n2258;
  assign n32507 = n2266 | n2267;
  assign n32508 = n2274 | ~n2275;
  assign n32509 = n2283 | n2284;
  assign n32510 = n2288 | n2289;
  assign n32511 = n2295 | n2296;
  assign n32512 = n2311 | n2312;
  assign n32513 = n2317 | n2318;
  assign n32514 = n2321 | n2322;
  assign n32515 = n2333 | n2334;
  assign n32516 = n2337 | n2338;
  assign n32517 = n2348 | n2349;
  assign n32518 = n2350 | n2351;
  assign n32519 = n2361 | n2362;
  assign n32520 = n2365 | n2366;
  assign n32521 = n2378 | n2379;
  assign n32522 = n2381 | ~n2382;
  assign n32523 = n2391 | n2392;
  assign n32524 = n2395 | n2396;
  assign n32525 = n2410 | ~n2411;
  assign n32526 = n2420 | n2421;
  assign n32527 = n2424 | n2425;
  assign n32528 = n2436 | n2437;
  assign n32529 = n2440 | ~n2441;
  assign n32530 = n2450 | n2451;
  assign n32531 = n2454 | n2455;
  assign n32532 = n2466 | n2467;
  assign n32533 = n2470 | ~n2471;
  assign n32534 = n2480 | n2481;
  assign n32535 = n2484 | n2485;
  assign n32536 = n2493 | n2494;
  assign n32537 = n2496 | n2497;
  assign n32538 = n2502 | ~n2503;
  assign n32539 = n2512 | n2513;
  assign n32540 = n2516 | n2517;
  assign n32541 = n2528 | n2529;
  assign n32542 = n2538 | n2539;
  assign n32543 = n2543 | n2544;
  assign n32544 = n2550 | n2551;
  assign n32545 = n2564 | n2565;
  assign n32546 = n2571 | n2572;
  assign n32547 = n2577 | n2578;
  assign n32548 = n2590 | n2591;
  assign n32549 = n2597 | n2598;
  assign n32550 = n2603 | n2604;
  assign n32551 = n2613 | n2614;
  assign n32552 = n2621 | ~n2622;
  assign n32553 = n2627 | n2628;
  assign n32554 = n2635 | n2636;
  assign n32555 = n2638 | ~n2639;
  assign n32556 = n2647 | n2648;
  assign n32557 = n2655 | ~n2656;
  assign n32558 = n2661 | n2662;
  assign n32559 = n2671 | ~n2672;
  assign n32560 = n2680 | n2681;
  assign n32561 = n2688 | ~n2689;
  assign n32562 = n2694 | n2695;
  assign n32563 = n2701 | n2702;
  assign n32564 = n2705 | ~n2706;
  assign n32565 = n2714 | n2715;
  assign n32566 = n2722 | ~n2723;
  assign n32567 = n2728 | n2729;
  assign n32568 = n2735 | n2736;
  assign n32569 = n2739 | ~n2740;
  assign n32570 = n2748 | n2749;
  assign n32571 = n2756 | ~n2757;
  assign n32572 = n2762 | n2763;
  assign n32573 = n2766 | n2767;
  assign n32574 = n2769 | n2770;
  assign n32575 = n2775 | ~n2776;
  assign n32576 = n2784 | n2785;
  assign n32577 = n2792 | ~n2793;
  assign n32578 = n2798 | n2799;
  assign n32579 = n2805 | n2806;
  assign n32580 = n2815 | n2816;
  assign n32581 = n2823 | ~n2824;
  assign n32582 = n2829 | n2830;
  assign n32583 = n2832 | n2833;
  assign n32584 = n2838 | ~n2839;
  assign n32585 = n2842 | n2843;
  assign n32586 = n2849 | n2850;
  assign n32587 = n2865 | n2866;
  assign n32588 = n2871 | n2872;
  assign n32589 = n2875 | n2876;
  assign n32590 = n2887 | n2888;
  assign n32591 = n2891 | n2892;
  assign n32592 = n2902 | n2903;
  assign n32593 = n2913 | n2914;
  assign n32594 = n2917 | n2918;
  assign n32595 = n2930 | n2931;
  assign n32596 = n2933 | ~n2934;
  assign n32597 = n2943 | n2944;
  assign n32598 = n2947 | n2948;
  assign n32599 = n2962 | ~n2963;
  assign n32600 = n2972 | n2973;
  assign n32601 = n2976 | n2977;
  assign n32602 = n2988 | n2989;
  assign n32603 = n2992 | ~n2993;
  assign n32604 = n3002 | n3003;
  assign n32605 = n3006 | n3007;
  assign n32606 = n3018 | n3019;
  assign n32607 = n3022 | ~n3023;
  assign n32608 = n3032 | n3033;
  assign n32609 = n3036 | n3037;
  assign n32610 = n3045 | n3046;
  assign n32611 = n3048 | n3049;
  assign n32612 = n3054 | ~n3055;
  assign n32613 = n3064 | n3065;
  assign n32614 = n3068 | n3069;
  assign n32615 = n3080 | n3081;
  assign n32616 = n3091 | n3092;
  assign n32617 = n3095 | n3096;
  assign n32618 = n3104 | n3105;
  assign n32619 = n3107 | n3108;
  assign n32620 = n3113 | ~n3114;
  assign n32621 = n3122 | n3123;
  assign n32622 = n3127 | n3128;
  assign n32623 = n3134 | n3135;
  assign n32624 = n3148 | n3149;
  assign n32625 = n3155 | n3156;
  assign n32626 = n3161 | n3162;
  assign n32627 = n3174 | n3175;
  assign n32628 = n3181 | n3182;
  assign n32629 = n3187 | n3188;
  assign n32630 = n3197 | n3198;
  assign n32631 = n3205 | ~n3206;
  assign n32632 = n3211 | n3212;
  assign n32633 = n3219 | n3220;
  assign n32634 = n3222 | ~n3223;
  assign n32635 = n3231 | n3232;
  assign n32636 = n3239 | ~n3240;
  assign n32637 = n3245 | n3246;
  assign n32638 = n3255 | ~n3256;
  assign n32639 = n3264 | n3265;
  assign n32640 = n3272 | ~n3273;
  assign n32641 = n3278 | n3279;
  assign n32642 = n3285 | n3286;
  assign n32643 = n3289 | ~n3290;
  assign n32644 = n3298 | n3299;
  assign n32645 = n3306 | ~n3307;
  assign n32646 = n3312 | n3313;
  assign n32647 = n3319 | n3320;
  assign n32648 = n3323 | ~n3324;
  assign n32649 = n3332 | n3333;
  assign n32650 = n3340 | ~n3341;
  assign n32651 = n3346 | n3347;
  assign n32652 = n3350 | n3351;
  assign n32653 = n3353 | n3354;
  assign n32654 = n3359 | ~n3360;
  assign n32655 = n3368 | n3369;
  assign n32656 = n3376 | ~n3377;
  assign n32657 = n3382 | n3383;
  assign n32658 = n3389 | n3390;
  assign n32659 = n3399 | n3400;
  assign n32660 = n3407 | ~n3408;
  assign n32661 = n3413 | n3414;
  assign n32662 = n3417 | n3418;
  assign n32663 = n3420 | n3421;
  assign n32664 = n3426 | ~n3427;
  assign n32665 = n3435 | n3436;
  assign n32666 = n3443 | ~n3444;
  assign n32667 = n3453 | n3454;
  assign n32668 = n3456 | ~n3457;
  assign n32669 = n3460 | n3461;
  assign n32670 = n3467 | n3468;
  assign n32671 = n3483 | n3484;
  assign n32672 = n3489 | n3490;
  assign n32673 = n3493 | n3494;
  assign n32674 = n3505 | n3506;
  assign n32675 = n3509 | n3510;
  assign n32676 = n3520 | n3521;
  assign n32677 = n3531 | n3532;
  assign n32678 = n3535 | n3536;
  assign n32679 = n3548 | n3549;
  assign n32680 = n3551 | ~n3552;
  assign n32681 = n3561 | n3562;
  assign n32682 = n3565 | n3566;
  assign n32683 = n3580 | ~n3581;
  assign n32684 = n3590 | n3591;
  assign n32685 = n3594 | n3595;
  assign n32686 = n3606 | n3607;
  assign n32687 = n3610 | ~n3611;
  assign n32688 = n3620 | n3621;
  assign n32689 = n3624 | n3625;
  assign n32690 = n3637 | n3638;
  assign n32691 = n3640 | ~n3641;
  assign n32692 = n3650 | n3651;
  assign n32693 = n3654 | n3655;
  assign n32694 = n3663 | n3664;
  assign n32695 = n3666 | n3667;
  assign n32696 = n3672 | ~n3673;
  assign n32697 = n3682 | n3683;
  assign n32698 = n3686 | n3687;
  assign n32699 = n3698 | n3699;
  assign n32700 = n3709 | n3710;
  assign n32701 = n3713 | n3714;
  assign n32702 = n3722 | n3723;
  assign n32703 = n3725 | n3726;
  assign n32704 = n3731 | ~n3732;
  assign n32705 = n3741 | n3742;
  assign n32706 = n3745 | n3746;
  assign n32707 = n3758 | n3759;
  assign n32708 = n3761 | ~n3762;
  assign n32709 = n3770 | n3771;
  assign n32710 = n3775 | n3776;
  assign n32711 = n3782 | n3783;
  assign n32712 = n3796 | n3797;
  assign n32713 = n3803 | n3804;
  assign n32714 = n3809 | n3810;
  assign n32715 = n3822 | n3823;
  assign n32716 = n3829 | n3830;
  assign n32717 = n3835 | n3836;
  assign n32718 = n3845 | n3846;
  assign n32719 = n3853 | ~n3854;
  assign n32720 = n3859 | n3860;
  assign n32721 = n3867 | n3868;
  assign n32722 = n3870 | ~n3871;
  assign n32723 = n3879 | n3880;
  assign n32724 = n3887 | ~n3888;
  assign n32725 = n3893 | n3894;
  assign n32726 = n3903 | ~n3904;
  assign n32727 = n3912 | n3913;
  assign n32728 = n3920 | ~n3921;
  assign n32729 = n3926 | n3927;
  assign n32730 = n3933 | n3934;
  assign n32731 = n3937 | ~n3938;
  assign n32732 = n3946 | n3947;
  assign n32733 = n3954 | ~n3955;
  assign n32734 = n3960 | n3961;
  assign n32735 = n3967 | n3968;
  assign n32736 = n3971 | ~n3972;
  assign n32737 = n3980 | n3981;
  assign n32738 = n3988 | ~n3989;
  assign n32739 = n3994 | n3995;
  assign n32740 = n4002 | n4003;
  assign n32741 = n4005 | ~n4006;
  assign n32742 = n4014 | n4015;
  assign n32743 = n4022 | ~n4023;
  assign n32744 = n4028 | n4029;
  assign n32745 = n4035 | n4036;
  assign n32746 = n4045 | n4046;
  assign n32747 = n4053 | ~n4054;
  assign n32748 = n4059 | n4060;
  assign n32749 = n4063 | n4064;
  assign n32750 = n4066 | n4067;
  assign n32751 = n4072 | ~n4073;
  assign n32752 = n4081 | n4082;
  assign n32753 = n4089 | ~n4090;
  assign n32754 = n4095 | n4096;
  assign n32755 = n4103 | n4104;
  assign n32756 = n4106 | ~n4107;
  assign n32757 = n4115 | n4116;
  assign n32758 = n4123 | ~n4124;
  assign n32759 = n4129 | n4130;
  assign n32760 = n4132 | n4133;
  assign n32761 = n4138 | ~n4139;
  assign n32762 = n4142 | n4143;
  assign n32763 = n4149 | n4150;
  assign n32764 = n4165 | n4166;
  assign n32765 = n4171 | n4172;
  assign n32766 = n4175 | n4176;
  assign n32767 = n4187 | n4188;
  assign n32768 = n4191 | n4192;
  assign n32769 = n4202 | n4203;
  assign n32770 = n4213 | n4214;
  assign n32771 = n4217 | n4218;
  assign n32772 = n4230 | n4231;
  assign n32773 = n4233 | ~n4234;
  assign n32774 = n4243 | n4244;
  assign n32775 = n4247 | n4248;
  assign n32776 = n4262 | ~n4263;
  assign n32777 = n4272 | n4273;
  assign n32778 = n4276 | n4277;
  assign n32779 = n4288 | n4289;
  assign n32780 = n4292 | ~n4293;
  assign n32781 = n4302 | n4303;
  assign n32782 = n4306 | n4307;
  assign n32783 = n4318 | n4319;
  assign n32784 = n4322 | ~n4323;
  assign n32785 = n4332 | n4333;
  assign n32786 = n4336 | n4337;
  assign n32787 = n4345 | n4346;
  assign n32788 = n4348 | n4349;
  assign n32789 = n4354 | ~n4355;
  assign n32790 = n4364 | n4365;
  assign n32791 = n4368 | n4369;
  assign n32792 = n4377 | n4378;
  assign n32793 = n4379 | n4380;
  assign n32794 = n4384 | n4385;
  assign n32795 = n4387 | ~n4388;
  assign n32796 = n4397 | n4398;
  assign n32797 = n4401 | n4402;
  assign n32798 = n4410 | n4411;
  assign n32799 = n4413 | n4414;
  assign n32800 = n4419 | ~n4420;
  assign n32801 = n4429 | n4430;
  assign n32802 = n4433 | n4434;
  assign n32803 = n4446 | n4447;
  assign n32804 = n4449 | ~n4450;
  assign n32805 = n4459 | n4460;
  assign n32806 = n4463 | n4464;
  assign n32807 = n4472 | n4473;
  assign n32808 = n4475 | n4476;
  assign n32809 = n4481 | ~n4482;
  assign n32810 = n4490 | n4491;
  assign n32811 = n4495 | n4496;
  assign n32812 = n4502 | n4503;
  assign n32813 = n4516 | n4517;
  assign n32814 = n4523 | n4524;
  assign n32815 = n4529 | n4530;
  assign n32816 = n4542 | n4543;
  assign n32817 = n4549 | n4550;
  assign n32818 = n4555 | n4556;
  assign n32819 = n4565 | n4566;
  assign n32820 = n4573 | ~n4574;
  assign n32821 = n4579 | n4580;
  assign n32822 = n4587 | n4588;
  assign n32823 = n4590 | ~n4591;
  assign n32824 = n4599 | n4600;
  assign n32825 = n4607 | ~n4608;
  assign n32826 = n4613 | n4614;
  assign n32827 = n4623 | ~n4624;
  assign n32828 = n4632 | n4633;
  assign n32829 = n4640 | ~n4641;
  assign n32830 = n4646 | n4647;
  assign n32831 = n4653 | n4654;
  assign n32832 = n4657 | ~n4658;
  assign n32833 = n4666 | n4667;
  assign n32834 = n4674 | ~n4675;
  assign n32835 = n4680 | n4681;
  assign n32836 = n4687 | n4688;
  assign n32837 = n4691 | ~n4692;
  assign n32838 = n4700 | n4701;
  assign n32839 = n4708 | ~n4709;
  assign n32840 = n4714 | n4715;
  assign n32841 = n4718 | n4719;
  assign n32842 = n4721 | n4722;
  assign n32843 = n4727 | ~n4728;
  assign n32844 = n4736 | n4737;
  assign n32845 = n4744 | ~n4745;
  assign n32846 = n4750 | n4751;
  assign n32847 = n4757 | n4758;
  assign n32848 = n4767 | n4768;
  assign n32849 = n4775 | ~n4776;
  assign n32850 = n4785 | n4786;
  assign n32851 = n4789 | n4790;
  assign n32852 = n4798 | n4799;
  assign n32853 = n4806 | ~n4807;
  assign n32854 = n4812 | n4813;
  assign n32855 = n4820 | n4821;
  assign n32856 = n4823 | ~n4824;
  assign n32857 = n4832 | n4833;
  assign n32858 = n4840 | ~n4841;
  assign n32859 = n4846 | n4847;
  assign n32860 = n4850 | n4851;
  assign n32861 = n4853 | n4854;
  assign n32862 = n4859 | ~n4860;
  assign n32863 = n4868 | n4869;
  assign n32864 = n4876 | ~n4877;
  assign n32865 = n4885 | n4886;
  assign n32866 = n4890 | n4891;
  assign n32867 = n4897 | n4898;
  assign n32868 = n4913 | n4914;
  assign n32869 = n4919 | n4920;
  assign n32870 = n4923 | n4924;
  assign n32871 = n4935 | n4936;
  assign n32872 = n4939 | n4940;
  assign n32873 = n4950 | n4951;
  assign n32874 = n4961 | n4962;
  assign n32875 = n4965 | n4966;
  assign n32876 = n4978 | n4979;
  assign n32877 = n4981 | ~n4982;
  assign n32878 = n4991 | n4992;
  assign n32879 = n4995 | n4996;
  assign n32880 = n5010 | ~n5011;
  assign n32881 = n5020 | n5021;
  assign n32882 = n5024 | n5025;
  assign n32883 = n5036 | n5037;
  assign n32884 = n5040 | ~n5041;
  assign n32885 = n5050 | n5051;
  assign n32886 = n5054 | n5055;
  assign n32887 = n5066 | n5067;
  assign n32888 = n5070 | ~n5071;
  assign n32889 = n5080 | n5081;
  assign n32890 = n5084 | n5085;
  assign n32891 = n5093 | n5094;
  assign n32892 = n5096 | n5097;
  assign n32893 = n5102 | ~n5103;
  assign n32894 = n5112 | n5113;
  assign n32895 = n5116 | n5117;
  assign n32896 = n5128 | n5129;
  assign n32897 = n5139 | n5140;
  assign n32898 = n5143 | n5144;
  assign n32899 = n5152 | n5153;
  assign n32900 = n5155 | n5156;
  assign n32901 = n5161 | ~n5162;
  assign n32902 = n5171 | n5172;
  assign n32903 = n5175 | n5176;
  assign n32904 = n5184 | n5185;
  assign n32905 = n5192 | ~n5193;
  assign n32906 = n5202 | n5203;
  assign n32907 = n5206 | n5207;
  assign n32908 = n5215 | n5216;
  assign n32909 = n5218 | n5219;
  assign n32910 = n5224 | ~n5225;
  assign n32911 = n5234 | n5235;
  assign n32912 = n5238 | n5239;
  assign n32913 = n5248 | n5249;
  assign n32914 = n5260 | n5261;
  assign n32915 = n5265 | n5266;
  assign n32916 = n5272 | n5273;
  assign n32917 = n5286 | n5287;
  assign n32918 = n5293 | n5294;
  assign n32919 = n5299 | n5300;
  assign n32920 = n5312 | n5313;
  assign n32921 = n5319 | n5320;
  assign n32922 = n5325 | n5326;
  assign n32923 = n5335 | n5336;
  assign n32924 = n5343 | ~n5344;
  assign n32925 = n5349 | n5350;
  assign n32926 = n5357 | n5358;
  assign n32927 = n5360 | ~n5361;
  assign n32928 = n5369 | n5370;
  assign n32929 = n5377 | ~n5378;
  assign n32930 = n5383 | n5384;
  assign n32931 = n5393 | ~n5394;
  assign n32932 = n5402 | n5403;
  assign n32933 = n5410 | ~n5411;
  assign n32934 = n5416 | n5417;
  assign n32935 = n5423 | n5424;
  assign n32936 = n5427 | ~n5428;
  assign n32937 = n5436 | n5437;
  assign n32938 = n5444 | ~n5445;
  assign n32939 = n5450 | n5451;
  assign n32940 = n5457 | n5458;
  assign n32941 = n5461 | ~n5462;
  assign n32942 = n5470 | n5471;
  assign n32943 = n5478 | ~n5479;
  assign n32944 = n5484 | n5485;
  assign n32945 = n5488 | n5489;
  assign n32946 = n5491 | n5492;
  assign n32947 = n5497 | ~n5498;
  assign n32948 = n5506 | n5507;
  assign n32949 = n5514 | ~n5515;
  assign n32950 = n5520 | n5521;
  assign n32951 = n5527 | n5528;
  assign n32952 = n5537 | n5538;
  assign n32953 = n5545 | ~n5546;
  assign n32954 = n5551 | n5552;
  assign n32955 = n5555 | n5556;
  assign n32956 = n5558 | n5559;
  assign n32957 = n5564 | ~n5565;
  assign n32958 = n5573 | n5574;
  assign n32959 = n5581 | ~n5582;
  assign n32960 = n5587 | n5588;
  assign n32961 = n5595 | n5596;
  assign n32962 = n5598 | ~n5599;
  assign n32963 = n5607 | n5608;
  assign n32964 = n5615 | ~n5616;
  assign n32965 = n5625 | n5626;
  assign n32966 = n5629 | n5630;
  assign n32967 = n5638 | n5639;
  assign n32968 = n5646 | ~n5647;
  assign n32969 = n5656 | n5657;
  assign n32970 = n5660 | n5661;
  assign n32971 = n5669 | n5670;
  assign n32972 = n5677 | ~n5678;
  assign n32973 = n5683 | n5684;
  assign n32974 = n5691 | ~n5692;
  assign n32975 = n5695 | n5696;
  assign n32976 = n5702 | n5703;
  assign n32977 = n5718 | n5719;
  assign n32978 = n5724 | n5725;
  assign n32979 = n5728 | n5729;
  assign n32980 = n5740 | n5741;
  assign n32981 = n5744 | n5745;
  assign n32982 = n5755 | n5756;
  assign n32983 = n5766 | n5767;
  assign n32984 = n5770 | n5771;
  assign n32985 = n5783 | n5784;
  assign n32986 = n5786 | ~n5787;
  assign n32987 = n5796 | n5797;
  assign n32988 = n5800 | n5801;
  assign n32989 = n5815 | ~n5816;
  assign n32990 = n5825 | n5826;
  assign n32991 = n5829 | n5830;
  assign n32992 = n5841 | n5842;
  assign n32993 = n5845 | ~n5846;
  assign n32994 = n5855 | n5856;
  assign n32995 = n5859 | n5860;
  assign n32996 = n5871 | n5872;
  assign n32997 = n5875 | ~n5876;
  assign n32998 = n5885 | n5886;
  assign n32999 = n5889 | n5890;
  assign n33000 = n5898 | n5899;
  assign n33001 = n5901 | n5902;
  assign n33002 = n5907 | ~n5908;
  assign n33003 = n5917 | n5918;
  assign n33004 = n5921 | n5922;
  assign n33005 = n5933 | n5934;
  assign n33006 = n5944 | n5945;
  assign n33007 = n5948 | n5949;
  assign n33008 = n5957 | n5958;
  assign n33009 = n5960 | n5961;
  assign n33010 = n5966 | ~n5967;
  assign n33011 = n5976 | n5977;
  assign n33012 = n5980 | n5981;
  assign n33013 = n5993 | n5994;
  assign n33014 = n5996 | ~n5997;
  assign n33015 = n6006 | n6007;
  assign n33016 = n6010 | n6011;
  assign n33017 = n6019 | n6020;
  assign n33018 = n6022 | n6023;
  assign n33019 = n6028 | ~n6029;
  assign n33020 = n6038 | n6039;
  assign n33021 = n6042 | n6043;
  assign n33022 = n6051 | n6052;
  assign n33023 = n6059 | ~n6060;
  assign n33024 = n6069 | n6070;
  assign n33025 = n6073 | n6074;
  assign n33026 = n6082 | n6083;
  assign n33027 = n6090 | ~n6091;
  assign n33028 = n6099 | n6100;
  assign n33029 = n6104 | n6105;
  assign n33030 = n6111 | n6112;
  assign n33031 = n6125 | n6126;
  assign n33032 = n6132 | n6133;
  assign n33033 = n6138 | n6139;
  assign n33034 = n6151 | n6152;
  assign n33035 = n6158 | n6159;
  assign n33036 = n6164 | n6165;
  assign n33037 = n6174 | n6175;
  assign n33038 = n6182 | ~n6183;
  assign n33039 = n6188 | n6189;
  assign n33040 = n6196 | n6197;
  assign n33041 = n6199 | ~n6200;
  assign n33042 = n6208 | n6209;
  assign n33043 = n6216 | ~n6217;
  assign n33044 = n6222 | n6223;
  assign n33045 = n6232 | ~n6233;
  assign n33046 = n6241 | n6242;
  assign n33047 = n6249 | ~n6250;
  assign n33048 = n6255 | n6256;
  assign n33049 = n6262 | n6263;
  assign n33050 = n6266 | ~n6267;
  assign n33051 = n6275 | n6276;
  assign n33052 = n6283 | ~n6284;
  assign n33053 = n6289 | n6290;
  assign n33054 = n6296 | n6297;
  assign n33055 = n6300 | ~n6301;
  assign n33056 = n6309 | n6310;
  assign n33057 = n6317 | ~n6318;
  assign n33058 = n6323 | n6324;
  assign n33059 = n6327 | n6328;
  assign n33060 = n6330 | n6331;
  assign n33061 = n6336 | ~n6337;
  assign n33062 = n6345 | n6346;
  assign n33063 = n6353 | ~n6354;
  assign n33064 = n6359 | n6360;
  assign n33065 = n6366 | n6367;
  assign n33066 = n6376 | n6377;
  assign n33067 = n6384 | ~n6385;
  assign n33068 = n6390 | n6391;
  assign n33069 = n6394 | n6395;
  assign n33070 = n6397 | n6398;
  assign n33071 = n6403 | ~n6404;
  assign n33072 = n6412 | n6413;
  assign n33073 = n6420 | ~n6421;
  assign n33074 = n6426 | n6427;
  assign n33075 = n6434 | n6435;
  assign n33076 = n6437 | ~n6438;
  assign n33077 = n6446 | n6447;
  assign n33078 = n6454 | ~n6455;
  assign n33079 = n6460 | n6461;
  assign n33080 = n6464 | n6465;
  assign n33081 = n6467 | n6468;
  assign n33082 = n6473 | ~n6474;
  assign n33083 = n6482 | n6483;
  assign n33084 = n6490 | ~n6491;
  assign n33085 = n6500 | n6501;
  assign n33086 = n6504 | n6505;
  assign n33087 = n6513 | n6514;
  assign n33088 = n6521 | ~n6522;
  assign n33089 = n6531 | n6532;
  assign n33090 = n6535 | n6536;
  assign n33091 = n6544 | n6545;
  assign n33092 = n6552 | ~n6553;
  assign n33093 = n6561 | n6562;
  assign n33094 = n6566 | n6567;
  assign n33095 = n6573 | n6574;
  assign n33096 = n6589 | n6590;
  assign n33097 = n6595 | n6596;
  assign n33098 = n6599 | n6600;
  assign n33099 = n6611 | n6612;
  assign n33100 = n6615 | n6616;
  assign n33101 = n6626 | n6627;
  assign n33102 = n6637 | n6638;
  assign n33103 = n6641 | n6642;
  assign n33104 = n6654 | n6655;
  assign n33105 = n6657 | ~n6658;
  assign n33106 = n6667 | n6668;
  assign n33107 = n6671 | n6672;
  assign n33108 = n6686 | ~n6687;
  assign n33109 = n6696 | n6697;
  assign n33110 = n6700 | n6701;
  assign n33111 = n6712 | n6713;
  assign n33112 = n6716 | ~n6717;
  assign n33113 = n6726 | n6727;
  assign n33114 = n6730 | n6731;
  assign n33115 = n6742 | n6743;
  assign n33116 = n6746 | ~n6747;
  assign n33117 = n6756 | n6757;
  assign n33118 = n6760 | n6761;
  assign n33119 = n6769 | n6770;
  assign n33120 = n6772 | n6773;
  assign n33121 = n6778 | ~n6779;
  assign n33122 = n6788 | n6789;
  assign n33123 = n6792 | n6793;
  assign n33124 = n6804 | n6805;
  assign n33125 = n6815 | n6816;
  assign n33126 = n6819 | n6820;
  assign n33127 = n6828 | n6829;
  assign n33128 = n6831 | n6832;
  assign n33129 = n6837 | ~n6838;
  assign n33130 = n6847 | n6848;
  assign n33131 = n6851 | n6852;
  assign n33132 = n6864 | n6865;
  assign n33133 = n6867 | ~n6868;
  assign n33134 = n6877 | n6878;
  assign n33135 = n6881 | n6882;
  assign n33136 = n6890 | n6891;
  assign n33137 = n6893 | n6894;
  assign n33138 = n6899 | ~n6900;
  assign n33139 = n6909 | n6910;
  assign n33140 = n6913 | n6914;
  assign n33141 = n6923 | n6924;
  assign n33142 = n6936 | n6937;
  assign n33143 = n6940 | n6941;
  assign n33144 = n6949 | n6950;
  assign n33145 = n6957 | ~n6958;
  assign n33146 = n6967 | n6968;
  assign n33147 = n6971 | n6972;
  assign n33148 = n6980 | n6981;
  assign n33149 = n6988 | ~n6989;
  assign n33150 = n6997 | n6998;
  assign n33151 = n7002 | n7003;
  assign n33152 = n7009 | n7010;
  assign n33153 = n7023 | n7024;
  assign n33154 = n7030 | n7031;
  assign n33155 = n7036 | n7037;
  assign n33156 = n7049 | n7050;
  assign n33157 = n7056 | n7057;
  assign n33158 = n7062 | n7063;
  assign n33159 = n7072 | n7073;
  assign n33160 = n7080 | ~n7081;
  assign n33161 = n7086 | n7087;
  assign n33162 = n7094 | n7095;
  assign n33163 = n7097 | ~n7098;
  assign n33164 = n7106 | n7107;
  assign n33165 = n7114 | ~n7115;
  assign n33166 = n7120 | n7121;
  assign n33167 = n7130 | ~n7131;
  assign n33168 = n7139 | n7140;
  assign n33169 = n7147 | ~n7148;
  assign n33170 = n7153 | n7154;
  assign n33171 = n7160 | n7161;
  assign n33172 = n7164 | ~n7165;
  assign n33173 = n7173 | n7174;
  assign n33174 = n7181 | ~n7182;
  assign n33175 = n7187 | n7188;
  assign n33176 = n7194 | n7195;
  assign n33177 = n7198 | ~n7199;
  assign n33178 = n7207 | n7208;
  assign n33179 = n7215 | ~n7216;
  assign n33180 = n7221 | n7222;
  assign n33181 = n7225 | n7226;
  assign n33182 = n7228 | n7229;
  assign n33183 = n7234 | ~n7235;
  assign n33184 = n7243 | n7244;
  assign n33185 = n7251 | ~n7252;
  assign n33186 = n7257 | n7258;
  assign n33187 = n7264 | n7265;
  assign n33188 = n7274 | n7275;
  assign n33189 = n7282 | ~n7283;
  assign n33190 = n7288 | n7289;
  assign n33191 = n7292 | n7293;
  assign n33192 = n7295 | n7296;
  assign n33193 = n7301 | ~n7302;
  assign n33194 = n7310 | n7311;
  assign n33195 = n7318 | ~n7319;
  assign n33196 = n7324 | n7325;
  assign n33197 = n7332 | n7333;
  assign n33198 = n7335 | ~n7336;
  assign n33199 = n7344 | n7345;
  assign n33200 = n7352 | ~n7353;
  assign n33201 = n7358 | n7359;
  assign n33202 = n7362 | n7363;
  assign n33203 = n7365 | n7366;
  assign n33204 = n7371 | ~n7372;
  assign n33205 = n7380 | n7381;
  assign n33206 = n7388 | ~n7389;
  assign n33207 = n7398 | n7399;
  assign n33208 = n7402 | n7403;
  assign n33209 = n7411 | n7412;
  assign n33210 = n7419 | ~n7420;
  assign n33211 = n7425 | n7426;
  assign n33212 = n7429 | n7430;
  assign n33213 = n7437 | ~n7438;
  assign n33214 = n7446 | n7447;
  assign n33215 = n7454 | ~n7455;
  assign n33216 = n7464 | n7465;
  assign n33217 = n7468 | n7469;
  assign n33218 = n7477 | n7478;
  assign n33219 = n7485 | ~n7486;
  assign n33220 = n7494 | n7495;
  assign n33221 = n7499 | n7500;
  assign n33222 = n7506 | n7507;
  assign n33223 = n7522 | n7523;
  assign n33224 = n7528 | n7529;
  assign n33225 = n7532 | n7533;
  assign n33226 = n7544 | n7545;
  assign n33227 = n7548 | n7549;
  assign n33228 = n7559 | n7560;
  assign n33229 = n7570 | n7571;
  assign n33230 = n7574 | n7575;
  assign n33231 = n7587 | n7588;
  assign n33232 = n7590 | ~n7591;
  assign n33233 = n7600 | n7601;
  assign n33234 = n7604 | n7605;
  assign n33235 = n7619 | ~n7620;
  assign n33236 = n7629 | n7630;
  assign n33237 = n7633 | n7634;
  assign n33238 = n7645 | n7646;
  assign n33239 = n7649 | ~n7650;
  assign n33240 = n7659 | n7660;
  assign n33241 = n7663 | n7664;
  assign n33242 = n7675 | n7676;
  assign n33243 = n7679 | ~n7680;
  assign n33244 = n7689 | n7690;
  assign n33245 = n7693 | n7694;
  assign n33246 = n7702 | n7703;
  assign n33247 = n7705 | n7706;
  assign n33248 = n7711 | ~n7712;
  assign n33249 = n7721 | n7722;
  assign n33250 = n7725 | n7726;
  assign n33251 = n7737 | n7738;
  assign n33252 = n7748 | n7749;
  assign n33253 = n7752 | n7753;
  assign n33254 = n7761 | n7762;
  assign n33255 = n7764 | n7765;
  assign n33256 = n7770 | ~n7771;
  assign n33257 = n7780 | n7781;
  assign n33258 = n7784 | n7785;
  assign n33259 = n7797 | n7798;
  assign n33260 = n7800 | ~n7801;
  assign n33261 = n7810 | n7811;
  assign n33262 = n7814 | n7815;
  assign n33263 = n7823 | n7824;
  assign n33264 = n7826 | n7827;
  assign n33265 = n7832 | ~n7833;
  assign n33266 = n7842 | n7843;
  assign n33267 = n7846 | n7847;
  assign n33268 = n7856 | n7857;
  assign n33269 = n7869 | n7870;
  assign n33270 = n7873 | n7874;
  assign n33271 = n7882 | n7883;
  assign n33272 = n7890 | ~n7891;
  assign n33273 = n7900 | n7901;
  assign n33274 = n7904 | n7905;
  assign n33275 = n7914 | n7915;
  assign n33276 = n7927 | n7928;
  assign n33277 = n7931 | n7932;
  assign n33278 = n7940 | n7941;
  assign n33279 = n7948 | ~n7949;
  assign n33280 = n7957 | n7958;
  assign n33281 = n7962 | n7963;
  assign n33282 = n7969 | n7970;
  assign n33283 = n7982 | n7983;
  assign n33284 = n7989 | n7990;
  assign n33285 = n7995 | n7996;
  assign n33286 = n8008 | n8009;
  assign n33287 = n8015 | n8016;
  assign n33288 = n8021 | n8022;
  assign n33289 = n8031 | n8032;
  assign n33290 = n8039 | ~n8040;
  assign n33291 = n8045 | n8046;
  assign n33292 = n8053 | n8054;
  assign n33293 = n8056 | ~n8057;
  assign n33294 = n8065 | n8066;
  assign n33295 = n8073 | ~n8074;
  assign n33296 = n8079 | n8080;
  assign n33297 = n8089 | ~n8090;
  assign n33298 = n8098 | n8099;
  assign n33299 = n8106 | ~n8107;
  assign n33300 = n8112 | n8113;
  assign n33301 = n8119 | n8120;
  assign n33302 = n8123 | ~n8124;
  assign n33303 = n8132 | n8133;
  assign n33304 = n8140 | ~n8141;
  assign n33305 = n8146 | n8147;
  assign n33306 = n8153 | n8154;
  assign n33307 = n8157 | ~n8158;
  assign n33308 = n8166 | n8167;
  assign n33309 = n8174 | ~n8175;
  assign n33310 = n8180 | n8181;
  assign n33311 = n8184 | n8185;
  assign n33312 = n8187 | n8188;
  assign n33313 = n8193 | ~n8194;
  assign n33314 = n8202 | n8203;
  assign n33315 = n8210 | ~n8211;
  assign n33316 = n8216 | n8217;
  assign n33317 = n8223 | n8224;
  assign n33318 = n8233 | n8234;
  assign n33319 = n8241 | ~n8242;
  assign n33320 = n8247 | n8248;
  assign n33321 = n8251 | n8252;
  assign n33322 = n8254 | n8255;
  assign n33323 = n8260 | ~n8261;
  assign n33324 = n8269 | n8270;
  assign n33325 = n8277 | ~n8278;
  assign n33326 = n8283 | n8284;
  assign n33327 = n8291 | n8292;
  assign n33328 = n8294 | ~n8295;
  assign n33329 = n8303 | n8304;
  assign n33330 = n8311 | ~n8312;
  assign n33331 = n8317 | n8318;
  assign n33332 = n8321 | n8322;
  assign n33333 = n8324 | n8325;
  assign n33334 = n8330 | ~n8331;
  assign n33335 = n8339 | n8340;
  assign n33336 = n8347 | ~n8348;
  assign n33337 = n8357 | n8358;
  assign n33338 = n8361 | n8362;
  assign n33339 = n8370 | n8371;
  assign n33340 = n8378 | ~n8379;
  assign n33341 = n8384 | n8385;
  assign n33342 = n8388 | n8389;
  assign n33343 = n8396 | ~n8397;
  assign n33344 = n8405 | n8406;
  assign n33345 = n8413 | ~n8414;
  assign n33346 = n8423 | n8424;
  assign n33347 = n8427 | n8428;
  assign n33348 = n8436 | n8437;
  assign n33349 = n8444 | ~n8445;
  assign n33350 = n8450 | n8451;
  assign n33351 = n8454 | n8455;
  assign n33352 = n8462 | ~n8463;
  assign n33353 = n8471 | n8472;
  assign n33354 = n8479 | ~n8480;
  assign n33355 = n8488 | n8489;
  assign n33356 = n8493 | n8494;
  assign n33357 = n8500 | n8501;
  assign n33358 = n8508 | n8509;
  assign n33359 = n8516 | n8517;
  assign n33360 = n8528 | n8529;
  assign n33361 = n8534 | n8535;
  assign n33362 = n8542 | n8543;
  assign n33363 = n8553 | n8554;
  assign n33364 = n8555 | n8556;
  assign n33365 = n8566 | n8567;
  assign n33366 = n8570 | n8571;
  assign n33367 = n8583 | n8584;
  assign n33368 = n8586 | ~n8587;
  assign n33369 = n8596 | n8597;
  assign n33370 = n8600 | n8601;
  assign n33371 = n8615 | ~n8616;
  assign n33372 = n8625 | n8626;
  assign n33373 = n8629 | n8630;
  assign n33374 = n8641 | n8642;
  assign n33375 = n8645 | ~n8646;
  assign n33376 = n8655 | n8656;
  assign n33377 = n8659 | n8660;
  assign n33378 = n8671 | n8672;
  assign n33379 = n8675 | ~n8676;
  assign n33380 = n8685 | n8686;
  assign n33381 = n8689 | n8690;
  assign n33382 = n8698 | n8699;
  assign n33383 = n8701 | n8702;
  assign n33384 = n8707 | ~n8708;
  assign n33385 = n8717 | n8718;
  assign n33386 = n8721 | n8722;
  assign n33387 = n8733 | n8734;
  assign n33388 = n8744 | n8745;
  assign n33389 = n8748 | n8749;
  assign n33390 = n8757 | n8758;
  assign n33391 = n8760 | n8761;
  assign n33392 = n8766 | ~n8767;
  assign n33393 = n8776 | n8777;
  assign n33394 = n8780 | n8781;
  assign n33395 = n8793 | n8794;
  assign n33396 = n8796 | ~n8797;
  assign n33397 = n8806 | n8807;
  assign n33398 = n8810 | n8811;
  assign n33399 = n8819 | n8820;
  assign n33400 = n8822 | n8823;
  assign n33401 = n8828 | ~n8829;
  assign n33402 = n8838 | n8839;
  assign n33403 = n8842 | n8843;
  assign n33404 = n8852 | n8853;
  assign n33405 = n8865 | n8866;
  assign n33406 = n8869 | n8870;
  assign n33407 = n8878 | n8879;
  assign n33408 = n8886 | ~n8887;
  assign n33409 = n8896 | n8897;
  assign n33410 = n8900 | n8901;
  assign n33411 = n8910 | n8911;
  assign n33412 = n8923 | n8924;
  assign n33413 = n8927 | n8928;
  assign n33414 = n8936 | n8937;
  assign n33415 = n8944 | ~n8945;
  assign n33416 = n8954 | n8955;
  assign n33417 = n8958 | n8959;
  assign n33418 = n8968 | n8969;
  assign n33419 = n8980 | n8981;
  assign n33420 = n8985 | n8986;
  assign n33421 = n8992 | n8993;
  assign n33422 = n9001 | n9002;
  assign n33423 = n9009 | ~n9010;
  assign n33424 = n9018 | n9019;
  assign n33425 = n9025 | n9026;
  assign n33426 = n9031 | n9032;
  assign n33427 = n9044 | n9045;
  assign n33428 = n9051 | n9052;
  assign n33429 = n9057 | n9058;
  assign n33430 = n9069 | n9070;
  assign n33431 = n9077 | n9078;
  assign n33432 = n9080 | ~n9081;
  assign n33433 = n9089 | n9090;
  assign n33434 = n9097 | ~n9098;
  assign n33435 = n9103 | n9104;
  assign n33436 = n9113 | ~n9114;
  assign n33437 = n9122 | n9123;
  assign n33438 = n9130 | ~n9131;
  assign n33439 = n9136 | n9137;
  assign n33440 = n9143 | n9144;
  assign n33441 = n9147 | ~n9148;
  assign n33442 = n9156 | n9157;
  assign n33443 = n9164 | ~n9165;
  assign n33444 = n9170 | n9171;
  assign n33445 = n9177 | n9178;
  assign n33446 = n9181 | ~n9182;
  assign n33447 = n9190 | n9191;
  assign n33448 = n9198 | ~n9199;
  assign n33449 = n9204 | n9205;
  assign n33450 = n9208 | n9209;
  assign n33451 = n9211 | n9212;
  assign n33452 = n9217 | ~n9218;
  assign n33453 = n9226 | n9227;
  assign n33454 = n9234 | ~n9235;
  assign n33455 = n9240 | n9241;
  assign n33456 = n9247 | n9248;
  assign n33457 = n9257 | n9258;
  assign n33458 = n9265 | ~n9266;
  assign n33459 = n9271 | n9272;
  assign n33460 = n9275 | n9276;
  assign n33461 = n9278 | n9279;
  assign n33462 = n9284 | ~n9285;
  assign n33463 = n9293 | n9294;
  assign n33464 = n9301 | ~n9302;
  assign n33465 = n9307 | n9308;
  assign n33466 = n9315 | n9316;
  assign n33467 = n9318 | ~n9319;
  assign n33468 = n9327 | n9328;
  assign n33469 = n9335 | ~n9336;
  assign n33470 = n9341 | n9342;
  assign n33471 = n9345 | n9346;
  assign n33472 = n9348 | n9349;
  assign n33473 = n9354 | ~n9355;
  assign n33474 = n9363 | n9364;
  assign n33475 = n9371 | ~n9372;
  assign n33476 = n9381 | n9382;
  assign n33477 = n9385 | n9386;
  assign n33478 = n9394 | n9395;
  assign n33479 = n9402 | ~n9403;
  assign n33480 = n9408 | n9409;
  assign n33481 = n9412 | n9413;
  assign n33482 = n9420 | ~n9421;
  assign n33483 = n9429 | n9430;
  assign n33484 = n9437 | ~n9438;
  assign n33485 = n9447 | n9448;
  assign n33486 = n9451 | n9452;
  assign n33487 = n9460 | n9461;
  assign n33488 = n9468 | ~n9469;
  assign n33489 = n9474 | n9475;
  assign n33490 = n9478 | n9479;
  assign n33491 = n9486 | ~n9487;
  assign n33492 = n9495 | n9496;
  assign n33493 = n9503 | ~n9504;
  assign n33494 = n9513 | n9514;
  assign n33495 = n9517 | n9518;
  assign n33496 = n9526 | n9527;
  assign n33497 = n9534 | ~n9535;
  assign n33498 = n9540 | n9541;
  assign n33499 = n9548 | ~n9549;
  assign n33500 = n9552 | n9553;
  assign n33501 = n9559 | n9560;
  assign n33502 = n9571 | n9572;
  assign n33503 = n9579 | n9580;
  assign n33504 = n9583 | n9584;
  assign n33505 = n9591 | n9592;
  assign n33506 = n9601 | n9602;
  assign n33507 = n9608 | n9609;
  assign n33508 = n9616 | n9617;
  assign n33509 = n9626 | n9627;
  assign n33510 = n9634 | n9635;
  assign n33511 = n9648 | n9649;
  assign n33512 = n9651 | ~n9652;
  assign n33513 = n9657 | n9658;
  assign n33514 = n9672 | ~n9673;
  assign n33515 = n9682 | n9683;
  assign n33516 = n9686 | n9687;
  assign n33517 = n9698 | n9699;
  assign n33518 = n9702 | ~n9703;
  assign n33519 = n9712 | n9713;
  assign n33520 = n9716 | n9717;
  assign n33521 = n9728 | n9729;
  assign n33522 = n9732 | ~n9733;
  assign n33523 = n9742 | n9743;
  assign n33524 = n9746 | n9747;
  assign n33525 = n9755 | n9756;
  assign n33526 = n9758 | n9759;
  assign n33527 = n9764 | ~n9765;
  assign n33528 = n9774 | n9775;
  assign n33529 = n9778 | n9779;
  assign n33530 = n9790 | n9791;
  assign n33531 = n9801 | n9802;
  assign n33532 = n9805 | n9806;
  assign n33533 = n9814 | n9815;
  assign n33534 = n9817 | n9818;
  assign n33535 = n9823 | ~n9824;
  assign n33536 = n9833 | n9834;
  assign n33537 = n9837 | n9838;
  assign n33538 = n9850 | n9851;
  assign n33539 = n9853 | ~n9854;
  assign n33540 = n9863 | n9864;
  assign n33541 = n9867 | n9868;
  assign n33542 = n9876 | n9877;
  assign n33543 = n9879 | n9880;
  assign n33544 = n9885 | ~n9886;
  assign n33545 = n9895 | n9896;
  assign n33546 = n9899 | n9900;
  assign n33547 = n9909 | n9910;
  assign n33548 = n9922 | n9923;
  assign n33549 = n9926 | n9927;
  assign n33550 = n9935 | n9936;
  assign n33551 = n9943 | ~n9944;
  assign n33552 = n9953 | n9954;
  assign n33553 = n9957 | n9958;
  assign n33554 = n9967 | n9968;
  assign n33555 = n9980 | n9981;
  assign n33556 = n9984 | n9985;
  assign n33557 = n9993 | n9994;
  assign n33558 = n10001 | ~n10002;
  assign n33559 = n10011 | n10012;
  assign n33560 = n10015 | n10016;
  assign n33561 = n10025 | n10026;
  assign n33562 = n10038 | n10039;
  assign n33563 = n10042 | n10043;
  assign n33564 = n10051 | n10052;
  assign n33565 = n10059 | ~n10060;
  assign n33566 = n10068 | n10069;
  assign n33567 = n10073 | n10074;
  assign n33568 = n10080 | n10081;
  assign n33569 = n10089 | n10090;
  assign n33570 = n10097 | ~n10098;
  assign n33571 = n10106 | n10107;
  assign n33572 = n10113 | n10114;
  assign n33573 = n10119 | n10120;
  assign n33574 = n10132 | n10133;
  assign n33575 = n10139 | n10140;
  assign n33576 = n10145 | n10146;
  assign n33577 = n10155 | n10156;
  assign n33578 = n10163 | ~n10164;
  assign n33579 = n10169 | n10170;
  assign n33580 = n10177 | n10178;
  assign n33581 = n10180 | ~n10181;
  assign n33582 = n10191 | n10192;
  assign n33583 = n10199 | n10200;
  assign n33584 = n10207 | n10208;
  assign n33585 = n10210 | ~n10211;
  assign n33586 = n10221 | n10222;
  assign n33587 = n10228 | n10229;
  assign n33588 = n10232 | ~n10233;
  assign n33589 = n10241 | n10242;
  assign n33590 = n10249 | ~n10250;
  assign n33591 = n10255 | n10256;
  assign n33592 = n10262 | n10263;
  assign n33593 = n10266 | ~n10267;
  assign n33594 = n10275 | n10276;
  assign n33595 = n10283 | ~n10284;
  assign n33596 = n10289 | n10290;
  assign n33597 = n10293 | n10294;
  assign n33598 = n10296 | n10297;
  assign n33599 = n10302 | ~n10303;
  assign n33600 = n10311 | n10312;
  assign n33601 = n10319 | ~n10320;
  assign n33602 = n10325 | n10326;
  assign n33603 = n10332 | n10333;
  assign n33604 = n10342 | n10343;
  assign n33605 = n10350 | ~n10351;
  assign n33606 = n10356 | n10357;
  assign n33607 = n10360 | n10361;
  assign n33608 = n10363 | n10364;
  assign n33609 = n10369 | ~n10370;
  assign n33610 = n10378 | n10379;
  assign n33611 = n10386 | ~n10387;
  assign n33612 = n10392 | n10393;
  assign n33613 = n10400 | n10401;
  assign n33614 = n10403 | ~n10404;
  assign n33615 = n10412 | n10413;
  assign n33616 = n10420 | ~n10421;
  assign n33617 = n10426 | n10427;
  assign n33618 = n10430 | n10431;
  assign n33619 = n10433 | n10434;
  assign n33620 = n10439 | ~n10440;
  assign n33621 = n10448 | n10449;
  assign n33622 = n10456 | ~n10457;
  assign n33623 = n10466 | n10467;
  assign n33624 = n10470 | n10471;
  assign n33625 = n10479 | n10480;
  assign n33626 = n10487 | ~n10488;
  assign n33627 = n10493 | n10494;
  assign n33628 = n10497 | n10498;
  assign n33629 = n10505 | ~n10506;
  assign n33630 = n10514 | n10515;
  assign n33631 = n10522 | ~n10523;
  assign n33632 = n10532 | n10533;
  assign n33633 = n10536 | n10537;
  assign n33634 = n10545 | n10546;
  assign n33635 = n10553 | ~n10554;
  assign n33636 = n10559 | n10560;
  assign n33637 = n10563 | n10564;
  assign n33638 = n10571 | ~n10572;
  assign n33639 = n10580 | n10581;
  assign n33640 = n10588 | ~n10589;
  assign n33641 = n10598 | n10599;
  assign n33642 = n10602 | n10603;
  assign n33643 = n10611 | n10612;
  assign n33644 = n10619 | ~n10620;
  assign n33645 = n10625 | n10626;
  assign n33646 = n10629 | n10630;
  assign n33647 = n10637 | ~n10638;
  assign n33648 = n10646 | n10647;
  assign n33649 = n10654 | ~n10655;
  assign n33650 = n10663 | n10664;
  assign n33651 = n10668 | n10669;
  assign n33652 = n10675 | n10676;
  assign n33653 = n10687 | n10688;
  assign n33654 = n10695 | n10696;
  assign n33655 = n10703 | n10704;
  assign n33656 = n10711 | n10712;
  assign n33657 = n10715 | n10716;
  assign n33658 = n10723 | n10724;
  assign n33659 = n10733 | n10734;
  assign n33660 = n10740 | n10741;
  assign n33661 = n10748 | n10749;
  assign n33662 = n10758 | n10759;
  assign n33663 = n10766 | n10767;
  assign n33664 = n10778 | n10779;
  assign n33665 = n10781 | ~n10782;
  assign n33666 = n10788 | n10789;
  assign n33667 = n10802 | ~n10803;
  assign n33668 = n10809 | n10810;
  assign n33669 = n10822 | n10823;
  assign n33670 = n10826 | ~n10827;
  assign n33671 = n10832 | n10833;
  assign n33672 = n10845 | n10846;
  assign n33673 = n10848 | ~n10849;
  assign n33674 = n10858 | n10859;
  assign n33675 = n10862 | n10863;
  assign n33676 = n10871 | n10872;
  assign n33677 = n10874 | n10875;
  assign n33678 = n10880 | ~n10881;
  assign n33679 = n10890 | n10891;
  assign n33680 = n10894 | n10895;
  assign n33681 = n10906 | n10907;
  assign n33682 = n10917 | n10918;
  assign n33683 = n10921 | n10922;
  assign n33684 = n10930 | n10931;
  assign n33685 = n10933 | n10934;
  assign n33686 = n10939 | ~n10940;
  assign n33687 = n10949 | n10950;
  assign n33688 = n10953 | n10954;
  assign n33689 = n10966 | n10967;
  assign n33690 = n10969 | ~n10970;
  assign n33691 = n10979 | n10980;
  assign n33692 = n10983 | n10984;
  assign n33693 = n10992 | n10993;
  assign n33694 = n10995 | n10996;
  assign n33695 = n11001 | ~n11002;
  assign n33696 = n11011 | n11012;
  assign n33697 = n11015 | n11016;
  assign n33698 = n11025 | n11026;
  assign n33699 = n11038 | n11039;
  assign n33700 = n11042 | n11043;
  assign n33701 = n11051 | n11052;
  assign n33702 = n11059 | ~n11060;
  assign n33703 = n11069 | n11070;
  assign n33704 = n11073 | n11074;
  assign n33705 = n11083 | n11084;
  assign n33706 = n11096 | n11097;
  assign n33707 = n11100 | n11101;
  assign n33708 = n11109 | n11110;
  assign n33709 = n11117 | ~n11118;
  assign n33710 = n11127 | n11128;
  assign n33711 = n11131 | n11132;
  assign n33712 = n11141 | n11142;
  assign n33713 = n11154 | n11155;
  assign n33714 = n11158 | n11159;
  assign n33715 = n11167 | n11168;
  assign n33716 = n11175 | ~n11176;
  assign n33717 = n11185 | n11186;
  assign n33718 = n11189 | n11190;
  assign n33719 = n11199 | n11200;
  assign n33720 = n11211 | n11212;
  assign n33721 = n11216 | n11217;
  assign n33722 = n11223 | n11224;
  assign n33723 = n11232 | n11233;
  assign n33724 = n11240 | ~n11241;
  assign n33725 = n11249 | n11250;
  assign n33726 = n11256 | n11257;
  assign n33727 = n11262 | n11263;
  assign n33728 = n11275 | n11276;
  assign n33729 = n11282 | n11283;
  assign n33730 = n11288 | n11289;
  assign n33731 = n11298 | n11299;
  assign n33732 = n11306 | ~n11307;
  assign n33733 = n11312 | n11313;
  assign n33734 = n11320 | n11321;
  assign n33735 = n11323 | ~n11324;
  assign n33736 = n11332 | n11333;
  assign n33737 = n11340 | ~n11341;
  assign n33738 = n11346 | n11347;
  assign n33739 = n11356 | ~n11357;
  assign n33740 = n11365 | n11366;
  assign n33741 = n11373 | ~n11374;
  assign n33742 = n11379 | n11380;
  assign n33743 = n11386 | n11387;
  assign n33744 = n11390 | ~n11391;
  assign n33745 = n11405 | ~n11406;
  assign n33746 = n11415 | n11416;
  assign n33747 = n11419 | ~n11420;
  assign n33748 = n11422 | n11423;
  assign n33749 = n11433 | n11434;
  assign n33750 = n11441 | n11442;
  assign n33751 = n11444 | ~n11445;
  assign n33752 = n11453 | n11454;
  assign n33753 = n11461 | ~n11462;
  assign n33754 = n11467 | n11468;
  assign n33755 = n11474 | n11475;
  assign n33756 = n11484 | n11485;
  assign n33757 = n11492 | ~n11493;
  assign n33758 = n11498 | n11499;
  assign n33759 = n11502 | n11503;
  assign n33760 = n11505 | n11506;
  assign n33761 = n11511 | ~n11512;
  assign n33762 = n11520 | n11521;
  assign n33763 = n11528 | ~n11529;
  assign n33764 = n11534 | n11535;
  assign n33765 = n11542 | n11543;
  assign n33766 = n11545 | ~n11546;
  assign n33767 = n11554 | n11555;
  assign n33768 = n11562 | ~n11563;
  assign n33769 = n11568 | n11569;
  assign n33770 = n11572 | n11573;
  assign n33771 = n11575 | n11576;
  assign n33772 = n11581 | ~n11582;
  assign n33773 = n11590 | n11591;
  assign n33774 = n11598 | ~n11599;
  assign n33775 = n11608 | n11609;
  assign n33776 = n11612 | n11613;
  assign n33777 = n11621 | n11622;
  assign n33778 = n11629 | ~n11630;
  assign n33779 = n11635 | n11636;
  assign n33780 = n11639 | n11640;
  assign n33781 = n11647 | ~n11648;
  assign n33782 = n11656 | n11657;
  assign n33783 = n11664 | ~n11665;
  assign n33784 = n11674 | n11675;
  assign n33785 = n11678 | n11679;
  assign n33786 = n11687 | n11688;
  assign n33787 = n11695 | ~n11696;
  assign n33788 = n11701 | n11702;
  assign n33789 = n11705 | n11706;
  assign n33790 = n11713 | ~n11714;
  assign n33791 = n11722 | n11723;
  assign n33792 = n11730 | ~n11731;
  assign n33793 = n11740 | n11741;
  assign n33794 = n11744 | n11745;
  assign n33795 = n11753 | n11754;
  assign n33796 = n11761 | ~n11762;
  assign n33797 = n11767 | n11768;
  assign n33798 = n11771 | n11772;
  assign n33799 = n11779 | ~n11780;
  assign n33800 = n11788 | n11789;
  assign n33801 = n11796 | ~n11797;
  assign n33802 = n11806 | n11807;
  assign n33803 = n11810 | n11811;
  assign n33804 = n11819 | n11820;
  assign n33805 = n11827 | ~n11828;
  assign n33806 = n11833 | n11834;
  assign n33807 = n11841 | ~n11842;
  assign n33808 = n11845 | n11846;
  assign n33809 = n11852 | n11853;
  assign n33810 = n11864 | n11865;
  assign n33811 = n11872 | n11873;
  assign n33812 = n11880 | n11881;
  assign n33813 = n11888 | n11889;
  assign n33814 = n11896 | n11897;
  assign n33815 = n11900 | n11901;
  assign n33816 = n11908 | n11909;
  assign n33817 = n11918 | n11919;
  assign n33818 = n11925 | n11926;
  assign n33819 = n11933 | n11934;
  assign n33820 = n11943 | n11944;
  assign n33821 = n11951 | n11952;
  assign n33822 = n11963 | n11964;
  assign n33823 = n11966 | ~n11967;
  assign n33824 = n11973 | n11974;
  assign n33825 = n11987 | ~n11988;
  assign n33826 = n11994 | n11995;
  assign n33827 = n12005 | n12006;
  assign n33828 = n12009 | ~n12010;
  assign n33829 = n12016 | n12017;
  assign n33830 = n12027 | n12028;
  assign n33831 = n12031 | ~n12032;
  assign n33832 = n12038 | n12039;
  assign n33833 = n12048 | ~n12049;
  assign n33834 = n12064 | ~n12065;
  assign n33835 = n12070 | n12071;
  assign n33836 = n12079 | n12080;
  assign n33837 = n12081 | n12082;
  assign n33838 = n12086 | n12087;
  assign n33839 = n12089 | ~n12090;
  assign n33840 = n12099 | n12100;
  assign n33841 = n12103 | n12104;
  assign n33842 = n12112 | n12113;
  assign n33843 = n12115 | n12116;
  assign n33844 = n12121 | ~n12122;
  assign n33845 = n12131 | n12132;
  assign n33846 = n12135 | n12136;
  assign n33847 = n12148 | n12149;
  assign n33848 = n12151 | ~n12152;
  assign n33849 = n12161 | n12162;
  assign n33850 = n12165 | n12166;
  assign n33851 = n12174 | n12175;
  assign n33852 = n12177 | n12178;
  assign n33853 = n12183 | ~n12184;
  assign n33854 = n12193 | n12194;
  assign n33855 = n12197 | n12198;
  assign n33856 = n12207 | n12208;
  assign n33857 = n12220 | n12221;
  assign n33858 = n12224 | n12225;
  assign n33859 = n12233 | n12234;
  assign n33860 = n12241 | ~n12242;
  assign n33861 = n12251 | n12252;
  assign n33862 = n12255 | n12256;
  assign n33863 = n12265 | n12266;
  assign n33864 = n12278 | n12279;
  assign n33865 = n12282 | n12283;
  assign n33866 = n12291 | n12292;
  assign n33867 = n12299 | ~n12300;
  assign n33868 = n12309 | n12310;
  assign n33869 = n12313 | n12314;
  assign n33870 = n12323 | n12324;
  assign n33871 = n12336 | n12337;
  assign n33872 = n12340 | n12341;
  assign n33873 = n12349 | n12350;
  assign n33874 = n12357 | ~n12358;
  assign n33875 = n12367 | n12368;
  assign n33876 = n12371 | n12372;
  assign n33877 = n12381 | n12382;
  assign n33878 = n12394 | n12395;
  assign n33879 = n12398 | n12399;
  assign n33880 = n12407 | n12408;
  assign n33881 = n12415 | ~n12416;
  assign n33882 = n12424 | n12425;
  assign n33883 = n12429 | n12430;
  assign n33884 = n12436 | n12437;
  assign n33885 = n12445 | n12446;
  assign n33886 = n12453 | ~n12454;
  assign n33887 = n12462 | n12463;
  assign n33888 = n12469 | n12470;
  assign n33889 = n12475 | n12476;
  assign n33890 = n12488 | n12489;
  assign n33891 = n12495 | n12496;
  assign n33892 = n12501 | n12502;
  assign n33893 = n12511 | n12512;
  assign n33894 = n12519 | ~n12520;
  assign n33895 = n12525 | n12526;
  assign n33896 = n12533 | n12534;
  assign n33897 = n12536 | ~n12537;
  assign n33898 = n12545 | n12546;
  assign n33899 = n12553 | ~n12554;
  assign n33900 = n12559 | n12560;
  assign n33901 = n12569 | ~n12570;
  assign n33902 = n12578 | n12579;
  assign n33903 = n12586 | ~n12587;
  assign n33904 = n12592 | n12593;
  assign n33905 = n12599 | n12600;
  assign n33906 = n12603 | ~n12604;
  assign n33907 = n12612 | n12613;
  assign n33908 = n12620 | ~n12621;
  assign n33909 = n12626 | n12627;
  assign n33910 = n12633 | n12634;
  assign n33911 = n12637 | ~n12638;
  assign n33912 = n12646 | n12647;
  assign n33913 = n12654 | ~n12655;
  assign n33914 = n12660 | n12661;
  assign n33915 = n12664 | n12665;
  assign n33916 = n12667 | n12668;
  assign n33917 = n12673 | ~n12674;
  assign n33918 = n12688 | ~n12689;
  assign n33919 = n12694 | n12695;
  assign n33920 = n12701 | n12702;
  assign n33921 = n12717 | n12718;
  assign n33922 = n12721 | n12722;
  assign n33923 = n12730 | n12731;
  assign n33924 = n12738 | ~n12739;
  assign n33925 = n12744 | n12745;
  assign n33926 = n12752 | n12753;
  assign n33927 = n12755 | ~n12756;
  assign n33928 = n12764 | n12765;
  assign n33929 = n12772 | ~n12773;
  assign n33930 = n12778 | n12779;
  assign n33931 = n12782 | n12783;
  assign n33932 = n12785 | n12786;
  assign n33933 = n12791 | ~n12792;
  assign n33934 = n12800 | n12801;
  assign n33935 = n12808 | ~n12809;
  assign n33936 = n12818 | n12819;
  assign n33937 = n12822 | n12823;
  assign n33938 = n12831 | n12832;
  assign n33939 = n12839 | ~n12840;
  assign n33940 = n12845 | n12846;
  assign n33941 = n12849 | n12850;
  assign n33942 = n12857 | ~n12858;
  assign n33943 = n12866 | n12867;
  assign n33944 = n12874 | ~n12875;
  assign n33945 = n12884 | n12885;
  assign n33946 = n12888 | n12889;
  assign n33947 = n12897 | n12898;
  assign n33948 = n12905 | ~n12906;
  assign n33949 = n12911 | n12912;
  assign n33950 = n12915 | n12916;
  assign n33951 = n12923 | ~n12924;
  assign n33952 = n12932 | n12933;
  assign n33953 = n12940 | ~n12941;
  assign n33954 = n12950 | n12951;
  assign n33955 = n12954 | n12955;
  assign n33956 = n12963 | n12964;
  assign n33957 = n12971 | ~n12972;
  assign n33958 = n12977 | n12978;
  assign n33959 = n12981 | n12982;
  assign n33960 = n12989 | ~n12990;
  assign n33961 = n12998 | n12999;
  assign n33962 = n13006 | ~n13007;
  assign n33963 = n13016 | n13017;
  assign n33964 = n13020 | n13021;
  assign n33965 = n13029 | n13030;
  assign n33966 = n13037 | ~n13038;
  assign n33967 = n13043 | n13044;
  assign n33968 = n13047 | n13048;
  assign n33969 = n13055 | ~n13056;
  assign n33970 = n13064 | n13065;
  assign n33971 = n13072 | ~n13073;
  assign n33972 = n13081 | n13082;
  assign n33973 = n13086 | n13087;
  assign n33974 = n13093 | n13094;
  assign n33975 = n13105 | n13106;
  assign n33976 = n13113 | n13114;
  assign n33977 = n13121 | n13122;
  assign n33978 = n13129 | n13130;
  assign n33979 = n13137 | n13138;
  assign n33980 = n13145 | n13146;
  assign n33981 = n13153 | n13154;
  assign n33982 = n13161 | n13162;
  assign n33983 = n13165 | n13166;
  assign n33984 = n13173 | n13174;
  assign n33985 = n13183 | n13184;
  assign n33986 = n13190 | n13191;
  assign n33987 = n13198 | n13199;
  assign n33988 = n13208 | n13209;
  assign n33989 = n13216 | n13217;
  assign n33990 = n13228 | n13229;
  assign n33991 = n13231 | ~n13232;
  assign n33992 = n13238 | n13239;
  assign n33993 = n13252 | ~n13253;
  assign n33994 = n13259 | n13260;
  assign n33995 = n13270 | n13271;
  assign n33996 = n13274 | ~n13275;
  assign n33997 = n13281 | n13282;
  assign n33998 = n13292 | n13293;
  assign n33999 = n13296 | ~n13297;
  assign n34000 = n13303 | n13304;
  assign n34001 = n13311 | n13312;
  assign n34002 = n13314 | n13315;
  assign n34003 = n13320 | ~n13321;
  assign n34004 = n13327 | n13328;
  assign n34005 = n13338 | n13339;
  assign n34006 = n13346 | n13347;
  assign n34007 = n13360 | n13361;
  assign n34008 = n13363 | ~n13364;
  assign n34009 = n13369 | n13370;
  assign n34010 = n13378 | n13379;
  assign n34011 = n13386 | ~n13387;
  assign n34012 = n13396 | n13397;
  assign n34013 = n13400 | n13401;
  assign n34014 = n13409 | n13410;
  assign n34015 = n13412 | n13413;
  assign n34016 = n13418 | ~n13419;
  assign n34017 = n13428 | n13429;
  assign n34018 = n13432 | n13433;
  assign n34019 = n13442 | n13443;
  assign n34020 = n13455 | n13456;
  assign n34021 = n13459 | n13460;
  assign n34022 = n13468 | n13469;
  assign n34023 = n13476 | ~n13477;
  assign n34024 = n13486 | n13487;
  assign n34025 = n13490 | n13491;
  assign n34026 = n13500 | n13501;
  assign n34027 = n13513 | n13514;
  assign n34028 = n13517 | n13518;
  assign n34029 = n13526 | n13527;
  assign n34030 = n13534 | ~n13535;
  assign n34031 = n13544 | n13545;
  assign n34032 = n13548 | n13549;
  assign n34033 = n13558 | n13559;
  assign n34034 = n13571 | n13572;
  assign n34035 = n13575 | n13576;
  assign n34036 = n13584 | n13585;
  assign n34037 = n13592 | ~n13593;
  assign n34038 = n13602 | n13603;
  assign n34039 = n13606 | n13607;
  assign n34040 = n13616 | n13617;
  assign n34041 = n13629 | n13630;
  assign n34042 = n13633 | n13634;
  assign n34043 = n13642 | n13643;
  assign n34044 = n13650 | ~n13651;
  assign n34045 = n13660 | n13661;
  assign n34046 = n13664 | n13665;
  assign n34047 = n13674 | n13675;
  assign n34048 = n13686 | n13687;
  assign n34049 = n13691 | n13692;
  assign n34050 = n13698 | n13699;
  assign n34051 = n13707 | n13708;
  assign n34052 = n13715 | ~n13716;
  assign n34053 = n13724 | n13725;
  assign n34054 = n13731 | n13732;
  assign n34055 = n13737 | n13738;
  assign n34056 = n13750 | n13751;
  assign n34057 = n13757 | n13758;
  assign n34058 = n13763 | n13764;
  assign n34059 = n13773 | n13774;
  assign n34060 = n13781 | ~n13782;
  assign n34061 = n13787 | n13788;
  assign n34062 = n13795 | n13796;
  assign n34063 = n13798 | ~n13799;
  assign n34064 = n13807 | n13808;
  assign n34065 = n13815 | ~n13816;
  assign n34066 = n13821 | n13822;
  assign n34067 = n13831 | ~n13832;
  assign n34068 = n13840 | n13841;
  assign n34069 = n13848 | ~n13849;
  assign n34070 = n13854 | n13855;
  assign n34071 = n13861 | n13862;
  assign n34072 = n13865 | ~n13866;
  assign n34073 = n13874 | n13875;
  assign n34074 = n13882 | ~n13883;
  assign n34075 = n13888 | n13889;
  assign n34076 = n13895 | n13896;
  assign n34077 = n13899 | ~n13900;
  assign n34078 = n13908 | n13909;
  assign n34079 = n13916 | ~n13917;
  assign n34080 = n13922 | n13923;
  assign n34081 = n13926 | n13927;
  assign n34082 = n13929 | n13930;
  assign n34083 = n13935 | ~n13936;
  assign n34084 = n13944 | n13945;
  assign n34085 = n13952 | ~n13953;
  assign n34086 = n13958 | n13959;
  assign n34087 = n13965 | n13966;
  assign n34088 = n13975 | n13976;
  assign n34089 = n13983 | ~n13984;
  assign n34090 = n13989 | n13990;
  assign n34091 = n13993 | n13994;
  assign n34092 = n13996 | n13997;
  assign n34093 = n14002 | ~n14003;
  assign n34094 = n14013 | n14014;
  assign n34095 = n14021 | n14022;
  assign n34096 = n14029 | n14030;
  assign n34097 = n14032 | ~n14033;
  assign n34098 = n14047 | n14048;
  assign n34099 = n14051 | n14052;
  assign n34100 = n14060 | n14061;
  assign n34101 = n14068 | ~n14069;
  assign n34102 = n14078 | n14079;
  assign n34103 = n14082 | n14083;
  assign n34104 = n14091 | n14092;
  assign n34105 = n14099 | ~n14100;
  assign n34106 = n14105 | n14106;
  assign n34107 = n14109 | n14110;
  assign n34108 = n14117 | ~n14118;
  assign n34109 = n14126 | n14127;
  assign n34110 = n14134 | ~n14135;
  assign n34111 = n14144 | n14145;
  assign n34112 = n14148 | n14149;
  assign n34113 = n14157 | n14158;
  assign n34114 = n14165 | ~n14166;
  assign n34115 = n14171 | n14172;
  assign n34116 = n14175 | n14176;
  assign n34117 = n14183 | ~n14184;
  assign n34118 = n14192 | n14193;
  assign n34119 = n14200 | ~n14201;
  assign n34120 = n14210 | n14211;
  assign n34121 = n14214 | n14215;
  assign n34122 = n14223 | n14224;
  assign n34123 = n14231 | ~n14232;
  assign n34124 = n14237 | n14238;
  assign n34125 = n14241 | n14242;
  assign n34126 = n14249 | ~n14250;
  assign n34127 = n14258 | n14259;
  assign n34128 = n14266 | ~n14267;
  assign n34129 = n14276 | n14277;
  assign n34130 = n14280 | n14281;
  assign n34131 = n14289 | n14290;
  assign n34132 = n14297 | ~n14298;
  assign n34133 = n14303 | n14304;
  assign n34134 = n14307 | n14308;
  assign n34135 = n14315 | ~n14316;
  assign n34136 = n14324 | n14325;
  assign n34137 = n14332 | ~n14333;
  assign n34138 = n14342 | n14343;
  assign n34139 = n14346 | n14347;
  assign n34140 = n14355 | n14356;
  assign n34141 = n14363 | ~n14364;
  assign n34142 = n14369 | n14370;
  assign n34143 = n14377 | ~n14378;
  assign n34144 = n14381 | n14382;
  assign n34145 = n14388 | n14389;
  assign n34146 = n14400 | n14401;
  assign n34147 = n14408 | n14409;
  assign n34148 = n14416 | n14417;
  assign n34149 = n14424 | n14425;
  assign n34150 = n14432 | n14433;
  assign n34151 = n14440 | n14441;
  assign n34152 = n14448 | n14449;
  assign n34153 = n14456 | n14457;
  assign n34154 = n14464 | n14465;
  assign n34155 = n14472 | n14473;
  assign n34156 = n14476 | n14477;
  assign n34157 = n14484 | n14485;
  assign n34158 = n14494 | n14495;
  assign n34159 = n14501 | n14502;
  assign n34160 = n14509 | n14510;
  assign n34161 = n14519 | n14520;
  assign n34162 = n14527 | n14528;
  assign n34163 = n14539 | n14540;
  assign n34164 = n14542 | ~n14543;
  assign n34165 = n14549 | n14550;
  assign n34166 = n14563 | ~n14564;
  assign n34167 = n14570 | n14571;
  assign n34168 = n14581 | n14582;
  assign n34169 = n14585 | ~n14586;
  assign n34170 = n14592 | n14593;
  assign n34171 = n14603 | n14604;
  assign n34172 = n14607 | ~n14608;
  assign n34173 = n14614 | n14615;
  assign n34174 = n14622 | n14623;
  assign n34175 = n14625 | n14626;
  assign n34176 = n14631 | ~n14632;
  assign n34177 = n14638 | n14639;
  assign n34178 = n14649 | n14650;
  assign n34179 = n14657 | n14658;
  assign n34180 = n14665 | n14666;
  assign n34181 = n14668 | n14669;
  assign n34182 = n14674 | ~n14675;
  assign n34183 = n14681 | n14682;
  assign n34184 = n14693 | n14694;
  assign n34185 = n14696 | ~n14697;
  assign n34186 = n14703 | n14704;
  assign n34187 = n14716 | n14717;
  assign n34188 = n14720 | ~n14721;
  assign n34189 = n14726 | n14727;
  assign n34190 = n14735 | n14736;
  assign n34191 = n14743 | ~n14744;
  assign n34192 = n14753 | n14754;
  assign n34193 = n14757 | n14758;
  assign n34194 = n14766 | n14767;
  assign n34195 = n14774 | ~n14775;
  assign n34196 = n14784 | n14785;
  assign n34197 = n14788 | n14789;
  assign n34198 = n14798 | n14799;
  assign n34199 = n14811 | n14812;
  assign n34200 = n14815 | n14816;
  assign n34201 = n14824 | n14825;
  assign n34202 = n14832 | ~n14833;
  assign n34203 = n14842 | n14843;
  assign n34204 = n14846 | n14847;
  assign n34205 = n14856 | n14857;
  assign n34206 = n14869 | n14870;
  assign n34207 = n14873 | n14874;
  assign n34208 = n14882 | n14883;
  assign n34209 = n14890 | ~n14891;
  assign n34210 = n14900 | n14901;
  assign n34211 = n14904 | n14905;
  assign n34212 = n14914 | n14915;
  assign n34213 = n14927 | n14928;
  assign n34214 = n14931 | n14932;
  assign n34215 = n14940 | n14941;
  assign n34216 = n14948 | ~n14949;
  assign n34217 = n14958 | n14959;
  assign n34218 = n14962 | n14963;
  assign n34219 = n14972 | n14973;
  assign n34220 = n14985 | n14986;
  assign n34221 = n14989 | n14990;
  assign n34222 = n14998 | n14999;
  assign n34223 = n15006 | ~n15007;
  assign n34224 = n15015 | n15016;
  assign n34225 = n15020 | n15021;
  assign n34226 = n15027 | n15028;
  assign n34227 = n15036 | n15037;
  assign n34228 = n15044 | ~n15045;
  assign n34229 = n15053 | n15054;
  assign n34230 = n15060 | n15061;
  assign n34231 = n15066 | n15067;
  assign n34232 = n15079 | n15080;
  assign n34233 = n15086 | n15087;
  assign n34234 = n15092 | n15093;
  assign n34235 = n15102 | n15103;
  assign n34236 = n15110 | ~n15111;
  assign n34237 = n15116 | n15117;
  assign n34238 = n15124 | n15125;
  assign n34239 = n15127 | ~n15128;
  assign n34240 = n15136 | n15137;
  assign n34241 = n15144 | ~n15145;
  assign n34242 = n15150 | n15151;
  assign n34243 = n15160 | ~n15161;
  assign n34244 = n15169 | n15170;
  assign n34245 = n15177 | ~n15178;
  assign n34246 = n15183 | n15184;
  assign n34247 = n15190 | n15191;
  assign n34248 = n15194 | ~n15195;
  assign n34249 = n15203 | n15204;
  assign n34250 = n15211 | ~n15212;
  assign n34251 = n15217 | n15218;
  assign n34252 = n15224 | n15225;
  assign n34253 = n15228 | ~n15229;
  assign n34254 = n15237 | n15238;
  assign n34255 = n15245 | ~n15246;
  assign n34256 = n15251 | n15252;
  assign n34257 = n15255 | n15256;
  assign n34258 = n15258 | n15259;
  assign n34259 = n15264 | ~n15265;
  assign n34260 = n15273 | n15274;
  assign n34261 = n15281 | ~n15282;
  assign n34262 = n15287 | n15288;
  assign n34263 = n15294 | n15295;
  assign n34264 = n15304 | n15305;
  assign n34265 = n15312 | ~n15313;
  assign n34266 = n15318 | n15319;
  assign n34267 = n15322 | n15323;
  assign n34268 = n15325 | n15326;
  assign n34269 = n15331 | ~n15332;
  assign n34270 = n15340 | n15341;
  assign n34271 = n15348 | ~n15349;
  assign n34272 = n15354 | n15355;
  assign n34273 = n15362 | n15363;
  assign n34274 = n15365 | ~n15366;
  assign n34275 = n15374 | n15375;
  assign n34276 = n15382 | ~n15383;
  assign n34277 = n15388 | n15389;
  assign n34278 = n15392 | n15393;
  assign n34279 = n15395 | n15396;
  assign n34280 = n15401 | ~n15402;
  assign n34281 = n15416 | ~n15417;
  assign n34282 = n15426 | n15427;
  assign n34283 = n15430 | ~n15431;
  assign n34284 = n15433 | n15434;
  assign n34285 = n15448 | n15449;
  assign n34286 = n15452 | n15453;
  assign n34287 = n15461 | n15462;
  assign n34288 = n15469 | ~n15470;
  assign n34289 = n15479 | n15480;
  assign n34290 = n15483 | n15484;
  assign n34291 = n15492 | n15493;
  assign n34292 = n15500 | ~n15501;
  assign n34293 = n15506 | n15507;
  assign n34294 = n15510 | n15511;
  assign n34295 = n15518 | ~n15519;
  assign n34296 = n15527 | n15528;
  assign n34297 = n15535 | ~n15536;
  assign n34298 = n15545 | n15546;
  assign n34299 = n15549 | n15550;
  assign n34300 = n15558 | n15559;
  assign n34301 = n15566 | ~n15567;
  assign n34302 = n15572 | n15573;
  assign n34303 = n15576 | n15577;
  assign n34304 = n15584 | ~n15585;
  assign n34305 = n15593 | n15594;
  assign n34306 = n15601 | ~n15602;
  assign n34307 = n15611 | n15612;
  assign n34308 = n15615 | n15616;
  assign n34309 = n15624 | n15625;
  assign n34310 = n15632 | ~n15633;
  assign n34311 = n15638 | n15639;
  assign n34312 = n15642 | n15643;
  assign n34313 = n15650 | ~n15651;
  assign n34314 = n15659 | n15660;
  assign n34315 = n15667 | ~n15668;
  assign n34316 = n15677 | n15678;
  assign n34317 = n15681 | n15682;
  assign n34318 = n15690 | n15691;
  assign n34319 = n15698 | ~n15699;
  assign n34320 = n15704 | n15705;
  assign n34321 = n15708 | n15709;
  assign n34322 = n15716 | ~n15717;
  assign n34323 = n15725 | n15726;
  assign n34324 = n15733 | ~n15734;
  assign n34325 = n15742 | n15743;
  assign n34326 = n15747 | n15748;
  assign n34327 = n15754 | n15755;
  assign n34328 = n15766 | n15767;
  assign n34329 = n15774 | n15775;
  assign n34330 = n15782 | n15783;
  assign n34331 = n15790 | n15791;
  assign n34332 = n15798 | n15799;
  assign n34333 = n15806 | n15807;
  assign n34334 = n15814 | n15815;
  assign n34335 = n15822 | n15823;
  assign n34336 = n15830 | n15831;
  assign n34337 = n15838 | n15839;
  assign n34338 = n15846 | n15847;
  assign n34339 = n15854 | n15855;
  assign n34340 = n15858 | n15859;
  assign n34341 = n15866 | n15867;
  assign n34342 = n15876 | n15877;
  assign n34343 = n15883 | n15884;
  assign n34344 = n15891 | n15892;
  assign n34345 = n15901 | n15902;
  assign n34346 = n15909 | n15910;
  assign n34347 = n15921 | n15922;
  assign n34348 = n15924 | ~n15925;
  assign n34349 = n15931 | n15932;
  assign n34350 = n15945 | ~n15946;
  assign n34351 = n15952 | n15953;
  assign n34352 = n15963 | n15964;
  assign n34353 = n15967 | ~n15968;
  assign n34354 = n15974 | n15975;
  assign n34355 = n15985 | n15986;
  assign n34356 = n15989 | ~n15990;
  assign n34357 = n15996 | n15997;
  assign n34358 = n16004 | n16005;
  assign n34359 = n16007 | n16008;
  assign n34360 = n16013 | ~n16014;
  assign n34361 = n16020 | n16021;
  assign n34362 = n16031 | n16032;
  assign n34363 = n16039 | n16040;
  assign n34364 = n16047 | n16048;
  assign n34365 = n16050 | n16051;
  assign n34366 = n16056 | ~n16057;
  assign n34367 = n16063 | n16064;
  assign n34368 = n16075 | n16076;
  assign n34369 = n16078 | ~n16079;
  assign n34370 = n16085 | n16086;
  assign n34371 = n16093 | n16094;
  assign n34372 = n16096 | n16097;
  assign n34373 = n16102 | ~n16103;
  assign n34374 = n16109 | n16110;
  assign n34375 = n16120 | n16121;
  assign n34376 = n16130 | ~n16131;
  assign n34377 = n16146 | ~n16147;
  assign n34378 = n16152 | n16153;
  assign n34379 = n16161 | n16162;
  assign n34380 = n16169 | ~n16170;
  assign n34381 = n16179 | n16180;
  assign n34382 = n16183 | n16184;
  assign n34383 = n16192 | n16193;
  assign n34384 = n16200 | ~n16201;
  assign n34385 = n16210 | n16211;
  assign n34386 = n16214 | n16215;
  assign n34387 = n16224 | n16225;
  assign n34388 = n16237 | n16238;
  assign n34389 = n16241 | n16242;
  assign n34390 = n16250 | n16251;
  assign n34391 = n16258 | ~n16259;
  assign n34392 = n16268 | n16269;
  assign n34393 = n16272 | n16273;
  assign n34394 = n16282 | n16283;
  assign n34395 = n16295 | n16296;
  assign n34396 = n16299 | n16300;
  assign n34397 = n16308 | n16309;
  assign n34398 = n16316 | ~n16317;
  assign n34399 = n16326 | n16327;
  assign n34400 = n16330 | n16331;
  assign n34401 = n16340 | n16341;
  assign n34402 = n16353 | n16354;
  assign n34403 = n16357 | n16358;
  assign n34404 = n16366 | n16367;
  assign n34405 = n16374 | ~n16375;
  assign n34406 = n16384 | n16385;
  assign n34407 = n16388 | n16389;
  assign n34408 = n16398 | n16399;
  assign n34409 = n16410 | n16411;
  assign n34410 = n16415 | n16416;
  assign n34411 = n16422 | n16423;
  assign n34412 = n16431 | n16432;
  assign n34413 = n16439 | ~n16440;
  assign n34414 = n16448 | n16449;
  assign n34415 = n16455 | n16456;
  assign n34416 = n16461 | n16462;
  assign n34417 = n16474 | n16475;
  assign n34418 = n16481 | n16482;
  assign n34419 = n16487 | n16488;
  assign n34420 = n16497 | n16498;
  assign n34421 = n16505 | ~n16506;
  assign n34422 = n16511 | n16512;
  assign n34423 = n16519 | n16520;
  assign n34424 = n16522 | ~n16523;
  assign n34425 = n16531 | n16532;
  assign n34426 = n16539 | ~n16540;
  assign n34427 = n16545 | n16546;
  assign n34428 = n16555 | ~n16556;
  assign n34429 = n16564 | n16565;
  assign n34430 = n16572 | ~n16573;
  assign n34431 = n16578 | n16579;
  assign n34432 = n16585 | n16586;
  assign n34433 = n16589 | ~n16590;
  assign n34434 = n16598 | n16599;
  assign n34435 = n16606 | ~n16607;
  assign n34436 = n16612 | n16613;
  assign n34437 = n16619 | n16620;
  assign n34438 = n16623 | ~n16624;
  assign n34439 = n16632 | n16633;
  assign n34440 = n16640 | ~n16641;
  assign n34441 = n16646 | n16647;
  assign n34442 = n16650 | n16651;
  assign n34443 = n16653 | n16654;
  assign n34444 = n16659 | ~n16660;
  assign n34445 = n16668 | n16669;
  assign n34446 = n16676 | ~n16677;
  assign n34447 = n16682 | n16683;
  assign n34448 = n16689 | n16690;
  assign n34449 = n16699 | n16700;
  assign n34450 = n16707 | ~n16708;
  assign n34451 = n16713 | n16714;
  assign n34452 = n16717 | n16718;
  assign n34453 = n16720 | n16721;
  assign n34454 = n16726 | ~n16727;
  assign n34455 = n16735 | n16736;
  assign n34456 = n16743 | ~n16744;
  assign n34457 = n16749 | n16750;
  assign n34458 = n16757 | n16758;
  assign n34459 = n16760 | ~n16761;
  assign n34460 = n16769 | n16770;
  assign n34461 = n16777 | ~n16778;
  assign n34462 = n16783 | n16784;
  assign n34463 = n16787 | n16788;
  assign n34464 = n16790 | n16791;
  assign n34465 = n16796 | ~n16797;
  assign n34466 = n16805 | n16806;
  assign n34467 = n16813 | ~n16814;
  assign n34468 = n16823 | n16824;
  assign n34469 = n16827 | n16828;
  assign n34470 = n16836 | n16837;
  assign n34471 = n16844 | ~n16845;
  assign n34472 = n16850 | n16851;
  assign n34473 = n16854 | n16855;
  assign n34474 = n16862 | ~n16863;
  assign n34475 = n16877 | ~n16878;
  assign n34476 = n16883 | n16884;
  assign n34477 = n16890 | n16891;
  assign n34478 = n16906 | n16907;
  assign n34479 = n16910 | n16911;
  assign n34480 = n16919 | n16920;
  assign n34481 = n16927 | ~n16928;
  assign n34482 = n16937 | n16938;
  assign n34483 = n16941 | n16942;
  assign n34484 = n16950 | n16951;
  assign n34485 = n16958 | ~n16959;
  assign n34486 = n16964 | n16965;
  assign n34487 = n16968 | n16969;
  assign n34488 = n16976 | ~n16977;
  assign n34489 = n16985 | n16986;
  assign n34490 = n16993 | ~n16994;
  assign n34491 = n17003 | n17004;
  assign n34492 = n17007 | n17008;
  assign n34493 = n17016 | n17017;
  assign n34494 = n17024 | ~n17025;
  assign n34495 = n17030 | n17031;
  assign n34496 = n17034 | n17035;
  assign n34497 = n17042 | ~n17043;
  assign n34498 = n17051 | n17052;
  assign n34499 = n17059 | ~n17060;
  assign n34500 = n17069 | n17070;
  assign n34501 = n17073 | n17074;
  assign n34502 = n17082 | n17083;
  assign n34503 = n17090 | ~n17091;
  assign n34504 = n17096 | n17097;
  assign n34505 = n17100 | n17101;
  assign n34506 = n17108 | ~n17109;
  assign n34507 = n17117 | n17118;
  assign n34508 = n17125 | ~n17126;
  assign n34509 = n17135 | n17136;
  assign n34510 = n17139 | n17140;
  assign n34511 = n17148 | n17149;
  assign n34512 = n17156 | ~n17157;
  assign n34513 = n17162 | n17163;
  assign n34514 = n17170 | ~n17171;
  assign n34515 = n17174 | n17175;
  assign n34516 = n17181 | n17182;
  assign n34517 = n17193 | n17194;
  assign n34518 = n17201 | n17202;
  assign n34519 = n17209 | n17210;
  assign n34520 = n17217 | n17218;
  assign n34521 = n17225 | n17226;
  assign n34522 = n17233 | n17234;
  assign n34523 = n17241 | n17242;
  assign n34524 = n17249 | n17250;
  assign n34525 = n17257 | n17258;
  assign n34526 = n17265 | n17266;
  assign n34527 = n17273 | n17274;
  assign n34528 = n17281 | n17282;
  assign n34529 = n17289 | n17290;
  assign n34530 = n17297 | n17298;
  assign n34531 = n17305 | n17306;
  assign n34532 = n17313 | n17314;
  assign n34533 = n17317 | n17318;
  assign n34534 = n17325 | n17326;
  assign n34535 = n17335 | n17336;
  assign n34536 = n17342 | n17343;
  assign n34537 = n17350 | n17351;
  assign n34538 = n17360 | n17361;
  assign n34539 = n17368 | n17369;
  assign n34540 = n17380 | n17381;
  assign n34541 = n17383 | ~n17384;
  assign n34542 = n17390 | n17391;
  assign n34543 = n17404 | ~n17405;
  assign n34544 = n17411 | n17412;
  assign n34545 = n17422 | n17423;
  assign n34546 = n17426 | ~n17427;
  assign n34547 = n17433 | n17434;
  assign n34548 = n17444 | n17445;
  assign n34549 = n17448 | ~n17449;
  assign n34550 = n17455 | n17456;
  assign n34551 = n17463 | n17464;
  assign n34552 = n17466 | n17467;
  assign n34553 = n17472 | ~n17473;
  assign n34554 = n17479 | n17480;
  assign n34555 = n17490 | n17491;
  assign n34556 = n17498 | n17499;
  assign n34557 = n17506 | n17507;
  assign n34558 = n17509 | n17510;
  assign n34559 = n17515 | ~n17516;
  assign n34560 = n17522 | n17523;
  assign n34561 = n17534 | n17535;
  assign n34562 = n17537 | ~n17538;
  assign n34563 = n17544 | n17545;
  assign n34564 = n17552 | n17553;
  assign n34565 = n17555 | n17556;
  assign n34566 = n17561 | ~n17562;
  assign n34567 = n17568 | n17569;
  assign n34568 = n17579 | n17580;
  assign n34569 = n17587 | n17588;
  assign n34570 = n17595 | ~n17596;
  assign n34571 = n17602 | n17603;
  assign n34572 = n17613 | n17614;
  assign n34573 = n17627 | n17628;
  assign n34574 = n17630 | ~n17631;
  assign n34575 = n17636 | n17637;
  assign n34576 = n17645 | n17646;
  assign n34577 = n17653 | ~n17654;
  assign n34578 = n17663 | n17664;
  assign n34579 = n17667 | n17668;
  assign n34580 = n17676 | n17677;
  assign n34581 = n17684 | ~n17685;
  assign n34582 = n17694 | n17695;
  assign n34583 = n17698 | n17699;
  assign n34584 = n17708 | n17709;
  assign n34585 = n17721 | n17722;
  assign n34586 = n17725 | n17726;
  assign n34587 = n17734 | n17735;
  assign n34588 = n17742 | ~n17743;
  assign n34589 = n17752 | n17753;
  assign n34590 = n17756 | n17757;
  assign n34591 = n17766 | n17767;
  assign n34592 = n17779 | n17780;
  assign n34593 = n17783 | n17784;
  assign n34594 = n17792 | n17793;
  assign n34595 = n17800 | ~n17801;
  assign n34596 = n17810 | n17811;
  assign n34597 = n17814 | n17815;
  assign n34598 = n17824 | n17825;
  assign n34599 = n17837 | n17838;
  assign n34600 = n17841 | n17842;
  assign n34601 = n17850 | n17851;
  assign n34602 = n17858 | ~n17859;
  assign n34603 = n17867 | n17868;
  assign n34604 = n17872 | n17873;
  assign n34605 = n17879 | n17880;
  assign n34606 = n17888 | n17889;
  assign n34607 = n17896 | ~n17897;
  assign n34608 = n17905 | n17906;
  assign n34609 = n17912 | n17913;
  assign n34610 = n17918 | n17919;
  assign n34611 = n17931 | n17932;
  assign n34612 = n17938 | n17939;
  assign n34613 = n17944 | n17945;
  assign n34614 = n17954 | n17955;
  assign n34615 = n17962 | ~n17963;
  assign n34616 = n17968 | n17969;
  assign n34617 = n17976 | n17977;
  assign n34618 = n17979 | ~n17980;
  assign n34619 = n17988 | n17989;
  assign n34620 = n17996 | ~n17997;
  assign n34621 = n18002 | n18003;
  assign n34622 = n18012 | ~n18013;
  assign n34623 = n18021 | n18022;
  assign n34624 = n18029 | ~n18030;
  assign n34625 = n18035 | n18036;
  assign n34626 = n18042 | n18043;
  assign n34627 = n18046 | ~n18047;
  assign n34628 = n18055 | n18056;
  assign n34629 = n18063 | ~n18064;
  assign n34630 = n18069 | n18070;
  assign n34631 = n18076 | n18077;
  assign n34632 = n18080 | ~n18081;
  assign n34633 = n18089 | n18090;
  assign n34634 = n18097 | ~n18098;
  assign n34635 = n18103 | n18104;
  assign n34636 = n18107 | n18108;
  assign n34637 = n18110 | n18111;
  assign n34638 = n18116 | ~n18117;
  assign n34639 = n18125 | n18126;
  assign n34640 = n18133 | ~n18134;
  assign n34641 = n18139 | n18140;
  assign n34642 = n18146 | n18147;
  assign n34643 = n18156 | n18157;
  assign n34644 = n18164 | ~n18165;
  assign n34645 = n18170 | n18171;
  assign n34646 = n18174 | n18175;
  assign n34647 = n18177 | n18178;
  assign n34648 = n18183 | ~n18184;
  assign n34649 = n18192 | n18193;
  assign n34650 = n18200 | ~n18201;
  assign n34651 = n18206 | n18207;
  assign n34652 = n18214 | n18215;
  assign n34653 = n18217 | ~n18218;
  assign n34654 = n18226 | n18227;
  assign n34655 = n18234 | ~n18235;
  assign n34656 = n18240 | n18241;
  assign n34657 = n18244 | n18245;
  assign n34658 = n18247 | n18248;
  assign n34659 = n18253 | ~n18254;
  assign n34660 = n18262 | n18263;
  assign n34661 = n18270 | ~n18271;
  assign n34662 = n18280 | n18281;
  assign n34663 = n18284 | n18285;
  assign n34664 = n18293 | n18294;
  assign n34665 = n18301 | ~n18302;
  assign n34666 = n18307 | n18308;
  assign n34667 = n18311 | n18312;
  assign n34668 = n18319 | ~n18320;
  assign n34669 = n18328 | n18329;
  assign n34670 = n18336 | ~n18337;
  assign n34671 = n18346 | n18347;
  assign n34672 = n18350 | n18351;
  assign n34673 = n18359 | n18360;
  assign n34674 = n18367 | ~n18368;
  assign n34675 = n18373 | n18374;
  assign n34676 = n18377 | n18378;
  assign n34677 = n18385 | ~n18386;
  assign n34678 = n18396 | n18397;
  assign n34679 = n18404 | n18405;
  assign n34680 = n18412 | n18413;
  assign n34681 = n18415 | ~n18416;
  assign n34682 = n18430 | n18431;
  assign n34683 = n18434 | n18435;
  assign n34684 = n18443 | n18444;
  assign n34685 = n18451 | ~n18452;
  assign n34686 = n18461 | n18462;
  assign n34687 = n18465 | n18466;
  assign n34688 = n18474 | n18475;
  assign n34689 = n18482 | ~n18483;
  assign n34690 = n18488 | n18489;
  assign n34691 = n18492 | n18493;
  assign n34692 = n18500 | ~n18501;
  assign n34693 = n18509 | n18510;
  assign n34694 = n18517 | ~n18518;
  assign n34695 = n18527 | n18528;
  assign n34696 = n18531 | n18532;
  assign n34697 = n18540 | n18541;
  assign n34698 = n18548 | ~n18549;
  assign n34699 = n18554 | n18555;
  assign n34700 = n18558 | n18559;
  assign n34701 = n18566 | ~n18567;
  assign n34702 = n18575 | n18576;
  assign n34703 = n18583 | ~n18584;
  assign n34704 = n18593 | n18594;
  assign n34705 = n18597 | n18598;
  assign n34706 = n18606 | n18607;
  assign n34707 = n18614 | ~n18615;
  assign n34708 = n18620 | n18621;
  assign n34709 = n18624 | n18625;
  assign n34710 = n18632 | ~n18633;
  assign n34711 = n18641 | n18642;
  assign n34712 = n18649 | ~n18650;
  assign n34713 = n18658 | n18659;
  assign n34714 = n18663 | n18664;
  assign n34715 = n18670 | n18671;
  assign n34716 = n18682 | n18683;
  assign n34717 = n18690 | n18691;
  assign n34718 = n18698 | n18699;
  assign n34719 = n18706 | n18707;
  assign n34720 = n18714 | n18715;
  assign n34721 = n18722 | n18723;
  assign n34722 = n18730 | n18731;
  assign n34723 = n18738 | n18739;
  assign n34724 = n18746 | n18747;
  assign n34725 = n18754 | n18755;
  assign n34726 = n18762 | n18763;
  assign n34727 = n18770 | n18771;
  assign n34728 = n18778 | n18779;
  assign n34729 = n18786 | n18787;
  assign n34730 = n18794 | n18795;
  assign n34731 = n18802 | n18803;
  assign n34732 = n18810 | n18811;
  assign n34733 = n18818 | n18819;
  assign n34734 = n18826 | n18827;
  assign n34735 = n18830 | n18831;
  assign n34736 = n18838 | n18839;
  assign n34737 = n18848 | n18849;
  assign n34738 = n18855 | n18856;
  assign n34739 = n18863 | n18864;
  assign n34740 = n18873 | n18874;
  assign n34741 = n18881 | n18882;
  assign n34742 = n18893 | n18894;
  assign n34743 = n18896 | ~n18897;
  assign n34744 = n18903 | n18904;
  assign n34745 = n18917 | ~n18918;
  assign n34746 = n18924 | n18925;
  assign n34747 = n18935 | n18936;
  assign n34748 = n18939 | ~n18940;
  assign n34749 = n18946 | n18947;
  assign n34750 = n18957 | n18958;
  assign n34751 = n18961 | ~n18962;
  assign n34752 = n18968 | n18969;
  assign n34753 = n18976 | n18977;
  assign n34754 = n18979 | n18980;
  assign n34755 = n18985 | ~n18986;
  assign n34756 = n18992 | n18993;
  assign n34757 = n19003 | n19004;
  assign n34758 = n19011 | n19012;
  assign n34759 = n19019 | n19020;
  assign n34760 = n19022 | n19023;
  assign n34761 = n19028 | ~n19029;
  assign n34762 = n19035 | n19036;
  assign n34763 = n19047 | n19048;
  assign n34764 = n19050 | ~n19051;
  assign n34765 = n19057 | n19058;
  assign n34766 = n19065 | n19066;
  assign n34767 = n19068 | n19069;
  assign n34768 = n19074 | ~n19075;
  assign n34769 = n19081 | n19082;
  assign n34770 = n19092 | n19093;
  assign n34771 = n19100 | n19101;
  assign n34772 = n19108 | ~n19109;
  assign n34773 = n19115 | n19116;
  assign n34774 = n19126 | n19127;
  assign n34775 = n19134 | n19135;
  assign n34776 = n19142 | ~n19143;
  assign n34777 = n19149 | n19150;
  assign n34778 = n19160 | n19161;
  assign n34779 = n19173 | n19174;
  assign n34780 = n19177 | ~n19178;
  assign n34781 = n19183 | n19184;
  assign n34782 = n19192 | n19193;
  assign n34783 = n19200 | ~n19201;
  assign n34784 = n19210 | n19211;
  assign n34785 = n19214 | n19215;
  assign n34786 = n19223 | n19224;
  assign n34787 = n19231 | ~n19232;
  assign n34788 = n19241 | n19242;
  assign n34789 = n19245 | n19246;
  assign n34790 = n19255 | n19256;
  assign n34791 = n19268 | n19269;
  assign n34792 = n19272 | n19273;
  assign n34793 = n19281 | n19282;
  assign n34794 = n19289 | ~n19290;
  assign n34795 = n19299 | n19300;
  assign n34796 = n19303 | n19304;
  assign n34797 = n19313 | n19314;
  assign n34798 = n19326 | n19327;
  assign n34799 = n19330 | n19331;
  assign n34800 = n19339 | n19340;
  assign n34801 = n19347 | ~n19348;
  assign n34802 = n19357 | n19358;
  assign n34803 = n19361 | n19362;
  assign n34804 = n19371 | n19372;
  assign n34805 = n19383 | n19384;
  assign n34806 = n19388 | n19389;
  assign n34807 = n19395 | n19396;
  assign n34808 = n19404 | n19405;
  assign n34809 = n19412 | ~n19413;
  assign n34810 = n19421 | n19422;
  assign n34811 = n19428 | n19429;
  assign n34812 = n19434 | n19435;
  assign n34813 = n19447 | n19448;
  assign n34814 = n19454 | n19455;
  assign n34815 = n19460 | n19461;
  assign n34816 = n19470 | n19471;
  assign n34817 = n19478 | ~n19479;
  assign n34818 = n19484 | n19485;
  assign n34819 = n19492 | n19493;
  assign n34820 = n19495 | ~n19496;
  assign n34821 = n19504 | n19505;
  assign n34822 = n19512 | ~n19513;
  assign n34823 = n19518 | n19519;
  assign n34824 = n19528 | ~n19529;
  assign n34825 = n19537 | n19538;
  assign n34826 = n19545 | ~n19546;
  assign n34827 = n19551 | n19552;
  assign n34828 = n19558 | n19559;
  assign n34829 = n19562 | ~n19563;
  assign n34830 = n19571 | n19572;
  assign n34831 = n19579 | ~n19580;
  assign n34832 = n19585 | n19586;
  assign n34833 = n19592 | n19593;
  assign n34834 = n19596 | ~n19597;
  assign n34835 = n19605 | n19606;
  assign n34836 = n19613 | ~n19614;
  assign n34837 = n19619 | n19620;
  assign n34838 = n19623 | n19624;
  assign n34839 = n19626 | n19627;
  assign n34840 = n19632 | ~n19633;
  assign n34841 = n19641 | n19642;
  assign n34842 = n19649 | ~n19650;
  assign n34843 = n19655 | n19656;
  assign n34844 = n19662 | n19663;
  assign n34845 = n19672 | n19673;
  assign n34846 = n19680 | ~n19681;
  assign n34847 = n19686 | n19687;
  assign n34848 = n19690 | n19691;
  assign n34849 = n19693 | n19694;
  assign n34850 = n19699 | ~n19700;
  assign n34851 = n19708 | n19709;
  assign n34852 = n19716 | ~n19717;
  assign n34853 = n19722 | n19723;
  assign n34854 = n19730 | n19731;
  assign n34855 = n19733 | ~n19734;
  assign n34856 = n19742 | n19743;
  assign n34857 = n19750 | ~n19751;
  assign n34858 = n19756 | n19757;
  assign n34859 = n19760 | n19761;
  assign n34860 = n19763 | n19764;
  assign n34861 = n19769 | ~n19770;
  assign n34862 = n19778 | n19779;
  assign n34863 = n19786 | ~n19787;
  assign n34864 = n19796 | n19797;
  assign n34865 = n19800 | n19801;
  assign n34866 = n19809 | n19810;
  assign n34867 = n19817 | ~n19818;
  assign n34868 = n19823 | n19824;
  assign n34869 = n19827 | n19828;
  assign n34870 = n19835 | ~n19836;
  assign n34871 = n19844 | n19845;
  assign n34872 = n19852 | ~n19853;
  assign n34873 = n19862 | n19863;
  assign n34874 = n19866 | n19867;
  assign n34875 = n19875 | n19876;
  assign n34876 = n19883 | ~n19884;
  assign n34877 = n19889 | n19890;
  assign n34878 = n19893 | n19894;
  assign n34879 = n19901 | ~n19902;
  assign n34880 = n19910 | n19911;
  assign n34881 = n19918 | ~n19919;
  assign n34882 = n19928 | n19929;
  assign n34883 = n19932 | n19933;
  assign n34884 = n19941 | n19942;
  assign n34885 = n19949 | ~n19950;
  assign n34886 = n19955 | n19956;
  assign n34887 = n19959 | n19960;
  assign n34888 = n19967 | ~n19968;
  assign n34889 = n19982 | ~n19983;
  assign n34890 = n19992 | n19993;
  assign n34891 = n19996 | ~n19997;
  assign n34892 = n19999 | n20000;
  assign n34893 = n20014 | n20015;
  assign n34894 = n20018 | n20019;
  assign n34895 = n20027 | n20028;
  assign n34896 = n20035 | ~n20036;
  assign n34897 = n20045 | n20046;
  assign n34898 = n20049 | n20050;
  assign n34899 = n20058 | n20059;
  assign n34900 = n20066 | ~n20067;
  assign n34901 = n20072 | n20073;
  assign n34902 = n20076 | n20077;
  assign n34903 = n20084 | ~n20085;
  assign n34904 = n20093 | n20094;
  assign n34905 = n20101 | ~n20102;
  assign n34906 = n20111 | n20112;
  assign n34907 = n20115 | n20116;
  assign n34908 = n20124 | n20125;
  assign n34909 = n20132 | ~n20133;
  assign n34910 = n20138 | n20139;
  assign n34911 = n20142 | n20143;
  assign n34912 = n20150 | ~n20151;
  assign n34913 = n20159 | n20160;
  assign n34914 = n20167 | ~n20168;
  assign n34915 = n20177 | n20178;
  assign n34916 = n20181 | n20182;
  assign n34917 = n20190 | n20191;
  assign n34918 = n20198 | ~n20199;
  assign n34919 = n20204 | n20205;
  assign n34920 = n20212 | ~n20213;
  assign n34921 = n20216 | n20217;
  assign n34922 = n20223 | n20224;
  assign n34923 = n20235 | n20236;
  assign n34924 = n20243 | n20244;
  assign n34925 = n20251 | n20252;
  assign n34926 = n20259 | n20260;
  assign n34927 = n20267 | n20268;
  assign n34928 = n20275 | n20276;
  assign n34929 = n20283 | n20284;
  assign n34930 = n20291 | n20292;
  assign n34931 = n20299 | n20300;
  assign n34932 = n20307 | n20308;
  assign n34933 = n20315 | n20316;
  assign n34934 = n20323 | n20324;
  assign n34935 = n20331 | n20332;
  assign n34936 = n20339 | n20340;
  assign n34937 = n20347 | n20348;
  assign n34938 = n20355 | n20356;
  assign n34939 = n20363 | n20364;
  assign n34940 = n20371 | n20372;
  assign n34941 = n20379 | n20380;
  assign n34942 = n20387 | n20388;
  assign n34943 = n20395 | n20396;
  assign n34944 = n20399 | n20400;
  assign n34945 = n20407 | n20408;
  assign n34946 = n20417 | n20418;
  assign n34947 = n20424 | n20425;
  assign n34948 = n20432 | n20433;
  assign n34949 = n20442 | n20443;
  assign n34950 = n20450 | n20451;
  assign n34951 = n20462 | n20463;
  assign n34952 = n20465 | ~n20466;
  assign n34953 = n20472 | n20473;
  assign n34954 = n20486 | ~n20487;
  assign n34955 = n20493 | n20494;
  assign n34956 = n20504 | n20505;
  assign n34957 = n20508 | ~n20509;
  assign n34958 = n20515 | n20516;
  assign n34959 = n20526 | n20527;
  assign n34960 = n20530 | ~n20531;
  assign n34961 = n20537 | n20538;
  assign n34962 = n20545 | n20546;
  assign n34963 = n20548 | n20549;
  assign n34964 = n20554 | ~n20555;
  assign n34965 = n20561 | n20562;
  assign n34966 = n20572 | n20573;
  assign n34967 = n20580 | n20581;
  assign n34968 = n20588 | n20589;
  assign n34969 = n20591 | n20592;
  assign n34970 = n20597 | ~n20598;
  assign n34971 = n20604 | n20605;
  assign n34972 = n20616 | n20617;
  assign n34973 = n20619 | ~n20620;
  assign n34974 = n20626 | n20627;
  assign n34975 = n20634 | n20635;
  assign n34976 = n20637 | n20638;
  assign n34977 = n20643 | ~n20644;
  assign n34978 = n20650 | n20651;
  assign n34979 = n20661 | n20662;
  assign n34980 = n20669 | n20670;
  assign n34981 = n20677 | ~n20678;
  assign n34982 = n20684 | n20685;
  assign n34983 = n20695 | n20696;
  assign n34984 = n20703 | n20704;
  assign n34985 = n20711 | ~n20712;
  assign n34986 = n20718 | n20719;
  assign n34987 = n20729 | n20730;
  assign n34988 = n20737 | n20738;
  assign n34989 = n20745 | ~n20746;
  assign n34990 = n20752 | n20753;
  assign n34991 = n20763 | n20764;
  assign n34992 = n20773 | ~n20774;
  assign n34993 = n20789 | ~n20790;
  assign n34994 = n20795 | n20796;
  assign n34995 = n20804 | n20805;
  assign n34996 = n20812 | ~n20813;
  assign n34997 = n20822 | n20823;
  assign n34998 = n20826 | n20827;
  assign n34999 = n20835 | n20836;
  assign n35000 = n20843 | ~n20844;
  assign n35001 = n20853 | n20854;
  assign n35002 = n20857 | n20858;
  assign n35003 = n20867 | n20868;
  assign n35004 = n20880 | n20881;
  assign n35005 = n20884 | n20885;
  assign n35006 = n20893 | n20894;
  assign n35007 = n20901 | ~n20902;
  assign n35008 = n20911 | n20912;
  assign n35009 = n20915 | n20916;
  assign n35010 = n20925 | n20926;
  assign n35011 = n20938 | n20939;
  assign n35012 = n20942 | n20943;
  assign n35013 = n20951 | n20952;
  assign n35014 = n20959 | ~n20960;
  assign n35015 = n20968 | n20969;
  assign n35016 = n20973 | n20974;
  assign n35017 = n20980 | n20981;
  assign n35018 = n20989 | n20990;
  assign n35019 = n20997 | ~n20998;
  assign n35020 = n21006 | n21007;
  assign n35021 = n21013 | n21014;
  assign n35022 = n21019 | n21020;
  assign n35023 = n21032 | n21033;
  assign n35024 = n21039 | n21040;
  assign n35025 = n21045 | n21046;
  assign n35026 = n21055 | n21056;
  assign n35027 = n21063 | ~n21064;
  assign n35028 = n21069 | n21070;
  assign n35029 = n21077 | n21078;
  assign n35030 = n21080 | ~n21081;
  assign n35031 = n21089 | n21090;
  assign n35032 = n21097 | ~n21098;
  assign n35033 = n21103 | n21104;
  assign n35034 = n21113 | ~n21114;
  assign n35035 = n21122 | n21123;
  assign n35036 = n21130 | ~n21131;
  assign n35037 = n21136 | n21137;
  assign n35038 = n21143 | n21144;
  assign n35039 = n21147 | ~n21148;
  assign n35040 = n21156 | n21157;
  assign n35041 = n21164 | ~n21165;
  assign n35042 = n21170 | n21171;
  assign n35043 = n21177 | n21178;
  assign n35044 = n21181 | ~n21182;
  assign n35045 = n21190 | n21191;
  assign n35046 = n21198 | ~n21199;
  assign n35047 = n21204 | n21205;
  assign n35048 = n21208 | n21209;
  assign n35049 = n21211 | n21212;
  assign n35050 = n21217 | ~n21218;
  assign n35051 = n21226 | n21227;
  assign n35052 = n21234 | ~n21235;
  assign n35053 = n21240 | n21241;
  assign n35054 = n21247 | n21248;
  assign n35055 = n21257 | n21258;
  assign n35056 = n21265 | ~n21266;
  assign n35057 = n21271 | n21272;
  assign n35058 = n21275 | n21276;
  assign n35059 = n21278 | n21279;
  assign n35060 = n21284 | ~n21285;
  assign n35061 = n21293 | n21294;
  assign n35062 = n21301 | ~n21302;
  assign n35063 = n21307 | n21308;
  assign n35064 = n21315 | n21316;
  assign n35065 = n21318 | ~n21319;
  assign n35066 = n21327 | n21328;
  assign n35067 = n21335 | ~n21336;
  assign n35068 = n21341 | n21342;
  assign n35069 = n21345 | n21346;
  assign n35070 = n21348 | n21349;
  assign n35071 = n21354 | ~n21355;
  assign n35072 = n21363 | n21364;
  assign n35073 = n21371 | ~n21372;
  assign n35074 = n21381 | n21382;
  assign n35075 = n21385 | n21386;
  assign n35076 = n21394 | n21395;
  assign n35077 = n21402 | ~n21403;
  assign n35078 = n21408 | n21409;
  assign n35079 = n21412 | n21413;
  assign n35080 = n21420 | ~n21421;
  assign n35081 = n21429 | n21430;
  assign n35082 = n21437 | ~n21438;
  assign n35083 = n21447 | n21448;
  assign n35084 = n21451 | n21452;
  assign n35085 = n21460 | n21461;
  assign n35086 = n21468 | ~n21469;
  assign n35087 = n21474 | n21475;
  assign n35088 = n21478 | n21479;
  assign n35089 = n21486 | ~n21487;
  assign n35090 = n21495 | n21496;
  assign n35091 = n21503 | ~n21504;
  assign n35092 = n21513 | n21514;
  assign n35093 = n21517 | n21518;
  assign n35094 = n21526 | n21527;
  assign n35095 = n21534 | ~n21535;
  assign n35096 = n21540 | n21541;
  assign n35097 = n21544 | n21545;
  assign n35098 = n21552 | ~n21553;
  assign n35099 = n21561 | n21562;
  assign n35100 = n21569 | ~n21570;
  assign n35101 = n21579 | n21580;
  assign n35102 = n21583 | n21584;
  assign n35103 = n21592 | n21593;
  assign n35104 = n21600 | ~n21601;
  assign n35105 = n21606 | n21607;
  assign n35106 = n21610 | n21611;
  assign n35107 = n21618 | ~n21619;
  assign n35108 = n21633 | ~n21634;
  assign n35109 = n21639 | n21640;
  assign n35110 = n21646 | n21647;
  assign n35111 = n21662 | n21663;
  assign n35112 = n21666 | n21667;
  assign n35113 = n21675 | n21676;
  assign n35114 = n21683 | ~n21684;
  assign n35115 = n21693 | n21694;
  assign n35116 = n21697 | n21698;
  assign n35117 = n21706 | n21707;
  assign n35118 = n21714 | ~n21715;
  assign n35119 = n21720 | n21721;
  assign n35120 = n21724 | n21725;
  assign n35121 = n21732 | ~n21733;
  assign n35122 = n21741 | n21742;
  assign n35123 = n21749 | ~n21750;
  assign n35124 = n21759 | n21760;
  assign n35125 = n21763 | n21764;
  assign n35126 = n21772 | n21773;
  assign n35127 = n21780 | ~n21781;
  assign n35128 = n21786 | n21787;
  assign n35129 = n21790 | n21791;
  assign n35130 = n21798 | ~n21799;
  assign n35131 = n21807 | n21808;
  assign n35132 = n21815 | ~n21816;
  assign n35133 = n21824 | n21825;
  assign n35134 = n21829 | n21830;
  assign n35135 = n21836 | n21837;
  assign n35136 = n21848 | n21849;
  assign n35137 = n21856 | n21857;
  assign n35138 = n21864 | n21865;
  assign n35139 = n21872 | n21873;
  assign n35140 = n21880 | n21881;
  assign n35141 = n21888 | n21889;
  assign n35142 = n21896 | n21897;
  assign n35143 = n21904 | n21905;
  assign n35144 = n21912 | n21913;
  assign n35145 = n21920 | n21921;
  assign n35146 = n21928 | n21929;
  assign n35147 = n21936 | n21937;
  assign n35148 = n21944 | n21945;
  assign n35149 = n21952 | n21953;
  assign n35150 = n21960 | n21961;
  assign n35151 = n21968 | n21969;
  assign n35152 = n21976 | n21977;
  assign n35153 = n21984 | n21985;
  assign n35154 = n21992 | n21993;
  assign n35155 = n22000 | n22001;
  assign n35156 = n22008 | n22009;
  assign n35157 = n22016 | n22017;
  assign n35158 = n22024 | n22025;
  assign n35159 = n22032 | n22033;
  assign n35160 = n22040 | n22041;
  assign n35161 = n22044 | n22045;
  assign n35162 = n22052 | n22053;
  assign n35163 = n22062 | n22063;
  assign n35164 = n22069 | n22070;
  assign n35165 = n22077 | n22078;
  assign n35166 = n22087 | n22088;
  assign n35167 = n22095 | n22096;
  assign n35168 = n22107 | n22108;
  assign n35169 = n22110 | ~n22111;
  assign n35170 = n22117 | n22118;
  assign n35171 = n22131 | ~n22132;
  assign n35172 = n22138 | n22139;
  assign n35173 = n22149 | n22150;
  assign n35174 = n22153 | ~n22154;
  assign n35175 = n22160 | n22161;
  assign n35176 = n22171 | n22172;
  assign n35177 = n22175 | ~n22176;
  assign n35178 = n22182 | n22183;
  assign n35179 = n22190 | n22191;
  assign n35180 = n22193 | n22194;
  assign n35181 = n22199 | ~n22200;
  assign n35182 = n22206 | n22207;
  assign n35183 = n22217 | n22218;
  assign n35184 = n22225 | n22226;
  assign n35185 = n22233 | n22234;
  assign n35186 = n22236 | n22237;
  assign n35187 = n22242 | ~n22243;
  assign n35188 = n22249 | n22250;
  assign n35189 = n22261 | n22262;
  assign n35190 = n22264 | ~n22265;
  assign n35191 = n22271 | n22272;
  assign n35192 = n22279 | n22280;
  assign n35193 = n22282 | n22283;
  assign n35194 = n22288 | ~n22289;
  assign n35195 = n22295 | n22296;
  assign n35196 = n22306 | n22307;
  assign n35197 = n22314 | n22315;
  assign n35198 = n22322 | ~n22323;
  assign n35199 = n22329 | n22330;
  assign n35200 = n22340 | n22341;
  assign n35201 = n22348 | n22349;
  assign n35202 = n22356 | ~n22357;
  assign n35203 = n22363 | n22364;
  assign n35204 = n22374 | n22375;
  assign n35205 = n22382 | n22383;
  assign n35206 = n22390 | ~n22391;
  assign n35207 = n22397 | n22398;
  assign n35208 = n22408 | n22409;
  assign n35209 = n22416 | n22417;
  assign n35210 = n22424 | ~n22425;
  assign n35211 = n22431 | n22432;
  assign n35212 = n22442 | n22443;
  assign n35213 = n22456 | n22457;
  assign n35214 = n22459 | ~n22460;
  assign n35215 = n22465 | n22466;
  assign n35216 = n22474 | n22475;
  assign n35217 = n22482 | ~n22483;
  assign n35218 = n22492 | n22493;
  assign n35219 = n22496 | n22497;
  assign n35220 = n22505 | n22506;
  assign n35221 = n22513 | ~n22514;
  assign n35222 = n22523 | n22524;
  assign n35223 = n22527 | n22528;
  assign n35224 = n22537 | n22538;
  assign n35225 = n22550 | n22551;
  assign n35226 = n22554 | n22555;
  assign n35227 = n22563 | n22564;
  assign n35228 = n22571 | ~n22572;
  assign n35229 = n22581 | n22582;
  assign n35230 = n22585 | n22586;
  assign n35231 = n22595 | n22596;
  assign n35232 = n22607 | n22608;
  assign n35233 = n22612 | n22613;
  assign n35234 = n22619 | n22620;
  assign n35235 = n22628 | n22629;
  assign n35236 = n22636 | ~n22637;
  assign n35237 = n22645 | n22646;
  assign n35238 = n22652 | n22653;
  assign n35239 = n22658 | n22659;
  assign n35240 = n22671 | n22672;
  assign n35241 = n22678 | n22679;
  assign n35242 = n22684 | n22685;
  assign n35243 = n22694 | n22695;
  assign n35244 = n22702 | ~n22703;
  assign n35245 = n22708 | n22709;
  assign n35246 = n22716 | n22717;
  assign n35247 = n22719 | ~n22720;
  assign n35248 = n22728 | n22729;
  assign n35249 = n22736 | ~n22737;
  assign n35250 = n22742 | n22743;
  assign n35251 = n22752 | ~n22753;
  assign n35252 = n22761 | n22762;
  assign n35253 = n22769 | ~n22770;
  assign n35254 = n22775 | n22776;
  assign n35255 = n22782 | n22783;
  assign n35256 = n22786 | ~n22787;
  assign n35257 = n22795 | n22796;
  assign n35258 = n22803 | ~n22804;
  assign n35259 = n22809 | n22810;
  assign n35260 = n22816 | n22817;
  assign n35261 = n22820 | ~n22821;
  assign n35262 = n22829 | n22830;
  assign n35263 = n22837 | ~n22838;
  assign n35264 = n22843 | n22844;
  assign n35265 = n22847 | n22848;
  assign n35266 = n22850 | n22851;
  assign n35267 = n22856 | ~n22857;
  assign n35268 = n22865 | n22866;
  assign n35269 = n22873 | ~n22874;
  assign n35270 = n22879 | n22880;
  assign n35271 = n22886 | n22887;
  assign n35272 = n22896 | n22897;
  assign n35273 = n22904 | ~n22905;
  assign n35274 = n22910 | n22911;
  assign n35275 = n22914 | n22915;
  assign n35276 = n22917 | n22918;
  assign n35277 = n22923 | ~n22924;
  assign n35278 = n22932 | n22933;
  assign n35279 = n22940 | ~n22941;
  assign n35280 = n22946 | n22947;
  assign n35281 = n22954 | n22955;
  assign n35282 = n22957 | ~n22958;
  assign n35283 = n22966 | n22967;
  assign n35284 = n22974 | ~n22975;
  assign n35285 = n22980 | n22981;
  assign n35286 = n22984 | n22985;
  assign n35287 = n22987 | n22988;
  assign n35288 = n22993 | ~n22994;
  assign n35289 = n23002 | n23003;
  assign n35290 = n23010 | ~n23011;
  assign n35291 = n23020 | n23021;
  assign n35292 = n23024 | n23025;
  assign n35293 = n23033 | n23034;
  assign n35294 = n23041 | ~n23042;
  assign n35295 = n23047 | n23048;
  assign n35296 = n23051 | n23052;
  assign n35297 = n23059 | ~n23060;
  assign n35298 = n23068 | n23069;
  assign n35299 = n23076 | ~n23077;
  assign n35300 = n23086 | n23087;
  assign n35301 = n23090 | n23091;
  assign n35302 = n23099 | n23100;
  assign n35303 = n23107 | ~n23108;
  assign n35304 = n23113 | n23114;
  assign n35305 = n23117 | n23118;
  assign n35306 = n23125 | ~n23126;
  assign n35307 = n23134 | n23135;
  assign n35308 = n23142 | ~n23143;
  assign n35309 = n23152 | n23153;
  assign n35310 = n23156 | n23157;
  assign n35311 = n23165 | n23166;
  assign n35312 = n23173 | ~n23174;
  assign n35313 = n23179 | n23180;
  assign n35314 = n23183 | n23184;
  assign n35315 = n23191 | ~n23192;
  assign n35316 = n23200 | n23201;
  assign n35317 = n23208 | ~n23209;
  assign n35318 = n23218 | n23219;
  assign n35319 = n23222 | n23223;
  assign n35320 = n23231 | n23232;
  assign n35321 = n23239 | ~n23240;
  assign n35322 = n23245 | n23246;
  assign n35323 = n23249 | n23250;
  assign n35324 = n23257 | ~n23258;
  assign n35325 = n23266 | n23267;
  assign n35326 = n23274 | ~n23275;
  assign n35327 = n23284 | n23285;
  assign n35328 = n23288 | n23289;
  assign n35329 = n23297 | n23298;
  assign n35330 = n23305 | ~n23306;
  assign n35331 = n23311 | n23312;
  assign n35332 = n23315 | n23316;
  assign n35333 = n23323 | ~n23324;
  assign n35334 = n23334 | n23335;
  assign n35335 = n23342 | n23343;
  assign n35336 = n23350 | n23351;
  assign n35337 = n23353 | ~n23354;
  assign n35338 = n23368 | n23369;
  assign n35339 = n23372 | n23373;
  assign n35340 = n23381 | n23382;
  assign n35341 = n23389 | ~n23390;
  assign n35342 = n23399 | n23400;
  assign n35343 = n23403 | n23404;
  assign n35344 = n23412 | n23413;
  assign n35345 = n23420 | ~n23421;
  assign n35346 = n23426 | n23427;
  assign n35347 = n23430 | n23431;
  assign n35348 = n23438 | ~n23439;
  assign n35349 = n23447 | n23448;
  assign n35350 = n23455 | ~n23456;
  assign n35351 = n23465 | n23466;
  assign n35352 = n23469 | n23470;
  assign n35353 = n23478 | n23479;
  assign n35354 = n23486 | ~n23487;
  assign n35355 = n23492 | n23493;
  assign n35356 = n23500 | ~n23501;
  assign n35357 = n23504 | n23505;
  assign n35358 = n23511 | n23512;
  assign n35359 = n23523 | n23524;
  assign n35360 = n23531 | n23532;
  assign n35361 = n23539 | n23540;
  assign n35362 = n23547 | n23548;
  assign n35363 = n23555 | n23556;
  assign n35364 = n23563 | n23564;
  assign n35365 = n23571 | n23572;
  assign n35366 = n23579 | n23580;
  assign n35367 = n23587 | n23588;
  assign n35368 = n23595 | n23596;
  assign n35369 = n23603 | n23604;
  assign n35370 = n23611 | n23612;
  assign n35371 = n23619 | n23620;
  assign n35372 = n23627 | n23628;
  assign n35373 = n23635 | n23636;
  assign n35374 = n23643 | n23644;
  assign n35375 = n23651 | n23652;
  assign n35376 = n23659 | n23660;
  assign n35377 = n23667 | n23668;
  assign n35378 = n23675 | n23676;
  assign n35379 = n23683 | n23684;
  assign n35380 = n23691 | n23692;
  assign n35381 = n23699 | n23700;
  assign n35382 = n23707 | n23708;
  assign n35383 = n23715 | n23716;
  assign n35384 = n23723 | n23724;
  assign n35385 = n23731 | n23732;
  assign n35386 = n23739 | n23740;
  assign n35387 = n23743 | n23744;
  assign n35388 = n23751 | n23752;
  assign n35389 = n23761 | n23762;
  assign n35390 = n23768 | n23769;
  assign n35391 = n23776 | n23777;
  assign n35392 = n23786 | n23787;
  assign n35393 = n23794 | n23795;
  assign n35394 = n23806 | n23807;
  assign n35395 = n23809 | ~n23810;
  assign n35396 = n23816 | n23817;
  assign n35397 = n23830 | ~n23831;
  assign n35398 = n23837 | n23838;
  assign n35399 = n23848 | n23849;
  assign n35400 = n23852 | ~n23853;
  assign n35401 = n23859 | n23860;
  assign n35402 = n23870 | n23871;
  assign n35403 = n23874 | ~n23875;
  assign n35404 = n23881 | n23882;
  assign n35405 = n23889 | n23890;
  assign n35406 = n23892 | n23893;
  assign n35407 = n23898 | ~n23899;
  assign n35408 = n23905 | n23906;
  assign n35409 = n23916 | n23917;
  assign n35410 = n23924 | n23925;
  assign n35411 = n23932 | n23933;
  assign n35412 = n23935 | n23936;
  assign n35413 = n23941 | ~n23942;
  assign n35414 = n23948 | n23949;
  assign n35415 = n23960 | n23961;
  assign n35416 = n23963 | ~n23964;
  assign n35417 = n23970 | n23971;
  assign n35418 = n23978 | n23979;
  assign n35419 = n23981 | n23982;
  assign n35420 = n23987 | ~n23988;
  assign n35421 = n23994 | n23995;
  assign n35422 = n24005 | n24006;
  assign n35423 = n24013 | n24014;
  assign n35424 = n24021 | ~n24022;
  assign n35425 = n24028 | n24029;
  assign n35426 = n24039 | n24040;
  assign n35427 = n24047 | n24048;
  assign n35428 = n24055 | ~n24056;
  assign n35429 = n24062 | n24063;
  assign n35430 = n24073 | n24074;
  assign n35431 = n24081 | n24082;
  assign n35432 = n24089 | ~n24090;
  assign n35433 = n24096 | n24097;
  assign n35434 = n24107 | n24108;
  assign n35435 = n24115 | n24116;
  assign n35436 = n24123 | ~n24124;
  assign n35437 = n24130 | n24131;
  assign n35438 = n24141 | n24142;
  assign n35439 = n24149 | n24150;
  assign n35440 = n24157 | ~n24158;
  assign n35441 = n24164 | n24165;
  assign n35442 = n24175 | n24176;
  assign n35443 = n24188 | n24189;
  assign n35444 = n24192 | ~n24193;
  assign n35445 = n24198 | n24199;
  assign n35446 = n24207 | n24208;
  assign n35447 = n24215 | ~n24216;
  assign n35448 = n24225 | n24226;
  assign n35449 = n24229 | n24230;
  assign n35450 = n24238 | n24239;
  assign n35451 = n24246 | ~n24247;
  assign n35452 = n24256 | n24257;
  assign n35453 = n24260 | n24261;
  assign n35454 = n24270 | n24271;
  assign n35455 = n24283 | n24284;
  assign n35456 = n24287 | n24288;
  assign n35457 = n24296 | n24297;
  assign n35458 = n24304 | ~n24305;
  assign n35459 = n24313 | n24314;
  assign n35460 = n24318 | n24319;
  assign n35461 = n24325 | n24326;
  assign n35462 = n24334 | n24335;
  assign n35463 = n24342 | ~n24343;
  assign n35464 = n24351 | n24352;
  assign n35465 = n24358 | n24359;
  assign n35466 = n24364 | n24365;
  assign n35467 = n24377 | n24378;
  assign n35468 = n24384 | n24385;
  assign n35469 = n24390 | n24391;
  assign n35470 = n24400 | n24401;
  assign n35471 = n24408 | ~n24409;
  assign n35472 = n24414 | n24415;
  assign n35473 = n24422 | n24423;
  assign n35474 = n24425 | ~n24426;
  assign n35475 = n24434 | n24435;
  assign n35476 = n24442 | ~n24443;
  assign n35477 = n24448 | n24449;
  assign n35478 = n24458 | ~n24459;
  assign n35479 = n24467 | n24468;
  assign n35480 = n24475 | ~n24476;
  assign n35481 = n24481 | n24482;
  assign n35482 = n24488 | n24489;
  assign n35483 = n24492 | ~n24493;
  assign n35484 = n24501 | n24502;
  assign n35485 = n24509 | ~n24510;
  assign n35486 = n24515 | n24516;
  assign n35487 = n24522 | n24523;
  assign n35488 = n24526 | ~n24527;
  assign n35489 = n24535 | n24536;
  assign n35490 = n24543 | ~n24544;
  assign n35491 = n24549 | n24550;
  assign n35492 = n24553 | n24554;
  assign n35493 = n24556 | n24557;
  assign n35494 = n24562 | ~n24563;
  assign n35495 = n24571 | n24572;
  assign n35496 = n24579 | ~n24580;
  assign n35497 = n24585 | n24586;
  assign n35498 = n24592 | n24593;
  assign n35499 = n24602 | n24603;
  assign n35500 = n24610 | ~n24611;
  assign n35501 = n24616 | n24617;
  assign n35502 = n24620 | n24621;
  assign n35503 = n24623 | n24624;
  assign n35504 = n24629 | ~n24630;
  assign n35505 = n24638 | n24639;
  assign n35506 = n24646 | ~n24647;
  assign n35507 = n24652 | n24653;
  assign n35508 = n24660 | n24661;
  assign n35509 = n24663 | ~n24664;
  assign n35510 = n24672 | n24673;
  assign n35511 = n24680 | ~n24681;
  assign n35512 = n24686 | n24687;
  assign n35513 = n24690 | n24691;
  assign n35514 = n24693 | n24694;
  assign n35515 = n24699 | ~n24700;
  assign n35516 = n24708 | n24709;
  assign n35517 = n24716 | ~n24717;
  assign n35518 = n24726 | n24727;
  assign n35519 = n24730 | n24731;
  assign n35520 = n24739 | n24740;
  assign n35521 = n24747 | ~n24748;
  assign n35522 = n24753 | n24754;
  assign n35523 = n24757 | n24758;
  assign n35524 = n24765 | ~n24766;
  assign n35525 = n24774 | n24775;
  assign n35526 = n24782 | ~n24783;
  assign n35527 = n24792 | n24793;
  assign n35528 = n24796 | n24797;
  assign n35529 = n24805 | n24806;
  assign n35530 = n24813 | ~n24814;
  assign n35531 = n24819 | n24820;
  assign n35532 = n24823 | n24824;
  assign n35533 = n24831 | ~n24832;
  assign n35534 = n24840 | n24841;
  assign n35535 = n24848 | ~n24849;
  assign n35536 = n24858 | n24859;
  assign n35537 = n24862 | n24863;
  assign n35538 = n24871 | n24872;
  assign n35539 = n24879 | ~n24880;
  assign n35540 = n24885 | n24886;
  assign n35541 = n24889 | n24890;
  assign n35542 = n24897 | ~n24898;
  assign n35543 = n24906 | n24907;
  assign n35544 = n24914 | ~n24915;
  assign n35545 = n24924 | n24925;
  assign n35546 = n24928 | n24929;
  assign n35547 = n24937 | n24938;
  assign n35548 = n24945 | ~n24946;
  assign n35549 = n24951 | n24952;
  assign n35550 = n24955 | n24956;
  assign n35551 = n24963 | ~n24964;
  assign n35552 = n24972 | n24973;
  assign n35553 = n24980 | ~n24981;
  assign n35554 = n24990 | n24991;
  assign n35555 = n24994 | n24995;
  assign n35556 = n25003 | n25004;
  assign n35557 = n25011 | ~n25012;
  assign n35558 = n25017 | n25018;
  assign n35559 = n25021 | n25022;
  assign n35560 = n25029 | ~n25030;
  assign n35561 = n25038 | n25039;
  assign n35562 = n25046 | ~n25047;
  assign n35563 = n25056 | n25057;
  assign n35564 = n25060 | n25061;
  assign n35565 = n25069 | n25070;
  assign n35566 = n25077 | ~n25078;
  assign n35567 = n25083 | n25084;
  assign n35568 = n25087 | n25088;
  assign n35569 = n25095 | ~n25096;
  assign n35570 = n25110 | ~n25111;
  assign n35571 = n25120 | n25121;
  assign n35572 = n25124 | ~n25125;
  assign n35573 = n25127 | n25128;
  assign n35574 = n25142 | n25143;
  assign n35575 = n25146 | n25147;
  assign n35576 = n25155 | n25156;
  assign n35577 = n25163 | ~n25164;
  assign n35578 = n25173 | n25174;
  assign n35579 = n25177 | n25178;
  assign n35580 = n25186 | n25187;
  assign n35581 = n25194 | ~n25195;
  assign n35582 = n25200 | n25201;
  assign n35583 = n25204 | n25205;
  assign n35584 = n25212 | ~n25213;
  assign n35585 = n25221 | n25222;
  assign n35586 = n25229 | ~n25230;
  assign n35587 = n25238 | n25239;
  assign n35588 = n25243 | n25244;
  assign n35589 = n25250 | n25251;
  assign n35590 = n25262 | n25263;
  assign n35591 = n25270 | n25271;
  assign n35592 = n25278 | n25279;
  assign n35593 = n25286 | n25287;
  assign n35594 = n25294 | n25295;
  assign n35595 = n25302 | n25303;
  assign n35596 = n25310 | n25311;
  assign n35597 = n25318 | n25319;
  assign n35598 = n25326 | n25327;
  assign n35599 = n25334 | n25335;
  assign n35600 = n25342 | n25343;
  assign n35601 = n25350 | n25351;
  assign n35602 = n25358 | n25359;
  assign n35603 = n25366 | n25367;
  assign n35604 = n25374 | n25375;
  assign n35605 = n25382 | n25383;
  assign n35606 = n25390 | n25391;
  assign n35607 = n25398 | n25399;
  assign n35608 = n25406 | n25407;
  assign n35609 = n25414 | n25415;
  assign n35610 = n25422 | n25423;
  assign n35611 = n25430 | n25431;
  assign n35612 = n25438 | n25439;
  assign n35613 = n25446 | n25447;
  assign n35614 = n25454 | n25455;
  assign n35615 = n25462 | n25463;
  assign n35616 = n25470 | n25471;
  assign n35617 = n25478 | n25479;
  assign n35618 = n25486 | n25487;
  assign n35619 = n25494 | n25495;
  assign n35620 = n25498 | n25499;
  assign n35621 = n25506 | n25507;
  assign n35622 = n25516 | n25517;
  assign n35623 = n25523 | n25524;
  assign n35624 = n25531 | n25532;
  assign n35625 = n25541 | n25542;
  assign n35626 = n25549 | n25550;
  assign n35627 = n25561 | n25562;
  assign n35628 = n25564 | ~n25565;
  assign n35629 = n25571 | n25572;
  assign n35630 = n25585 | ~n25586;
  assign n35631 = n25592 | n25593;
  assign n35632 = n25603 | n25604;
  assign n35633 = n25607 | ~n25608;
  assign n35634 = n25614 | n25615;
  assign n35635 = n25625 | n25626;
  assign n35636 = n25629 | ~n25630;
  assign n35637 = n25636 | n25637;
  assign n35638 = n25644 | n25645;
  assign n35639 = n25647 | n25648;
  assign n35640 = n25653 | ~n25654;
  assign n35641 = n25660 | n25661;
  assign n35642 = n25671 | n25672;
  assign n35643 = n25679 | n25680;
  assign n35644 = n25687 | n25688;
  assign n35645 = n25690 | n25691;
  assign n35646 = n25696 | ~n25697;
  assign n35647 = n25703 | n25704;
  assign n35648 = n25715 | n25716;
  assign n35649 = n25718 | ~n25719;
  assign n35650 = n25725 | n25726;
  assign n35651 = n25733 | n25734;
  assign n35652 = n25736 | n25737;
  assign n35653 = n25742 | ~n25743;
  assign n35654 = n25749 | n25750;
  assign n35655 = n25760 | n25761;
  assign n35656 = n25768 | n25769;
  assign n35657 = n25776 | ~n25777;
  assign n35658 = n25783 | n25784;
  assign n35659 = n25794 | n25795;
  assign n35660 = n25802 | n25803;
  assign n35661 = n25810 | ~n25811;
  assign n35662 = n25817 | n25818;
  assign n35663 = n25828 | n25829;
  assign n35664 = n25836 | n25837;
  assign n35665 = n25844 | ~n25845;
  assign n35666 = n25851 | n25852;
  assign n35667 = n25862 | n25863;
  assign n35668 = n25870 | n25871;
  assign n35669 = n25878 | ~n25879;
  assign n35670 = n25885 | n25886;
  assign n35671 = n25896 | n25897;
  assign n35672 = n25904 | n25905;
  assign n35673 = n25912 | ~n25913;
  assign n35674 = n25919 | n25920;
  assign n35675 = n25930 | n25931;
  assign n35676 = n25938 | n25939;
  assign n35677 = n25946 | ~n25947;
  assign n35678 = n25953 | n25954;
  assign n35679 = n25964 | n25965;
  assign n35680 = n25974 | ~n25975;
  assign n35681 = n25990 | ~n25991;
  assign n35682 = n25996 | n25997;
  assign n35683 = n26005 | n26006;
  assign n35684 = n26013 | ~n26014;
  assign n35685 = n26023 | n26024;
  assign n35686 = n26027 | n26028;
  assign n35687 = n26036 | n26037;
  assign n35688 = n26044 | ~n26045;
  assign n35689 = n26054 | n26055;
  assign n35690 = n26058 | n26059;
  assign n35691 = n26068 | n26069;
  assign n35692 = n26080 | n26081;
  assign n35693 = n26085 | n26086;
  assign n35694 = n26092 | n26093;
  assign n35695 = n26101 | n26102;
  assign n35696 = n26109 | ~n26110;
  assign n35697 = n26118 | n26119;
  assign n35698 = n26125 | n26126;
  assign n35699 = n26131 | n26132;
  assign n35700 = n26144 | n26145;
  assign n35701 = n26151 | n26152;
  assign n35702 = n26157 | n26158;
  assign n35703 = n26167 | n26168;
  assign n35704 = n26175 | ~n26176;
  assign n35705 = n26181 | n26182;
  assign n35706 = n26189 | n26190;
  assign n35707 = n26192 | ~n26193;
  assign n35708 = n26201 | n26202;
  assign n35709 = n26209 | ~n26210;
  assign n35710 = n26215 | n26216;
  assign n35711 = n26225 | ~n26226;
  assign n35712 = n26234 | n26235;
  assign n35713 = n26242 | ~n26243;
  assign n35714 = n26248 | n26249;
  assign n35715 = n26255 | n26256;
  assign n35716 = n26259 | ~n26260;
  assign n35717 = n26268 | n26269;
  assign n35718 = n26276 | ~n26277;
  assign n35719 = n26282 | n26283;
  assign n35720 = n26289 | n26290;
  assign n35721 = n26293 | ~n26294;
  assign n35722 = n26302 | n26303;
  assign n35723 = n26310 | ~n26311;
  assign n35724 = n26316 | n26317;
  assign n35725 = n26320 | n26321;
  assign n35726 = n26323 | n26324;
  assign n35727 = n26329 | ~n26330;
  assign n35728 = n26338 | n26339;
  assign n35729 = n26346 | ~n26347;
  assign n35730 = n26352 | n26353;
  assign n35731 = n26359 | n26360;
  assign n35732 = n26369 | n26370;
  assign n35733 = n26377 | ~n26378;
  assign n35734 = n26383 | n26384;
  assign n35735 = n26387 | n26388;
  assign n35736 = n26390 | n26391;
  assign n35737 = n26396 | ~n26397;
  assign n35738 = n26405 | n26406;
  assign n35739 = n26413 | ~n26414;
  assign n35740 = n26419 | n26420;
  assign n35741 = n26427 | n26428;
  assign n35742 = n26430 | ~n26431;
  assign n35743 = n26439 | n26440;
  assign n35744 = n26447 | ~n26448;
  assign n35745 = n26453 | n26454;
  assign n35746 = n26457 | n26458;
  assign n35747 = n26460 | n26461;
  assign n35748 = n26466 | ~n26467;
  assign n35749 = n26475 | n26476;
  assign n35750 = n26483 | ~n26484;
  assign n35751 = n26493 | n26494;
  assign n35752 = n26497 | n26498;
  assign n35753 = n26506 | n26507;
  assign n35754 = n26514 | ~n26515;
  assign n35755 = n26520 | n26521;
  assign n35756 = n26524 | n26525;
  assign n35757 = n26532 | ~n26533;
  assign n35758 = n26541 | n26542;
  assign n35759 = n26549 | ~n26550;
  assign n35760 = n26559 | n26560;
  assign n35761 = n26563 | n26564;
  assign n35762 = n26572 | n26573;
  assign n35763 = n26580 | ~n26581;
  assign n35764 = n26586 | n26587;
  assign n35765 = n26590 | n26591;
  assign n35766 = n26598 | ~n26599;
  assign n35767 = n26607 | n26608;
  assign n35768 = n26615 | ~n26616;
  assign n35769 = n26625 | n26626;
  assign n35770 = n26629 | n26630;
  assign n35771 = n26638 | n26639;
  assign n35772 = n26646 | ~n26647;
  assign n35773 = n26652 | n26653;
  assign n35774 = n26656 | n26657;
  assign n35775 = n26664 | ~n26665;
  assign n35776 = n26673 | n26674;
  assign n35777 = n26681 | ~n26682;
  assign n35778 = n26691 | n26692;
  assign n35779 = n26695 | n26696;
  assign n35780 = n26704 | n26705;
  assign n35781 = n26712 | ~n26713;
  assign n35782 = n26718 | n26719;
  assign n35783 = n26722 | n26723;
  assign n35784 = n26730 | ~n26731;
  assign n35785 = n26739 | n26740;
  assign n35786 = n26747 | ~n26748;
  assign n35787 = n26757 | n26758;
  assign n35788 = n26761 | n26762;
  assign n35789 = n26770 | n26771;
  assign n35790 = n26778 | ~n26779;
  assign n35791 = n26784 | n26785;
  assign n35792 = n26788 | n26789;
  assign n35793 = n26796 | ~n26797;
  assign n35794 = n26805 | n26806;
  assign n35795 = n26813 | ~n26814;
  assign n35796 = n26823 | n26824;
  assign n35797 = n26827 | n26828;
  assign n35798 = n26836 | n26837;
  assign n35799 = n26844 | ~n26845;
  assign n35800 = n26850 | n26851;
  assign n35801 = n26854 | n26855;
  assign n35802 = n26862 | ~n26863;
  assign n35803 = n26871 | n26872;
  assign n35804 = n26879 | ~n26880;
  assign n35805 = n26889 | n26890;
  assign n35806 = n26893 | n26894;
  assign n35807 = n26902 | n26903;
  assign n35808 = n26910 | ~n26911;
  assign n35809 = n26916 | n26917;
  assign n35810 = n26920 | n26921;
  assign n35811 = n26928 | ~n26929;
  assign n35812 = n26943 | ~n26944;
  assign n35813 = n26949 | n26950;
  assign n35814 = n26956 | n26957;
  assign n35815 = n26972 | n26973;
  assign n35816 = n26976 | n26977;
  assign n35817 = n26985 | n26986;
  assign n35818 = n26993 | ~n26994;
  assign n35819 = n27003 | n27004;
  assign n35820 = n27007 | n27008;
  assign n35821 = n27016 | n27017;
  assign n35822 = n27024 | ~n27025;
  assign n35823 = n27030 | n27031;
  assign n35824 = n27038 | ~n27039;
  assign n35825 = n27042 | n27043;
  assign n35826 = n27049 | n27050;
  assign n35827 = n27061 | n27062;
  assign n35828 = n27069 | n27070;
  assign n35829 = n27077 | n27078;
  assign n35830 = n27085 | n27086;
  assign n35831 = n27093 | n27094;
  assign n35832 = n27101 | n27102;
  assign n35833 = n27109 | n27110;
  assign n35834 = n27117 | n27118;
  assign n35835 = n27125 | n27126;
  assign n35836 = n27133 | n27134;
  assign n35837 = n27141 | n27142;
  assign n35838 = n27149 | n27150;
  assign n35839 = n27157 | n27158;
  assign n35840 = n27165 | n27166;
  assign n35841 = n27173 | n27174;
  assign n35842 = n27181 | n27182;
  assign n35843 = n27189 | n27190;
  assign n35844 = n27197 | n27198;
  assign n35845 = n27205 | n27206;
  assign n35846 = n27213 | n27214;
  assign n35847 = n27221 | n27222;
  assign n35848 = n27229 | n27230;
  assign n35849 = n27237 | n27238;
  assign n35850 = n27245 | n27246;
  assign n35851 = n27253 | n27254;
  assign n35852 = n27261 | n27262;
  assign n35853 = n27269 | n27270;
  assign n35854 = n27277 | n27278;
  assign n35855 = n27285 | n27286;
  assign n35856 = n27293 | n27294;
  assign n35857 = n27301 | n27302;
  assign n35858 = n27309 | n27310;
  assign n35859 = n27317 | n27318;
  assign n35860 = n27325 | n27326;
  assign n35861 = n27329 | n27330;
  assign n35862 = n27333 | n27334;
  assign n35863 = n27338 | n27339;
  assign n35864 = n27348 | n27349;
  assign n35865 = n27356 | ~n27357;
  assign n35866 = n27358 | n27359;
  assign n35867 = n27366 | n27367;
  assign n35868 = n27376 | n27377;
  assign n35869 = n27384 | n27385;
  assign n35870 = n27396 | n27397;
  assign n35871 = n27399 | ~n27400;
  assign n35872 = n27406 | n27407;
  assign n35873 = n27420 | ~n27421;
  assign n35874 = n27427 | n27428;
  assign n35875 = n27438 | n27439;
  assign n35876 = n27442 | ~n27443;
  assign n35877 = n27449 | n27450;
  assign n35878 = n27460 | n27461;
  assign n35879 = n27464 | ~n27465;
  assign n35880 = n27471 | n27472;
  assign n35881 = n27479 | n27480;
  assign n35882 = n27482 | n27483;
  assign n35883 = n27488 | ~n27489;
  assign n35884 = n27495 | n27496;
  assign n35885 = n27506 | n27507;
  assign n35886 = n27514 | n27515;
  assign n35887 = n27522 | n27523;
  assign n35888 = n27525 | n27526;
  assign n35889 = n27531 | ~n27532;
  assign n35890 = n27538 | n27539;
  assign n35891 = n27550 | n27551;
  assign n35892 = n27553 | ~n27554;
  assign n35893 = n27560 | n27561;
  assign n35894 = n27568 | n27569;
  assign n35895 = n27571 | n27572;
  assign n35896 = n27577 | ~n27578;
  assign n35897 = n27584 | n27585;
  assign n35898 = n27595 | n27596;
  assign n35899 = n27603 | n27604;
  assign n35900 = n27611 | ~n27612;
  assign n35901 = n27618 | n27619;
  assign n35902 = n27629 | n27630;
  assign n35903 = n27637 | n27638;
  assign n35904 = n27645 | ~n27646;
  assign n35905 = n27652 | n27653;
  assign n35906 = n27663 | n27664;
  assign n35907 = n27671 | n27672;
  assign n35908 = n27679 | ~n27680;
  assign n35909 = n27686 | n27687;
  assign n35910 = n27697 | n27698;
  assign n35911 = n27705 | n27706;
  assign n35912 = n27713 | ~n27714;
  assign n35913 = n27720 | n27721;
  assign n35914 = n27731 | n27732;
  assign n35915 = n27739 | n27740;
  assign n35916 = n27747 | ~n27748;
  assign n35917 = n27754 | n27755;
  assign n35918 = n27765 | n27766;
  assign n35919 = n27773 | n27774;
  assign n35920 = n27781 | ~n27782;
  assign n35921 = n27788 | n27789;
  assign n35922 = n27799 | n27800;
  assign n35923 = n27807 | n27808;
  assign n35924 = n27815 | ~n27816;
  assign n35925 = n27822 | n27823;
  assign n35926 = n27833 | n27834;
  assign n35927 = n27847 | n27848;
  assign n35928 = n27850 | ~n27851;
  assign n35929 = n27856 | n27857;
  assign n35930 = n27865 | n27866;
  assign n35931 = n27873 | ~n27874;
  assign n35932 = n27883 | n27884;
  assign n35933 = n27887 | n27888;
  assign n35934 = n27896 | n27897;
  assign n35935 = n27904 | ~n27905;
  assign n35936 = n27913 | n27914;
  assign n35937 = n27918 | n27919;
  assign n35938 = n27925 | n27926;
  assign n35939 = n27934 | n27935;
  assign n35940 = n27942 | ~n27943;
  assign n35941 = n27949 | ~n27950;
  assign n35942 = n27954 | n27955;
  assign n35943 = n27960 | n27961;
  assign n35944 = n27969 | n27970;
  assign n35945 = n27974 | n27975;
  assign n35946 = n27981 | n27982;
  assign n35947 = n27987 | n27988;
  assign n35948 = n27997 | n27998;
  assign n35949 = n28005 | ~n28006;
  assign n35950 = n28011 | n28012;
  assign n35951 = n28019 | n28020;
  assign n35952 = n28022 | ~n28023;
  assign n35953 = n28031 | n28032;
  assign n35954 = n28039 | ~n28040;
  assign n35955 = n28045 | n28046;
  assign n35956 = n28055 | ~n28056;
  assign n35957 = n28064 | n28065;
  assign n35958 = n28072 | ~n28073;
  assign n35959 = n28078 | n28079;
  assign n35960 = n28085 | n28086;
  assign n35961 = n28089 | ~n28090;
  assign n35962 = n28098 | n28099;
  assign n35963 = n28106 | ~n28107;
  assign n35964 = n28112 | n28113;
  assign n35965 = n28119 | n28120;
  assign n35966 = n28123 | ~n28124;
  assign n35967 = n28132 | n28133;
  assign n35968 = n28140 | ~n28141;
  assign n35969 = n28146 | n28147;
  assign n35970 = n28150 | n28151;
  assign n35971 = n28153 | n28154;
  assign n35972 = n28159 | ~n28160;
  assign n35973 = n28168 | n28169;
  assign n35974 = n28176 | ~n28177;
  assign n35975 = n28182 | n28183;
  assign n35976 = n28189 | n28190;
  assign n35977 = n28199 | n28200;
  assign n35978 = n28207 | ~n28208;
  assign n35979 = n28213 | n28214;
  assign n35980 = n28217 | n28218;
  assign n35981 = n28220 | n28221;
  assign n35982 = n28226 | ~n28227;
  assign n35983 = n28235 | n28236;
  assign n35984 = n28243 | ~n28244;
  assign n35985 = n28249 | n28250;
  assign n35986 = n28257 | n28258;
  assign n35987 = n28260 | ~n28261;
  assign n35988 = n28269 | n28270;
  assign n35989 = n28277 | ~n28278;
  assign n35990 = n28283 | n28284;
  assign n35991 = n28287 | n28288;
  assign n35992 = n28290 | n28291;
  assign n35993 = n28296 | ~n28297;
  assign n35994 = n28305 | n28306;
  assign n35995 = n28313 | ~n28314;
  assign n35996 = n28323 | n28324;
  assign n35997 = n28327 | n28328;
  assign n35998 = n28336 | n28337;
  assign n35999 = n28344 | ~n28345;
  assign n36000 = n28350 | n28351;
  assign n36001 = n28354 | n28355;
  assign n36002 = n28362 | ~n28363;
  assign n36003 = n28371 | n28372;
  assign n36004 = n28379 | ~n28380;
  assign n36005 = n28389 | n28390;
  assign n36006 = n28393 | n28394;
  assign n36007 = n28402 | n28403;
  assign n36008 = n28410 | ~n28411;
  assign n36009 = n28416 | n28417;
  assign n36010 = n28420 | n28421;
  assign n36011 = n28428 | ~n28429;
  assign n36012 = n28437 | n28438;
  assign n36013 = n28445 | ~n28446;
  assign n36014 = n28455 | n28456;
  assign n36015 = n28459 | n28460;
  assign n36016 = n28468 | n28469;
  assign n36017 = n28476 | ~n28477;
  assign n36018 = n28482 | n28483;
  assign n36019 = n28486 | n28487;
  assign n36020 = n28494 | ~n28495;
  assign n36021 = n28503 | n28504;
  assign n36022 = n28511 | ~n28512;
  assign n36023 = n28521 | n28522;
  assign n36024 = n28525 | n28526;
  assign n36025 = n28534 | n28535;
  assign n36026 = n28542 | ~n28543;
  assign n36027 = n28548 | n28549;
  assign n36028 = n28552 | n28553;
  assign n36029 = n28560 | ~n28561;
  assign n36030 = n28569 | n28570;
  assign n36031 = n28577 | ~n28578;
  assign n36032 = n28587 | n28588;
  assign n36033 = n28591 | n28592;
  assign n36034 = n28600 | n28601;
  assign n36035 = n28608 | ~n28609;
  assign n36036 = n28614 | n28615;
  assign n36037 = n28618 | n28619;
  assign n36038 = n28626 | ~n28627;
  assign n36039 = n28635 | n28636;
  assign n36040 = n28643 | ~n28644;
  assign n36041 = n28653 | n28654;
  assign n36042 = n28657 | n28658;
  assign n36043 = n28666 | n28667;
  assign n36044 = n28674 | ~n28675;
  assign n36045 = n28680 | n28681;
  assign n36046 = n28684 | n28685;
  assign n36047 = n28692 | ~n28693;
  assign n36048 = n28701 | n28702;
  assign n36049 = n28709 | ~n28710;
  assign n36050 = n28719 | n28720;
  assign n36051 = n28723 | n28724;
  assign n36052 = n28732 | n28733;
  assign n36053 = n28740 | ~n28741;
  assign n36054 = n28746 | n28747;
  assign n36055 = n28750 | n28751;
  assign n36056 = n28758 | ~n28759;
  assign n36057 = n28767 | n28768;
  assign n36058 = n28775 | ~n28776;
  assign n36059 = n28785 | n28786;
  assign n36060 = n28789 | n28790;
  assign n36061 = n28798 | n28799;
  assign n36062 = n28806 | ~n28807;
  assign n36063 = n28812 | n28813;
  assign n36064 = n28816 | n28817;
  assign n36065 = n28824 | ~n28825;
  assign n36066 = n28835 | n28836;
  assign n36067 = n28843 | n28844;
  assign n36068 = n28851 | n28852;
  assign n36069 = n28854 | ~n28855;
  assign n36070 = n28869 | n28870;
  assign n36071 = n28873 | n28874;
  assign n36072 = n28882 | n28883;
  assign n36073 = n28890 | ~n28891;
  assign n36074 = n28899 | n28900;
  assign n36075 = n28904 | n28905;
  assign n36076 = n28911 | n28912;
  assign n36077 = n28923 | n28924;
  assign n36078 = n28931 | n28932;
  assign n36079 = n28939 | n28940;
  assign n36080 = n28947 | n28948;
  assign n36081 = n28955 | n28956;
  assign n36082 = n28963 | n28964;
  assign n36083 = n28971 | n28972;
  assign n36084 = n28979 | n28980;
  assign n36085 = n28987 | n28988;
  assign n36086 = n28995 | n28996;
  assign n36087 = n29003 | n29004;
  assign n36088 = n29011 | n29012;
  assign n36089 = n29019 | n29020;
  assign n36090 = n29027 | n29028;
  assign n36091 = n29035 | n29036;
  assign n36092 = n29043 | n29044;
  assign n36093 = n29051 | n29052;
  assign n36094 = n29059 | n29060;
  assign n36095 = n29067 | n29068;
  assign n36096 = n29075 | n29076;
  assign n36097 = n29083 | n29084;
  assign n36098 = n29091 | n29092;
  assign n36099 = n29099 | n29100;
  assign n36100 = n29107 | n29108;
  assign n36101 = n29115 | n29116;
  assign n36102 = n29123 | n29124;
  assign n36103 = n29131 | n29132;
  assign n36104 = n29139 | n29140;
  assign n36105 = n29147 | n29148;
  assign n36106 = n29155 | n29156;
  assign n36107 = n29163 | n29164;
  assign n36108 = n29171 | n29172;
  assign n36109 = n29179 | n29180;
  assign n36110 = n29187 | n29188;
  assign n36111 = n29195 | n29196;
  assign n36112 = n29203 | n29204;
  assign n36113 = n29211 | n29212;
  assign n36114 = n29215 | n29216;
  assign n36115 = n29219 | n29220;
  assign n36116 = n29224 | n29225;
  assign n36117 = n29235 | ~n29236;
  assign n36118 = n29237 | n29238;
  assign n36119 = n29245 | n29246;
  assign n36120 = n29255 | n29256;
  assign n36121 = n29263 | n29264;
  assign n36122 = n29275 | n29276;
  assign n36123 = n29278 | ~n29279;
  assign n36124 = n29285 | n29286;
  assign n36125 = n29299 | ~n29300;
  assign n36126 = n29306 | n29307;
  assign n36127 = n29317 | n29318;
  assign n36128 = n29321 | ~n29322;
  assign n36129 = n29328 | n29329;
  assign n36130 = n29339 | n29340;
  assign n36131 = n29343 | ~n29344;
  assign n36132 = n29350 | n29351;
  assign n36133 = n29358 | n29359;
  assign n36134 = n29361 | n29362;
  assign n36135 = n29367 | ~n29368;
  assign n36136 = n29374 | n29375;
  assign n36137 = n29385 | n29386;
  assign n36138 = n29393 | n29394;
  assign n36139 = n29401 | n29402;
  assign n36140 = n29404 | n29405;
  assign n36141 = n29410 | ~n29411;
  assign n36142 = n29417 | n29418;
  assign n36143 = n29429 | n29430;
  assign n36144 = n29432 | ~n29433;
  assign n36145 = n29439 | n29440;
  assign n36146 = n29447 | n29448;
  assign n36147 = n29450 | n29451;
  assign n36148 = n29456 | ~n29457;
  assign n36149 = n29463 | n29464;
  assign n36150 = n29474 | n29475;
  assign n36151 = n29482 | n29483;
  assign n36152 = n29490 | ~n29491;
  assign n36153 = n29497 | n29498;
  assign n36154 = n29508 | n29509;
  assign n36155 = n29516 | n29517;
  assign n36156 = n29524 | ~n29525;
  assign n36157 = n29531 | n29532;
  assign n36158 = n29542 | n29543;
  assign n36159 = n29550 | n29551;
  assign n36160 = n29558 | ~n29559;
  assign n36161 = n29565 | n29566;
  assign n36162 = n29576 | n29577;
  assign n36163 = n29584 | n29585;
  assign n36164 = n29592 | ~n29593;
  assign n36165 = n29599 | n29600;
  assign n36166 = n29610 | n29611;
  assign n36167 = n29618 | n29619;
  assign n36168 = n29626 | ~n29627;
  assign n36169 = n29633 | n29634;
  assign n36170 = n29644 | n29645;
  assign n36171 = n29652 | n29653;
  assign n36172 = n29660 | ~n29661;
  assign n36173 = n29667 | n29668;
  assign n36174 = n29678 | n29679;
  assign n36175 = n29686 | n29687;
  assign n36176 = n29694 | ~n29695;
  assign n36177 = n29701 | n29702;
  assign n36178 = n29712 | n29713;
  assign n36179 = n29720 | n29721;
  assign n36180 = n29728 | ~n29729;
  assign n36181 = n29735 | n29736;
  assign n36182 = n29746 | n29747;
  assign n36183 = n29759 | n29760;
  assign n36184 = n29763 | ~n29764;
  assign n36185 = n29769 | n29770;
  assign n36186 = n29778 | n29779;
  assign n36187 = n29786 | ~n29787;
  assign n36188 = n29795 | n29796;
  assign n36189 = n29800 | n29801;
  assign n36190 = n29807 | n29808;
  assign n36191 = n29816 | n29817;
  assign n36192 = n29824 | ~n29825;
  assign n36193 = n29831 | ~n29832;
  assign n36194 = n29836 | n29837;
  assign n36195 = n29842 | n29843;
  assign n36196 = n29851 | n29852;
  assign n36197 = n29856 | n29857;
  assign n36198 = n29863 | n29864;
  assign n36199 = n29869 | n29870;
  assign n36200 = n29879 | n29880;
  assign n36201 = n29887 | ~n29888;
  assign n36202 = n29893 | n29894;
  assign n36203 = n29901 | n29902;
  assign n36204 = n29904 | ~n29905;
  assign n36205 = n29913 | n29914;
  assign n36206 = n29921 | ~n29922;
  assign n36207 = n29927 | n29928;
  assign n36208 = n29937 | ~n29938;
  assign n36209 = n29946 | n29947;
  assign n36210 = n29954 | ~n29955;
  assign n36211 = n29960 | n29961;
  assign n36212 = n29967 | n29968;
  assign n36213 = n29971 | ~n29972;
  assign n36214 = n29980 | n29981;
  assign n36215 = n29988 | ~n29989;
  assign n36216 = n29994 | n29995;
  assign n36217 = n30001 | n30002;
  assign n36218 = n30005 | ~n30006;
  assign n36219 = n30014 | n30015;
  assign n36220 = n30022 | ~n30023;
  assign n36221 = n30028 | n30029;
  assign n36222 = n30032 | n30033;
  assign n36223 = n30035 | n30036;
  assign n36224 = n30041 | ~n30042;
  assign n36225 = n30050 | n30051;
  assign n36226 = n30058 | ~n30059;
  assign n36227 = n30064 | n30065;
  assign n36228 = n30071 | n30072;
  assign n36229 = n30081 | n30082;
  assign n36230 = n30089 | ~n30090;
  assign n36231 = n30095 | n30096;
  assign n36232 = n30099 | n30100;
  assign n36233 = n30102 | n30103;
  assign n36234 = n30108 | ~n30109;
  assign n36235 = n30117 | n30118;
  assign n36236 = n30125 | ~n30126;
  assign n36237 = n30131 | n30132;
  assign n36238 = n30139 | n30140;
  assign n36239 = n30142 | ~n30143;
  assign n36240 = n30151 | n30152;
  assign n36241 = n30159 | ~n30160;
  assign n36242 = n30165 | n30166;
  assign n36243 = n30169 | n30170;
  assign n36244 = n30172 | n30173;
  assign n36245 = n30178 | ~n30179;
  assign n36246 = n30187 | n30188;
  assign n36247 = n30195 | ~n30196;
  assign n36248 = n30205 | n30206;
  assign n36249 = n30209 | n30210;
  assign n36250 = n30218 | n30219;
  assign n36251 = n30226 | ~n30227;
  assign n36252 = n30232 | n30233;
  assign n36253 = n30236 | n30237;
  assign n36254 = n30244 | ~n30245;
  assign n36255 = n30253 | n30254;
  assign n36256 = n30261 | ~n30262;
  assign n36257 = n30271 | n30272;
  assign n36258 = n30275 | n30276;
  assign n36259 = n30284 | n30285;
  assign n36260 = n30292 | ~n30293;
  assign n36261 = n30298 | n30299;
  assign n36262 = n30302 | n30303;
  assign n36263 = n30310 | ~n30311;
  assign n36264 = n30319 | n30320;
  assign n36265 = n30327 | ~n30328;
  assign n36266 = n30337 | n30338;
  assign n36267 = n30341 | n30342;
  assign n36268 = n30350 | n30351;
  assign n36269 = n30358 | ~n30359;
  assign n36270 = n30364 | n30365;
  assign n36271 = n30368 | n30369;
  assign n36272 = n30376 | ~n30377;
  assign n36273 = n30385 | n30386;
  assign n36274 = n30393 | ~n30394;
  assign n36275 = n30403 | n30404;
  assign n36276 = n30407 | n30408;
  assign n36277 = n30416 | n30417;
  assign n36278 = n30424 | ~n30425;
  assign n36279 = n30430 | n30431;
  assign n36280 = n30434 | n30435;
  assign n36281 = n30442 | ~n30443;
  assign n36282 = n30451 | n30452;
  assign n36283 = n30459 | ~n30460;
  assign n36284 = n30469 | n30470;
  assign n36285 = n30473 | n30474;
  assign n36286 = n30482 | n30483;
  assign n36287 = n30490 | ~n30491;
  assign n36288 = n30496 | n30497;
  assign n36289 = n30500 | n30501;
  assign n36290 = n30508 | ~n30509;
  assign n36291 = n30517 | n30518;
  assign n36292 = n30525 | ~n30526;
  assign n36293 = n30535 | n30536;
  assign n36294 = n30539 | n30540;
  assign n36295 = n30548 | n30549;
  assign n36296 = n30556 | ~n30557;
  assign n36297 = n30562 | n30563;
  assign n36298 = n30566 | n30567;
  assign n36299 = n30574 | ~n30575;
  assign n36300 = n30583 | n30584;
  assign n36301 = n30591 | ~n30592;
  assign n36302 = n30601 | n30602;
  assign n36303 = n30605 | n30606;
  assign n36304 = n30614 | n30615;
  assign n36305 = n30622 | ~n30623;
  assign n36306 = n30628 | n30629;
  assign n36307 = n30632 | n30633;
  assign n36308 = n30640 | ~n30641;
  assign n36309 = n30649 | n30650;
  assign n36310 = n30657 | ~n30658;
  assign n36311 = n30667 | n30668;
  assign n36312 = n30671 | n30672;
  assign n36313 = n30680 | n30681;
  assign n36314 = n30688 | ~n30689;
  assign n36315 = n30694 | n30695;
  assign n36316 = n30698 | n30699;
  assign n36317 = n30706 | ~n30707;
  assign n36318 = n30715 | n30716;
  assign n36319 = n30723 | ~n30724;
  assign n36320 = n30733 | n30734;
  assign n36321 = n30737 | n30738;
  assign n36322 = n30746 | n30747;
  assign n36323 = n30754 | ~n30755;
  assign n36324 = n30760 | n30761;
  assign n36325 = n30764 | n30765;
  assign n36326 = n30772 | ~n30773;
  assign n36327 = n30787 | ~n30788;
  assign n36328 = n30797 | n30798;
  assign n36329 = n30801 | ~n30802;
  assign n36330 = n30804 | n30805;
  assign n36331 = n30818 | n30819;
  assign n36332 = n30823 | n30824;
  assign n36333 = n30830 | n30831;
  assign n36334 = n30842 | n30843;
  assign n36335 = n30854 | ~n30855;
  assign n36336 = n30866 | ~n30867;
  assign n36337 = n30874 | n30875;
  assign n36338 = n30880 | n30881;
  assign n36339 = n30888 | ~n30889;
  assign n36340 = n30896 | n30897;
  assign n36341 = n30902 | n30903;
  assign n36342 = n30910 | ~n30911;
  assign n36343 = n30918 | n30919;
  assign n36344 = n30924 | n30925;
  assign n36345 = n30932 | ~n30933;
  assign n36346 = n30940 | n30941;
  assign n36347 = n30946 | n30947;
  assign n36348 = n30954 | ~n30955;
  assign n36349 = n30962 | n30963;
  assign n36350 = n30968 | n30969;
  assign n36351 = n30976 | ~n30977;
  assign n36352 = n30984 | n30985;
  assign n36353 = n30990 | n30991;
  assign n36354 = n30998 | ~n30999;
  assign n36355 = n31006 | n31007;
  assign n36356 = n31012 | n31013;
  assign n36357 = n31020 | ~n31021;
  assign n36358 = n31028 | n31029;
  assign n36359 = n31034 | n31035;
  assign n36360 = n31042 | ~n31043;
  assign n36361 = n31050 | n31051;
  assign n36362 = n31056 | n31057;
  assign n36363 = n31059 | n31060;
  assign n36364 = n31065 | ~n31066;
  assign n36365 = n31075 | n31076;
  assign n36366 = n31077 | ~n31078;
  assign n36367 = n31082 | n31083;
  assign n36368 = n31085 | n31086;
  assign n36369 = n31091 | ~n31092;
  assign n36370 = n31099 | n31100;
  assign n36371 = n31105 | n31106;
  assign n36372 = n31108 | n31109;
  assign n36373 = n31114 | ~n31115;
  assign n36374 = n31122 | n31123;
  assign n36375 = n31126 | ~n31127;
  assign n36376 = n31134 | n31135;
  assign n36377 = n31138 | ~n31139;
  assign n36378 = n31149 | ~n31150;
  assign n36379 = n31158 | n31159;
  assign n36380 = n31161 | ~n31162;
  assign n36381 = n31170 | n31171;
  assign n36382 = n31178 | n31179;
  assign n36383 = n31183 | n31184;
  assign n36384 = n31190 | n31191;
  assign n36385 = ~n31197 | n31194 | ~n31196;
  assign n36386 = n31201 | n31202;
  assign n36387 = n31206 | n31207;
  assign n36388 = n31214 | n31215;
  assign n36389 = n31231 | n31232;
  assign n36390 = n31236 | n31237;
  assign n36391 = ~n31242 | n31240 | n31241;
  assign n36392 = n31249 | n31244 | n31248;
  assign n36393 = ~n31259 | n31253 | ~n31258;
  assign n36394 = n31266 | n31267;
  assign n36395 = n31279 | n31280;
  assign n36396 = n31285 | n31283 | n31284;
  assign n36397 = ~n31293 | n31287 | n31292;
  assign n36398 = n31300 | n31301;
  assign n36399 = n31313 | n31314;
  assign n36400 = n31319 | n31317 | n31318;
  assign n36401 = ~n31327 | n31321 | n31326;
  assign n36402 = n31334 | n31335;
  assign n36403 = n31347 | n31348;
  assign n36404 = n31353 | n31351 | n31352;
  assign n36405 = ~n31361 | n31355 | n31360;
  assign n36406 = n31368 | n31369;
  assign n36407 = n31381 | n31382;
  assign n36408 = n31387 | n31385 | n31386;
  assign n36409 = ~n31395 | n31389 | n31394;
  assign n36410 = n31402 | n31403;
  assign n36411 = n31415 | n31416;
  assign n36412 = n31421 | n31419 | n31420;
  assign n36413 = ~n31429 | n31423 | n31428;
  assign n36414 = n31436 | n31437;
  assign n36415 = n31449 | n31450;
  assign n36416 = n31455 | n31453 | n31454;
  assign n36417 = ~n31463 | n31457 | n31462;
  assign n36418 = n31470 | n31471;
  assign n36419 = n31483 | n31484;
  assign n36420 = n31489 | n31487 | n31488;
  assign n36421 = ~n31497 | n31491 | n31496;
  assign n36422 = n31504 | n31505;
  assign n36423 = n31517 | n31518;
  assign n36424 = n31523 | n31521 | n31522;
  assign n36425 = ~n31531 | n31525 | n31530;
  assign n36426 = n31538 | n31539;
  assign n36427 = n31551 | n31552;
  assign n36428 = n31557 | n31555 | n31556;
  assign n36429 = ~n31565 | n31559 | n31564;
  assign n36430 = n31572 | n31573;
  assign n36431 = n31585 | n31586;
  assign n36432 = n31591 | n31589 | n31590;
  assign n36433 = ~n31599 | n31593 | n31598;
  assign n36434 = n31606 | n31607;
  assign n36435 = n31619 | n31620;
  assign n36436 = n31625 | n31623 | n31624;
  assign n36437 = ~n31633 | n31627 | n31632;
  assign n36438 = n31640 | n31641;
  assign n36439 = n31653 | n31654;
  assign n36440 = n31659 | n31657 | n31658;
  assign n36441 = ~n31667 | n31661 | n31666;
  assign n36442 = n31674 | n31675;
  assign n36443 = n31687 | n31688;
  assign n36444 = n31693 | n31691 | n31692;
  assign n36445 = ~n31701 | n31695 | n31700;
  assign n36446 = n31708 | n31709;
  assign n36447 = n31721 | n31722;
  assign n36448 = n31727 | n31725 | n31726;
  assign n36449 = ~n31735 | n31729 | n31734;
  assign n36450 = n31742 | n31743;
  assign n36451 = n31755 | n31756;
  assign n36452 = n31761 | n31759 | n31760;
  assign n36453 = ~n31769 | n31763 | n31768;
  assign n36454 = n31776 | n31777;
  assign n36455 = n31789 | n31790;
  assign n36456 = n31795 | n31793 | n31794;
  assign n36457 = ~n31803 | n31797 | n31802;
  assign n36458 = n31810 | n31811;
  assign n36459 = n31823 | n31824;
  assign n36460 = n31829 | n31827 | n31828;
  assign n36461 = ~n31837 | n31831 | n31836;
  assign n36462 = n31844 | n31845;
  assign n36463 = n31857 | n31858;
  assign n36464 = n31863 | n31861 | n31862;
  assign n36465 = ~n31871 | n31865 | n31870;
  assign n36466 = n31878 | n31879;
  assign n36467 = n31891 | n31892;
  assign n36468 = n31897 | n31895 | n31896;
  assign n36469 = ~n31905 | n31899 | n31904;
  assign n36470 = n31912 | n31913;
  assign n36471 = n31925 | n31926;
  assign n36472 = n31931 | n31929 | n31930;
  assign n36473 = ~n31939 | n31933 | n31938;
  assign n36474 = n31946 | n31947;
  assign n36475 = n31959 | n31960;
  assign n36476 = n31965 | n31963 | n31964;
  assign n36477 = ~n31973 | n31967 | n31972;
  assign n36478 = n31980 | n31981;
  assign n36479 = n31993 | n31994;
  assign n36480 = n31999 | n31997 | n31998;
  assign n36481 = ~n32007 | n32001 | n32006;
  assign n36482 = n32014 | n32015;
  assign n36483 = n32027 | n32028;
  assign n36484 = n32033 | n32031 | n32032;
  assign n36485 = ~n32041 | n32035 | n32040;
  assign n36486 = n32048 | n32049;
  assign n36487 = n32061 | n32062;
  assign n36488 = n32067 | n32065 | n32066;
  assign n36489 = ~n32075 | n32069 | n32074;
  assign n36490 = n32082 | n32083;
  assign n36491 = n32095 | n32096;
  assign n36492 = n32101 | n32099 | n32100;
  assign n36493 = ~n32109 | n32103 | n32108;
  assign n36494 = n32116 | n32117;
  assign n36495 = n32122 | n32123;
  assign n36496 = n32130 | ~n32131;
  assign n36497 = n32142 | n32143;
  assign n36498 = n32152 | n32153;
  assign n36499 = n32158 | n32156 | n32157;
  assign n36500 = n32164 | n32165;
  assign n36501 = n32166 | n32167;
  assign n36502 = n32174 | n32175;
  assign n36503 = n32189 | n32190;
  assign n36504 = n32193 | n32194;
  assign n36505 = n32200 | n32201;
  assign n36506 = n32206 | n32203 | n32205;
  assign n36507 = n32209 | n32210;
  assign n36508 = n32216 | n32217;
  assign n36509 = n32224 | n32225;
  assign n36510 = n32234 | n32231 | n32233;
  assign n36511 = n32238 | n32239;
  assign po0  = ~n36511;
  assign po1  = ~n30836;
  assign po2  = ~n29813;
  assign po3  = ~n28917;
  assign po4  = ~n27931;
  assign po5  = ~n27055;
  assign po6  = ~n26098;
  assign po7  = ~n25256;
  assign po8  = ~n24331;
  assign po9  = ~n23517;
  assign po10  = ~n22625;
  assign po11  = ~n21842;
  assign po12  = ~n20986;
  assign po13  = ~n20229;
  assign po14  = ~n19401;
  assign po15  = ~n18676;
  assign po16  = ~n17885;
  assign po17  = ~n17187;
  assign po18  = ~n16428;
  assign po19  = ~n15760;
  assign po20  = ~n15033;
  assign po21  = ~n14394;
  assign po22  = ~n13704;
  assign po23  = ~n13099;
  assign po24  = ~n12442;
  assign po25  = ~n11858;
  assign po26  = ~n11229;
  assign po27  = ~n10681;
  assign po28  = ~n10086;
  assign po29  = ~n9565;
  assign po30  = ~n8998;
  assign po31  = ~n8506;
  assign po32  = ~n7975;
  assign po33  = ~n7512;
  assign po34  = ~n7015;
  assign po35  = ~n6579;
  assign po36  = ~n6117;
  assign po37  = ~n5708;
  assign po38  = ~n5278;
  assign po39  = ~n4903;
  assign po40  = ~n4508;
  assign po41  = ~n4155;
  assign po42  = ~n3788;
  assign po43  = ~n3473;
  assign po44  = ~n3140;
  assign po45  = ~n2855;
  assign po46  = ~n2556;
  assign po47  = ~n2301;
  assign po48  = ~n2038;
  assign po49  = ~n1812;
  assign po50  = ~n1582;
  assign po51  = ~n1388;
  assign po52  = ~n1192;
  assign po53  = ~n1028;
  assign po54  = ~n866;
  assign po55  = ~n730;
  assign po56  = ~n602;
  assign po57  = ~n497;
  assign po58  = ~n403;
  assign po59  = ~n330;
  assign po60  = ~n271;
  assign po61  = ~n217;
  assign po62  = ~n198;
  assign po63  = ~n193;
endmodule
