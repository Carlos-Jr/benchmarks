module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10   );
  input  pi0 , pi1 , pi2 ,
    pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 ;
  output po0 , po1 , po2 ,
    po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 ;
  wire n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n414, n415, n416, n417, n418,
    n419, n420, n422, n423, n424, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589,
    n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n646, n647,
    n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n682, n683,
    n684, n685, n686, n687;
  assign n22 = ~pi3  & ~pi5 ;
  assign n23 = ~pi1  & pi9 ;
  assign n24 = ~pi0  & pi9 ;
  assign n25 = pi1  & ~n24;
  assign n26 = n22 & ~n23;
  assign n27 = ~n25 & n26;
  assign n28 = pi0  & ~pi9 ;
  assign n29 = ~pi1  & ~n28;
  assign n30 = pi1  & ~pi9 ;
  assign n31 = ~pi7  & ~n30;
  assign n32 = ~n29 & n31;
  assign n33 = ~n27 & ~n32;
  assign n34 = ~pi2  & ~n33;
  assign n35 = ~pi0  & pi5 ;
  assign n36 = pi0  & ~pi1 ;
  assign n37 = pi2  & ~n36;
  assign n38 = ~n35 & ~n37;
  assign n39 = ~pi9  & ~n38;
  assign n40 = ~pi2  & ~pi3 ;
  assign n41 = pi9  & ~n40;
  assign n42 = pi0  & pi3 ;
  assign n43 = ~n41 & ~n42;
  assign n44 = ~pi1  & ~n43;
  assign n45 = pi1  & ~pi3 ;
  assign n46 = ~n39 & ~n45;
  assign n47 = ~n44 & n46;
  assign n48 = ~pi7  & ~n47;
  assign n49 = ~n34 & ~n48;
  assign n50 = ~pi8  & ~n49;
  assign n51 = ~pi5  & pi7 ;
  assign n52 = pi8  & n51;
  assign n53 = ~pi7  & pi9 ;
  assign n54 = ~n52 & ~n53;
  assign n55 = pi1  & ~n54;
  assign n56 = pi1  & ~pi7 ;
  assign n57 = ~pi5  & ~pi9 ;
  assign n58 = ~n56 & n57;
  assign n59 = ~n55 & ~n58;
  assign n60 = pi0  & ~pi2 ;
  assign n61 = ~n59 & n60;
  assign n62 = ~pi0  & ~pi1 ;
  assign n63 = pi2  & ~pi9 ;
  assign n64 = n62 & n63;
  assign n65 = n52 & n64;
  assign n66 = ~n61 & ~n65;
  assign n67 = ~pi3  & ~n66;
  assign n68 = ~n50 & ~n67;
  assign n69 = ~pi6  & ~n68;
  assign n70 = ~pi1  & ~pi9 ;
  assign n71 = ~pi8  & n70;
  assign n72 = ~pi0  & n40;
  assign n73 = n71 & n72;
  assign n74 = ~pi0  & ~pi2 ;
  assign n75 = n23 & n74;
  assign n76 = ~pi5  & ~n75;
  assign n77 = pi6  & ~n76;
  assign n78 = ~pi0  & ~pi9 ;
  assign n79 = pi0  & pi9 ;
  assign n80 = ~n78 & ~n79;
  assign n81 = pi1  & pi5 ;
  assign n82 = pi2  & n81;
  assign n83 = ~n80 & n82;
  assign n84 = ~n77 & ~n83;
  assign n85 = pi8  & ~n84;
  assign n86 = ~pi1  & ~n24;
  assign n87 = ~pi8  & ~n86;
  assign n88 = n36 & n63;
  assign n89 = ~n87 & ~n88;
  assign n90 = ~pi5  & ~n89;
  assign n91 = ~n85 & ~n90;
  assign n92 = pi3  & ~n91;
  assign n93 = ~pi2  & ~n28;
  assign n94 = pi6  & ~n93;
  assign n95 = pi1  & n40;
  assign n96 = ~n80 & n95;
  assign n97 = ~n94 & ~n96;
  assign n98 = pi5  & ~n97;
  assign n99 = pi2  & pi9 ;
  assign n100 = ~pi2  & n30;
  assign n101 = ~n99 & ~n100;
  assign n102 = ~pi0  & ~pi3 ;
  assign n103 = pi6  & n102;
  assign n104 = ~n101 & n103;
  assign n105 = ~n98 & ~n104;
  assign n106 = pi8  & ~n105;
  assign n107 = pi1  & ~pi8 ;
  assign n108 = pi2  & ~pi3 ;
  assign n109 = n23 & n108;
  assign n110 = ~n107 & ~n109;
  assign n111 = ~pi0  & ~n110;
  assign n112 = ~pi2  & pi6 ;
  assign n113 = pi3  & ~n112;
  assign n114 = n70 & ~n113;
  assign n115 = ~n99 & ~n114;
  assign n116 = ~pi8  & ~n115;
  assign n117 = ~n111 & ~n116;
  assign n118 = ~pi5  & ~n117;
  assign n119 = ~n73 & ~n106;
  assign n120 = ~n118 & n119;
  assign n121 = ~n92 & n120;
  assign n122 = ~pi7  & ~n121;
  assign n123 = ~n69 & ~n122;
  assign n124 = ~pi4  & ~n123;
  assign n125 = ~pi1  & ~pi3 ;
  assign n126 = ~pi6  & pi8 ;
  assign n127 = pi5  & ~n126;
  assign n128 = pi4  & pi8 ;
  assign n129 = ~pi6  & ~pi9 ;
  assign n130 = ~n128 & ~n129;
  assign n131 = n127 & ~n130;
  assign n132 = pi6  & ~pi9 ;
  assign n133 = pi4  & pi9 ;
  assign n134 = ~n132 & ~n133;
  assign n135 = pi5  & pi6 ;
  assign n136 = ~pi8  & ~n135;
  assign n137 = ~n134 & n136;
  assign n138 = ~n131 & ~n137;
  assign n139 = ~pi7  & n74;
  assign n140 = n125 & n139;
  assign n141 = ~n138 & n140;
  assign po0  = n124 | n141;
  assign n143 = ~pi2  & ~pi8 ;
  assign n144 = n78 & n143;
  assign n145 = pi8  & n79;
  assign n146 = pi2  & n145;
  assign n147 = ~n144 & ~n146;
  assign n148 = pi5  & ~n147;
  assign n149 = ~pi5  & pi8 ;
  assign n150 = pi6  & pi9 ;
  assign n151 = ~n149 & ~n150;
  assign n152 = ~pi0  & ~n151;
  assign n153 = ~pi8  & n57;
  assign n154 = pi8  & n150;
  assign n155 = ~n153 & ~n154;
  assign n156 = ~n152 & n155;
  assign n157 = pi2  & ~n156;
  assign n158 = ~n148 & ~n157;
  assign n159 = ~pi4  & ~n158;
  assign n160 = ~pi6  & pi9 ;
  assign n161 = pi5  & ~pi8 ;
  assign n162 = ~n128 & ~n161;
  assign n163 = ~pi6  & ~n162;
  assign n164 = ~n133 & ~n163;
  assign n165 = n74 & ~n160;
  assign n166 = ~n164 & n165;
  assign n167 = ~n159 & ~n166;
  assign n168 = ~pi1  & ~n167;
  assign n169 = ~pi8  & pi9 ;
  assign n170 = n35 & n169;
  assign n171 = pi6  & pi8 ;
  assign n172 = pi0  & ~n171;
  assign n173 = ~n151 & n172;
  assign n174 = ~n170 & ~n173;
  assign n175 = ~pi2  & ~n174;
  assign n176 = ~pi6  & ~pi8 ;
  assign n177 = ~pi0  & pi6 ;
  assign n178 = ~pi2  & ~n177;
  assign n179 = n149 & ~n178;
  assign n180 = ~n176 & ~n179;
  assign n181 = ~pi9  & ~n180;
  assign n182 = ~n175 & ~n181;
  assign n183 = pi1  & ~n182;
  assign n184 = n63 & n126;
  assign n185 = ~n183 & ~n184;
  assign n186 = ~pi4  & ~n185;
  assign n187 = ~n168 & ~n186;
  assign n188 = ~pi3  & ~n187;
  assign n189 = pi1  & pi2 ;
  assign n190 = pi3  & n189;
  assign n191 = n161 & n190;
  assign n192 = ~pi1  & pi3 ;
  assign n193 = n143 & n192;
  assign n194 = ~n81 & ~n193;
  assign n195 = pi0  & ~n194;
  assign n196 = pi5  & ~n40;
  assign n197 = ~n190 & ~n196;
  assign n198 = ~n195 & n197;
  assign n199 = pi6  & ~n198;
  assign n200 = pi9  & ~n191;
  assign n201 = ~n199 & n200;
  assign n202 = ~pi1  & ~pi8 ;
  assign n203 = ~pi1  & pi6 ;
  assign n204 = pi2  & ~n203;
  assign n205 = pi3  & ~n202;
  assign n206 = ~n204 & n205;
  assign n207 = ~pi0  & pi8 ;
  assign n208 = ~pi1  & ~pi6 ;
  assign n209 = pi0  & pi1 ;
  assign n210 = ~pi2  & ~n207;
  assign n211 = ~n208 & ~n209;
  assign n212 = n210 & n211;
  assign n213 = ~n206 & ~n212;
  assign n214 = ~pi5  & ~n213;
  assign n215 = pi3  & pi8 ;
  assign n216 = ~pi2  & ~n215;
  assign n217 = ~pi0  & ~n216;
  assign n218 = pi5  & n143;
  assign n219 = ~pi3  & ~pi8 ;
  assign n220 = ~n149 & ~n219;
  assign n221 = pi0  & n220;
  assign n222 = ~n218 & ~n221;
  assign n223 = ~pi1  & ~n222;
  assign n224 = ~pi2  & pi8 ;
  assign n225 = pi0  & n224;
  assign n226 = pi0  & ~pi5 ;
  assign n227 = ~n35 & ~n226;
  assign n228 = ~n225 & n227;
  assign n229 = pi1  & ~n228;
  assign n230 = ~n217 & ~n229;
  assign n231 = ~n223 & n230;
  assign n232 = ~pi6  & ~n231;
  assign n233 = ~pi9  & ~n214;
  assign n234 = ~n232 & n233;
  assign n235 = ~pi4  & ~n201;
  assign n236 = ~n234 & n235;
  assign n237 = ~n188 & ~n236;
  assign n238 = ~pi7  & ~n237;
  assign n239 = n30 & n224;
  assign n240 = n93 & ~n209;
  assign n241 = pi2  & ~n62;
  assign n242 = ~pi8  & ~n241;
  assign n243 = ~n240 & n242;
  assign n244 = ~n239 & ~n243;
  assign n245 = pi7  & ~n244;
  assign n246 = ~n64 & ~n245;
  assign n247 = ~pi6  & n22;
  assign n248 = ~pi4  & n247;
  assign n249 = ~n246 & n248;
  assign po1  = n238 | n249;
  assign n251 = pi6  & ~pi8 ;
  assign n252 = ~pi3  & pi9 ;
  assign n253 = pi1  & n252;
  assign n254 = n251 & n253;
  assign n255 = pi3  & ~n224;
  assign n256 = pi5  & ~n255;
  assign n257 = pi2  & ~pi5 ;
  assign n258 = pi3  & ~n257;
  assign n259 = pi8  & ~n258;
  assign n260 = ~n256 & ~n259;
  assign n261 = pi1  & ~n260;
  assign n262 = ~pi5  & pi6 ;
  assign n263 = ~pi3  & n262;
  assign n264 = n202 & n263;
  assign n265 = ~n261 & ~n264;
  assign n266 = ~pi9  & ~n265;
  assign n267 = pi1  & pi8 ;
  assign n268 = pi6  & ~n267;
  assign n269 = ~pi9  & ~n268;
  assign n270 = ~pi2  & ~n269;
  assign n271 = ~pi8  & n23;
  assign n272 = ~n270 & ~n271;
  assign n273 = pi3  & ~n272;
  assign n274 = pi2  & ~n126;
  assign n275 = pi1  & ~n274;
  assign n276 = pi5  & ~n216;
  assign n277 = ~n275 & n276;
  assign n278 = ~n45 & ~n169;
  assign n279 = ~pi6  & ~n252;
  assign n280 = ~n278 & n279;
  assign n281 = ~n254 & ~n280;
  assign n282 = ~n277 & n281;
  assign n283 = ~n273 & n282;
  assign n284 = ~n266 & n283;
  assign n285 = ~pi4  & ~n284;
  assign n286 = pi8  & ~pi9 ;
  assign n287 = ~pi5  & ~n176;
  assign n288 = ~n286 & n287;
  assign n289 = ~pi3  & pi4 ;
  assign n290 = ~pi2  & n289;
  assign n291 = ~pi1  & n290;
  assign n292 = ~n288 & n291;
  assign n293 = ~n285 & ~n292;
  assign n294 = ~pi0  & ~n293;
  assign n295 = ~pi5  & n99;
  assign n296 = ~n169 & ~n286;
  assign n297 = pi5  & ~n207;
  assign n298 = n296 & n297;
  assign n299 = ~n295 & ~n298;
  assign n300 = pi1  & ~n299;
  assign n301 = ~n70 & n296;
  assign n302 = pi2  & ~n301;
  assign n303 = ~n300 & ~n302;
  assign n304 = ~pi3  & ~n303;
  assign n305 = ~pi1  & pi8 ;
  assign n306 = n41 & n305;
  assign n307 = pi5  & ~n192;
  assign n308 = ~pi8  & ~pi9 ;
  assign n309 = ~pi2  & n308;
  assign n310 = ~n307 & n309;
  assign n311 = ~n306 & ~n310;
  assign n312 = pi0  & ~n311;
  assign n313 = ~n304 & ~n312;
  assign n314 = ~pi6  & ~n313;
  assign n315 = pi6  & ~n23;
  assign n316 = ~n30 & ~n315;
  assign n317 = pi8  & ~n316;
  assign n318 = pi1  & pi9 ;
  assign n319 = ~n70 & ~n318;
  assign n320 = n219 & ~n319;
  assign n321 = ~n317 & ~n320;
  assign n322 = ~pi2  & ~n321;
  assign n323 = pi2  & n318;
  assign n324 = ~n305 & ~n323;
  assign n325 = pi6  & ~n324;
  assign n326 = pi8  & ~n63;
  assign n327 = pi2  & n308;
  assign n328 = ~n326 & ~n327;
  assign n329 = ~n325 & n328;
  assign n330 = pi3  & ~n329;
  assign n331 = ~n322 & ~n330;
  assign n332 = n226 & ~n331;
  assign n333 = ~n314 & ~n332;
  assign n334 = ~pi4  & ~n333;
  assign n335 = ~n294 & ~n334;
  assign n336 = ~pi7  & ~n335;
  assign n337 = pi8  & pi9 ;
  assign n338 = pi7  & n337;
  assign n339 = pi0  & ~n338;
  assign n340 = n25 & ~n339;
  assign n341 = n28 & n202;
  assign n342 = ~n340 & ~n341;
  assign n343 = ~pi5  & ~pi6 ;
  assign n344 = ~pi4  & n40;
  assign n345 = n343 & n344;
  assign n346 = ~n342 & n345;
  assign po2  = n336 | n346;
  assign n348 = pi6  & ~n40;
  assign n349 = pi3  & ~pi9 ;
  assign n350 = ~n348 & ~n349;
  assign n351 = ~pi4  & ~n350;
  assign n352 = ~pi5  & ~n337;
  assign n353 = ~n135 & ~n343;
  assign n354 = n290 & ~n352;
  assign n355 = ~n353 & n354;
  assign n356 = ~n351 & ~n355;
  assign n357 = ~pi1  & ~n356;
  assign n358 = pi6  & n257;
  assign n359 = pi5  & pi9 ;
  assign n360 = ~n308 & ~n359;
  assign n361 = pi2  & ~n360;
  assign n362 = ~pi3  & ~n251;
  assign n363 = ~n361 & n362;
  assign n364 = pi1  & ~n127;
  assign n365 = ~n363 & n364;
  assign n366 = ~n358 & ~n365;
  assign n367 = ~pi4  & ~n366;
  assign n368 = ~n357 & ~n367;
  assign n369 = ~pi0  & ~n368;
  assign n370 = ~pi9  & n262;
  assign n371 = n267 & n370;
  assign n372 = pi2  & ~n220;
  assign n373 = pi5  & n224;
  assign n374 = ~n372 & ~n373;
  assign n375 = ~pi9  & ~n374;
  assign n376 = pi5  & n169;
  assign n377 = ~pi3  & ~n376;
  assign n378 = ~pi2  & ~n377;
  assign n379 = pi3  & ~pi8 ;
  assign n380 = ~pi6  & ~n379;
  assign n381 = pi3  & ~pi5 ;
  assign n382 = ~n380 & ~n381;
  assign n383 = ~n378 & ~n382;
  assign n384 = ~n375 & n383;
  assign n385 = pi1  & ~n384;
  assign n386 = n208 & n218;
  assign n387 = ~n263 & ~n386;
  assign n388 = ~pi9  & ~n387;
  assign n389 = ~n385 & ~n388;
  assign n390 = pi0  & ~n389;
  assign n391 = pi3  & ~pi6 ;
  assign n392 = pi2  & n391;
  assign n393 = ~n40 & n262;
  assign n394 = ~n392 & ~n393;
  assign n395 = pi9  & ~n394;
  assign n396 = ~n370 & ~n391;
  assign n397 = ~pi8  & ~n396;
  assign n398 = ~n395 & ~n397;
  assign n399 = ~pi1  & ~n398;
  assign n400 = ~n57 & ~n176;
  assign n401 = ~pi2  & ~n400;
  assign n402 = ~pi6  & ~n359;
  assign n403 = pi5  & pi8 ;
  assign n404 = ~n318 & ~n403;
  assign n405 = n402 & ~n404;
  assign n406 = ~n401 & ~n405;
  assign n407 = pi3  & ~n406;
  assign n408 = ~n371 & ~n407;
  assign n409 = ~n399 & n408;
  assign n410 = ~n390 & n409;
  assign n411 = ~pi4  & ~n410;
  assign n412 = ~n369 & ~n411;
  assign po3  = ~pi7  & ~n412;
  assign n414 = ~pi4  & n241;
  assign n415 = pi3  & ~pi4 ;
  assign n416 = ~n289 & ~n415;
  assign n417 = ~pi2  & n62;
  assign n418 = ~n416 & n417;
  assign n419 = ~n414 & ~n418;
  assign n420 = ~pi7  & n135;
  assign po4  = ~n419 & n420;
  assign n422 = n415 & ~n417;
  assign n423 = n62 & n290;
  assign n424 = ~n422 & ~n423;
  assign po5  = n420 & ~n424;
  assign n426 = ~pi1  & ~pi5 ;
  assign n427 = pi2  & ~n426;
  assign n428 = n129 & ~n427;
  assign n429 = pi5  & n318;
  assign n430 = ~n428 & ~n429;
  assign n431 = pi0  & ~n430;
  assign n432 = ~pi0  & pi2 ;
  assign n433 = ~n57 & n432;
  assign n434 = ~n431 & ~n433;
  assign n435 = pi8  & ~n434;
  assign n436 = pi9  & n432;
  assign n437 = ~n71 & ~n436;
  assign n438 = pi5  & ~n437;
  assign n439 = ~pi2  & pi9 ;
  assign n440 = ~n63 & ~n439;
  assign n441 = pi2  & pi8 ;
  assign n442 = ~n143 & ~n441;
  assign n443 = pi6  & n440;
  assign n444 = ~n442 & n443;
  assign n445 = ~n438 & ~n444;
  assign n446 = ~n435 & n445;
  assign n447 = ~pi7  & ~n446;
  assign n448 = pi7  & ~pi9 ;
  assign n449 = pi8  & ~n448;
  assign n450 = ~pi1  & pi2 ;
  assign n451 = ~n449 & n450;
  assign n452 = ~n100 & ~n451;
  assign n453 = ~pi0  & ~n452;
  assign n454 = pi1  & n145;
  assign n455 = ~n308 & ~n454;
  assign n456 = ~pi2  & pi7 ;
  assign n457 = ~n455 & n456;
  assign n458 = ~n453 & ~n457;
  assign n459 = n343 & ~n458;
  assign n460 = ~n447 & ~n459;
  assign n461 = ~pi3  & ~n460;
  assign n462 = n107 & ~n432;
  assign n463 = pi0  & n171;
  assign n464 = ~pi2  & n463;
  assign n465 = ~n462 & ~n464;
  assign n466 = pi9  & ~n465;
  assign n467 = ~pi0  & ~pi6 ;
  assign n468 = ~n202 & n467;
  assign n469 = ~n189 & ~n468;
  assign n470 = n319 & ~n469;
  assign n471 = ~pi1  & ~n308;
  assign n472 = pi0  & ~n30;
  assign n473 = ~n471 & n472;
  assign n474 = ~n470 & ~n473;
  assign n475 = ~pi5  & ~n474;
  assign n476 = ~pi0  & ~pi8 ;
  assign n477 = n30 & ~n226;
  assign n478 = ~n476 & n477;
  assign n479 = ~n466 & ~n478;
  assign n480 = ~n475 & n479;
  assign n481 = pi3  & ~n480;
  assign n482 = ~pi2  & pi5 ;
  assign n483 = ~n80 & n482;
  assign n484 = ~pi6  & ~n257;
  assign n485 = n24 & ~n484;
  assign n486 = ~n483 & ~n485;
  assign n487 = ~pi8  & ~n486;
  assign n488 = pi2  & ~n308;
  assign n489 = ~n145 & ~n488;
  assign n490 = pi6  & ~n489;
  assign n491 = ~n487 & ~n490;
  assign n492 = pi1  & ~n491;
  assign n493 = n24 & n441;
  assign n494 = pi8  & ~n226;
  assign n495 = ~pi2  & ~pi9 ;
  assign n496 = ~n467 & n495;
  assign n497 = ~n494 & n496;
  assign n498 = ~n493 & ~n497;
  assign n499 = ~pi1  & ~n498;
  assign n500 = ~n492 & ~n499;
  assign n501 = ~n481 & n500;
  assign n502 = ~pi7  & ~n501;
  assign n503 = ~n461 & ~n502;
  assign n504 = ~pi4  & ~n503;
  assign n505 = pi4  & n40;
  assign n506 = n62 & n505;
  assign n507 = ~n135 & ~n506;
  assign n508 = ~pi7  & ~n507;
  assign po6  = ~n504 & ~n508;
  assign n510 = n129 & n219;
  assign n511 = n207 & n391;
  assign n512 = ~n251 & ~n511;
  assign n513 = pi9  & ~n512;
  assign n514 = ~pi8  & ~n150;
  assign n515 = pi0  & ~n391;
  assign n516 = ~n132 & ~n515;
  assign n517 = ~n514 & ~n516;
  assign n518 = ~n513 & ~n517;
  assign n519 = ~pi2  & ~n518;
  assign n520 = pi0  & pi8 ;
  assign n521 = pi3  & ~n337;
  assign n522 = ~n520 & ~n521;
  assign n523 = ~pi6  & ~n522;
  assign n524 = ~pi3  & n337;
  assign n525 = ~n523 & ~n524;
  assign n526 = pi2  & ~n525;
  assign n527 = ~n510 & ~n519;
  assign n528 = ~n526 & n527;
  assign n529 = pi1  & ~n528;
  assign n530 = n177 & n296;
  assign n531 = ~n78 & ~n169;
  assign n532 = ~pi2  & ~pi6 ;
  assign n533 = ~n531 & n532;
  assign n534 = ~n530 & ~n533;
  assign n535 = pi3  & ~n534;
  assign n536 = ~pi0  & n143;
  assign n537 = ~n463 & ~n536;
  assign n538 = ~pi9  & ~n537;
  assign n539 = ~pi6  & ~n219;
  assign n540 = n488 & ~n539;
  assign n541 = ~n538 & ~n540;
  assign n542 = ~n535 & n541;
  assign n543 = ~pi1  & ~n542;
  assign n544 = pi3  & n143;
  assign n545 = n132 & n544;
  assign n546 = ~n543 & ~n545;
  assign n547 = ~n529 & n546;
  assign n548 = ~pi5  & ~n547;
  assign n549 = pi0  & ~n440;
  assign n550 = ~pi9  & n35;
  assign n551 = ~n549 & ~n550;
  assign n552 = pi8  & ~n551;
  assign n553 = n99 & n161;
  assign n554 = ~n552 & ~n553;
  assign n555 = ~pi3  & ~n554;
  assign n556 = pi3  & n482;
  assign n557 = pi3  & pi5 ;
  assign n558 = ~n63 & ~n557;
  assign n559 = n476 & ~n558;
  assign n560 = ~n556 & ~n559;
  assign n561 = ~n337 & ~n560;
  assign n562 = ~n555 & ~n561;
  assign n563 = pi1  & ~n562;
  assign n564 = n42 & n327;
  assign n565 = pi2  & pi3 ;
  assign n566 = ~n296 & ~n565;
  assign n567 = ~pi2  & ~n42;
  assign n568 = pi5  & ~n567;
  assign n569 = ~n566 & n568;
  assign n570 = ~n564 & ~n569;
  assign n571 = ~pi1  & ~n570;
  assign n572 = pi8  & n359;
  assign n573 = n565 & n572;
  assign n574 = ~n571 & ~n573;
  assign n575 = ~n563 & n574;
  assign n576 = ~pi6  & ~n575;
  assign n577 = ~n548 & ~n576;
  assign n578 = ~pi7  & ~n577;
  assign n579 = ~n296 & n432;
  assign n580 = n225 & n448;
  assign n581 = ~n579 & ~n580;
  assign n582 = n22 & n208;
  assign n583 = ~n581 & n582;
  assign n584 = ~n578 & ~n583;
  assign n585 = ~pi4  & ~n584;
  assign n586 = pi4  & ~pi7 ;
  assign n587 = n22 & n586;
  assign n588 = n417 & n587;
  assign n589 = ~pi6  & n588;
  assign po7  = ~n585 & ~n589;
  assign n591 = ~pi2  & ~n81;
  assign n592 = ~n381 & n591;
  assign n593 = ~n102 & n592;
  assign n594 = n22 & n36;
  assign n595 = ~n593 & ~n594;
  assign n596 = pi8  & ~n595;
  assign n597 = ~pi5  & ~n207;
  assign n598 = n189 & ~n557;
  assign n599 = ~n597 & n598;
  assign n600 = ~n596 & ~n599;
  assign n601 = ~pi9  & ~n600;
  assign n602 = n319 & ~n426;
  assign n603 = n108 & ~n602;
  assign n604 = n70 & n482;
  assign n605 = ~n253 & ~n604;
  assign n606 = ~pi0  & ~n605;
  assign n607 = ~n70 & ~n252;
  assign n608 = n592 & n607;
  assign n609 = ~n603 & ~n606;
  assign n610 = ~n608 & n609;
  assign n611 = ~pi8  & ~n610;
  assign n612 = ~n257 & ~n557;
  assign n613 = pi1  & ~n255;
  assign n614 = ~n612 & n613;
  assign n615 = ~n35 & n192;
  assign n616 = n224 & n615;
  assign n617 = ~n614 & ~n616;
  assign n618 = pi9  & ~n617;
  assign n619 = ~n611 & ~n618;
  assign n620 = ~n601 & n619;
  assign n621 = ~pi6  & ~n620;
  assign n622 = pi2  & ~n471;
  assign n623 = ~n315 & ~n622;
  assign n624 = pi0  & ~n623;
  assign n625 = ~pi6  & ~n107;
  assign n626 = pi2  & ~n625;
  assign n627 = pi6  & ~n337;
  assign n628 = ~n471 & n627;
  assign n629 = ~n626 & ~n628;
  assign n630 = ~n624 & n629;
  assign n631 = n381 & ~n630;
  assign n632 = ~n621 & ~n631;
  assign n633 = ~pi7  & ~n632;
  assign n634 = ~pi0  & ~n442;
  assign n635 = ~n225 & ~n634;
  assign n636 = ~pi9  & ~n635;
  assign n637 = ~pi8  & n436;
  assign n638 = ~n636 & ~n637;
  assign n639 = ~pi1  & ~n638;
  assign n640 = n318 & n536;
  assign n641 = ~n639 & ~n640;
  assign n642 = n247 & ~n641;
  assign n643 = ~n633 & ~n642;
  assign n644 = ~pi4  & ~n643;
  assign po8  = ~n588 & ~n644;
  assign n646 = ~pi2  & n125;
  assign n647 = pi4  & ~n646;
  assign n648 = n352 & n392;
  assign n649 = ~pi3  & ~n57;
  assign n650 = pi3  & ~n150;
  assign n651 = n207 & ~n650;
  assign n652 = ~n649 & ~n651;
  assign n653 = ~pi2  & ~n652;
  assign n654 = ~pi6  & ~n572;
  assign n655 = ~pi3  & ~n654;
  assign n656 = ~n648 & ~n655;
  assign n657 = ~n653 & n656;
  assign n658 = pi1  & ~n657;
  assign n659 = n289 & ~n343;
  assign n660 = n207 & ~n402;
  assign n661 = n650 & ~n660;
  assign n662 = ~pi2  & ~n659;
  assign n663 = ~n661 & n662;
  assign n664 = n108 & ~n308;
  assign n665 = ~n352 & n664;
  assign n666 = ~n663 & ~n665;
  assign n667 = ~pi1  & ~n666;
  assign n668 = n226 & n392;
  assign n669 = ~pi7  & ~n668;
  assign n670 = ~n471 & ~n669;
  assign n671 = ~pi7  & ~n646;
  assign n672 = pi0  & ~n671;
  assign n673 = pi7  & ~n108;
  assign n674 = ~pi5  & ~n108;
  assign n675 = pi6  & ~n674;
  assign n676 = ~n647 & ~n673;
  assign n677 = ~n675 & n676;
  assign n678 = ~n672 & n677;
  assign n679 = ~n670 & n678;
  assign n680 = ~n658 & n679;
  assign po9  = ~n667 & n680;
  assign n682 = pi8  & ~n25;
  assign n683 = pi2  & n415;
  assign n684 = ~n29 & n683;
  assign n685 = ~n682 & n684;
  assign n686 = ~n423 & ~n685;
  assign n687 = ~pi7  & n343;
  assign po10  = ~n686 & n687;
endmodule
