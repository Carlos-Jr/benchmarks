module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 , pi10 , pi11 , pi12 ,
    pi13 , pi14 , pi15 , pi16 , pi17 , pi18 ,
    pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 ,
    pi31 , pi32 , pi33 , pi34 , pi35 , pi36 ,
    pi37 , pi38 , pi39 , pi40 , pi41 , pi42 ,
    pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 , pi60 ,
    pi61 , pi62 , pi63 , pi64 , pi65 , pi66 ,
    pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 ,
    pi79 , pi80 , pi81 , pi82 , pi83 , pi84 ,
    pi85 , pi86 , pi87 , pi88 , pi89 , pi90 ,
    pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 ,
    pi109 , pi110 , pi111 , pi112 , pi113 , pi114 ,
    pi115 , pi116 , pi117 , pi118 , pi119 , pi120 ,
    pi121 , pi122 , pi123 , pi124 , pi125 , pi126 ,
    pi127 , pi128 , pi129 , pi130 , pi131 , pi132 , pi133 ,
    pi134 , pi135 , pi136 , pi137 , pi138 , pi139 ,
    pi140 , pi141 , pi142 , pi143 , pi144 , pi145 ,
    pi146 , pi147 , pi148 , pi149 , pi150 , pi151 ,
    pi152 , pi153 , pi154 , pi155 , pi156 , pi157 ,
    pi158 , pi159 , pi160 , pi161 , pi162 , pi163 ,
    pi164 , pi165 , pi166 , pi167 , pi168 , pi169 ,
    pi170 , pi171 , pi172 , pi173 , pi174 , pi175 ,
    pi176 , pi177 , pi178 , pi179 , pi180 , pi181 ,
    pi182 , pi183 , pi184 , pi185 , pi186 , pi187 ,
    pi188 , pi189 , pi190 , pi191 , pi192 , pi193 ,
    pi194 , pi195 , pi196 , pi197 , pi198 , pi199 ,
    pi200 , pi201 , pi202 , pi203 , pi204 , pi205 ,
    pi206 , pi207 , pi208 , pi209 , pi210 , pi211 ,
    pi212 , pi213 , pi214 , pi215 , pi216 , pi217 ,
    pi218 , pi219 , pi220 , pi221 , pi222 , pi223 ,
    pi224 , pi225 , pi226 , pi227 , pi228 , pi229 ,
    pi230 , pi231 , pi232 , pi233 , pi234 , pi235 ,
    pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 ,
    pi248 , pi249 , pi250 , pi251 , pi252 , pi253 ,
    pi254 , pi255 , pi256 , pi257 , pi258 , pi259 ,
    pi260 , pi261 , pi262 , pi263 , pi264 , pi265 , pi266 ,
    pi267 , pi268 , pi269 , pi270 , pi271 , pi272 ,
    pi273 , pi274 , pi275 , pi276 , pi277 , pi278 ,
    pi279 , pi280 , pi281 , pi282 , pi283 , pi284 ,
    pi285 , pi286 , pi287 , pi288 , pi289 , pi290 ,
    pi291 , pi292 , pi293 , pi294 , pi295 , pi296 ,
    pi297 , pi298 , pi299 , pi300 , pi301 , pi302 ,
    pi303 , pi304 , pi305 , pi306 , pi307 , pi308 ,
    pi309 , pi310 , pi311 , pi312 , pi313 , pi314 ,
    pi315 , pi316 , pi317 , pi318 , pi319 , pi320 ,
    pi321 , pi322 , pi323 , pi324 , pi325 , pi326 ,
    pi327 , pi328 , pi329 , pi330 , pi331 , pi332 ,
    pi333 , pi334 , pi335 , pi336 , pi337 , pi338 ,
    pi339 , pi340 , pi341 , pi342 , pi343 , pi344 ,
    pi345 , pi346 , pi347 , pi348 , pi349 , pi350 ,
    pi351 , pi352 , pi353 , pi354 , pi355 , pi356 ,
    pi357 , pi358 , pi359 , pi360 , pi361 , pi362 ,
    pi363 , pi364 , pi365 , pi366 , pi367 , pi368 ,
    pi369 , pi370 , pi371 , pi372 , pi373 , pi374 ,
    pi375 , pi376 , pi377 , pi378 , pi379 , pi380 ,
    pi381 , pi382 , pi383 , pi384 , pi385 , pi386 ,
    pi387 , pi388 , pi389 , pi390 , pi391 , pi392 , pi393 ,
    pi394 , pi395 , pi396 , pi397 , pi398 , pi399 ,
    pi400 , pi401 , pi402 , pi403 , pi404 , pi405 ,
    pi406 , pi407 , pi408 , pi409 , pi410 , pi411 ,
    pi412 , pi413 , pi414 , pi415 , pi416 , pi417 ,
    pi418 , pi419 , pi420 , pi421 , pi422 , pi423 ,
    pi424 , pi425 , pi426 , pi427 , pi428 , pi429 ,
    pi430 , pi431 , pi432 , pi433 , pi434 , pi435 ,
    pi436 , pi437 , pi438 , pi439 , pi440 , pi441 ,
    pi442 , pi443 , pi444 , pi445 , pi446 , pi447 ,
    pi448 , pi449 , pi450 , pi451 , pi452 , pi453 ,
    pi454 , pi455 , pi456 , pi457 , pi458 , pi459 ,
    pi460 , pi461 , pi462 , pi463 , pi464 , pi465 ,
    pi466 , pi467 , pi468 , pi469 , pi470 , pi471 ,
    pi472 , pi473 , pi474 , pi475 , pi476 , pi477 ,
    pi478 , pi479 , pi480 , pi481 , pi482 , pi483 ,
    pi484 , pi485 , pi486 , pi487 , pi488 , pi489 ,
    pi490 , pi491 , pi492 , pi493 , pi494 , pi495 ,
    pi496 , pi497 , pi498 , pi499 , pi500 , pi501 ,
    pi502 , pi503 , pi504 , pi505 , pi506 , pi507 ,
    pi508 , pi509 , pi510 , pi511 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ,
    po128 , po129   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 ,
    pi6 , pi7 , pi8 , pi9 , pi10 , pi11 ,
    pi12 , pi13 , pi14 , pi15 , pi16 , pi17 ,
    pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 , pi35 ,
    pi36 , pi37 , pi38 , pi39 , pi40 , pi41 ,
    pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 ,
    pi54 , pi55 , pi56 , pi57 , pi58 , pi59 ,
    pi60 , pi61 , pi62 , pi63 , pi64 , pi65 ,
    pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 ,
    pi78 , pi79 , pi80 , pi81 , pi82 , pi83 ,
    pi84 , pi85 , pi86 , pi87 , pi88 , pi89 ,
    pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 ,
    pi102 , pi103 , pi104 , pi105 , pi106 , pi107 ,
    pi108 , pi109 , pi110 , pi111 , pi112 , pi113 ,
    pi114 , pi115 , pi116 , pi117 , pi118 , pi119 ,
    pi120 , pi121 , pi122 , pi123 , pi124 , pi125 ,
    pi126 , pi127 , pi128 , pi129 , pi130 , pi131 ,
    pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 ,
    pi139 , pi140 , pi141 , pi142 , pi143 , pi144 ,
    pi145 , pi146 , pi147 , pi148 , pi149 , pi150 ,
    pi151 , pi152 , pi153 , pi154 , pi155 , pi156 ,
    pi157 , pi158 , pi159 , pi160 , pi161 , pi162 ,
    pi163 , pi164 , pi165 , pi166 , pi167 , pi168 ,
    pi169 , pi170 , pi171 , pi172 , pi173 , pi174 ,
    pi175 , pi176 , pi177 , pi178 , pi179 , pi180 ,
    pi181 , pi182 , pi183 , pi184 , pi185 , pi186 ,
    pi187 , pi188 , pi189 , pi190 , pi191 , pi192 ,
    pi193 , pi194 , pi195 , pi196 , pi197 , pi198 ,
    pi199 , pi200 , pi201 , pi202 , pi203 , pi204 ,
    pi205 , pi206 , pi207 , pi208 , pi209 , pi210 ,
    pi211 , pi212 , pi213 , pi214 , pi215 , pi216 ,
    pi217 , pi218 , pi219 , pi220 , pi221 , pi222 ,
    pi223 , pi224 , pi225 , pi226 , pi227 , pi228 ,
    pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 ,
    pi241 , pi242 , pi243 , pi244 , pi245 , pi246 ,
    pi247 , pi248 , pi249 , pi250 , pi251 , pi252 ,
    pi253 , pi254 , pi255 , pi256 , pi257 , pi258 ,
    pi259 , pi260 , pi261 , pi262 , pi263 , pi264 , pi265 ,
    pi266 , pi267 , pi268 , pi269 , pi270 , pi271 ,
    pi272 , pi273 , pi274 , pi275 , pi276 , pi277 ,
    pi278 , pi279 , pi280 , pi281 , pi282 , pi283 ,
    pi284 , pi285 , pi286 , pi287 , pi288 , pi289 ,
    pi290 , pi291 , pi292 , pi293 , pi294 , pi295 ,
    pi296 , pi297 , pi298 , pi299 , pi300 , pi301 ,
    pi302 , pi303 , pi304 , pi305 , pi306 , pi307 ,
    pi308 , pi309 , pi310 , pi311 , pi312 , pi313 ,
    pi314 , pi315 , pi316 , pi317 , pi318 , pi319 ,
    pi320 , pi321 , pi322 , pi323 , pi324 , pi325 ,
    pi326 , pi327 , pi328 , pi329 , pi330 , pi331 ,
    pi332 , pi333 , pi334 , pi335 , pi336 , pi337 ,
    pi338 , pi339 , pi340 , pi341 , pi342 , pi343 ,
    pi344 , pi345 , pi346 , pi347 , pi348 , pi349 ,
    pi350 , pi351 , pi352 , pi353 , pi354 , pi355 ,
    pi356 , pi357 , pi358 , pi359 , pi360 , pi361 ,
    pi362 , pi363 , pi364 , pi365 , pi366 , pi367 ,
    pi368 , pi369 , pi370 , pi371 , pi372 , pi373 ,
    pi374 , pi375 , pi376 , pi377 , pi378 , pi379 ,
    pi380 , pi381 , pi382 , pi383 , pi384 , pi385 ,
    pi386 , pi387 , pi388 , pi389 , pi390 , pi391 , pi392 ,
    pi393 , pi394 , pi395 , pi396 , pi397 , pi398 ,
    pi399 , pi400 , pi401 , pi402 , pi403 , pi404 ,
    pi405 , pi406 , pi407 , pi408 , pi409 , pi410 ,
    pi411 , pi412 , pi413 , pi414 , pi415 , pi416 ,
    pi417 , pi418 , pi419 , pi420 , pi421 , pi422 ,
    pi423 , pi424 , pi425 , pi426 , pi427 , pi428 ,
    pi429 , pi430 , pi431 , pi432 , pi433 , pi434 ,
    pi435 , pi436 , pi437 , pi438 , pi439 , pi440 ,
    pi441 , pi442 , pi443 , pi444 , pi445 , pi446 ,
    pi447 , pi448 , pi449 , pi450 , pi451 , pi452 ,
    pi453 , pi454 , pi455 , pi456 , pi457 , pi458 ,
    pi459 , pi460 , pi461 , pi462 , pi463 , pi464 ,
    pi465 , pi466 , pi467 , pi468 , pi469 , pi470 ,
    pi471 , pi472 , pi473 , pi474 , pi475 , pi476 ,
    pi477 , pi478 , pi479 , pi480 , pi481 , pi482 ,
    pi483 , pi484 , pi485 , pi486 , pi487 , pi488 ,
    pi489 , pi490 , pi491 , pi492 , pi493 , pi494 ,
    pi495 , pi496 , pi497 , pi498 , pi499 , pi500 ,
    pi501 , pi502 , pi503 , pi504 , pi505 , pi506 ,
    pi507 , pi508 , pi509 , pi510 , pi511 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ,
    po128 , po129 ;
  wire n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061,
    n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331,
    n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231,
    n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3296, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321,
    n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561,
    n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591,
    n3592, n3593, n3594, n3595, n3596, n3597,
    n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621,
    n3622, n3623, n3624, n3625, n3626, n3627,
    n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651,
    n3652, n3653, n3654, n3655, n3656, n3657,
    n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681,
    n3682, n3683, n3684, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927,
    n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951,
    n3952, n3953, n3954, n3955, n3956, n3957,
    n3958, n3959, n3960, n3961, n3962, n3963,
    n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981,
    n3982, n3983, n3984, n3985, n3986, n3987,
    n3988, n3989, n3990, n3991, n3992, n3993,
    n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011,
    n4012, n4013, n4014, n4015, n4016, n4017,
    n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4047,
    n4048, n4049, n4050, n4051, n4052, n4053,
    n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4076, n4077,
    n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101,
    n4102, n4103, n4104, n4105, n4106, n4107,
    n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131,
    n4132, n4133, n4134, n4135, n4136, n4137,
    n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161,
    n4162, n4163, n4164, n4165, n4166, n4167,
    n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191,
    n4192, n4193, n4194, n4195, n4196, n4197,
    n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227,
    n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4249, n4250, n4251,
    n4252, n4253, n4254, n4255, n4256, n4257,
    n4258, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317,
    n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341,
    n4342, n4343, n4344, n4345, n4346, n4347,
    n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371,
    n4372, n4373, n4374, n4375, n4376, n4377,
    n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4394, n4395,
    n4396, n4397, n4398, n4399, n4400, n4401,
    n4402, n4403, n4404, n4405, n4406, n4407,
    n4408, n4409, n4410, n4411, n4412, n4413,
    n4414, n4415, n4416, n4417, n4418, n4419,
    n4420, n4421, n4422, n4423, n4424, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431,
    n4432, n4433, n4434, n4435, n4436, n4437,
    n4438, n4439, n4440, n4441, n4442, n4443,
    n4444, n4445, n4446, n4447, n4448, n4449,
    n4450, n4451, n4452, n4453, n4454, n4455,
    n4456, n4457, n4458, n4459, n4460, n4461,
    n4462, n4463, n4464, n4465, n4466, n4467,
    n4468, n4469, n4470, n4471, n4472, n4473,
    n4474, n4475, n4476, n4477, n4478, n4479,
    n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491,
    n4492, n4493, n4494, n4495, n4496, n4497,
    n4498, n4499, n4500, n4501, n4502, n4503,
    n4504, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515,
    n4516, n4517, n4518, n4519, n4520, n4521,
    n4522, n4523, n4524, n4525, n4526, n4527,
    n4528, n4529, n4530, n4531, n4532, n4533,
    n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551,
    n4552, n4553, n4554, n4555, n4556, n4557,
    n4558, n4559, n4560, n4561, n4562, n4563,
    n4564, n4565, n4566, n4567, n4568, n4569,
    n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581,
    n4582, n4583, n4584, n4585, n4586, n4587,
    n4588, n4589, n4590, n4591, n4592, n4593,
    n4594, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611,
    n4612, n4613, n4614, n4615, n4616, n4617,
    n4618, n4619, n4620, n4621, n4622, n4623,
    n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641,
    n4642, n4643, n4644, n4645, n4646, n4647,
    n4648, n4649, n4650, n4651, n4652, n4653,
    n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665,
    n4666, n4667, n4668, n4669, n4670, n4671,
    n4672, n4673, n4674, n4675, n4676, n4677,
    n4678, n4679, n4680, n4681, n4682, n4683,
    n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707,
    n4708, n4709, n4710, n4711, n4712, n4713,
    n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737,
    n4738, n4739, n4740, n4741, n4742, n4743,
    n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761,
    n4762, n4763, n4764, n4765, n4766, n4767,
    n4768, n4769, n4770, n4771, n4773, n4774,
    n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786,
    n4787, n4788, n4789, n4790, n4791, n4792,
    n4793, n4794, n4795, n4796, n4797, n4798,
    n4799, n4800, n4801, n4802, n4803, n4804,
    n4805, n4806, n4807, n4808, n4809, n4810,
    n4811, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822,
    n4823, n4824, n4825, n4826, n4827, n4828,
    n4829, n4830, n4831, n4832, n4833, n4834,
    n4835, n4836, n4837, n4838, n4839, n4840,
    n4841, n4842, n4843, n4844, n4845, n4846,
    n4847, n4848, n4849, n4850, n4851, n4852,
    n4853, n4854, n4855, n4856, n4857, n4858,
    n4859, n4860, n4861, n4862, n4863, n4864,
    n4865, n4866, n4867, n4868, n4869, n4870,
    n4871, n4872, n4873, n4874, n4875, n4876,
    n4877, n4878, n4879, n4880, n4881, n4882,
    n4883, n4884, n4885, n4886, n4887, n4888,
    n4889, n4890, n4891, n4892, n4893, n4894,
    n4895, n4896;
  assign n643 = ~pi28  & pi156 ;
  assign n644 = pi27  & ~pi155 ;
  assign n645 = ~pi27  & pi155 ;
  assign n646 = pi26  & ~pi154 ;
  assign n647 = ~pi26  & pi154 ;
  assign n648 = pi25  & ~pi153 ;
  assign n649 = ~pi25  & pi153 ;
  assign n650 = pi24  & ~pi152 ;
  assign n651 = ~pi24  & pi152 ;
  assign n652 = pi23  & ~pi151 ;
  assign n653 = ~pi23  & pi151 ;
  assign n654 = pi22  & ~pi150 ;
  assign n655 = ~pi22  & pi150 ;
  assign n656 = pi21  & ~pi149 ;
  assign n657 = ~pi21  & pi149 ;
  assign n658 = pi20  & ~pi148 ;
  assign n659 = ~pi20  & pi148 ;
  assign n660 = pi19  & ~pi147 ;
  assign n661 = ~pi19  & pi147 ;
  assign n662 = pi18  & ~pi146 ;
  assign n663 = ~pi18  & pi146 ;
  assign n664 = pi17  & ~pi145 ;
  assign n665 = ~pi17  & pi145 ;
  assign n666 = pi16  & ~pi144 ;
  assign n667 = ~pi16  & pi144 ;
  assign n668 = pi15  & ~pi143 ;
  assign n669 = ~pi15  & pi143 ;
  assign n670 = pi14  & ~pi142 ;
  assign n671 = ~pi14  & pi142 ;
  assign n672 = pi13  & ~pi141 ;
  assign n673 = ~pi13  & pi141 ;
  assign n674 = pi12  & ~pi140 ;
  assign n675 = ~pi12  & pi140 ;
  assign n676 = pi11  & ~pi139 ;
  assign n677 = ~pi11  & pi139 ;
  assign n678 = pi10  & ~pi138 ;
  assign n679 = ~pi10  & pi138 ;
  assign n680 = pi9  & ~pi137 ;
  assign n681 = ~pi9  & pi137 ;
  assign n682 = pi8  & ~pi136 ;
  assign n683 = ~pi8  & pi136 ;
  assign n684 = pi7  & ~pi135 ;
  assign n685 = ~pi7  & pi135 ;
  assign n686 = pi6  & ~pi134 ;
  assign n687 = ~pi6  & pi134 ;
  assign n688 = pi5  & ~pi133 ;
  assign n689 = ~pi5  & pi133 ;
  assign n690 = pi4  & ~pi132 ;
  assign n691 = ~pi4  & pi132 ;
  assign n692 = pi3  & ~pi131 ;
  assign n693 = ~pi3  & pi131 ;
  assign n694 = pi2  & ~pi130 ;
  assign n695 = pi1  & ~pi129 ;
  assign n696 = pi0  & ~pi128 ;
  assign n697 = ~n695 & ~n696;
  assign n698 = ~pi2  & pi130 ;
  assign n699 = ~pi1  & pi129 ;
  assign n700 = ~n698 & ~n699;
  assign n701 = n696 & ~n699;
  assign n702 = ~n695 & ~n701;
  assign n703 = ~n698 & ~n702;
  assign n704 = ~n697 & n700;
  assign n705 = ~n694 & ~n4553;
  assign n706 = ~n693 & ~n705;
  assign n707 = ~n692 & ~n706;
  assign n708 = ~n691 & ~n707;
  assign n709 = ~pi4  & n707;
  assign n710 = ~pi132  & ~n709;
  assign n711 = pi4  & ~n707;
  assign n712 = ~n710 & ~n711;
  assign n713 = ~n690 & ~n708;
  assign n714 = ~n689 & ~n4554;
  assign n715 = ~pi5  & n4554;
  assign n716 = ~pi133  & ~n715;
  assign n717 = pi5  & ~n4554;
  assign n718 = ~n716 & ~n717;
  assign n719 = ~n688 & ~n714;
  assign n720 = ~n687 & ~n4555;
  assign n721 = ~n686 & ~n720;
  assign n722 = ~n685 & ~n721;
  assign n723 = ~n684 & ~n722;
  assign n724 = ~n683 & ~n723;
  assign n725 = ~pi8  & n723;
  assign n726 = ~pi136  & ~n725;
  assign n727 = pi8  & ~n723;
  assign n728 = ~n726 & ~n727;
  assign n729 = ~n682 & ~n724;
  assign n730 = ~n681 & ~n4556;
  assign n731 = ~pi9  & n4556;
  assign n732 = ~pi137  & ~n731;
  assign n733 = pi9  & ~n4556;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~n680 & ~n730;
  assign n736 = ~n679 & ~n4557;
  assign n737 = ~n678 & ~n736;
  assign n738 = ~n677 & ~n737;
  assign n739 = ~n676 & ~n738;
  assign n740 = ~n675 & ~n739;
  assign n741 = ~n674 & ~n740;
  assign n742 = ~n673 & ~n741;
  assign n743 = ~n672 & ~n742;
  assign n744 = ~n671 & ~n743;
  assign n745 = ~n670 & ~n744;
  assign n746 = ~n669 & ~n745;
  assign n747 = ~n668 & ~n746;
  assign n748 = ~n667 & ~n747;
  assign n749 = ~pi16  & n747;
  assign n750 = ~pi144  & ~n749;
  assign n751 = pi16  & ~n747;
  assign n752 = ~n750 & ~n751;
  assign n753 = ~n666 & ~n748;
  assign n754 = ~n665 & ~n4558;
  assign n755 = ~pi17  & n4558;
  assign n756 = ~pi145  & ~n755;
  assign n757 = pi17  & ~n4558;
  assign n758 = ~n756 & ~n757;
  assign n759 = ~n664 & ~n754;
  assign n760 = ~n663 & ~n4559;
  assign n761 = ~n662 & ~n760;
  assign n762 = ~n661 & ~n761;
  assign n763 = ~n660 & ~n762;
  assign n764 = ~n659 & ~n763;
  assign n765 = ~n658 & ~n764;
  assign n766 = ~n657 & ~n765;
  assign n767 = ~n656 & ~n766;
  assign n768 = ~n655 & ~n767;
  assign n769 = ~n654 & ~n768;
  assign n770 = ~n653 & ~n769;
  assign n771 = ~n652 & ~n770;
  assign n772 = ~n651 & ~n771;
  assign n773 = ~pi24  & n771;
  assign n774 = ~pi152  & ~n773;
  assign n775 = pi24  & ~n771;
  assign n776 = ~n774 & ~n775;
  assign n777 = ~n650 & ~n772;
  assign n778 = ~n649 & ~n4560;
  assign n779 = ~pi25  & n4560;
  assign n780 = ~pi153  & ~n779;
  assign n781 = pi25  & ~n4560;
  assign n782 = ~n780 & ~n781;
  assign n783 = ~n648 & ~n778;
  assign n784 = ~n647 & ~n4561;
  assign n785 = ~n646 & ~n784;
  assign n786 = ~n645 & ~n785;
  assign n787 = ~n644 & ~n786;
  assign n788 = ~n643 & ~n787;
  assign n789 = pi28  & ~pi156 ;
  assign n790 = pi29  & ~pi157 ;
  assign n791 = ~n789 & ~n790;
  assign n792 = ~n788 & n791;
  assign n793 = ~pi29  & pi157 ;
  assign n794 = ~pi30  & pi158 ;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~n788 & ~n789;
  assign n797 = ~n793 & ~n796;
  assign n798 = ~n790 & ~n797;
  assign n799 = ~n794 & ~n798;
  assign n800 = ~n792 & n795;
  assign n801 = pi30  & ~pi158 ;
  assign n802 = pi31  & ~pi159 ;
  assign n803 = ~n801 & ~n802;
  assign n804 = ~n4562 & n803;
  assign n805 = ~pi39  & pi167 ;
  assign n806 = ~pi38  & pi166 ;
  assign n807 = ~n805 & ~n806;
  assign n808 = ~pi37  & pi165 ;
  assign n809 = ~pi36  & pi164 ;
  assign n810 = ~n808 & ~n809;
  assign n811 = n807 & n810;
  assign n812 = ~pi35  & pi163 ;
  assign n813 = ~pi34  & pi162 ;
  assign n814 = ~n812 & ~n813;
  assign n815 = ~pi33  & pi161 ;
  assign n816 = ~pi32  & pi160 ;
  assign n817 = ~pi31  & pi159 ;
  assign n818 = ~n816 & ~n817;
  assign n819 = ~n815 & ~n817;
  assign n820 = ~n816 & n819;
  assign n821 = ~n815 & n818;
  assign n822 = n814 & n4563;
  assign n823 = n811 & n822;
  assign n824 = ~n4562 & ~n801;
  assign n825 = ~n817 & ~n824;
  assign n826 = ~n802 & ~n825;
  assign n827 = n814 & ~n815;
  assign n828 = n811 & n827;
  assign n829 = ~n826 & n828;
  assign n830 = ~n816 & n829;
  assign n831 = ~n804 & n823;
  assign n832 = pi35  & ~pi163 ;
  assign n833 = pi32  & ~pi160 ;
  assign n834 = ~pi160  & ~n815;
  assign n835 = pi32  & n834;
  assign n836 = ~n815 & n833;
  assign n837 = pi33  & ~pi161 ;
  assign n838 = pi34  & ~pi162 ;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~n4565 & ~n837;
  assign n841 = ~n838 & n840;
  assign n842 = ~n4565 & n839;
  assign n843 = n814 & ~n4566;
  assign n844 = ~n832 & ~n843;
  assign n845 = n811 & ~n844;
  assign n846 = pi39  & ~pi167 ;
  assign n847 = pi36  & ~pi164 ;
  assign n848 = ~n808 & n847;
  assign n849 = pi38  & ~pi166 ;
  assign n850 = pi37  & ~pi165 ;
  assign n851 = ~n849 & ~n850;
  assign n852 = ~n848 & n851;
  assign n853 = n807 & ~n852;
  assign n854 = ~n848 & ~n850;
  assign n855 = n807 & ~n854;
  assign n856 = ~pi166  & ~n805;
  assign n857 = pi38  & n856;
  assign n858 = ~n805 & n849;
  assign n859 = ~n846 & ~n4567;
  assign n860 = ~n855 & n859;
  assign n861 = ~n846 & ~n853;
  assign n862 = ~n845 & ~n4567;
  assign n863 = ~n855 & n862;
  assign n864 = ~n846 & n863;
  assign n865 = ~n845 & n4568;
  assign n866 = ~n4564 & n4569;
  assign n867 = ~pi47  & pi175 ;
  assign n868 = ~pi46  & pi174 ;
  assign n869 = ~n867 & ~n868;
  assign n870 = ~pi45  & pi173 ;
  assign n871 = ~pi44  & pi172 ;
  assign n872 = ~n870 & ~n871;
  assign n873 = n869 & n872;
  assign n874 = ~pi43  & pi171 ;
  assign n875 = ~pi42  & pi170 ;
  assign n876 = ~n874 & ~n875;
  assign n877 = ~pi40  & pi168 ;
  assign n878 = ~pi41  & pi169 ;
  assign n879 = ~n877 & ~n878;
  assign n880 = n876 & n879;
  assign n881 = n873 & n880;
  assign n882 = ~n866 & n881;
  assign n883 = pi43  & ~pi171 ;
  assign n884 = pi40  & ~pi168 ;
  assign n885 = ~n878 & n884;
  assign n886 = pi41  & ~pi169 ;
  assign n887 = pi42  & ~pi170 ;
  assign n888 = ~n886 & ~n887;
  assign n889 = ~n885 & ~n886;
  assign n890 = ~n887 & n889;
  assign n891 = ~n885 & n888;
  assign n892 = n876 & ~n4570;
  assign n893 = ~n883 & ~n892;
  assign n894 = n873 & ~n893;
  assign n895 = pi47  & ~pi175 ;
  assign n896 = pi44  & ~pi172 ;
  assign n897 = ~n870 & n896;
  assign n898 = pi46  & ~pi174 ;
  assign n899 = pi45  & ~pi173 ;
  assign n900 = ~n898 & ~n899;
  assign n901 = ~n897 & n900;
  assign n902 = n869 & ~n901;
  assign n903 = ~n897 & ~n899;
  assign n904 = n869 & ~n903;
  assign n905 = ~pi174  & ~n867;
  assign n906 = pi46  & n905;
  assign n907 = ~n867 & n898;
  assign n908 = ~n895 & ~n4571;
  assign n909 = ~n904 & n908;
  assign n910 = ~n895 & ~n902;
  assign n911 = ~n894 & n4572;
  assign n912 = ~n882 & ~n4571;
  assign n913 = ~n904 & n912;
  assign n914 = ~n894 & n913;
  assign n915 = ~n895 & n914;
  assign n916 = ~n882 & n911;
  assign n917 = ~pi53  & pi181 ;
  assign n918 = ~pi52  & pi180 ;
  assign n919 = ~pi180  & ~n917;
  assign n920 = pi52  & ~n917;
  assign n921 = ~n919 & ~n920;
  assign n922 = ~n917 & ~n918;
  assign n923 = ~pi55  & pi183 ;
  assign n924 = ~pi54  & pi182 ;
  assign n925 = ~n923 & ~n924;
  assign n926 = ~n4574 & n925;
  assign n927 = ~pi51  & pi179 ;
  assign n928 = ~pi50  & pi178 ;
  assign n929 = ~n927 & ~n928;
  assign n930 = ~pi48  & pi176 ;
  assign n931 = ~pi49  & pi177 ;
  assign n932 = ~n930 & ~n931;
  assign n933 = n929 & n932;
  assign n934 = n925 & n932;
  assign n935 = n929 & n934;
  assign n936 = ~n4574 & n935;
  assign n937 = n929 & ~n931;
  assign n938 = n926 & n937;
  assign n939 = ~n930 & n938;
  assign n940 = n926 & n933;
  assign n941 = ~n4573 & n4575;
  assign n942 = pi51  & ~pi179 ;
  assign n943 = pi48  & ~pi176 ;
  assign n944 = ~pi176  & ~n931;
  assign n945 = pi48  & n944;
  assign n946 = ~n931 & n943;
  assign n947 = pi49  & ~pi177 ;
  assign n948 = pi50  & ~pi178 ;
  assign n949 = ~n947 & ~n948;
  assign n950 = ~n4576 & ~n947;
  assign n951 = ~n948 & n950;
  assign n952 = ~n4576 & n949;
  assign n953 = n929 & ~n4577;
  assign n954 = ~n942 & ~n953;
  assign n955 = n926 & ~n954;
  assign n956 = pi55  & ~pi183 ;
  assign n957 = pi52  & ~pi180 ;
  assign n958 = pi52  & n919;
  assign n959 = ~n917 & n957;
  assign n960 = pi53  & ~pi181 ;
  assign n961 = pi54  & ~pi182 ;
  assign n962 = ~n960 & ~n961;
  assign n963 = ~n4578 & ~n960;
  assign n964 = ~n961 & n963;
  assign n965 = ~n4578 & n962;
  assign n966 = n925 & ~n4579;
  assign n967 = ~n956 & ~n966;
  assign n968 = ~n4574 & ~n954;
  assign n969 = n4579 & ~n968;
  assign n970 = n925 & ~n969;
  assign n971 = ~n955 & ~n966;
  assign n972 = ~n956 & ~n4580;
  assign n973 = ~n955 & n967;
  assign n974 = ~n941 & n4581;
  assign n975 = ~pi63  & pi191 ;
  assign n976 = ~pi62  & pi190 ;
  assign n977 = ~n975 & ~n976;
  assign n978 = ~pi61  & pi189 ;
  assign n979 = ~pi60  & pi188 ;
  assign n980 = ~n978 & ~n979;
  assign n981 = n977 & n980;
  assign n982 = ~pi59  & pi187 ;
  assign n983 = ~pi58  & pi186 ;
  assign n984 = ~n982 & ~n983;
  assign n985 = ~pi56  & pi184 ;
  assign n986 = ~pi57  & pi185 ;
  assign n987 = ~n985 & ~n986;
  assign n988 = n984 & n987;
  assign n989 = n981 & n987;
  assign n990 = n984 & n989;
  assign n991 = n981 & n988;
  assign n992 = ~n974 & n4582;
  assign n993 = pi59  & ~pi187 ;
  assign n994 = pi56  & ~pi184 ;
  assign n995 = ~n986 & n994;
  assign n996 = pi57  & ~pi185 ;
  assign n997 = pi58  & ~pi186 ;
  assign n998 = ~n996 & ~n997;
  assign n999 = ~n995 & ~n996;
  assign n1000 = ~n997 & n999;
  assign n1001 = ~n995 & n998;
  assign n1002 = n984 & ~n4583;
  assign n1003 = ~n993 & ~n1002;
  assign n1004 = n981 & ~n1003;
  assign n1005 = pi63  & ~pi191 ;
  assign n1006 = pi60  & ~pi188 ;
  assign n1007 = ~n978 & n1006;
  assign n1008 = pi62  & ~pi190 ;
  assign n1009 = pi61  & ~pi189 ;
  assign n1010 = ~n1008 & ~n1009;
  assign n1011 = ~n1007 & n1010;
  assign n1012 = n977 & ~n1011;
  assign n1013 = ~n1007 & ~n1009;
  assign n1014 = n977 & ~n1013;
  assign n1015 = ~pi190  & ~n975;
  assign n1016 = pi62  & n1015;
  assign n1017 = ~n975 & n1008;
  assign n1018 = ~n1005 & ~n4584;
  assign n1019 = ~n1014 & n1018;
  assign n1020 = ~n1005 & ~n1012;
  assign n1021 = ~n1004 & n4585;
  assign n1022 = ~n992 & ~n4584;
  assign n1023 = ~n1014 & n1022;
  assign n1024 = ~n1004 & n1023;
  assign n1025 = ~n1005 & n1024;
  assign n1026 = ~n992 & n1021;
  assign n1027 = ~pi67  & pi195 ;
  assign n1028 = ~pi66  & pi194 ;
  assign n1029 = ~n1027 & ~n1028;
  assign n1030 = ~pi65  & pi193 ;
  assign n1031 = ~pi64  & pi192 ;
  assign n1032 = ~n1030 & ~n1031;
  assign n1033 = n1029 & n1032;
  assign n1034 = ~n4586 & ~n1031;
  assign n1035 = ~n1030 & n1034;
  assign n1036 = n1029 & n1035;
  assign n1037 = ~n4586 & n1033;
  assign n1038 = pi67  & ~pi195 ;
  assign n1039 = pi64  & ~pi192 ;
  assign n1040 = ~n1030 & n1039;
  assign n1041 = pi65  & ~pi193 ;
  assign n1042 = pi66  & ~pi194 ;
  assign n1043 = ~n1041 & ~n1042;
  assign n1044 = ~n1040 & ~n1041;
  assign n1045 = ~n1042 & n1044;
  assign n1046 = ~n1040 & n1043;
  assign n1047 = n1029 & ~n4588;
  assign n1048 = ~n1038 & ~n1047;
  assign n1049 = ~n4587 & n1048;
  assign n1050 = ~pi71  & pi199 ;
  assign n1051 = ~pi70  & pi198 ;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = ~pi69  & pi197 ;
  assign n1054 = ~pi68  & pi196 ;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = n1052 & n1055;
  assign n1057 = ~n1049 & n1056;
  assign n1058 = pi71  & ~pi199 ;
  assign n1059 = pi68  & ~pi196 ;
  assign n1060 = ~n1053 & n1059;
  assign n1061 = pi70  & ~pi198 ;
  assign n1062 = pi69  & ~pi197 ;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = ~n1060 & n1063;
  assign n1065 = n1052 & ~n1064;
  assign n1066 = ~n1060 & ~n1062;
  assign n1067 = n1052 & ~n1066;
  assign n1068 = ~pi198  & ~n1050;
  assign n1069 = pi70  & n1068;
  assign n1070 = ~n1050 & n1061;
  assign n1071 = ~n1058 & ~n4589;
  assign n1072 = ~n1067 & n1071;
  assign n1073 = ~n1058 & ~n1065;
  assign n1074 = ~n1057 & ~n4589;
  assign n1075 = ~n1067 & n1074;
  assign n1076 = ~n1058 & n1075;
  assign n1077 = ~n1057 & n4590;
  assign n1078 = ~pi75  & pi203 ;
  assign n1079 = ~pi74  & pi202 ;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = ~pi73  & pi201 ;
  assign n1082 = ~pi72  & pi200 ;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = n1080 & n1083;
  assign n1085 = ~n4591 & n1084;
  assign n1086 = pi75  & ~pi203 ;
  assign n1087 = pi72  & ~pi200 ;
  assign n1088 = ~n1081 & n1087;
  assign n1089 = pi73  & ~pi201 ;
  assign n1090 = pi74  & ~pi202 ;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = ~n1088 & ~n1089;
  assign n1093 = ~n1090 & n1092;
  assign n1094 = ~n1088 & n1091;
  assign n1095 = n1080 & ~n4592;
  assign n1096 = ~n1086 & ~n1095;
  assign n1097 = ~n1085 & n1096;
  assign n1098 = ~pi79  & pi207 ;
  assign n1099 = ~pi78  & pi206 ;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = ~pi77  & pi205 ;
  assign n1102 = ~pi76  & pi204 ;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = n1100 & n1103;
  assign n1105 = ~n1097 & n1104;
  assign n1106 = pi79  & ~pi207 ;
  assign n1107 = pi76  & ~pi204 ;
  assign n1108 = ~n1101 & n1107;
  assign n1109 = pi78  & ~pi206 ;
  assign n1110 = pi77  & ~pi205 ;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = ~n1108 & n1111;
  assign n1113 = n1100 & ~n1112;
  assign n1114 = ~n1108 & ~n1110;
  assign n1115 = n1100 & ~n1114;
  assign n1116 = ~pi206  & ~n1098;
  assign n1117 = pi78  & n1116;
  assign n1118 = ~n1098 & n1109;
  assign n1119 = ~n1106 & ~n4593;
  assign n1120 = ~n1115 & n1119;
  assign n1121 = ~n1106 & ~n1113;
  assign n1122 = ~n1105 & ~n4593;
  assign n1123 = ~n1115 & n1122;
  assign n1124 = ~n1106 & n1123;
  assign n1125 = ~n1105 & n4594;
  assign n1126 = ~pi83  & pi211 ;
  assign n1127 = ~pi82  & pi210 ;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = ~pi81  & pi209 ;
  assign n1130 = ~pi80  & pi208 ;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = n1128 & n1131;
  assign n1133 = ~n4595 & ~n1129;
  assign n1134 = n1128 & n1133;
  assign n1135 = ~n1130 & n1134;
  assign n1136 = ~n4595 & n1132;
  assign n1137 = pi83  & ~pi211 ;
  assign n1138 = pi80  & ~pi208 ;
  assign n1139 = ~pi208  & ~n1129;
  assign n1140 = pi80  & n1139;
  assign n1141 = ~n1129 & n1138;
  assign n1142 = pi81  & ~pi209 ;
  assign n1143 = pi82  & ~pi210 ;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = ~n4597 & ~n1142;
  assign n1146 = ~n1143 & n1145;
  assign n1147 = ~n4597 & n1144;
  assign n1148 = n1128 & ~n4598;
  assign n1149 = ~n1137 & ~n1148;
  assign n1150 = ~n4596 & n1149;
  assign n1151 = ~pi87  & pi215 ;
  assign n1152 = ~pi86  & pi214 ;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~pi85  & pi213 ;
  assign n1155 = ~pi84  & pi212 ;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = n1153 & n1156;
  assign n1158 = ~n1150 & n1157;
  assign n1159 = pi87  & ~pi215 ;
  assign n1160 = pi84  & ~pi212 ;
  assign n1161 = ~n1154 & n1160;
  assign n1162 = pi86  & ~pi214 ;
  assign n1163 = pi85  & ~pi213 ;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = ~n1161 & n1164;
  assign n1166 = n1153 & ~n1165;
  assign n1167 = ~n1161 & ~n1163;
  assign n1168 = n1153 & ~n1167;
  assign n1169 = ~pi214  & ~n1151;
  assign n1170 = pi86  & n1169;
  assign n1171 = ~n1151 & n1162;
  assign n1172 = ~n1159 & ~n4599;
  assign n1173 = ~n1168 & n1172;
  assign n1174 = ~n1159 & ~n1166;
  assign n1175 = ~n1158 & ~n4599;
  assign n1176 = ~n1168 & n1175;
  assign n1177 = ~n1159 & n1176;
  assign n1178 = ~n1158 & n4600;
  assign n1179 = ~pi91  & pi219 ;
  assign n1180 = ~pi90  & pi218 ;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = ~pi89  & pi217 ;
  assign n1183 = ~pi88  & pi216 ;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = n1181 & n1184;
  assign n1186 = ~n4601 & n1185;
  assign n1187 = pi91  & ~pi219 ;
  assign n1188 = pi88  & ~pi216 ;
  assign n1189 = ~n1182 & n1188;
  assign n1190 = pi89  & ~pi217 ;
  assign n1191 = pi90  & ~pi218 ;
  assign n1192 = ~n1190 & ~n1191;
  assign n1193 = ~n1189 & ~n1190;
  assign n1194 = ~n1191 & n1193;
  assign n1195 = ~n1189 & n1192;
  assign n1196 = n1181 & ~n4602;
  assign n1197 = ~n1187 & ~n1196;
  assign n1198 = ~n1186 & n1197;
  assign n1199 = ~pi95  & pi223 ;
  assign n1200 = ~pi94  & pi222 ;
  assign n1201 = ~n1199 & ~n1200;
  assign n1202 = ~pi93  & pi221 ;
  assign n1203 = ~pi92  & pi220 ;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = n1201 & n1204;
  assign n1206 = ~n1198 & n1205;
  assign n1207 = pi95  & ~pi223 ;
  assign n1208 = pi92  & ~pi220 ;
  assign n1209 = ~n1202 & n1208;
  assign n1210 = pi94  & ~pi222 ;
  assign n1211 = pi93  & ~pi221 ;
  assign n1212 = ~n1210 & ~n1211;
  assign n1213 = ~n1209 & n1212;
  assign n1214 = n1201 & ~n1213;
  assign n1215 = ~n1209 & ~n1211;
  assign n1216 = n1201 & ~n1215;
  assign n1217 = ~pi222  & ~n1199;
  assign n1218 = pi94  & n1217;
  assign n1219 = ~n1199 & n1210;
  assign n1220 = ~n1207 & ~n4603;
  assign n1221 = ~n1216 & n1220;
  assign n1222 = ~n1207 & ~n1214;
  assign n1223 = ~n1206 & ~n4603;
  assign n1224 = ~n1216 & n1223;
  assign n1225 = ~n1207 & n1224;
  assign n1226 = ~n1206 & n4604;
  assign n1227 = ~pi99  & pi227 ;
  assign n1228 = ~pi98  & pi226 ;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~pi97  & pi225 ;
  assign n1231 = ~pi96  & pi224 ;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = n1229 & n1232;
  assign n1234 = ~n4605 & ~n1230;
  assign n1235 = n1229 & n1234;
  assign n1236 = ~n1231 & n1235;
  assign n1237 = ~n4605 & n1233;
  assign n1238 = pi99  & ~pi227 ;
  assign n1239 = pi96  & ~pi224 ;
  assign n1240 = ~pi224  & ~n1230;
  assign n1241 = pi96  & n1240;
  assign n1242 = ~n1230 & n1239;
  assign n1243 = pi97  & ~pi225 ;
  assign n1244 = pi98  & ~pi226 ;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = ~n4607 & ~n1243;
  assign n1247 = ~n1244 & n1246;
  assign n1248 = ~n4607 & n1245;
  assign n1249 = n1229 & ~n4608;
  assign n1250 = ~n1238 & ~n1249;
  assign n1251 = ~n4606 & n1250;
  assign n1252 = ~pi103  & pi231 ;
  assign n1253 = ~pi102  & pi230 ;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = ~pi101  & pi229 ;
  assign n1256 = ~pi100  & pi228 ;
  assign n1257 = ~n1255 & ~n1256;
  assign n1258 = n1254 & n1257;
  assign n1259 = ~n1251 & n1258;
  assign n1260 = pi103  & ~pi231 ;
  assign n1261 = pi100  & ~pi228 ;
  assign n1262 = ~n1255 & n1261;
  assign n1263 = pi102  & ~pi230 ;
  assign n1264 = pi101  & ~pi229 ;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = ~n1262 & n1265;
  assign n1267 = n1254 & ~n1266;
  assign n1268 = ~n1262 & ~n1264;
  assign n1269 = n1254 & ~n1268;
  assign n1270 = ~pi230  & ~n1252;
  assign n1271 = pi102  & n1270;
  assign n1272 = ~n1252 & n1263;
  assign n1273 = ~n1260 & ~n4609;
  assign n1274 = ~n1269 & n1273;
  assign n1275 = ~n1260 & ~n1267;
  assign n1276 = ~n1259 & ~n4609;
  assign n1277 = ~n1269 & n1276;
  assign n1278 = ~n1260 & n1277;
  assign n1279 = ~n1259 & n4610;
  assign n1280 = ~pi107  & pi235 ;
  assign n1281 = ~pi106  & pi234 ;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = ~pi105  & pi233 ;
  assign n1284 = ~pi104  & pi232 ;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = n1282 & n1285;
  assign n1287 = ~n4611 & n1286;
  assign n1288 = pi107  & ~pi235 ;
  assign n1289 = pi104  & ~pi232 ;
  assign n1290 = ~n1283 & n1289;
  assign n1291 = pi105  & ~pi233 ;
  assign n1292 = pi106  & ~pi234 ;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = ~n1290 & ~n1291;
  assign n1295 = ~n1292 & n1294;
  assign n1296 = ~n1290 & n1293;
  assign n1297 = n1282 & ~n4612;
  assign n1298 = ~n1288 & ~n1297;
  assign n1299 = ~n1287 & n1298;
  assign n1300 = ~pi111  & pi239 ;
  assign n1301 = ~pi110  & pi238 ;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = ~pi109  & pi237 ;
  assign n1304 = ~pi108  & pi236 ;
  assign n1305 = ~n1303 & ~n1304;
  assign n1306 = n1302 & n1305;
  assign n1307 = ~n1299 & n1306;
  assign n1308 = pi111  & ~pi239 ;
  assign n1309 = pi108  & ~pi236 ;
  assign n1310 = ~n1303 & n1309;
  assign n1311 = pi110  & ~pi238 ;
  assign n1312 = pi109  & ~pi237 ;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = ~n1310 & n1313;
  assign n1315 = n1302 & ~n1314;
  assign n1316 = ~n1310 & ~n1312;
  assign n1317 = n1302 & ~n1316;
  assign n1318 = ~pi238  & ~n1300;
  assign n1319 = pi110  & n1318;
  assign n1320 = ~n1300 & n1311;
  assign n1321 = ~n1308 & ~n4613;
  assign n1322 = ~n1317 & n1321;
  assign n1323 = ~n1308 & ~n1315;
  assign n1324 = ~n1307 & ~n4613;
  assign n1325 = ~n1317 & n1324;
  assign n1326 = ~n1308 & n1325;
  assign n1327 = ~n1307 & n4614;
  assign n1328 = ~pi115  & pi243 ;
  assign n1329 = ~pi114  & pi242 ;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = ~pi113  & pi241 ;
  assign n1332 = ~pi112  & pi240 ;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = n1330 & n1333;
  assign n1335 = ~n4615 & ~n1331;
  assign n1336 = n1330 & n1335;
  assign n1337 = ~n1332 & n1336;
  assign n1338 = ~n4615 & n1334;
  assign n1339 = pi115  & ~pi243 ;
  assign n1340 = pi112  & ~pi240 ;
  assign n1341 = ~pi240  & ~n1331;
  assign n1342 = pi112  & n1341;
  assign n1343 = ~n1331 & n1340;
  assign n1344 = pi113  & ~pi241 ;
  assign n1345 = pi114  & ~pi242 ;
  assign n1346 = ~n1344 & ~n1345;
  assign n1347 = ~n4617 & ~n1344;
  assign n1348 = ~n1345 & n1347;
  assign n1349 = ~n4617 & n1346;
  assign n1350 = n1330 & ~n4618;
  assign n1351 = ~n1339 & ~n1350;
  assign n1352 = ~n4616 & n1351;
  assign n1353 = ~pi119  & pi247 ;
  assign n1354 = ~pi118  & pi246 ;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = ~pi117  & pi245 ;
  assign n1357 = ~pi116  & pi244 ;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = n1355 & n1358;
  assign n1360 = ~n1352 & n1359;
  assign n1361 = pi119  & ~pi247 ;
  assign n1362 = pi116  & ~pi244 ;
  assign n1363 = ~n1356 & n1362;
  assign n1364 = pi118  & ~pi246 ;
  assign n1365 = pi117  & ~pi245 ;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~n1363 & n1366;
  assign n1368 = n1355 & ~n1367;
  assign n1369 = ~n1363 & ~n1365;
  assign n1370 = n1355 & ~n1369;
  assign n1371 = ~pi246  & ~n1353;
  assign n1372 = pi118  & n1371;
  assign n1373 = ~n1353 & n1364;
  assign n1374 = ~n1361 & ~n4619;
  assign n1375 = ~n1370 & n1374;
  assign n1376 = ~n1361 & ~n1368;
  assign n1377 = ~n1360 & ~n4619;
  assign n1378 = ~n1370 & n1377;
  assign n1379 = ~n1361 & n1378;
  assign n1380 = ~n1360 & n4620;
  assign n1381 = ~pi123  & pi251 ;
  assign n1382 = ~pi122  & pi250 ;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = ~pi121  & pi249 ;
  assign n1385 = ~pi120  & pi248 ;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = n1383 & n1386;
  assign n1388 = ~n4621 & n1387;
  assign n1389 = pi123  & ~pi251 ;
  assign n1390 = pi120  & ~pi248 ;
  assign n1391 = ~n1384 & n1390;
  assign n1392 = pi121  & ~pi249 ;
  assign n1393 = pi122  & ~pi250 ;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = ~n1391 & ~n1392;
  assign n1396 = ~n1393 & n1395;
  assign n1397 = ~n1391 & n1394;
  assign n1398 = n1383 & ~n4622;
  assign n1399 = ~n1389 & ~n1398;
  assign n1400 = ~n1388 & n1399;
  assign n1401 = ~pi126  & pi254 ;
  assign n1402 = ~pi125  & pi253 ;
  assign n1403 = ~n1401 & ~n1402;
  assign n1404 = pi127  & ~pi255 ;
  assign n1405 = ~pi124  & pi252 ;
  assign n1406 = ~n1404 & ~n1405;
  assign n1407 = n1403 & ~n1404;
  assign n1408 = ~n1405 & n1407;
  assign n1409 = n1403 & n1406;
  assign n1410 = ~n1400 & n4623;
  assign n1411 = pi124  & ~pi252 ;
  assign n1412 = pi125  & ~pi253 ;
  assign n1413 = ~n1411 & ~n1412;
  assign n1414 = n1403 & ~n1413;
  assign n1415 = pi126  & ~pi254 ;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = ~n1404 & ~n1416;
  assign n1418 = ~pi127  & pi255 ;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = ~n1410 & ~n1417;
  assign n1421 = ~n1418 & n1420;
  assign n1422 = ~n1410 & n1419;
  assign n1423 = pi28  & ~n4624;
  assign n1424 = pi156  & n4624;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = ~pi284  & pi412 ;
  assign n1427 = pi283  & ~pi411 ;
  assign n1428 = ~pi283  & pi411 ;
  assign n1429 = pi282  & ~pi410 ;
  assign n1430 = ~pi282  & pi410 ;
  assign n1431 = pi281  & ~pi409 ;
  assign n1432 = ~pi281  & pi409 ;
  assign n1433 = pi280  & ~pi408 ;
  assign n1434 = ~pi280  & pi408 ;
  assign n1435 = pi279  & ~pi407 ;
  assign n1436 = ~pi279  & pi407 ;
  assign n1437 = pi278  & ~pi406 ;
  assign n1438 = ~pi278  & pi406 ;
  assign n1439 = pi277  & ~pi405 ;
  assign n1440 = ~pi277  & pi405 ;
  assign n1441 = pi276  & ~pi404 ;
  assign n1442 = ~pi276  & pi404 ;
  assign n1443 = pi275  & ~pi403 ;
  assign n1444 = ~pi275  & pi403 ;
  assign n1445 = pi274  & ~pi402 ;
  assign n1446 = ~pi274  & pi402 ;
  assign n1447 = pi273  & ~pi401 ;
  assign n1448 = ~pi273  & pi401 ;
  assign n1449 = pi272  & ~pi400 ;
  assign n1450 = ~pi272  & pi400 ;
  assign n1451 = pi271  & ~pi399 ;
  assign n1452 = ~pi271  & pi399 ;
  assign n1453 = pi270  & ~pi398 ;
  assign n1454 = ~pi270  & pi398 ;
  assign n1455 = pi269  & ~pi397 ;
  assign n1456 = ~pi269  & pi397 ;
  assign n1457 = pi268  & ~pi396 ;
  assign n1458 = ~pi268  & pi396 ;
  assign n1459 = pi267  & ~pi395 ;
  assign n1460 = ~pi267  & pi395 ;
  assign n1461 = pi266  & ~pi394 ;
  assign n1462 = ~pi266  & pi394 ;
  assign n1463 = pi265  & ~pi393 ;
  assign n1464 = ~pi265  & pi393 ;
  assign n1465 = pi264  & ~pi392 ;
  assign n1466 = ~pi264  & pi392 ;
  assign n1467 = pi263  & ~pi391 ;
  assign n1468 = ~pi263  & pi391 ;
  assign n1469 = pi262  & ~pi390 ;
  assign n1470 = ~pi262  & pi390 ;
  assign n1471 = pi261  & ~pi389 ;
  assign n1472 = ~pi261  & pi389 ;
  assign n1473 = pi260  & ~pi388 ;
  assign n1474 = ~pi260  & pi388 ;
  assign n1475 = pi259  & ~pi387 ;
  assign n1476 = ~pi259  & pi387 ;
  assign n1477 = pi258  & ~pi386 ;
  assign n1478 = ~pi258  & pi386 ;
  assign n1479 = pi257  & ~pi385 ;
  assign n1480 = ~pi257  & pi385 ;
  assign n1481 = pi256  & ~pi384 ;
  assign n1482 = ~n1480 & n1481;
  assign n1483 = ~n1479 & ~n1482;
  assign n1484 = pi257  & n1481;
  assign n1485 = pi385  & ~n1484;
  assign n1486 = ~pi257  & ~n1481;
  assign n1487 = ~n1478 & ~n1486;
  assign n1488 = ~n1485 & n1487;
  assign n1489 = ~n1478 & ~n1483;
  assign n1490 = ~n1477 & ~n4625;
  assign n1491 = ~n1476 & ~n1490;
  assign n1492 = ~n1475 & ~n1491;
  assign n1493 = ~n1474 & ~n1492;
  assign n1494 = ~pi260  & n1492;
  assign n1495 = ~pi388  & ~n1494;
  assign n1496 = pi260  & ~n1492;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = ~n1473 & ~n1493;
  assign n1499 = ~n1472 & ~n4626;
  assign n1500 = ~pi261  & n4626;
  assign n1501 = ~pi389  & ~n1500;
  assign n1502 = pi261  & ~n4626;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = ~n1471 & ~n1499;
  assign n1505 = ~n1470 & ~n4627;
  assign n1506 = ~n1469 & ~n1505;
  assign n1507 = ~n1468 & ~n1506;
  assign n1508 = ~n1467 & ~n1507;
  assign n1509 = ~n1466 & ~n1508;
  assign n1510 = ~pi264  & n1508;
  assign n1511 = ~pi392  & ~n1510;
  assign n1512 = pi264  & ~n1508;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = ~n1465 & ~n1509;
  assign n1515 = ~n1464 & ~n4628;
  assign n1516 = ~pi265  & n4628;
  assign n1517 = ~pi393  & ~n1516;
  assign n1518 = pi265  & ~n4628;
  assign n1519 = ~n1517 & ~n1518;
  assign n1520 = ~n1463 & ~n1515;
  assign n1521 = ~n1462 & ~n4629;
  assign n1522 = ~n1461 & ~n1521;
  assign n1523 = ~n1460 & ~n1522;
  assign n1524 = ~n1459 & ~n1523;
  assign n1525 = ~n1458 & ~n1524;
  assign n1526 = ~n1457 & ~n1525;
  assign n1527 = ~n1456 & ~n1526;
  assign n1528 = ~n1455 & ~n1527;
  assign n1529 = ~n1454 & ~n1528;
  assign n1530 = ~n1453 & ~n1529;
  assign n1531 = ~n1452 & ~n1530;
  assign n1532 = ~n1451 & ~n1531;
  assign n1533 = ~n1450 & ~n1532;
  assign n1534 = ~pi272  & n1532;
  assign n1535 = ~pi400  & ~n1534;
  assign n1536 = pi272  & ~n1532;
  assign n1537 = ~n1535 & ~n1536;
  assign n1538 = ~n1449 & ~n1533;
  assign n1539 = ~n1448 & ~n4630;
  assign n1540 = ~pi273  & n4630;
  assign n1541 = ~pi401  & ~n1540;
  assign n1542 = pi273  & ~n4630;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = ~n1447 & ~n1539;
  assign n1545 = ~n1446 & ~n4631;
  assign n1546 = ~n1445 & ~n1545;
  assign n1547 = ~n1444 & ~n1546;
  assign n1548 = ~n1443 & ~n1547;
  assign n1549 = ~n1442 & ~n1548;
  assign n1550 = ~n1441 & ~n1549;
  assign n1551 = ~n1440 & ~n1550;
  assign n1552 = ~n1439 & ~n1551;
  assign n1553 = ~n1438 & ~n1552;
  assign n1554 = ~n1437 & ~n1553;
  assign n1555 = ~n1436 & ~n1554;
  assign n1556 = ~n1435 & ~n1555;
  assign n1557 = ~n1434 & ~n1556;
  assign n1558 = ~pi280  & n1556;
  assign n1559 = ~pi408  & ~n1558;
  assign n1560 = pi280  & ~n1556;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = ~n1433 & ~n1557;
  assign n1563 = ~n1432 & ~n4632;
  assign n1564 = ~pi281  & n4632;
  assign n1565 = ~pi409  & ~n1564;
  assign n1566 = pi281  & ~n4632;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = ~n1431 & ~n1563;
  assign n1569 = ~n1430 & ~n4633;
  assign n1570 = ~n1429 & ~n1569;
  assign n1571 = ~n1428 & ~n1570;
  assign n1572 = ~n1427 & ~n1571;
  assign n1573 = ~n1426 & ~n1572;
  assign n1574 = pi284  & ~pi412 ;
  assign n1575 = pi285  & ~pi413 ;
  assign n1576 = ~n1574 & ~n1575;
  assign n1577 = ~n1573 & n1576;
  assign n1578 = ~pi285  & pi413 ;
  assign n1579 = ~pi286  & pi414 ;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = ~n1573 & ~n1574;
  assign n1582 = ~n1578 & ~n1581;
  assign n1583 = ~n1575 & ~n1582;
  assign n1584 = ~n1579 & ~n1583;
  assign n1585 = ~n1577 & n1580;
  assign n1586 = pi286  & ~pi414 ;
  assign n1587 = pi287  & ~pi415 ;
  assign n1588 = ~n1586 & ~n1587;
  assign n1589 = ~n4634 & n1588;
  assign n1590 = ~pi295  & pi423 ;
  assign n1591 = ~pi294  & pi422 ;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = ~pi293  & pi421 ;
  assign n1594 = ~pi292  & pi420 ;
  assign n1595 = ~n1593 & ~n1594;
  assign n1596 = n1592 & n1595;
  assign n1597 = ~pi291  & pi419 ;
  assign n1598 = ~pi290  & pi418 ;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = ~pi289  & pi417 ;
  assign n1601 = ~pi288  & pi416 ;
  assign n1602 = ~pi287  & pi415 ;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = ~n1600 & ~n1602;
  assign n1605 = ~n1601 & n1604;
  assign n1606 = ~n1600 & n1603;
  assign n1607 = n1599 & n4635;
  assign n1608 = n1596 & n1607;
  assign n1609 = ~n4634 & ~n1586;
  assign n1610 = ~n1602 & ~n1609;
  assign n1611 = ~n1587 & ~n1610;
  assign n1612 = n1599 & ~n1600;
  assign n1613 = n1596 & n1612;
  assign n1614 = ~n1611 & n1613;
  assign n1615 = ~n1601 & n1614;
  assign n1616 = ~n1589 & n1608;
  assign n1617 = pi291  & ~pi419 ;
  assign n1618 = pi288  & ~pi416 ;
  assign n1619 = ~pi416  & ~n1600;
  assign n1620 = pi288  & n1619;
  assign n1621 = ~n1600 & n1618;
  assign n1622 = pi289  & ~pi417 ;
  assign n1623 = pi290  & ~pi418 ;
  assign n1624 = ~n1622 & ~n1623;
  assign n1625 = ~n4637 & ~n1622;
  assign n1626 = ~n1623 & n1625;
  assign n1627 = ~n4637 & n1624;
  assign n1628 = n1599 & ~n4638;
  assign n1629 = ~n1617 & ~n1628;
  assign n1630 = n1596 & ~n1629;
  assign n1631 = pi295  & ~pi423 ;
  assign n1632 = pi292  & ~pi420 ;
  assign n1633 = ~n1593 & n1632;
  assign n1634 = pi294  & ~pi422 ;
  assign n1635 = pi293  & ~pi421 ;
  assign n1636 = ~n1634 & ~n1635;
  assign n1637 = ~n1633 & n1636;
  assign n1638 = n1592 & ~n1637;
  assign n1639 = ~n1633 & ~n1635;
  assign n1640 = n1592 & ~n1639;
  assign n1641 = ~pi422  & ~n1590;
  assign n1642 = pi294  & n1641;
  assign n1643 = ~n1590 & n1634;
  assign n1644 = ~n1631 & ~n4639;
  assign n1645 = ~n1640 & n1644;
  assign n1646 = ~n1631 & ~n1638;
  assign n1647 = ~n1630 & ~n4639;
  assign n1648 = ~n1640 & n1647;
  assign n1649 = ~n1631 & n1648;
  assign n1650 = ~n1630 & n4640;
  assign n1651 = ~n4636 & n4641;
  assign n1652 = ~pi303  & pi431 ;
  assign n1653 = ~pi302  & pi430 ;
  assign n1654 = ~n1652 & ~n1653;
  assign n1655 = ~pi301  & pi429 ;
  assign n1656 = ~pi300  & pi428 ;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = n1654 & n1657;
  assign n1659 = ~pi299  & pi427 ;
  assign n1660 = ~pi298  & pi426 ;
  assign n1661 = ~n1659 & ~n1660;
  assign n1662 = ~pi296  & pi424 ;
  assign n1663 = ~pi297  & pi425 ;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = n1661 & n1664;
  assign n1666 = n1658 & n1665;
  assign n1667 = ~n1651 & n1666;
  assign n1668 = pi299  & ~pi427 ;
  assign n1669 = pi296  & ~pi424 ;
  assign n1670 = ~n1663 & n1669;
  assign n1671 = pi297  & ~pi425 ;
  assign n1672 = pi298  & ~pi426 ;
  assign n1673 = ~n1671 & ~n1672;
  assign n1674 = ~n1670 & ~n1671;
  assign n1675 = ~n1672 & n1674;
  assign n1676 = ~n1670 & n1673;
  assign n1677 = n1661 & ~n4642;
  assign n1678 = ~n1668 & ~n1677;
  assign n1679 = n1658 & ~n1678;
  assign n1680 = pi303  & ~pi431 ;
  assign n1681 = pi300  & ~pi428 ;
  assign n1682 = ~n1655 & n1681;
  assign n1683 = pi302  & ~pi430 ;
  assign n1684 = pi301  & ~pi429 ;
  assign n1685 = ~n1683 & ~n1684;
  assign n1686 = ~n1682 & n1685;
  assign n1687 = n1654 & ~n1686;
  assign n1688 = ~n1682 & ~n1684;
  assign n1689 = n1654 & ~n1688;
  assign n1690 = ~pi430  & ~n1652;
  assign n1691 = pi302  & n1690;
  assign n1692 = ~n1652 & n1683;
  assign n1693 = ~n1680 & ~n4643;
  assign n1694 = ~n1689 & n1693;
  assign n1695 = ~n1680 & ~n1687;
  assign n1696 = ~n1679 & n4644;
  assign n1697 = ~n1667 & ~n4643;
  assign n1698 = ~n1689 & n1697;
  assign n1699 = ~n1679 & n1698;
  assign n1700 = ~n1680 & n1699;
  assign n1701 = ~n1667 & n1696;
  assign n1702 = ~pi309  & pi437 ;
  assign n1703 = ~pi308  & pi436 ;
  assign n1704 = ~pi436  & ~n1702;
  assign n1705 = pi308  & ~n1702;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = ~n1702 & ~n1703;
  assign n1708 = ~pi311  & pi439 ;
  assign n1709 = ~pi310  & pi438 ;
  assign n1710 = ~n1708 & ~n1709;
  assign n1711 = ~n4646 & n1710;
  assign n1712 = ~pi307  & pi435 ;
  assign n1713 = ~pi306  & pi434 ;
  assign n1714 = ~n1712 & ~n1713;
  assign n1715 = ~pi304  & pi432 ;
  assign n1716 = ~pi305  & pi433 ;
  assign n1717 = ~n1715 & ~n1716;
  assign n1718 = n1714 & n1717;
  assign n1719 = n1710 & n1717;
  assign n1720 = n1714 & n1719;
  assign n1721 = ~n4646 & n1720;
  assign n1722 = n1714 & ~n1716;
  assign n1723 = n1711 & n1722;
  assign n1724 = ~n1715 & n1723;
  assign n1725 = n1711 & n1718;
  assign n1726 = ~n4645 & n4647;
  assign n1727 = pi307  & ~pi435 ;
  assign n1728 = pi304  & ~pi432 ;
  assign n1729 = ~pi432  & ~n1716;
  assign n1730 = pi304  & n1729;
  assign n1731 = ~n1716 & n1728;
  assign n1732 = pi305  & ~pi433 ;
  assign n1733 = pi306  & ~pi434 ;
  assign n1734 = ~n1732 & ~n1733;
  assign n1735 = ~n4648 & ~n1732;
  assign n1736 = ~n1733 & n1735;
  assign n1737 = ~n4648 & n1734;
  assign n1738 = n1714 & ~n4649;
  assign n1739 = ~n1727 & ~n1738;
  assign n1740 = n1711 & ~n1739;
  assign n1741 = pi311  & ~pi439 ;
  assign n1742 = pi308  & ~pi436 ;
  assign n1743 = pi308  & n1704;
  assign n1744 = ~n1702 & n1742;
  assign n1745 = pi309  & ~pi437 ;
  assign n1746 = pi310  & ~pi438 ;
  assign n1747 = ~n1745 & ~n1746;
  assign n1748 = ~n4650 & ~n1745;
  assign n1749 = ~n1746 & n1748;
  assign n1750 = ~n4650 & n1747;
  assign n1751 = n1710 & ~n4651;
  assign n1752 = ~n1741 & ~n1751;
  assign n1753 = ~n4646 & ~n1739;
  assign n1754 = n4651 & ~n1753;
  assign n1755 = n1710 & ~n1754;
  assign n1756 = ~n1740 & ~n1751;
  assign n1757 = ~n1741 & ~n4652;
  assign n1758 = ~n1740 & n1752;
  assign n1759 = ~n1726 & n4653;
  assign n1760 = ~pi319  & pi447 ;
  assign n1761 = ~pi318  & pi446 ;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = ~pi317  & pi445 ;
  assign n1764 = ~pi316  & pi444 ;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = n1762 & n1765;
  assign n1767 = ~pi315  & pi443 ;
  assign n1768 = ~pi314  & pi442 ;
  assign n1769 = ~n1767 & ~n1768;
  assign n1770 = ~pi312  & pi440 ;
  assign n1771 = ~pi313  & pi441 ;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = n1769 & n1772;
  assign n1774 = n1766 & n1772;
  assign n1775 = n1769 & n1774;
  assign n1776 = n1766 & n1773;
  assign n1777 = ~n1759 & n4654;
  assign n1778 = pi315  & ~pi443 ;
  assign n1779 = pi312  & ~pi440 ;
  assign n1780 = ~n1771 & n1779;
  assign n1781 = pi313  & ~pi441 ;
  assign n1782 = pi314  & ~pi442 ;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = ~n1780 & ~n1781;
  assign n1785 = ~n1782 & n1784;
  assign n1786 = ~n1780 & n1783;
  assign n1787 = n1769 & ~n4655;
  assign n1788 = ~n1778 & ~n1787;
  assign n1789 = n1766 & ~n1788;
  assign n1790 = pi319  & ~pi447 ;
  assign n1791 = pi316  & ~pi444 ;
  assign n1792 = ~n1763 & n1791;
  assign n1793 = pi318  & ~pi446 ;
  assign n1794 = pi317  & ~pi445 ;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = ~n1792 & n1795;
  assign n1797 = n1762 & ~n1796;
  assign n1798 = ~n1792 & ~n1794;
  assign n1799 = n1762 & ~n1798;
  assign n1800 = ~pi446  & ~n1760;
  assign n1801 = pi318  & n1800;
  assign n1802 = ~n1760 & n1793;
  assign n1803 = ~n1790 & ~n4656;
  assign n1804 = ~n1799 & n1803;
  assign n1805 = ~n1790 & ~n1797;
  assign n1806 = ~n1789 & n4657;
  assign n1807 = ~n1777 & ~n4656;
  assign n1808 = ~n1799 & n1807;
  assign n1809 = ~n1789 & n1808;
  assign n1810 = ~n1790 & n1809;
  assign n1811 = ~n1777 & n1806;
  assign n1812 = ~pi323  & pi451 ;
  assign n1813 = ~pi322  & pi450 ;
  assign n1814 = ~n1812 & ~n1813;
  assign n1815 = ~pi321  & pi449 ;
  assign n1816 = ~pi320  & pi448 ;
  assign n1817 = ~n1815 & ~n1816;
  assign n1818 = n1814 & n1817;
  assign n1819 = ~n4658 & ~n1816;
  assign n1820 = ~n1815 & n1819;
  assign n1821 = n1814 & n1820;
  assign n1822 = ~n4658 & n1818;
  assign n1823 = pi323  & ~pi451 ;
  assign n1824 = pi320  & ~pi448 ;
  assign n1825 = ~n1815 & n1824;
  assign n1826 = pi321  & ~pi449 ;
  assign n1827 = pi322  & ~pi450 ;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = ~n1825 & ~n1826;
  assign n1830 = ~n1827 & n1829;
  assign n1831 = ~n1825 & n1828;
  assign n1832 = n1814 & ~n4660;
  assign n1833 = ~n1823 & ~n1832;
  assign n1834 = ~n4659 & n1833;
  assign n1835 = ~pi327  & pi455 ;
  assign n1836 = ~pi326  & pi454 ;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = ~pi325  & pi453 ;
  assign n1839 = ~pi324  & pi452 ;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = n1837 & n1840;
  assign n1842 = ~n1834 & n1841;
  assign n1843 = pi327  & ~pi455 ;
  assign n1844 = pi324  & ~pi452 ;
  assign n1845 = ~n1838 & n1844;
  assign n1846 = pi326  & ~pi454 ;
  assign n1847 = pi325  & ~pi453 ;
  assign n1848 = ~n1846 & ~n1847;
  assign n1849 = ~n1845 & n1848;
  assign n1850 = n1837 & ~n1849;
  assign n1851 = ~n1845 & ~n1847;
  assign n1852 = n1837 & ~n1851;
  assign n1853 = ~pi454  & ~n1835;
  assign n1854 = pi326  & n1853;
  assign n1855 = ~n1835 & n1846;
  assign n1856 = ~n1843 & ~n4661;
  assign n1857 = ~n1852 & n1856;
  assign n1858 = ~n1843 & ~n1850;
  assign n1859 = ~n1842 & ~n4661;
  assign n1860 = ~n1852 & n1859;
  assign n1861 = ~n1843 & n1860;
  assign n1862 = ~n1842 & n4662;
  assign n1863 = ~pi331  & pi459 ;
  assign n1864 = ~pi330  & pi458 ;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = ~pi329  & pi457 ;
  assign n1867 = ~pi328  & pi456 ;
  assign n1868 = ~n1866 & ~n1867;
  assign n1869 = n1865 & n1868;
  assign n1870 = ~n4663 & n1869;
  assign n1871 = pi331  & ~pi459 ;
  assign n1872 = pi328  & ~pi456 ;
  assign n1873 = ~n1866 & n1872;
  assign n1874 = pi329  & ~pi457 ;
  assign n1875 = pi330  & ~pi458 ;
  assign n1876 = ~n1874 & ~n1875;
  assign n1877 = ~n1873 & ~n1874;
  assign n1878 = ~n1875 & n1877;
  assign n1879 = ~n1873 & n1876;
  assign n1880 = n1865 & ~n4664;
  assign n1881 = ~n1871 & ~n1880;
  assign n1882 = ~n1870 & n1881;
  assign n1883 = ~pi335  & pi463 ;
  assign n1884 = ~pi334  & pi462 ;
  assign n1885 = ~n1883 & ~n1884;
  assign n1886 = ~pi333  & pi461 ;
  assign n1887 = ~pi332  & pi460 ;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = n1885 & n1888;
  assign n1890 = ~n1882 & n1889;
  assign n1891 = pi335  & ~pi463 ;
  assign n1892 = pi332  & ~pi460 ;
  assign n1893 = ~n1886 & n1892;
  assign n1894 = pi334  & ~pi462 ;
  assign n1895 = pi333  & ~pi461 ;
  assign n1896 = ~n1894 & ~n1895;
  assign n1897 = ~n1893 & n1896;
  assign n1898 = n1885 & ~n1897;
  assign n1899 = ~n1893 & ~n1895;
  assign n1900 = n1885 & ~n1899;
  assign n1901 = ~pi462  & ~n1883;
  assign n1902 = pi334  & n1901;
  assign n1903 = ~n1883 & n1894;
  assign n1904 = ~n1891 & ~n4665;
  assign n1905 = ~n1900 & n1904;
  assign n1906 = ~n1891 & ~n1898;
  assign n1907 = ~n1890 & ~n4665;
  assign n1908 = ~n1900 & n1907;
  assign n1909 = ~n1891 & n1908;
  assign n1910 = ~n1890 & n4666;
  assign n1911 = ~pi339  & pi467 ;
  assign n1912 = ~pi338  & pi466 ;
  assign n1913 = ~n1911 & ~n1912;
  assign n1914 = ~pi337  & pi465 ;
  assign n1915 = ~pi336  & pi464 ;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = n1913 & n1916;
  assign n1918 = ~n4667 & ~n1914;
  assign n1919 = n1913 & n1918;
  assign n1920 = ~n1915 & n1919;
  assign n1921 = ~n4667 & n1917;
  assign n1922 = pi339  & ~pi467 ;
  assign n1923 = pi336  & ~pi464 ;
  assign n1924 = ~pi464  & ~n1914;
  assign n1925 = pi336  & n1924;
  assign n1926 = ~n1914 & n1923;
  assign n1927 = pi337  & ~pi465 ;
  assign n1928 = pi338  & ~pi466 ;
  assign n1929 = ~n1927 & ~n1928;
  assign n1930 = ~n4669 & ~n1927;
  assign n1931 = ~n1928 & n1930;
  assign n1932 = ~n4669 & n1929;
  assign n1933 = n1913 & ~n4670;
  assign n1934 = ~n1922 & ~n1933;
  assign n1935 = ~n4668 & n1934;
  assign n1936 = ~pi343  & pi471 ;
  assign n1937 = ~pi342  & pi470 ;
  assign n1938 = ~n1936 & ~n1937;
  assign n1939 = ~pi341  & pi469 ;
  assign n1940 = ~pi340  & pi468 ;
  assign n1941 = ~n1939 & ~n1940;
  assign n1942 = n1938 & n1941;
  assign n1943 = ~n1935 & n1942;
  assign n1944 = pi343  & ~pi471 ;
  assign n1945 = pi340  & ~pi468 ;
  assign n1946 = ~n1939 & n1945;
  assign n1947 = pi342  & ~pi470 ;
  assign n1948 = pi341  & ~pi469 ;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = ~n1946 & n1949;
  assign n1951 = n1938 & ~n1950;
  assign n1952 = ~n1946 & ~n1948;
  assign n1953 = n1938 & ~n1952;
  assign n1954 = ~pi470  & ~n1936;
  assign n1955 = pi342  & n1954;
  assign n1956 = ~n1936 & n1947;
  assign n1957 = ~n1944 & ~n4671;
  assign n1958 = ~n1953 & n1957;
  assign n1959 = ~n1944 & ~n1951;
  assign n1960 = ~n1943 & ~n4671;
  assign n1961 = ~n1953 & n1960;
  assign n1962 = ~n1944 & n1961;
  assign n1963 = ~n1943 & n4672;
  assign n1964 = ~pi347  & pi475 ;
  assign n1965 = ~pi346  & pi474 ;
  assign n1966 = ~n1964 & ~n1965;
  assign n1967 = ~pi345  & pi473 ;
  assign n1968 = ~pi344  & pi472 ;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = n1966 & n1969;
  assign n1971 = ~n4673 & n1970;
  assign n1972 = pi347  & ~pi475 ;
  assign n1973 = pi344  & ~pi472 ;
  assign n1974 = ~n1967 & n1973;
  assign n1975 = pi345  & ~pi473 ;
  assign n1976 = pi346  & ~pi474 ;
  assign n1977 = ~n1975 & ~n1976;
  assign n1978 = ~n1974 & ~n1975;
  assign n1979 = ~n1976 & n1978;
  assign n1980 = ~n1974 & n1977;
  assign n1981 = n1966 & ~n4674;
  assign n1982 = ~n1972 & ~n1981;
  assign n1983 = ~n1971 & n1982;
  assign n1984 = ~pi351  & pi479 ;
  assign n1985 = ~pi350  & pi478 ;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = ~pi349  & pi477 ;
  assign n1988 = ~pi348  & pi476 ;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = n1986 & n1989;
  assign n1991 = ~n1983 & n1990;
  assign n1992 = pi351  & ~pi479 ;
  assign n1993 = pi348  & ~pi476 ;
  assign n1994 = ~n1987 & n1993;
  assign n1995 = pi350  & ~pi478 ;
  assign n1996 = pi349  & ~pi477 ;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = ~n1994 & n1997;
  assign n1999 = n1986 & ~n1998;
  assign n2000 = ~n1994 & ~n1996;
  assign n2001 = n1986 & ~n2000;
  assign n2002 = ~pi478  & ~n1984;
  assign n2003 = pi350  & n2002;
  assign n2004 = ~n1984 & n1995;
  assign n2005 = ~n1992 & ~n4675;
  assign n2006 = ~n2001 & n2005;
  assign n2007 = ~n1992 & ~n1999;
  assign n2008 = ~n1991 & ~n4675;
  assign n2009 = ~n2001 & n2008;
  assign n2010 = ~n1992 & n2009;
  assign n2011 = ~n1991 & n4676;
  assign n2012 = ~pi355  & pi483 ;
  assign n2013 = ~pi354  & pi482 ;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = ~pi353  & pi481 ;
  assign n2016 = ~pi352  & pi480 ;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = n2014 & n2017;
  assign n2019 = ~n4677 & ~n2015;
  assign n2020 = n2014 & n2019;
  assign n2021 = ~n2016 & n2020;
  assign n2022 = ~n4677 & n2018;
  assign n2023 = pi355  & ~pi483 ;
  assign n2024 = pi352  & ~pi480 ;
  assign n2025 = ~pi480  & ~n2015;
  assign n2026 = pi352  & n2025;
  assign n2027 = ~n2015 & n2024;
  assign n2028 = pi353  & ~pi481 ;
  assign n2029 = pi354  & ~pi482 ;
  assign n2030 = ~n2028 & ~n2029;
  assign n2031 = ~n4679 & ~n2028;
  assign n2032 = ~n2029 & n2031;
  assign n2033 = ~n4679 & n2030;
  assign n2034 = n2014 & ~n4680;
  assign n2035 = ~n2023 & ~n2034;
  assign n2036 = ~n4678 & n2035;
  assign n2037 = ~pi359  & pi487 ;
  assign n2038 = ~pi358  & pi486 ;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = ~pi357  & pi485 ;
  assign n2041 = ~pi356  & pi484 ;
  assign n2042 = ~n2040 & ~n2041;
  assign n2043 = n2039 & n2042;
  assign n2044 = ~n2036 & n2043;
  assign n2045 = pi359  & ~pi487 ;
  assign n2046 = pi356  & ~pi484 ;
  assign n2047 = ~n2040 & n2046;
  assign n2048 = pi358  & ~pi486 ;
  assign n2049 = pi357  & ~pi485 ;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = ~n2047 & n2050;
  assign n2052 = n2039 & ~n2051;
  assign n2053 = ~n2047 & ~n2049;
  assign n2054 = n2039 & ~n2053;
  assign n2055 = ~pi486  & ~n2037;
  assign n2056 = pi358  & n2055;
  assign n2057 = ~n2037 & n2048;
  assign n2058 = ~n2045 & ~n4681;
  assign n2059 = ~n2054 & n2058;
  assign n2060 = ~n2045 & ~n2052;
  assign n2061 = ~n2044 & ~n4681;
  assign n2062 = ~n2054 & n2061;
  assign n2063 = ~n2045 & n2062;
  assign n2064 = ~n2044 & n4682;
  assign n2065 = ~pi363  & pi491 ;
  assign n2066 = ~pi362  & pi490 ;
  assign n2067 = ~n2065 & ~n2066;
  assign n2068 = ~pi361  & pi489 ;
  assign n2069 = ~pi360  & pi488 ;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = n2067 & n2070;
  assign n2072 = ~n4683 & n2071;
  assign n2073 = pi363  & ~pi491 ;
  assign n2074 = pi360  & ~pi488 ;
  assign n2075 = ~n2068 & n2074;
  assign n2076 = pi361  & ~pi489 ;
  assign n2077 = pi362  & ~pi490 ;
  assign n2078 = ~n2076 & ~n2077;
  assign n2079 = ~n2075 & ~n2076;
  assign n2080 = ~n2077 & n2079;
  assign n2081 = ~n2075 & n2078;
  assign n2082 = n2067 & ~n4684;
  assign n2083 = ~n2073 & ~n2082;
  assign n2084 = ~n2072 & n2083;
  assign n2085 = ~pi367  & pi495 ;
  assign n2086 = ~pi366  & pi494 ;
  assign n2087 = ~n2085 & ~n2086;
  assign n2088 = ~pi365  & pi493 ;
  assign n2089 = ~pi364  & pi492 ;
  assign n2090 = ~n2088 & ~n2089;
  assign n2091 = n2087 & n2090;
  assign n2092 = ~n2084 & n2091;
  assign n2093 = pi367  & ~pi495 ;
  assign n2094 = pi364  & ~pi492 ;
  assign n2095 = ~n2088 & n2094;
  assign n2096 = pi366  & ~pi494 ;
  assign n2097 = pi365  & ~pi493 ;
  assign n2098 = ~n2096 & ~n2097;
  assign n2099 = ~n2095 & n2098;
  assign n2100 = n2087 & ~n2099;
  assign n2101 = ~n2095 & ~n2097;
  assign n2102 = n2087 & ~n2101;
  assign n2103 = ~pi494  & ~n2085;
  assign n2104 = pi366  & n2103;
  assign n2105 = ~n2085 & n2096;
  assign n2106 = ~n2093 & ~n4685;
  assign n2107 = ~n2102 & n2106;
  assign n2108 = ~n2093 & ~n2100;
  assign n2109 = ~n2092 & ~n4685;
  assign n2110 = ~n2102 & n2109;
  assign n2111 = ~n2093 & n2110;
  assign n2112 = ~n2092 & n4686;
  assign n2113 = ~pi371  & pi499 ;
  assign n2114 = ~pi370  & pi498 ;
  assign n2115 = ~n2113 & ~n2114;
  assign n2116 = ~pi369  & pi497 ;
  assign n2117 = ~pi368  & pi496 ;
  assign n2118 = ~n2116 & ~n2117;
  assign n2119 = n2115 & n2118;
  assign n2120 = ~n4687 & ~n2116;
  assign n2121 = n2115 & n2120;
  assign n2122 = ~n2117 & n2121;
  assign n2123 = ~n4687 & n2119;
  assign n2124 = pi371  & ~pi499 ;
  assign n2125 = pi368  & ~pi496 ;
  assign n2126 = ~pi496  & ~n2116;
  assign n2127 = pi368  & n2126;
  assign n2128 = ~n2116 & n2125;
  assign n2129 = pi369  & ~pi497 ;
  assign n2130 = pi370  & ~pi498 ;
  assign n2131 = ~n2129 & ~n2130;
  assign n2132 = ~n4689 & ~n2129;
  assign n2133 = ~n2130 & n2132;
  assign n2134 = ~n4689 & n2131;
  assign n2135 = n2115 & ~n4690;
  assign n2136 = ~n2124 & ~n2135;
  assign n2137 = ~n4688 & n2136;
  assign n2138 = ~pi375  & pi503 ;
  assign n2139 = ~pi374  & pi502 ;
  assign n2140 = ~n2138 & ~n2139;
  assign n2141 = ~pi373  & pi501 ;
  assign n2142 = ~pi372  & pi500 ;
  assign n2143 = ~n2141 & ~n2142;
  assign n2144 = n2140 & n2143;
  assign n2145 = ~n2137 & n2144;
  assign n2146 = pi375  & ~pi503 ;
  assign n2147 = pi372  & ~pi500 ;
  assign n2148 = ~n2141 & n2147;
  assign n2149 = pi374  & ~pi502 ;
  assign n2150 = pi373  & ~pi501 ;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = ~n2148 & n2151;
  assign n2153 = n2140 & ~n2152;
  assign n2154 = ~n2148 & ~n2150;
  assign n2155 = n2140 & ~n2154;
  assign n2156 = ~pi502  & ~n2138;
  assign n2157 = pi374  & n2156;
  assign n2158 = ~n2138 & n2149;
  assign n2159 = ~n2146 & ~n4691;
  assign n2160 = ~n2155 & n2159;
  assign n2161 = ~n2146 & ~n2153;
  assign n2162 = ~n2145 & ~n4691;
  assign n2163 = ~n2155 & n2162;
  assign n2164 = ~n2146 & n2163;
  assign n2165 = ~n2145 & n4692;
  assign n2166 = ~pi379  & pi507 ;
  assign n2167 = ~pi378  & pi506 ;
  assign n2168 = ~n2166 & ~n2167;
  assign n2169 = ~pi377  & pi505 ;
  assign n2170 = ~pi376  & pi504 ;
  assign n2171 = ~n2169 & ~n2170;
  assign n2172 = n2168 & n2171;
  assign n2173 = ~n4693 & n2172;
  assign n2174 = pi379  & ~pi507 ;
  assign n2175 = pi376  & ~pi504 ;
  assign n2176 = ~n2169 & n2175;
  assign n2177 = pi377  & ~pi505 ;
  assign n2178 = pi378  & ~pi506 ;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = ~n2176 & ~n2177;
  assign n2181 = ~n2178 & n2180;
  assign n2182 = ~n2176 & n2179;
  assign n2183 = n2168 & ~n4694;
  assign n2184 = ~n2174 & ~n2183;
  assign n2185 = ~n2173 & n2184;
  assign n2186 = ~pi382  & pi510 ;
  assign n2187 = ~pi381  & pi509 ;
  assign n2188 = ~n2186 & ~n2187;
  assign n2189 = pi383  & ~pi511 ;
  assign n2190 = ~pi380  & pi508 ;
  assign n2191 = ~n2189 & ~n2190;
  assign n2192 = n2188 & ~n2189;
  assign n2193 = ~n2190 & n2192;
  assign n2194 = n2188 & n2191;
  assign n2195 = ~n2185 & n4695;
  assign n2196 = pi380  & ~pi508 ;
  assign n2197 = pi381  & ~pi509 ;
  assign n2198 = ~n2196 & ~n2197;
  assign n2199 = n2188 & ~n2198;
  assign n2200 = pi382  & ~pi510 ;
  assign n2201 = ~n2199 & ~n2200;
  assign n2202 = ~n2189 & ~n2201;
  assign n2203 = ~pi383  & pi511 ;
  assign n2204 = ~n2202 & ~n2203;
  assign n2205 = ~n2195 & ~n2202;
  assign n2206 = ~n2203 & n2205;
  assign n2207 = ~n2195 & n2204;
  assign n2208 = pi284  & ~n4696;
  assign n2209 = pi412  & n4696;
  assign n2210 = ~n2208 & ~n2209;
  assign n2211 = n1425 & ~n2210;
  assign n2212 = pi27  & ~n4624;
  assign n2213 = pi155  & n4624;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = pi283  & ~n4696;
  assign n2216 = pi411  & n4696;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = ~n2214 & n2217;
  assign n2219 = n2214 & ~n2217;
  assign n2220 = pi26  & ~n4624;
  assign n2221 = pi154  & n4624;
  assign n2222 = ~n2220 & ~n2221;
  assign n2223 = pi282  & ~n4696;
  assign n2224 = pi410  & n4696;
  assign n2225 = ~n2223 & ~n2224;
  assign n2226 = ~n2222 & n2225;
  assign n2227 = n2222 & ~n2225;
  assign n2228 = pi25  & ~n4624;
  assign n2229 = pi153  & n4624;
  assign n2230 = ~n2228 & ~n2229;
  assign n2231 = pi281  & ~n4696;
  assign n2232 = pi409  & n4696;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = ~n2230 & n2233;
  assign n2235 = pi21  & ~n4624;
  assign n2236 = pi149  & n4624;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = pi277  & ~n4696;
  assign n2239 = pi405  & n4696;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = n2237 & ~n2240;
  assign n2242 = pi20  & ~n4624;
  assign n2243 = pi148  & n4624;
  assign n2244 = ~n2242 & ~n2243;
  assign n2245 = pi276  & ~n4696;
  assign n2246 = pi404  & n4696;
  assign n2247 = ~n2245 & ~n2246;
  assign n2248 = ~n2244 & n2247;
  assign n2249 = n2244 & ~n2247;
  assign n2250 = pi19  & ~n4624;
  assign n2251 = pi147  & n4624;
  assign n2252 = ~n2250 & ~n2251;
  assign n2253 = pi275  & ~n4696;
  assign n2254 = pi403  & n4696;
  assign n2255 = ~n2253 & ~n2254;
  assign n2256 = ~n2252 & n2255;
  assign n2257 = n2252 & ~n2255;
  assign n2258 = pi18  & ~n4624;
  assign n2259 = pi146  & n4624;
  assign n2260 = ~n2258 & ~n2259;
  assign n2261 = pi274  & ~n4696;
  assign n2262 = pi402  & n4696;
  assign n2263 = ~n2261 & ~n2262;
  assign n2264 = ~n2260 & n2263;
  assign n2265 = n2260 & ~n2263;
  assign n2266 = pi17  & ~n4624;
  assign n2267 = pi145  & n4624;
  assign n2268 = ~n2266 & ~n2267;
  assign n2269 = pi273  & ~n4696;
  assign n2270 = pi401  & n4696;
  assign n2271 = ~n2269 & ~n2270;
  assign n2272 = ~n2268 & n2271;
  assign n2273 = pi13  & ~n4624;
  assign n2274 = pi141  & n4624;
  assign n2275 = ~n2273 & ~n2274;
  assign n2276 = pi269  & ~n4696;
  assign n2277 = pi397  & n4696;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = n2275 & ~n2278;
  assign n2280 = pi12  & ~n4624;
  assign n2281 = pi140  & n4624;
  assign n2282 = ~n2280 & ~n2281;
  assign n2283 = pi268  & ~n4696;
  assign n2284 = pi396  & n4696;
  assign n2285 = ~n2283 & ~n2284;
  assign n2286 = ~n2282 & n2285;
  assign n2287 = n2282 & ~n2285;
  assign n2288 = pi11  & ~n4624;
  assign n2289 = pi139  & n4624;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = pi267  & ~n4696;
  assign n2292 = pi395  & n4696;
  assign n2293 = ~n2291 & ~n2292;
  assign n2294 = ~n2290 & n2293;
  assign n2295 = n2290 & ~n2293;
  assign n2296 = pi10  & ~n4624;
  assign n2297 = pi138  & n4624;
  assign n2298 = ~n2296 & ~n2297;
  assign n2299 = pi266  & ~n4696;
  assign n2300 = pi394  & n4696;
  assign n2301 = ~n2299 & ~n2300;
  assign n2302 = ~n2298 & n2301;
  assign n2303 = pi7  & ~n4624;
  assign n2304 = pi135  & n4624;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = pi263  & ~n4696;
  assign n2307 = pi391  & n4696;
  assign n2308 = ~n2306 & ~n2307;
  assign n2309 = ~n2305 & n2308;
  assign n2310 = pi261  & ~n4696;
  assign n2311 = pi389  & n4696;
  assign n2312 = ~n2310 & ~n2311;
  assign n2313 = pi260  & ~n4696;
  assign n2314 = pi388  & n4696;
  assign n2315 = ~n2313 & ~n2314;
  assign n2316 = pi3  & ~n4624;
  assign n2317 = pi131  & n4624;
  assign n2318 = ~n2316 & ~n2317;
  assign n2319 = pi259  & ~n4696;
  assign n2320 = pi387  & n4696;
  assign n2321 = ~n2319 & ~n2320;
  assign n2322 = n2318 & ~n2321;
  assign n2323 = ~n2318 & n2321;
  assign n2324 = pi2  & ~n4624;
  assign n2325 = pi130  & n4624;
  assign n2326 = ~n2324 & ~n2325;
  assign n2327 = pi258  & ~n4696;
  assign n2328 = pi386  & n4696;
  assign n2329 = ~n2327 & ~n2328;
  assign n2330 = n2326 & ~n2329;
  assign n2331 = ~n2326 & n2329;
  assign n2332 = pi257  & ~n4696;
  assign n2333 = pi385  & n4696;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = pi1  & ~n4624;
  assign n2336 = pi129  & n4624;
  assign n2337 = ~n2335 & ~n2336;
  assign n2338 = ~n2334 & n2337;
  assign n2339 = pi256  & ~n4696;
  assign n2340 = pi384  & n4696;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = pi0  & ~n4624;
  assign n2343 = pi128  & n4624;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = n2341 & ~n2344;
  assign n2346 = n2334 & ~n2337;
  assign n2347 = ~n2345 & ~n2346;
  assign n2348 = ~n2338 & ~n2347;
  assign n2349 = n2337 & ~n2345;
  assign n2350 = n2334 & ~n2349;
  assign n2351 = ~n2337 & n2345;
  assign n2352 = ~n2331 & ~n2351;
  assign n2353 = ~n2350 & n2352;
  assign n2354 = ~n2331 & ~n2348;
  assign n2355 = n2334 & n2345;
  assign n2356 = n2337 & ~n2355;
  assign n2357 = ~n2334 & ~n2345;
  assign n2358 = ~n2330 & ~n2357;
  assign n2359 = ~n2356 & n2358;
  assign n2360 = ~n2331 & ~n2359;
  assign n2361 = ~n2330 & ~n4697;
  assign n2362 = ~n2323 & n4698;
  assign n2363 = ~n2322 & ~n4698;
  assign n2364 = ~n2323 & ~n2363;
  assign n2365 = ~n2322 & ~n2362;
  assign n2366 = pi4  & ~n4624;
  assign n2367 = pi132  & n4624;
  assign n2368 = ~n2366 & ~n2367;
  assign n2369 = n4699 & n2368;
  assign n2370 = n2315 & ~n2369;
  assign n2371 = ~n4699 & ~n2368;
  assign n2372 = n2315 & ~n4699;
  assign n2373 = n2368 & ~n2372;
  assign n2374 = ~n2315 & n4699;
  assign n2375 = ~n2373 & ~n2374;
  assign n2376 = ~n2370 & ~n2371;
  assign n2377 = pi5  & ~n4624;
  assign n2378 = pi133  & n4624;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = ~n4700 & n2379;
  assign n2381 = n2312 & ~n2380;
  assign n2382 = n4700 & ~n2379;
  assign n2383 = n2312 & n4700;
  assign n2384 = n2379 & ~n2383;
  assign n2385 = ~n2312 & ~n4700;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = ~n2381 & ~n2382;
  assign n2388 = pi262  & ~n4696;
  assign n2389 = pi390  & n4696;
  assign n2390 = ~n2388 & ~n2389;
  assign n2391 = ~n4701 & ~n2390;
  assign n2392 = n4701 & n2390;
  assign n2393 = pi6  & ~n4624;
  assign n2394 = pi134  & n4624;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = ~n2392 & n2395;
  assign n2397 = ~n4701 & n2395;
  assign n2398 = n2390 & ~n2397;
  assign n2399 = n4701 & ~n2395;
  assign n2400 = ~n2398 & ~n2399;
  assign n2401 = ~n2391 & ~n2396;
  assign n2402 = ~n2309 & n4702;
  assign n2403 = n2305 & ~n2308;
  assign n2404 = pi8  & ~n4624;
  assign n2405 = pi136  & n4624;
  assign n2406 = ~n2404 & ~n2405;
  assign n2407 = pi264  & ~n4696;
  assign n2408 = pi392  & n4696;
  assign n2409 = ~n2407 & ~n2408;
  assign n2410 = n2406 & ~n2409;
  assign n2411 = ~n2403 & ~n2410;
  assign n2412 = ~n2402 & n2411;
  assign n2413 = ~n2406 & n2409;
  assign n2414 = pi9  & ~n4624;
  assign n2415 = pi137  & n4624;
  assign n2416 = ~n2414 & ~n2415;
  assign n2417 = pi265  & ~n4696;
  assign n2418 = pi393  & n4696;
  assign n2419 = ~n2417 & ~n2418;
  assign n2420 = ~n2416 & n2419;
  assign n2421 = ~n2413 & ~n2420;
  assign n2422 = ~n2412 & n2421;
  assign n2423 = n2298 & ~n2301;
  assign n2424 = n2416 & ~n2419;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = ~n4702 & ~n2403;
  assign n2427 = ~n2309 & ~n2413;
  assign n2428 = ~n2426 & n2427;
  assign n2429 = ~n2309 & ~n2426;
  assign n2430 = n2406 & n2429;
  assign n2431 = n2409 & ~n2430;
  assign n2432 = ~n2406 & ~n2429;
  assign n2433 = ~n2431 & ~n2432;
  assign n2434 = ~n2410 & ~n2428;
  assign n2435 = n2416 & n4703;
  assign n2436 = n2419 & ~n2435;
  assign n2437 = ~n2416 & ~n4703;
  assign n2438 = ~n2436 & ~n2437;
  assign n2439 = ~n2423 & ~n2438;
  assign n2440 = ~n2422 & n2425;
  assign n2441 = ~n2302 & ~n4704;
  assign n2442 = ~n2295 & ~n2441;
  assign n2443 = ~n2294 & ~n2442;
  assign n2444 = ~n2287 & ~n2443;
  assign n2445 = ~n2286 & ~n2444;
  assign n2446 = ~n2279 & ~n2445;
  assign n2447 = ~n2275 & n2278;
  assign n2448 = pi14  & ~n4624;
  assign n2449 = pi142  & n4624;
  assign n2450 = ~n2448 & ~n2449;
  assign n2451 = pi270  & ~n4696;
  assign n2452 = pi398  & n4696;
  assign n2453 = ~n2451 & ~n2452;
  assign n2454 = ~n2450 & n2453;
  assign n2455 = ~n2447 & ~n2454;
  assign n2456 = ~n2446 & n2455;
  assign n2457 = n2450 & ~n2453;
  assign n2458 = pi15  & ~n4624;
  assign n2459 = pi143  & n4624;
  assign n2460 = ~n2458 & ~n2459;
  assign n2461 = pi271  & ~n4696;
  assign n2462 = pi399  & n4696;
  assign n2463 = ~n2461 & ~n2462;
  assign n2464 = n2460 & ~n2463;
  assign n2465 = ~n2457 & ~n2464;
  assign n2466 = ~n2446 & ~n2447;
  assign n2467 = ~n2457 & ~n2466;
  assign n2468 = ~n2454 & ~n2467;
  assign n2469 = ~n2464 & ~n2468;
  assign n2470 = ~n2456 & n2465;
  assign n2471 = ~n2460 & n2463;
  assign n2472 = pi16  & ~n4624;
  assign n2473 = pi144  & n4624;
  assign n2474 = ~n2472 & ~n2473;
  assign n2475 = pi272  & ~n4696;
  assign n2476 = pi400  & n4696;
  assign n2477 = ~n2475 & ~n2476;
  assign n2478 = ~n2474 & n2477;
  assign n2479 = ~n2471 & ~n2478;
  assign n2480 = ~n4705 & n2479;
  assign n2481 = n2474 & ~n2477;
  assign n2482 = n2268 & ~n2271;
  assign n2483 = ~n2481 & ~n2482;
  assign n2484 = ~n2480 & n2483;
  assign n2485 = ~n4705 & ~n2471;
  assign n2486 = n2474 & n2485;
  assign n2487 = n2477 & ~n2486;
  assign n2488 = ~n2474 & ~n2485;
  assign n2489 = ~n2487 & ~n2488;
  assign n2490 = ~n2480 & ~n2481;
  assign n2491 = n2268 & n4706;
  assign n2492 = n2271 & ~n2491;
  assign n2493 = ~n2268 & ~n4706;
  assign n2494 = ~n2492 & ~n2493;
  assign n2495 = ~n2272 & ~n2484;
  assign n2496 = ~n2265 & ~n4707;
  assign n2497 = ~n2264 & ~n2496;
  assign n2498 = ~n2257 & ~n2497;
  assign n2499 = ~n2256 & ~n2498;
  assign n2500 = ~n2249 & ~n2499;
  assign n2501 = ~n2248 & ~n2500;
  assign n2502 = ~n2241 & ~n2501;
  assign n2503 = ~n2237 & n2240;
  assign n2504 = pi22  & ~n4624;
  assign n2505 = pi150  & n4624;
  assign n2506 = ~n2504 & ~n2505;
  assign n2507 = pi278  & ~n4696;
  assign n2508 = pi406  & n4696;
  assign n2509 = ~n2507 & ~n2508;
  assign n2510 = ~n2506 & n2509;
  assign n2511 = ~n2503 & ~n2510;
  assign n2512 = ~n2502 & n2511;
  assign n2513 = n2506 & ~n2509;
  assign n2514 = pi23  & ~n4624;
  assign n2515 = pi151  & n4624;
  assign n2516 = ~n2514 & ~n2515;
  assign n2517 = pi279  & ~n4696;
  assign n2518 = pi407  & n4696;
  assign n2519 = ~n2517 & ~n2518;
  assign n2520 = n2516 & ~n2519;
  assign n2521 = ~n2513 & ~n2520;
  assign n2522 = ~n2502 & ~n2503;
  assign n2523 = ~n2513 & ~n2522;
  assign n2524 = ~n2510 & ~n2523;
  assign n2525 = ~n2520 & ~n2524;
  assign n2526 = ~n2512 & n2521;
  assign n2527 = ~n2516 & n2519;
  assign n2528 = pi24  & ~n4624;
  assign n2529 = pi152  & n4624;
  assign n2530 = ~n2528 & ~n2529;
  assign n2531 = pi280  & ~n4696;
  assign n2532 = pi408  & n4696;
  assign n2533 = ~n2531 & ~n2532;
  assign n2534 = ~n2530 & n2533;
  assign n2535 = ~n2527 & ~n2534;
  assign n2536 = ~n4708 & n2535;
  assign n2537 = n2530 & ~n2533;
  assign n2538 = n2230 & ~n2233;
  assign n2539 = ~n2537 & ~n2538;
  assign n2540 = ~n2536 & n2539;
  assign n2541 = ~n4708 & ~n2527;
  assign n2542 = n2530 & n2541;
  assign n2543 = n2533 & ~n2542;
  assign n2544 = ~n2530 & ~n2541;
  assign n2545 = ~n2543 & ~n2544;
  assign n2546 = ~n2536 & ~n2537;
  assign n2547 = n2230 & n4709;
  assign n2548 = n2233 & ~n2547;
  assign n2549 = ~n2230 & ~n4709;
  assign n2550 = ~n2548 & ~n2549;
  assign n2551 = ~n2234 & ~n2540;
  assign n2552 = ~n2227 & ~n4710;
  assign n2553 = ~n2226 & ~n2552;
  assign n2554 = ~n2219 & ~n2553;
  assign n2555 = ~n2218 & ~n2554;
  assign n2556 = ~n2211 & ~n2555;
  assign n2557 = ~n1425 & n2210;
  assign n2558 = pi29  & ~n4624;
  assign n2559 = pi157  & n4624;
  assign n2560 = ~n2558 & ~n2559;
  assign n2561 = pi285  & ~n4696;
  assign n2562 = pi413  & n4696;
  assign n2563 = ~n2561 & ~n2562;
  assign n2564 = ~n2560 & n2563;
  assign n2565 = ~n2557 & ~n2564;
  assign n2566 = ~n2556 & n2565;
  assign n2567 = n2560 & ~n2563;
  assign n2568 = pi30  & ~n4624;
  assign n2569 = pi158  & n4624;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = pi286  & ~n4696;
  assign n2572 = pi414  & n4696;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = n2570 & ~n2573;
  assign n2575 = ~n2567 & ~n2574;
  assign n2576 = ~n2556 & ~n2557;
  assign n2577 = ~n2567 & ~n2576;
  assign n2578 = ~n2564 & ~n2577;
  assign n2579 = ~n2574 & ~n2578;
  assign n2580 = ~n2566 & n2575;
  assign n2581 = ~n2570 & n2573;
  assign n2582 = pi31  & ~n4624;
  assign n2583 = pi159  & n4624;
  assign n2584 = ~n2582 & ~n2583;
  assign n2585 = pi287  & ~n4696;
  assign n2586 = pi415  & n4696;
  assign n2587 = ~n2585 & ~n2586;
  assign n2588 = ~n2584 & n2587;
  assign n2589 = ~n2581 & ~n2588;
  assign n2590 = ~n4711 & n2589;
  assign n2591 = pi33  & ~n4624;
  assign n2592 = pi161  & n4624;
  assign n2593 = ~n2591 & ~n2592;
  assign n2594 = pi289  & ~n4696;
  assign n2595 = pi417  & n4696;
  assign n2596 = ~n2594 & ~n2595;
  assign n2597 = n2593 & ~n2596;
  assign n2598 = pi35  & ~n4624;
  assign n2599 = pi163  & n4624;
  assign n2600 = ~n2598 & ~n2599;
  assign n2601 = pi291  & ~n4696;
  assign n2602 = pi419  & n4696;
  assign n2603 = ~n2601 & ~n2602;
  assign n2604 = n2600 & ~n2603;
  assign n2605 = pi290  & ~n4696;
  assign n2606 = pi418  & n4696;
  assign n2607 = ~n2605 & ~n2606;
  assign n2608 = pi34  & ~n4624;
  assign n2609 = pi162  & n4624;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = ~n2607 & n2610;
  assign n2612 = ~n2604 & ~n2611;
  assign n2613 = ~n2597 & n2612;
  assign n2614 = pi39  & ~n4624;
  assign n2615 = pi167  & n4624;
  assign n2616 = ~n2614 & ~n2615;
  assign n2617 = pi295  & ~n4696;
  assign n2618 = pi423  & n4696;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = n2616 & ~n2619;
  assign n2621 = pi37  & ~n4624;
  assign n2622 = pi165  & n4624;
  assign n2623 = ~n2621 & ~n2622;
  assign n2624 = pi293  & ~n4696;
  assign n2625 = pi421  & n4696;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = n2623 & ~n2626;
  assign n2628 = pi294  & ~n4696;
  assign n2629 = pi422  & n4696;
  assign n2630 = ~n2628 & ~n2629;
  assign n2631 = pi38  & ~n4624;
  assign n2632 = pi166  & n4624;
  assign n2633 = ~n2631 & ~n2632;
  assign n2634 = ~n2630 & n2633;
  assign n2635 = ~n2627 & ~n2634;
  assign n2636 = ~n2620 & n2635;
  assign n2637 = pi288  & ~n4696;
  assign n2638 = pi416  & n4696;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = pi32  & ~n4624;
  assign n2641 = pi160  & n4624;
  assign n2642 = ~n2640 & ~n2641;
  assign n2643 = ~n2639 & n2642;
  assign n2644 = n2584 & ~n2587;
  assign n2645 = pi36  & ~n4624;
  assign n2646 = pi164  & n4624;
  assign n2647 = ~n2645 & ~n2646;
  assign n2648 = pi292  & ~n4696;
  assign n2649 = pi420  & n4696;
  assign n2650 = ~n2648 & ~n2649;
  assign n2651 = n2647 & ~n2650;
  assign n2652 = ~n2644 & ~n2651;
  assign n2653 = ~n2643 & n2652;
  assign n2654 = n2636 & n2653;
  assign n2655 = ~n2620 & ~n2634;
  assign n2656 = ~n2627 & ~n2651;
  assign n2657 = n2636 & ~n2651;
  assign n2658 = n2655 & n2656;
  assign n2659 = ~n2643 & ~n2644;
  assign n2660 = n2613 & n2659;
  assign n2661 = n4712 & n2660;
  assign n2662 = n2613 & n2654;
  assign n2663 = ~n4711 & ~n2581;
  assign n2664 = ~n2644 & ~n2663;
  assign n2665 = ~n2588 & ~n2664;
  assign n2666 = n2613 & n4712;
  assign n2667 = ~n2665 & n2666;
  assign n2668 = ~n2643 & n2667;
  assign n2669 = ~n2590 & n4713;
  assign n2670 = n2639 & ~n2642;
  assign n2671 = ~n2593 & n2596;
  assign n2672 = ~n2670 & ~n2671;
  assign n2673 = n2613 & ~n2672;
  assign n2674 = n2607 & ~n2610;
  assign n2675 = ~n2604 & n2607;
  assign n2676 = ~n2610 & n2675;
  assign n2677 = ~n2604 & n2674;
  assign n2678 = ~n2600 & n2603;
  assign n2679 = ~n4715 & ~n2678;
  assign n2680 = ~n2673 & ~n4715;
  assign n2681 = ~n2678 & n2680;
  assign n2682 = ~n2673 & n2679;
  assign n2683 = n4712 & ~n4716;
  assign n2684 = n2630 & ~n2633;
  assign n2685 = ~n2620 & n2630;
  assign n2686 = ~n2633 & n2685;
  assign n2687 = ~n2620 & n2684;
  assign n2688 = ~n2616 & n2619;
  assign n2689 = ~n4717 & ~n2688;
  assign n2690 = ~n2647 & n2650;
  assign n2691 = ~n2623 & n2626;
  assign n2692 = ~n2690 & ~n2691;
  assign n2693 = ~n2627 & n2690;
  assign n2694 = ~n2691 & ~n2693;
  assign n2695 = n2655 & ~n2694;
  assign n2696 = n2636 & ~n2692;
  assign n2697 = n2689 & ~n4718;
  assign n2698 = ~n2651 & ~n4716;
  assign n2699 = n2692 & ~n2698;
  assign n2700 = n2636 & ~n2699;
  assign n2701 = n2689 & ~n2700;
  assign n2702 = ~n2683 & ~n4717;
  assign n2703 = ~n4718 & n2702;
  assign n2704 = ~n2688 & n2703;
  assign n2705 = ~n2683 & n2697;
  assign n2706 = ~n4714 & n4719;
  assign n2707 = pi47  & ~n4624;
  assign n2708 = pi175  & n4624;
  assign n2709 = ~n2707 & ~n2708;
  assign n2710 = pi303  & ~n4696;
  assign n2711 = pi431  & n4696;
  assign n2712 = ~n2710 & ~n2711;
  assign n2713 = n2709 & ~n2712;
  assign n2714 = pi302  & ~n4696;
  assign n2715 = pi430  & n4696;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = pi46  & ~n4624;
  assign n2718 = pi174  & n4624;
  assign n2719 = ~n2717 & ~n2718;
  assign n2720 = ~n2716 & n2719;
  assign n2721 = ~n2713 & ~n2720;
  assign n2722 = pi45  & ~n4624;
  assign n2723 = pi173  & n4624;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = pi301  & ~n4696;
  assign n2726 = pi429  & n4696;
  assign n2727 = ~n2725 & ~n2726;
  assign n2728 = n2724 & ~n2727;
  assign n2729 = pi44  & ~n4624;
  assign n2730 = pi172  & n4624;
  assign n2731 = ~n2729 & ~n2730;
  assign n2732 = pi300  & ~n4696;
  assign n2733 = pi428  & n4696;
  assign n2734 = ~n2732 & ~n2733;
  assign n2735 = n2731 & ~n2734;
  assign n2736 = ~n2728 & ~n2735;
  assign n2737 = ~n2720 & ~n2728;
  assign n2738 = ~n2713 & n2737;
  assign n2739 = ~n2735 & n2738;
  assign n2740 = n2721 & n2736;
  assign n2741 = pi43  & ~n4624;
  assign n2742 = pi171  & n4624;
  assign n2743 = ~n2741 & ~n2742;
  assign n2744 = pi299  & ~n4696;
  assign n2745 = pi427  & n4696;
  assign n2746 = ~n2744 & ~n2745;
  assign n2747 = n2743 & ~n2746;
  assign n2748 = pi42  & ~n4624;
  assign n2749 = pi170  & n4624;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = pi298  & ~n4696;
  assign n2752 = pi426  & n4696;
  assign n2753 = ~n2751 & ~n2752;
  assign n2754 = n2750 & ~n2753;
  assign n2755 = ~n2747 & ~n2754;
  assign n2756 = pi41  & ~n4624;
  assign n2757 = pi169  & n4624;
  assign n2758 = ~n2756 & ~n2757;
  assign n2759 = pi297  & ~n4696;
  assign n2760 = pi425  & n4696;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = n2758 & ~n2761;
  assign n2763 = pi40  & ~n4624;
  assign n2764 = pi168  & n4624;
  assign n2765 = ~n2763 & ~n2764;
  assign n2766 = pi296  & ~n4696;
  assign n2767 = pi424  & n4696;
  assign n2768 = ~n2766 & ~n2767;
  assign n2769 = n2765 & ~n2768;
  assign n2770 = ~n2762 & ~n2769;
  assign n2771 = n2755 & n2770;
  assign n2772 = ~n2735 & ~n2769;
  assign n2773 = ~n2762 & n2772;
  assign n2774 = n2755 & n2773;
  assign n2775 = n2738 & n2774;
  assign n2776 = n4720 & n2771;
  assign n2777 = ~n2706 & n4721;
  assign n2778 = ~n2743 & n2746;
  assign n2779 = ~n2765 & n2768;
  assign n2780 = ~n2762 & n2779;
  assign n2781 = ~n2758 & n2761;
  assign n2782 = ~n2750 & n2753;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = ~n2780 & ~n2781;
  assign n2785 = ~n2782 & n2784;
  assign n2786 = ~n2780 & n2783;
  assign n2787 = n2755 & ~n4722;
  assign n2788 = ~n2778 & ~n2787;
  assign n2789 = n4720 & ~n2788;
  assign n2790 = n2716 & ~n2719;
  assign n2791 = ~n2713 & n2790;
  assign n2792 = ~n2709 & n2712;
  assign n2793 = ~n2791 & ~n2792;
  assign n2794 = ~n2731 & n2734;
  assign n2795 = ~n2724 & n2727;
  assign n2796 = ~n2794 & ~n2795;
  assign n2797 = ~n2728 & n2794;
  assign n2798 = ~n2795 & ~n2797;
  assign n2799 = n2721 & ~n2798;
  assign n2800 = n2738 & ~n2796;
  assign n2801 = n2793 & ~n4723;
  assign n2802 = ~n2735 & ~n2788;
  assign n2803 = n2796 & ~n2802;
  assign n2804 = n2738 & ~n2803;
  assign n2805 = n2793 & ~n2804;
  assign n2806 = ~n2789 & n2801;
  assign n2807 = ~n2777 & ~n2791;
  assign n2808 = ~n4723 & n2807;
  assign n2809 = ~n2789 & n2808;
  assign n2810 = ~n2792 & n2809;
  assign n2811 = ~n2777 & n4724;
  assign n2812 = pi55  & ~n4624;
  assign n2813 = pi183  & n4624;
  assign n2814 = ~n2812 & ~n2813;
  assign n2815 = pi311  & ~n4696;
  assign n2816 = pi439  & n4696;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = n2814 & ~n2817;
  assign n2819 = pi310  & ~n4696;
  assign n2820 = pi438  & n4696;
  assign n2821 = ~n2819 & ~n2820;
  assign n2822 = pi54  & ~n4624;
  assign n2823 = pi182  & n4624;
  assign n2824 = ~n2822 & ~n2823;
  assign n2825 = ~n2821 & n2824;
  assign n2826 = ~n2818 & ~n2825;
  assign n2827 = pi53  & ~n4624;
  assign n2828 = pi181  & n4624;
  assign n2829 = ~n2827 & ~n2828;
  assign n2830 = pi309  & ~n4696;
  assign n2831 = pi437  & n4696;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = n2829 & ~n2832;
  assign n2834 = pi308  & ~n4696;
  assign n2835 = pi436  & n4696;
  assign n2836 = ~n2834 & ~n2835;
  assign n2837 = pi52  & ~n4624;
  assign n2838 = pi180  & n4624;
  assign n2839 = ~n2837 & ~n2838;
  assign n2840 = ~n2836 & n2839;
  assign n2841 = ~n2833 & ~n2840;
  assign n2842 = n2826 & n2841;
  assign n2843 = pi49  & ~n4624;
  assign n2844 = pi177  & n4624;
  assign n2845 = ~n2843 & ~n2844;
  assign n2846 = pi305  & ~n4696;
  assign n2847 = pi433  & n4696;
  assign n2848 = ~n2846 & ~n2847;
  assign n2849 = n2845 & ~n2848;
  assign n2850 = pi51  & ~n4624;
  assign n2851 = pi179  & n4624;
  assign n2852 = ~n2850 & ~n2851;
  assign n2853 = pi307  & ~n4696;
  assign n2854 = pi435  & n4696;
  assign n2855 = ~n2853 & ~n2854;
  assign n2856 = n2852 & ~n2855;
  assign n2857 = pi306  & ~n4696;
  assign n2858 = pi434  & n4696;
  assign n2859 = ~n2857 & ~n2858;
  assign n2860 = pi50  & ~n4624;
  assign n2861 = pi178  & n4624;
  assign n2862 = ~n2860 & ~n2861;
  assign n2863 = ~n2859 & n2862;
  assign n2864 = ~n2856 & ~n2863;
  assign n2865 = ~n2849 & n2864;
  assign n2866 = pi304  & ~n4696;
  assign n2867 = pi432  & n4696;
  assign n2868 = ~n2866 & ~n2867;
  assign n2869 = pi48  & ~n4624;
  assign n2870 = pi176  & n4624;
  assign n2871 = ~n2869 & ~n2870;
  assign n2872 = ~n2868 & n2871;
  assign n2873 = n2865 & ~n2872;
  assign n2874 = n2842 & n2865;
  assign n2875 = ~n2872 & n2874;
  assign n2876 = n2842 & ~n2872;
  assign n2877 = n2865 & n2876;
  assign n2878 = n2842 & n2873;
  assign n2879 = ~n4725 & n4726;
  assign n2880 = n2868 & ~n2871;
  assign n2881 = ~n2845 & n2848;
  assign n2882 = ~n2880 & ~n2881;
  assign n2883 = n2865 & ~n2882;
  assign n2884 = ~n2852 & n2855;
  assign n2885 = n2859 & ~n2862;
  assign n2886 = ~n2856 & n2859;
  assign n2887 = ~n2862 & n2886;
  assign n2888 = ~n2856 & n2885;
  assign n2889 = ~n2884 & ~n4727;
  assign n2890 = ~n2883 & ~n4727;
  assign n2891 = ~n2884 & n2890;
  assign n2892 = ~n2883 & n2889;
  assign n2893 = n2842 & ~n4728;
  assign n2894 = ~n2814 & n2817;
  assign n2895 = n2836 & ~n2839;
  assign n2896 = ~n2833 & n2895;
  assign n2897 = ~n2829 & n2832;
  assign n2898 = n2821 & ~n2824;
  assign n2899 = ~n2897 & ~n2898;
  assign n2900 = ~n2896 & ~n2897;
  assign n2901 = ~n2898 & n2900;
  assign n2902 = ~n2896 & n2899;
  assign n2903 = n2826 & ~n4729;
  assign n2904 = ~n2894 & ~n2903;
  assign n2905 = ~n2893 & ~n2903;
  assign n2906 = ~n2894 & n2905;
  assign n2907 = ~n2893 & n2904;
  assign n2908 = ~n2879 & n4730;
  assign n2909 = pi63  & ~n4624;
  assign n2910 = pi191  & n4624;
  assign n2911 = ~n2909 & ~n2910;
  assign n2912 = pi319  & ~n4696;
  assign n2913 = pi447  & n4696;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = n2911 & ~n2914;
  assign n2916 = pi318  & ~n4696;
  assign n2917 = pi446  & n4696;
  assign n2918 = ~n2916 & ~n2917;
  assign n2919 = pi62  & ~n4624;
  assign n2920 = pi190  & n4624;
  assign n2921 = ~n2919 & ~n2920;
  assign n2922 = ~n2918 & n2921;
  assign n2923 = ~n2915 & ~n2922;
  assign n2924 = pi61  & ~n4624;
  assign n2925 = pi189  & n4624;
  assign n2926 = ~n2924 & ~n2925;
  assign n2927 = pi317  & ~n4696;
  assign n2928 = pi445  & n4696;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = n2926 & ~n2929;
  assign n2931 = pi60  & ~n4624;
  assign n2932 = pi188  & n4624;
  assign n2933 = ~n2931 & ~n2932;
  assign n2934 = pi316  & ~n4696;
  assign n2935 = pi444  & n4696;
  assign n2936 = ~n2934 & ~n2935;
  assign n2937 = n2933 & ~n2936;
  assign n2938 = ~n2930 & ~n2937;
  assign n2939 = ~n2922 & ~n2930;
  assign n2940 = ~n2915 & n2939;
  assign n2941 = ~n2937 & n2940;
  assign n2942 = n2923 & n2938;
  assign n2943 = pi59  & ~n4624;
  assign n2944 = pi187  & n4624;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = pi315  & ~n4696;
  assign n2947 = pi443  & n4696;
  assign n2948 = ~n2946 & ~n2947;
  assign n2949 = n2945 & ~n2948;
  assign n2950 = pi58  & ~n4624;
  assign n2951 = pi186  & n4624;
  assign n2952 = ~n2950 & ~n2951;
  assign n2953 = pi314  & ~n4696;
  assign n2954 = pi442  & n4696;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = n2952 & ~n2955;
  assign n2957 = ~n2949 & ~n2956;
  assign n2958 = pi57  & ~n4624;
  assign n2959 = pi185  & n4624;
  assign n2960 = ~n2958 & ~n2959;
  assign n2961 = pi313  & ~n4696;
  assign n2962 = pi441  & n4696;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = n2960 & ~n2963;
  assign n2965 = pi56  & ~n4624;
  assign n2966 = pi184  & n4624;
  assign n2967 = ~n2965 & ~n2966;
  assign n2968 = pi312  & ~n4696;
  assign n2969 = pi440  & n4696;
  assign n2970 = ~n2968 & ~n2969;
  assign n2971 = n2967 & ~n2970;
  assign n2972 = ~n2964 & ~n2971;
  assign n2973 = n2957 & n2972;
  assign n2974 = ~n2937 & ~n2971;
  assign n2975 = ~n2964 & n2974;
  assign n2976 = n2957 & n2975;
  assign n2977 = n2940 & n2976;
  assign n2978 = n4731 & n2972;
  assign n2979 = n2957 & n2978;
  assign n2980 = n4731 & n2973;
  assign n2981 = ~n2908 & n4732;
  assign n2982 = ~n2945 & n2948;
  assign n2983 = ~n2967 & n2970;
  assign n2984 = ~n2964 & n2983;
  assign n2985 = ~n2960 & n2963;
  assign n2986 = ~n2952 & n2955;
  assign n2987 = ~n2985 & ~n2986;
  assign n2988 = ~n2984 & ~n2985;
  assign n2989 = ~n2986 & n2988;
  assign n2990 = ~n2984 & n2987;
  assign n2991 = n2957 & ~n4733;
  assign n2992 = ~n2982 & ~n2991;
  assign n2993 = n4731 & ~n2992;
  assign n2994 = n2918 & ~n2921;
  assign n2995 = ~n2915 & n2994;
  assign n2996 = ~n2911 & n2914;
  assign n2997 = ~n2995 & ~n2996;
  assign n2998 = ~n2933 & n2936;
  assign n2999 = ~n2926 & n2929;
  assign n3000 = ~n2998 & ~n2999;
  assign n3001 = ~n2930 & n2998;
  assign n3002 = ~n2999 & ~n3001;
  assign n3003 = n2923 & ~n3002;
  assign n3004 = n2940 & ~n3000;
  assign n3005 = n2997 & ~n4734;
  assign n3006 = ~n2937 & ~n2992;
  assign n3007 = n3000 & ~n3006;
  assign n3008 = n2940 & ~n3007;
  assign n3009 = n2997 & ~n3008;
  assign n3010 = ~n2993 & n3005;
  assign n3011 = ~n2981 & ~n2995;
  assign n3012 = ~n4734 & n3011;
  assign n3013 = ~n2993 & n3012;
  assign n3014 = ~n2996 & n3013;
  assign n3015 = ~n2981 & n4735;
  assign n3016 = pi67  & ~n4624;
  assign n3017 = pi195  & n4624;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = pi323  & ~n4696;
  assign n3020 = pi451  & n4696;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = n3018 & ~n3021;
  assign n3023 = pi322  & ~n4696;
  assign n3024 = pi450  & n4696;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = pi66  & ~n4624;
  assign n3027 = pi194  & n4624;
  assign n3028 = ~n3026 & ~n3027;
  assign n3029 = ~n3025 & n3028;
  assign n3030 = ~n3022 & ~n3029;
  assign n3031 = pi65  & ~n4624;
  assign n3032 = pi193  & n4624;
  assign n3033 = ~n3031 & ~n3032;
  assign n3034 = pi321  & ~n4696;
  assign n3035 = pi449  & n4696;
  assign n3036 = ~n3034 & ~n3035;
  assign n3037 = n3033 & ~n3036;
  assign n3038 = pi320  & ~n4696;
  assign n3039 = pi448  & n4696;
  assign n3040 = ~n3038 & ~n3039;
  assign n3041 = pi64  & ~n4624;
  assign n3042 = pi192  & n4624;
  assign n3043 = ~n3041 & ~n3042;
  assign n3044 = ~n3040 & n3043;
  assign n3045 = ~n3037 & ~n3044;
  assign n3046 = n3030 & n3045;
  assign n3047 = ~n4736 & ~n3037;
  assign n3048 = ~n3044 & n3047;
  assign n3049 = n3030 & n3048;
  assign n3050 = ~n4736 & n3046;
  assign n3051 = ~n3018 & n3021;
  assign n3052 = n3040 & ~n3043;
  assign n3053 = ~n3037 & n3040;
  assign n3054 = ~n3043 & n3053;
  assign n3055 = ~n3037 & n3052;
  assign n3056 = ~n3033 & n3036;
  assign n3057 = n3025 & ~n3028;
  assign n3058 = ~n3056 & ~n3057;
  assign n3059 = ~n4738 & ~n3056;
  assign n3060 = ~n3057 & n3059;
  assign n3061 = ~n4738 & n3058;
  assign n3062 = n3030 & ~n4739;
  assign n3063 = ~n3051 & ~n3062;
  assign n3064 = ~n4737 & n3063;
  assign n3065 = pi71  & ~n4624;
  assign n3066 = pi199  & n4624;
  assign n3067 = ~n3065 & ~n3066;
  assign n3068 = pi327  & ~n4696;
  assign n3069 = pi455  & n4696;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = n3067 & ~n3070;
  assign n3072 = pi326  & ~n4696;
  assign n3073 = pi454  & n4696;
  assign n3074 = ~n3072 & ~n3073;
  assign n3075 = pi70  & ~n4624;
  assign n3076 = pi198  & n4624;
  assign n3077 = ~n3075 & ~n3076;
  assign n3078 = ~n3074 & n3077;
  assign n3079 = ~n3071 & ~n3078;
  assign n3080 = pi69  & ~n4624;
  assign n3081 = pi197  & n4624;
  assign n3082 = ~n3080 & ~n3081;
  assign n3083 = pi325  & ~n4696;
  assign n3084 = pi453  & n4696;
  assign n3085 = ~n3083 & ~n3084;
  assign n3086 = n3082 & ~n3085;
  assign n3087 = pi68  & ~n4624;
  assign n3088 = pi196  & n4624;
  assign n3089 = ~n3087 & ~n3088;
  assign n3090 = pi324  & ~n4696;
  assign n3091 = pi452  & n4696;
  assign n3092 = ~n3090 & ~n3091;
  assign n3093 = n3089 & ~n3092;
  assign n3094 = ~n3086 & ~n3093;
  assign n3095 = n3079 & n3094;
  assign n3096 = ~n3064 & n3095;
  assign n3097 = ~n3067 & n3070;
  assign n3098 = ~n3089 & n3092;
  assign n3099 = ~n3086 & n3098;
  assign n3100 = n3074 & ~n3077;
  assign n3101 = ~n3082 & n3085;
  assign n3102 = ~n3100 & ~n3101;
  assign n3103 = ~n3099 & n3102;
  assign n3104 = n3079 & ~n3103;
  assign n3105 = ~n3099 & ~n3101;
  assign n3106 = n3079 & ~n3105;
  assign n3107 = ~n3071 & n3100;
  assign n3108 = ~n3097 & ~n3107;
  assign n3109 = ~n3106 & n3108;
  assign n3110 = ~n3097 & ~n3104;
  assign n3111 = ~n3096 & ~n3107;
  assign n3112 = ~n3106 & n3111;
  assign n3113 = ~n3097 & n3112;
  assign n3114 = ~n3096 & n4740;
  assign n3115 = pi75  & ~n4624;
  assign n3116 = pi203  & n4624;
  assign n3117 = ~n3115 & ~n3116;
  assign n3118 = pi331  & ~n4696;
  assign n3119 = pi459  & n4696;
  assign n3120 = ~n3118 & ~n3119;
  assign n3121 = n3117 & ~n3120;
  assign n3122 = pi330  & ~n4696;
  assign n3123 = pi458  & n4696;
  assign n3124 = ~n3122 & ~n3123;
  assign n3125 = pi74  & ~n4624;
  assign n3126 = pi202  & n4624;
  assign n3127 = ~n3125 & ~n3126;
  assign n3128 = ~n3124 & n3127;
  assign n3129 = ~n3121 & ~n3128;
  assign n3130 = pi73  & ~n4624;
  assign n3131 = pi201  & n4624;
  assign n3132 = ~n3130 & ~n3131;
  assign n3133 = pi329  & ~n4696;
  assign n3134 = pi457  & n4696;
  assign n3135 = ~n3133 & ~n3134;
  assign n3136 = n3132 & ~n3135;
  assign n3137 = pi328  & ~n4696;
  assign n3138 = pi456  & n4696;
  assign n3139 = ~n3137 & ~n3138;
  assign n3140 = pi72  & ~n4624;
  assign n3141 = pi200  & n4624;
  assign n3142 = ~n3140 & ~n3141;
  assign n3143 = ~n3139 & n3142;
  assign n3144 = ~n3136 & ~n3143;
  assign n3145 = n3129 & n3144;
  assign n3146 = ~n4741 & n3145;
  assign n3147 = ~n3117 & n3120;
  assign n3148 = n3139 & ~n3142;
  assign n3149 = ~n3136 & n3148;
  assign n3150 = ~n3132 & n3135;
  assign n3151 = n3124 & ~n3127;
  assign n3152 = ~n3150 & ~n3151;
  assign n3153 = ~n3149 & ~n3150;
  assign n3154 = ~n3151 & n3153;
  assign n3155 = ~n3149 & n3152;
  assign n3156 = n3129 & ~n4742;
  assign n3157 = ~n3147 & ~n3156;
  assign n3158 = ~n3146 & n3157;
  assign n3159 = pi79  & ~n4624;
  assign n3160 = pi207  & n4624;
  assign n3161 = ~n3159 & ~n3160;
  assign n3162 = pi335  & ~n4696;
  assign n3163 = pi463  & n4696;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = n3161 & ~n3164;
  assign n3166 = pi334  & ~n4696;
  assign n3167 = pi462  & n4696;
  assign n3168 = ~n3166 & ~n3167;
  assign n3169 = pi78  & ~n4624;
  assign n3170 = pi206  & n4624;
  assign n3171 = ~n3169 & ~n3170;
  assign n3172 = ~n3168 & n3171;
  assign n3173 = ~n3165 & ~n3172;
  assign n3174 = pi77  & ~n4624;
  assign n3175 = pi205  & n4624;
  assign n3176 = ~n3174 & ~n3175;
  assign n3177 = pi333  & ~n4696;
  assign n3178 = pi461  & n4696;
  assign n3179 = ~n3177 & ~n3178;
  assign n3180 = n3176 & ~n3179;
  assign n3181 = pi76  & ~n4624;
  assign n3182 = pi204  & n4624;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = pi332  & ~n4696;
  assign n3185 = pi460  & n4696;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = n3183 & ~n3186;
  assign n3188 = ~n3180 & ~n3187;
  assign n3189 = n3173 & n3188;
  assign n3190 = ~n3158 & n3189;
  assign n3191 = ~n3161 & n3164;
  assign n3192 = ~n3183 & n3186;
  assign n3193 = ~n3180 & n3192;
  assign n3194 = n3168 & ~n3171;
  assign n3195 = ~n3176 & n3179;
  assign n3196 = ~n3194 & ~n3195;
  assign n3197 = ~n3193 & n3196;
  assign n3198 = n3173 & ~n3197;
  assign n3199 = ~n3193 & ~n3195;
  assign n3200 = n3173 & ~n3199;
  assign n3201 = ~n3165 & n3194;
  assign n3202 = ~n3191 & ~n3201;
  assign n3203 = ~n3200 & n3202;
  assign n3204 = ~n3191 & ~n3198;
  assign n3205 = ~n3190 & ~n3201;
  assign n3206 = ~n3200 & n3205;
  assign n3207 = ~n3191 & n3206;
  assign n3208 = ~n3190 & n4743;
  assign n3209 = pi83  & ~n4624;
  assign n3210 = pi211  & n4624;
  assign n3211 = ~n3209 & ~n3210;
  assign n3212 = pi339  & ~n4696;
  assign n3213 = pi467  & n4696;
  assign n3214 = ~n3212 & ~n3213;
  assign n3215 = n3211 & ~n3214;
  assign n3216 = pi338  & ~n4696;
  assign n3217 = pi466  & n4696;
  assign n3218 = ~n3216 & ~n3217;
  assign n3219 = pi82  & ~n4624;
  assign n3220 = pi210  & n4624;
  assign n3221 = ~n3219 & ~n3220;
  assign n3222 = ~n3218 & n3221;
  assign n3223 = ~n3215 & ~n3222;
  assign n3224 = pi81  & ~n4624;
  assign n3225 = pi209  & n4624;
  assign n3226 = ~n3224 & ~n3225;
  assign n3227 = pi337  & ~n4696;
  assign n3228 = pi465  & n4696;
  assign n3229 = ~n3227 & ~n3228;
  assign n3230 = n3226 & ~n3229;
  assign n3231 = pi336  & ~n4696;
  assign n3232 = pi464  & n4696;
  assign n3233 = ~n3231 & ~n3232;
  assign n3234 = pi80  & ~n4624;
  assign n3235 = pi208  & n4624;
  assign n3236 = ~n3234 & ~n3235;
  assign n3237 = ~n3233 & n3236;
  assign n3238 = ~n3230 & ~n3237;
  assign n3239 = n3223 & n3238;
  assign n3240 = ~n4744 & ~n3230;
  assign n3241 = n3223 & n3240;
  assign n3242 = ~n3237 & n3241;
  assign n3243 = ~n4744 & n3239;
  assign n3244 = ~n3211 & n3214;
  assign n3245 = n3233 & ~n3236;
  assign n3246 = ~n3230 & n3233;
  assign n3247 = ~n3236 & n3246;
  assign n3248 = ~n3230 & n3245;
  assign n3249 = ~n3226 & n3229;
  assign n3250 = n3218 & ~n3221;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = ~n4746 & ~n3249;
  assign n3253 = ~n3250 & n3252;
  assign n3254 = ~n4746 & n3251;
  assign n3255 = n3223 & ~n4747;
  assign n3256 = ~n3244 & ~n3255;
  assign n3257 = ~n4745 & n3256;
  assign n3258 = pi87  & ~n4624;
  assign n3259 = pi215  & n4624;
  assign n3260 = ~n3258 & ~n3259;
  assign n3261 = pi343  & ~n4696;
  assign n3262 = pi471  & n4696;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = n3260 & ~n3263;
  assign n3265 = pi342  & ~n4696;
  assign n3266 = pi470  & n4696;
  assign n3267 = ~n3265 & ~n3266;
  assign n3268 = pi86  & ~n4624;
  assign n3269 = pi214  & n4624;
  assign n3270 = ~n3268 & ~n3269;
  assign n3271 = ~n3267 & n3270;
  assign n3272 = ~n3264 & ~n3271;
  assign n3273 = pi85  & ~n4624;
  assign n3274 = pi213  & n4624;
  assign n3275 = ~n3273 & ~n3274;
  assign n3276 = pi341  & ~n4696;
  assign n3277 = pi469  & n4696;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = n3275 & ~n3278;
  assign n3280 = pi84  & ~n4624;
  assign n3281 = pi212  & n4624;
  assign n3282 = ~n3280 & ~n3281;
  assign n3283 = pi340  & ~n4696;
  assign n3284 = pi468  & n4696;
  assign n3285 = ~n3283 & ~n3284;
  assign n3286 = n3282 & ~n3285;
  assign n3287 = ~n3279 & ~n3286;
  assign n3288 = n3272 & n3287;
  assign n3289 = ~n3257 & n3288;
  assign n3290 = ~n3260 & n3263;
  assign n3291 = ~n3282 & n3285;
  assign n3292 = ~n3279 & n3291;
  assign n3293 = n3267 & ~n3270;
  assign n3294 = ~n3275 & n3278;
  assign n3295 = ~n3293 & ~n3294;
  assign n3296 = ~n3292 & n3295;
  assign n3297 = n3272 & ~n3296;
  assign n3298 = ~n3292 & ~n3294;
  assign n3299 = n3272 & ~n3298;
  assign n3300 = ~n3264 & n3293;
  assign n3301 = ~n3290 & ~n3300;
  assign n3302 = ~n3299 & n3301;
  assign n3303 = ~n3290 & ~n3297;
  assign n3304 = ~n3289 & ~n3300;
  assign n3305 = ~n3299 & n3304;
  assign n3306 = ~n3290 & n3305;
  assign n3307 = ~n3289 & n4748;
  assign n3308 = pi91  & ~n4624;
  assign n3309 = pi219  & n4624;
  assign n3310 = ~n3308 & ~n3309;
  assign n3311 = pi347  & ~n4696;
  assign n3312 = pi475  & n4696;
  assign n3313 = ~n3311 & ~n3312;
  assign n3314 = n3310 & ~n3313;
  assign n3315 = pi346  & ~n4696;
  assign n3316 = pi474  & n4696;
  assign n3317 = ~n3315 & ~n3316;
  assign n3318 = pi90  & ~n4624;
  assign n3319 = pi218  & n4624;
  assign n3320 = ~n3318 & ~n3319;
  assign n3321 = ~n3317 & n3320;
  assign n3322 = ~n3314 & ~n3321;
  assign n3323 = pi89  & ~n4624;
  assign n3324 = pi217  & n4624;
  assign n3325 = ~n3323 & ~n3324;
  assign n3326 = pi345  & ~n4696;
  assign n3327 = pi473  & n4696;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = n3325 & ~n3328;
  assign n3330 = pi344  & ~n4696;
  assign n3331 = pi472  & n4696;
  assign n3332 = ~n3330 & ~n3331;
  assign n3333 = pi88  & ~n4624;
  assign n3334 = pi216  & n4624;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = ~n3332 & n3335;
  assign n3337 = ~n3329 & ~n3336;
  assign n3338 = n3322 & n3337;
  assign n3339 = ~n4749 & n3338;
  assign n3340 = ~n3310 & n3313;
  assign n3341 = n3332 & ~n3335;
  assign n3342 = ~n3329 & n3341;
  assign n3343 = ~n3325 & n3328;
  assign n3344 = n3317 & ~n3320;
  assign n3345 = ~n3343 & ~n3344;
  assign n3346 = ~n3342 & ~n3343;
  assign n3347 = ~n3344 & n3346;
  assign n3348 = ~n3342 & n3345;
  assign n3349 = n3322 & ~n4750;
  assign n3350 = ~n3340 & ~n3349;
  assign n3351 = ~n3339 & n3350;
  assign n3352 = pi95  & ~n4624;
  assign n3353 = pi223  & n4624;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355 = pi351  & ~n4696;
  assign n3356 = pi479  & n4696;
  assign n3357 = ~n3355 & ~n3356;
  assign n3358 = n3354 & ~n3357;
  assign n3359 = pi350  & ~n4696;
  assign n3360 = pi478  & n4696;
  assign n3361 = ~n3359 & ~n3360;
  assign n3362 = pi94  & ~n4624;
  assign n3363 = pi222  & n4624;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = ~n3361 & n3364;
  assign n3366 = ~n3358 & ~n3365;
  assign n3367 = pi93  & ~n4624;
  assign n3368 = pi221  & n4624;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = pi349  & ~n4696;
  assign n3371 = pi477  & n4696;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = n3369 & ~n3372;
  assign n3374 = pi92  & ~n4624;
  assign n3375 = pi220  & n4624;
  assign n3376 = ~n3374 & ~n3375;
  assign n3377 = pi348  & ~n4696;
  assign n3378 = pi476  & n4696;
  assign n3379 = ~n3377 & ~n3378;
  assign n3380 = n3376 & ~n3379;
  assign n3381 = ~n3373 & ~n3380;
  assign n3382 = n3366 & n3381;
  assign n3383 = ~n3351 & n3382;
  assign n3384 = ~n3354 & n3357;
  assign n3385 = ~n3376 & n3379;
  assign n3386 = ~n3373 & n3385;
  assign n3387 = n3361 & ~n3364;
  assign n3388 = ~n3369 & n3372;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = ~n3386 & n3389;
  assign n3391 = n3366 & ~n3390;
  assign n3392 = ~n3386 & ~n3388;
  assign n3393 = n3366 & ~n3392;
  assign n3394 = ~n3358 & n3387;
  assign n3395 = ~n3384 & ~n3394;
  assign n3396 = ~n3393 & n3395;
  assign n3397 = ~n3384 & ~n3391;
  assign n3398 = ~n3383 & ~n3394;
  assign n3399 = ~n3393 & n3398;
  assign n3400 = ~n3384 & n3399;
  assign n3401 = ~n3383 & n4751;
  assign n3402 = pi99  & ~n4624;
  assign n3403 = pi227  & n4624;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = pi355  & ~n4696;
  assign n3406 = pi483  & n4696;
  assign n3407 = ~n3405 & ~n3406;
  assign n3408 = n3404 & ~n3407;
  assign n3409 = pi354  & ~n4696;
  assign n3410 = pi482  & n4696;
  assign n3411 = ~n3409 & ~n3410;
  assign n3412 = pi98  & ~n4624;
  assign n3413 = pi226  & n4624;
  assign n3414 = ~n3412 & ~n3413;
  assign n3415 = ~n3411 & n3414;
  assign n3416 = ~n3408 & ~n3415;
  assign n3417 = pi97  & ~n4624;
  assign n3418 = pi225  & n4624;
  assign n3419 = ~n3417 & ~n3418;
  assign n3420 = pi353  & ~n4696;
  assign n3421 = pi481  & n4696;
  assign n3422 = ~n3420 & ~n3421;
  assign n3423 = n3419 & ~n3422;
  assign n3424 = pi352  & ~n4696;
  assign n3425 = pi480  & n4696;
  assign n3426 = ~n3424 & ~n3425;
  assign n3427 = pi96  & ~n4624;
  assign n3428 = pi224  & n4624;
  assign n3429 = ~n3427 & ~n3428;
  assign n3430 = ~n3426 & n3429;
  assign n3431 = ~n3423 & ~n3430;
  assign n3432 = n3416 & n3431;
  assign n3433 = ~n4752 & ~n3423;
  assign n3434 = n3416 & n3433;
  assign n3435 = ~n3430 & n3434;
  assign n3436 = ~n4752 & n3432;
  assign n3437 = ~n3404 & n3407;
  assign n3438 = n3426 & ~n3429;
  assign n3439 = ~n3423 & n3426;
  assign n3440 = ~n3429 & n3439;
  assign n3441 = ~n3423 & n3438;
  assign n3442 = ~n3419 & n3422;
  assign n3443 = n3411 & ~n3414;
  assign n3444 = ~n3442 & ~n3443;
  assign n3445 = ~n4754 & ~n3442;
  assign n3446 = ~n3443 & n3445;
  assign n3447 = ~n4754 & n3444;
  assign n3448 = n3416 & ~n4755;
  assign n3449 = ~n3437 & ~n3448;
  assign n3450 = ~n4753 & n3449;
  assign n3451 = pi103  & ~n4624;
  assign n3452 = pi231  & n4624;
  assign n3453 = ~n3451 & ~n3452;
  assign n3454 = pi359  & ~n4696;
  assign n3455 = pi487  & n4696;
  assign n3456 = ~n3454 & ~n3455;
  assign n3457 = n3453 & ~n3456;
  assign n3458 = pi358  & ~n4696;
  assign n3459 = pi486  & n4696;
  assign n3460 = ~n3458 & ~n3459;
  assign n3461 = pi102  & ~n4624;
  assign n3462 = pi230  & n4624;
  assign n3463 = ~n3461 & ~n3462;
  assign n3464 = ~n3460 & n3463;
  assign n3465 = ~n3457 & ~n3464;
  assign n3466 = pi101  & ~n4624;
  assign n3467 = pi229  & n4624;
  assign n3468 = ~n3466 & ~n3467;
  assign n3469 = pi357  & ~n4696;
  assign n3470 = pi485  & n4696;
  assign n3471 = ~n3469 & ~n3470;
  assign n3472 = n3468 & ~n3471;
  assign n3473 = pi100  & ~n4624;
  assign n3474 = pi228  & n4624;
  assign n3475 = ~n3473 & ~n3474;
  assign n3476 = pi356  & ~n4696;
  assign n3477 = pi484  & n4696;
  assign n3478 = ~n3476 & ~n3477;
  assign n3479 = n3475 & ~n3478;
  assign n3480 = ~n3472 & ~n3479;
  assign n3481 = n3465 & n3480;
  assign n3482 = ~n3450 & n3481;
  assign n3483 = ~n3453 & n3456;
  assign n3484 = ~n3475 & n3478;
  assign n3485 = ~n3472 & n3484;
  assign n3486 = n3460 & ~n3463;
  assign n3487 = ~n3468 & n3471;
  assign n3488 = ~n3486 & ~n3487;
  assign n3489 = ~n3485 & n3488;
  assign n3490 = n3465 & ~n3489;
  assign n3491 = ~n3485 & ~n3487;
  assign n3492 = n3465 & ~n3491;
  assign n3493 = ~n3457 & n3486;
  assign n3494 = ~n3483 & ~n3493;
  assign n3495 = ~n3492 & n3494;
  assign n3496 = ~n3483 & ~n3490;
  assign n3497 = ~n3482 & ~n3493;
  assign n3498 = ~n3492 & n3497;
  assign n3499 = ~n3483 & n3498;
  assign n3500 = ~n3482 & n4756;
  assign n3501 = pi107  & ~n4624;
  assign n3502 = pi235  & n4624;
  assign n3503 = ~n3501 & ~n3502;
  assign n3504 = pi363  & ~n4696;
  assign n3505 = pi491  & n4696;
  assign n3506 = ~n3504 & ~n3505;
  assign n3507 = n3503 & ~n3506;
  assign n3508 = pi362  & ~n4696;
  assign n3509 = pi490  & n4696;
  assign n3510 = ~n3508 & ~n3509;
  assign n3511 = pi106  & ~n4624;
  assign n3512 = pi234  & n4624;
  assign n3513 = ~n3511 & ~n3512;
  assign n3514 = ~n3510 & n3513;
  assign n3515 = ~n3507 & ~n3514;
  assign n3516 = pi105  & ~n4624;
  assign n3517 = pi233  & n4624;
  assign n3518 = ~n3516 & ~n3517;
  assign n3519 = pi361  & ~n4696;
  assign n3520 = pi489  & n4696;
  assign n3521 = ~n3519 & ~n3520;
  assign n3522 = n3518 & ~n3521;
  assign n3523 = pi360  & ~n4696;
  assign n3524 = pi488  & n4696;
  assign n3525 = ~n3523 & ~n3524;
  assign n3526 = pi104  & ~n4624;
  assign n3527 = pi232  & n4624;
  assign n3528 = ~n3526 & ~n3527;
  assign n3529 = ~n3525 & n3528;
  assign n3530 = ~n3522 & ~n3529;
  assign n3531 = n3515 & n3530;
  assign n3532 = ~n4757 & n3531;
  assign n3533 = ~n3503 & n3506;
  assign n3534 = n3525 & ~n3528;
  assign n3535 = ~n3522 & n3534;
  assign n3536 = ~n3518 & n3521;
  assign n3537 = n3510 & ~n3513;
  assign n3538 = ~n3536 & ~n3537;
  assign n3539 = ~n3535 & ~n3536;
  assign n3540 = ~n3537 & n3539;
  assign n3541 = ~n3535 & n3538;
  assign n3542 = n3515 & ~n4758;
  assign n3543 = ~n3533 & ~n3542;
  assign n3544 = ~n3532 & n3543;
  assign n3545 = pi111  & ~n4624;
  assign n3546 = pi239  & n4624;
  assign n3547 = ~n3545 & ~n3546;
  assign n3548 = pi367  & ~n4696;
  assign n3549 = pi495  & n4696;
  assign n3550 = ~n3548 & ~n3549;
  assign n3551 = n3547 & ~n3550;
  assign n3552 = pi366  & ~n4696;
  assign n3553 = pi494  & n4696;
  assign n3554 = ~n3552 & ~n3553;
  assign n3555 = pi110  & ~n4624;
  assign n3556 = pi238  & n4624;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = ~n3554 & n3557;
  assign n3559 = ~n3551 & ~n3558;
  assign n3560 = pi109  & ~n4624;
  assign n3561 = pi237  & n4624;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = pi365  & ~n4696;
  assign n3564 = pi493  & n4696;
  assign n3565 = ~n3563 & ~n3564;
  assign n3566 = n3562 & ~n3565;
  assign n3567 = pi108  & ~n4624;
  assign n3568 = pi236  & n4624;
  assign n3569 = ~n3567 & ~n3568;
  assign n3570 = pi364  & ~n4696;
  assign n3571 = pi492  & n4696;
  assign n3572 = ~n3570 & ~n3571;
  assign n3573 = n3569 & ~n3572;
  assign n3574 = ~n3566 & ~n3573;
  assign n3575 = n3559 & n3574;
  assign n3576 = ~n3544 & n3575;
  assign n3577 = ~n3547 & n3550;
  assign n3578 = ~n3569 & n3572;
  assign n3579 = ~n3566 & n3578;
  assign n3580 = n3554 & ~n3557;
  assign n3581 = ~n3562 & n3565;
  assign n3582 = ~n3580 & ~n3581;
  assign n3583 = ~n3579 & n3582;
  assign n3584 = n3559 & ~n3583;
  assign n3585 = ~n3579 & ~n3581;
  assign n3586 = n3559 & ~n3585;
  assign n3587 = ~n3551 & n3580;
  assign n3588 = ~n3577 & ~n3587;
  assign n3589 = ~n3586 & n3588;
  assign n3590 = ~n3577 & ~n3584;
  assign n3591 = ~n3576 & ~n3587;
  assign n3592 = ~n3586 & n3591;
  assign n3593 = ~n3577 & n3592;
  assign n3594 = ~n3576 & n4759;
  assign n3595 = pi115  & ~n4624;
  assign n3596 = pi243  & n4624;
  assign n3597 = ~n3595 & ~n3596;
  assign n3598 = pi371  & ~n4696;
  assign n3599 = pi499  & n4696;
  assign n3600 = ~n3598 & ~n3599;
  assign n3601 = n3597 & ~n3600;
  assign n3602 = pi370  & ~n4696;
  assign n3603 = pi498  & n4696;
  assign n3604 = ~n3602 & ~n3603;
  assign n3605 = pi114  & ~n4624;
  assign n3606 = pi242  & n4624;
  assign n3607 = ~n3605 & ~n3606;
  assign n3608 = ~n3604 & n3607;
  assign n3609 = ~n3601 & ~n3608;
  assign n3610 = pi113  & ~n4624;
  assign n3611 = pi241  & n4624;
  assign n3612 = ~n3610 & ~n3611;
  assign n3613 = pi369  & ~n4696;
  assign n3614 = pi497  & n4696;
  assign n3615 = ~n3613 & ~n3614;
  assign n3616 = n3612 & ~n3615;
  assign n3617 = pi368  & ~n4696;
  assign n3618 = pi496  & n4696;
  assign n3619 = ~n3617 & ~n3618;
  assign n3620 = pi112  & ~n4624;
  assign n3621 = pi240  & n4624;
  assign n3622 = ~n3620 & ~n3621;
  assign n3623 = ~n3619 & n3622;
  assign n3624 = ~n3616 & ~n3623;
  assign n3625 = n3609 & n3624;
  assign n3626 = ~n4760 & ~n3616;
  assign n3627 = n3609 & n3626;
  assign n3628 = ~n3623 & n3627;
  assign n3629 = ~n4760 & n3625;
  assign n3630 = ~n3597 & n3600;
  assign n3631 = n3619 & ~n3622;
  assign n3632 = ~n3616 & n3619;
  assign n3633 = ~n3622 & n3632;
  assign n3634 = ~n3616 & n3631;
  assign n3635 = ~n3612 & n3615;
  assign n3636 = n3604 & ~n3607;
  assign n3637 = ~n3635 & ~n3636;
  assign n3638 = ~n4762 & ~n3635;
  assign n3639 = ~n3636 & n3638;
  assign n3640 = ~n4762 & n3637;
  assign n3641 = n3609 & ~n4763;
  assign n3642 = ~n3630 & ~n3641;
  assign n3643 = ~n4761 & n3642;
  assign n3644 = pi119  & ~n4624;
  assign n3645 = pi247  & n4624;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = pi375  & ~n4696;
  assign n3648 = pi503  & n4696;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650 = n3646 & ~n3649;
  assign n3651 = pi374  & ~n4696;
  assign n3652 = pi502  & n4696;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = pi118  & ~n4624;
  assign n3655 = pi246  & n4624;
  assign n3656 = ~n3654 & ~n3655;
  assign n3657 = ~n3653 & n3656;
  assign n3658 = ~n3650 & ~n3657;
  assign n3659 = pi117  & ~n4624;
  assign n3660 = pi245  & n4624;
  assign n3661 = ~n3659 & ~n3660;
  assign n3662 = pi373  & ~n4696;
  assign n3663 = pi501  & n4696;
  assign n3664 = ~n3662 & ~n3663;
  assign n3665 = n3661 & ~n3664;
  assign n3666 = pi116  & ~n4624;
  assign n3667 = pi244  & n4624;
  assign n3668 = ~n3666 & ~n3667;
  assign n3669 = pi372  & ~n4696;
  assign n3670 = pi500  & n4696;
  assign n3671 = ~n3669 & ~n3670;
  assign n3672 = n3668 & ~n3671;
  assign n3673 = ~n3665 & ~n3672;
  assign n3674 = n3658 & n3673;
  assign n3675 = ~n3643 & n3674;
  assign n3676 = ~n3646 & n3649;
  assign n3677 = ~n3668 & n3671;
  assign n3678 = ~n3665 & n3671;
  assign n3679 = ~n3668 & n3678;
  assign n3680 = ~n3665 & n3677;
  assign n3681 = n3653 & ~n3656;
  assign n3682 = ~n3661 & n3664;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = ~n4764 & n3683;
  assign n3685 = n3658 & ~n3684;
  assign n3686 = ~n4764 & ~n3682;
  assign n3687 = n3658 & ~n3686;
  assign n3688 = ~n3650 & n3681;
  assign n3689 = ~n3676 & ~n3688;
  assign n3690 = ~n3687 & n3689;
  assign n3691 = ~n3676 & ~n3685;
  assign n3692 = ~n3675 & ~n3688;
  assign n3693 = ~n3687 & n3692;
  assign n3694 = ~n3676 & n3693;
  assign n3695 = ~n3675 & n4765;
  assign n3696 = pi123  & ~n4624;
  assign n3697 = pi251  & n4624;
  assign n3698 = ~n3696 & ~n3697;
  assign n3699 = pi379  & ~n4696;
  assign n3700 = pi507  & n4696;
  assign n3701 = ~n3699 & ~n3700;
  assign n3702 = n3698 & ~n3701;
  assign n3703 = pi378  & ~n4696;
  assign n3704 = pi506  & n4696;
  assign n3705 = ~n3703 & ~n3704;
  assign n3706 = pi122  & ~n4624;
  assign n3707 = pi250  & n4624;
  assign n3708 = ~n3706 & ~n3707;
  assign n3709 = ~n3705 & n3708;
  assign n3710 = ~n3702 & ~n3709;
  assign n3711 = pi121  & ~n4624;
  assign n3712 = pi249  & n4624;
  assign n3713 = ~n3711 & ~n3712;
  assign n3714 = pi377  & ~n4696;
  assign n3715 = pi505  & n4696;
  assign n3716 = ~n3714 & ~n3715;
  assign n3717 = n3713 & ~n3716;
  assign n3718 = pi376  & ~n4696;
  assign n3719 = pi504  & n4696;
  assign n3720 = ~n3718 & ~n3719;
  assign n3721 = pi120  & ~n4624;
  assign n3722 = pi248  & n4624;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = ~n3720 & n3723;
  assign n3725 = ~n3717 & ~n3724;
  assign n3726 = n3710 & n3725;
  assign n3727 = ~n4766 & n3726;
  assign n3728 = ~n3698 & n3701;
  assign n3729 = n3720 & ~n3723;
  assign n3730 = ~n3717 & n3720;
  assign n3731 = ~n3723 & n3730;
  assign n3732 = ~n3717 & n3729;
  assign n3733 = ~n3713 & n3716;
  assign n3734 = n3705 & ~n3708;
  assign n3735 = ~n3733 & ~n3734;
  assign n3736 = ~n4767 & ~n3733;
  assign n3737 = ~n3734 & n3736;
  assign n3738 = ~n4767 & n3735;
  assign n3739 = n3710 & ~n4768;
  assign n3740 = ~n3728 & ~n3739;
  assign n3741 = ~n3727 & n3740;
  assign n3742 = pi126  & ~n4624;
  assign n3743 = pi254  & n4624;
  assign n3744 = ~n3742 & ~n3743;
  assign n3745 = pi382  & ~n4696;
  assign n3746 = pi510  & n4696;
  assign n3747 = ~n3745 & ~n3746;
  assign n3748 = n3744 & ~n3747;
  assign n3749 = pi125  & ~n4624;
  assign n3750 = pi253  & n4624;
  assign n3751 = ~n3749 & ~n3750;
  assign n3752 = pi381  & ~n4696;
  assign n3753 = pi509  & n4696;
  assign n3754 = ~n3752 & ~n3753;
  assign n3755 = n3751 & ~n3754;
  assign n3756 = ~n3748 & ~n3755;
  assign n3757 = ~pi511  & n2205;
  assign n3758 = pi383  & ~n3757;
  assign n3759 = ~pi511  & ~n2195;
  assign n3760 = pi383  & ~n3759;
  assign n3761 = pi383  & pi511 ;
  assign n3762 = ~pi255  & n1420;
  assign n3763 = pi127  & ~n3762;
  assign n3764 = ~pi255  & ~n1410;
  assign n3765 = pi127  & ~n3764;
  assign n3766 = pi127  & pi255 ;
  assign n3767 = ~n4769 & n4770;
  assign n3768 = pi124  & ~n4624;
  assign n3769 = pi252  & n4624;
  assign n3770 = ~n3768 & ~n3769;
  assign n3771 = pi380  & ~n4696;
  assign n3772 = pi508  & n4696;
  assign n3773 = ~n3771 & ~n3772;
  assign n3774 = n3770 & ~n3773;
  assign n3775 = ~n3767 & ~n3774;
  assign n3776 = n3756 & ~n3767;
  assign n3777 = ~n3774 & n3776;
  assign n3778 = n3756 & n3775;
  assign n3779 = ~n3741 & n4771;
  assign n3780 = ~n3770 & n3773;
  assign n3781 = ~n3751 & n3754;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = n3756 & ~n3782;
  assign n3784 = n4769 & ~n4770;
  assign n3785 = ~n3744 & n3747;
  assign n3786 = ~n3784 & ~n3785;
  assign n3787 = ~n3783 & n3786;
  assign n3788 = ~n3767 & ~n3787;
  assign n3789 = ~n3783 & ~n3785;
  assign n3790 = ~n3767 & ~n3789;
  assign n3791 = ~n3779 & ~n3790;
  assign n3792 = ~n3784 & n3791;
  assign n3793 = ~n3779 & ~n3788;
  assign n3794 = ~n2341 & po129 ;
  assign n3795 = ~n2344 & ~po129 ;
  assign n3796 = ~n3794 & ~n3795;
  assign n3797 = n2337 & ~po129 ;
  assign n3798 = n2334 & po129 ;
  assign n3799 = ~n2334 & po129 ;
  assign n3800 = ~n2337 & ~po129 ;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = ~n3797 & ~n3798;
  assign n3803 = n2326 & ~po129 ;
  assign n3804 = n2329 & po129 ;
  assign n3805 = ~n2329 & po129 ;
  assign n3806 = ~n2326 & ~po129 ;
  assign n3807 = ~n3805 & ~n3806;
  assign n3808 = ~n3803 & ~n3804;
  assign n3809 = n2318 & ~po129 ;
  assign n3810 = n2321 & po129 ;
  assign n3811 = ~n2321 & po129 ;
  assign n3812 = ~n2318 & ~po129 ;
  assign n3813 = ~n3811 & ~n3812;
  assign n3814 = ~n3809 & ~n3810;
  assign n3815 = ~n2315 & po129 ;
  assign n3816 = ~n2368 & ~po129 ;
  assign n3817 = ~n3815 & ~n3816;
  assign n3818 = ~n2312 & po129 ;
  assign n3819 = ~n2379 & ~po129 ;
  assign n3820 = ~n3818 & ~n3819;
  assign n3821 = ~n2390 & po129 ;
  assign n3822 = ~n2395 & ~po129 ;
  assign n3823 = ~n3821 & ~n3822;
  assign n3824 = n2305 & ~po129 ;
  assign n3825 = n2308 & po129 ;
  assign n3826 = ~n2308 & po129 ;
  assign n3827 = ~n2305 & ~po129 ;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = ~n3824 & ~n3825;
  assign n3830 = n2406 & ~po129 ;
  assign n3831 = n2409 & po129 ;
  assign n3832 = ~n2409 & po129 ;
  assign n3833 = ~n2406 & ~po129 ;
  assign n3834 = ~n3832 & ~n3833;
  assign n3835 = ~n3830 & ~n3831;
  assign n3836 = n2416 & ~po129 ;
  assign n3837 = n2419 & po129 ;
  assign n3838 = ~n2419 & po129 ;
  assign n3839 = ~n2416 & ~po129 ;
  assign n3840 = ~n3838 & ~n3839;
  assign n3841 = ~n3836 & ~n3837;
  assign n3842 = n2298 & ~po129 ;
  assign n3843 = n2301 & po129 ;
  assign n3844 = ~n2301 & po129 ;
  assign n3845 = ~n2298 & ~po129 ;
  assign n3846 = ~n3844 & ~n3845;
  assign n3847 = ~n3842 & ~n3843;
  assign n3848 = n2290 & ~po129 ;
  assign n3849 = n2293 & po129 ;
  assign n3850 = ~n2293 & po129 ;
  assign n3851 = ~n2290 & ~po129 ;
  assign n3852 = ~n3850 & ~n3851;
  assign n3853 = ~n3848 & ~n3849;
  assign n3854 = n2282 & ~po129 ;
  assign n3855 = n2285 & po129 ;
  assign n3856 = ~n2285 & po129 ;
  assign n3857 = ~n2282 & ~po129 ;
  assign n3858 = ~n3856 & ~n3857;
  assign n3859 = ~n3854 & ~n3855;
  assign n3860 = n2275 & ~po129 ;
  assign n3861 = n2278 & po129 ;
  assign n3862 = ~n2278 & po129 ;
  assign n3863 = ~n2275 & ~po129 ;
  assign n3864 = ~n3862 & ~n3863;
  assign n3865 = ~n3860 & ~n3861;
  assign n3866 = n2450 & ~po129 ;
  assign n3867 = n2453 & po129 ;
  assign n3868 = ~n2453 & po129 ;
  assign n3869 = ~n2450 & ~po129 ;
  assign n3870 = ~n3868 & ~n3869;
  assign n3871 = ~n3866 & ~n3867;
  assign n3872 = n2460 & ~po129 ;
  assign n3873 = n2463 & po129 ;
  assign n3874 = ~n2463 & po129 ;
  assign n3875 = ~n2460 & ~po129 ;
  assign n3876 = ~n3874 & ~n3875;
  assign n3877 = ~n3872 & ~n3873;
  assign n3878 = n2474 & ~po129 ;
  assign n3879 = n2477 & po129 ;
  assign n3880 = ~n2477 & po129 ;
  assign n3881 = ~n2474 & ~po129 ;
  assign n3882 = ~n3880 & ~n3881;
  assign n3883 = ~n3878 & ~n3879;
  assign n3884 = n2268 & ~po129 ;
  assign n3885 = n2271 & po129 ;
  assign n3886 = ~n2271 & po129 ;
  assign n3887 = ~n2268 & ~po129 ;
  assign n3888 = ~n3886 & ~n3887;
  assign n3889 = ~n3884 & ~n3885;
  assign n3890 = n2260 & ~po129 ;
  assign n3891 = n2263 & po129 ;
  assign n3892 = ~n2263 & po129 ;
  assign n3893 = ~n2260 & ~po129 ;
  assign n3894 = ~n3892 & ~n3893;
  assign n3895 = ~n3890 & ~n3891;
  assign n3896 = n2252 & ~po129 ;
  assign n3897 = n2255 & po129 ;
  assign n3898 = ~n2255 & po129 ;
  assign n3899 = ~n2252 & ~po129 ;
  assign n3900 = ~n3898 & ~n3899;
  assign n3901 = ~n3896 & ~n3897;
  assign n3902 = n2244 & ~po129 ;
  assign n3903 = n2247 & po129 ;
  assign n3904 = ~n2247 & po129 ;
  assign n3905 = ~n2244 & ~po129 ;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = ~n3902 & ~n3903;
  assign n3908 = n2237 & ~po129 ;
  assign n3909 = n2240 & po129 ;
  assign n3910 = ~n2240 & po129 ;
  assign n3911 = ~n2237 & ~po129 ;
  assign n3912 = ~n3910 & ~n3911;
  assign n3913 = ~n3908 & ~n3909;
  assign n3914 = n2506 & ~po129 ;
  assign n3915 = n2509 & po129 ;
  assign n3916 = ~n2509 & po129 ;
  assign n3917 = ~n2506 & ~po129 ;
  assign n3918 = ~n3916 & ~n3917;
  assign n3919 = ~n3914 & ~n3915;
  assign n3920 = n2516 & ~po129 ;
  assign n3921 = n2519 & po129 ;
  assign n3922 = ~n2519 & po129 ;
  assign n3923 = ~n2516 & ~po129 ;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = ~n3920 & ~n3921;
  assign n3926 = n2530 & ~po129 ;
  assign n3927 = n2533 & po129 ;
  assign n3928 = ~n2533 & po129 ;
  assign n3929 = ~n2530 & ~po129 ;
  assign n3930 = ~n3928 & ~n3929;
  assign n3931 = ~n3926 & ~n3927;
  assign n3932 = n2230 & ~po129 ;
  assign n3933 = n2233 & po129 ;
  assign n3934 = ~n2233 & po129 ;
  assign n3935 = ~n2230 & ~po129 ;
  assign n3936 = ~n3934 & ~n3935;
  assign n3937 = ~n3932 & ~n3933;
  assign n3938 = n2222 & ~po129 ;
  assign n3939 = n2225 & po129 ;
  assign n3940 = ~n2225 & po129 ;
  assign n3941 = ~n2222 & ~po129 ;
  assign n3942 = ~n3940 & ~n3941;
  assign n3943 = ~n3938 & ~n3939;
  assign n3944 = n2214 & ~po129 ;
  assign n3945 = n2217 & po129 ;
  assign n3946 = ~n2217 & po129 ;
  assign n3947 = ~n2214 & ~po129 ;
  assign n3948 = ~n3946 & ~n3947;
  assign n3949 = ~n3944 & ~n3945;
  assign n3950 = n1425 & ~po129 ;
  assign n3951 = n2210 & po129 ;
  assign n3952 = ~n2210 & po129 ;
  assign n3953 = ~n1425 & ~po129 ;
  assign n3954 = ~n3952 & ~n3953;
  assign n3955 = ~n3950 & ~n3951;
  assign n3956 = n2560 & ~po129 ;
  assign n3957 = n2563 & po129 ;
  assign n3958 = ~n2563 & po129 ;
  assign n3959 = ~n2560 & ~po129 ;
  assign n3960 = ~n3958 & ~n3959;
  assign n3961 = ~n3956 & ~n3957;
  assign n3962 = n2570 & ~po129 ;
  assign n3963 = n2573 & po129 ;
  assign n3964 = ~n2573 & po129 ;
  assign n3965 = ~n2570 & ~po129 ;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = ~n3962 & ~n3963;
  assign n3968 = n2584 & ~po129 ;
  assign n3969 = n2587 & po129 ;
  assign n3970 = ~n2587 & po129 ;
  assign n3971 = ~n2584 & ~po129 ;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = ~n3968 & ~n3969;
  assign n3974 = n2642 & ~po129 ;
  assign n3975 = n2639 & po129 ;
  assign n3976 = ~n2639 & po129 ;
  assign n3977 = ~n2642 & ~po129 ;
  assign n3978 = ~n3976 & ~n3977;
  assign n3979 = ~n3974 & ~n3975;
  assign n3980 = n2593 & ~po129 ;
  assign n3981 = n2596 & po129 ;
  assign n3982 = ~n2596 & po129 ;
  assign n3983 = ~n2593 & ~po129 ;
  assign n3984 = ~n3982 & ~n3983;
  assign n3985 = ~n3980 & ~n3981;
  assign n3986 = n2610 & ~po129 ;
  assign n3987 = n2607 & po129 ;
  assign n3988 = ~n2607 & po129 ;
  assign n3989 = ~n2610 & ~po129 ;
  assign n3990 = ~n3988 & ~n3989;
  assign n3991 = ~n3986 & ~n3987;
  assign n3992 = n2600 & ~po129 ;
  assign n3993 = n2603 & po129 ;
  assign n3994 = ~n2603 & po129 ;
  assign n3995 = ~n2600 & ~po129 ;
  assign n3996 = ~n3994 & ~n3995;
  assign n3997 = ~n3992 & ~n3993;
  assign n3998 = n2647 & ~po129 ;
  assign n3999 = n2650 & po129 ;
  assign n4000 = ~n2650 & po129 ;
  assign n4001 = ~n2647 & ~po129 ;
  assign n4002 = ~n4000 & ~n4001;
  assign n4003 = ~n3998 & ~n3999;
  assign n4004 = n2623 & ~po129 ;
  assign n4005 = n2626 & po129 ;
  assign n4006 = ~n2626 & po129 ;
  assign n4007 = ~n2623 & ~po129 ;
  assign n4008 = ~n4006 & ~n4007;
  assign n4009 = ~n4004 & ~n4005;
  assign n4010 = n2633 & ~po129 ;
  assign n4011 = n2630 & po129 ;
  assign n4012 = ~n2630 & po129 ;
  assign n4013 = ~n2633 & ~po129 ;
  assign n4014 = ~n4012 & ~n4013;
  assign n4015 = ~n4010 & ~n4011;
  assign n4016 = n2616 & ~po129 ;
  assign n4017 = n2619 & po129 ;
  assign n4018 = ~n2619 & po129 ;
  assign n4019 = ~n2616 & ~po129 ;
  assign n4020 = ~n4018 & ~n4019;
  assign n4021 = ~n4016 & ~n4017;
  assign n4022 = n2765 & ~po129 ;
  assign n4023 = n2768 & po129 ;
  assign n4024 = ~n2768 & po129 ;
  assign n4025 = ~n2765 & ~po129 ;
  assign n4026 = ~n4024 & ~n4025;
  assign n4027 = ~n4022 & ~n4023;
  assign n4028 = n2758 & ~po129 ;
  assign n4029 = n2761 & po129 ;
  assign n4030 = ~n2761 & po129 ;
  assign n4031 = ~n2758 & ~po129 ;
  assign n4032 = ~n4030 & ~n4031;
  assign n4033 = ~n4028 & ~n4029;
  assign n4034 = n2750 & ~po129 ;
  assign n4035 = n2753 & po129 ;
  assign n4036 = ~n2753 & po129 ;
  assign n4037 = ~n2750 & ~po129 ;
  assign n4038 = ~n4036 & ~n4037;
  assign n4039 = ~n4034 & ~n4035;
  assign n4040 = n2743 & ~po129 ;
  assign n4041 = n2746 & po129 ;
  assign n4042 = ~n2746 & po129 ;
  assign n4043 = ~n2743 & ~po129 ;
  assign n4044 = ~n4042 & ~n4043;
  assign n4045 = ~n4040 & ~n4041;
  assign n4046 = n2731 & ~po129 ;
  assign n4047 = n2734 & po129 ;
  assign n4048 = ~n2734 & po129 ;
  assign n4049 = ~n2731 & ~po129 ;
  assign n4050 = ~n4048 & ~n4049;
  assign n4051 = ~n4046 & ~n4047;
  assign n4052 = n2724 & ~po129 ;
  assign n4053 = n2727 & po129 ;
  assign n4054 = ~n2727 & po129 ;
  assign n4055 = ~n2724 & ~po129 ;
  assign n4056 = ~n4054 & ~n4055;
  assign n4057 = ~n4052 & ~n4053;
  assign n4058 = n2719 & ~po129 ;
  assign n4059 = n2716 & po129 ;
  assign n4060 = ~n2716 & po129 ;
  assign n4061 = ~n2719 & ~po129 ;
  assign n4062 = ~n4060 & ~n4061;
  assign n4063 = ~n4058 & ~n4059;
  assign n4064 = n2709 & ~po129 ;
  assign n4065 = n2712 & po129 ;
  assign n4066 = ~n2712 & po129 ;
  assign n4067 = ~n2709 & ~po129 ;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = ~n4064 & ~n4065;
  assign n4070 = n2871 & ~po129 ;
  assign n4071 = n2868 & po129 ;
  assign n4072 = ~n2868 & po129 ;
  assign n4073 = ~n2871 & ~po129 ;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = ~n4070 & ~n4071;
  assign n4076 = n2845 & ~po129 ;
  assign n4077 = n2848 & po129 ;
  assign n4078 = ~n2848 & po129 ;
  assign n4079 = ~n2845 & ~po129 ;
  assign n4080 = ~n4078 & ~n4079;
  assign n4081 = ~n4076 & ~n4077;
  assign n4082 = n2862 & ~po129 ;
  assign n4083 = n2859 & po129 ;
  assign n4084 = ~n2859 & po129 ;
  assign n4085 = ~n2862 & ~po129 ;
  assign n4086 = ~n4084 & ~n4085;
  assign n4087 = ~n4082 & ~n4083;
  assign n4088 = n2852 & ~po129 ;
  assign n4089 = n2855 & po129 ;
  assign n4090 = ~n2855 & po129 ;
  assign n4091 = ~n2852 & ~po129 ;
  assign n4092 = ~n4090 & ~n4091;
  assign n4093 = ~n4088 & ~n4089;
  assign n4094 = n2839 & ~po129 ;
  assign n4095 = n2836 & po129 ;
  assign n4096 = ~n2836 & po129 ;
  assign n4097 = ~n2839 & ~po129 ;
  assign n4098 = ~n4096 & ~n4097;
  assign n4099 = ~n4094 & ~n4095;
  assign n4100 = n2829 & ~po129 ;
  assign n4101 = n2832 & po129 ;
  assign n4102 = ~n2832 & po129 ;
  assign n4103 = ~n2829 & ~po129 ;
  assign n4104 = ~n4102 & ~n4103;
  assign n4105 = ~n4100 & ~n4101;
  assign n4106 = n2824 & ~po129 ;
  assign n4107 = n2821 & po129 ;
  assign n4108 = ~n2821 & po129 ;
  assign n4109 = ~n2824 & ~po129 ;
  assign n4110 = ~n4108 & ~n4109;
  assign n4111 = ~n4106 & ~n4107;
  assign n4112 = n2814 & ~po129 ;
  assign n4113 = n2817 & po129 ;
  assign n4114 = ~n2817 & po129 ;
  assign n4115 = ~n2814 & ~po129 ;
  assign n4116 = ~n4114 & ~n4115;
  assign n4117 = ~n4112 & ~n4113;
  assign n4118 = n2967 & ~po129 ;
  assign n4119 = n2970 & po129 ;
  assign n4120 = ~n2970 & po129 ;
  assign n4121 = ~n2967 & ~po129 ;
  assign n4122 = ~n4120 & ~n4121;
  assign n4123 = ~n4118 & ~n4119;
  assign n4124 = n2960 & ~po129 ;
  assign n4125 = n2963 & po129 ;
  assign n4126 = ~n2963 & po129 ;
  assign n4127 = ~n2960 & ~po129 ;
  assign n4128 = ~n4126 & ~n4127;
  assign n4129 = ~n4124 & ~n4125;
  assign n4130 = n2952 & ~po129 ;
  assign n4131 = n2955 & po129 ;
  assign n4132 = ~n2955 & po129 ;
  assign n4133 = ~n2952 & ~po129 ;
  assign n4134 = ~n4132 & ~n4133;
  assign n4135 = ~n4130 & ~n4131;
  assign n4136 = n2945 & ~po129 ;
  assign n4137 = n2948 & po129 ;
  assign n4138 = ~n2948 & po129 ;
  assign n4139 = ~n2945 & ~po129 ;
  assign n4140 = ~n4138 & ~n4139;
  assign n4141 = ~n4136 & ~n4137;
  assign n4142 = n2933 & ~po129 ;
  assign n4143 = n2936 & po129 ;
  assign n4144 = ~n2936 & po129 ;
  assign n4145 = ~n2933 & ~po129 ;
  assign n4146 = ~n4144 & ~n4145;
  assign n4147 = ~n4142 & ~n4143;
  assign n4148 = n2926 & ~po129 ;
  assign n4149 = n2929 & po129 ;
  assign n4150 = ~n2929 & po129 ;
  assign n4151 = ~n2926 & ~po129 ;
  assign n4152 = ~n4150 & ~n4151;
  assign n4153 = ~n4148 & ~n4149;
  assign n4154 = n2921 & ~po129 ;
  assign n4155 = n2918 & po129 ;
  assign n4156 = ~n2918 & po129 ;
  assign n4157 = ~n2921 & ~po129 ;
  assign n4158 = ~n4156 & ~n4157;
  assign n4159 = ~n4154 & ~n4155;
  assign n4160 = n2911 & ~po129 ;
  assign n4161 = n2914 & po129 ;
  assign n4162 = ~n2914 & po129 ;
  assign n4163 = ~n2911 & ~po129 ;
  assign n4164 = ~n4162 & ~n4163;
  assign n4165 = ~n4160 & ~n4161;
  assign n4166 = n3043 & ~po129 ;
  assign n4167 = n3040 & po129 ;
  assign n4168 = ~n3040 & po129 ;
  assign n4169 = ~n3043 & ~po129 ;
  assign n4170 = ~n4168 & ~n4169;
  assign n4171 = ~n4166 & ~n4167;
  assign n4172 = n3033 & ~po129 ;
  assign n4173 = n3036 & po129 ;
  assign n4174 = ~n3036 & po129 ;
  assign n4175 = ~n3033 & ~po129 ;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = ~n4172 & ~n4173;
  assign n4178 = n3028 & ~po129 ;
  assign n4179 = n3025 & po129 ;
  assign n4180 = ~n3025 & po129 ;
  assign n4181 = ~n3028 & ~po129 ;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = ~n4178 & ~n4179;
  assign n4184 = n3018 & ~po129 ;
  assign n4185 = n3021 & po129 ;
  assign n4186 = ~n3021 & po129 ;
  assign n4187 = ~n3018 & ~po129 ;
  assign n4188 = ~n4186 & ~n4187;
  assign n4189 = ~n4184 & ~n4185;
  assign n4190 = n3089 & ~po129 ;
  assign n4191 = n3092 & po129 ;
  assign n4192 = ~n3092 & po129 ;
  assign n4193 = ~n3089 & ~po129 ;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = ~n4190 & ~n4191;
  assign n4196 = n3082 & ~po129 ;
  assign n4197 = n3085 & po129 ;
  assign n4198 = ~n3085 & po129 ;
  assign n4199 = ~n3082 & ~po129 ;
  assign n4200 = ~n4198 & ~n4199;
  assign n4201 = ~n4196 & ~n4197;
  assign n4202 = n3077 & ~po129 ;
  assign n4203 = n3074 & po129 ;
  assign n4204 = ~n3074 & po129 ;
  assign n4205 = ~n3077 & ~po129 ;
  assign n4206 = ~n4204 & ~n4205;
  assign n4207 = ~n4202 & ~n4203;
  assign n4208 = n3067 & ~po129 ;
  assign n4209 = n3070 & po129 ;
  assign n4210 = ~n3070 & po129 ;
  assign n4211 = ~n3067 & ~po129 ;
  assign n4212 = ~n4210 & ~n4211;
  assign n4213 = ~n4208 & ~n4209;
  assign n4214 = n3142 & ~po129 ;
  assign n4215 = n3139 & po129 ;
  assign n4216 = ~n3139 & po129 ;
  assign n4217 = ~n3142 & ~po129 ;
  assign n4218 = ~n4216 & ~n4217;
  assign n4219 = ~n4214 & ~n4215;
  assign n4220 = n3132 & ~po129 ;
  assign n4221 = n3135 & po129 ;
  assign n4222 = ~n3135 & po129 ;
  assign n4223 = ~n3132 & ~po129 ;
  assign n4224 = ~n4222 & ~n4223;
  assign n4225 = ~n4220 & ~n4221;
  assign n4226 = n3127 & ~po129 ;
  assign n4227 = n3124 & po129 ;
  assign n4228 = ~n3124 & po129 ;
  assign n4229 = ~n3127 & ~po129 ;
  assign n4230 = ~n4228 & ~n4229;
  assign n4231 = ~n4226 & ~n4227;
  assign n4232 = n3117 & ~po129 ;
  assign n4233 = n3120 & po129 ;
  assign n4234 = ~n3120 & po129 ;
  assign n4235 = ~n3117 & ~po129 ;
  assign n4236 = ~n4234 & ~n4235;
  assign n4237 = ~n4232 & ~n4233;
  assign n4238 = n3183 & ~po129 ;
  assign n4239 = n3186 & po129 ;
  assign n4240 = ~n3186 & po129 ;
  assign n4241 = ~n3183 & ~po129 ;
  assign n4242 = ~n4240 & ~n4241;
  assign n4243 = ~n4238 & ~n4239;
  assign n4244 = n3176 & ~po129 ;
  assign n4245 = n3179 & po129 ;
  assign n4246 = ~n3179 & po129 ;
  assign n4247 = ~n3176 & ~po129 ;
  assign n4248 = ~n4246 & ~n4247;
  assign n4249 = ~n4244 & ~n4245;
  assign n4250 = n3171 & ~po129 ;
  assign n4251 = n3168 & po129 ;
  assign n4252 = ~n3168 & po129 ;
  assign n4253 = ~n3171 & ~po129 ;
  assign n4254 = ~n4252 & ~n4253;
  assign n4255 = ~n4250 & ~n4251;
  assign n4256 = n3161 & ~po129 ;
  assign n4257 = n3164 & po129 ;
  assign n4258 = ~n3164 & po129 ;
  assign n4259 = ~n3161 & ~po129 ;
  assign n4260 = ~n4258 & ~n4259;
  assign n4261 = ~n4256 & ~n4257;
  assign n4262 = n3236 & ~po129 ;
  assign n4263 = n3233 & po129 ;
  assign n4264 = ~n3233 & po129 ;
  assign n4265 = ~n3236 & ~po129 ;
  assign n4266 = ~n4264 & ~n4265;
  assign n4267 = ~n4262 & ~n4263;
  assign n4268 = n3226 & ~po129 ;
  assign n4269 = n3229 & po129 ;
  assign n4270 = ~n3229 & po129 ;
  assign n4271 = ~n3226 & ~po129 ;
  assign n4272 = ~n4270 & ~n4271;
  assign n4273 = ~n4268 & ~n4269;
  assign n4274 = n3221 & ~po129 ;
  assign n4275 = n3218 & po129 ;
  assign n4276 = ~n3218 & po129 ;
  assign n4277 = ~n3221 & ~po129 ;
  assign n4278 = ~n4276 & ~n4277;
  assign n4279 = ~n4274 & ~n4275;
  assign n4280 = n3211 & ~po129 ;
  assign n4281 = n3214 & po129 ;
  assign n4282 = ~n3214 & po129 ;
  assign n4283 = ~n3211 & ~po129 ;
  assign n4284 = ~n4282 & ~n4283;
  assign n4285 = ~n4280 & ~n4281;
  assign n4286 = n3282 & ~po129 ;
  assign n4287 = n3285 & po129 ;
  assign n4288 = ~n3285 & po129 ;
  assign n4289 = ~n3282 & ~po129 ;
  assign n4290 = ~n4288 & ~n4289;
  assign n4291 = ~n4286 & ~n4287;
  assign n4292 = n3275 & ~po129 ;
  assign n4293 = n3278 & po129 ;
  assign n4294 = ~n3278 & po129 ;
  assign n4295 = ~n3275 & ~po129 ;
  assign n4296 = ~n4294 & ~n4295;
  assign n4297 = ~n4292 & ~n4293;
  assign n4298 = n3270 & ~po129 ;
  assign n4299 = n3267 & po129 ;
  assign n4300 = ~n3267 & po129 ;
  assign n4301 = ~n3270 & ~po129 ;
  assign n4302 = ~n4300 & ~n4301;
  assign n4303 = ~n4298 & ~n4299;
  assign n4304 = n3260 & ~po129 ;
  assign n4305 = n3263 & po129 ;
  assign n4306 = ~n3263 & po129 ;
  assign n4307 = ~n3260 & ~po129 ;
  assign n4308 = ~n4306 & ~n4307;
  assign n4309 = ~n4304 & ~n4305;
  assign n4310 = n3335 & ~po129 ;
  assign n4311 = n3332 & po129 ;
  assign n4312 = ~n3332 & po129 ;
  assign n4313 = ~n3335 & ~po129 ;
  assign n4314 = ~n4312 & ~n4313;
  assign n4315 = ~n4310 & ~n4311;
  assign n4316 = n3325 & ~po129 ;
  assign n4317 = n3328 & po129 ;
  assign n4318 = ~n3328 & po129 ;
  assign n4319 = ~n3325 & ~po129 ;
  assign n4320 = ~n4318 & ~n4319;
  assign n4321 = ~n4316 & ~n4317;
  assign n4322 = n3320 & ~po129 ;
  assign n4323 = n3317 & po129 ;
  assign n4324 = ~n3317 & po129 ;
  assign n4325 = ~n3320 & ~po129 ;
  assign n4326 = ~n4324 & ~n4325;
  assign n4327 = ~n4322 & ~n4323;
  assign n4328 = n3310 & ~po129 ;
  assign n4329 = n3313 & po129 ;
  assign n4330 = ~n3313 & po129 ;
  assign n4331 = ~n3310 & ~po129 ;
  assign n4332 = ~n4330 & ~n4331;
  assign n4333 = ~n4328 & ~n4329;
  assign n4334 = n3376 & ~po129 ;
  assign n4335 = n3379 & po129 ;
  assign n4336 = ~n3379 & po129 ;
  assign n4337 = ~n3376 & ~po129 ;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = ~n4334 & ~n4335;
  assign n4340 = n3369 & ~po129 ;
  assign n4341 = n3372 & po129 ;
  assign n4342 = ~n3372 & po129 ;
  assign n4343 = ~n3369 & ~po129 ;
  assign n4344 = ~n4342 & ~n4343;
  assign n4345 = ~n4340 & ~n4341;
  assign n4346 = n3364 & ~po129 ;
  assign n4347 = n3361 & po129 ;
  assign n4348 = ~n3361 & po129 ;
  assign n4349 = ~n3364 & ~po129 ;
  assign n4350 = ~n4348 & ~n4349;
  assign n4351 = ~n4346 & ~n4347;
  assign n4352 = n3354 & ~po129 ;
  assign n4353 = n3357 & po129 ;
  assign n4354 = ~n3357 & po129 ;
  assign n4355 = ~n3354 & ~po129 ;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = ~n4352 & ~n4353;
  assign n4358 = n3429 & ~po129 ;
  assign n4359 = n3426 & po129 ;
  assign n4360 = ~n3426 & po129 ;
  assign n4361 = ~n3429 & ~po129 ;
  assign n4362 = ~n4360 & ~n4361;
  assign n4363 = ~n4358 & ~n4359;
  assign n4364 = n3419 & ~po129 ;
  assign n4365 = n3422 & po129 ;
  assign n4366 = ~n3422 & po129 ;
  assign n4367 = ~n3419 & ~po129 ;
  assign n4368 = ~n4366 & ~n4367;
  assign n4369 = ~n4364 & ~n4365;
  assign n4370 = n3414 & ~po129 ;
  assign n4371 = n3411 & po129 ;
  assign n4372 = ~n3411 & po129 ;
  assign n4373 = ~n3414 & ~po129 ;
  assign n4374 = ~n4372 & ~n4373;
  assign n4375 = ~n4370 & ~n4371;
  assign n4376 = n3404 & ~po129 ;
  assign n4377 = n3407 & po129 ;
  assign n4378 = ~n3407 & po129 ;
  assign n4379 = ~n3404 & ~po129 ;
  assign n4380 = ~n4378 & ~n4379;
  assign n4381 = ~n4376 & ~n4377;
  assign n4382 = n3475 & ~po129 ;
  assign n4383 = n3478 & po129 ;
  assign n4384 = ~n3478 & po129 ;
  assign n4385 = ~n3475 & ~po129 ;
  assign n4386 = ~n4384 & ~n4385;
  assign n4387 = ~n4382 & ~n4383;
  assign n4388 = n3468 & ~po129 ;
  assign n4389 = n3471 & po129 ;
  assign n4390 = ~n3471 & po129 ;
  assign n4391 = ~n3468 & ~po129 ;
  assign n4392 = ~n4390 & ~n4391;
  assign n4393 = ~n4388 & ~n4389;
  assign n4394 = n3463 & ~po129 ;
  assign n4395 = n3460 & po129 ;
  assign n4396 = ~n3460 & po129 ;
  assign n4397 = ~n3463 & ~po129 ;
  assign n4398 = ~n4396 & ~n4397;
  assign n4399 = ~n4394 & ~n4395;
  assign n4400 = n3453 & ~po129 ;
  assign n4401 = n3456 & po129 ;
  assign n4402 = ~n3456 & po129 ;
  assign n4403 = ~n3453 & ~po129 ;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = ~n4400 & ~n4401;
  assign n4406 = n3528 & ~po129 ;
  assign n4407 = n3525 & po129 ;
  assign n4408 = ~n3525 & po129 ;
  assign n4409 = ~n3528 & ~po129 ;
  assign n4410 = ~n4408 & ~n4409;
  assign n4411 = ~n4406 & ~n4407;
  assign n4412 = n3518 & ~po129 ;
  assign n4413 = n3521 & po129 ;
  assign n4414 = ~n3521 & po129 ;
  assign n4415 = ~n3518 & ~po129 ;
  assign n4416 = ~n4414 & ~n4415;
  assign n4417 = ~n4412 & ~n4413;
  assign n4418 = n3513 & ~po129 ;
  assign n4419 = n3510 & po129 ;
  assign n4420 = ~n3510 & po129 ;
  assign n4421 = ~n3513 & ~po129 ;
  assign n4422 = ~n4420 & ~n4421;
  assign n4423 = ~n4418 & ~n4419;
  assign n4424 = n3503 & ~po129 ;
  assign n4425 = n3506 & po129 ;
  assign n4426 = ~n3506 & po129 ;
  assign n4427 = ~n3503 & ~po129 ;
  assign n4428 = ~n4426 & ~n4427;
  assign n4429 = ~n4424 & ~n4425;
  assign n4430 = n3569 & ~po129 ;
  assign n4431 = n3572 & po129 ;
  assign n4432 = ~n3572 & po129 ;
  assign n4433 = ~n3569 & ~po129 ;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = ~n4430 & ~n4431;
  assign n4436 = n3562 & ~po129 ;
  assign n4437 = n3565 & po129 ;
  assign n4438 = ~n3565 & po129 ;
  assign n4439 = ~n3562 & ~po129 ;
  assign n4440 = ~n4438 & ~n4439;
  assign n4441 = ~n4436 & ~n4437;
  assign n4442 = n3557 & ~po129 ;
  assign n4443 = n3554 & po129 ;
  assign n4444 = ~n3554 & po129 ;
  assign n4445 = ~n3557 & ~po129 ;
  assign n4446 = ~n4444 & ~n4445;
  assign n4447 = ~n4442 & ~n4443;
  assign n4448 = n3547 & ~po129 ;
  assign n4449 = n3550 & po129 ;
  assign n4450 = ~n3550 & po129 ;
  assign n4451 = ~n3547 & ~po129 ;
  assign n4452 = ~n4450 & ~n4451;
  assign n4453 = ~n4448 & ~n4449;
  assign n4454 = n3622 & ~po129 ;
  assign n4455 = n3619 & po129 ;
  assign n4456 = ~n3619 & po129 ;
  assign n4457 = ~n3622 & ~po129 ;
  assign n4458 = ~n4456 & ~n4457;
  assign n4459 = ~n4454 & ~n4455;
  assign n4460 = n3612 & ~po129 ;
  assign n4461 = n3615 & po129 ;
  assign n4462 = ~n3615 & po129 ;
  assign n4463 = ~n3612 & ~po129 ;
  assign n4464 = ~n4462 & ~n4463;
  assign n4465 = ~n4460 & ~n4461;
  assign n4466 = n3607 & ~po129 ;
  assign n4467 = n3604 & po129 ;
  assign n4468 = ~n3604 & po129 ;
  assign n4469 = ~n3607 & ~po129 ;
  assign n4470 = ~n4468 & ~n4469;
  assign n4471 = ~n4466 & ~n4467;
  assign n4472 = n3597 & ~po129 ;
  assign n4473 = n3600 & po129 ;
  assign n4474 = ~n3600 & po129 ;
  assign n4475 = ~n3597 & ~po129 ;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = ~n4472 & ~n4473;
  assign n4478 = n3668 & ~po129 ;
  assign n4479 = n3671 & po129 ;
  assign n4480 = ~n3671 & po129 ;
  assign n4481 = ~n3668 & ~po129 ;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = ~n4478 & ~n4479;
  assign n4484 = n3661 & ~po129 ;
  assign n4485 = n3664 & po129 ;
  assign n4486 = ~n3664 & po129 ;
  assign n4487 = ~n3661 & ~po129 ;
  assign n4488 = ~n4486 & ~n4487;
  assign n4489 = ~n4484 & ~n4485;
  assign n4490 = n3656 & ~po129 ;
  assign n4491 = n3653 & po129 ;
  assign n4492 = ~n3653 & po129 ;
  assign n4493 = ~n3656 & ~po129 ;
  assign n4494 = ~n4492 & ~n4493;
  assign n4495 = ~n4490 & ~n4491;
  assign n4496 = n3646 & ~po129 ;
  assign n4497 = n3649 & po129 ;
  assign n4498 = ~n3649 & po129 ;
  assign n4499 = ~n3646 & ~po129 ;
  assign n4500 = ~n4498 & ~n4499;
  assign n4501 = ~n4496 & ~n4497;
  assign n4502 = n3723 & ~po129 ;
  assign n4503 = n3720 & po129 ;
  assign n4504 = ~n3720 & po129 ;
  assign n4505 = ~n3723 & ~po129 ;
  assign n4506 = ~n4504 & ~n4505;
  assign n4507 = ~n4502 & ~n4503;
  assign n4508 = n3713 & ~po129 ;
  assign n4509 = n3716 & po129 ;
  assign n4510 = ~n3716 & po129 ;
  assign n4511 = ~n3713 & ~po129 ;
  assign n4512 = ~n4510 & ~n4511;
  assign n4513 = ~n4508 & ~n4509;
  assign n4514 = n3708 & ~po129 ;
  assign n4515 = n3705 & po129 ;
  assign n4516 = ~n3705 & po129 ;
  assign n4517 = ~n3708 & ~po129 ;
  assign n4518 = ~n4516 & ~n4517;
  assign n4519 = ~n4514 & ~n4515;
  assign n4520 = n3698 & ~po129 ;
  assign n4521 = n3701 & po129 ;
  assign n4522 = ~n3701 & po129 ;
  assign n4523 = ~n3698 & ~po129 ;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = ~n4520 & ~n4521;
  assign n4526 = n3770 & ~po129 ;
  assign n4527 = n3773 & po129 ;
  assign n4528 = ~n3773 & po129 ;
  assign n4529 = ~n3770 & ~po129 ;
  assign n4530 = ~n4528 & ~n4529;
  assign n4531 = ~n4526 & ~n4527;
  assign n4532 = n3751 & ~po129 ;
  assign n4533 = n3754 & po129 ;
  assign n4534 = ~n3754 & po129 ;
  assign n4535 = ~n3751 & ~po129 ;
  assign n4536 = ~n4534 & ~n4535;
  assign n4537 = ~n4532 & ~n4533;
  assign n4538 = n3744 & ~po129 ;
  assign n4539 = n3747 & po129 ;
  assign n4540 = ~n3747 & po129 ;
  assign n4541 = ~n3744 & ~po129 ;
  assign n4542 = ~n4540 & ~n4541;
  assign n4543 = ~n4538 & ~n4539;
  assign n4544 = ~n4696 & po129 ;
  assign n4545 = ~n4624 & ~po129 ;
  assign n4546 = n4624 & ~po129 ;
  assign n4547 = n4696 & po129 ;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = ~n4544 & ~n4545;
  assign n4550 = ~n4769 & n3791;
  assign n4551 = n4770 & ~n4550;
  assign n4552 = n4769 & n4770;
  assign n4553 = n703 | n704;
  assign n4554 = n712 | n713;
  assign n4555 = n718 | n719;
  assign n4556 = n728 | n729;
  assign n4557 = n734 | n735;
  assign n4558 = n752 | n753;
  assign n4559 = n758 | n759;
  assign n4560 = n776 | n777;
  assign n4561 = n782 | n783;
  assign n4562 = n799 | n800;
  assign n4563 = n820 | n821;
  assign n4564 = n830 | n831;
  assign n4565 = n835 | n836;
  assign n4566 = n841 | n842;
  assign n4567 = n857 | n858;
  assign n4568 = n860 | n861;
  assign n4569 = n864 | n865;
  assign n4570 = n890 | n891;
  assign n4571 = n906 | n907;
  assign n4572 = n909 | n910;
  assign n4573 = n915 | n916;
  assign n4574 = n921 | ~n922;
  assign n4575 = n940 | n936 | n939;
  assign n4576 = n945 | n946;
  assign n4577 = n951 | n952;
  assign n4578 = n958 | n959;
  assign n4579 = n964 | n965;
  assign n4580 = n970 | ~n971;
  assign n4581 = n972 | n973;
  assign n4582 = n990 | n991;
  assign n4583 = n1000 | n1001;
  assign n4584 = n1016 | n1017;
  assign n4585 = n1019 | n1020;
  assign n4586 = n1025 | n1026;
  assign n4587 = n1036 | n1037;
  assign n4588 = n1045 | n1046;
  assign n4589 = n1069 | n1070;
  assign n4590 = n1072 | n1073;
  assign n4591 = n1076 | n1077;
  assign n4592 = n1093 | n1094;
  assign n4593 = n1117 | n1118;
  assign n4594 = n1120 | n1121;
  assign n4595 = n1124 | n1125;
  assign n4596 = n1135 | n1136;
  assign n4597 = n1140 | n1141;
  assign n4598 = n1146 | n1147;
  assign n4599 = n1170 | n1171;
  assign n4600 = n1173 | n1174;
  assign n4601 = n1177 | n1178;
  assign n4602 = n1194 | n1195;
  assign n4603 = n1218 | n1219;
  assign n4604 = n1221 | n1222;
  assign n4605 = n1225 | n1226;
  assign n4606 = n1236 | n1237;
  assign n4607 = n1241 | n1242;
  assign n4608 = n1247 | n1248;
  assign n4609 = n1271 | n1272;
  assign n4610 = n1274 | n1275;
  assign n4611 = n1278 | n1279;
  assign n4612 = n1295 | n1296;
  assign n4613 = n1319 | n1320;
  assign n4614 = n1322 | n1323;
  assign n4615 = n1326 | n1327;
  assign n4616 = n1337 | n1338;
  assign n4617 = n1342 | n1343;
  assign n4618 = n1348 | n1349;
  assign n4619 = n1372 | n1373;
  assign n4620 = n1375 | n1376;
  assign n4621 = n1379 | n1380;
  assign n4622 = n1396 | n1397;
  assign n4623 = n1408 | n1409;
  assign n4624 = n1421 | n1422;
  assign n4625 = n1488 | n1489;
  assign n4626 = n1497 | n1498;
  assign n4627 = n1503 | n1504;
  assign n4628 = n1513 | n1514;
  assign n4629 = n1519 | n1520;
  assign n4630 = n1537 | n1538;
  assign n4631 = n1543 | n1544;
  assign n4632 = n1561 | n1562;
  assign n4633 = n1567 | n1568;
  assign n4634 = n1584 | n1585;
  assign n4635 = n1605 | n1606;
  assign n4636 = n1615 | n1616;
  assign n4637 = n1620 | n1621;
  assign n4638 = n1626 | n1627;
  assign n4639 = n1642 | n1643;
  assign n4640 = n1645 | n1646;
  assign n4641 = n1649 | n1650;
  assign n4642 = n1675 | n1676;
  assign n4643 = n1691 | n1692;
  assign n4644 = n1694 | n1695;
  assign n4645 = n1700 | n1701;
  assign n4646 = n1706 | ~n1707;
  assign n4647 = n1725 | n1721 | n1724;
  assign n4648 = n1730 | n1731;
  assign n4649 = n1736 | n1737;
  assign n4650 = n1743 | n1744;
  assign n4651 = n1749 | n1750;
  assign n4652 = n1755 | ~n1756;
  assign n4653 = n1757 | n1758;
  assign n4654 = n1775 | n1776;
  assign n4655 = n1785 | n1786;
  assign n4656 = n1801 | n1802;
  assign n4657 = n1804 | n1805;
  assign n4658 = n1810 | n1811;
  assign n4659 = n1821 | n1822;
  assign n4660 = n1830 | n1831;
  assign n4661 = n1854 | n1855;
  assign n4662 = n1857 | n1858;
  assign n4663 = n1861 | n1862;
  assign n4664 = n1878 | n1879;
  assign n4665 = n1902 | n1903;
  assign n4666 = n1905 | n1906;
  assign n4667 = n1909 | n1910;
  assign n4668 = n1920 | n1921;
  assign n4669 = n1925 | n1926;
  assign n4670 = n1931 | n1932;
  assign n4671 = n1955 | n1956;
  assign n4672 = n1958 | n1959;
  assign n4673 = n1962 | n1963;
  assign n4674 = n1979 | n1980;
  assign n4675 = n2003 | n2004;
  assign n4676 = n2006 | n2007;
  assign n4677 = n2010 | n2011;
  assign n4678 = n2021 | n2022;
  assign n4679 = n2026 | n2027;
  assign n4680 = n2032 | n2033;
  assign n4681 = n2056 | n2057;
  assign n4682 = n2059 | n2060;
  assign n4683 = n2063 | n2064;
  assign n4684 = n2080 | n2081;
  assign n4685 = n2104 | n2105;
  assign n4686 = n2107 | n2108;
  assign n4687 = n2111 | n2112;
  assign n4688 = n2122 | n2123;
  assign n4689 = n2127 | n2128;
  assign n4690 = n2133 | n2134;
  assign n4691 = n2157 | n2158;
  assign n4692 = n2160 | n2161;
  assign n4693 = n2164 | n2165;
  assign n4694 = n2181 | n2182;
  assign n4695 = n2193 | n2194;
  assign n4696 = n2206 | n2207;
  assign n4697 = n2353 | n2354;
  assign n4698 = n2360 | ~n2361;
  assign n4699 = n2364 | ~n2365;
  assign n4700 = n2375 | ~n2376;
  assign n4701 = n2386 | ~n2387;
  assign n4702 = n2400 | ~n2401;
  assign n4703 = n2433 | ~n2434;
  assign n4704 = n2439 | n2440;
  assign n4705 = n2469 | n2470;
  assign n4706 = n2489 | ~n2490;
  assign n4707 = n2494 | n2495;
  assign n4708 = n2525 | n2526;
  assign n4709 = n2545 | ~n2546;
  assign n4710 = n2550 | n2551;
  assign n4711 = n2579 | n2580;
  assign n4712 = n2657 | n2658;
  assign n4713 = n2661 | n2662;
  assign n4714 = n2668 | n2669;
  assign n4715 = n2676 | n2677;
  assign n4716 = n2681 | n2682;
  assign n4717 = n2686 | n2687;
  assign n4718 = n2695 | n2696;
  assign n4719 = n2705 | n2701 | n2704;
  assign n4720 = n2739 | n2740;
  assign n4721 = n2775 | n2776;
  assign n4722 = n2785 | n2786;
  assign n4723 = n2799 | n2800;
  assign n4724 = n2805 | n2806;
  assign n4725 = n2810 | n2811;
  assign n4726 = n2878 | n2875 | n2877;
  assign n4727 = n2887 | n2888;
  assign n4728 = n2891 | n2892;
  assign n4729 = n2901 | n2902;
  assign n4730 = n2906 | n2907;
  assign n4731 = n2941 | n2942;
  assign n4732 = n2980 | n2977 | n2979;
  assign n4733 = n2989 | n2990;
  assign n4734 = n3003 | n3004;
  assign n4735 = n3009 | n3010;
  assign n4736 = n3014 | n3015;
  assign n4737 = n3049 | n3050;
  assign n4738 = n3054 | n3055;
  assign n4739 = n3060 | n3061;
  assign n4740 = n3109 | n3110;
  assign n4741 = n3113 | n3114;
  assign n4742 = n3154 | n3155;
  assign n4743 = n3203 | n3204;
  assign n4744 = n3207 | n3208;
  assign n4745 = n3242 | n3243;
  assign n4746 = n3247 | n3248;
  assign n4747 = n3253 | n3254;
  assign n4748 = n3302 | n3303;
  assign n4749 = n3306 | n3307;
  assign n4750 = n3347 | n3348;
  assign n4751 = n3396 | n3397;
  assign n4752 = n3400 | n3401;
  assign n4753 = n3435 | n3436;
  assign n4754 = n3440 | n3441;
  assign n4755 = n3446 | n3447;
  assign n4756 = n3495 | n3496;
  assign n4757 = n3499 | n3500;
  assign n4758 = n3540 | n3541;
  assign n4759 = n3589 | n3590;
  assign n4760 = n3593 | n3594;
  assign n4761 = n3628 | n3629;
  assign n4762 = n3633 | n3634;
  assign n4763 = n3639 | n3640;
  assign n4764 = n3679 | n3680;
  assign n4765 = n3690 | n3691;
  assign n4766 = n3694 | n3695;
  assign n4767 = n3731 | n3732;
  assign n4768 = n3737 | n3738;
  assign n4769 = n3761 | n3758 | n3760;
  assign n4770 = n3766 | n3763 | n3765;
  assign n4771 = n3777 | n3778;
  assign po129  = n3792 | n3793;
  assign n4773 = n3801 | ~n3802;
  assign n4774 = n3807 | ~n3808;
  assign n4775 = n3813 | ~n3814;
  assign n4776 = n3828 | ~n3829;
  assign n4777 = n3834 | ~n3835;
  assign n4778 = n3840 | ~n3841;
  assign n4779 = n3846 | ~n3847;
  assign n4780 = n3852 | ~n3853;
  assign n4781 = n3858 | ~n3859;
  assign n4782 = n3864 | ~n3865;
  assign n4783 = n3870 | ~n3871;
  assign n4784 = n3876 | ~n3877;
  assign n4785 = n3882 | ~n3883;
  assign n4786 = n3888 | ~n3889;
  assign n4787 = n3894 | ~n3895;
  assign n4788 = n3900 | ~n3901;
  assign n4789 = n3906 | ~n3907;
  assign n4790 = n3912 | ~n3913;
  assign n4791 = n3918 | ~n3919;
  assign n4792 = n3924 | ~n3925;
  assign n4793 = n3930 | ~n3931;
  assign n4794 = n3936 | ~n3937;
  assign n4795 = n3942 | ~n3943;
  assign n4796 = n3948 | ~n3949;
  assign n4797 = n3954 | ~n3955;
  assign n4798 = n3960 | ~n3961;
  assign n4799 = n3966 | ~n3967;
  assign n4800 = n3972 | ~n3973;
  assign n4801 = n3978 | ~n3979;
  assign n4802 = n3984 | ~n3985;
  assign n4803 = n3990 | ~n3991;
  assign n4804 = n3996 | ~n3997;
  assign n4805 = n4002 | ~n4003;
  assign n4806 = n4008 | ~n4009;
  assign n4807 = n4014 | ~n4015;
  assign n4808 = n4020 | ~n4021;
  assign n4809 = n4026 | ~n4027;
  assign n4810 = n4032 | ~n4033;
  assign n4811 = n4038 | ~n4039;
  assign n4812 = n4044 | ~n4045;
  assign n4813 = n4050 | ~n4051;
  assign n4814 = n4056 | ~n4057;
  assign n4815 = n4062 | ~n4063;
  assign n4816 = n4068 | ~n4069;
  assign n4817 = n4074 | ~n4075;
  assign n4818 = n4080 | ~n4081;
  assign n4819 = n4086 | ~n4087;
  assign n4820 = n4092 | ~n4093;
  assign n4821 = n4098 | ~n4099;
  assign n4822 = n4104 | ~n4105;
  assign n4823 = n4110 | ~n4111;
  assign n4824 = n4116 | ~n4117;
  assign n4825 = n4122 | ~n4123;
  assign n4826 = n4128 | ~n4129;
  assign n4827 = n4134 | ~n4135;
  assign n4828 = n4140 | ~n4141;
  assign n4829 = n4146 | ~n4147;
  assign n4830 = n4152 | ~n4153;
  assign n4831 = n4158 | ~n4159;
  assign n4832 = n4164 | ~n4165;
  assign n4833 = n4170 | ~n4171;
  assign n4834 = n4176 | ~n4177;
  assign n4835 = n4182 | ~n4183;
  assign n4836 = n4188 | ~n4189;
  assign n4837 = n4194 | ~n4195;
  assign n4838 = n4200 | ~n4201;
  assign n4839 = n4206 | ~n4207;
  assign n4840 = n4212 | ~n4213;
  assign n4841 = n4218 | ~n4219;
  assign n4842 = n4224 | ~n4225;
  assign n4843 = n4230 | ~n4231;
  assign n4844 = n4236 | ~n4237;
  assign n4845 = n4242 | ~n4243;
  assign n4846 = n4248 | ~n4249;
  assign n4847 = n4254 | ~n4255;
  assign n4848 = n4260 | ~n4261;
  assign n4849 = n4266 | ~n4267;
  assign n4850 = n4272 | ~n4273;
  assign n4851 = n4278 | ~n4279;
  assign n4852 = n4284 | ~n4285;
  assign n4853 = n4290 | ~n4291;
  assign n4854 = n4296 | ~n4297;
  assign n4855 = n4302 | ~n4303;
  assign n4856 = n4308 | ~n4309;
  assign n4857 = n4314 | ~n4315;
  assign n4858 = n4320 | ~n4321;
  assign n4859 = n4326 | ~n4327;
  assign n4860 = n4332 | ~n4333;
  assign n4861 = n4338 | ~n4339;
  assign n4862 = n4344 | ~n4345;
  assign n4863 = n4350 | ~n4351;
  assign n4864 = n4356 | ~n4357;
  assign n4865 = n4362 | ~n4363;
  assign n4866 = n4368 | ~n4369;
  assign n4867 = n4374 | ~n4375;
  assign n4868 = n4380 | ~n4381;
  assign n4869 = n4386 | ~n4387;
  assign n4870 = n4392 | ~n4393;
  assign n4871 = n4398 | ~n4399;
  assign n4872 = n4404 | ~n4405;
  assign n4873 = n4410 | ~n4411;
  assign n4874 = n4416 | ~n4417;
  assign n4875 = n4422 | ~n4423;
  assign n4876 = n4428 | ~n4429;
  assign n4877 = n4434 | ~n4435;
  assign n4878 = n4440 | ~n4441;
  assign n4879 = n4446 | ~n4447;
  assign n4880 = n4452 | ~n4453;
  assign n4881 = n4458 | ~n4459;
  assign n4882 = n4464 | ~n4465;
  assign n4883 = n4470 | ~n4471;
  assign n4884 = n4476 | ~n4477;
  assign n4885 = n4482 | ~n4483;
  assign n4886 = n4488 | ~n4489;
  assign n4887 = n4494 | ~n4495;
  assign n4888 = n4500 | ~n4501;
  assign n4889 = n4506 | ~n4507;
  assign n4890 = n4512 | ~n4513;
  assign n4891 = n4518 | ~n4519;
  assign n4892 = n4524 | ~n4525;
  assign n4893 = n4530 | ~n4531;
  assign n4894 = n4536 | ~n4537;
  assign n4895 = n4542 | ~n4543;
  assign n4896 = n4548 | ~n4549;
  assign po127  = n4551 | n4552;
  assign po0  = ~n3796;
  assign po1  = ~n4773;
  assign po2  = ~n4774;
  assign po3  = ~n4775;
  assign po4  = ~n3817;
  assign po5  = ~n3820;
  assign po6  = ~n3823;
  assign po7  = ~n4776;
  assign po8  = ~n4777;
  assign po9  = ~n4778;
  assign po10  = ~n4779;
  assign po11  = ~n4780;
  assign po12  = ~n4781;
  assign po13  = ~n4782;
  assign po14  = ~n4783;
  assign po15  = ~n4784;
  assign po16  = ~n4785;
  assign po17  = ~n4786;
  assign po18  = ~n4787;
  assign po19  = ~n4788;
  assign po20  = ~n4789;
  assign po21  = ~n4790;
  assign po22  = ~n4791;
  assign po23  = ~n4792;
  assign po24  = ~n4793;
  assign po25  = ~n4794;
  assign po26  = ~n4795;
  assign po27  = ~n4796;
  assign po28  = ~n4797;
  assign po29  = ~n4798;
  assign po30  = ~n4799;
  assign po31  = ~n4800;
  assign po32  = ~n4801;
  assign po33  = ~n4802;
  assign po34  = ~n4803;
  assign po35  = ~n4804;
  assign po36  = ~n4805;
  assign po37  = ~n4806;
  assign po38  = ~n4807;
  assign po39  = ~n4808;
  assign po40  = ~n4809;
  assign po41  = ~n4810;
  assign po42  = ~n4811;
  assign po43  = ~n4812;
  assign po44  = ~n4813;
  assign po45  = ~n4814;
  assign po46  = ~n4815;
  assign po47  = ~n4816;
  assign po48  = ~n4817;
  assign po49  = ~n4818;
  assign po50  = ~n4819;
  assign po51  = ~n4820;
  assign po52  = ~n4821;
  assign po53  = ~n4822;
  assign po54  = ~n4823;
  assign po55  = ~n4824;
  assign po56  = ~n4825;
  assign po57  = ~n4826;
  assign po58  = ~n4827;
  assign po59  = ~n4828;
  assign po60  = ~n4829;
  assign po61  = ~n4830;
  assign po62  = ~n4831;
  assign po63  = ~n4832;
  assign po64  = ~n4833;
  assign po65  = ~n4834;
  assign po66  = ~n4835;
  assign po67  = ~n4836;
  assign po68  = ~n4837;
  assign po69  = ~n4838;
  assign po70  = ~n4839;
  assign po71  = ~n4840;
  assign po72  = ~n4841;
  assign po73  = ~n4842;
  assign po74  = ~n4843;
  assign po75  = ~n4844;
  assign po76  = ~n4845;
  assign po77  = ~n4846;
  assign po78  = ~n4847;
  assign po79  = ~n4848;
  assign po80  = ~n4849;
  assign po81  = ~n4850;
  assign po82  = ~n4851;
  assign po83  = ~n4852;
  assign po84  = ~n4853;
  assign po85  = ~n4854;
  assign po86  = ~n4855;
  assign po87  = ~n4856;
  assign po88  = ~n4857;
  assign po89  = ~n4858;
  assign po90  = ~n4859;
  assign po91  = ~n4860;
  assign po92  = ~n4861;
  assign po93  = ~n4862;
  assign po94  = ~n4863;
  assign po95  = ~n4864;
  assign po96  = ~n4865;
  assign po97  = ~n4866;
  assign po98  = ~n4867;
  assign po99  = ~n4868;
  assign po100  = ~n4869;
  assign po101  = ~n4870;
  assign po102  = ~n4871;
  assign po103  = ~n4872;
  assign po104  = ~n4873;
  assign po105  = ~n4874;
  assign po106  = ~n4875;
  assign po107  = ~n4876;
  assign po108  = ~n4877;
  assign po109  = ~n4878;
  assign po110  = ~n4879;
  assign po111  = ~n4880;
  assign po112  = ~n4881;
  assign po113  = ~n4882;
  assign po114  = ~n4883;
  assign po115  = ~n4884;
  assign po116  = ~n4885;
  assign po117  = ~n4886;
  assign po118  = ~n4887;
  assign po119  = ~n4888;
  assign po120  = ~n4889;
  assign po121  = ~n4890;
  assign po122  = ~n4891;
  assign po123  = ~n4892;
  assign po124  = ~n4893;
  assign po125  = ~n4894;
  assign po126  = ~n4895;
  assign po128  = ~n4896;
endmodule
